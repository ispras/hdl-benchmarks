module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
 n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
 n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
 n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
 n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
 n271 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 ;
output n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
 n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
 n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
 n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
 n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
 n271 ;
wire n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , 
 n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , 
 n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , 
 n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , 
 n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , 
 n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , 
 n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , 
 n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , 
 n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , 
 n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , 
 n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , 
 n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , 
 n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , 
 n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , 
 n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , 
 n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , 
 n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , 
 n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , 
 n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , 
 n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , 
 n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , 
 n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , 
 n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , 
 n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , 
 n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , 
 n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , 
 n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , 
 n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , 
 n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , 
 n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , 
 n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , 
 n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , 
 n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , 
 n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , 
 n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , 
 n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , 
 n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , 
 n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , 
 n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , 
 n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , 
 n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , 
 n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , 
 n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , 
 n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , 
 n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , 
 n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , 
 n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , 
 n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , 
 n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , 
 n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , 
 n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , 
 n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , 
 n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , 
 n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , 
 n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , 
 n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , 
 n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , 
 n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , 
 n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , 
 n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , 
 n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , 
 n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , 
 n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , 
 n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , 
 n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , 
 n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , 
 n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , 
 n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , 
 n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , 
 n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , 
 n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , 
 n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , 
 n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , 
 n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , 
 n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , 
 n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , 
 n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , 
 n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , 
 n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , 
 n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , 
 n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , 
 n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , 
 n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , 
 n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , 
 n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , 
 n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , 
 n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , 
 n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , 
 n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , 
 n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , 
 n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , 
 n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , 
 n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , 
 n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , 
 n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , 
 n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , 
 n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , 
 n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , 
 n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , 
 n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , 
 n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , 
 n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , 
 n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , 
 n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , 
 n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , 
 n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , 
 n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , 
 n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , 
 n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , 
 n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , 
 n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , 
 n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , 
 n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , 
 n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , 
 n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , 
 n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , 
 n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , 
 n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , 
 n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , 
 n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , 
 n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , 
 n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , 
 n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , 
 n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , 
 n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , 
 n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , 
 n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , 
 n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , 
 n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , 
 n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , 
 n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , 
 n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , 
 n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , 
 n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , 
 n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , 
 n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , 
 n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , 
 n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , 
 n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , 
 n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , 
 n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , 
 n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , 
 n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , 
 n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , 
 n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , 
 n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , 
 n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , 
 n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , 
 n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , 
 n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , 
 n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , 
 n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , 
 n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , 
 n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , 
 n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , 
 n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , 
 n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , 
 n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , 
 n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , 
 n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , 
 n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , 
 n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , 
 n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , 
 n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , 
 n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , 
 n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , 
 n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , 
 n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , 
 n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , 
 n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , 
 n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , 
 n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , 
 n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , 
 n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , 
 n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , 
 n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , 
 n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , 
 n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , 
 n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , 
 n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , 
 n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , 
 n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , 
 n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , 
 n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , 
 n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , 
 n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , 
 n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , 
 n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , 
 n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , 
 n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , 
 n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , 
 n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , 
 n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , 
 n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , 
 n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , 
 n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , 
 n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , 
 n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , 
 n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , 
 n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , 
 n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , 
 n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , 
 n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , 
 n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , 
 n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , 
 n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , 
 n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , 
 n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , 
 n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , 
 n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , 
 n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , 
 n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , 
 n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , 
 n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , 
 n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , 
 n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , 
 n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , 
 n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , 
 n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , 
 n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , 
 n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , 
 n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , 
 n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , 
 n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , 
 n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , 
 n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , 
 n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , 
 n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , 
 n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , 
 n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , 
 n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , 
 n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , 
 n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , 
 n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , 
 n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , 
 n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , 
 n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , 
 n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , 
 n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , 
 n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , 
 n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , 
 n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , 
 n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , 
 n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , 
 n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , 
 n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , 
 n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , 
 n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , 
 n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , 
 n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , 
 n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , 
 n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , 
 n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , 
 n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , 
 n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , 
 n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , 
 n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , 
 n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , 
 n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , 
 n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , 
 n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , 
 n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , 
 n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , 
 n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , 
 n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , 
 n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , 
 n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , 
 n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , 
 n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , 
 n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , 
 n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , 
 n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , 
 n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , 
 n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , 
 n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , 
 n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , 
 n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , 
 n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , 
 n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , 
 n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , 
 n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , 
 n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , 
 n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , 
 n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , 
 n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , 
 n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , 
 n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , 
 n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , 
 n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , 
 n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , 
 n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , 
 n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , 
 n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , 
 n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , 
 n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , 
 n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , 
 n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , 
 n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , 
 n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , 
 n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , 
 n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , 
 n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , 
 n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , 
 n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , 
 n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , 
 n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , 
 n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , 
 n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , 
 n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , 
 n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , 
 n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , 
 n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , 
 n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , 
 n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , 
 n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , 
 n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , 
 n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , 
 n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , 
 n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , 
 n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , 
 n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , 
 n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , 
 n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , 
 n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , 
 n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , 
 n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , 
 n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , 
 n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , 
 n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , 
 n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , 
 n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , 
 n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , 
 n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , 
 n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , 
 n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , 
 n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , 
 n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , 
 n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , 
 n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , 
 n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , 
 n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , 
 n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , 
 n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , 
 n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , 
 n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , 
 n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , 
 n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , 
 n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , 
 n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , 
 n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , 
 n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , 
 n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , 
 n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , 
 n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , 
 n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , 
 n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , 
 n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , 
 n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , 
 n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , 
 n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , 
 n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , 
 n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , 
 n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , 
 n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , 
 n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , 
 n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , 
 n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , 
 n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , 
 n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , 
 n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , 
 n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , 
 n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , 
 n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , 
 n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , 
 n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , 
 n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , 
 n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , 
 n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , 
 n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , 
 n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , 
 n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , 
 n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , 
 n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , 
 n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , 
 n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , 
 n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , 
 n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , 
 n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , 
 n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , 
 n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , 
 n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , 
 n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , 
 n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , 
 n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , 
 n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , 
 n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , 
 n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , 
 n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , 
 n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , 
 n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , 
 n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , 
 n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , 
 n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , 
 n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , 
 n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , 
 n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , 
 n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , 
 n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , 
 n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , 
 n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , 
 n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , 
 n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , 
 n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , 
 n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , 
 n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , 
 n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , 
 n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , 
 n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , 
 n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , 
 n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , 
 n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , 
 n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , 
 n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , 
 n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , 
 n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , 
 n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , 
 n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , 
 n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , 
 n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , 
 n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , 
 n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , 
 n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , 
 n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , 
 n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , 
 n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , 
 n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , 
 n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , 
 n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , 
 n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , 
 n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , 
 n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , 
 n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , 
 n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , 
 n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , 
 n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , 
 n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , 
 n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , 
 n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , 
 n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , 
 n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , 
 n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , 
 n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , 
 n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , 
 n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , 
 n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , 
 n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , 
 n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , 
 n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , 
 n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , 
 n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , 
 n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , 
 n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , 
 n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , 
 n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , 
 n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , 
 n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , 
 n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , 
 n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , 
 n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , 
 n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , 
 n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , 
 n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , 
 n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , 
 n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , 
 n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , 
 n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , 
 n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , 
 n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , 
 n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , 
 n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , 
 n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , 
 n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , 
 n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , 
 n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , 
 n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , 
 n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , 
 n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , 
 n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , 
 n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , 
 n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , 
 n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , 
 n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , 
 n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , 
 n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , 
 n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , 
 n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , 
 n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , 
 n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , 
 n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , 
 n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , 
 n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , 
 n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , 
 n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , 
 n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , 
 n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , 
 n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , 
 n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , 
 n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , 
 n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , 
 n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , 
 n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , 
 n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , 
 n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , 
 n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , 
 n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , 
 n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , 
 n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , 
 n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , 
 n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , 
 n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , 
 n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , 
 n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , 
 n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , 
 n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , 
 n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , 
 n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , 
 n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , 
 n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , 
 n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , 
 n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , 
 n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , 
 n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , 
 n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , 
 n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , 
 n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , 
 n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , 
 n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , 
 n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , 
 n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , 
 n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , 
 n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , 
 n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , 
 n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , 
 n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , 
 n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , 
 n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , 
 n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , 
 n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , 
 n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , 
 n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , 
 n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , 
 n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , 
 n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , 
 n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , 
 n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , 
 n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , 
 n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , 
 n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , 
 n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , 
 n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , 
 n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , 
 n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , 
 n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , 
 n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , 
 n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , 
 n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , 
 n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , 
 n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , 
 n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , 
 n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , 
 n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , 
 n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , 
 n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , 
 n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , 
 n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , 
 n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , 
 n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , 
 n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , 
 n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , 
 n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , 
 n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , 
 n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , 
 n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , 
 n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , 
 n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , 
 n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , 
 n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , 
 n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , 
 n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , 
 n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , 
 n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , 
 n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , 
 n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , 
 n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , 
 n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , 
 n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , 
 n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , 
 n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , 
 n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , 
 n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , 
 n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , 
 n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , 
 n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , 
 n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , 
 n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , 
 n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , 
 n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , 
 n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , 
 n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , 
 n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , 
 n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , 
 n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , 
 n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , 
 n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , 
 n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , 
 n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , 
 n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , 
 n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , 
 n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , 
 n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , 
 n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , 
 n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , 
 n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , 
 n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , 
 n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , 
 n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , 
 n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , 
 n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , 
 n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , 
 n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , 
 n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , 
 n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , 
 n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , 
 n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , 
 n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , 
 n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , 
 n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , 
 n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , 
 n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , 
 n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , 
 n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , 
 n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , 
 n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , 
 n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , 
 n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , 
 n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , 
 n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , 
 n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , 
 n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , 
 n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , 
 n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , 
 n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , 
 n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , 
 n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , 
 n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , 
 n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , 
 n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , 
 n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , 
 n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , 
 n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , 
 n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , 
 n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , 
 n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , 
 n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , 
 n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , 
 n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , 
 n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , 
 n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , 
 n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , 
 n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , 
 n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , 
 n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , 
 n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , 
 n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , 
 n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , 
 n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , 
 n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , 
 n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , 
 n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , 
 n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , 
 n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , 
 n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , 
 n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , 
 n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , 
 n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , 
 n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , 
 n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , 
 n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , 
 n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , 
 n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , 
 n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , 
 n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , 
 n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , 
 n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , 
 n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , 
 n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , 
 n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , 
 n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , 
 n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , 
 n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , 
 n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , 
 n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , 
 n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , 
 n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , 
 n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , 
 n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , 
 n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , 
 n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , 
 n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , 
 n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , 
 n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , 
 n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , 
 n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , 
 n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , 
 n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , 
 n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , 
 n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , 
 n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , 
 n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , 
 n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , 
 n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , 
 n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , 
 n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , 
 n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , 
 n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , 
 n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , 
 n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , 
 n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , 
 n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , 
 n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , 
 n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , 
 n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , 
 n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , 
 n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , 
 n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , 
 n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , 
 n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , 
 n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , 
 n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , 
 n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , 
 n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , 
 n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , 
 n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , 
 n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , 
 n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , 
 n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , 
 n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , 
 n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , 
 n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , 
 n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , 
 n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , 
 n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , 
 n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , 
 n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , 
 n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , 
 n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , 
 n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , 
 n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , 
 n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , 
 n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , 
 n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , 
 n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , 
 n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , 
 n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , 
 n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , 
 n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , 
 n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , 
 n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , 
 n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , 
 n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , 
 n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , 
 n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , 
 n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , 
 n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , 
 n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , 
 n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , 
 n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , 
 n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , 
 n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , 
 n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , 
 n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , 
 n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , 
 n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , 
 n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , 
 n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , 
 n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , 
 n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , 
 n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , 
 n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , 
 n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , 
 n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , 
 n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , 
 n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , 
 n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , 
 n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , 
 n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , 
 n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , 
 n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , 
 n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , 
 n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , 
 n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , 
 n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , 
 n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , 
 n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , 
 n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , 
 n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , 
 n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , 
 n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , 
 n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , 
 n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , 
 n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , 
 n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , 
 n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , 
 n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , 
 n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , 
 n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , 
 n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , 
 n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , 
 n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , 
 n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , 
 n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , 
 n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , 
 n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , 
 n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , 
 n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , 
 n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , 
 n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , 
 n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , 
 n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , 
 n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , 
 n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , 
 n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , 
 n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , 
 n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , 
 n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , 
 n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , 
 n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , 
 n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , 
 n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , 
 n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , 
 n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , 
 n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , 
 n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , 
 n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , 
 n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , 
 n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , 
 n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , 
 n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , 
 n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , 
 n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , 
 n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , 
 n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , 
 n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , 
 n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , 
 n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , 
 n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , 
 n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , 
 n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , 
 n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , 
 n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , 
 n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , 
 n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , 
 n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , 
 n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , 
 n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , 
 n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , 
 n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , 
 n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , 
 n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , 
 n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , 
 n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , 
 n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , 
 n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , 
 n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , 
 n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , 
 n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , 
 n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , 
 n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , 
 n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , 
 n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , 
 n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , 
 n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , 
 n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , 
 n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , 
 n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , 
 n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , 
 n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , 
 n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , 
 n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , 
 n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , 
 n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , 
 n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , 
 n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , 
 n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , 
 n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , 
 n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , 
 n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , 
 n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , 
 n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , 
 n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , 
 n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , 
 n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , 
 n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , 
 n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , 
 n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , 
 n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , 
 n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , 
 n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , 
 n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , 
 n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , 
 n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , 
 n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , 
 n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , 
 n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , 
 n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , 
 n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , 
 n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , 
 n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , 
 n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , 
 n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , 
 n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , 
 n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , 
 n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , 
 n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , 
 n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , 
 n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , 
 n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , 
 n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , 
 n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , 
 n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , 
 n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , 
 n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , 
 n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , 
 n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , 
 n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , 
 n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , 
 n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , 
 n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , 
 n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , 
 n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , 
 n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , 
 n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , 
 n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , 
 n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , 
 n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , 
 n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , 
 n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , 
 n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , 
 n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , 
 n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , 
 n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , 
 n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , 
 n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , 
 n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , 
 n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , 
 n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , 
 n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , 
 n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , 
 n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , 
 n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , 
 n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , 
 n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , 
 n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , 
 n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , 
 n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , 
 n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , 
 n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , 
 n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , 
 n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , 
 n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , 
 n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , 
 n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , 
 n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , 
 n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , 
 n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , 
 n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , 
 n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , 
 n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , 
 n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , 
 n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , 
 n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , 
 n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , 
 n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , 
 n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , 
 n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , 
 n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , 
 n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , 
 n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , 
 n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , 
 n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , 
 n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , 
 n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , 
 n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , 
 n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , 
 n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , 
 n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , 
 n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , 
 n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , 
 n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , 
 n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , 
 n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , 
 n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , 
 n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , 
 n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , 
 n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , 
 n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , 
 n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , 
 n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , 
 n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , 
 n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , 
 n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , 
 n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , 
 n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , 
 n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , 
 n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , 
 n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , 
 n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , 
 n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , 
 n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , 
 n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , 
 n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , 
 n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , 
 n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , 
 n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , 
 n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , 
 n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , 
 n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , 
 n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , 
 n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , 
 n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , 
 n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , 
 n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , 
 n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , 
 n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , 
 n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , 
 n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , 
 n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , 
 n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , 
 n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , 
 n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , 
 n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , 
 n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , 
 n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , 
 n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , 
 n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , 
 n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , 
 n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , 
 n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , 
 n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , 
 n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , 
 n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , 
 n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , 
 n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , 
 n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , 
 n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , 
 n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , 
 n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , 
 n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , 
 n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , 
 n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , 
 n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , 
 n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , 
 n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , 
 n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , 
 n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , 
 n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , 
 n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , 
 n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , 
 n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , 
 n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , 
 n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , 
 n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , 
 n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , 
 n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , 
 n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , 
 n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , 
 n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , 
 n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , 
 n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , 
 n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , 
 n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , 
 n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , 
 n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , 
 n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , 
 n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , 
 n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , 
 n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , 
 n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , 
 n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , 
 n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , 
 n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , 
 n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , 
 n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , 
 n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , 
 n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , 
 n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , 
 n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , 
 n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , 
 n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , 
 n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , 
 n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , 
 n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , 
 n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , 
 n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , 
 n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , 
 n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , 
 n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , 
 n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , 
 n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , 
 n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , 
 n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , 
 n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , 
 n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , 
 n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , 
 n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , 
 n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , 
 n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , 
 n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , 
 n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , 
 n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , 
 n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , 
 n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , 
 n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , 
 n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , 
 n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , 
 n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , 
 n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , 
 n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , 
 n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , 
 n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , 
 n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , 
 n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , 
 n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , 
 n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , 
 n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , 
 n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , 
 n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , 
 n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , 
 n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , 
 n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , 
 n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , 
 n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , 
 n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , 
 n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , 
 n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , 
 n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , 
 n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , 
 n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , 
 n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , 
 n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , 
 n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , 
 n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , 
 n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , 
 n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , 
 n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , 
 n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , 
 n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , 
 n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , 
 n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , 
 n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , 
 n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , 
 n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , 
 n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , 
 n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , 
 n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , 
 n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , 
 n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , 
 n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , 
 n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , 
 n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , 
 n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , 
 n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , 
 n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , 
 n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , 
 n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , 
 n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , 
 n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , 
 n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , 
 n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , 
 n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , 
 n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , 
 n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , 
 n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , 
 n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , 
 n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , 
 n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , 
 n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , 
 n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , 
 n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , 
 n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , 
 n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , 
 n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , 
 n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , 
 n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , 
 n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , 
 n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , 
 n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , 
 n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , 
 n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , 
 n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , 
 n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , 
 n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , 
 n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , 
 n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , 
 n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , 
 n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , 
 n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , 
 n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , 
 n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , 
 n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , 
 n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , 
 n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , 
 n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , 
 n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , 
 n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , 
 n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , 
 n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , 
 n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , 
 n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , 
 n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , 
 n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , 
 n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , 
 n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , 
 n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , 
 n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , 
 n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , 
 n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , 
 n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , 
 n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , 
 n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , 
 n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , 
 n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , 
 n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , 
 n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , 
 n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , 
 n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , 
 n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , 
 n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , 
 n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , 
 n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , 
 n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , 
 n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , 
 n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , 
 n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , 
 n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , 
 n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , 
 n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , 
 n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , 
 n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , 
 n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , 
 n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , 
 n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , 
 n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , 
 n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , 
 n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , 
 n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , 
 n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , 
 n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , 
 n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , 
 n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , 
 n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , 
 n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , 
 n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , 
 n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , 
 n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , 
 n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , 
 n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , 
 n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , 
 n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , 
 n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , 
 n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , 
 n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , 
 n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , 
 n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , 
 n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , 
 n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , 
 n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , 
 n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , 
 n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , 
 n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , 
 n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , 
 n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , 
 n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , 
 n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , 
 n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , 
 n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , 
 n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , 
 n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , 
 n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , 
 n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , 
 n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , 
 n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , 
 n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , 
 n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , 
 n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , 
 n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , 
 n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , 
 n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , 
 n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , 
 n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , 
 n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , 
 n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , 
 n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , 
 n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , 
 n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , 
 n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , 
 n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , 
 n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , 
 n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , 
 n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , 
 n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , 
 n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , 
 n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , 
 n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , 
 n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , 
 n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , 
 n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , 
 n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , 
 n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , 
 n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , 
 n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , 
 n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , 
 n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , 
 n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , 
 n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , 
 n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , 
 n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , 
 n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , 
 n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , 
 n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , 
 n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , 
 n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , 
 n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , 
 n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , 
 n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , 
 n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , 
 n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , 
 n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , 
 n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , 
 n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , 
 n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , 
 n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , 
 n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , 
 n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , 
 n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , 
 n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , 
 n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , 
 n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , 
 n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , 
 n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , 
 n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , 
 n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , 
 n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , 
 n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , 
 n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , 
 n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , 
 n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , 
 n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , 
 n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , 
 n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , 
 n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , 
 n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , 
 n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , 
 n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , 
 n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , 
 n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , 
 n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , 
 n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , 
 n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , 
 n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , 
 n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , 
 n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , 
 n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , 
 n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , 
 n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , 
 n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , 
 n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , 
 n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , 
 n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , 
 n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , 
 n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , 
 n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , 
 n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , 
 n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , 
 n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , 
 n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , 
 n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , 
 n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , 
 n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , 
 n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , 
 n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , 
 n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , 
 n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , 
 n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , 
 n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , 
 n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , 
 n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , 
 n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , 
 n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , 
 n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , 
 n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , 
 n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , 
 n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , 
 n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , 
 n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , 
 n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , 
 n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , 
 n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , 
 n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , 
 n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , 
 n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , 
 n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , 
 n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , 
 n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , 
 n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , 
 n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , 
 n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , 
 n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , 
 n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , 
 n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , 
 n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , 
 n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , 
 n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , 
 n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , 
 n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , 
 n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , 
 n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , 
 n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , 
 n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , 
 n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , 
 n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , 
 n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , 
 n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , 
 n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , 
 n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , 
 n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , 
 n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , 
 n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , 
 n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , 
 n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , 
 n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , 
 n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , 
 n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , 
 n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , 
 n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , 
 n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , 
 n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , 
 n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , 
 n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , 
 n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , 
 n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , 
 n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , 
 n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , 
 n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , 
 n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , 
 n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , 
 n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , 
 n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , 
 n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , 
 n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , 
 n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , 
 n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , 
 n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , 
 n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , 
 n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , 
 n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , 
 n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , 
 n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , 
 n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , 
 n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , 
 n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , 
 n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , 
 n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , 
 n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , 
 n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , 
 n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , 
 n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , 
 n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , 
 n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , 
 n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , 
 n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , 
 n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , 
 n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , 
 n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , 
 n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , 
 n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , 
 n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , 
 n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , 
 n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , 
 n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , 
 n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , 
 n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , 
 n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , 
 n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , 
 n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , 
 n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , 
 n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , 
 n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , 
 n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , 
 n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , 
 n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , 
 n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , 
 n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , 
 n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , 
 n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , 
 n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , 
 n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , 
 n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , 
 n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , 
 n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , 
 n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , 
 n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , 
 n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , 
 n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , 
 n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , 
 n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , 
 n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , 
 n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , 
 n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , 
 n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , 
 n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , 
 n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , 
 n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , 
 n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , 
 n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , 
 n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , 
 n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , 
 n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , 
 n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , 
 n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , 
 n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , 
 n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , 
 n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , 
 n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , 
 n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , 
 n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , 
 n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , 
 n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , 
 n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , 
 n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , 
 n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , 
 n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , 
 n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , 
 n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , 
 n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , 
 n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , 
 n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , 
 n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , 
 n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , 
 n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , 
 n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , 
 n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , 
 n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , 
 n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , 
 n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , 
 n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , 
 n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , 
 n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , 
 n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , 
 n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , 
 n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , 
 n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , 
 n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , 
 n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , 
 n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , 
 n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , 
 n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , 
 n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , 
 n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , 
 n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , 
 n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , 
 n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , 
 n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , 
 n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , 
 n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , 
 n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , 
 n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , 
 n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , 
 n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , 
 n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , 
 n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , 
 n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , 
 n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , 
 n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , 
 n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , 
 n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , 
 n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , 
 n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , 
 n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , 
 n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , 
 n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , 
 n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , 
 n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , 
 n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , 
 n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , 
 n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , 
 n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , 
 n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , 
 n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , 
 n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , 
 n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , 
 n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , 
 n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , 
 n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , 
 n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , 
 n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , 
 n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , 
 n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , 
 n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , 
 n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , 
 n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , 
 n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , 
 n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , 
 n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , 
 n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , 
 n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , 
 n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , 
 n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , 
 n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , 
 n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , 
 n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , 
 n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , 
 n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , 
 n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , 
 n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , 
 n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , 
 n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , 
 n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , 
 n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , 
 n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , 
 n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , 
 n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , 
 n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , 
 n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , 
 n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , 
 n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , 
 n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , 
 n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , 
 n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , 
 n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , 
 n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , 
 n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , 
 n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , 
 n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , 
 n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , 
 n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , 
 n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , 
 n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , 
 n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , 
 n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , 
 n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , 
 n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , 
 n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , 
 n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , 
 n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , 
 n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , 
 n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , 
 n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , 
 n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , 
 n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , 
 n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , 
 n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , 
 n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , 
 n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , 
 n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , 
 n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , 
 n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , 
 n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , 
 n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , 
 n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , 
 n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , 
 n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , 
 n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , 
 n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , 
 n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , 
 n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , 
 n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , 
 n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , 
 n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , 
 n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , 
 n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , 
 n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , 
 n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , 
 n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , 
 n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , 
 n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , 
 n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , 
 n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , 
 n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , 
 n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , 
 n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , 
 n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , 
 n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , 
 n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , 
 n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , 
 n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , 
 n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , 
 n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , 
 n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , 
 n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , 
 n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , 
 n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , 
 n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , 
 n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , 
 n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , 
 n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , 
 n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , 
 n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , 
 n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , 
 n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , 
 n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , 
 n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , 
 n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , 
 n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , 
 n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , 
 n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , 
 n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , 
 n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , 
 n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , 
 n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , 
 n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , 
 n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , 
 n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , 
 n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , 
 n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , 
 n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , 
 n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , 
 n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , 
 n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , 
 n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , 
 n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , 
 n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , 
 n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , 
 n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , 
 n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , 
 n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , 
 n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , 
 n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , 
 n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , 
 n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , 
 n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , 
 n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , 
 n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , 
 n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , 
 n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , 
 n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , 
 n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , 
 n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , 
 n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , 
 n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , 
 n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , 
 n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , 
 n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , 
 n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , 
 n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , 
 n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , 
 n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , 
 n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , 
 n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , 
 n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , 
 n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , 
 n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , 
 n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , 
 n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , 
 n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , 
 n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , 
 n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , 
 n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , 
 n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , 
 n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , 
 n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , 
 n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , 
 n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , 
 n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , 
 n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , 
 n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , 
 n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , 
 n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , 
 n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , 
 n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , 
 n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , 
 n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , 
 n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , 
 n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , 
 n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , 
 n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , 
 n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , 
 n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , 
 n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , 
 n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , 
 n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , 
 n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , 
 n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , 
 n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , 
 n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , 
 n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , 
 n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , 
 n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , 
 n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , 
 n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , 
 n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , 
 n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , 
 n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , 
 n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , 
 n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , 
 n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , 
 n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , 
 n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , 
 n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , 
 n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , 
 n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , 
 n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , 
 n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , 
 n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , 
 n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , 
 n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , 
 n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , 
 n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , 
 n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , 
 n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , 
 n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , 
 n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , 
 n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , 
 n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , 
 n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , 
 n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , 
 n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , 
 n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , 
 n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , 
 n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , 
 n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , 
 n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , 
 n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , 
 n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , 
 n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , 
 n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , 
 n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , 
 n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , 
 n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , 
 n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , 
 n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , 
 n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , 
 n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , 
 n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , 
 n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , 
 n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , 
 n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , 
 n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , 
 n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , 
 n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , 
 n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , 
 n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , 
 n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , 
 n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , 
 n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , 
 n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , 
 n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , 
 n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , 
 n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , 
 n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , 
 n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , 
 n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , 
 n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , 
 n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , 
 n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , 
 n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , 
 n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , 
 n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , 
 n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , 
 n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , 
 n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , 
 n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , 
 n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , 
 n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , 
 n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , 
 n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , 
 n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , 
 n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , 
 n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , 
 n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , 
 n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , 
 n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , 
 n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , 
 n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , 
 n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , 
 n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , 
 n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , 
 n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , 
 n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , 
 n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , 
 n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , 
 n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , 
 n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , 
 n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , 
 n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , 
 n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , 
 n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , 
 n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , 
 n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , 
 n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , 
 n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , 
 n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , 
 n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , 
 n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , 
 n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , 
 n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , 
 n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , 
 n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , 
 n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , 
 n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , 
 n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , 
 n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , 
 n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , 
 n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , 
 n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , 
 n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , 
 n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , 
 n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , 
 n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , 
 n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , 
 n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , 
 n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , 
 n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , 
 n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , 
 n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , 
 n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , 
 n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , 
 n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , 
 n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , 
 n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , 
 n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , 
 n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , 
 n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , 
 n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , 
 n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , 
 n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , 
 n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , 
 n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , 
 n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , 
 n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , 
 n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , 
 n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , 
 n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , 
 n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , 
 n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , 
 n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , 
 n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , 
 n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , 
 n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , 
 n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , 
 n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , 
 n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , 
 n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , 
 n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , 
 n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , 
 n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , 
 n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , 
 n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , 
 n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , 
 n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , 
 n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , 
 n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , 
 n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , 
 n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , 
 n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , 
 n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , 
 n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , 
 n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , 
 n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , 
 n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , 
 n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , 
 n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , 
 n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , 
 n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , 
 n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , 
 n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , 
 n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , 
 n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , 
 n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , 
 n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , 
 n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , 
 n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , 
 n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , 
 n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , 
 n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , 
 n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , 
 n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , 
 n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , 
 n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , 
 n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , 
 n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , 
 n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , 
 n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , 
 n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , 
 n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , 
 n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , 
 n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , 
 n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , 
 n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , 
 n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , 
 n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , 
 n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , 
 n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , 
 n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , 
 n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , 
 n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , 
 n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , 
 n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , 
 n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , 
 n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , 
 n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , 
 n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , 
 n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , 
 n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , 
 n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , 
 n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , 
 n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , 
 n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , 
 n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , 
 n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , 
 n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , 
 n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , 
 n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , 
 n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , 
 n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , 
 n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , 
 n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , 
 n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , 
 n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , 
 n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , 
 n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , 
 n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , 
 n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , 
 n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , 
 n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , 
 n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , 
 n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , 
 n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , 
 n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , 
 n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , 
 n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , 
 n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , 
 n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , 
 n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , 
 n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , 
 n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , 
 n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , 
 n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , 
 n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , 
 n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , 
 n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , 
 n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , 
 n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , 
 n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , 
 n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , 
 n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , 
 n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , 
 n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , 
 n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , 
 n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , 
 n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , 
 n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , 
 n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , 
 n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , 
 n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , 
 n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , 
 n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , 
 n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , 
 n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , 
 n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , 
 n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , 
 n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , 
 n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , 
 n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , 
 n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , 
 n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , 
 n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , 
 n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , 
 n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , 
 n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , 
 n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , 
 n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , 
 n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , 
 n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , 
 n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , 
 n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , 
 n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , 
 n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , 
 n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , 
 n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , 
 n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , 
 n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , 
 n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , 
 n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , 
 n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , 
 n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , 
 n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , 
 n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , 
 n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , 
 n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , 
 n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , 
 n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , 
 n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , 
 n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , 
 n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , 
 n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , 
 n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , 
 n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , 
 n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , 
 n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , 
 n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , 
 n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , 
 n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , 
 n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , 
 n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , 
 n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , 
 n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , 
 n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , 
 n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , 
 n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , 
 n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , 
 n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , 
 n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , 
 n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , 
 n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , 
 n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , 
 n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , 
 n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , 
 n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , 
 n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , 
 n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , 
 n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , 
 n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , 
 n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , 
 n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , 
 n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , 
 n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , 
 n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , 
 n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , 
 n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , 
 n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , 
 n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , 
 n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , 
 n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , 
 n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , 
 n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , 
 n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , 
 n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , 
 n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , 
 n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , 
 n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , 
 n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , 
 n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , 
 n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , 
 n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , 
 n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , 
 n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , 
 n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , 
 n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , 
 n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , 
 n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , 
 n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , 
 n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , 
 n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , 
 n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , 
 n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , 
 n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , 
 n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , 
 n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , 
 n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , 
 n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , 
 n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , 
 n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , 
 n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , 
 n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , 
 n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , 
 n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , 
 n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , 
 n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , 
 n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , 
 n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , 
 n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , 
 n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , 
 n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , 
 n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , 
 n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , 
 n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , 
 n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , 
 n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , 
 n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , 
 n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , 
 n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , 
 n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , 
 n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , 
 n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , 
 n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , 
 n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , 
 n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , 
 n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , 
 n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , 
 n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , 
 n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , 
 n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , 
 n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , 
 n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , 
 n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , 
 n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , 
 n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , 
 n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , 
 n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , 
 n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , 
 n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , 
 n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , 
 n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , 
 n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , 
 n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , 
 n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , 
 n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , 
 n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , 
 n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , 
 n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , 
 n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , 
 n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , 
 n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , 
 n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , 
 n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , 
 n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , 
 n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , 
 n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , 
 n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , 
 n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , 
 n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , 
 n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , 
 n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , 
 n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , 
 n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , 
 n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , 
 n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , 
 n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , 
 n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , 
 n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , 
 n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , 
 n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , 
 n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , 
 n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , 
 n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , 
 n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , 
 n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , 
 n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , 
 n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , 
 n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , 
 n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , 
 n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , 
 n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , 
 n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , 
 n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , 
 n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , 
 n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , 
 n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , 
 n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , 
 n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , 
 n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , 
 n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , 
 n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , 
 n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , 
 n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , 
 n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , 
 n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , 
 n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , 
 n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , 
 n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , 
 n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , 
 n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , 
 n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , 
 n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , 
 n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , 
 n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , 
 n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , 
 n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , 
 n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , 
 n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , 
 n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , 
 n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , 
 n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , 
 n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , 
 n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , 
 n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , 
 n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , 
 n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , 
 n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , 
 n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , 
 n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , 
 n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , 
 n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , 
 n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , 
 n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , 
 n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , 
 n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , 
 n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , 
 n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , 
 n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , 
 n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , 
 n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , 
 n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , 
 n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , 
 n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , 
 n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , 
 n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , 
 n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , 
 n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , 
 n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , 
 n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , 
 n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , 
 n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , 
 n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , 
 n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , 
 n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , 
 n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , 
 n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , 
 n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , 
 n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , 
 n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , 
 n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , 
 n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , 
 n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , 
 n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , 
 n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , 
 n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , 
 n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , 
 n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , 
 n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , 
 n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , 
 n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , 
 n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , 
 n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , 
 n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , 
 n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , 
 n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , 
 n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , 
 n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , 
 n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , 
 n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , 
 n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , 
 n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , 
 n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , 
 n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , 
 n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , 
 n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , 
 n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , 
 n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , 
 n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , 
 n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , 
 n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , 
 n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , 
 n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , 
 n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , 
 n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , 
 n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , 
 n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , 
 n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , 
 n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , 
 n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , 
 n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , 
 n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , 
 n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , 
 n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , 
 n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , 
 n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , 
 n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , 
 n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , 
 n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , 
 n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , 
 n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , 
 n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , 
 n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , 
 n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , 
 n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , 
 n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , 
 n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , 
 n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , 
 n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , 
 n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , 
 n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , 
 n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , 
 n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , 
 n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , 
 n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , 
 n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , 
 n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , 
 n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , 
 n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , 
 n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , 
 n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , 
 n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , 
 n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , 
 n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , 
 n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , 
 n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , 
 n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , 
 n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , 
 n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , 
 n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , 
 n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , 
 n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , 
 n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , 
 n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , 
 n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , 
 n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , 
 n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , 
 n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , 
 n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , 
 n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , 
 n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , 
 n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , 
 n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , 
 n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , 
 n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , 
 n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , 
 n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , 
 n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , 
 n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , 
 n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , 
 n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , 
 n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , 
 n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , 
 n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , 
 n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , 
 n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , 
 n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , 
 n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , 
 n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , 
 n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , 
 n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , 
 n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , 
 n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , 
 n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , 
 n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , 
 n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , 
 n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , 
 n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , 
 n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , 
 n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , 
 n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , 
 n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , 
 n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , 
 n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , 
 n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , 
 n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , 
 n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , 
 n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , 
 n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , 
 n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , 
 n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , 
 n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , 
 n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , 
 n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , 
 n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , 
 n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , 
 n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , 
 n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , 
 n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , 
 n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , 
 n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , 
 n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , 
 n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , 
 n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , 
 n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , 
 n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , 
 n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , 
 n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , 
 n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , 
 n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , 
 n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , 
 n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , 
 n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , 
 n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , 
 n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , 
 n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , 
 n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , 
 n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , 
 n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , 
 n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , 
 n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , 
 n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , 
 n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , 
 n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , 
 n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , 
 n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , 
 n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , 
 n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , 
 n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , 
 n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , 
 n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , 
 n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , 
 n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , 
 n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , 
 n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , 
 n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , 
 n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , 
 n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , 
 n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , 
 n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , 
 n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , 
 n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , 
 n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , 
 n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , 
 n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , 
 n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , 
 n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , 
 n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , 
 n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , 
 n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , 
 n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , 
 n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , 
 n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , 
 n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , 
 n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , 
 n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , 
 n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , 
 n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , 
 n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , 
 n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , 
 n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , 
 n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , 
 n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , 
 n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , 
 n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , 
 n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , 
 n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , 
 n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , 
 n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , 
 n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , 
 n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , 
 n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , 
 n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , 
 n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , 
 n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , 
 n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , 
 n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , 
 n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , 
 n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , 
 n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , 
 n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , 
 n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , 
 n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , 
 n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , 
 n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , 
 n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , 
 n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , 
 n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , 
 n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , 
 n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , 
 n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , 
 n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , 
 n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , 
 n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , 
 n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , 
 n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , 
 n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , 
 n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , 
 n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , 
 n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , 
 n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , 
 n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , 
 n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , 
 n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , 
 n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , 
 n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , 
 n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , 
 n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , 
 n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , 
 n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , 
 n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , 
 n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , 
 n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , 
 n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , 
 n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , 
 n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , 
 n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , 
 n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , 
 n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , 
 n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , 
 n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , 
 n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , 
 n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , 
 n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , 
 n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , 
 n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , 
 n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , 
 n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , 
 n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , 
 n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , 
 n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , 
 n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , 
 n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , 
 n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , 
 n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , 
 n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , 
 n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , 
 n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , 
 n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , 
 n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , 
 n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , 
 n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , 
 n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , 
 n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , 
 n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , 
 n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , 
 n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , 
 n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , 
 n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , 
 n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , 
 n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , 
 n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , 
 n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , 
 n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , 
 n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , 
 n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , 
 n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , 
 n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , 
 n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , 
 n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , 
 n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , 
 n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , 
 n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , 
 n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , 
 n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , 
 n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , 
 n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , 
 n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , 
 n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , 
 n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , 
 n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , 
 n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , 
 n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , 
 n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , 
 n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , 
 n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , 
 n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , 
 n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , 
 n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , 
 n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , 
 n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , 
 n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , 
 n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , 
 n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , 
 n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , 
 n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , 
 n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , 
 n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , 
 n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , 
 n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , 
 n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , 
 n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , 
 n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , 
 n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , 
 n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , 
 n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , 
 n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , 
 n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , 
 n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , 
 n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , 
 n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , 
 n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , 
 n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , 
 n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , 
 n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , 
 n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , 
 n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , 
 n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , 
 n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , 
 n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , 
 n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , 
 n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , 
 n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , 
 n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , 
 n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , 
 n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , 
 n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , 
 n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , 
 n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , 
 n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , 
 n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , 
 n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , 
 n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , 
 n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , 
 n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , 
 n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , 
 n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , 
 n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , 
 n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , 
 n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , 
 n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , 
 n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , 
 n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , 
 n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , 
 n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , 
 n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , 
 n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , 
 n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , 
 n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , 
 n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , 
 n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , 
 n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , 
 n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , 
 n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , 
 n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , 
 n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , 
 n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , 
 n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , 
 n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , 
 n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , 
 n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , 
 n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , 
 n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , 
 n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , 
 n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , 
 n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , 
 n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , 
 n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , 
 n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , 
 n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , 
 n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , 
 n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , 
 n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , 
 n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , 
 n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , 
 n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , 
 n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , 
 n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , 
 n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , 
 n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , 
 n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , 
 n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , 
 n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , 
 n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , 
 n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , 
 n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , 
 n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , 
 n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , 
 n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , 
 n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , 
 n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , 
 n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , 
 n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , 
 n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , 
 n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , 
 n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , 
 n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , 
 n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , 
 n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , 
 n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , 
 n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , 
 n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , 
 n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , 
 n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , 
 n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , 
 n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , 
 n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , 
 n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , 
 n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , 
 n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , 
 n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , 
 n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , 
 n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , 
 n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , 
 n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , 
 n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , 
 n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , 
 n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , 
 n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , 
 n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , 
 n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , 
 n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , 
 n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , 
 n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , 
 n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , 
 n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , 
 n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , 
 n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , 
 n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , 
 n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , 
 n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , 
 n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , 
 n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , 
 n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , 
 n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , 
 n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , 
 n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , 
 n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , 
 n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , 
 n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , 
 n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , 
 n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , 
 n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , 
 n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , 
 n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , 
 n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , 
 n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , 
 n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , 
 n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , 
 n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , 
 n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , 
 n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , 
 n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , 
 n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , 
 n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , 
 n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , 
 n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , 
 n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , 
 n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , 
 n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , 
 n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , 
 n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , 
 n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , 
 n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , 
 n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , 
 n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , 
 n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , 
 n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , 
 n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , 
 n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , 
 n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , 
 n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , 
 n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , 
 n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , 
 n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , 
 n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , 
 n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , 
 n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , 
 n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , 
 n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , 
 n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , 
 n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , 
 n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , 
 n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , 
 n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , 
 n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , 
 n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , 
 n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , 
 n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , 
 n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , 
 n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , 
 n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , 
 n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , 
 n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , 
 n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , 
 n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , 
 n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , 
 n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , 
 n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , 
 n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , 
 n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , 
 n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , 
 n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , 
 n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , 
 n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , 
 n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , 
 n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , 
 n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , 
 n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , 
 n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , 
 n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , 
 n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , 
 n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , 
 n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , 
 n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , 
 n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , 
 n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , 
 n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , 
 n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , 
 n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , 
 n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , 
 n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , 
 n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , 
 n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , 
 n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , 
 n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , 
 n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , 
 n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , 
 n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , 
 n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , 
 n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , 
 n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , 
 n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , 
 n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , 
 n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , 
 n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , 
 n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , 
 n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , 
 n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , 
 n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , 
 n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , 
 n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , 
 n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , 
 n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , 
 n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , 
 n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , 
 n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , 
 n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , 
 n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , 
 n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , 
 n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , 
 n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , 
 n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , 
 n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , 
 n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , 
 n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , 
 n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , 
 n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , 
 n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , 
 n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , 
 n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , 
 n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , 
 n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , 
 n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , 
 n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , 
 n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , 
 n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , 
 n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , 
 n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , 
 n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , 
 n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , 
 n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , 
 n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , 
 n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , 
 n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , 
 n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , 
 n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , 
 n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , 
 n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , 
 n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , 
 n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , 
 n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , 
 n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , 
 n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , 
 n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , 
 n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , 
 n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , 
 n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , 
 n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , 
 n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , 
 n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , 
 n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , 
 n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , 
 n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , 
 n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , 
 n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , 
 n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , 
 n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , 
 n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , 
 n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , 
 n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , 
 n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , 
 n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , 
 n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , 
 n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , 
 n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , 
 n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , 
 n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , 
 n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , 
 n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , 
 n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , 
 n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , 
 n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , 
 n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , 
 n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , 
 n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , 
 n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , 
 n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , 
 n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , 
 n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , 
 n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , 
 n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , 
 n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , 
 n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , 
 n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , 
 n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , 
 n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , 
 n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , 
 n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , 
 n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , 
 n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , 
 n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , 
 n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , 
 n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , 
 n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , 
 n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , 
 n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , 
 n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , 
 n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , 
 n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , 
 n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , 
 n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , 
 n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , 
 n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , 
 n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , 
 n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , 
 n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , 
 n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , 
 n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , 
 n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , 
 n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , 
 n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , 
 n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , 
 n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , 
 n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , 
 n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , 
 n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , 
 n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , 
 n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , 
 n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , 
 n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , 
 n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , 
 n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , 
 n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , 
 n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , 
 n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , 
 n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , 
 n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , 
 n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , 
 n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , 
 n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , 
 n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , 
 n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , 
 n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , 
 n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , 
 n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , 
 n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , 
 n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , 
 n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , 
 n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , 
 n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , 
 n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , 
 n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , 
 n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , 
 n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , 
 n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , 
 n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , 
 n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , 
 n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , 
 n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , 
 n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , 
 n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , 
 n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , 
 n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , 
 n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , 
 n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , 
 n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , 
 n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , 
 n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , 
 n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , 
 n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , 
 n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , 
 n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , 
 n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , 
 n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , 
 n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , 
 n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , 
 n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , 
 n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , 
 n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , 
 n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , 
 n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , 
 n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , 
 n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , 
 n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , 
 n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , 
 n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , 
 n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , 
 n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , 
 n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , 
 n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , 
 n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , 
 n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , 
 n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , 
 n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , 
 n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , 
 n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , 
 n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , 
 n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , 
 n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , 
 n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , 
 n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , 
 n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , 
 n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , 
 n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , 
 n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , 
 n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , 
 n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , 
 n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , 
 n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , 
 n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , 
 n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , 
 n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , 
 n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , 
 n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , 
 n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , 
 n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , 
 n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , 
 n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , 
 n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , 
 n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , 
 n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , 
 n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , 
 n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , 
 n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , 
 n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , 
 n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , 
 n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , 
 n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , 
 n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , 
 n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , 
 n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , 
 n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , 
 n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , 
 n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , 
 n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , 
 n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , 
 n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , 
 n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , 
 n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , 
 n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , 
 n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , 
 n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , 
 n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , 
 n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , 
 n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , 
 n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , 
 n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , 
 n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , 
 n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , 
 n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , 
 n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , 
 n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , 
 n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , 
 n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , 
 n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , 
 n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , 
 n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , 
 n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , 
 n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , 
 n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , 
 n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , 
 n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , 
 n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , 
 n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , 
 n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , 
 n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , 
 n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , 
 n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , 
 n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , 
 n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , 
 n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , 
 n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , 
 n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , 
 n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , 
 n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , 
 n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , 
 n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , 
 n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , 
 n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , 
 n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , 
 n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , 
 n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , 
 n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , 
 n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , 
 n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , 
 n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , 
 n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , 
 n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , 
 n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , 
 n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , 
 n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , 
 n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , 
 n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , 
 n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , 
 n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , 
 n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , 
 n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , 
 n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , 
 n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , 
 n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , 
 n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , 
 n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , 
 n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , 
 n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , 
 n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , 
 n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , 
 n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , 
 n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , 
 n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , 
 n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , 
 n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , 
 n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , 
 n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , 
 n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , 
 n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , 
 n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , 
 n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , 
 n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , 
 n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , 
 n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , 
 n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , 
 n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , 
 n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , 
 n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , 
 n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , 
 n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , 
 n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , 
 n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , 
 n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , 
 n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , 
 n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , 
 n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , 
 n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , 
 n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , 
 n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , 
 n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , 
 n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , 
 n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , 
 n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , 
 n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , 
 n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , 
 n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , 
 n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , 
 n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , 
 n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , 
 n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , 
 n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , 
 n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , 
 n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , 
 n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , 
 n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , 
 n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , 
 n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , 
 n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , 
 n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , 
 n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , 
 n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , 
 n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , 
 n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , 
 n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , 
 n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , 
 n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , 
 n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , 
 n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , 
 n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , 
 n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , 
 n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , 
 n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , 
 n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , 
 n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , 
 n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , 
 n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , 
 n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , 
 n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , 
 n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , 
 n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , 
 n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , 
 n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , 
 n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , 
 n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , 
 n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , 
 n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , 
 n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , 
 n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , 
 n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , 
 n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , 
 n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , 
 n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , 
 n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , 
 n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , 
 n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , 
 n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , 
 n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , 
 n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , 
 n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , 
 n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , 
 n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , 
 n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , 
 n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , 
 n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , 
 n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , 
 n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , 
 n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , 
 n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , 
 n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , 
 n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , 
 n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , 
 n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , 
 n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , 
 n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , 
 n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , 
 n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , 
 n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , 
 n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , 
 n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , 
 n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , 
 n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , 
 n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , 
 n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , 
 n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , 
 n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , 
 n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , 
 n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , 
 n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , 
 n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , 
 n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , 
 n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , 
 n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , 
 n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , 
 n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , 
 n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , 
 n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , 
 n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , 
 n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , 
 n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , 
 n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , 
 n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , 
 n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , 
 n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , 
 n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , 
 n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , 
 n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , 
 n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , 
 n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , 
 n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , 
 n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , 
 n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , 
 n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , 
 n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , 
 n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , 
 n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , 
 n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , 
 n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , 
 n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , 
 n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , 
 n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , 
 n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , 
 n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , 
 n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , 
 n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , 
 n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , 
 n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , 
 n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , 
 n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , 
 n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , 
 n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , 
 n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , 
 n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , 
 n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , 
 n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , 
 n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , 
 n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , 
 n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , 
 n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , 
 n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , 
 n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , 
 n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , 
 n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , 
 n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , 
 n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , 
 n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , 
 n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , 
 n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , 
 n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , 
 n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , 
 n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , 
 n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , 
 n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , 
 n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , 
 n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , 
 n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , 
 n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , 
 n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , 
 n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , 
 n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , 
 n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , 
 n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , 
 n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , 
 n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , 
 n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , 
 n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , 
 n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , 
 n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , 
 n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , 
 n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , 
 n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , 
 n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , 
 n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , 
 n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , 
 n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , 
 n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , 
 n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , 
 n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , 
 n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , 
 n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , 
 n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , 
 n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , 
 n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , 
 n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , 
 n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , 
 n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , 
 n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , 
 n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , 
 n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , 
 n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , 
 n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , 
 n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , 
 n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , 
 n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , 
 n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , 
 n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , 
 n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , 
 n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , 
 n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , 
 n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , 
 n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , 
 n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , 
 n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , 
 n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , 
 n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , 
 n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , 
 n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , 
 n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , 
 n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , 
 n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , 
 n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , 
 n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , 
 n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , 
 n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , 
 n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , 
 n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , 
 n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , 
 n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , 
 n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , 
 n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , 
 n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , 
 n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , 
 n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , 
 n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , 
 n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , 
 n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , 
 n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , 
 n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , 
 n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , 
 n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , 
 n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , 
 n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , 
 n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , 
 n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , 
 n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , 
 n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , 
 n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , 
 n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , 
 n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , 
 n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , 
 n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , 
 n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , 
 n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , 
 n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , 
 n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , 
 n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , 
 n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , 
 n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , 
 n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , 
 n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , 
 n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , 
 n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , 
 n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , 
 n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , 
 n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , 
 n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , 
 n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , 
 n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , 
 n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , 
 n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , 
 n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , 
 n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , 
 n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , 
 n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , 
 n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , 
 n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , 
 n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , 
 n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , 
 n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , 
 n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , 
 n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , 
 n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , 
 n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , 
 n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , 
 n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , 
 n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , 
 n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , 
 n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , 
 n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , 
 n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , 
 n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , 
 n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , 
 n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , 
 n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , 
 n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , 
 n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , 
 n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , 
 n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , 
 n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , 
 n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , 
 n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , 
 n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , 
 n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , 
 n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , 
 n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , 
 n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , 
 n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , 
 n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , 
 n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , 
 n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , 
 n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , 
 n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , 
 n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , 
 n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , 
 n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , 
 n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , 
 n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , 
 n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , 
 n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , 
 n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , 
 n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , 
 n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , 
 n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , 
 n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , 
 n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , 
 n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , 
 n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , 
 n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , 
 n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , 
 n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , 
 n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , 
 n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , 
 n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , 
 n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , 
 n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , 
 n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , 
 n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , 
 n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , 
 n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , 
 n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , 
 n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , 
 n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , 
 n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , 
 n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , 
 n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , 
 n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , 
 n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , 
 n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , 
 n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , 
 n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , 
 n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , 
 n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , 
 n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , 
 n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , 
 n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , 
 n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , 
 n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , 
 n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , 
 n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , 
 n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , 
 n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , 
 n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , 
 n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , 
 n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , 
 n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , 
 n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , 
 n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , 
 n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , 
 n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , 
 n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , 
 n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , 
 n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , 
 n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , 
 n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , 
 n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , 
 n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , 
 n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , 
 n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , 
 n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , 
 n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , 
 n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , 
 n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , 
 n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , 
 n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , 
 n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , 
 n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , 
 n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , 
 n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , 
 n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , 
 n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , 
 n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , 
 n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , 
 n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , 
 n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , 
 n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , 
 n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , 
 n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , 
 n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , 
 n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , 
 n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , 
 n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , 
 n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , 
 n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , 
 n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , 
 n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , 
 n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , 
 n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , 
 n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , 
 n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , 
 n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , 
 n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , 
 n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , 
 n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , 
 n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , 
 n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , 
 n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , 
 n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , 
 n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , 
 n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , 
 n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , 
 n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , 
 n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , 
 n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , 
 n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , 
 n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , 
 n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , 
 n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , 
 n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , 
 n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , 
 n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , 
 n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , 
 n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , 
 n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , 
 n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , 
 n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , 
 n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , 
 n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , 
 n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , 
 n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , 
 n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , 
 n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , 
 n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , 
 n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , 
 n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , 
 n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , 
 n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , 
 n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , 
 n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , 
 n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , 
 n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , 
 n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , 
 n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , 
 n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , 
 n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , 
 n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , 
 n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , 
 n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , 
 n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , 
 n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , 
 n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , 
 n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , 
 n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , 
 n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , 
 n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , 
 n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , 
 n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , 
 n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , 
 n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , 
 n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , 
 n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , 
 n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , 
 n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , 
 n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , 
 n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , 
 n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , 
 n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , 
 n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , 
 n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , 
 n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , 
 n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , 
 n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , 
 n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , 
 n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , 
 n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , 
 n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , 
 n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , 
 n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , 
 n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , 
 n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , 
 n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , 
 n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , 
 n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , 
 n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , 
 n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , 
 n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , 
 n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , 
 n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , 
 n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , 
 n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , 
 n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , 
 n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , 
 n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , 
 n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , 
 n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , 
 n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , 
 n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , 
 n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , 
 n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , 
 n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , 
 n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , 
 n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , 
 n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , 
 n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , 
 n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , 
 n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , 
 n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , 
 n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , 
 n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , 
 n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , 
 n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , 
 n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , 
 n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , 
 n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , 
 n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , 
 n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , 
 n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , 
 n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , 
 n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , 
 n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , 
 n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , 
 n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , 
 n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , 
 n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , 
 n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , 
 n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , 
 n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , 
 n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , 
 n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , 
 n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , 
 n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , 
 n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , 
 n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , 
 n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , 
 n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , 
 n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , 
 n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , 
 n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , 
 n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , 
 n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , 
 n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , 
 n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , 
 n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , 
 n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , 
 n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , 
 n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , 
 n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , 
 n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , 
 n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , 
 n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , 
 n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , 
 n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , 
 n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , 
 n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , 
 n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , 
 n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , 
 n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , 
 n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , 
 n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , 
 n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , 
 n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , 
 n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , 
 n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , 
 n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , 
 n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , 
 n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , 
 n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , 
 n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , 
 n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , 
 n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , 
 n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , 
 n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , 
 n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , 
 n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , 
 n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , 
 n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , 
 n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , 
 n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , 
 n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , 
 n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , 
 n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , 
 n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , 
 n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , 
 n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , 
 n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , 
 n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , 
 n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , 
 n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , 
 n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , 
 n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , 
 n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , 
 n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , 
 n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , 
 n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , 
 n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , 
 n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , 
 n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , 
 n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , 
 n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , 
 n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , 
 n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , 
 n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , 
 n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , 
 n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , 
 n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , 
 n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , 
 n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , 
 n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , 
 n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , 
 n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , 
 n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , 
 n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , 
 n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , 
 n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , 
 n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , 
 n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , 
 n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , 
 n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , 
 n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , 
 n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , 
 n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , 
 n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , 
 n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , 
 n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , 
 n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , 
 n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , 
 n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , 
 n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , 
 n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , 
 n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , 
 n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , 
 n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , 
 n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , 
 n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , 
 n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , 
 n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , 
 n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , 
 n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , 
 n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , 
 n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , 
 n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , 
 n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , 
 n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , 
 n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , 
 n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , 
 n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , 
 n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , 
 n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , 
 n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , 
 n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , 
 n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , 
 n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , 
 n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , 
 n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , 
 n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , 
 n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , 
 n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , 
 n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , 
 n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , 
 n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , 
 n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , 
 n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , 
 n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , 
 n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , 
 n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , 
 n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , 
 n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , 
 n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , 
 n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , 
 n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , 
 n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , 
 n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , 
 n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , 
 n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , 
 n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , 
 n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , 
 n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , 
 n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , 
 n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , 
 n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , 
 n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , 
 n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , 
 n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , 
 n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , 
 n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , 
 n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , 
 n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , 
 n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , 
 n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , 
 n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , 
 n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , 
 n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , 
 n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , 
 n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , 
 n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , 
 n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , 
 n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , 
 n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , 
 n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , 
 n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , 
 n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , 
 n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , 
 n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , 
 n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , 
 n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , 
 n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , 
 n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , 
 n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , 
 n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , 
 n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , 
 n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , 
 n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , 
 n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , 
 n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , 
 n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , 
 n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , 
 n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , 
 n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , 
 n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , 
 n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , 
 n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , 
 n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , 
 n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , 
 n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , 
 n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , 
 n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , 
 n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , 
 n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , 
 n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , 
 n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , 
 n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , 
 n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , 
 n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , 
 n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , 
 n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , 
 n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , 
 n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , 
 n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , 
 n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , 
 n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , 
 n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , 
 n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , 
 n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , 
 n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , 
 n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , 
 n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , 
 n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , 
 n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , 
 n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , 
 n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , 
 n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , 
 n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , 
 n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , 
 n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , 
 n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , 
 n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , 
 n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , 
 n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , 
 n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , 
 n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , 
 n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , 
 n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , 
 n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , 
 n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , 
 n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , 
 n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , 
 n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , 
 n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , 
 n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , 
 n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , 
 n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , 
 n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , 
 n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , 
 n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , 
 n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , 
 n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , 
 n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , 
 n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , 
 n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , 
 n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , 
 n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , 
 n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , 
 n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , 
 n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , 
 n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , 
 n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , 
 n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , 
 n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , 
 n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , 
 n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , 
 n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , 
 n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , 
 n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , 
 n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , 
 n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , 
 n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , 
 n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , 
 n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , 
 n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , 
 n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , 
 n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , 
 n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , 
 n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , 
 n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , 
 n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , 
 n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , 
 n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , 
 n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , 
 n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , 
 n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , 
 n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , 
 n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , 
 n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , 
 n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , 
 n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , 
 n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , 
 n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , 
 n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , 
 n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , 
 n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , 
 n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , 
 n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , 
 n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , 
 n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , 
 n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , 
 n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , 
 n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , 
 n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , 
 n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , 
 n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , 
 n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , 
 n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , 
 n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , 
 n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , 
 n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , 
 n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , 
 n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , 
 n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , 
 n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , 
 n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , 
 n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , 
 n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , 
 n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , 
 n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , 
 n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , 
 n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , 
 n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , 
 n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , 
 n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , 
 n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , 
 n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , 
 n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , 
 n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , 
 n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , 
 n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , 
 n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , 
 n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , 
 n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , 
 n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , 
 n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , 
 n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , 
 n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , 
 n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , 
 n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , 
 n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , 
 n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , 
 n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , 
 n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , 
 n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , 
 n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , 
 n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , 
 n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , 
 n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , 
 n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , 
 n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , 
 n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , 
 n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , 
 n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , 
 n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , 
 n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , 
 n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , 
 n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , 
 n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , 
 n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , 
 n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , 
 n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , 
 n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , 
 n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , 
 n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , 
 n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , 
 n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , 
 n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , 
 n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , 
 n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , 
 n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , 
 n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , 
 n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , 
 n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , 
 n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , 
 n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , 
 n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , 
 n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , 
 n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , 
 n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , 
 n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , 
 n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , 
 n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , 
 n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , 
 n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , 
 n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , 
 n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , 
 n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , 
 n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , 
 n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , 
 n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , 
 n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , 
 n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , 
 n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , 
 n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , 
 n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , 
 n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , 
 n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , 
 n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , 
 n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , 
 n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , 
 n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , 
 n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , 
 n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , 
 n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , 
 n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , 
 n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , 
 n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , 
 n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , 
 n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , 
 n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , 
 n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , 
 n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , 
 n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , 
 n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , 
 n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , 
 n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , 
 n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , 
 n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , 
 n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , 
 n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , 
 n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , 
 n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , 
 n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , 
 n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , 
 n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , 
 n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , 
 n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , 
 n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , 
 n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , 
 n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , 
 n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , 
 n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , 
 n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , 
 n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , 
 n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , 
 n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , 
 n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , 
 n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , 
 n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , 
 n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , 
 n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , 
 n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , 
 n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , 
 n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , 
 n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , 
 n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , 
 n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , 
 n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , 
 n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , 
 n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , 
 n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , 
 n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , 
 n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , 
 n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , 
 n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , 
 n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , 
 n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , 
 n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , 
 n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , 
 n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , 
 n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , 
 n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , 
 n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , 
 n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , 
 n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , 
 n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , 
 n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , 
 n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , 
 n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , 
 n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , 
 n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , 
 n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , 
 n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , 
 n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , 
 n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , 
 n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , 
 n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , 
 n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , 
 n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , 
 n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , 
 n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , 
 n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , 
 n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , 
 n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , 
 n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , 
 n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , 
 n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , 
 n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , 
 n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , 
 n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , 
 n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , 
 n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , 
 n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , 
 n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , 
 n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , 
 n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , 
 n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , 
 n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , 
 n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , 
 n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , 
 n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , 
 n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , 
 n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , 
 n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , 
 n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , 
 n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , 
 n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , 
 n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , 
 n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , 
 n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , 
 n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , 
 n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , 
 n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , 
 n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , 
 n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , 
 n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , 
 n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , 
 n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , 
 n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , 
 n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , 
 n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , 
 n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , 
 n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , 
 n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , 
 n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , 
 n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , 
 n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , 
 n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , 
 n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , 
 n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , 
 n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , 
 n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , 
 n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , 
 n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , 
 n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , 
 n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , 
 n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , 
 n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , 
 n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , 
 n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , 
 n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , 
 n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , 
 n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , 
 n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , 
 n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , 
 n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , 
 n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , 
 n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , 
 n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , 
 n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , 
 n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , 
 n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , 
 n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , 
 n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , 
 n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , 
 n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , 
 n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , 
 n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , 
 n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , 
 n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , 
 n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , 
 n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , 
 n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , 
 n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , 
 n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , 
 n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , 
 n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , 
 n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , 
 n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , 
 n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , 
 n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , 
 n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , 
 n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , 
 n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , 
 n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , 
 n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , 
 n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , 
 n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , 
 n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , 
 n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , 
 n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , 
 n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , 
 n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , 
 n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , 
 n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , 
 n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , 
 n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , 
 n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , 
 n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , 
 n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , 
 n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , 
 n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , 
 n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , 
 n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , 
 n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , 
 n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , 
 n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , 
 n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , 
 n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , 
 n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , 
 n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , 
 n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , 
 n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , 
 n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , 
 n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , 
 n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , 
 n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , 
 n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , 
 n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , 
 n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , 
 n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , 
 n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , 
 n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , 
 n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , 
 n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , 
 n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , 
 n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , 
 n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , 
 n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , 
 n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , 
 n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , 
 n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , 
 n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , 
 n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , 
 n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , 
 n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , 
 n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , 
 n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , 
 n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , 
 n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , 
 n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , 
 n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , 
 n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , 
 n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , 
 n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , 
 n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , 
 n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , 
 n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , 
 n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , 
 n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , 
 n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , 
 n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , 
 n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , 
 n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , 
 n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , 
 n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , 
 n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , 
 n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , 
 n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , 
 n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , 
 n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , 
 n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , 
 n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , 
 n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , 
 n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , 
 n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , 
 n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , 
 n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , 
 n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , 
 n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , 
 n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , 
 n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , 
 n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , 
 n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , 
 n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , 
 n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , 
 n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , 
 n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , 
 n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , 
 n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , 
 n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , 
 n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , 
 n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , 
 n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , 
 n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , 
 n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , 
 n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , 
 n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , 
 n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , 
 n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , 
 n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , 
 n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , 
 n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , 
 n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , 
 n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , 
 n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , 
 n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , 
 n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , 
 n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , 
 n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , 
 n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , 
 n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , 
 n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , 
 n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , 
 n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , 
 n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , 
 n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , 
 n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , 
 n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , 
 n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , 
 n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , 
 n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , 
 n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , 
 n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , 
 n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , 
 n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , 
 n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , 
 n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , 
 n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , 
 n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , 
 n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , 
 n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , 
 n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , 
 n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , 
 n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , 
 n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , 
 n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , 
 n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , 
 n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , 
 n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , 
 n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , 
 n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , 
 n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , 
 n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , 
 n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , 
 n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , 
 n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , 
 n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , 
 n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , 
 n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , 
 n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , 
 n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , 
 n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , 
 n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , 
 n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , 
 n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , 
 n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , 
 n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , 
 n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , 
 n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , 
 n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , 
 n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , 
 n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , 
 n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , 
 n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , 
 n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , 
 n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , 
 n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , 
 n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , 
 n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , 
 n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , 
 n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , 
 n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , 
 n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , 
 n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , 
 n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , 
 n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , 
 n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , 
 n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , 
 n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , 
 n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , 
 n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , 
 n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , 
 n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , 
 n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , 
 n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , 
 n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , 
 n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , 
 n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , 
 n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , 
 n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , 
 n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , 
 n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , 
 n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , 
 n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , 
 n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , 
 n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , 
 n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , 
 n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , 
 n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , 
 n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , 
 n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , 
 n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , 
 n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , 
 n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , 
 n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , 
 n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , 
 n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , 
 n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , 
 n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , 
 n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , 
 n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , 
 n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , 
 n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , 
 n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , 
 n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , 
 n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , 
 n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , 
 n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , 
 n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , 
 n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , 
 n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , 
 n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , 
 n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , 
 n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , 
 n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , 
 n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , 
 n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , 
 n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , 
 n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , 
 n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , 
 n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , 
 n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , 
 n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , 
 n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , 
 n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , 
 n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , 
 n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , 
 n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , 
 n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , 
 n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , 
 n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , 
 n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , 
 n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , 
 n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , 
 n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , 
 n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , 
 n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , 
 n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , 
 n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , 
 n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , 
 n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , 
 n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , 
 n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , 
 n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , 
 n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , 
 n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , 
 n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , 
 n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , 
 n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , 
 n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , 
 n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , 
 n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , 
 n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , 
 n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , 
 n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , 
 n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , 
 n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , 
 n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , 
 n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , 
 n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , 
 n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , 
 n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , 
 n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , 
 n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , 
 n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , 
 n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , 
 n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , 
 n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , 
 n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , 
 n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , 
 n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , 
 n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , 
 n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , 
 n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , 
 n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , 
 n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , 
 n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , 
 n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , 
 n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , 
 n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , 
 n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , 
 n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , 
 n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , 
 n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , 
 n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , 
 n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , 
 n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , 
 n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , 
 n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , 
 n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , 
 n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , 
 n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , 
 n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , 
 n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , 
 n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , 
 n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , 
 n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , 
 n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , 
 n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , 
 n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , 
 n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , 
 n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , 
 n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , 
 n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , 
 n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , 
 n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , 
 n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , 
 n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , 
 n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , 
 n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , 
 n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , 
 n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , 
 n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , 
 n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , 
 n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , 
 n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , 
 n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , 
 n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , 
 n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , 
 n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , 
 n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , 
 n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , 
 n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , 
 n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , 
 n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , 
 n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , 
 n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , 
 n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , 
 n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , 
 n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , 
 n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , 
 n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , 
 n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , 
 n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , 
 n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , 
 n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , 
 n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , 
 n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , 
 n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , 
 n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , 
 n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , 
 n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , 
 n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , 
 n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , 
 n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , 
 n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , 
 n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , 
 n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , 
 n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , 
 n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , 
 n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , 
 n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , 
 n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , 
 n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , 
 n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , 
 n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , 
 n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , 
 n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , 
 n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , 
 n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , 
 n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , 
 n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , 
 n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , 
 n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , 
 n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , 
 n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , 
 n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , 
 n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , 
 n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , 
 n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , 
 n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , 
 n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , 
 n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , 
 n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , 
 n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , 
 n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , 
 n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , 
 n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , 
 n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , 
 n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , 
 n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , 
 n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , 
 n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , 
 n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , 
 n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , 
 n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , 
 n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , 
 n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , 
 n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , 
 n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , 
 n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , 
 n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , 
 n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , 
 n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , 
 n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , 
 n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , 
 n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , 
 n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , 
 n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , 
 n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , 
 n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , 
 n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , 
 n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , 
 n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , 
 n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , 
 n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , 
 n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , 
 n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , 
 n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , 
 n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , 
 n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , 
 n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , 
 n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , 
 n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , 
 n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , 
 n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , 
 n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , 
 n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , 
 n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , 
 n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , 
 n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , 
 n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , 
 n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , 
 n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , 
 n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , 
 n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , 
 n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , 
 n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , 
 n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , 
 n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , 
 n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , 
 n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , 
 n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , 
 n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , 
 n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , 
 n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , 
 n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , 
 n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , 
 n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , 
 n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , 
 n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , 
 n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , 
 n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , 
 n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , 
 n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , 
 n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , 
 n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , 
 n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , 
 n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , 
 n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , 
 n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , 
 n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , 
 n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , 
 n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , 
 n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , 
 n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , 
 n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , 
 n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , 
 n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , 
 n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , 
 n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , 
 n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , 
 n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , 
 n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , 
 n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , 
 n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , 
 n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , 
 n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , 
 n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , 
 n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , 
 n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , 
 n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , 
 n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , 
 n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , 
 n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , 
 n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , 
 n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , 
 n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , 
 n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , 
 n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , 
 n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , 
 n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , 
 n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , 
 n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , 
 n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , 
 n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , 
 n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , 
 n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , 
 n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , 
 n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , 
 n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , 
 n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , 
 n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , 
 n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , 
 n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , 
 n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , 
 n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , 
 n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , 
 n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , 
 n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , 
 n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , 
 n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , 
 n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , 
 n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , 
 n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , 
 n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , 
 n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , 
 n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , 
 n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , 
 n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , 
 n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , 
 n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , 
 n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , 
 n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , 
 n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , 
 n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , 
 n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , 
 n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , 
 n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , 
 n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , 
 n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , 
 n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , 
 n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , 
 n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , 
 n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , 
 n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , 
 n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , 
 n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , 
 n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , 
 n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , 
 n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , 
 n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , 
 n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , 
 n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , 
 n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , 
 n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , 
 n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , 
 n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , 
 n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , 
 n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , 
 n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , 
 n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , 
 n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , 
 n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , 
 n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , 
 n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , 
 n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , 
 n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , 
 n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , 
 n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , 
 n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , 
 n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , 
 n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , 
 n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , 
 n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , 
 n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , 
 n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , 
 n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , 
 n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , 
 n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , 
 n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , 
 n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , 
 n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , 
 n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , 
 n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , 
 n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , 
 n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , 
 n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , 
 n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , 
 n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , 
 n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , 
 n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , 
 n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , 
 n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , 
 n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , 
 n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , 
 n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , 
 n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , 
 n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , 
 n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , 
 n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , 
 n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , 
 n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , 
 n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , 
 n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , 
 n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , 
 n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , 
 n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , 
 n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , 
 n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , 
 n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , 
 n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , 
 n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , 
 n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , 
 n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , 
 n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , 
 n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , 
 n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , 
 n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , 
 n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , 
 n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , 
 n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , 
 n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , 
 n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , 
 n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , 
 n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , 
 n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , 
 n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , 
 n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , 
 n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , 
 n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , 
 n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , 
 n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , 
 n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , 
 n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , 
 n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , 
 n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , 
 n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , 
 n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , 
 n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , 
 n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , 
 n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , 
 n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , 
 n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , 
 n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , 
 n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , 
 n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , 
 n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , 
 n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , 
 n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , 
 n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , 
 n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , 
 n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , 
 n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , 
 n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , 
 n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , 
 n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , 
 n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , 
 n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , 
 n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , 
 n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , 
 n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , 
 n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , 
 n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , 
 n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , 
 n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , 
 n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , 
 n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , 
 n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , 
 n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , 
 n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , 
 n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , 
 n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , 
 n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , 
 n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , 
 n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , 
 n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , 
 n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , 
 n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , 
 n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , 
 n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , 
 n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , 
 n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , 
 n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , 
 n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , 
 n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , 
 n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , 
 n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , 
 n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , 
 n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , 
 n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , 
 n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , 
 n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , 
 n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , 
 n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , 
 n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , 
 n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , 
 n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , 
 n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , 
 n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , 
 n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , 
 n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , 
 n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , 
 n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , 
 n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , 
 n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , 
 n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , 
 n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , 
 n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , 
 n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , 
 n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , 
 n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , 
 n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , 
 n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , 
 n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , 
 n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , 
 n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , 
 n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , 
 n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , 
 n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , 
 n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , 
 n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , 
 n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , 
 n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , 
 n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , 
 n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , 
 n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , 
 n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , 
 n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , 
 n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , 
 n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , 
 n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , 
 n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , 
 n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , 
 n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , 
 n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , 
 n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , 
 n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , 
 n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , 
 n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , 
 n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , 
 n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , 
 n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , 
 n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , 
 n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , 
 n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , 
 n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , 
 n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , 
 n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , 
 n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , 
 n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , 
 n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , 
 n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , 
 n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , 
 n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , 
 n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , 
 n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , 
 n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , 
 n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , 
 n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , 
 n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , 
 n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , 
 n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , 
 n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , 
 n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , 
 n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , 
 n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , 
 n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , 
 n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , 
 n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , 
 n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , 
 n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , 
 n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , 
 n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , 
 n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , 
 n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , 
 n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , 
 n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , 
 n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , 
 n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , 
 n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , 
 n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , 
 n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , 
 n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , 
 n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , 
 n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , 
 n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , 
 n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , 
 n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , 
 n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , 
 n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , 
 n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , 
 n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , 
 n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , 
 n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , 
 n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , 
 n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , 
 n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , 
 n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , 
 n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , 
 n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , 
 n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , 
 n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , 
 n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , 
 n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , 
 n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , 
 n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , 
 n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , 
 n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , 
 n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , 
 n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , 
 n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , 
 n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , 
 n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , 
 n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , 
 n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , 
 n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , 
 n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , 
 n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , 
 n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , 
 n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , 
 n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , 
 n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , 
 n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , 
 n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , 
 n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , 
 n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , 
 n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , 
 n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , 
 n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , 
 n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , 
 n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , 
 n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , 
 n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , 
 n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , 
 n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , 
 n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , 
 n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , 
 n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , 
 n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , 
 n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , 
 n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , 
 n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , 
 n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , 
 n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , 
 n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , 
 n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , 
 n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , 
 n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , 
 n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , 
 n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , 
 n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , 
 n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , 
 n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , 
 n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , 
 n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , 
 n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , 
 n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , 
 n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , 
 n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , 
 n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , 
 n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , 
 n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , 
 n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , 
 n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , 
 n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , 
 n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , 
 n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , 
 n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , 
 n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , 
 n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , 
 n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , 
 n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , 
 n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , 
 n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , 
 n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , 
 n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , 
 n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , 
 n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , 
 n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , 
 n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , 
 n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , 
 n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , 
 n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , 
 n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , 
 n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , 
 n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , 
 n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , 
 n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , 
 n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , 
 n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , 
 n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , 
 n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , 
 n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , 
 n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , 
 n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , 
 n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , 
 n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , 
 n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , 
 n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , 
 n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , 
 n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , 
 n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , 
 n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , 
 n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , 
 n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , 
 n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , 
 n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , 
 n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , 
 n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , 
 n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , 
 n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , 
 n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , 
 n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , 
 n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , 
 n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , 
 n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , 
 n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , 
 n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , 
 n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , 
 n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , 
 n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , 
 n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , 
 n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , 
 n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , 
 n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , 
 n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , 
 n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , 
 n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , 
 n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , 
 n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , 
 n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , 
 n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , 
 n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , 
 n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , 
 n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , 
 n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , 
 n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , 
 n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , 
 n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , 
 n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , 
 n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , 
 n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , 
 n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , 
 n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , 
 n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , 
 n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , 
 n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , 
 n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , 
 n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , 
 n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , 
 n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , 
 n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , 
 n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , 
 n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , 
 n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , 
 n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , 
 n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , 
 n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , 
 n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , 
 n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , 
 n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , 
 n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , 
 n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , 
 n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , 
 n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , 
 n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , 
 n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , 
 n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , 
 n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , 
 n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , 
 n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , 
 n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , 
 n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , 
 n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , 
 n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , 
 n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , 
 n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , 
 n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , 
 n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , 
 n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , 
 n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , 
 n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , 
 n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , 
 n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , 
 n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , 
 n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , 
 n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , 
 n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , 
 n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , 
 n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , 
 n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , 
 n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , 
 n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , 
 n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , 
 n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , 
 n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , 
 n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , 
 n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , 
 n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , 
 n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , 
 n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , 
 n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , 
 n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , 
 n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , 
 n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , 
 n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , 
 n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , 
 n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , 
 n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , 
 n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , 
 n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , 
 n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , 
 n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , 
 n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , 
 n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , 
 n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , 
 n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , 
 n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , 
 n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , 
 n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , 
 n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , 
 n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , 
 n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , 
 n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , 
 n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , 
 n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , 
 n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , 
 n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , 
 n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , 
 n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , 
 n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , 
 n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , 
 n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , 
 n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , 
 n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , 
 n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , 
 n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , 
 n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , 
 n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , 
 n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , 
 n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , 
 n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , 
 n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , 
 n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , 
 n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , 
 n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , 
 n54145 , n54146 , n54147 , n54148 , n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , 
 n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , 
 n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , 
 n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , 
 n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , 
 n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , 
 n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , 
 n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , 
 n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , 
 n54235 , n54236 , n54237 , n54238 , n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , 
 n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , 
 n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , 
 n54265 , n54266 , n54267 , n54268 , n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , 
 n54275 , n54276 , n54277 , n54278 , n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , 
 n54285 , n54286 , n54287 , n54288 , n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , 
 n54295 , n54296 , n54297 , n54298 , n54299 , n54300 , n54301 , n54302 , n54303 , n54304 , 
 n54305 , n54306 , n54307 , n54308 , n54309 , n54310 , n54311 , n54312 , n54313 , n54314 , 
 n54315 , n54316 , n54317 , n54318 , n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , 
 n54325 , n54326 , n54327 , n54328 , n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , 
 n54335 , n54336 , n54337 , n54338 , n54339 , n54340 , n54341 , n54342 , n54343 , n54344 , 
 n54345 , n54346 , n54347 , n54348 , n54349 , n54350 , n54351 , n54352 , n54353 , n54354 , 
 n54355 , n54356 , n54357 , n54358 , n54359 , n54360 , n54361 , n54362 , n54363 , n54364 , 
 n54365 , n54366 , n54367 , n54368 , n54369 , n54370 , n54371 , n54372 , n54373 , n54374 , 
 n54375 , n54376 , n54377 , n54378 , n54379 , n54380 , n54381 , n54382 , n54383 , n54384 , 
 n54385 , n54386 , n54387 , n54388 , n54389 , n54390 , n54391 , n54392 , n54393 , n54394 , 
 n54395 , n54396 , n54397 , n54398 , n54399 , n54400 , n54401 , n54402 , n54403 , n54404 , 
 n54405 , n54406 , n54407 , n54408 , n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , 
 n54415 , n54416 , n54417 , n54418 , n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , 
 n54425 , n54426 , n54427 , n54428 , n54429 , n54430 , n54431 , n54432 , n54433 , n54434 , 
 n54435 , n54436 , n54437 , n54438 , n54439 , n54440 , n54441 , n54442 , n54443 , n54444 , 
 n54445 , n54446 , n54447 , n54448 , n54449 , n54450 , n54451 , n54452 , n54453 , n54454 , 
 n54455 , n54456 , n54457 , n54458 , n54459 , n54460 , n54461 , n54462 , n54463 , n54464 , 
 n54465 , n54466 , n54467 , n54468 , n54469 , n54470 , n54471 , n54472 , n54473 , n54474 , 
 n54475 , n54476 , n54477 , n54478 , n54479 , n54480 , n54481 , n54482 , n54483 , n54484 , 
 n54485 , n54486 , n54487 , n54488 , n54489 , n54490 , n54491 , n54492 , n54493 , n54494 , 
 n54495 , n54496 , n54497 , n54498 , n54499 , n54500 , n54501 , n54502 , n54503 , n54504 , 
 n54505 , n54506 , n54507 , n54508 , n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , 
 n54515 , n54516 , n54517 , n54518 , n54519 , n54520 , n54521 , n54522 , n54523 , n54524 , 
 n54525 , n54526 , n54527 , n54528 , n54529 , n54530 , n54531 , n54532 , n54533 , n54534 , 
 n54535 , n54536 , n54537 , n54538 , n54539 , n54540 , n54541 , n54542 , n54543 , n54544 , 
 n54545 , n54546 , n54547 , n54548 , n54549 , n54550 , n54551 , n54552 , n54553 , n54554 , 
 n54555 , n54556 , n54557 , n54558 , n54559 , n54560 , n54561 , n54562 , n54563 , n54564 , 
 n54565 , n54566 , n54567 , n54568 , n54569 , n54570 , n54571 , n54572 , n54573 , n54574 , 
 n54575 , n54576 , n54577 , n54578 , n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , 
 n54585 , n54586 , n54587 , n54588 , n54589 , n54590 , n54591 , n54592 , n54593 , n54594 , 
 n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , n54601 , n54602 , n54603 , n54604 , 
 n54605 , n54606 , n54607 , n54608 , n54609 , n54610 , n54611 , n54612 , n54613 , n54614 , 
 n54615 , n54616 , n54617 , n54618 , n54619 , n54620 , n54621 , n54622 , n54623 , n54624 , 
 n54625 , n54626 , n54627 , n54628 , n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , 
 n54635 , n54636 , n54637 , n54638 , n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , 
 n54645 , n54646 , n54647 , n54648 , n54649 , n54650 , n54651 , n54652 , n54653 , n54654 , 
 n54655 , n54656 , n54657 , n54658 , n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , 
 n54665 , n54666 , n54667 , n54668 , n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , 
 n54675 , n54676 , n54677 , n54678 , n54679 , n54680 , n54681 , n54682 , n54683 , n54684 , 
 n54685 , n54686 , n54687 , n54688 , n54689 , n54690 , n54691 , n54692 , n54693 , n54694 , 
 n54695 , n54696 , n54697 , n54698 , n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , 
 n54705 , n54706 , n54707 , n54708 , n54709 , n54710 , n54711 , n54712 , n54713 , n54714 , 
 n54715 , n54716 , n54717 , n54718 , n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , 
 n54725 , n54726 , n54727 , n54728 , n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , 
 n54735 , n54736 , n54737 , n54738 , n54739 , n54740 , n54741 , n54742 , n54743 , n54744 , 
 n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , n54751 , n54752 , n54753 , n54754 , 
 n54755 , n54756 , n54757 , n54758 , n54759 , n54760 , n54761 , n54762 , n54763 , n54764 , 
 n54765 , n54766 , n54767 , n54768 , n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , 
 n54775 , n54776 , n54777 , n54778 , n54779 , n54780 , n54781 , n54782 , n54783 , n54784 , 
 n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , 
 n54795 , n54796 , n54797 , n54798 , n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , 
 n54805 , n54806 , n54807 , n54808 , n54809 , n54810 , n54811 , n54812 , n54813 , n54814 , 
 n54815 , n54816 , n54817 , n54818 , n54819 , n54820 , n54821 , n54822 , n54823 , n54824 , 
 n54825 , n54826 , n54827 , n54828 , n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , 
 n54835 , n54836 , n54837 , n54838 , n54839 , n54840 , n54841 , n54842 , n54843 , n54844 , 
 n54845 , n54846 , n54847 , n54848 , n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , 
 n54855 , n54856 , n54857 , n54858 , n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , 
 n54865 , n54866 , n54867 , n54868 , n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , 
 n54875 , n54876 , n54877 , n54878 , n54879 , n54880 , n54881 , n54882 , n54883 , n54884 , 
 n54885 , n54886 , n54887 , n54888 , n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , 
 n54895 , n54896 , n54897 , n54898 , n54899 , n54900 , n54901 , n54902 , n54903 , n54904 , 
 n54905 , n54906 , n54907 , n54908 , n54909 , n54910 , n54911 , n54912 , n54913 , n54914 , 
 n54915 , n54916 , n54917 , n54918 , n54919 , n54920 , n54921 , n54922 , n54923 , n54924 , 
 n54925 , n54926 , n54927 , n54928 , n54929 , n54930 , n54931 , n54932 , n54933 , n54934 , 
 n54935 , n54936 , n54937 , n54938 , n54939 , n54940 , n54941 , n54942 , n54943 , n54944 , 
 n54945 , n54946 , n54947 , n54948 , n54949 , n54950 , n54951 , n54952 , n54953 , n54954 , 
 n54955 , n54956 , n54957 , n54958 , n54959 , n54960 , n54961 , n54962 , n54963 , n54964 , 
 n54965 , n54966 , n54967 , n54968 , n54969 , n54970 , n54971 , n54972 , n54973 , n54974 , 
 n54975 , n54976 , n54977 , n54978 , n54979 , n54980 , n54981 , n54982 , n54983 , n54984 , 
 n54985 , n54986 , n54987 , n54988 , n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , 
 n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , n55001 , n55002 , n55003 , n55004 , 
 n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , n55011 , n55012 , n55013 , n55014 , 
 n55015 , n55016 , n55017 , n55018 , n55019 , n55020 , n55021 , n55022 , n55023 , n55024 , 
 n55025 , n55026 , n55027 , n55028 , n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , 
 n55035 , n55036 , n55037 , n55038 , n55039 , n55040 , n55041 , n55042 , n55043 , n55044 , 
 n55045 , n55046 , n55047 , n55048 , n55049 , n55050 , n55051 , n55052 , n55053 , n55054 , 
 n55055 , n55056 , n55057 , n55058 , n55059 , n55060 , n55061 , n55062 , n55063 , n55064 , 
 n55065 , n55066 , n55067 , n55068 , n55069 , n55070 , n55071 , n55072 , n55073 , n55074 , 
 n55075 , n55076 , n55077 , n55078 , n55079 , n55080 , n55081 , n55082 , n55083 , n55084 , 
 n55085 , n55086 , n55087 , n55088 , n55089 , n55090 , n55091 , n55092 , n55093 , n55094 , 
 n55095 , n55096 , n55097 , n55098 , n55099 , n55100 , n55101 , n55102 , n55103 , n55104 , 
 n55105 , n55106 , n55107 , n55108 , n55109 , n55110 , n55111 , n55112 , n55113 , n55114 , 
 n55115 , n55116 , n55117 , n55118 , n55119 , n55120 , n55121 , n55122 , n55123 , n55124 , 
 n55125 , n55126 , n55127 , n55128 , n55129 , n55130 , n55131 , n55132 , n55133 , n55134 , 
 n55135 , n55136 , n55137 , n55138 , n55139 , n55140 , n55141 , n55142 , n55143 , n55144 , 
 n55145 , n55146 , n55147 , n55148 , n55149 , n55150 , n55151 , n55152 , n55153 , n55154 , 
 n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , n55161 , n55162 , n55163 , n55164 , 
 n55165 , n55166 , n55167 , n55168 , n55169 , n55170 , n55171 , n55172 , n55173 , n55174 , 
 n55175 , n55176 , n55177 , n55178 , n55179 , n55180 , n55181 , n55182 , n55183 , n55184 , 
 n55185 , n55186 , n55187 , n55188 , n55189 , n55190 , n55191 , n55192 , n55193 , n55194 , 
 n55195 , n55196 , n55197 , n55198 , n55199 , n55200 , n55201 , n55202 , n55203 , n55204 , 
 n55205 , n55206 , n55207 , n55208 , n55209 , n55210 , n55211 , n55212 , n55213 , n55214 , 
 n55215 , n55216 , n55217 , n55218 , n55219 , n55220 , n55221 , n55222 , n55223 , n55224 , 
 n55225 , n55226 , n55227 , n55228 , n55229 , n55230 , n55231 , n55232 , n55233 , n55234 , 
 n55235 , n55236 , n55237 , n55238 , n55239 , n55240 , n55241 , n55242 , n55243 , n55244 , 
 n55245 , n55246 , n55247 , n55248 , n55249 , n55250 , n55251 , n55252 , n55253 , n55254 , 
 n55255 , n55256 , n55257 , n55258 , n55259 , n55260 , n55261 , n55262 , n55263 , n55264 , 
 n55265 , n55266 , n55267 , n55268 , n55269 , n55270 , n55271 , n55272 , n55273 , n55274 , 
 n55275 , n55276 , n55277 , n55278 , n55279 , n55280 , n55281 , n55282 , n55283 , n55284 , 
 n55285 , n55286 , n55287 , n55288 , n55289 , n55290 , n55291 , n55292 , n55293 , n55294 , 
 n55295 , n55296 , n55297 , n55298 , n55299 , n55300 , n55301 , n55302 , n55303 , n55304 , 
 n55305 , n55306 , n55307 , n55308 , n55309 , n55310 , n55311 , n55312 , n55313 , n55314 , 
 n55315 , n55316 , n55317 , n55318 , n55319 , n55320 , n55321 , n55322 , n55323 , n55324 , 
 n55325 , n55326 , n55327 , n55328 , n55329 , n55330 , n55331 , n55332 , n55333 , n55334 , 
 n55335 , n55336 , n55337 , n55338 , n55339 , n55340 , n55341 , n55342 , n55343 , n55344 , 
 n55345 , n55346 , n55347 , n55348 , n55349 , n55350 , n55351 , n55352 , n55353 , n55354 , 
 n55355 , n55356 , n55357 , n55358 , n55359 , n55360 , n55361 , n55362 , n55363 , n55364 , 
 n55365 , n55366 , n55367 , n55368 , n55369 , n55370 , n55371 , n55372 , n55373 , n55374 , 
 n55375 , n55376 , n55377 , n55378 , n55379 , n55380 , n55381 , n55382 , n55383 , n55384 , 
 n55385 , n55386 , n55387 , n55388 , n55389 , n55390 , n55391 , n55392 , n55393 , n55394 , 
 n55395 , n55396 , n55397 , n55398 , n55399 , n55400 , n55401 , n55402 , n55403 , n55404 , 
 n55405 , n55406 , n55407 , n55408 , n55409 , n55410 , n55411 , n55412 , n55413 , n55414 , 
 n55415 , n55416 , n55417 , n55418 , n55419 , n55420 , n55421 , n55422 , n55423 , n55424 , 
 n55425 , n55426 , n55427 , n55428 , n55429 , n55430 , n55431 , n55432 , n55433 , n55434 , 
 n55435 , n55436 , n55437 , n55438 , n55439 , n55440 , n55441 , n55442 , n55443 , n55444 , 
 n55445 , n55446 , n55447 , n55448 , n55449 , n55450 , n55451 , n55452 , n55453 , n55454 , 
 n55455 , n55456 , n55457 , n55458 , n55459 , n55460 , n55461 , n55462 , n55463 , n55464 , 
 n55465 , n55466 , n55467 , n55468 , n55469 , n55470 , n55471 , n55472 , n55473 , n55474 , 
 n55475 , n55476 , n55477 , n55478 , n55479 , n55480 , n55481 , n55482 , n55483 , n55484 , 
 n55485 , n55486 , n55487 , n55488 , n55489 , n55490 , n55491 , n55492 , n55493 , n55494 , 
 n55495 , n55496 , n55497 , n55498 , n55499 , n55500 , n55501 , n55502 , n55503 , n55504 , 
 n55505 , n55506 , n55507 , n55508 , n55509 , n55510 , n55511 , n55512 , n55513 , n55514 , 
 n55515 , n55516 , n55517 , n55518 , n55519 , n55520 , n55521 , n55522 , n55523 , n55524 , 
 n55525 , n55526 , n55527 , n55528 , n55529 , n55530 , n55531 , n55532 , n55533 , n55534 , 
 n55535 , n55536 , n55537 , n55538 , n55539 , n55540 , n55541 , n55542 , n55543 , n55544 , 
 n55545 , n55546 , n55547 , n55548 , n55549 , n55550 , n55551 , n55552 , n55553 , n55554 , 
 n55555 , n55556 , n55557 , n55558 , n55559 , n55560 , n55561 , n55562 , n55563 , n55564 , 
 n55565 , n55566 , n55567 , n55568 , n55569 , n55570 , n55571 , n55572 , n55573 , n55574 , 
 n55575 , n55576 , n55577 , n55578 , n55579 , n55580 , n55581 , n55582 , n55583 , n55584 , 
 n55585 , n55586 , n55587 , n55588 , n55589 , n55590 , n55591 , n55592 , n55593 , n55594 , 
 n55595 , n55596 , n55597 , n55598 , n55599 , n55600 , n55601 , n55602 , n55603 , n55604 , 
 n55605 , n55606 , n55607 , n55608 , n55609 , n55610 , n55611 , n55612 , n55613 , n55614 , 
 n55615 , n55616 , n55617 , n55618 , n55619 , n55620 , n55621 , n55622 , n55623 , n55624 , 
 n55625 , n55626 , n55627 , n55628 , n55629 , n55630 , n55631 , n55632 , n55633 , n55634 , 
 n55635 , n55636 , n55637 , n55638 , n55639 , n55640 , n55641 , n55642 , n55643 , n55644 , 
 n55645 , n55646 , n55647 , n55648 , n55649 , n55650 , n55651 , n55652 , n55653 , n55654 , 
 n55655 , n55656 , n55657 , n55658 , n55659 , n55660 , n55661 , n55662 , n55663 , n55664 , 
 n55665 , n55666 , n55667 , n55668 , n55669 , n55670 , n55671 , n55672 , n55673 , n55674 , 
 n55675 , n55676 , n55677 , n55678 , n55679 , n55680 , n55681 , n55682 , n55683 , n55684 , 
 n55685 , n55686 , n55687 , n55688 , n55689 , n55690 , n55691 , n55692 , n55693 , n55694 , 
 n55695 , n55696 , n55697 , n55698 , n55699 , n55700 , n55701 , n55702 , n55703 , n55704 , 
 n55705 , n55706 , n55707 , n55708 , n55709 , n55710 , n55711 , n55712 , n55713 , n55714 , 
 n55715 , n55716 , n55717 , n55718 , n55719 , n55720 , n55721 , n55722 , n55723 , n55724 , 
 n55725 , n55726 , n55727 , n55728 , n55729 , n55730 , n55731 , n55732 , n55733 , n55734 , 
 n55735 , n55736 , n55737 , n55738 , n55739 , n55740 , n55741 , n55742 , n55743 , n55744 , 
 n55745 , n55746 , n55747 , n55748 , n55749 , n55750 , n55751 , n55752 , n55753 , n55754 , 
 n55755 , n55756 , n55757 , n55758 , n55759 , n55760 , n55761 , n55762 , n55763 , n55764 , 
 n55765 , n55766 , n55767 , n55768 , n55769 , n55770 , n55771 , n55772 , n55773 , n55774 , 
 n55775 , n55776 , n55777 , n55778 , n55779 , n55780 , n55781 , n55782 , n55783 , n55784 , 
 n55785 , n55786 , n55787 , n55788 , n55789 , n55790 , n55791 , n55792 , n55793 , n55794 , 
 n55795 , n55796 , n55797 , n55798 , n55799 , n55800 , n55801 , n55802 , n55803 , n55804 , 
 n55805 , n55806 , n55807 , n55808 , n55809 , n55810 , n55811 , n55812 , n55813 , n55814 , 
 n55815 , n55816 , n55817 , n55818 , n55819 , n55820 , n55821 , n55822 , n55823 , n55824 , 
 n55825 , n55826 , n55827 , n55828 , n55829 , n55830 , n55831 , n55832 , n55833 , n55834 , 
 n55835 , n55836 , n55837 , n55838 , n55839 , n55840 , n55841 , n55842 , n55843 , n55844 , 
 n55845 , n55846 , n55847 , n55848 , n55849 , n55850 , n55851 , n55852 , n55853 , n55854 , 
 n55855 , n55856 , n55857 , n55858 , n55859 , n55860 , n55861 , n55862 , n55863 , n55864 , 
 n55865 , n55866 , n55867 , n55868 , n55869 , n55870 , n55871 , n55872 , n55873 , n55874 , 
 n55875 , n55876 , n55877 , n55878 , n55879 , n55880 , n55881 , n55882 , n55883 , n55884 , 
 n55885 , n55886 , n55887 , n55888 , n55889 , n55890 , n55891 , n55892 , n55893 , n55894 , 
 n55895 , n55896 , n55897 , n55898 , n55899 , n55900 , n55901 , n55902 , n55903 , n55904 , 
 n55905 , n55906 , n55907 , n55908 , n55909 , n55910 , n55911 , n55912 , n55913 , n55914 , 
 n55915 , n55916 , n55917 , n55918 , n55919 , n55920 , n55921 , n55922 , n55923 , n55924 , 
 n55925 , n55926 , n55927 , n55928 , n55929 , n55930 , n55931 , n55932 , n55933 , n55934 , 
 n55935 , n55936 , n55937 , n55938 , n55939 , n55940 , n55941 , n55942 , n55943 , n55944 , 
 n55945 , n55946 , n55947 , n55948 , n55949 , n55950 , n55951 , n55952 , n55953 , n55954 , 
 n55955 , n55956 , n55957 , n55958 , n55959 , n55960 , n55961 , n55962 , n55963 , n55964 , 
 n55965 , n55966 , n55967 , n55968 , n55969 , n55970 , n55971 , n55972 , n55973 , n55974 , 
 n55975 , n55976 , n55977 , n55978 , n55979 , n55980 , n55981 , n55982 , n55983 , n55984 , 
 n55985 , n55986 , n55987 , n55988 , n55989 , n55990 , n55991 , n55992 , n55993 , n55994 , 
 n55995 , n55996 , n55997 , n55998 , n55999 , n56000 , n56001 , n56002 , n56003 , n56004 , 
 n56005 , n56006 , n56007 , n56008 , n56009 , n56010 , n56011 , n56012 , n56013 , n56014 , 
 n56015 , n56016 , n56017 , n56018 , n56019 , n56020 , n56021 , n56022 , n56023 , n56024 , 
 n56025 , n56026 , n56027 , n56028 , n56029 , n56030 , n56031 , n56032 , n56033 , n56034 , 
 n56035 , n56036 , n56037 , n56038 , n56039 , n56040 , n56041 , n56042 , n56043 , n56044 , 
 n56045 , n56046 , n56047 , n56048 , n56049 , n56050 , n56051 , n56052 , n56053 , n56054 , 
 n56055 , n56056 , n56057 , n56058 , n56059 , n56060 , n56061 , n56062 , n56063 , n56064 , 
 n56065 , n56066 , n56067 , n56068 , n56069 , n56070 , n56071 , n56072 , n56073 , n56074 , 
 n56075 , n56076 , n56077 , n56078 , n56079 , n56080 , n56081 , n56082 , n56083 , n56084 , 
 n56085 , n56086 , n56087 , n56088 , n56089 , n56090 , n56091 , n56092 , n56093 , n56094 , 
 n56095 , n56096 , n56097 , n56098 , n56099 , n56100 , n56101 , n56102 , n56103 , n56104 , 
 n56105 , n56106 , n56107 , n56108 , n56109 , n56110 , n56111 , n56112 , n56113 , n56114 , 
 n56115 , n56116 , n56117 , n56118 , n56119 , n56120 , n56121 , n56122 , n56123 , n56124 , 
 n56125 , n56126 , n56127 , n56128 , n56129 , n56130 , n56131 , n56132 , n56133 , n56134 , 
 n56135 , n56136 , n56137 , n56138 , n56139 , n56140 , n56141 , n56142 , n56143 , n56144 , 
 n56145 , n56146 , n56147 , n56148 , n56149 , n56150 , n56151 , n56152 , n56153 , n56154 , 
 n56155 , n56156 , n56157 , n56158 , n56159 , n56160 , n56161 , n56162 , n56163 , n56164 , 
 n56165 , n56166 , n56167 , n56168 , n56169 , n56170 , n56171 , n56172 , n56173 , n56174 , 
 n56175 , n56176 , n56177 , n56178 , n56179 , n56180 , n56181 , n56182 , n56183 , n56184 , 
 n56185 , n56186 , n56187 , n56188 , n56189 , n56190 , n56191 , n56192 , n56193 , n56194 , 
 n56195 , n56196 , n56197 , n56198 , n56199 , n56200 , n56201 , n56202 , n56203 , n56204 , 
 n56205 , n56206 , n56207 , n56208 , n56209 , n56210 , n56211 , n56212 , n56213 , n56214 , 
 n56215 , n56216 , n56217 , n56218 , n56219 , n56220 , n56221 , n56222 , n56223 , n56224 , 
 n56225 , n56226 , n56227 , n56228 , n56229 , n56230 , n56231 , n56232 , n56233 , n56234 , 
 n56235 , n56236 , n56237 , n56238 , n56239 , n56240 , n56241 , n56242 , n56243 , n56244 , 
 n56245 , n56246 , n56247 , n56248 , n56249 , n56250 , n56251 , n56252 , n56253 , n56254 , 
 n56255 , n56256 , n56257 , n56258 , n56259 , n56260 , n56261 , n56262 , n56263 , n56264 , 
 n56265 , n56266 , n56267 , n56268 , n56269 , n56270 , n56271 , n56272 , n56273 , n56274 , 
 n56275 , n56276 , n56277 , n56278 , n56279 , n56280 , n56281 , n56282 , n56283 , n56284 , 
 n56285 , n56286 , n56287 , n56288 , n56289 , n56290 , n56291 , n56292 , n56293 , n56294 , 
 n56295 , n56296 , n56297 , n56298 , n56299 , n56300 , n56301 , n56302 , n56303 , n56304 , 
 n56305 , n56306 , n56307 , n56308 , n56309 , n56310 , n56311 , n56312 , n56313 , n56314 , 
 n56315 , n56316 , n56317 , n56318 , n56319 , n56320 , n56321 , n56322 , n56323 , n56324 , 
 n56325 , n56326 , n56327 , n56328 , n56329 , n56330 , n56331 , n56332 , n56333 , n56334 , 
 n56335 , n56336 , n56337 , n56338 , n56339 , n56340 , n56341 , n56342 , n56343 , n56344 , 
 n56345 , n56346 , n56347 , n56348 , n56349 , n56350 , n56351 , n56352 , n56353 , n56354 , 
 n56355 , n56356 , n56357 , n56358 , n56359 , n56360 , n56361 , n56362 , n56363 , n56364 , 
 n56365 , n56366 , n56367 , n56368 , n56369 , n56370 , n56371 , n56372 , n56373 , n56374 , 
 n56375 , n56376 , n56377 , n56378 , n56379 , n56380 , n56381 , n56382 , n56383 , n56384 , 
 n56385 , n56386 , n56387 , n56388 , n56389 , n56390 , n56391 , n56392 , n56393 , n56394 , 
 n56395 , n56396 , n56397 , n56398 , n56399 , n56400 , n56401 , n56402 , n56403 , n56404 , 
 n56405 , n56406 , n56407 , n56408 , n56409 , n56410 , n56411 , n56412 , n56413 , n56414 , 
 n56415 , n56416 , n56417 , n56418 , n56419 , n56420 , n56421 , n56422 , n56423 , n56424 , 
 n56425 , n56426 , n56427 , n56428 , n56429 , n56430 , n56431 , n56432 , n56433 , n56434 , 
 n56435 , n56436 , n56437 , n56438 , n56439 , n56440 , n56441 , n56442 , n56443 , n56444 , 
 n56445 , n56446 , n56447 , n56448 , n56449 , n56450 , n56451 , n56452 , n56453 , n56454 , 
 n56455 , n56456 , n56457 , n56458 , n56459 , n56460 , n56461 , n56462 , n56463 , n56464 , 
 n56465 , n56466 , n56467 , n56468 , n56469 , n56470 , n56471 , n56472 , n56473 , n56474 , 
 n56475 , n56476 , n56477 , n56478 , n56479 , n56480 , n56481 , n56482 , n56483 , n56484 , 
 n56485 , n56486 , n56487 , n56488 , n56489 , n56490 , n56491 , n56492 , n56493 , n56494 , 
 n56495 , n56496 , n56497 , n56498 , n56499 , n56500 , n56501 , n56502 , n56503 , n56504 , 
 n56505 , n56506 , n56507 , n56508 , n56509 , n56510 , n56511 , n56512 , n56513 , n56514 , 
 n56515 , n56516 , n56517 , n56518 , n56519 , n56520 , n56521 , n56522 , n56523 , n56524 , 
 n56525 , n56526 , n56527 , n56528 , n56529 , n56530 , n56531 , n56532 , n56533 , n56534 , 
 n56535 , n56536 , n56537 , n56538 , n56539 , n56540 , n56541 , n56542 , n56543 , n56544 , 
 n56545 , n56546 , n56547 , n56548 , n56549 , n56550 , n56551 , n56552 , n56553 , n56554 , 
 n56555 , n56556 , n56557 , n56558 , n56559 , n56560 , n56561 , n56562 , n56563 , n56564 , 
 n56565 , n56566 , n56567 , n56568 , n56569 , n56570 , n56571 , n56572 , n56573 , n56574 , 
 n56575 , n56576 , n56577 , n56578 , n56579 , n56580 , n56581 , n56582 , n56583 , n56584 , 
 n56585 , n56586 , n56587 , n56588 , n56589 , n56590 , n56591 , n56592 , n56593 , n56594 , 
 n56595 , n56596 , n56597 , n56598 , n56599 , n56600 , n56601 , n56602 , n56603 , n56604 , 
 n56605 , n56606 , n56607 , n56608 , n56609 , n56610 , n56611 , n56612 , n56613 , n56614 , 
 n56615 , n56616 , n56617 , n56618 , n56619 , n56620 , n56621 , n56622 , n56623 , n56624 , 
 n56625 , n56626 , n56627 , n56628 , n56629 , n56630 , n56631 , n56632 , n56633 , n56634 , 
 n56635 , n56636 , n56637 , n56638 , n56639 , n56640 , n56641 , n56642 , n56643 , n56644 , 
 n56645 , n56646 , n56647 , n56648 , n56649 , n56650 , n56651 , n56652 , n56653 , n56654 , 
 n56655 , n56656 , n56657 , n56658 , n56659 , n56660 , n56661 , n56662 , n56663 , n56664 , 
 n56665 , n56666 , n56667 , n56668 , n56669 , n56670 , n56671 , n56672 , n56673 , n56674 , 
 n56675 , n56676 , n56677 , n56678 , n56679 , n56680 , n56681 , n56682 , n56683 , n56684 , 
 n56685 , n56686 , n56687 , n56688 , n56689 , n56690 , n56691 , n56692 , n56693 , n56694 , 
 n56695 , n56696 , n56697 , n56698 , n56699 , n56700 , n56701 , n56702 , n56703 , n56704 , 
 n56705 , n56706 , n56707 , n56708 , n56709 , n56710 , n56711 , n56712 , n56713 , n56714 , 
 n56715 , n56716 , n56717 , n56718 , n56719 , n56720 , n56721 , n56722 , n56723 , n56724 , 
 n56725 , n56726 , n56727 , n56728 , n56729 , n56730 , n56731 , n56732 , n56733 , n56734 , 
 n56735 , n56736 , n56737 , n56738 , n56739 , n56740 , n56741 , n56742 , n56743 , n56744 , 
 n56745 , n56746 , n56747 , n56748 , n56749 , n56750 , n56751 , n56752 , n56753 , n56754 , 
 n56755 , n56756 , n56757 , n56758 , n56759 , n56760 , n56761 , n56762 , n56763 , n56764 , 
 n56765 , n56766 , n56767 , n56768 , n56769 , n56770 , n56771 , n56772 , n56773 , n56774 , 
 n56775 , n56776 , n56777 , n56778 , n56779 , n56780 , n56781 , n56782 , n56783 , n56784 , 
 n56785 , n56786 , n56787 , n56788 , n56789 , n56790 , n56791 , n56792 , n56793 , n56794 , 
 n56795 , n56796 , n56797 , n56798 , n56799 , n56800 , n56801 , n56802 , n56803 , n56804 , 
 n56805 , n56806 , n56807 , n56808 , n56809 , n56810 , n56811 , n56812 , n56813 , n56814 , 
 n56815 , n56816 , n56817 , n56818 , n56819 , n56820 , n56821 , n56822 , n56823 , n56824 , 
 n56825 , n56826 , n56827 , n56828 , n56829 , n56830 , n56831 , n56832 , n56833 , n56834 , 
 n56835 , n56836 , n56837 , n56838 , n56839 , n56840 , n56841 , n56842 , n56843 , n56844 , 
 n56845 , n56846 , n56847 , n56848 , n56849 , n56850 , n56851 , n56852 , n56853 , n56854 , 
 n56855 , n56856 , n56857 , n56858 , n56859 , n56860 , n56861 , n56862 , n56863 , n56864 , 
 n56865 , n56866 , n56867 , n56868 , n56869 , n56870 , n56871 , n56872 , n56873 , n56874 , 
 n56875 , n56876 , n56877 , n56878 , n56879 , n56880 , n56881 , n56882 , n56883 , n56884 , 
 n56885 , n56886 , n56887 , n56888 , n56889 , n56890 , n56891 , n56892 , n56893 , n56894 , 
 n56895 , n56896 , n56897 , n56898 , n56899 , n56900 , n56901 , n56902 , n56903 , n56904 , 
 n56905 , n56906 , n56907 , n56908 , n56909 , n56910 , n56911 , n56912 , n56913 , n56914 , 
 n56915 , n56916 , n56917 , n56918 , n56919 , n56920 , n56921 , n56922 , n56923 , n56924 , 
 n56925 , n56926 , n56927 , n56928 , n56929 , n56930 , n56931 , n56932 , n56933 , n56934 , 
 n56935 , n56936 , n56937 , n56938 , n56939 , n56940 , n56941 , n56942 , n56943 , n56944 , 
 n56945 , n56946 , n56947 , n56948 , n56949 , n56950 , n56951 , n56952 , n56953 , n56954 , 
 n56955 , n56956 , n56957 , n56958 , n56959 , n56960 , n56961 , n56962 , n56963 , n56964 , 
 n56965 , n56966 , n56967 , n56968 , n56969 , n56970 , n56971 , n56972 , n56973 , n56974 , 
 n56975 , n56976 , n56977 , n56978 , n56979 , n56980 , n56981 , n56982 , n56983 , n56984 , 
 n56985 , n56986 , n56987 , n56988 , n56989 , n56990 , n56991 , n56992 , n56993 , n56994 , 
 n56995 , n56996 , n56997 , n56998 , n56999 , n57000 , n57001 , n57002 , n57003 , n57004 , 
 n57005 , n57006 , n57007 , n57008 , n57009 , n57010 , n57011 , n57012 , n57013 , n57014 , 
 n57015 , n57016 , n57017 , n57018 , n57019 , n57020 , n57021 , n57022 , n57023 , n57024 , 
 n57025 , n57026 , n57027 , n57028 , n57029 , n57030 , n57031 , n57032 , n57033 , n57034 , 
 n57035 , n57036 , n57037 , n57038 , n57039 , n57040 , n57041 , n57042 , n57043 , n57044 , 
 n57045 , n57046 , n57047 , n57048 , n57049 , n57050 , n57051 , n57052 , n57053 , n57054 , 
 n57055 , n57056 , n57057 , n57058 , n57059 , n57060 , n57061 , n57062 , n57063 , n57064 , 
 n57065 , n57066 , n57067 , n57068 , n57069 , n57070 , n57071 , n57072 , n57073 , n57074 , 
 n57075 , n57076 , n57077 , n57078 , n57079 , n57080 , n57081 , n57082 , n57083 , n57084 , 
 n57085 , n57086 , n57087 , n57088 , n57089 , n57090 , n57091 , n57092 , n57093 , n57094 , 
 n57095 , n57096 , n57097 , n57098 , n57099 , n57100 , n57101 , n57102 , n57103 , n57104 , 
 n57105 , n57106 , n57107 , n57108 , n57109 , n57110 , n57111 , n57112 , n57113 , n57114 , 
 n57115 , n57116 , n57117 , n57118 , n57119 , n57120 , n57121 , n57122 , n57123 , n57124 , 
 n57125 , n57126 , n57127 , n57128 , n57129 , n57130 , n57131 , n57132 , n57133 , n57134 , 
 n57135 , n57136 , n57137 , n57138 , n57139 , n57140 , n57141 , n57142 , n57143 , n57144 , 
 n57145 , n57146 , n57147 , n57148 , n57149 , n57150 , n57151 , n57152 , n57153 , n57154 , 
 n57155 , n57156 , n57157 , n57158 , n57159 , n57160 , n57161 , n57162 , n57163 , n57164 , 
 n57165 , n57166 , n57167 , n57168 , n57169 , n57170 , n57171 , n57172 , n57173 , n57174 , 
 n57175 , n57176 , n57177 , n57178 , n57179 , n57180 , n57181 , n57182 , n57183 , n57184 , 
 n57185 , n57186 , n57187 , n57188 , n57189 , n57190 , n57191 , n57192 , n57193 , n57194 , 
 n57195 , n57196 , n57197 , n57198 , n57199 , n57200 , n57201 , n57202 , n57203 , n57204 , 
 n57205 , n57206 , n57207 , n57208 , n57209 , n57210 , n57211 , n57212 , n57213 , n57214 , 
 n57215 , n57216 , n57217 , n57218 , n57219 , n57220 , n57221 , n57222 , n57223 , n57224 , 
 n57225 , n57226 , n57227 , n57228 , n57229 , n57230 , n57231 , n57232 , n57233 , n57234 , 
 n57235 , n57236 , n57237 , n57238 , n57239 , n57240 , n57241 , n57242 , n57243 , n57244 , 
 n57245 , n57246 , n57247 , n57248 , n57249 , n57250 , n57251 , n57252 , n57253 , n57254 , 
 n57255 , n57256 , n57257 , n57258 , n57259 , n57260 , n57261 , n57262 , n57263 , n57264 , 
 n57265 , n57266 , n57267 , n57268 , n57269 , n57270 , n57271 , n57272 , n57273 , n57274 , 
 n57275 , n57276 , n57277 , n57278 , n57279 , n57280 , n57281 , n57282 , n57283 , n57284 , 
 n57285 , n57286 , n57287 , n57288 , n57289 , n57290 , n57291 , n57292 , n57293 , n57294 , 
 n57295 , n57296 , n57297 , n57298 , n57299 , n57300 , n57301 , n57302 , n57303 , n57304 , 
 n57305 , n57306 , n57307 , n57308 , n57309 , n57310 , n57311 , n57312 , n57313 , n57314 , 
 n57315 , n57316 , n57317 , n57318 , n57319 , n57320 , n57321 , n57322 , n57323 , n57324 , 
 n57325 , n57326 , n57327 , n57328 , n57329 , n57330 , n57331 , n57332 , n57333 , n57334 , 
 n57335 , n57336 , n57337 , n57338 , n57339 , n57340 , n57341 , n57342 , n57343 , n57344 , 
 n57345 , n57346 , n57347 , n57348 , n57349 , n57350 , n57351 , n57352 , n57353 , n57354 , 
 n57355 , n57356 , n57357 , n57358 , n57359 , n57360 , n57361 , n57362 , n57363 , n57364 , 
 n57365 , n57366 , n57367 , n57368 , n57369 , n57370 , n57371 , n57372 , n57373 , n57374 , 
 n57375 , n57376 , n57377 , n57378 , n57379 , n57380 , n57381 , n57382 , n57383 , n57384 , 
 n57385 , n57386 , n57387 , n57388 , n57389 , n57390 , n57391 , n57392 , n57393 , n57394 , 
 n57395 , n57396 , n57397 , n57398 , n57399 , n57400 , n57401 , n57402 , n57403 , n57404 , 
 n57405 , n57406 , n57407 , n57408 , n57409 , n57410 , n57411 , n57412 , n57413 , n57414 , 
 n57415 , n57416 , n57417 , n57418 , n57419 , n57420 , n57421 , n57422 , n57423 , n57424 , 
 n57425 , n57426 , n57427 , n57428 , n57429 , n57430 , n57431 , n57432 , n57433 , n57434 , 
 n57435 , n57436 , n57437 , n57438 , n57439 , n57440 , n57441 , n57442 , n57443 , n57444 , 
 n57445 , n57446 , n57447 , n57448 , n57449 , n57450 , n57451 , n57452 , n57453 , n57454 , 
 n57455 , n57456 , n57457 , n57458 , n57459 , n57460 , n57461 , n57462 , n57463 , n57464 , 
 n57465 , n57466 , n57467 , n57468 , n57469 , n57470 , n57471 , n57472 , n57473 , n57474 , 
 n57475 , n57476 , n57477 , n57478 , n57479 , n57480 , n57481 , n57482 , n57483 , n57484 , 
 n57485 , n57486 , n57487 , n57488 , n57489 , n57490 , n57491 , n57492 , n57493 , n57494 , 
 n57495 , n57496 , n57497 , n57498 , n57499 , n57500 , n57501 , n57502 , n57503 , n57504 , 
 n57505 , n57506 , n57507 , n57508 , n57509 , n57510 , n57511 , n57512 , n57513 , n57514 , 
 n57515 , n57516 , n57517 , n57518 , n57519 , n57520 , n57521 , n57522 , n57523 , n57524 , 
 n57525 , n57526 , n57527 , n57528 , n57529 , n57530 , n57531 , n57532 , n57533 , n57534 , 
 n57535 , n57536 , n57537 , n57538 , n57539 , n57540 , n57541 , n57542 , n57543 , n57544 , 
 n57545 , n57546 , n57547 , n57548 , n57549 , n57550 , n57551 , n57552 , n57553 , n57554 , 
 n57555 , n57556 , n57557 , n57558 , n57559 , n57560 , n57561 , n57562 , n57563 , n57564 , 
 n57565 , n57566 , n57567 , n57568 , n57569 , n57570 , n57571 , n57572 , n57573 , n57574 , 
 n57575 , n57576 , n57577 , n57578 , n57579 , n57580 , n57581 , n57582 , n57583 , n57584 , 
 n57585 , n57586 , n57587 , n57588 , n57589 , n57590 , n57591 , n57592 , n57593 , n57594 , 
 n57595 , n57596 , n57597 , n57598 , n57599 , n57600 , n57601 , n57602 , n57603 , n57604 , 
 n57605 , n57606 , n57607 , n57608 , n57609 , n57610 , n57611 , n57612 , n57613 , n57614 , 
 n57615 , n57616 , n57617 , n57618 , n57619 , n57620 , n57621 , n57622 , n57623 , n57624 , 
 n57625 , n57626 , n57627 , n57628 , n57629 , n57630 , n57631 , n57632 , n57633 , n57634 , 
 n57635 , n57636 , n57637 , n57638 , n57639 , n57640 , n57641 , n57642 , n57643 , n57644 , 
 n57645 , n57646 , n57647 , n57648 , n57649 , n57650 , n57651 , n57652 , n57653 , n57654 , 
 n57655 , n57656 , n57657 , n57658 , n57659 , n57660 , n57661 , n57662 , n57663 , n57664 , 
 n57665 , n57666 , n57667 , n57668 , n57669 , n57670 , n57671 , n57672 , n57673 , n57674 , 
 n57675 , n57676 , n57677 , n57678 , n57679 , n57680 , n57681 , n57682 , n57683 , n57684 , 
 n57685 , n57686 , n57687 , n57688 , n57689 , n57690 , n57691 , n57692 , n57693 , n57694 , 
 n57695 , n57696 , n57697 , n57698 , n57699 , n57700 , n57701 , n57702 , n57703 , n57704 , 
 n57705 , n57706 , n57707 , n57708 , n57709 , n57710 , n57711 , n57712 , n57713 , n57714 , 
 n57715 , n57716 , n57717 , n57718 , n57719 , n57720 , n57721 , n57722 , n57723 , n57724 , 
 n57725 , n57726 , n57727 , n57728 , n57729 , n57730 , n57731 , n57732 , n57733 , n57734 , 
 n57735 , n57736 , n57737 , n57738 , n57739 , n57740 , n57741 , n57742 , n57743 , n57744 , 
 n57745 , n57746 , n57747 , n57748 , n57749 , n57750 , n57751 , n57752 , n57753 , n57754 , 
 n57755 , n57756 , n57757 , n57758 , n57759 , n57760 , n57761 , n57762 , n57763 , n57764 , 
 n57765 , n57766 , n57767 , n57768 , n57769 , n57770 , n57771 , n57772 , n57773 , n57774 , 
 n57775 , n57776 , n57777 , n57778 , n57779 , n57780 , n57781 , n57782 , n57783 , n57784 , 
 n57785 , n57786 , n57787 , n57788 , n57789 , n57790 , n57791 , n57792 , n57793 , n57794 , 
 n57795 , n57796 , n57797 , n57798 , n57799 , n57800 , n57801 , n57802 , n57803 , n57804 , 
 n57805 , n57806 , n57807 , n57808 , n57809 , n57810 , n57811 , n57812 , n57813 , n57814 , 
 n57815 , n57816 , n57817 , n57818 , n57819 , n57820 , n57821 , n57822 , n57823 , n57824 , 
 n57825 , n57826 , n57827 , n57828 , n57829 , n57830 , n57831 , n57832 , n57833 , n57834 , 
 n57835 , n57836 , n57837 , n57838 , n57839 , n57840 , n57841 , n57842 , n57843 , n57844 , 
 n57845 , n57846 , n57847 , n57848 , n57849 , n57850 , n57851 , n57852 , n57853 , n57854 , 
 n57855 , n57856 , n57857 , n57858 , n57859 , n57860 , n57861 , n57862 , n57863 , n57864 , 
 n57865 , n57866 , n57867 , n57868 , n57869 , n57870 , n57871 , n57872 , n57873 , n57874 , 
 n57875 , n57876 , n57877 , n57878 , n57879 , n57880 , n57881 , n57882 , n57883 , n57884 , 
 n57885 , n57886 , n57887 , n57888 , n57889 , n57890 , n57891 , n57892 , n57893 , n57894 , 
 n57895 , n57896 , n57897 , n57898 , n57899 , n57900 , n57901 , n57902 , n57903 , n57904 , 
 n57905 , n57906 , n57907 , n57908 , n57909 , n57910 , n57911 , n57912 , n57913 , n57914 , 
 n57915 , n57916 , n57917 , n57918 , n57919 , n57920 , n57921 , n57922 , n57923 , n57924 , 
 n57925 , n57926 , n57927 , n57928 , n57929 , n57930 , n57931 , n57932 , n57933 , n57934 , 
 n57935 , n57936 , n57937 , n57938 , n57939 , n57940 , n57941 , n57942 , n57943 , n57944 , 
 n57945 , n57946 , n57947 , n57948 , n57949 , n57950 , n57951 , n57952 , n57953 , n57954 , 
 n57955 , n57956 , n57957 , n57958 , n57959 , n57960 , n57961 , n57962 , n57963 , n57964 , 
 n57965 , n57966 , n57967 , n57968 , n57969 , n57970 , n57971 , n57972 , n57973 , n57974 , 
 n57975 , n57976 , n57977 , n57978 , n57979 , n57980 , n57981 , n57982 , n57983 , n57984 , 
 n57985 , n57986 , n57987 , n57988 , n57989 , n57990 , n57991 , n57992 , n57993 , n57994 , 
 n57995 , n57996 , n57997 , n57998 , n57999 , n58000 , n58001 , n58002 , n58003 , n58004 , 
 n58005 , n58006 , n58007 , n58008 , n58009 , n58010 , n58011 , n58012 , n58013 , n58014 , 
 n58015 , n58016 , n58017 , n58018 , n58019 , n58020 , n58021 , n58022 , n58023 , n58024 , 
 n58025 , n58026 , n58027 , n58028 , n58029 , n58030 , n58031 , n58032 , n58033 , n58034 , 
 n58035 , n58036 , n58037 , n58038 , n58039 , n58040 , n58041 , n58042 , n58043 , n58044 , 
 n58045 , n58046 , n58047 , n58048 , n58049 , n58050 , n58051 , n58052 , n58053 , n58054 , 
 n58055 , n58056 , n58057 , n58058 , n58059 , n58060 , n58061 , n58062 , n58063 , n58064 , 
 n58065 , n58066 , n58067 , n58068 , n58069 , n58070 , n58071 , n58072 , n58073 , n58074 , 
 n58075 , n58076 , n58077 , n58078 , n58079 , n58080 , n58081 , n58082 , n58083 , n58084 , 
 n58085 , n58086 , n58087 , n58088 , n58089 , n58090 , n58091 , n58092 , n58093 , n58094 , 
 n58095 , n58096 , n58097 , n58098 , n58099 , n58100 , n58101 , n58102 , n58103 , n58104 , 
 n58105 , n58106 , n58107 , n58108 , n58109 , n58110 , n58111 , n58112 , n58113 , n58114 , 
 n58115 , n58116 , n58117 , n58118 , n58119 , n58120 , n58121 , n58122 , n58123 , n58124 , 
 n58125 , n58126 , n58127 , n58128 , n58129 , n58130 , n58131 , n58132 , n58133 , n58134 , 
 n58135 , n58136 , n58137 , n58138 , n58139 , n58140 , n58141 , n58142 , n58143 , n58144 , 
 n58145 , n58146 , n58147 , n58148 , n58149 , n58150 , n58151 , n58152 , n58153 , n58154 , 
 n58155 , n58156 , n58157 , n58158 , n58159 , n58160 , n58161 , n58162 , n58163 , n58164 , 
 n58165 , n58166 , n58167 , n58168 , n58169 , n58170 , n58171 , n58172 , n58173 , n58174 , 
 n58175 , n58176 , n58177 , n58178 , n58179 , n58180 , n58181 , n58182 , n58183 , n58184 , 
 n58185 , n58186 , n58187 , n58188 , n58189 , n58190 , n58191 , n58192 , n58193 , n58194 , 
 n58195 , n58196 , n58197 , n58198 , n58199 , n58200 , n58201 , n58202 , n58203 , n58204 , 
 n58205 , n58206 , n58207 , n58208 , n58209 , n58210 , n58211 , n58212 , n58213 , n58214 , 
 n58215 , n58216 , n58217 , n58218 , n58219 , n58220 , n58221 , n58222 , n58223 , n58224 , 
 n58225 , n58226 , n58227 , n58228 , n58229 , n58230 , n58231 , n58232 , n58233 , n58234 , 
 n58235 , n58236 , n58237 , n58238 , n58239 , n58240 , n58241 , n58242 , n58243 , n58244 , 
 n58245 , n58246 , n58247 , n58248 , n58249 , n58250 , n58251 , n58252 , n58253 , n58254 , 
 n58255 , n58256 , n58257 , n58258 , n58259 , n58260 , n58261 , n58262 , n58263 , n58264 , 
 n58265 , n58266 , n58267 , n58268 , n58269 , n58270 , n58271 , n58272 , n58273 , n58274 , 
 n58275 , n58276 , n58277 , n58278 , n58279 , n58280 , n58281 , n58282 , n58283 , n58284 , 
 n58285 , n58286 , n58287 , n58288 , n58289 , n58290 , n58291 , n58292 , n58293 , n58294 , 
 n58295 , n58296 , n58297 , n58298 , n58299 , n58300 , n58301 , n58302 , n58303 , n58304 , 
 n58305 , n58306 , n58307 , n58308 , n58309 , n58310 , n58311 , n58312 , n58313 , n58314 , 
 n58315 , n58316 , n58317 , n58318 , n58319 , n58320 , n58321 , n58322 , n58323 , n58324 , 
 n58325 , n58326 , n58327 , n58328 , n58329 , n58330 , n58331 , n58332 , n58333 , n58334 , 
 n58335 , n58336 , n58337 , n58338 , n58339 , n58340 , n58341 , n58342 , n58343 , n58344 , 
 n58345 , n58346 , n58347 , n58348 , n58349 , n58350 , n58351 , n58352 , n58353 , n58354 , 
 n58355 , n58356 , n58357 , n58358 , n58359 , n58360 , n58361 , n58362 , n58363 , n58364 , 
 n58365 , n58366 , n58367 , n58368 , n58369 , n58370 , n58371 , n58372 , n58373 , n58374 , 
 n58375 , n58376 , n58377 , n58378 , n58379 , n58380 , n58381 , n58382 , n58383 , n58384 , 
 n58385 , n58386 , n58387 , n58388 , n58389 , n58390 , n58391 , n58392 , n58393 , n58394 , 
 n58395 , n58396 , n58397 , n58398 , n58399 , n58400 , n58401 , n58402 , n58403 , n58404 , 
 n58405 , n58406 , n58407 , n58408 , n58409 , n58410 , n58411 , n58412 , n58413 , n58414 , 
 n58415 , n58416 , n58417 , n58418 , n58419 , n58420 , n58421 , n58422 , n58423 , n58424 , 
 n58425 , n58426 , n58427 , n58428 , n58429 , n58430 , n58431 , n58432 , n58433 , n58434 , 
 n58435 , n58436 , n58437 , n58438 , n58439 , n58440 , n58441 , n58442 , n58443 , n58444 , 
 n58445 , n58446 , n58447 , n58448 , n58449 , n58450 , n58451 , n58452 , n58453 , n58454 , 
 n58455 , n58456 , n58457 , n58458 , n58459 , n58460 , n58461 , n58462 , n58463 , n58464 , 
 n58465 , n58466 , n58467 , n58468 , n58469 , n58470 , n58471 , n58472 , n58473 , n58474 , 
 n58475 , n58476 , n58477 , n58478 , n58479 , n58480 , n58481 , n58482 , n58483 , n58484 , 
 n58485 , n58486 , n58487 , n58488 , n58489 , n58490 , n58491 , n58492 , n58493 , n58494 , 
 n58495 , n58496 , n58497 , n58498 , n58499 , n58500 , n58501 , n58502 , n58503 , n58504 , 
 n58505 , n58506 , n58507 , n58508 , n58509 , n58510 , n58511 , n58512 , n58513 , n58514 , 
 n58515 , n58516 , n58517 , n58518 , n58519 , n58520 , n58521 , n58522 , n58523 , n58524 , 
 n58525 , n58526 , n58527 , n58528 , n58529 , n58530 , n58531 , n58532 , n58533 , n58534 , 
 n58535 , n58536 , n58537 , n58538 , n58539 , n58540 , n58541 , n58542 , n58543 , n58544 , 
 n58545 , n58546 , n58547 , n58548 , n58549 , n58550 , n58551 , n58552 , n58553 , n58554 , 
 n58555 , n58556 , n58557 , n58558 , n58559 , n58560 , n58561 , n58562 , n58563 , n58564 , 
 n58565 , n58566 , n58567 , n58568 , n58569 , n58570 , n58571 , n58572 , n58573 , n58574 , 
 n58575 , n58576 , n58577 , n58578 , n58579 , n58580 , n58581 , n58582 , n58583 , n58584 , 
 n58585 , n58586 , n58587 , n58588 , n58589 , n58590 , n58591 , n58592 , n58593 , n58594 , 
 n58595 , n58596 , n58597 , n58598 , n58599 , n58600 , n58601 , n58602 , n58603 , n58604 , 
 n58605 , n58606 , n58607 , n58608 , n58609 , n58610 , n58611 , n58612 , n58613 , n58614 , 
 n58615 , n58616 , n58617 , n58618 , n58619 , n58620 , n58621 , n58622 , n58623 , n58624 , 
 n58625 , n58626 , n58627 , n58628 , n58629 , n58630 , n58631 , n58632 , n58633 , n58634 , 
 n58635 , n58636 , n58637 , n58638 , n58639 , n58640 , n58641 , n58642 , n58643 , n58644 , 
 n58645 , n58646 , n58647 , n58648 , n58649 , n58650 , n58651 , n58652 , n58653 , n58654 , 
 n58655 , n58656 , n58657 , n58658 , n58659 , n58660 , n58661 , n58662 , n58663 , n58664 , 
 n58665 , n58666 , n58667 , n58668 , n58669 , n58670 , n58671 , n58672 , n58673 , n58674 , 
 n58675 , n58676 , n58677 , n58678 , n58679 , n58680 , n58681 , n58682 , n58683 , n58684 , 
 n58685 , n58686 , n58687 , n58688 , n58689 , n58690 , n58691 , n58692 , n58693 , n58694 , 
 n58695 , n58696 , n58697 , n58698 , n58699 , n58700 , n58701 , n58702 , n58703 , n58704 , 
 n58705 , n58706 , n58707 , n58708 , n58709 , n58710 , n58711 , n58712 , n58713 , n58714 , 
 n58715 , n58716 , n58717 , n58718 , n58719 , n58720 , n58721 , n58722 , n58723 , n58724 , 
 n58725 , n58726 , n58727 , n58728 , n58729 , n58730 , n58731 , n58732 , n58733 , n58734 , 
 n58735 , n58736 , n58737 , n58738 , n58739 , n58740 , n58741 , n58742 , n58743 , n58744 , 
 n58745 , n58746 , n58747 , n58748 , n58749 , n58750 , n58751 , n58752 , n58753 , n58754 , 
 n58755 , n58756 , n58757 , n58758 , n58759 , n58760 , n58761 , n58762 , n58763 , n58764 , 
 n58765 , n58766 , n58767 , n58768 , n58769 , n58770 , n58771 , n58772 , n58773 , n58774 , 
 n58775 , n58776 , n58777 , n58778 , n58779 , n58780 , n58781 , n58782 , n58783 , n58784 , 
 n58785 , n58786 , n58787 , n58788 , n58789 , n58790 , n58791 , n58792 , n58793 , n58794 , 
 n58795 , n58796 , n58797 , n58798 , n58799 , n58800 , n58801 , n58802 , n58803 , n58804 , 
 n58805 , n58806 , n58807 , n58808 , n58809 , n58810 , n58811 , n58812 , n58813 , n58814 , 
 n58815 , n58816 , n58817 , n58818 , n58819 , n58820 , n58821 , n58822 , n58823 , n58824 , 
 n58825 , n58826 , n58827 , n58828 , n58829 , n58830 , n58831 , n58832 , n58833 , n58834 , 
 n58835 , n58836 , n58837 , n58838 , n58839 , n58840 , n58841 , n58842 , n58843 , n58844 , 
 n58845 , n58846 , n58847 , n58848 , n58849 , n58850 , n58851 , n58852 , n58853 , n58854 , 
 n58855 , n58856 , n58857 , n58858 , n58859 , n58860 , n58861 , n58862 , n58863 , n58864 , 
 n58865 , n58866 , n58867 , n58868 , n58869 , n58870 , n58871 , n58872 , n58873 , n58874 , 
 n58875 , n58876 , n58877 , n58878 , n58879 , n58880 , n58881 , n58882 , n58883 , n58884 , 
 n58885 , n58886 , n58887 , n58888 , n58889 , n58890 , n58891 , n58892 , n58893 , n58894 , 
 n58895 , n58896 , n58897 , n58898 , n58899 , n58900 , n58901 , n58902 , n58903 , n58904 , 
 n58905 , n58906 , n58907 , n58908 , n58909 , n58910 , n58911 , n58912 , n58913 , n58914 , 
 n58915 , n58916 , n58917 , n58918 , n58919 , n58920 , n58921 , n58922 , n58923 , n58924 , 
 n58925 , n58926 , n58927 , n58928 , n58929 , n58930 , n58931 , n58932 , n58933 , n58934 , 
 n58935 , n58936 , n58937 , n58938 , n58939 , n58940 , n58941 , n58942 , n58943 , n58944 , 
 n58945 , n58946 , n58947 , n58948 , n58949 , n58950 , n58951 , n58952 , n58953 , n58954 , 
 n58955 , n58956 , n58957 , n58958 , n58959 , n58960 , n58961 , n58962 , n58963 , n58964 , 
 n58965 , n58966 , n58967 , n58968 , n58969 , n58970 , n58971 , n58972 , n58973 , n58974 , 
 n58975 , n58976 , n58977 , n58978 , n58979 , n58980 , n58981 , n58982 , n58983 , n58984 , 
 n58985 , n58986 , n58987 , n58988 , n58989 , n58990 , n58991 , n58992 , n58993 , n58994 , 
 n58995 , n58996 , n58997 , n58998 , n58999 , n59000 , n59001 , n59002 , n59003 , n59004 , 
 n59005 , n59006 , n59007 , n59008 , n59009 , n59010 , n59011 , n59012 , n59013 , n59014 , 
 n59015 , n59016 , n59017 , n59018 , n59019 , n59020 , n59021 , n59022 , n59023 , n59024 , 
 n59025 , n59026 , n59027 , n59028 , n59029 , n59030 , n59031 , n59032 , n59033 , n59034 , 
 n59035 , n59036 , n59037 , n59038 , n59039 , n59040 , n59041 , n59042 , n59043 , n59044 , 
 n59045 , n59046 , n59047 , n59048 , n59049 , n59050 , n59051 , n59052 , n59053 , n59054 , 
 n59055 , n59056 , n59057 , n59058 , n59059 , n59060 , n59061 , n59062 , n59063 , n59064 , 
 n59065 , n59066 , n59067 , n59068 , n59069 , n59070 , n59071 , n59072 , n59073 , n59074 , 
 n59075 , n59076 , n59077 , n59078 , n59079 , n59080 , n59081 , n59082 , n59083 , n59084 , 
 n59085 , n59086 , n59087 , n59088 , n59089 , n59090 , n59091 , n59092 , n59093 , n59094 , 
 n59095 , n59096 , n59097 , n59098 , n59099 , n59100 , n59101 , n59102 , n59103 , n59104 , 
 n59105 , n59106 , n59107 , n59108 , n59109 , n59110 , n59111 , n59112 , n59113 , n59114 , 
 n59115 , n59116 , n59117 , n59118 , n59119 , n59120 , n59121 , n59122 , n59123 , n59124 , 
 n59125 , n59126 , n59127 , n59128 , n59129 , n59130 , n59131 , n59132 , n59133 , n59134 , 
 n59135 , n59136 , n59137 , n59138 , n59139 , n59140 , n59141 , n59142 , n59143 , n59144 , 
 n59145 , n59146 , n59147 , n59148 , n59149 , n59150 , n59151 , n59152 , n59153 , n59154 , 
 n59155 , n59156 , n59157 , n59158 , n59159 , n59160 , n59161 , n59162 , n59163 , n59164 , 
 n59165 , n59166 , n59167 , n59168 , n59169 , n59170 , n59171 , n59172 , n59173 , n59174 , 
 n59175 , n59176 , n59177 , n59178 , n59179 , n59180 , n59181 , n59182 , n59183 , n59184 , 
 n59185 , n59186 , n59187 , n59188 , n59189 , n59190 , n59191 , n59192 , n59193 , n59194 , 
 n59195 , n59196 , n59197 , n59198 , n59199 , n59200 , n59201 , n59202 , n59203 , n59204 , 
 n59205 , n59206 , n59207 , n59208 , n59209 , n59210 , n59211 , n59212 , n59213 , n59214 , 
 n59215 , n59216 , n59217 , n59218 , n59219 , n59220 , n59221 , n59222 , n59223 , n59224 , 
 n59225 , n59226 , n59227 , n59228 , n59229 , n59230 , n59231 , n59232 , n59233 , n59234 , 
 n59235 , n59236 , n59237 , n59238 , n59239 , n59240 , n59241 , n59242 , n59243 , n59244 , 
 n59245 , n59246 , n59247 , n59248 , n59249 , n59250 , n59251 , n59252 , n59253 , n59254 , 
 n59255 , n59256 , n59257 , n59258 , n59259 , n59260 , n59261 , n59262 , n59263 , n59264 , 
 n59265 , n59266 , n59267 , n59268 , n59269 , n59270 , n59271 , n59272 , n59273 , n59274 , 
 n59275 , n59276 , n59277 , n59278 , n59279 , n59280 , n59281 , n59282 , n59283 , n59284 , 
 n59285 , n59286 , n59287 , n59288 , n59289 , n59290 , n59291 , n59292 , n59293 , n59294 , 
 n59295 , n59296 , n59297 , n59298 , n59299 , n59300 , n59301 , n59302 , n59303 , n59304 , 
 n59305 , n59306 , n59307 , n59308 , n59309 , n59310 , n59311 , n59312 , n59313 , n59314 , 
 n59315 , n59316 , n59317 , n59318 , n59319 , n59320 , n59321 , n59322 , n59323 , n59324 , 
 n59325 , n59326 , n59327 , n59328 , n59329 , n59330 , n59331 , n59332 , n59333 , n59334 , 
 n59335 , n59336 , n59337 , n59338 , n59339 , n59340 , n59341 , n59342 , n59343 , n59344 , 
 n59345 , n59346 , n59347 , n59348 , n59349 , n59350 , n59351 , n59352 , n59353 , n59354 , 
 n59355 , n59356 , n59357 , n59358 , n59359 , n59360 , n59361 , n59362 , n59363 , n59364 , 
 n59365 , n59366 , n59367 , n59368 , n59369 , n59370 , n59371 , n59372 , n59373 , n59374 , 
 n59375 , n59376 , n59377 , n59378 , n59379 , n59380 , n59381 , n59382 , n59383 , n59384 , 
 n59385 , n59386 , n59387 , n59388 , n59389 , n59390 , n59391 , n59392 , n59393 , n59394 , 
 n59395 , n59396 , n59397 , n59398 , n59399 , n59400 , n59401 , n59402 , n59403 , n59404 , 
 n59405 , n59406 , n59407 , n59408 , n59409 , n59410 , n59411 , n59412 , n59413 , n59414 , 
 n59415 , n59416 , n59417 , n59418 , n59419 , n59420 , n59421 , n59422 , n59423 , n59424 , 
 n59425 , n59426 , n59427 , n59428 , n59429 , n59430 , n59431 , n59432 , n59433 , n59434 , 
 n59435 , n59436 , n59437 , n59438 , n59439 , n59440 , n59441 , n59442 , n59443 , n59444 , 
 n59445 , n59446 , n59447 , n59448 , n59449 , n59450 , n59451 , n59452 , n59453 , n59454 , 
 n59455 , n59456 , n59457 , n59458 , n59459 , n59460 , n59461 , n59462 , n59463 , n59464 , 
 n59465 , n59466 , n59467 , n59468 , n59469 , n59470 , n59471 , n59472 , n59473 , n59474 , 
 n59475 , n59476 , n59477 , n59478 , n59479 , n59480 , n59481 , n59482 , n59483 , n59484 , 
 n59485 , n59486 , n59487 , n59488 , n59489 , n59490 , n59491 , n59492 , n59493 , n59494 , 
 n59495 , n59496 , n59497 , n59498 , n59499 , n59500 , n59501 , n59502 , n59503 , n59504 , 
 n59505 , n59506 , n59507 , n59508 , n59509 , n59510 , n59511 , n59512 , n59513 , n59514 , 
 n59515 , n59516 , n59517 , n59518 , n59519 , n59520 , n59521 , n59522 , n59523 , n59524 , 
 n59525 , n59526 , n59527 , n59528 , n59529 , n59530 , n59531 , n59532 , n59533 , n59534 , 
 n59535 , n59536 , n59537 , n59538 , n59539 , n59540 , n59541 , n59542 , n59543 , n59544 , 
 n59545 , n59546 , n59547 , n59548 , n59549 , n59550 , n59551 , n59552 , n59553 , n59554 , 
 n59555 , n59556 , n59557 , n59558 , n59559 , n59560 , n59561 , n59562 , n59563 , n59564 , 
 n59565 , n59566 , n59567 , n59568 , n59569 , n59570 , n59571 , n59572 , n59573 , n59574 , 
 n59575 , n59576 , n59577 , n59578 , n59579 , n59580 , n59581 , n59582 , n59583 , n59584 , 
 n59585 , n59586 , n59587 , n59588 , n59589 , n59590 , n59591 , n59592 , n59593 , n59594 , 
 n59595 , n59596 , n59597 , n59598 , n59599 , n59600 , n59601 , n59602 , n59603 , n59604 , 
 n59605 , n59606 , n59607 , n59608 , n59609 , n59610 , n59611 , n59612 , n59613 , n59614 , 
 n59615 , n59616 , n59617 , n59618 , n59619 , n59620 , n59621 , n59622 , n59623 , n59624 , 
 n59625 , n59626 , n59627 , n59628 , n59629 , n59630 , n59631 , n59632 , n59633 , n59634 , 
 n59635 , n59636 , n59637 , n59638 , n59639 , n59640 , n59641 , n59642 , n59643 , n59644 , 
 n59645 , n59646 , n59647 , n59648 , n59649 , n59650 , n59651 , n59652 , n59653 , n59654 , 
 n59655 , n59656 , n59657 , n59658 , n59659 , n59660 , n59661 , n59662 , n59663 , n59664 , 
 n59665 , n59666 , n59667 , n59668 , n59669 , n59670 , n59671 , n59672 , n59673 , n59674 , 
 n59675 , n59676 , n59677 , n59678 , n59679 , n59680 , n59681 , n59682 , n59683 , n59684 , 
 n59685 , n59686 , n59687 , n59688 , n59689 , n59690 , n59691 , n59692 , n59693 , n59694 , 
 n59695 , n59696 , n59697 , n59698 , n59699 , n59700 , n59701 , n59702 , n59703 , n59704 , 
 n59705 , n59706 , n59707 , n59708 , n59709 , n59710 , n59711 , n59712 , n59713 , n59714 , 
 n59715 , n59716 , n59717 , n59718 , n59719 , n59720 , n59721 , n59722 , n59723 , n59724 , 
 n59725 , n59726 , n59727 , n59728 , n59729 , n59730 , n59731 , n59732 , n59733 , n59734 , 
 n59735 , n59736 , n59737 , n59738 , n59739 , n59740 , n59741 , n59742 , n59743 , n59744 , 
 n59745 , n59746 , n59747 , n59748 , n59749 , n59750 , n59751 , n59752 , n59753 , n59754 , 
 n59755 , n59756 , n59757 , n59758 , n59759 , n59760 , n59761 , n59762 , n59763 , n59764 , 
 n59765 , n59766 , n59767 , n59768 , n59769 , n59770 , n59771 , n59772 , n59773 , n59774 , 
 n59775 , n59776 , n59777 , n59778 , n59779 , n59780 , n59781 , n59782 , n59783 , n59784 , 
 n59785 , n59786 , n59787 , n59788 , n59789 , n59790 , n59791 , n59792 , n59793 , n59794 , 
 n59795 , n59796 , n59797 , n59798 , n59799 , n59800 , n59801 , n59802 , n59803 , n59804 , 
 n59805 , n59806 , n59807 , n59808 , n59809 , n59810 , n59811 , n59812 , n59813 , n59814 , 
 n59815 , n59816 , n59817 , n59818 , n59819 , n59820 , n59821 , n59822 , n59823 , n59824 , 
 n59825 , n59826 , n59827 , n59828 , n59829 , n59830 , n59831 , n59832 , n59833 , n59834 , 
 n59835 , n59836 , n59837 , n59838 , n59839 , n59840 , n59841 , n59842 , n59843 , n59844 , 
 n59845 , n59846 , n59847 , n59848 , n59849 , n59850 , n59851 , n59852 , n59853 , n59854 , 
 n59855 , n59856 , n59857 , n59858 , n59859 , n59860 , n59861 , n59862 , n59863 , n59864 , 
 n59865 , n59866 , n59867 , n59868 , n59869 , n59870 , n59871 , n59872 , n59873 , n59874 , 
 n59875 , n59876 , n59877 , n59878 , n59879 , n59880 , n59881 , n59882 , n59883 , n59884 , 
 n59885 , n59886 , n59887 , n59888 , n59889 , n59890 , n59891 , n59892 , n59893 , n59894 , 
 n59895 , n59896 , n59897 , n59898 , n59899 , n59900 , n59901 , n59902 , n59903 , n59904 , 
 n59905 , n59906 , n59907 , n59908 , n59909 , n59910 , n59911 , n59912 , n59913 , n59914 , 
 n59915 , n59916 , n59917 , n59918 , n59919 , n59920 , n59921 , n59922 , n59923 , n59924 , 
 n59925 , n59926 , n59927 , n59928 , n59929 , n59930 , n59931 , n59932 , n59933 , n59934 , 
 n59935 , n59936 , n59937 , n59938 , n59939 , n59940 , n59941 , n59942 , n59943 , n59944 , 
 n59945 , n59946 , n59947 , n59948 , n59949 , n59950 , n59951 , n59952 , n59953 , n59954 , 
 n59955 , n59956 , n59957 , n59958 , n59959 , n59960 , n59961 , n59962 , n59963 , n59964 , 
 n59965 , n59966 , n59967 , n59968 , n59969 , n59970 , n59971 , n59972 , n59973 , n59974 , 
 n59975 , n59976 , n59977 , n59978 , n59979 , n59980 , n59981 , n59982 , n59983 , n59984 , 
 n59985 , n59986 , n59987 , n59988 , n59989 , n59990 , n59991 , n59992 , n59993 , n59994 , 
 n59995 , n59996 , n59997 , n59998 , n59999 , n60000 , n60001 , n60002 , n60003 , n60004 , 
 n60005 , n60006 , n60007 , n60008 , n60009 , n60010 , n60011 , n60012 , n60013 , n60014 , 
 n60015 , n60016 , n60017 , n60018 , n60019 , n60020 , n60021 , n60022 , n60023 , n60024 , 
 n60025 , n60026 , n60027 , n60028 , n60029 , n60030 , n60031 , n60032 , n60033 , n60034 , 
 n60035 , n60036 , n60037 , n60038 , n60039 , n60040 , n60041 , n60042 , n60043 , n60044 , 
 n60045 , n60046 , n60047 , n60048 , n60049 , n60050 , n60051 , n60052 , n60053 , n60054 , 
 n60055 , n60056 , n60057 , n60058 , n60059 , n60060 , n60061 , n60062 , n60063 , n60064 , 
 n60065 , n60066 , n60067 , n60068 , n60069 , n60070 , n60071 , n60072 , n60073 , n60074 , 
 n60075 , n60076 , n60077 , n60078 , n60079 , n60080 , n60081 , n60082 , n60083 , n60084 , 
 n60085 , n60086 , n60087 , n60088 , n60089 , n60090 , n60091 , n60092 , n60093 , n60094 , 
 n60095 , n60096 , n60097 , n60098 , n60099 , n60100 , n60101 , n60102 , n60103 , n60104 , 
 n60105 , n60106 , n60107 , n60108 , n60109 , n60110 , n60111 , n60112 , n60113 , n60114 , 
 n60115 , n60116 , n60117 , n60118 , n60119 , n60120 , n60121 , n60122 , n60123 , n60124 , 
 n60125 , n60126 , n60127 , n60128 , n60129 , n60130 , n60131 , n60132 , n60133 , n60134 , 
 n60135 , n60136 , n60137 , n60138 , n60139 , n60140 , n60141 , n60142 , n60143 , n60144 , 
 n60145 , n60146 , n60147 , n60148 , n60149 , n60150 , n60151 , n60152 , n60153 , n60154 , 
 n60155 , n60156 , n60157 , n60158 , n60159 , n60160 , n60161 , n60162 , n60163 , n60164 , 
 n60165 , n60166 , n60167 , n60168 , n60169 , n60170 , n60171 , n60172 , n60173 , n60174 , 
 n60175 , n60176 , n60177 , n60178 , n60179 , n60180 , n60181 , n60182 , n60183 , n60184 , 
 n60185 , n60186 , n60187 , n60188 , n60189 , n60190 , n60191 , n60192 , n60193 , n60194 , 
 n60195 , n60196 , n60197 , n60198 , n60199 , n60200 , n60201 , n60202 , n60203 , n60204 , 
 n60205 , n60206 , n60207 , n60208 , n60209 , n60210 , n60211 , n60212 , n60213 , n60214 , 
 n60215 , n60216 , n60217 , n60218 , n60219 , n60220 , n60221 , n60222 , n60223 , n60224 , 
 n60225 , n60226 , n60227 , n60228 , n60229 , n60230 , n60231 , n60232 , n60233 , n60234 , 
 n60235 , n60236 , n60237 , n60238 , n60239 , n60240 , n60241 , n60242 , n60243 , n60244 , 
 n60245 , n60246 , n60247 , n60248 , n60249 , n60250 , n60251 , n60252 , n60253 , n60254 , 
 n60255 , n60256 , n60257 , n60258 , n60259 , n60260 , n60261 , n60262 , n60263 , n60264 , 
 n60265 , n60266 , n60267 , n60268 , n60269 , n60270 , n60271 , n60272 , n60273 , n60274 , 
 n60275 , n60276 , n60277 , n60278 , n60279 , n60280 , n60281 , n60282 , n60283 , n60284 , 
 n60285 , n60286 , n60287 , n60288 , n60289 , n60290 , n60291 , n60292 , n60293 , n60294 , 
 n60295 , n60296 , n60297 , n60298 , n60299 , n60300 , n60301 , n60302 , n60303 , n60304 , 
 n60305 , n60306 , n60307 , n60308 , n60309 , n60310 , n60311 , n60312 , n60313 , n60314 , 
 n60315 , n60316 , n60317 , n60318 , n60319 , n60320 , n60321 , n60322 , n60323 , n60324 , 
 n60325 , n60326 , n60327 , n60328 , n60329 , n60330 , n60331 , n60332 , n60333 , n60334 , 
 n60335 , n60336 , n60337 , n60338 , n60339 , n60340 , n60341 , n60342 , n60343 , n60344 , 
 n60345 , n60346 , n60347 , n60348 , n60349 , n60350 , n60351 , n60352 , n60353 , n60354 , 
 n60355 , n60356 , n60357 , n60358 , n60359 , n60360 , n60361 , n60362 , n60363 , n60364 , 
 n60365 , n60366 , n60367 , n60368 , n60369 , n60370 , n60371 , n60372 , n60373 , n60374 , 
 n60375 , n60376 , n60377 , n60378 , n60379 , n60380 , n60381 , n60382 , n60383 , n60384 , 
 n60385 , n60386 , n60387 , n60388 , n60389 , n60390 , n60391 , n60392 , n60393 , n60394 , 
 n60395 , n60396 , n60397 , n60398 , n60399 , n60400 , n60401 , n60402 , n60403 , n60404 , 
 n60405 , n60406 , n60407 , n60408 , n60409 , n60410 , n60411 , n60412 , n60413 , n60414 , 
 n60415 , n60416 , n60417 , n60418 , n60419 , n60420 , n60421 , n60422 , n60423 , n60424 , 
 n60425 , n60426 , n60427 , n60428 , n60429 , n60430 , n60431 , n60432 , n60433 , n60434 , 
 n60435 , n60436 , n60437 , n60438 , n60439 , n60440 , n60441 , n60442 , n60443 , n60444 , 
 n60445 , n60446 , n60447 , n60448 , n60449 , n60450 , n60451 , n60452 , n60453 , n60454 , 
 n60455 , n60456 , n60457 , n60458 , n60459 , n60460 , n60461 , n60462 , n60463 , n60464 , 
 n60465 , n60466 , n60467 , n60468 , n60469 , n60470 , n60471 , n60472 , n60473 , n60474 , 
 n60475 , n60476 , n60477 , n60478 , n60479 , n60480 , n60481 , n60482 , n60483 , n60484 , 
 n60485 , n60486 , n60487 , n60488 , n60489 , n60490 , n60491 , n60492 , n60493 , n60494 , 
 n60495 , n60496 , n60497 , n60498 , n60499 , n60500 , n60501 , n60502 , n60503 , n60504 , 
 n60505 , n60506 , n60507 , n60508 , n60509 , n60510 , n60511 , n60512 , n60513 , n60514 , 
 n60515 , n60516 , n60517 , n60518 , n60519 , n60520 , n60521 , n60522 , n60523 , n60524 , 
 n60525 , n60526 , n60527 , n60528 , n60529 , n60530 , n60531 , n60532 , n60533 , n60534 , 
 n60535 , n60536 , n60537 , n60538 , n60539 , n60540 , n60541 , n60542 , n60543 , n60544 , 
 n60545 , n60546 , n60547 , n60548 , n60549 , n60550 , n60551 , n60552 , n60553 , n60554 , 
 n60555 , n60556 , n60557 , n60558 , n60559 , n60560 , n60561 , n60562 , n60563 , n60564 , 
 n60565 , n60566 , n60567 , n60568 , n60569 , n60570 , n60571 , n60572 , n60573 , n60574 , 
 n60575 , n60576 , n60577 , n60578 , n60579 , n60580 , n60581 , n60582 , n60583 , n60584 , 
 n60585 , n60586 , n60587 , n60588 , n60589 , n60590 , n60591 , n60592 , n60593 , n60594 , 
 n60595 , n60596 , n60597 , n60598 , n60599 , n60600 , n60601 , n60602 , n60603 , n60604 , 
 n60605 , n60606 , n60607 , n60608 , n60609 , n60610 , n60611 , n60612 , n60613 , n60614 , 
 n60615 , n60616 , n60617 , n60618 , n60619 , n60620 , n60621 , n60622 , n60623 , n60624 , 
 n60625 , n60626 , n60627 , n60628 , n60629 , n60630 , n60631 , n60632 , n60633 , n60634 , 
 n60635 , n60636 , n60637 , n60638 , n60639 , n60640 , n60641 , n60642 , n60643 , n60644 , 
 n60645 , n60646 , n60647 , n60648 , n60649 , n60650 , n60651 , n60652 , n60653 , n60654 , 
 n60655 , n60656 , n60657 , n60658 , n60659 , n60660 , n60661 , n60662 , n60663 , n60664 , 
 n60665 , n60666 , n60667 , n60668 , n60669 , n60670 , n60671 , n60672 , n60673 , n60674 , 
 n60675 , n60676 , n60677 , n60678 , n60679 , n60680 , n60681 , n60682 , n60683 , n60684 , 
 n60685 , n60686 , n60687 , n60688 , n60689 , n60690 , n60691 , n60692 , n60693 , n60694 , 
 n60695 , n60696 , n60697 , n60698 , n60699 , n60700 , n60701 , n60702 , n60703 , n60704 , 
 n60705 , n60706 , n60707 , n60708 , n60709 , n60710 , n60711 , n60712 , n60713 , n60714 , 
 n60715 , n60716 , n60717 , n60718 , n60719 , n60720 , n60721 , n60722 , n60723 , n60724 , 
 n60725 , n60726 , n60727 , n60728 , n60729 , n60730 , n60731 , n60732 , n60733 , n60734 , 
 n60735 , n60736 , n60737 , n60738 , n60739 , n60740 , n60741 , n60742 , n60743 , n60744 , 
 n60745 , n60746 , n60747 , n60748 , n60749 , n60750 , n60751 , n60752 , n60753 , n60754 , 
 n60755 , n60756 , n60757 , n60758 , n60759 , n60760 , n60761 , n60762 , n60763 , n60764 , 
 n60765 , n60766 , n60767 , n60768 , n60769 , n60770 , n60771 , n60772 , n60773 , n60774 , 
 n60775 , n60776 , n60777 , n60778 , n60779 , n60780 , n60781 , n60782 , n60783 , n60784 , 
 n60785 , n60786 , n60787 , n60788 , n60789 , n60790 , n60791 , n60792 , n60793 , n60794 , 
 n60795 , n60796 , n60797 , n60798 , n60799 , n60800 , n60801 , n60802 , n60803 , n60804 , 
 n60805 , n60806 , n60807 , n60808 , n60809 , n60810 , n60811 , n60812 , n60813 , n60814 , 
 n60815 , n60816 , n60817 , n60818 , n60819 , n60820 , n60821 , n60822 , n60823 , n60824 , 
 n60825 , n60826 , n60827 , n60828 , n60829 , n60830 , n60831 , n60832 , n60833 , n60834 , 
 n60835 , n60836 , n60837 , n60838 , n60839 , n60840 , n60841 , n60842 , n60843 , n60844 , 
 n60845 , n60846 , n60847 , n60848 , n60849 , n60850 , n60851 , n60852 , n60853 , n60854 , 
 n60855 , n60856 , n60857 , n60858 , n60859 , n60860 , n60861 , n60862 , n60863 , n60864 , 
 n60865 , n60866 , n60867 , n60868 , n60869 , n60870 , n60871 , n60872 , n60873 , n60874 , 
 n60875 , n60876 , n60877 , n60878 , n60879 , n60880 , n60881 , n60882 , n60883 , n60884 , 
 n60885 , n60886 , n60887 , n60888 , n60889 , n60890 , n60891 , n60892 , n60893 , n60894 , 
 n60895 , n60896 , n60897 , n60898 , n60899 , n60900 , n60901 , n60902 , n60903 , n60904 , 
 n60905 , n60906 , n60907 , n60908 , n60909 , n60910 , n60911 , n60912 , n60913 , n60914 , 
 n60915 , n60916 , n60917 , n60918 , n60919 , n60920 , n60921 , n60922 , n60923 , n60924 , 
 n60925 , n60926 , n60927 , n60928 , n60929 , n60930 , n60931 , n60932 , n60933 , n60934 , 
 n60935 , n60936 , n60937 , n60938 , n60939 , n60940 , n60941 , n60942 , n60943 , n60944 , 
 n60945 , n60946 , n60947 , n60948 , n60949 , n60950 , n60951 , n60952 , n60953 , n60954 , 
 n60955 , n60956 , n60957 , n60958 , n60959 , n60960 , n60961 , n60962 , n60963 , n60964 , 
 n60965 , n60966 , n60967 , n60968 , n60969 , n60970 , n60971 , n60972 , n60973 , n60974 , 
 n60975 , n60976 , n60977 , n60978 , n60979 , n60980 , n60981 , n60982 , n60983 , n60984 , 
 n60985 , n60986 , n60987 , n60988 , n60989 , n60990 , n60991 , n60992 , n60993 , n60994 , 
 n60995 , n60996 , n60997 , n60998 , n60999 , n61000 , n61001 , n61002 , n61003 , n61004 , 
 n61005 , n61006 , n61007 , n61008 , n61009 , n61010 , n61011 , n61012 , n61013 , n61014 , 
 n61015 , n61016 , n61017 , n61018 , n61019 , n61020 , n61021 , n61022 , n61023 , n61024 , 
 n61025 , n61026 , n61027 , n61028 , n61029 , n61030 , n61031 , n61032 , n61033 , n61034 , 
 n61035 , n61036 , n61037 , n61038 , n61039 , n61040 , n61041 , n61042 , n61043 , n61044 , 
 n61045 , n61046 , n61047 , n61048 , n61049 , n61050 , n61051 , n61052 , n61053 , n61054 , 
 n61055 , n61056 , n61057 , n61058 , n61059 , n61060 , n61061 , n61062 , n61063 , n61064 , 
 n61065 , n61066 , n61067 , n61068 , n61069 , n61070 , n61071 , n61072 , n61073 , n61074 , 
 n61075 , n61076 , n61077 , n61078 , n61079 , n61080 , n61081 , n61082 , n61083 , n61084 , 
 n61085 , n61086 , n61087 , n61088 , n61089 , n61090 , n61091 , n61092 , n61093 , n61094 , 
 n61095 , n61096 , n61097 , n61098 , n61099 , n61100 , n61101 , n61102 , n61103 , n61104 , 
 n61105 , n61106 , n61107 , n61108 , n61109 , n61110 , n61111 , n61112 , n61113 , n61114 , 
 n61115 , n61116 , n61117 , n61118 , n61119 , n61120 , n61121 , n61122 , n61123 , n61124 , 
 n61125 , n61126 , n61127 , n61128 , n61129 , n61130 , n61131 , n61132 , n61133 , n61134 , 
 n61135 , n61136 , n61137 , n61138 , n61139 , n61140 , n61141 , n61142 , n61143 , n61144 , 
 n61145 , n61146 , n61147 , n61148 , n61149 , n61150 , n61151 , n61152 , n61153 , n61154 , 
 n61155 , n61156 , n61157 , n61158 , n61159 , n61160 , n61161 , n61162 , n61163 , n61164 , 
 n61165 , n61166 , n61167 , n61168 , n61169 , n61170 , n61171 , n61172 , n61173 , n61174 , 
 n61175 , n61176 , n61177 , n61178 , n61179 , n61180 , n61181 , n61182 , n61183 , n61184 , 
 n61185 , n61186 , n61187 , n61188 , n61189 , n61190 , n61191 , n61192 , n61193 , n61194 , 
 n61195 , n61196 , n61197 , n61198 , n61199 , n61200 , n61201 , n61202 , n61203 , n61204 , 
 n61205 , n61206 , n61207 , n61208 , n61209 , n61210 , n61211 , n61212 , n61213 , n61214 , 
 n61215 , n61216 , n61217 , n61218 , n61219 , n61220 , n61221 , n61222 , n61223 , n61224 , 
 n61225 , n61226 , n61227 , n61228 , n61229 , n61230 , n61231 , n61232 , n61233 , n61234 , 
 n61235 , n61236 , n61237 , n61238 , n61239 , n61240 , n61241 , n61242 , n61243 , n61244 , 
 n61245 , n61246 , n61247 , n61248 , n61249 , n61250 , n61251 , n61252 , n61253 , n61254 , 
 n61255 , n61256 , n61257 , n61258 , n61259 , n61260 , n61261 , n61262 , n61263 , n61264 , 
 n61265 , n61266 , n61267 , n61268 , n61269 , n61270 , n61271 , n61272 , n61273 , n61274 , 
 n61275 , n61276 , n61277 , n61278 , n61279 , n61280 , n61281 , n61282 , n61283 , n61284 , 
 n61285 , n61286 , n61287 , n61288 , n61289 , n61290 , n61291 , n61292 , n61293 , n61294 , 
 n61295 , n61296 , n61297 , n61298 , n61299 , n61300 , n61301 , n61302 , n61303 , n61304 , 
 n61305 , n61306 , n61307 , n61308 , n61309 , n61310 , n61311 , n61312 , n61313 , n61314 , 
 n61315 , n61316 , n61317 , n61318 , n61319 , n61320 , n61321 , n61322 , n61323 , n61324 , 
 n61325 , n61326 , n61327 , n61328 , n61329 , n61330 , n61331 , n61332 , n61333 , n61334 , 
 n61335 , n61336 , n61337 , n61338 , n61339 , n61340 , n61341 , n61342 , n61343 , n61344 , 
 n61345 , n61346 , n61347 , n61348 , n61349 , n61350 , n61351 , n61352 , n61353 , n61354 , 
 n61355 , n61356 , n61357 , n61358 , n61359 , n61360 , n61361 , n61362 , n61363 , n61364 , 
 n61365 , n61366 , n61367 , n61368 , n61369 , n61370 , n61371 , n61372 , n61373 , n61374 , 
 n61375 , n61376 , n61377 , n61378 , n61379 , n61380 , n61381 , n61382 , n61383 , n61384 , 
 n61385 , n61386 , n61387 , n61388 , n61389 , n61390 , n61391 , n61392 , n61393 , n61394 , 
 n61395 , n61396 , n61397 , n61398 , n61399 , n61400 , n61401 , n61402 , n61403 , n61404 , 
 n61405 , n61406 , n61407 , n61408 , n61409 , n61410 , n61411 , n61412 , n61413 , n61414 , 
 n61415 , n61416 , n61417 , n61418 , n61419 , n61420 , n61421 , n61422 , n61423 , n61424 , 
 n61425 , n61426 , n61427 , n61428 , n61429 , n61430 , n61431 , n61432 , n61433 , n61434 , 
 n61435 , n61436 , n61437 , n61438 , n61439 , n61440 , n61441 , n61442 , n61443 , n61444 , 
 n61445 , n61446 , n61447 , n61448 , n61449 , n61450 , n61451 , n61452 , n61453 , n61454 , 
 n61455 , n61456 , n61457 , n61458 , n61459 , n61460 , n61461 , n61462 , n61463 , n61464 , 
 n61465 , n61466 , n61467 , n61468 , n61469 , n61470 , n61471 , n61472 , n61473 , n61474 , 
 n61475 , n61476 , n61477 , n61478 , n61479 , n61480 , n61481 , n61482 , n61483 , n61484 , 
 n61485 , n61486 , n61487 , n61488 , n61489 , n61490 , n61491 , n61492 , n61493 , n61494 , 
 n61495 , n61496 , n61497 , n61498 , n61499 , n61500 , n61501 , n61502 , n61503 , n61504 , 
 n61505 , n61506 , n61507 , n61508 , n61509 , n61510 , n61511 , n61512 , n61513 , n61514 , 
 n61515 , n61516 , n61517 , n61518 , n61519 , n61520 , n61521 , n61522 , n61523 , n61524 , 
 n61525 , n61526 , n61527 , n61528 , n61529 , n61530 , n61531 , n61532 , n61533 , n61534 , 
 n61535 , n61536 , n61537 , n61538 , n61539 , n61540 , n61541 , n61542 , n61543 , n61544 , 
 n61545 , n61546 , n61547 , n61548 , n61549 , n61550 , n61551 , n61552 , n61553 , n61554 , 
 n61555 , n61556 , n61557 , n61558 , n61559 , n61560 , n61561 , n61562 , n61563 , n61564 , 
 n61565 , n61566 , n61567 , n61568 , n61569 , n61570 , n61571 , n61572 , n61573 , n61574 , 
 n61575 , n61576 , n61577 , n61578 , n61579 , n61580 , n61581 , n61582 , n61583 , n61584 , 
 n61585 , n61586 , n61587 , n61588 , n61589 , n61590 , n61591 , n61592 , n61593 , n61594 , 
 n61595 , n61596 , n61597 , n61598 , n61599 , n61600 , n61601 , n61602 , n61603 , n61604 , 
 n61605 , n61606 , n61607 , n61608 , n61609 , n61610 , n61611 , n61612 , n61613 , n61614 , 
 n61615 , n61616 , n61617 , n61618 , n61619 , n61620 , n61621 , n61622 , n61623 , n61624 , 
 n61625 , n61626 , n61627 , n61628 , n61629 , n61630 , n61631 , n61632 , n61633 , n61634 , 
 n61635 , n61636 , n61637 , n61638 , n61639 , n61640 , n61641 , n61642 , n61643 , n61644 , 
 n61645 , n61646 , n61647 , n61648 , n61649 , n61650 , n61651 , n61652 , n61653 , n61654 , 
 n61655 , n61656 , n61657 , n61658 , n61659 , n61660 , n61661 , n61662 , n61663 , n61664 , 
 n61665 , n61666 , n61667 , n61668 , n61669 , n61670 , n61671 , n61672 , n61673 , n61674 , 
 n61675 , n61676 , n61677 , n61678 , n61679 , n61680 , n61681 , n61682 , n61683 , n61684 , 
 n61685 , n61686 , n61687 , n61688 , n61689 , n61690 , n61691 , n61692 , n61693 , n61694 , 
 n61695 , n61696 , n61697 , n61698 , n61699 , n61700 , n61701 , n61702 , n61703 , n61704 , 
 n61705 , n61706 , n61707 , n61708 , n61709 , n61710 , n61711 , n61712 , n61713 , n61714 , 
 n61715 , n61716 , n61717 , n61718 , n61719 , n61720 , n61721 , n61722 , n61723 , n61724 , 
 n61725 , n61726 , n61727 , n61728 , n61729 , n61730 , n61731 , n61732 , n61733 , n61734 , 
 n61735 , n61736 , n61737 , n61738 , n61739 , n61740 , n61741 , n61742 , n61743 , n61744 , 
 n61745 , n61746 , n61747 , n61748 , n61749 , n61750 , n61751 , n61752 , n61753 , n61754 , 
 n61755 , n61756 , n61757 , n61758 , n61759 , n61760 , n61761 , n61762 , n61763 , n61764 , 
 n61765 , n61766 , n61767 , n61768 , n61769 , n61770 , n61771 , n61772 , n61773 , n61774 , 
 n61775 , n61776 , n61777 , n61778 , n61779 , n61780 , n61781 , n61782 , n61783 , n61784 , 
 n61785 , n61786 , n61787 , n61788 , n61789 , n61790 , n61791 , n61792 , n61793 , n61794 , 
 n61795 , n61796 , n61797 , n61798 , n61799 , n61800 , n61801 , n61802 , n61803 , n61804 , 
 n61805 , n61806 , n61807 , n61808 , n61809 , n61810 , n61811 , n61812 , n61813 , n61814 , 
 n61815 , n61816 , n61817 , n61818 , n61819 , n61820 , n61821 , n61822 , n61823 , n61824 , 
 n61825 , n61826 , n61827 , n61828 , n61829 , n61830 , n61831 , n61832 , n61833 , n61834 , 
 n61835 , n61836 , n61837 , n61838 , n61839 , n61840 , n61841 , n61842 , n61843 , n61844 , 
 n61845 , n61846 , n61847 , n61848 , n61849 , n61850 , n61851 , n61852 , n61853 , n61854 , 
 n61855 , n61856 , n61857 , n61858 , n61859 , n61860 , n61861 , n61862 , n61863 , n61864 , 
 n61865 , n61866 , n61867 , n61868 , n61869 , n61870 , n61871 , n61872 , n61873 , n61874 , 
 n61875 , n61876 , n61877 , n61878 , n61879 , n61880 , n61881 , n61882 , n61883 , n61884 , 
 n61885 , n61886 , n61887 , n61888 , n61889 , n61890 , n61891 , n61892 , n61893 , n61894 , 
 n61895 , n61896 , n61897 , n61898 , n61899 , n61900 , n61901 , n61902 , n61903 , n61904 , 
 n61905 , n61906 , n61907 , n61908 , n61909 , n61910 , n61911 , n61912 , n61913 , n61914 , 
 n61915 , n61916 , n61917 , n61918 , n61919 , n61920 , n61921 , n61922 , n61923 , n61924 , 
 n61925 , n61926 , n61927 , n61928 , n61929 , n61930 , n61931 , n61932 , n61933 , n61934 , 
 n61935 , n61936 , n61937 , n61938 , n61939 , n61940 , n61941 , n61942 , n61943 , n61944 , 
 n61945 , n61946 , n61947 , n61948 , n61949 , n61950 , n61951 , n61952 , n61953 , n61954 , 
 n61955 , n61956 , n61957 , n61958 , n61959 , n61960 , n61961 , n61962 , n61963 , n61964 , 
 n61965 , n61966 , n61967 , n61968 , n61969 , n61970 , n61971 , n61972 , n61973 , n61974 , 
 n61975 , n61976 , n61977 , n61978 , n61979 , n61980 , n61981 , n61982 , n61983 , n61984 , 
 n61985 , n61986 , n61987 , n61988 , n61989 , n61990 , n61991 , n61992 , n61993 , n61994 , 
 n61995 , n61996 , n61997 , n61998 , n61999 , n62000 , n62001 , n62002 , n62003 , n62004 , 
 n62005 , n62006 , n62007 , n62008 , n62009 , n62010 , n62011 , n62012 , n62013 , n62014 , 
 n62015 , n62016 , n62017 , n62018 , n62019 , n62020 , n62021 , n62022 , n62023 , n62024 , 
 n62025 , n62026 , n62027 , n62028 , n62029 , n62030 , n62031 , n62032 , n62033 , n62034 , 
 n62035 , n62036 , n62037 , n62038 , n62039 , n62040 , n62041 , n62042 , n62043 , n62044 , 
 n62045 , n62046 , n62047 , n62048 , n62049 , n62050 , n62051 , n62052 , n62053 , n62054 , 
 n62055 , n62056 , n62057 , n62058 , n62059 , n62060 , n62061 , n62062 , n62063 , n62064 , 
 n62065 , n62066 , n62067 , n62068 , n62069 , n62070 , n62071 , n62072 , n62073 , n62074 , 
 n62075 , n62076 , n62077 , n62078 , n62079 , n62080 , n62081 , n62082 , n62083 , n62084 , 
 n62085 , n62086 , n62087 , n62088 , n62089 , n62090 , n62091 , n62092 , n62093 , n62094 , 
 n62095 , n62096 , n62097 , n62098 , n62099 , n62100 , n62101 , n62102 , n62103 , n62104 , 
 n62105 , n62106 , n62107 , n62108 , n62109 , n62110 , n62111 , n62112 , n62113 , n62114 , 
 n62115 , n62116 , n62117 , n62118 , n62119 , n62120 , n62121 , n62122 , n62123 , n62124 , 
 n62125 , n62126 , n62127 , n62128 , n62129 , n62130 , n62131 , n62132 , n62133 , n62134 , 
 n62135 , n62136 , n62137 , n62138 , n62139 , n62140 , n62141 , n62142 , n62143 , n62144 , 
 n62145 , n62146 , n62147 , n62148 , n62149 , n62150 , n62151 , n62152 , n62153 , n62154 , 
 n62155 , n62156 , n62157 , n62158 , n62159 , n62160 , n62161 , n62162 , n62163 , n62164 , 
 n62165 , n62166 , n62167 , n62168 , n62169 , n62170 , n62171 , n62172 , n62173 , n62174 , 
 n62175 , n62176 , n62177 , n62178 , n62179 , n62180 , n62181 , n62182 , n62183 , n62184 , 
 n62185 , n62186 , n62187 , n62188 , n62189 , n62190 , n62191 , n62192 , n62193 , n62194 , 
 n62195 , n62196 , n62197 , n62198 , n62199 , n62200 , n62201 , n62202 , n62203 , n62204 , 
 n62205 , n62206 , n62207 , n62208 , n62209 , n62210 , n62211 , n62212 , n62213 , n62214 , 
 n62215 , n62216 , n62217 , n62218 , n62219 , n62220 , n62221 , n62222 , n62223 , n62224 , 
 n62225 , n62226 , n62227 , n62228 , n62229 , n62230 , n62231 , n62232 , n62233 , n62234 , 
 n62235 , n62236 , n62237 , n62238 , n62239 , n62240 , n62241 , n62242 , n62243 , n62244 , 
 n62245 , n62246 , n62247 , n62248 , n62249 , n62250 , n62251 , n62252 , n62253 , n62254 , 
 n62255 , n62256 , n62257 , n62258 , n62259 , n62260 , n62261 , n62262 , n62263 , n62264 , 
 n62265 , n62266 , n62267 , n62268 , n62269 , n62270 , n62271 , n62272 , n62273 , n62274 , 
 n62275 , n62276 , n62277 , n62278 , n62279 , n62280 , n62281 , n62282 , n62283 , n62284 , 
 n62285 , n62286 , n62287 , n62288 , n62289 , n62290 , n62291 , n62292 , n62293 , n62294 , 
 n62295 , n62296 , n62297 , n62298 , n62299 , n62300 , n62301 , n62302 , n62303 , n62304 , 
 n62305 , n62306 , n62307 , n62308 , n62309 , n62310 , n62311 , n62312 , n62313 , n62314 , 
 n62315 , n62316 , n62317 , n62318 , n62319 , n62320 , n62321 , n62322 , n62323 , n62324 , 
 n62325 , n62326 , n62327 , n62328 , n62329 , n62330 , n62331 , n62332 , n62333 , n62334 , 
 n62335 , n62336 , n62337 , n62338 , n62339 , n62340 , n62341 , n62342 , n62343 , n62344 , 
 n62345 , n62346 , n62347 , n62348 , n62349 , n62350 , n62351 , n62352 , n62353 , n62354 , 
 n62355 , n62356 , n62357 , n62358 , n62359 , n62360 , n62361 , n62362 , n62363 , n62364 , 
 n62365 , n62366 , n62367 , n62368 , n62369 , n62370 , n62371 , n62372 , n62373 , n62374 , 
 n62375 , n62376 , n62377 , n62378 , n62379 , n62380 , n62381 , n62382 , n62383 , n62384 , 
 n62385 , n62386 , n62387 , n62388 , n62389 , n62390 , n62391 , n62392 , n62393 , n62394 , 
 n62395 , n62396 , n62397 , n62398 , n62399 , n62400 , n62401 , n62402 , n62403 , n62404 , 
 n62405 , n62406 , n62407 , n62408 , n62409 , n62410 , n62411 , n62412 , n62413 , n62414 , 
 n62415 , n62416 , n62417 , n62418 , n62419 , n62420 , n62421 , n62422 , n62423 , n62424 , 
 n62425 , n62426 , n62427 , n62428 , n62429 , n62430 , n62431 , n62432 , n62433 , n62434 , 
 n62435 , n62436 , n62437 , n62438 , n62439 , n62440 , n62441 , n62442 , n62443 , n62444 , 
 n62445 , n62446 , n62447 , n62448 , n62449 , n62450 , n62451 , n62452 , n62453 , n62454 , 
 n62455 , n62456 , n62457 , n62458 , n62459 , n62460 , n62461 , n62462 , n62463 , n62464 , 
 n62465 , n62466 , n62467 , n62468 , n62469 , n62470 , n62471 , n62472 , n62473 , n62474 , 
 n62475 , n62476 , n62477 , n62478 , n62479 , n62480 , n62481 , n62482 , n62483 , n62484 , 
 n62485 , n62486 , n62487 , n62488 , n62489 , n62490 , n62491 , n62492 , n62493 , n62494 , 
 n62495 , n62496 , n62497 , n62498 , n62499 , n62500 , n62501 , n62502 , n62503 , n62504 , 
 n62505 , n62506 , n62507 , n62508 , n62509 , n62510 , n62511 , n62512 , n62513 , n62514 , 
 n62515 , n62516 , n62517 , n62518 , n62519 , n62520 , n62521 , n62522 , n62523 , n62524 , 
 n62525 , n62526 , n62527 , n62528 , n62529 , n62530 , n62531 , n62532 , n62533 , n62534 , 
 n62535 , n62536 , n62537 , n62538 , n62539 , n62540 , n62541 , n62542 , n62543 , n62544 , 
 n62545 , n62546 , n62547 , n62548 , n62549 , n62550 , n62551 , n62552 , n62553 , n62554 , 
 n62555 , n62556 , n62557 , n62558 , n62559 , n62560 , n62561 , n62562 , n62563 , n62564 , 
 n62565 , n62566 , n62567 , n62568 , n62569 , n62570 , n62571 , n62572 , n62573 , n62574 , 
 n62575 , n62576 , n62577 , n62578 , n62579 , n62580 , n62581 , n62582 , n62583 , n62584 , 
 n62585 , n62586 , n62587 , n62588 , n62589 , n62590 , n62591 , n62592 , n62593 , n62594 , 
 n62595 , n62596 , n62597 , n62598 , n62599 , n62600 , n62601 , n62602 , n62603 , n62604 , 
 n62605 , n62606 , n62607 , n62608 , n62609 , n62610 , n62611 , n62612 , n62613 , n62614 , 
 n62615 , n62616 , n62617 , n62618 , n62619 , n62620 , n62621 , n62622 , n62623 , n62624 , 
 n62625 , n62626 , n62627 , n62628 , n62629 , n62630 , n62631 , n62632 , n62633 , n62634 , 
 n62635 , n62636 , n62637 , n62638 , n62639 , n62640 , n62641 , n62642 , n62643 , n62644 , 
 n62645 , n62646 , n62647 , n62648 , n62649 , n62650 , n62651 , n62652 , n62653 , n62654 , 
 n62655 , n62656 , n62657 , n62658 , n62659 , n62660 , n62661 , n62662 , n62663 , n62664 , 
 n62665 , n62666 , n62667 , n62668 , n62669 , n62670 , n62671 , n62672 , n62673 , n62674 , 
 n62675 , n62676 , n62677 , n62678 , n62679 , n62680 , n62681 , n62682 , n62683 , n62684 , 
 n62685 , n62686 , n62687 , n62688 , n62689 , n62690 , n62691 , n62692 , n62693 , n62694 , 
 n62695 , n62696 , n62697 , n62698 , n62699 , n62700 , n62701 , n62702 , n62703 , n62704 , 
 n62705 , n62706 , n62707 , n62708 , n62709 , n62710 , n62711 , n62712 , n62713 , n62714 , 
 n62715 , n62716 , n62717 , n62718 , n62719 , n62720 , n62721 , n62722 , n62723 , n62724 , 
 n62725 , n62726 , n62727 , n62728 , n62729 , n62730 , n62731 , n62732 , n62733 , n62734 , 
 n62735 , n62736 , n62737 , n62738 , n62739 , n62740 , n62741 , n62742 , n62743 , n62744 , 
 n62745 , n62746 , n62747 , n62748 , n62749 , n62750 , n62751 , n62752 , n62753 , n62754 , 
 n62755 , n62756 , n62757 , n62758 , n62759 , n62760 , n62761 , n62762 , n62763 , n62764 , 
 n62765 , n62766 , n62767 , n62768 , n62769 , n62770 , n62771 , n62772 , n62773 , n62774 , 
 n62775 , n62776 , n62777 , n62778 , n62779 , n62780 , n62781 , n62782 , n62783 , n62784 , 
 n62785 , n62786 , n62787 , n62788 , n62789 , n62790 , n62791 , n62792 , n62793 , n62794 , 
 n62795 , n62796 , n62797 , n62798 , n62799 , n62800 , n62801 , n62802 , n62803 , n62804 , 
 n62805 , n62806 , n62807 , n62808 , n62809 , n62810 , n62811 , n62812 , n62813 , n62814 , 
 n62815 , n62816 , n62817 , n62818 , n62819 , n62820 , n62821 , n62822 , n62823 , n62824 , 
 n62825 , n62826 , n62827 , n62828 , n62829 , n62830 , n62831 , n62832 , n62833 , n62834 , 
 n62835 , n62836 , n62837 , n62838 , n62839 , n62840 , n62841 , n62842 , n62843 , n62844 , 
 n62845 , n62846 , n62847 , n62848 , n62849 , n62850 , n62851 , n62852 , n62853 , n62854 , 
 n62855 , n62856 , n62857 , n62858 , n62859 , n62860 , n62861 , n62862 , n62863 , n62864 , 
 n62865 , n62866 , n62867 , n62868 , n62869 , n62870 , n62871 , n62872 , n62873 , n62874 , 
 n62875 , n62876 , n62877 , n62878 , n62879 , n62880 , n62881 , n62882 , n62883 , n62884 , 
 n62885 , n62886 , n62887 , n62888 , n62889 , n62890 , n62891 , n62892 , n62893 , n62894 , 
 n62895 , n62896 , n62897 , n62898 , n62899 , n62900 , n62901 , n62902 , n62903 , n62904 , 
 n62905 , n62906 , n62907 , n62908 , n62909 , n62910 , n62911 , n62912 , n62913 , n62914 , 
 n62915 , n62916 , n62917 , n62918 , n62919 , n62920 , n62921 , n62922 , n62923 , n62924 , 
 n62925 , n62926 , n62927 , n62928 , n62929 , n62930 , n62931 , n62932 , n62933 , n62934 , 
 n62935 , n62936 , n62937 , n62938 , n62939 , n62940 , n62941 , n62942 , n62943 , n62944 , 
 n62945 , n62946 , n62947 , n62948 , n62949 , n62950 , n62951 , n62952 , n62953 , n62954 , 
 n62955 , n62956 , n62957 , n62958 , n62959 , n62960 , n62961 , n62962 , n62963 , n62964 , 
 n62965 , n62966 , n62967 , n62968 , n62969 , n62970 , n62971 , n62972 , n62973 , n62974 , 
 n62975 , n62976 , n62977 , n62978 , n62979 , n62980 , n62981 , n62982 , n62983 , n62984 , 
 n62985 , n62986 , n62987 , n62988 , n62989 , n62990 , n62991 , n62992 , n62993 , n62994 , 
 n62995 , n62996 , n62997 , n62998 , n62999 , n63000 , n63001 , n63002 , n63003 , n63004 , 
 n63005 , n63006 , n63007 , n63008 , n63009 , n63010 , n63011 , n63012 , n63013 , n63014 , 
 n63015 , n63016 , n63017 , n63018 , n63019 , n63020 , n63021 , n63022 , n63023 , n63024 , 
 n63025 , n63026 , n63027 , n63028 , n63029 , n63030 , n63031 , n63032 , n63033 , n63034 , 
 n63035 , n63036 , n63037 , n63038 , n63039 , n63040 , n63041 , n63042 , n63043 , n63044 , 
 n63045 , n63046 , n63047 , n63048 , n63049 , n63050 , n63051 , n63052 , n63053 , n63054 , 
 n63055 , n63056 , n63057 , n63058 , n63059 , n63060 , n63061 , n63062 , n63063 , n63064 , 
 n63065 , n63066 , n63067 , n63068 , n63069 , n63070 , n63071 , n63072 , n63073 , n63074 , 
 n63075 , n63076 , n63077 , n63078 , n63079 , n63080 , n63081 , n63082 , n63083 , n63084 , 
 n63085 , n63086 , n63087 , n63088 , n63089 , n63090 , n63091 , n63092 , n63093 , n63094 , 
 n63095 , n63096 , n63097 , n63098 , n63099 , n63100 , n63101 , n63102 , n63103 , n63104 , 
 n63105 , n63106 , n63107 , n63108 , n63109 , n63110 , n63111 , n63112 , n63113 , n63114 , 
 n63115 , n63116 , n63117 , n63118 , n63119 , n63120 , n63121 , n63122 , n63123 , n63124 , 
 n63125 , n63126 , n63127 , n63128 , n63129 , n63130 , n63131 , n63132 , n63133 , n63134 , 
 n63135 , n63136 , n63137 , n63138 , n63139 , n63140 , n63141 , n63142 , n63143 , n63144 , 
 n63145 , n63146 , n63147 , n63148 , n63149 , n63150 , n63151 , n63152 , n63153 , n63154 , 
 n63155 , n63156 , n63157 , n63158 , n63159 , n63160 , n63161 , n63162 , n63163 , n63164 , 
 n63165 , n63166 , n63167 , n63168 , n63169 , n63170 , n63171 , n63172 , n63173 , n63174 , 
 n63175 , n63176 , n63177 , n63178 , n63179 , n63180 , n63181 , n63182 , n63183 , n63184 , 
 n63185 , n63186 , n63187 , n63188 , n63189 , n63190 , n63191 , n63192 , n63193 , n63194 , 
 n63195 , n63196 , n63197 , n63198 , n63199 , n63200 , n63201 , n63202 , n63203 , n63204 , 
 n63205 , n63206 , n63207 , n63208 , n63209 , n63210 , n63211 , n63212 , n63213 , n63214 , 
 n63215 , n63216 , n63217 , n63218 , n63219 , n63220 , n63221 , n63222 , n63223 , n63224 , 
 n63225 , n63226 , n63227 , n63228 , n63229 , n63230 , n63231 , n63232 , n63233 , n63234 , 
 n63235 , n63236 , n63237 , n63238 , n63239 , n63240 , n63241 , n63242 , n63243 , n63244 , 
 n63245 , n63246 , n63247 , n63248 , n63249 , n63250 , n63251 , n63252 , n63253 , n63254 , 
 n63255 , n63256 , n63257 , n63258 , n63259 , n63260 , n63261 , n63262 , n63263 , n63264 , 
 n63265 , n63266 , n63267 , n63268 , n63269 , n63270 , n63271 , n63272 , n63273 , n63274 , 
 n63275 , n63276 , n63277 , n63278 , n63279 , n63280 , n63281 , n63282 , n63283 , n63284 , 
 n63285 , n63286 , n63287 , n63288 , n63289 , n63290 , n63291 , n63292 , n63293 , n63294 , 
 n63295 , n63296 , n63297 , n63298 , n63299 , n63300 , n63301 , n63302 , n63303 , n63304 , 
 n63305 , n63306 , n63307 , n63308 , n63309 , n63310 , n63311 , n63312 , n63313 , n63314 , 
 n63315 , n63316 , n63317 , n63318 , n63319 , n63320 , n63321 , n63322 , n63323 , n63324 , 
 n63325 , n63326 , n63327 , n63328 , n63329 , n63330 , n63331 , n63332 , n63333 , n63334 , 
 n63335 , n63336 , n63337 , n63338 , n63339 , n63340 , n63341 , n63342 , n63343 , n63344 , 
 n63345 , n63346 , n63347 , n63348 , n63349 , n63350 , n63351 , n63352 , n63353 , n63354 , 
 n63355 , n63356 , n63357 , n63358 , n63359 , n63360 , n63361 , n63362 , n63363 , n63364 , 
 n63365 , n63366 , n63367 , n63368 , n63369 , n63370 , n63371 , n63372 , n63373 , n63374 , 
 n63375 , n63376 , n63377 , n63378 , n63379 , n63380 , n63381 , n63382 , n63383 , n63384 , 
 n63385 , n63386 , n63387 , n63388 , n63389 , n63390 , n63391 , n63392 , n63393 , n63394 , 
 n63395 , n63396 , n63397 , n63398 , n63399 , n63400 , n63401 , n63402 , n63403 , n63404 , 
 n63405 , n63406 , n63407 , n63408 , n63409 , n63410 , n63411 , n63412 , n63413 , n63414 , 
 n63415 , n63416 , n63417 , n63418 , n63419 , n63420 , n63421 , n63422 , n63423 , n63424 , 
 n63425 , n63426 , n63427 , n63428 , n63429 , n63430 , n63431 , n63432 , n63433 , n63434 , 
 n63435 , n63436 , n63437 , n63438 , n63439 , n63440 , n63441 , n63442 , n63443 , n63444 , 
 n63445 , n63446 , n63447 , n63448 , n63449 , n63450 , n63451 , n63452 , n63453 , n63454 , 
 n63455 , n63456 , n63457 , n63458 , n63459 , n63460 , n63461 , n63462 , n63463 , n63464 , 
 n63465 , n63466 , n63467 , n63468 , n63469 , n63470 , n63471 , n63472 , n63473 , n63474 , 
 n63475 , n63476 , n63477 , n63478 , n63479 , n63480 , n63481 , n63482 , n63483 , n63484 , 
 n63485 , n63486 , n63487 , n63488 , n63489 , n63490 , n63491 , n63492 , n63493 , n63494 , 
 n63495 , n63496 , n63497 , n63498 , n63499 , n63500 , n63501 , n63502 , n63503 , n63504 , 
 n63505 , n63506 , n63507 , n63508 , n63509 , n63510 , n63511 , n63512 , n63513 , n63514 , 
 n63515 , n63516 , n63517 , n63518 , n63519 , n63520 , n63521 , n63522 , n63523 , n63524 , 
 n63525 , n63526 , n63527 , n63528 , n63529 , n63530 , n63531 , n63532 , n63533 , n63534 , 
 n63535 , n63536 , n63537 , n63538 , n63539 , n63540 , n63541 , n63542 , n63543 , n63544 , 
 n63545 , n63546 , n63547 , n63548 , n63549 , n63550 , n63551 , n63552 , n63553 , n63554 , 
 n63555 , n63556 , n63557 , n63558 , n63559 , n63560 , n63561 , n63562 , n63563 , n63564 , 
 n63565 , n63566 , n63567 , n63568 , n63569 , n63570 , n63571 , n63572 , n63573 , n63574 , 
 n63575 , n63576 , n63577 , n63578 , n63579 , n63580 , n63581 , n63582 , n63583 , n63584 , 
 n63585 , n63586 , n63587 , n63588 , n63589 , n63590 , n63591 , n63592 , n63593 , n63594 , 
 n63595 , n63596 , n63597 , n63598 , n63599 , n63600 , n63601 , n63602 , n63603 , n63604 , 
 n63605 , n63606 , n63607 , n63608 , n63609 , n63610 , n63611 , n63612 , n63613 , n63614 , 
 n63615 , n63616 , n63617 , n63618 , n63619 , n63620 , n63621 , n63622 , n63623 , n63624 , 
 n63625 , n63626 , n63627 , n63628 , n63629 , n63630 , n63631 , n63632 , n63633 , n63634 , 
 n63635 , n63636 , n63637 , n63638 , n63639 , n63640 , n63641 , n63642 , n63643 , n63644 , 
 n63645 , n63646 , n63647 , n63648 , n63649 , n63650 , n63651 , n63652 , n63653 , n63654 , 
 n63655 , n63656 , n63657 , n63658 , n63659 , n63660 , n63661 , n63662 , n63663 , n63664 , 
 n63665 , n63666 , n63667 , n63668 , n63669 , n63670 , n63671 , n63672 , n63673 , n63674 , 
 n63675 , n63676 , n63677 , n63678 , n63679 , n63680 , n63681 , n63682 , n63683 , n63684 , 
 n63685 , n63686 , n63687 , n63688 , n63689 , n63690 , n63691 , n63692 , n63693 , n63694 , 
 n63695 , n63696 , n63697 , n63698 , n63699 , n63700 , n63701 , n63702 , n63703 , n63704 , 
 n63705 , n63706 , n63707 , n63708 , n63709 , n63710 , n63711 , n63712 , n63713 , n63714 , 
 n63715 , n63716 , n63717 , n63718 , n63719 , n63720 , n63721 , n63722 , n63723 , n63724 , 
 n63725 , n63726 , n63727 , n63728 , n63729 , n63730 , n63731 , n63732 , n63733 , n63734 , 
 n63735 , n63736 , n63737 , n63738 , n63739 , n63740 , n63741 , n63742 , n63743 , n63744 , 
 n63745 , n63746 , n63747 , n63748 , n63749 , n63750 , n63751 , n63752 , n63753 , n63754 , 
 n63755 , n63756 , n63757 , n63758 , n63759 , n63760 , n63761 , n63762 , n63763 , n63764 , 
 n63765 , n63766 , n63767 , n63768 , n63769 , n63770 , n63771 , n63772 , n63773 , n63774 , 
 n63775 , n63776 , n63777 , n63778 , n63779 , n63780 , n63781 , n63782 , n63783 , n63784 , 
 n63785 , n63786 , n63787 , n63788 , n63789 , n63790 , n63791 , n63792 , n63793 , n63794 , 
 n63795 , n63796 , n63797 , n63798 , n63799 , n63800 , n63801 , n63802 , n63803 , n63804 , 
 n63805 , n63806 , n63807 , n63808 , n63809 , n63810 , n63811 , n63812 , n63813 , n63814 , 
 n63815 , n63816 , n63817 , n63818 , n63819 , n63820 , n63821 , n63822 , n63823 , n63824 , 
 n63825 , n63826 , n63827 , n63828 , n63829 , n63830 , n63831 , n63832 , n63833 , n63834 , 
 n63835 , n63836 , n63837 , n63838 , n63839 , n63840 , n63841 , n63842 , n63843 , n63844 , 
 n63845 , n63846 , n63847 , n63848 , n63849 , n63850 , n63851 , n63852 , n63853 , n63854 , 
 n63855 , n63856 , n63857 , n63858 , n63859 , n63860 , n63861 , n63862 , n63863 , n63864 , 
 n63865 , n63866 , n63867 , n63868 , n63869 , n63870 , n63871 , n63872 , n63873 , n63874 , 
 n63875 , n63876 , n63877 , n63878 , n63879 , n63880 , n63881 , n63882 , n63883 , n63884 , 
 n63885 , n63886 , n63887 , n63888 , n63889 , n63890 , n63891 , n63892 , n63893 , n63894 , 
 n63895 , n63896 , n63897 , n63898 , n63899 , n63900 , n63901 , n63902 , n63903 , n63904 , 
 n63905 , n63906 , n63907 , n63908 , n63909 , n63910 , n63911 , n63912 , n63913 , n63914 , 
 n63915 , n63916 , n63917 , n63918 , n63919 , n63920 , n63921 , n63922 , n63923 , n63924 , 
 n63925 , n63926 , n63927 , n63928 , n63929 , n63930 , n63931 , n63932 , n63933 , n63934 , 
 n63935 , n63936 , n63937 , n63938 , n63939 , n63940 , n63941 , n63942 , n63943 , n63944 , 
 n63945 , n63946 , n63947 , n63948 , n63949 , n63950 , n63951 , n63952 , n63953 , n63954 , 
 n63955 , n63956 , n63957 , n63958 , n63959 , n63960 , n63961 , n63962 , n63963 , n63964 , 
 n63965 , n63966 , n63967 , n63968 , n63969 , n63970 , n63971 , n63972 , n63973 , n63974 , 
 n63975 , n63976 , n63977 , n63978 , n63979 , n63980 , n63981 , n63982 , n63983 , n63984 , 
 n63985 , n63986 , n63987 , n63988 , n63989 , n63990 , n63991 , n63992 , n63993 , n63994 , 
 n63995 , n63996 , n63997 , n63998 , n63999 , n64000 , n64001 , n64002 , n64003 , n64004 , 
 n64005 , n64006 , n64007 , n64008 , n64009 , n64010 , n64011 , n64012 , n64013 , n64014 , 
 n64015 , n64016 , n64017 , n64018 , n64019 , n64020 , n64021 , n64022 , n64023 , n64024 , 
 n64025 , n64026 , n64027 , n64028 , n64029 , n64030 , n64031 , n64032 , n64033 , n64034 , 
 n64035 , n64036 , n64037 , n64038 , n64039 , n64040 , n64041 , n64042 , n64043 , n64044 , 
 n64045 , n64046 , n64047 , n64048 , n64049 , n64050 , n64051 , n64052 , n64053 , n64054 , 
 n64055 , n64056 , n64057 , n64058 , n64059 , n64060 , n64061 , n64062 , n64063 , n64064 , 
 n64065 , n64066 , n64067 , n64068 , n64069 , n64070 , n64071 , n64072 , n64073 , n64074 , 
 n64075 , n64076 , n64077 , n64078 , n64079 , n64080 , n64081 , n64082 , n64083 , n64084 , 
 n64085 , n64086 , n64087 , n64088 , n64089 , n64090 , n64091 , n64092 , n64093 , n64094 , 
 n64095 , n64096 , n64097 , n64098 , n64099 , n64100 , n64101 , n64102 , n64103 , n64104 , 
 n64105 , n64106 , n64107 , n64108 , n64109 , n64110 , n64111 , n64112 , n64113 , n64114 , 
 n64115 , n64116 , n64117 , n64118 , n64119 , n64120 , n64121 , n64122 , n64123 , n64124 , 
 n64125 , n64126 , n64127 , n64128 , n64129 , n64130 , n64131 , n64132 , n64133 , n64134 , 
 n64135 , n64136 , n64137 , n64138 , n64139 , n64140 , n64141 , n64142 , n64143 , n64144 , 
 n64145 , n64146 , n64147 , n64148 , n64149 , n64150 , n64151 , n64152 , n64153 , n64154 , 
 n64155 , n64156 , n64157 , n64158 , n64159 , n64160 , n64161 , n64162 , n64163 , n64164 , 
 n64165 , n64166 , n64167 , n64168 , n64169 , n64170 , n64171 , n64172 , n64173 , n64174 , 
 n64175 , n64176 , n64177 , n64178 , n64179 , n64180 , n64181 , n64182 , n64183 , n64184 , 
 n64185 , n64186 , n64187 , n64188 , n64189 , n64190 , n64191 , n64192 , n64193 , n64194 , 
 n64195 , n64196 , n64197 , n64198 , n64199 , n64200 , n64201 , n64202 , n64203 , n64204 , 
 n64205 , n64206 , n64207 , n64208 , n64209 , n64210 , n64211 , n64212 , n64213 , n64214 , 
 n64215 , n64216 , n64217 , n64218 , n64219 , n64220 , n64221 , n64222 , n64223 , n64224 , 
 n64225 , n64226 , n64227 , n64228 , n64229 , n64230 , n64231 , n64232 , n64233 , n64234 , 
 n64235 , n64236 , n64237 , n64238 , n64239 , n64240 , n64241 , n64242 , n64243 , n64244 , 
 n64245 , n64246 , n64247 , n64248 , n64249 , n64250 , n64251 , n64252 , n64253 , n64254 , 
 n64255 , n64256 , n64257 , n64258 , n64259 , n64260 , n64261 , n64262 , n64263 , n64264 , 
 n64265 , n64266 , n64267 , n64268 , n64269 , n64270 , n64271 , n64272 , n64273 , n64274 , 
 n64275 , n64276 , n64277 , n64278 , n64279 , n64280 , n64281 , n64282 , n64283 , n64284 , 
 n64285 , n64286 , n64287 , n64288 , n64289 , n64290 , n64291 , n64292 , n64293 , n64294 , 
 n64295 , n64296 , n64297 , n64298 , n64299 , n64300 , n64301 , n64302 , n64303 , n64304 , 
 n64305 , n64306 , n64307 , n64308 , n64309 , n64310 , n64311 , n64312 , n64313 , n64314 , 
 n64315 , n64316 , n64317 , n64318 , n64319 , n64320 , n64321 , n64322 , n64323 , n64324 , 
 n64325 , n64326 , n64327 , n64328 , n64329 , n64330 , n64331 , n64332 , n64333 , n64334 , 
 n64335 , n64336 , n64337 , n64338 , n64339 , n64340 , n64341 , n64342 , n64343 , n64344 , 
 n64345 , n64346 , n64347 , n64348 , n64349 , n64350 , n64351 , n64352 , n64353 , n64354 , 
 n64355 , n64356 , n64357 , n64358 , n64359 , n64360 , n64361 , n64362 , n64363 , n64364 , 
 n64365 , n64366 , n64367 , n64368 , n64369 , n64370 , n64371 , n64372 , n64373 , n64374 , 
 n64375 , n64376 , n64377 , n64378 , n64379 , n64380 , n64381 , n64382 , n64383 , n64384 , 
 n64385 , n64386 , n64387 , n64388 , n64389 , n64390 , n64391 , n64392 , n64393 , n64394 , 
 n64395 , n64396 , n64397 , n64398 , n64399 , n64400 , n64401 , n64402 , n64403 , n64404 , 
 n64405 , n64406 , n64407 , n64408 , n64409 , n64410 , n64411 , n64412 , n64413 , n64414 , 
 n64415 , n64416 , n64417 , n64418 , n64419 , n64420 , n64421 , n64422 , n64423 , n64424 , 
 n64425 , n64426 , n64427 , n64428 , n64429 , n64430 , n64431 , n64432 , n64433 , n64434 , 
 n64435 , n64436 , n64437 , n64438 , n64439 , n64440 , n64441 , n64442 , n64443 , n64444 , 
 n64445 , n64446 , n64447 , n64448 , n64449 , n64450 , n64451 , n64452 , n64453 , n64454 , 
 n64455 , n64456 , n64457 , n64458 , n64459 , n64460 , n64461 , n64462 , n64463 , n64464 , 
 n64465 , n64466 , n64467 , n64468 , n64469 , n64470 , n64471 , n64472 , n64473 , n64474 , 
 n64475 , n64476 , n64477 , n64478 , n64479 , n64480 , n64481 , n64482 , n64483 , n64484 , 
 n64485 , n64486 , n64487 , n64488 , n64489 , n64490 , n64491 , n64492 , n64493 , n64494 , 
 n64495 , n64496 , n64497 , n64498 , n64499 , n64500 , n64501 , n64502 , n64503 , n64504 , 
 n64505 , n64506 , n64507 , n64508 , n64509 , n64510 , n64511 , n64512 , n64513 , n64514 , 
 n64515 , n64516 , n64517 , n64518 , n64519 , n64520 , n64521 , n64522 , n64523 , n64524 , 
 n64525 , n64526 , n64527 , n64528 , n64529 , n64530 , n64531 , n64532 , n64533 , n64534 , 
 n64535 , n64536 , n64537 , n64538 , n64539 , n64540 , n64541 , n64542 , n64543 , n64544 , 
 n64545 , n64546 , n64547 , n64548 , n64549 , n64550 , n64551 , n64552 , n64553 , n64554 , 
 n64555 , n64556 , n64557 , n64558 , n64559 , n64560 , n64561 , n64562 , n64563 , n64564 , 
 n64565 , n64566 , n64567 , n64568 , n64569 , n64570 , n64571 , n64572 , n64573 , n64574 , 
 n64575 , n64576 , n64577 , n64578 , n64579 , n64580 , n64581 , n64582 , n64583 , n64584 , 
 n64585 , n64586 , n64587 , n64588 , n64589 , n64590 , n64591 , n64592 , n64593 , n64594 , 
 n64595 , n64596 , n64597 , n64598 , n64599 , n64600 , n64601 , n64602 , n64603 , n64604 , 
 n64605 , n64606 , n64607 , n64608 , n64609 , n64610 , n64611 , n64612 , n64613 , n64614 , 
 n64615 , n64616 , n64617 , n64618 , n64619 , n64620 , n64621 , n64622 , n64623 , n64624 , 
 n64625 , n64626 , n64627 , n64628 , n64629 , n64630 , n64631 , n64632 , n64633 , n64634 , 
 n64635 , n64636 , n64637 , n64638 , n64639 , n64640 , n64641 , n64642 , n64643 , n64644 , 
 n64645 , n64646 , n64647 , n64648 , n64649 , n64650 , n64651 , n64652 , n64653 , n64654 , 
 n64655 , n64656 , n64657 , n64658 , n64659 , n64660 , n64661 , n64662 , n64663 , n64664 , 
 n64665 , n64666 , n64667 , n64668 , n64669 , n64670 , n64671 , n64672 , n64673 , n64674 , 
 n64675 , n64676 , n64677 , n64678 , n64679 , n64680 , n64681 , n64682 , n64683 , n64684 , 
 n64685 , n64686 , n64687 , n64688 , n64689 , n64690 , n64691 , n64692 , n64693 , n64694 , 
 n64695 , n64696 , n64697 , n64698 , n64699 , n64700 , n64701 , n64702 , n64703 , n64704 , 
 n64705 , n64706 , n64707 , n64708 , n64709 , n64710 , n64711 , n64712 , n64713 , n64714 , 
 n64715 , n64716 , n64717 , n64718 , n64719 , n64720 , n64721 , n64722 , n64723 , n64724 , 
 n64725 , n64726 , n64727 , n64728 , n64729 , n64730 , n64731 , n64732 , n64733 , n64734 , 
 n64735 , n64736 , n64737 , n64738 , n64739 , n64740 , n64741 , n64742 , n64743 , n64744 , 
 n64745 , n64746 , n64747 , n64748 , n64749 , n64750 , n64751 , n64752 , n64753 , n64754 , 
 n64755 , n64756 , n64757 , n64758 , n64759 , n64760 , n64761 , n64762 , n64763 , n64764 , 
 n64765 , n64766 , n64767 , n64768 , n64769 , n64770 , n64771 , n64772 , n64773 , n64774 , 
 n64775 , n64776 , n64777 , n64778 , n64779 , n64780 , n64781 , n64782 , n64783 , n64784 , 
 n64785 , n64786 , n64787 , n64788 , n64789 , n64790 , n64791 , n64792 , n64793 , n64794 , 
 n64795 , n64796 , n64797 , n64798 , n64799 , n64800 , n64801 , n64802 , n64803 , n64804 , 
 n64805 , n64806 , n64807 , n64808 , n64809 , n64810 , n64811 , n64812 , n64813 , n64814 , 
 n64815 , n64816 , n64817 , n64818 , n64819 , n64820 , n64821 , n64822 , n64823 , n64824 , 
 n64825 , n64826 , n64827 , n64828 , n64829 , n64830 , n64831 , n64832 , n64833 , n64834 , 
 n64835 , n64836 , n64837 , n64838 , n64839 , n64840 , n64841 , n64842 , n64843 , n64844 , 
 n64845 , n64846 , n64847 , n64848 , n64849 , n64850 , n64851 , n64852 , n64853 , n64854 , 
 n64855 , n64856 , n64857 , n64858 , n64859 , n64860 , n64861 , n64862 , n64863 , n64864 , 
 n64865 , n64866 , n64867 , n64868 , n64869 , n64870 , n64871 , n64872 , n64873 , n64874 , 
 n64875 , n64876 , n64877 , n64878 , n64879 , n64880 , n64881 , n64882 , n64883 , n64884 , 
 n64885 , n64886 , n64887 , n64888 , n64889 , n64890 , n64891 , n64892 , n64893 , n64894 , 
 n64895 , n64896 , n64897 , n64898 , n64899 , n64900 , n64901 , n64902 , n64903 , n64904 , 
 n64905 , n64906 , n64907 , n64908 , n64909 , n64910 , n64911 , n64912 , n64913 , n64914 , 
 n64915 , n64916 , n64917 , n64918 , n64919 , n64920 , n64921 , n64922 , n64923 , n64924 , 
 n64925 , n64926 , n64927 , n64928 , n64929 , n64930 , n64931 , n64932 , n64933 , n64934 , 
 n64935 , n64936 , n64937 , n64938 , n64939 , n64940 , n64941 , n64942 , n64943 , n64944 , 
 n64945 , n64946 , n64947 , n64948 , n64949 , n64950 , n64951 , n64952 , n64953 , n64954 , 
 n64955 , n64956 , n64957 , n64958 , n64959 , n64960 , n64961 , n64962 , n64963 , n64964 , 
 n64965 , n64966 , n64967 , n64968 , n64969 , n64970 , n64971 , n64972 , n64973 , n64974 , 
 n64975 , n64976 , n64977 , n64978 , n64979 , n64980 , n64981 , n64982 , n64983 , n64984 , 
 n64985 , n64986 , n64987 , n64988 , n64989 , n64990 , n64991 , n64992 , n64993 , n64994 , 
 n64995 , n64996 , n64997 , n64998 , n64999 , n65000 , n65001 , n65002 , n65003 , n65004 , 
 n65005 , n65006 , n65007 , n65008 , n65009 , n65010 , n65011 , n65012 , n65013 , n65014 , 
 n65015 , n65016 , n65017 , n65018 , n65019 , n65020 , n65021 , n65022 , n65023 , n65024 , 
 n65025 , n65026 , n65027 , n65028 , n65029 , n65030 , n65031 , n65032 , n65033 , n65034 , 
 n65035 , n65036 , n65037 , n65038 , n65039 , n65040 , n65041 , n65042 , n65043 , n65044 , 
 n65045 , n65046 , n65047 , n65048 , n65049 , n65050 , n65051 , n65052 , n65053 , n65054 , 
 n65055 , n65056 , n65057 , n65058 , n65059 , n65060 , n65061 , n65062 , n65063 , n65064 , 
 n65065 , n65066 , n65067 , n65068 , n65069 , n65070 , n65071 , n65072 , n65073 , n65074 , 
 n65075 , n65076 , n65077 , n65078 , n65079 , n65080 , n65081 , n65082 , n65083 , n65084 , 
 n65085 , n65086 , n65087 , n65088 , n65089 , n65090 , n65091 , n65092 , n65093 , n65094 , 
 n65095 , n65096 , n65097 , n65098 , n65099 , n65100 , n65101 , n65102 , n65103 , n65104 , 
 n65105 , n65106 , n65107 , n65108 , n65109 , n65110 , n65111 , n65112 , n65113 , n65114 , 
 n65115 , n65116 , n65117 , n65118 , n65119 , n65120 , n65121 , n65122 , n65123 , n65124 , 
 n65125 , n65126 , n65127 , n65128 , n65129 , n65130 , n65131 , n65132 , n65133 , n65134 , 
 n65135 , n65136 , n65137 , n65138 , n65139 , n65140 , n65141 , n65142 , n65143 , n65144 , 
 n65145 , n65146 , n65147 , n65148 , n65149 , n65150 , n65151 , n65152 , n65153 , n65154 , 
 n65155 , n65156 , n65157 , n65158 , n65159 , n65160 , n65161 , n65162 , n65163 , n65164 , 
 n65165 , n65166 , n65167 , n65168 , n65169 , n65170 , n65171 , n65172 , n65173 , n65174 , 
 n65175 , n65176 , n65177 , n65178 , n65179 , n65180 , n65181 , n65182 , n65183 , n65184 , 
 n65185 , n65186 , n65187 , n65188 , n65189 , n65190 , n65191 , n65192 , n65193 , n65194 , 
 n65195 , n65196 , n65197 , n65198 , n65199 , n65200 , n65201 , n65202 , n65203 , n65204 , 
 n65205 , n65206 , n65207 , n65208 , n65209 , n65210 , n65211 , n65212 , n65213 , n65214 , 
 n65215 , n65216 , n65217 , n65218 , n65219 , n65220 , n65221 , n65222 , n65223 , n65224 , 
 n65225 , n65226 , n65227 , n65228 , n65229 , n65230 , n65231 , n65232 , n65233 , n65234 , 
 n65235 , n65236 , n65237 , n65238 , n65239 , n65240 , n65241 , n65242 , n65243 , n65244 , 
 n65245 , n65246 , n65247 , n65248 , n65249 , n65250 , n65251 , n65252 , n65253 , n65254 , 
 n65255 , n65256 , n65257 , n65258 , n65259 , n65260 , n65261 , n65262 , n65263 , n65264 , 
 n65265 , n65266 , n65267 , n65268 , n65269 , n65270 , n65271 , n65272 , n65273 , n65274 , 
 n65275 , n65276 , n65277 , n65278 , n65279 , n65280 , n65281 , n65282 , n65283 , n65284 , 
 n65285 , n65286 , n65287 , n65288 , n65289 , n65290 , n65291 , n65292 , n65293 , n65294 , 
 n65295 , n65296 , n65297 , n65298 , n65299 , n65300 , n65301 , n65302 , n65303 , n65304 , 
 n65305 , n65306 , n65307 , n65308 , n65309 , n65310 , n65311 , n65312 , n65313 , n65314 , 
 n65315 , n65316 , n65317 , n65318 , n65319 , n65320 , n65321 , n65322 , n65323 , n65324 , 
 n65325 , n65326 , n65327 , n65328 , n65329 , n65330 , n65331 , n65332 , n65333 , n65334 , 
 n65335 , n65336 , n65337 , n65338 , n65339 , n65340 , n65341 , n65342 , n65343 , n65344 , 
 n65345 , n65346 , n65347 , n65348 , n65349 , n65350 , n65351 , n65352 , n65353 , n65354 , 
 n65355 , n65356 , n65357 , n65358 , n65359 , n65360 , n65361 , n65362 , n65363 , n65364 , 
 n65365 , n65366 , n65367 , n65368 , n65369 , n65370 , n65371 , n65372 , n65373 , n65374 , 
 n65375 , n65376 , n65377 , n65378 , n65379 , n65380 , n65381 , n65382 , n65383 , n65384 , 
 n65385 , n65386 , n65387 , n65388 , n65389 , n65390 , n65391 , n65392 , n65393 , n65394 , 
 n65395 , n65396 , n65397 , n65398 , n65399 , n65400 , n65401 , n65402 , n65403 , n65404 , 
 n65405 , n65406 , n65407 , n65408 , n65409 , n65410 , n65411 , n65412 , n65413 , n65414 , 
 n65415 , n65416 , n65417 , n65418 , n65419 , n65420 , n65421 , n65422 , n65423 , n65424 , 
 n65425 , n65426 , n65427 , n65428 , n65429 , n65430 , n65431 , n65432 , n65433 , n65434 , 
 n65435 , n65436 , n65437 , n65438 , n65439 , n65440 , n65441 , n65442 , n65443 , n65444 , 
 n65445 , n65446 , n65447 , n65448 , n65449 , n65450 , n65451 , n65452 , n65453 , n65454 , 
 n65455 , n65456 , n65457 , n65458 , n65459 , n65460 , n65461 , n65462 , n65463 , n65464 , 
 n65465 , n65466 , n65467 , n65468 , n65469 , n65470 , n65471 , n65472 , n65473 , n65474 , 
 n65475 , n65476 , n65477 , n65478 , n65479 , n65480 , n65481 , n65482 , n65483 , n65484 , 
 n65485 , n65486 , n65487 , n65488 , n65489 , n65490 , n65491 , n65492 , n65493 , n65494 , 
 n65495 , n65496 , n65497 , n65498 , n65499 , n65500 , n65501 , n65502 , n65503 , n65504 , 
 n65505 , n65506 , n65507 , n65508 , n65509 , n65510 , n65511 , n65512 , n65513 , n65514 , 
 n65515 , n65516 , n65517 , n65518 , n65519 , n65520 , n65521 , n65522 , n65523 , n65524 , 
 n65525 , n65526 , n65527 , n65528 , n65529 , n65530 , n65531 , n65532 , n65533 , n65534 , 
 n65535 , n65536 , n65537 , n65538 , n65539 , n65540 , n65541 , n65542 , n65543 , n65544 , 
 n65545 , n65546 , n65547 , n65548 , n65549 , n65550 , n65551 , n65552 , n65553 , n65554 , 
 n65555 , n65556 , n65557 , n65558 , n65559 , n65560 , n65561 , n65562 , n65563 , n65564 , 
 n65565 , n65566 , n65567 , n65568 , n65569 , n65570 , n65571 , n65572 , n65573 , n65574 , 
 n65575 , n65576 , n65577 , n65578 , n65579 , n65580 , n65581 , n65582 , n65583 , n65584 , 
 n65585 , n65586 , n65587 , n65588 , n65589 , n65590 , n65591 , n65592 , n65593 , n65594 , 
 n65595 , n65596 , n65597 , n65598 , n65599 , n65600 , n65601 , n65602 , n65603 , n65604 , 
 n65605 , n65606 , n65607 , n65608 , n65609 , n65610 , n65611 , n65612 , n65613 , n65614 , 
 n65615 , n65616 , n65617 , n65618 , n65619 , n65620 , n65621 , n65622 , n65623 , n65624 , 
 n65625 , n65626 , n65627 , n65628 , n65629 , n65630 , n65631 , n65632 , n65633 , n65634 , 
 n65635 , n65636 , n65637 , n65638 , n65639 , n65640 , n65641 , n65642 , n65643 , n65644 , 
 n65645 , n65646 , n65647 , n65648 , n65649 , n65650 , n65651 , n65652 , n65653 , n65654 , 
 n65655 , n65656 , n65657 , n65658 , n65659 , n65660 , n65661 , n65662 , n65663 , n65664 , 
 n65665 , n65666 , n65667 , n65668 , n65669 , n65670 , n65671 , n65672 , n65673 , n65674 , 
 n65675 , n65676 , n65677 , n65678 , n65679 , n65680 , n65681 , n65682 , n65683 , n65684 , 
 n65685 , n65686 , n65687 , n65688 , n65689 , n65690 , n65691 , n65692 , n65693 , n65694 , 
 n65695 , n65696 , n65697 , n65698 , n65699 , n65700 , n65701 , n65702 , n65703 , n65704 , 
 n65705 , n65706 , n65707 , n65708 , n65709 , n65710 , n65711 , n65712 , n65713 , n65714 , 
 n65715 , n65716 , n65717 , n65718 , n65719 , n65720 , n65721 , n65722 , n65723 , n65724 , 
 n65725 , n65726 , n65727 , n65728 , n65729 , n65730 , n65731 , n65732 , n65733 , n65734 , 
 n65735 , n65736 , n65737 , n65738 , n65739 , n65740 , n65741 , n65742 , n65743 , n65744 , 
 n65745 , n65746 , n65747 , n65748 , n65749 , n65750 , n65751 , n65752 , n65753 , n65754 , 
 n65755 , n65756 , n65757 , n65758 , n65759 , n65760 , n65761 , n65762 , n65763 , n65764 , 
 n65765 , n65766 , n65767 , n65768 , n65769 , n65770 , n65771 , n65772 , n65773 , n65774 , 
 n65775 , n65776 , n65777 , n65778 , n65779 , n65780 , n65781 , n65782 , n65783 , n65784 , 
 n65785 , n65786 , n65787 , n65788 , n65789 , n65790 , n65791 , n65792 , n65793 , n65794 , 
 n65795 , n65796 , n65797 , n65798 , n65799 , n65800 , n65801 , n65802 , n65803 , n65804 , 
 n65805 , n65806 , n65807 , n65808 , n65809 , n65810 , n65811 , n65812 , n65813 , n65814 , 
 n65815 , n65816 , n65817 , n65818 , n65819 , n65820 , n65821 , n65822 , n65823 , n65824 , 
 n65825 , n65826 , n65827 , n65828 , n65829 , n65830 , n65831 , n65832 , n65833 , n65834 , 
 n65835 , n65836 , n65837 , n65838 , n65839 , n65840 , n65841 , n65842 , n65843 , n65844 , 
 n65845 , n65846 , n65847 , n65848 , n65849 , n65850 , n65851 , n65852 , n65853 , n65854 , 
 n65855 , n65856 , n65857 , n65858 , n65859 , n65860 , n65861 , n65862 , n65863 , n65864 , 
 n65865 , n65866 , n65867 , n65868 , n65869 , n65870 , n65871 , n65872 , n65873 , n65874 , 
 n65875 , n65876 , n65877 , n65878 , n65879 , n65880 , n65881 , n65882 , n65883 , n65884 , 
 n65885 , n65886 , n65887 , n65888 , n65889 , n65890 , n65891 , n65892 , n65893 , n65894 , 
 n65895 , n65896 , n65897 , n65898 , n65899 , n65900 , n65901 , n65902 , n65903 , n65904 , 
 n65905 , n65906 , n65907 , n65908 , n65909 , n65910 , n65911 , n65912 , n65913 , n65914 , 
 n65915 , n65916 , n65917 , n65918 , n65919 , n65920 , n65921 , n65922 , n65923 , n65924 , 
 n65925 , n65926 , n65927 , n65928 , n65929 , n65930 , n65931 , n65932 , n65933 , n65934 , 
 n65935 , n65936 , n65937 , n65938 , n65939 , n65940 , n65941 , n65942 , n65943 , n65944 , 
 n65945 , n65946 , n65947 , n65948 , n65949 , n65950 , n65951 , n65952 , n65953 , n65954 , 
 n65955 , n65956 , n65957 , n65958 , n65959 , n65960 , n65961 , n65962 , n65963 , n65964 , 
 n65965 , n65966 , n65967 , n65968 , n65969 , n65970 , n65971 , n65972 , n65973 , n65974 , 
 n65975 , n65976 , n65977 , n65978 , n65979 , n65980 , n65981 , n65982 , n65983 , n65984 , 
 n65985 , n65986 , n65987 , n65988 , n65989 , n65990 , n65991 , n65992 , n65993 , n65994 , 
 n65995 , n65996 , n65997 , n65998 , n65999 , n66000 , n66001 , n66002 , n66003 , n66004 , 
 n66005 , n66006 , n66007 , n66008 , n66009 , n66010 , n66011 , n66012 , n66013 , n66014 , 
 n66015 , n66016 , n66017 , n66018 , n66019 , n66020 , n66021 , n66022 , n66023 , n66024 , 
 n66025 , n66026 , n66027 , n66028 , n66029 , n66030 , n66031 , n66032 , n66033 , n66034 , 
 n66035 , n66036 , n66037 , n66038 , n66039 , n66040 , n66041 , n66042 , n66043 , n66044 , 
 n66045 , n66046 , n66047 , n66048 , n66049 , n66050 , n66051 , n66052 , n66053 , n66054 , 
 n66055 , n66056 , n66057 , n66058 , n66059 , n66060 , n66061 , n66062 , n66063 , n66064 , 
 n66065 , n66066 , n66067 , n66068 , n66069 , n66070 , n66071 , n66072 , n66073 , n66074 , 
 n66075 , n66076 , n66077 , n66078 , n66079 , n66080 , n66081 , n66082 , n66083 , n66084 , 
 n66085 , n66086 , n66087 , n66088 , n66089 , n66090 , n66091 , n66092 , n66093 , n66094 , 
 n66095 , n66096 , n66097 , n66098 , n66099 , n66100 , n66101 , n66102 , n66103 , n66104 , 
 n66105 , n66106 , n66107 , n66108 , n66109 , n66110 , n66111 , n66112 , n66113 , n66114 , 
 n66115 , n66116 , n66117 , n66118 , n66119 , n66120 , n66121 , n66122 , n66123 , n66124 , 
 n66125 , n66126 , n66127 , n66128 , n66129 , n66130 , n66131 , n66132 , n66133 , n66134 , 
 n66135 , n66136 , n66137 , n66138 , n66139 , n66140 , n66141 , n66142 , n66143 , n66144 , 
 n66145 , n66146 , n66147 , n66148 , n66149 , n66150 , n66151 , n66152 , n66153 , n66154 , 
 n66155 , n66156 , n66157 , n66158 , n66159 , n66160 , n66161 , n66162 , n66163 , n66164 , 
 n66165 , n66166 , n66167 , n66168 , n66169 , n66170 , n66171 , n66172 , n66173 , n66174 , 
 n66175 , n66176 , n66177 , n66178 , n66179 , n66180 , n66181 , n66182 , n66183 , n66184 , 
 n66185 , n66186 , n66187 , n66188 , n66189 , n66190 , n66191 , n66192 , n66193 , n66194 , 
 n66195 , n66196 , n66197 , n66198 , n66199 , n66200 , n66201 , n66202 , n66203 , n66204 , 
 n66205 , n66206 , n66207 , n66208 , n66209 , n66210 , n66211 , n66212 , n66213 , n66214 , 
 n66215 , n66216 , n66217 , n66218 , n66219 , n66220 , n66221 , n66222 , n66223 , n66224 , 
 n66225 , n66226 , n66227 , n66228 , n66229 , n66230 , n66231 , n66232 , n66233 , n66234 , 
 n66235 , n66236 , n66237 , n66238 , n66239 , n66240 , n66241 , n66242 , n66243 , n66244 , 
 n66245 , n66246 , n66247 , n66248 , n66249 , n66250 , n66251 , n66252 , n66253 , n66254 , 
 n66255 , n66256 , n66257 , n66258 , n66259 , n66260 , n66261 , n66262 , n66263 , n66264 , 
 n66265 , n66266 , n66267 , n66268 , n66269 , n66270 , n66271 , n66272 , n66273 , n66274 , 
 n66275 , n66276 , n66277 , n66278 , n66279 , n66280 , n66281 , n66282 , n66283 , n66284 , 
 n66285 , n66286 , n66287 , n66288 , n66289 , n66290 , n66291 , n66292 , n66293 , n66294 , 
 n66295 , n66296 , n66297 , n66298 , n66299 , n66300 , n66301 , n66302 , n66303 , n66304 , 
 n66305 , n66306 , n66307 , n66308 , n66309 , n66310 , n66311 , n66312 , n66313 , n66314 , 
 n66315 , n66316 , n66317 , n66318 , n66319 , n66320 , n66321 , n66322 , n66323 , n66324 , 
 n66325 , n66326 , n66327 , n66328 , n66329 , n66330 , n66331 , n66332 , n66333 , n66334 , 
 n66335 , n66336 , n66337 , n66338 , n66339 , n66340 , n66341 , n66342 , n66343 , n66344 , 
 n66345 , n66346 , n66347 , n66348 , n66349 , n66350 , n66351 , n66352 , n66353 , n66354 , 
 n66355 , n66356 , n66357 , n66358 , n66359 , n66360 , n66361 , n66362 , n66363 , n66364 , 
 n66365 , n66366 , n66367 , n66368 , n66369 , n66370 , n66371 , n66372 , n66373 , n66374 , 
 n66375 , n66376 , n66377 , n66378 , n66379 , n66380 , n66381 , n66382 , n66383 , n66384 , 
 n66385 , n66386 , n66387 , n66388 , n66389 , n66390 , n66391 , n66392 , n66393 , n66394 , 
 n66395 , n66396 , n66397 , n66398 , n66399 , n66400 , n66401 , n66402 , n66403 , n66404 , 
 n66405 , n66406 , n66407 , n66408 , n66409 , n66410 , n66411 , n66412 , n66413 , n66414 , 
 n66415 , n66416 , n66417 , n66418 , n66419 , n66420 , n66421 , n66422 , n66423 , n66424 , 
 n66425 , n66426 , n66427 , n66428 , n66429 , n66430 , n66431 , n66432 , n66433 , n66434 , 
 n66435 , n66436 , n66437 , n66438 , n66439 , n66440 , n66441 , n66442 , n66443 , n66444 , 
 n66445 , n66446 , n66447 , n66448 , n66449 , n66450 , n66451 , n66452 , n66453 , n66454 , 
 n66455 , n66456 , n66457 , n66458 , n66459 , n66460 , n66461 , n66462 , n66463 , n66464 , 
 n66465 , n66466 , n66467 , n66468 , n66469 , n66470 , n66471 , n66472 , n66473 , n66474 , 
 n66475 , n66476 , n66477 , n66478 , n66479 , n66480 , n66481 , n66482 , n66483 , n66484 , 
 n66485 , n66486 , n66487 , n66488 , n66489 , n66490 , n66491 , n66492 , n66493 , n66494 , 
 n66495 , n66496 , n66497 , n66498 , n66499 , n66500 , n66501 , n66502 , n66503 , n66504 , 
 n66505 , n66506 , n66507 , n66508 , n66509 , n66510 , n66511 , n66512 , n66513 , n66514 , 
 n66515 , n66516 , n66517 , n66518 , n66519 , n66520 , n66521 , n66522 , n66523 , n66524 , 
 n66525 , n66526 , n66527 , n66528 , n66529 , n66530 , n66531 , n66532 , n66533 , n66534 , 
 n66535 , n66536 , n66537 , n66538 , n66539 , n66540 , n66541 , n66542 , n66543 , n66544 , 
 n66545 , n66546 , n66547 , n66548 , n66549 , n66550 , n66551 , n66552 , n66553 , n66554 , 
 n66555 , n66556 , n66557 , n66558 , n66559 , n66560 , n66561 , n66562 , n66563 , n66564 , 
 n66565 , n66566 , n66567 , n66568 , n66569 , n66570 , n66571 , n66572 , n66573 , n66574 , 
 n66575 , n66576 , n66577 , n66578 , n66579 , n66580 , n66581 , n66582 , n66583 , n66584 , 
 n66585 , n66586 , n66587 , n66588 , n66589 , n66590 , n66591 , n66592 , n66593 , n66594 , 
 n66595 , n66596 , n66597 , n66598 , n66599 , n66600 , n66601 , n66602 , n66603 , n66604 , 
 n66605 , n66606 , n66607 , n66608 , n66609 , n66610 , n66611 , n66612 , n66613 , n66614 , 
 n66615 , n66616 , n66617 , n66618 , n66619 , n66620 , n66621 , n66622 , n66623 , n66624 , 
 n66625 , n66626 , n66627 , n66628 , n66629 , n66630 , n66631 , n66632 , n66633 , n66634 , 
 n66635 , n66636 , n66637 , n66638 , n66639 , n66640 , n66641 , n66642 , n66643 , n66644 , 
 n66645 , n66646 , n66647 , n66648 , n66649 , n66650 , n66651 , n66652 , n66653 , n66654 , 
 n66655 , n66656 , n66657 , n66658 , n66659 , n66660 , n66661 , n66662 , n66663 , n66664 , 
 n66665 , n66666 , n66667 , n66668 , n66669 , n66670 , n66671 , n66672 , n66673 , n66674 , 
 n66675 , n66676 , n66677 , n66678 , n66679 , n66680 , n66681 , n66682 , n66683 , n66684 , 
 n66685 , n66686 , n66687 , n66688 , n66689 , n66690 , n66691 , n66692 , n66693 , n66694 , 
 n66695 , n66696 , n66697 , n66698 , n66699 , n66700 , n66701 , n66702 , n66703 , n66704 , 
 n66705 , n66706 , n66707 , n66708 , n66709 , n66710 , n66711 , n66712 , n66713 , n66714 , 
 n66715 , n66716 , n66717 , n66718 , n66719 , n66720 , n66721 , n66722 , n66723 , n66724 , 
 n66725 , n66726 , n66727 , n66728 , n66729 , n66730 , n66731 , n66732 , n66733 , n66734 , 
 n66735 , n66736 , n66737 , n66738 , n66739 , n66740 , n66741 , n66742 , n66743 , n66744 , 
 n66745 , n66746 , n66747 , n66748 , n66749 , n66750 , n66751 , n66752 , n66753 , n66754 , 
 n66755 , n66756 , n66757 , n66758 , n66759 , n66760 , n66761 , n66762 , n66763 , n66764 , 
 n66765 , n66766 , n66767 , n66768 , n66769 , n66770 , n66771 , n66772 , n66773 , n66774 , 
 n66775 , n66776 , n66777 , n66778 , n66779 , n66780 , n66781 , n66782 , n66783 , n66784 , 
 n66785 , n66786 , n66787 , n66788 , n66789 , n66790 , n66791 , n66792 , n66793 , n66794 , 
 n66795 , n66796 , n66797 , n66798 , n66799 , n66800 , n66801 , n66802 , n66803 , n66804 , 
 n66805 , n66806 , n66807 , n66808 , n66809 , n66810 , n66811 , n66812 , n66813 , n66814 , 
 n66815 , n66816 , n66817 , n66818 , n66819 , n66820 , n66821 , n66822 , n66823 , n66824 , 
 n66825 , n66826 , n66827 , n66828 , n66829 , n66830 , n66831 , n66832 , n66833 , n66834 , 
 n66835 , n66836 , n66837 , n66838 , n66839 , n66840 , n66841 , n66842 , n66843 , n66844 , 
 n66845 , n66846 , n66847 , n66848 , n66849 , n66850 , n66851 , n66852 , n66853 , n66854 , 
 n66855 , n66856 , n66857 , n66858 , n66859 , n66860 , n66861 , n66862 , n66863 , n66864 , 
 n66865 , n66866 , n66867 , n66868 , n66869 , n66870 , n66871 , n66872 , n66873 , n66874 , 
 n66875 , n66876 , n66877 , n66878 , n66879 , n66880 , n66881 , n66882 , n66883 , n66884 , 
 n66885 , n66886 , n66887 , n66888 , n66889 , n66890 , n66891 , n66892 , n66893 , n66894 , 
 n66895 , n66896 , n66897 , n66898 , n66899 , n66900 , n66901 , n66902 , n66903 , n66904 , 
 n66905 , n66906 , n66907 , n66908 , n66909 , n66910 , n66911 , n66912 , n66913 , n66914 , 
 n66915 , n66916 , n66917 , n66918 , n66919 , n66920 , n66921 , n66922 , n66923 , n66924 , 
 n66925 , n66926 , n66927 , n66928 , n66929 , n66930 , n66931 , n66932 , n66933 , n66934 , 
 n66935 , n66936 , n66937 , n66938 , n66939 , n66940 , n66941 , n66942 , n66943 , n66944 , 
 n66945 , n66946 , n66947 , n66948 , n66949 , n66950 , n66951 , n66952 , n66953 , n66954 , 
 n66955 , n66956 , n66957 , n66958 , n66959 , n66960 , n66961 , n66962 , n66963 , n66964 , 
 n66965 , n66966 , n66967 , n66968 , n66969 , n66970 , n66971 , n66972 , n66973 , n66974 , 
 n66975 , n66976 , n66977 , n66978 , n66979 , n66980 , n66981 , n66982 , n66983 , n66984 , 
 n66985 , n66986 , n66987 , n66988 , n66989 , n66990 , n66991 , n66992 , n66993 , n66994 , 
 n66995 , n66996 , n66997 , n66998 , n66999 , n67000 , n67001 , n67002 , n67003 , n67004 , 
 n67005 , n67006 , n67007 , n67008 , n67009 , n67010 , n67011 , n67012 , n67013 , n67014 , 
 n67015 , n67016 , n67017 , n67018 , n67019 , n67020 , n67021 , n67022 , n67023 , n67024 , 
 n67025 , n67026 , n67027 , n67028 , n67029 , n67030 , n67031 , n67032 , n67033 , n67034 , 
 n67035 , n67036 , n67037 , n67038 , n67039 , n67040 , n67041 , n67042 , n67043 , n67044 , 
 n67045 , n67046 , n67047 , n67048 , n67049 , n67050 , n67051 , n67052 , n67053 , n67054 , 
 n67055 , n67056 , n67057 , n67058 , n67059 , n67060 , n67061 , n67062 , n67063 , n67064 , 
 n67065 , n67066 , n67067 , n67068 , n67069 , n67070 , n67071 , n67072 , n67073 , n67074 , 
 n67075 , n67076 , n67077 , n67078 , n67079 , n67080 , n67081 , n67082 , n67083 , n67084 , 
 n67085 , n67086 , n67087 , n67088 , n67089 , n67090 , n67091 , n67092 , n67093 , n67094 , 
 n67095 , n67096 , n67097 , n67098 , n67099 , n67100 , n67101 , n67102 , n67103 , n67104 , 
 n67105 , n67106 , n67107 , n67108 , n67109 , n67110 , n67111 , n67112 , n67113 , n67114 , 
 n67115 , n67116 , n67117 , n67118 , n67119 , n67120 , n67121 , n67122 , n67123 , n67124 , 
 n67125 , n67126 , n67127 , n67128 , n67129 , n67130 , n67131 , n67132 , n67133 , n67134 , 
 n67135 , n67136 , n67137 , n67138 , n67139 , n67140 , n67141 , n67142 , n67143 , n67144 , 
 n67145 , n67146 , n67147 , n67148 , n67149 , n67150 , n67151 , n67152 , n67153 , n67154 , 
 n67155 , n67156 , n67157 , n67158 , n67159 , n67160 , n67161 , n67162 , n67163 , n67164 , 
 n67165 , n67166 , n67167 , n67168 , n67169 , n67170 , n67171 , n67172 , n67173 , n67174 , 
 n67175 , n67176 , n67177 , n67178 , n67179 , n67180 , n67181 , n67182 , n67183 , n67184 , 
 n67185 , n67186 , n67187 , n67188 , n67189 , n67190 , n67191 , n67192 , n67193 , n67194 , 
 n67195 , n67196 , n67197 , n67198 , n67199 , n67200 , n67201 , n67202 , n67203 , n67204 , 
 n67205 , n67206 , n67207 , n67208 , n67209 , n67210 , n67211 , n67212 , n67213 , n67214 , 
 n67215 , n67216 , n67217 , n67218 , n67219 , n67220 , n67221 , n67222 , n67223 , n67224 , 
 n67225 , n67226 , n67227 , n67228 , n67229 , n67230 , n67231 , n67232 , n67233 , n67234 , 
 n67235 , n67236 , n67237 , n67238 , n67239 , n67240 , n67241 , n67242 , n67243 , n67244 , 
 n67245 , n67246 , n67247 , n67248 , n67249 , n67250 , n67251 , n67252 , n67253 , n67254 , 
 n67255 , n67256 , n67257 , n67258 , n67259 , n67260 , n67261 , n67262 , n67263 , n67264 , 
 n67265 , n67266 , n67267 , n67268 , n67269 , n67270 , n67271 , n67272 , n67273 , n67274 , 
 n67275 , n67276 , n67277 , n67278 , n67279 , n67280 , n67281 , n67282 , n67283 , n67284 , 
 n67285 , n67286 , n67287 , n67288 , n67289 , n67290 , n67291 , n67292 , n67293 , n67294 , 
 n67295 , n67296 , n67297 , n67298 , n67299 , n67300 , n67301 , n67302 , n67303 , n67304 , 
 n67305 , n67306 , n67307 , n67308 , n67309 , n67310 , n67311 , n67312 , n67313 , n67314 , 
 n67315 , n67316 , n67317 , n67318 , n67319 , n67320 , n67321 , n67322 , n67323 , n67324 , 
 n67325 , n67326 , n67327 , n67328 , n67329 , n67330 , n67331 , n67332 , n67333 , n67334 , 
 n67335 , n67336 , n67337 , n67338 , n67339 , n67340 , n67341 , n67342 , n67343 , n67344 , 
 n67345 , n67346 , n67347 , n67348 , n67349 , n67350 , n67351 , n67352 , n67353 , n67354 , 
 n67355 , n67356 , n67357 , n67358 , n67359 , n67360 , n67361 , n67362 , n67363 , n67364 , 
 n67365 , n67366 , n67367 , n67368 , n67369 , n67370 , n67371 , n67372 , n67373 , n67374 , 
 n67375 , n67376 , n67377 , n67378 , n67379 , n67380 , n67381 , n67382 , n67383 , n67384 , 
 n67385 , n67386 , n67387 , n67388 , n67389 , n67390 , n67391 , n67392 , n67393 , n67394 , 
 n67395 , n67396 , n67397 , n67398 , n67399 , n67400 , n67401 , n67402 , n67403 , n67404 , 
 n67405 , n67406 , n67407 , n67408 , n67409 , n67410 , n67411 , n67412 , n67413 , n67414 , 
 n67415 , n67416 , n67417 , n67418 , n67419 , n67420 , n67421 , n67422 , n67423 , n67424 , 
 n67425 , n67426 , n67427 , n67428 , n67429 , n67430 , n67431 , n67432 , n67433 , n67434 , 
 n67435 , n67436 , n67437 , n67438 , n67439 , n67440 , n67441 , n67442 , n67443 , n67444 , 
 n67445 , n67446 , n67447 , n67448 , n67449 , n67450 , n67451 , n67452 , n67453 , n67454 , 
 n67455 , n67456 , n67457 , n67458 , n67459 , n67460 , n67461 , n67462 , n67463 , n67464 , 
 n67465 , n67466 , n67467 , n67468 , n67469 , n67470 , n67471 , n67472 , n67473 , n67474 , 
 n67475 , n67476 , n67477 , n67478 , n67479 , n67480 , n67481 , n67482 , n67483 , n67484 , 
 n67485 , n67486 , n67487 , n67488 , n67489 , n67490 , n67491 , n67492 , n67493 , n67494 , 
 n67495 , n67496 , n67497 , n67498 , n67499 , n67500 , n67501 , n67502 , n67503 , n67504 , 
 n67505 , n67506 , n67507 , n67508 , n67509 , n67510 , n67511 , n67512 , n67513 , n67514 , 
 n67515 , n67516 , n67517 , n67518 , n67519 , n67520 , n67521 , n67522 , n67523 , n67524 , 
 n67525 , n67526 , n67527 , n67528 , n67529 , n67530 , n67531 , n67532 , n67533 , n67534 , 
 n67535 , n67536 , n67537 , n67538 , n67539 , n67540 , n67541 , n67542 , n67543 , n67544 , 
 n67545 , n67546 , n67547 , n67548 , n67549 , n67550 , n67551 , n67552 , n67553 , n67554 , 
 n67555 , n67556 , n67557 , n67558 , n67559 , n67560 , n67561 , n67562 , n67563 , n67564 , 
 n67565 , n67566 , n67567 , n67568 , n67569 , n67570 , n67571 , n67572 , n67573 , n67574 , 
 n67575 , n67576 , n67577 , n67578 , n67579 , n67580 , n67581 , n67582 , n67583 , n67584 , 
 n67585 , n67586 , n67587 , n67588 , n67589 , n67590 , n67591 , n67592 , n67593 , n67594 , 
 n67595 , n67596 , n67597 , n67598 , n67599 , n67600 , n67601 , n67602 , n67603 , n67604 , 
 n67605 , n67606 , n67607 , n67608 , n67609 , n67610 , n67611 , n67612 , n67613 , n67614 , 
 n67615 , n67616 , n67617 , n67618 , n67619 , n67620 , n67621 , n67622 , n67623 , n67624 , 
 n67625 , n67626 , n67627 , n67628 , n67629 , n67630 , n67631 , n67632 , n67633 , n67634 , 
 n67635 , n67636 , n67637 , n67638 , n67639 , n67640 , n67641 , n67642 , n67643 , n67644 , 
 n67645 , n67646 , n67647 , n67648 , n67649 , n67650 , n67651 , n67652 , n67653 , n67654 , 
 n67655 , n67656 , n67657 , n67658 , n67659 , n67660 , n67661 , n67662 , n67663 , n67664 , 
 n67665 , n67666 , n67667 , n67668 , n67669 , n67670 , n67671 , n67672 , n67673 , n67674 , 
 n67675 , n67676 , n67677 , n67678 , n67679 , n67680 , n67681 , n67682 , n67683 , n67684 , 
 n67685 , n67686 , n67687 , n67688 , n67689 , n67690 , n67691 , n67692 , n67693 , n67694 , 
 n67695 , n67696 , n67697 , n67698 , n67699 , n67700 , n67701 , n67702 , n67703 , n67704 , 
 n67705 , n67706 , n67707 , n67708 , n67709 , n67710 , n67711 , n67712 , n67713 , n67714 , 
 n67715 , n67716 , n67717 , n67718 , n67719 , n67720 , n67721 , n67722 , n67723 , n67724 , 
 n67725 , n67726 , n67727 , n67728 , n67729 , n67730 , n67731 , n67732 , n67733 , n67734 , 
 n67735 , n67736 , n67737 , n67738 , n67739 , n67740 , n67741 , n67742 , n67743 , n67744 , 
 n67745 , n67746 , n67747 , n67748 , n67749 , n67750 , n67751 , n67752 , n67753 , n67754 , 
 n67755 , n67756 , n67757 , n67758 , n67759 , n67760 , n67761 , n67762 , n67763 , n67764 , 
 n67765 , n67766 , n67767 , n67768 , n67769 , n67770 , n67771 , n67772 , n67773 , n67774 , 
 n67775 , n67776 , n67777 , n67778 , n67779 , n67780 , n67781 , n67782 , n67783 , n67784 , 
 n67785 , n67786 , n67787 , n67788 , n67789 , n67790 , n67791 , n67792 , n67793 , n67794 , 
 n67795 , n67796 , n67797 , n67798 , n67799 , n67800 , n67801 , n67802 , n67803 , n67804 , 
 n67805 , n67806 , n67807 , n67808 , n67809 , n67810 , n67811 , n67812 , n67813 , n67814 , 
 n67815 , n67816 , n67817 , n67818 , n67819 , n67820 , n67821 , n67822 , n67823 , n67824 , 
 n67825 , n67826 , n67827 , n67828 , n67829 , n67830 , n67831 , n67832 , n67833 , n67834 , 
 n67835 , n67836 , n67837 , n67838 , n67839 , n67840 , n67841 , n67842 , n67843 , n67844 , 
 n67845 , n67846 , n67847 , n67848 , n67849 , n67850 , n67851 , n67852 , n67853 , n67854 , 
 n67855 , n67856 , n67857 , n67858 , n67859 , n67860 , n67861 , n67862 , n67863 , n67864 , 
 n67865 , n67866 , n67867 , n67868 , n67869 , n67870 , n67871 , n67872 , n67873 , n67874 , 
 n67875 , n67876 , n67877 , n67878 , n67879 , n67880 , n67881 , n67882 , n67883 , n67884 , 
 n67885 , n67886 , n67887 , n67888 , n67889 , n67890 , n67891 , n67892 , n67893 , n67894 , 
 n67895 , n67896 , n67897 , n67898 , n67899 , n67900 , n67901 , n67902 , n67903 , n67904 , 
 n67905 , n67906 , n67907 , n67908 , n67909 , n67910 , n67911 , n67912 , n67913 , n67914 , 
 n67915 , n67916 , n67917 , n67918 , n67919 , n67920 , n67921 , n67922 , n67923 , n67924 , 
 n67925 , n67926 , n67927 , n67928 , n67929 , n67930 , n67931 , n67932 , n67933 , n67934 , 
 n67935 , n67936 , n67937 , n67938 , n67939 , n67940 , n67941 , n67942 , n67943 , n67944 , 
 n67945 , n67946 , n67947 , n67948 , n67949 , n67950 , n67951 , n67952 , n67953 , n67954 , 
 n67955 , n67956 , n67957 , n67958 , n67959 , n67960 , n67961 , n67962 , n67963 , n67964 , 
 n67965 , n67966 , n67967 , n67968 , n67969 , n67970 , n67971 , n67972 , n67973 , n67974 , 
 n67975 , n67976 , n67977 , n67978 , n67979 , n67980 , n67981 , n67982 , n67983 , n67984 , 
 n67985 , n67986 , n67987 , n67988 , n67989 , n67990 , n67991 , n67992 , n67993 , n67994 , 
 n67995 , n67996 , n67997 , n67998 , n67999 , n68000 , n68001 , n68002 , n68003 , n68004 , 
 n68005 , n68006 , n68007 , n68008 , n68009 , n68010 , n68011 , n68012 , n68013 , n68014 , 
 n68015 , n68016 , n68017 , n68018 , n68019 , n68020 , n68021 , n68022 , n68023 , n68024 , 
 n68025 , n68026 , n68027 , n68028 , n68029 , n68030 , n68031 , n68032 , n68033 , n68034 , 
 n68035 , n68036 , n68037 , n68038 , n68039 , n68040 , n68041 , n68042 , n68043 , n68044 , 
 n68045 , n68046 , n68047 , n68048 , n68049 , n68050 , n68051 , n68052 , n68053 , n68054 , 
 n68055 , n68056 , n68057 , n68058 , n68059 , n68060 , n68061 , n68062 , n68063 , n68064 , 
 n68065 , n68066 , n68067 , n68068 , n68069 , n68070 , n68071 , n68072 , n68073 , n68074 , 
 n68075 , n68076 , n68077 , n68078 , n68079 , n68080 , n68081 , n68082 , n68083 , n68084 , 
 n68085 , n68086 , n68087 , n68088 , n68089 , n68090 , n68091 , n68092 , n68093 , n68094 , 
 n68095 , n68096 , n68097 , n68098 , n68099 , n68100 , n68101 , n68102 , n68103 , n68104 , 
 n68105 , n68106 , n68107 , n68108 , n68109 , n68110 , n68111 , n68112 , n68113 , n68114 , 
 n68115 , n68116 , n68117 , n68118 , n68119 , n68120 , n68121 , n68122 , n68123 , n68124 , 
 n68125 , n68126 , n68127 , n68128 , n68129 , n68130 , n68131 , n68132 , n68133 , n68134 , 
 n68135 , n68136 , n68137 , n68138 , n68139 , n68140 , n68141 , n68142 , n68143 , n68144 , 
 n68145 , n68146 , n68147 , n68148 , n68149 , n68150 , n68151 , n68152 , n68153 , n68154 , 
 n68155 , n68156 , n68157 , n68158 , n68159 , n68160 , n68161 , n68162 , n68163 , n68164 , 
 n68165 , n68166 , n68167 , n68168 , n68169 , n68170 , n68171 , n68172 , n68173 , n68174 , 
 n68175 , n68176 , n68177 , n68178 , n68179 , n68180 , n68181 , n68182 , n68183 , n68184 , 
 n68185 , n68186 , n68187 , n68188 , n68189 , n68190 , n68191 , n68192 , n68193 , n68194 , 
 n68195 , n68196 , n68197 , n68198 , n68199 , n68200 , n68201 , n68202 , n68203 , n68204 , 
 n68205 , n68206 , n68207 , n68208 , n68209 , n68210 , n68211 , n68212 , n68213 , n68214 , 
 n68215 , n68216 , n68217 , n68218 , n68219 , n68220 , n68221 , n68222 , n68223 , n68224 , 
 n68225 , n68226 , n68227 , n68228 , n68229 , n68230 , n68231 , n68232 , n68233 , n68234 , 
 n68235 , n68236 , n68237 , n68238 , n68239 , n68240 , n68241 , n68242 , n68243 , n68244 , 
 n68245 , n68246 , n68247 , n68248 , n68249 , n68250 , n68251 , n68252 , n68253 , n68254 , 
 n68255 , n68256 , n68257 , n68258 , n68259 , n68260 , n68261 , n68262 , n68263 , n68264 , 
 n68265 , n68266 , n68267 , n68268 , n68269 , n68270 , n68271 , n68272 , n68273 , n68274 , 
 n68275 , n68276 , n68277 , n68278 , n68279 , n68280 , n68281 , n68282 , n68283 , n68284 , 
 n68285 , n68286 , n68287 , n68288 , n68289 , n68290 , n68291 , n68292 , n68293 , n68294 , 
 n68295 , n68296 , n68297 , n68298 , n68299 , n68300 , n68301 , n68302 , n68303 , n68304 , 
 n68305 , n68306 , n68307 , n68308 , n68309 , n68310 , n68311 , n68312 , n68313 , n68314 , 
 n68315 , n68316 , n68317 , n68318 , n68319 , n68320 , n68321 , n68322 , n68323 , n68324 , 
 n68325 , n68326 , n68327 , n68328 , n68329 , n68330 , n68331 , n68332 , n68333 , n68334 , 
 n68335 , n68336 , n68337 , n68338 , n68339 , n68340 , n68341 , n68342 , n68343 , n68344 , 
 n68345 , n68346 , n68347 , n68348 , n68349 , n68350 , n68351 , n68352 , n68353 , n68354 , 
 n68355 , n68356 , n68357 , n68358 , n68359 , n68360 , n68361 , n68362 , n68363 , n68364 , 
 n68365 , n68366 , n68367 , n68368 , n68369 , n68370 , n68371 , n68372 , n68373 , n68374 , 
 n68375 , n68376 , n68377 , n68378 , n68379 , n68380 , n68381 , n68382 , n68383 , n68384 , 
 n68385 , n68386 , n68387 , n68388 , n68389 , n68390 , n68391 , n68392 , n68393 , n68394 , 
 n68395 , n68396 , n68397 , n68398 , n68399 , n68400 , n68401 , n68402 , n68403 , n68404 , 
 n68405 , n68406 , n68407 , n68408 , n68409 , n68410 , n68411 , n68412 , n68413 , n68414 , 
 n68415 , n68416 , n68417 , n68418 , n68419 , n68420 , n68421 , n68422 , n68423 , n68424 , 
 n68425 , n68426 , n68427 , n68428 , n68429 , n68430 , n68431 , n68432 , n68433 , n68434 , 
 n68435 , n68436 , n68437 , n68438 , n68439 , n68440 , n68441 , n68442 , n68443 , n68444 , 
 n68445 , n68446 , n68447 , n68448 , n68449 , n68450 , n68451 , n68452 , n68453 , n68454 , 
 n68455 , n68456 , n68457 , n68458 , n68459 , n68460 , n68461 , n68462 , n68463 , n68464 , 
 n68465 , n68466 , n68467 , n68468 , n68469 , n68470 , n68471 , n68472 , n68473 , n68474 , 
 n68475 , n68476 , n68477 , n68478 , n68479 , n68480 , n68481 , n68482 , n68483 , n68484 , 
 n68485 , n68486 , n68487 , n68488 , n68489 , n68490 , n68491 , n68492 , n68493 , n68494 , 
 n68495 , n68496 , n68497 , n68498 , n68499 , n68500 , n68501 , n68502 , n68503 , n68504 , 
 n68505 , n68506 , n68507 , n68508 , n68509 , n68510 , n68511 , n68512 , n68513 , n68514 , 
 n68515 , n68516 , n68517 , n68518 , n68519 , n68520 , n68521 , n68522 , n68523 , n68524 , 
 n68525 , n68526 , n68527 , n68528 , n68529 , n68530 , n68531 , n68532 , n68533 , n68534 , 
 n68535 , n68536 , n68537 , n68538 , n68539 , n68540 , n68541 , n68542 , n68543 , n68544 , 
 n68545 , n68546 , n68547 , n68548 , n68549 , n68550 , n68551 , n68552 , n68553 , n68554 , 
 n68555 , n68556 , n68557 , n68558 , n68559 , n68560 , n68561 , n68562 , n68563 , n68564 , 
 n68565 , n68566 , n68567 , n68568 , n68569 , n68570 , n68571 , n68572 , n68573 , n68574 , 
 n68575 , n68576 , n68577 , n68578 , n68579 , n68580 , n68581 , n68582 , n68583 , n68584 , 
 n68585 , n68586 , n68587 , n68588 , n68589 , n68590 , n68591 , n68592 , n68593 , n68594 , 
 n68595 , n68596 , n68597 , n68598 , n68599 , n68600 , n68601 , n68602 , n68603 , n68604 , 
 n68605 , n68606 , n68607 , n68608 , n68609 , n68610 , n68611 , n68612 , n68613 , n68614 , 
 n68615 , n68616 , n68617 , n68618 , n68619 , n68620 , n68621 , n68622 , n68623 , n68624 , 
 n68625 , n68626 , n68627 , n68628 , n68629 , n68630 , n68631 , n68632 , n68633 , n68634 , 
 n68635 , n68636 , n68637 , n68638 , n68639 , n68640 , n68641 , n68642 , n68643 , n68644 , 
 n68645 , n68646 , n68647 , n68648 , n68649 , n68650 , n68651 , n68652 , n68653 , n68654 , 
 n68655 , n68656 , n68657 , n68658 , n68659 , n68660 , n68661 , n68662 , n68663 , n68664 , 
 n68665 , n68666 , n68667 , n68668 , n68669 , n68670 , n68671 , n68672 , n68673 , n68674 , 
 n68675 , n68676 , n68677 , n68678 , n68679 , n68680 , n68681 , n68682 , n68683 , n68684 , 
 n68685 , n68686 , n68687 , n68688 , n68689 , n68690 , n68691 , n68692 , n68693 , n68694 , 
 n68695 , n68696 , n68697 , n68698 , n68699 , n68700 , n68701 , n68702 , n68703 , n68704 , 
 n68705 , n68706 , n68707 , n68708 , n68709 , n68710 , n68711 , n68712 , n68713 , n68714 , 
 n68715 , n68716 , n68717 , n68718 , n68719 , n68720 , n68721 , n68722 , n68723 , n68724 , 
 n68725 , n68726 , n68727 , n68728 , n68729 , n68730 , n68731 , n68732 , n68733 , n68734 , 
 n68735 , n68736 , n68737 , n68738 , n68739 , n68740 , n68741 , n68742 , n68743 , n68744 , 
 n68745 , n68746 , n68747 , n68748 , n68749 , n68750 , n68751 , n68752 , n68753 , n68754 , 
 n68755 , n68756 , n68757 , n68758 , n68759 , n68760 , n68761 , n68762 , n68763 , n68764 , 
 n68765 , n68766 , n68767 , n68768 , n68769 , n68770 , n68771 , n68772 , n68773 , n68774 , 
 n68775 , n68776 , n68777 , n68778 , n68779 , n68780 , n68781 , n68782 , n68783 , n68784 , 
 n68785 , n68786 , n68787 , n68788 , n68789 , n68790 , n68791 , n68792 , n68793 , n68794 , 
 n68795 , n68796 , n68797 , n68798 , n68799 , n68800 , n68801 , n68802 , n68803 , n68804 , 
 n68805 , n68806 , n68807 , n68808 , n68809 , n68810 , n68811 , n68812 , n68813 , n68814 , 
 n68815 , n68816 , n68817 , n68818 , n68819 , n68820 , n68821 , n68822 , n68823 , n68824 , 
 n68825 , n68826 , n68827 , n68828 , n68829 , n68830 , n68831 , n68832 , n68833 , n68834 , 
 n68835 , n68836 , n68837 , n68838 , n68839 , n68840 , n68841 , n68842 , n68843 , n68844 , 
 n68845 , n68846 , n68847 , n68848 , n68849 , n68850 , n68851 , n68852 , n68853 , n68854 , 
 n68855 , n68856 , n68857 , n68858 , n68859 , n68860 , n68861 , n68862 , n68863 , n68864 , 
 n68865 , n68866 , n68867 , n68868 , n68869 , n68870 , n68871 , n68872 , n68873 , n68874 , 
 n68875 , n68876 , n68877 , n68878 , n68879 , n68880 , n68881 , n68882 , n68883 , n68884 , 
 n68885 , n68886 , n68887 , n68888 , n68889 , n68890 , n68891 , n68892 , n68893 , n68894 , 
 n68895 , n68896 , n68897 , n68898 , n68899 , n68900 , n68901 , n68902 , n68903 , n68904 , 
 n68905 , n68906 , n68907 , n68908 , n68909 , n68910 , n68911 , n68912 , n68913 , n68914 , 
 n68915 , n68916 , n68917 , n68918 , n68919 , n68920 , n68921 , n68922 , n68923 , n68924 , 
 n68925 , n68926 , n68927 , n68928 , n68929 , n68930 , n68931 , n68932 , n68933 , n68934 , 
 n68935 , n68936 , n68937 , n68938 , n68939 , n68940 , n68941 , n68942 , n68943 , n68944 , 
 n68945 , n68946 , n68947 , n68948 , n68949 , n68950 , n68951 , n68952 , n68953 , n68954 , 
 n68955 , n68956 , n68957 , n68958 , n68959 , n68960 , n68961 , n68962 , n68963 , n68964 , 
 n68965 , n68966 , n68967 , n68968 , n68969 , n68970 , n68971 , n68972 , n68973 , n68974 , 
 n68975 , n68976 , n68977 , n68978 , n68979 , n68980 , n68981 , n68982 , n68983 , n68984 , 
 n68985 , n68986 , n68987 , n68988 , n68989 , n68990 , n68991 , n68992 , n68993 , n68994 , 
 n68995 , n68996 , n68997 , n68998 , n68999 , n69000 , n69001 , n69002 , n69003 , n69004 , 
 n69005 , n69006 , n69007 , n69008 , n69009 , n69010 , n69011 , n69012 , n69013 , n69014 , 
 n69015 , n69016 , n69017 , n69018 , n69019 , n69020 , n69021 , n69022 , n69023 , n69024 , 
 n69025 , n69026 , n69027 , n69028 , n69029 , n69030 , n69031 , n69032 , n69033 , n69034 , 
 n69035 , n69036 , n69037 , n69038 , n69039 , n69040 , n69041 , n69042 , n69043 , n69044 , 
 n69045 , n69046 , n69047 , n69048 , n69049 , n69050 , n69051 , n69052 , n69053 , n69054 , 
 n69055 , n69056 , n69057 , n69058 , n69059 , n69060 , n69061 , n69062 , n69063 , n69064 , 
 n69065 , n69066 , n69067 , n69068 , n69069 , n69070 , n69071 , n69072 , n69073 , n69074 , 
 n69075 , n69076 , n69077 , n69078 , n69079 , n69080 , n69081 , n69082 , n69083 , n69084 , 
 n69085 , n69086 , n69087 , n69088 , n69089 , n69090 , n69091 , n69092 , n69093 , n69094 , 
 n69095 , n69096 , n69097 , n69098 , n69099 , n69100 , n69101 , n69102 , n69103 , n69104 , 
 n69105 , n69106 , n69107 , n69108 , n69109 , n69110 , n69111 , n69112 , n69113 , n69114 , 
 n69115 , n69116 , n69117 , n69118 , n69119 , n69120 , n69121 , n69122 , n69123 , n69124 , 
 n69125 , n69126 , n69127 , n69128 , n69129 , n69130 , n69131 , n69132 , n69133 , n69134 , 
 n69135 , n69136 , n69137 , n69138 , n69139 , n69140 , n69141 , n69142 , n69143 , n69144 , 
 n69145 , n69146 , n69147 , n69148 , n69149 , n69150 , n69151 , n69152 , n69153 , n69154 , 
 n69155 , n69156 , n69157 , n69158 , n69159 , n69160 , n69161 , n69162 , n69163 , n69164 , 
 n69165 , n69166 , n69167 , n69168 , n69169 , n69170 , n69171 , n69172 , n69173 , n69174 , 
 n69175 , n69176 , n69177 , n69178 , n69179 , n69180 , n69181 , n69182 , n69183 , n69184 , 
 n69185 , n69186 , n69187 , n69188 , n69189 , n69190 , n69191 , n69192 , n69193 , n69194 , 
 n69195 , n69196 , n69197 , n69198 , n69199 , n69200 , n69201 , n69202 , n69203 , n69204 , 
 n69205 , n69206 , n69207 , n69208 , n69209 , n69210 , n69211 , n69212 , n69213 , n69214 , 
 n69215 , n69216 , n69217 , n69218 , n69219 , n69220 , n69221 , n69222 , n69223 , n69224 , 
 n69225 , n69226 , n69227 , n69228 , n69229 , n69230 , n69231 , n69232 , n69233 , n69234 , 
 n69235 , n69236 , n69237 , n69238 , n69239 , n69240 , n69241 , n69242 , n69243 , n69244 , 
 n69245 , n69246 , n69247 , n69248 , n69249 , n69250 , n69251 , n69252 , n69253 , n69254 , 
 n69255 , n69256 , n69257 , n69258 , n69259 , n69260 , n69261 , n69262 , n69263 , n69264 , 
 n69265 , n69266 , n69267 , n69268 , n69269 , n69270 , n69271 , n69272 , n69273 , n69274 , 
 n69275 , n69276 , n69277 , n69278 , n69279 , n69280 , n69281 , n69282 , n69283 , n69284 , 
 n69285 , n69286 , n69287 , n69288 , n69289 , n69290 , n69291 , n69292 , n69293 , n69294 , 
 n69295 , n69296 , n69297 , n69298 , n69299 , n69300 , n69301 , n69302 , n69303 , n69304 , 
 n69305 , n69306 , n69307 , n69308 , n69309 , n69310 , n69311 , n69312 , n69313 , n69314 , 
 n69315 , n69316 , n69317 , n69318 , n69319 , n69320 , n69321 , n69322 , n69323 , n69324 , 
 n69325 , n69326 , n69327 , n69328 , n69329 , n69330 , n69331 , n69332 , n69333 , n69334 , 
 n69335 , n69336 , n69337 , n69338 , n69339 , n69340 , n69341 , n69342 , n69343 , n69344 , 
 n69345 , n69346 , n69347 , n69348 , n69349 , n69350 , n69351 , n69352 , n69353 , n69354 , 
 n69355 , n69356 , n69357 , n69358 , n69359 , n69360 , n69361 , n69362 , n69363 , n69364 , 
 n69365 , n69366 , n69367 , n69368 , n69369 , n69370 , n69371 , n69372 , n69373 , n69374 , 
 n69375 , n69376 , n69377 , n69378 , n69379 , n69380 , n69381 , n69382 , n69383 , n69384 , 
 n69385 , n69386 , n69387 , n69388 , n69389 , n69390 , n69391 , n69392 , n69393 , n69394 , 
 n69395 , n69396 , n69397 , n69398 , n69399 , n69400 , n69401 , n69402 , n69403 , n69404 , 
 n69405 , n69406 , n69407 , n69408 , n69409 , n69410 , n69411 , n69412 , n69413 , n69414 , 
 n69415 , n69416 , n69417 , n69418 , n69419 , n69420 , n69421 , n69422 , n69423 , n69424 , 
 n69425 , n69426 , n69427 , n69428 , n69429 , n69430 , n69431 , n69432 , n69433 , n69434 , 
 n69435 , n69436 , n69437 , n69438 , n69439 , n69440 , n69441 , n69442 , n69443 , n69444 , 
 n69445 , n69446 , n69447 , n69448 , n69449 , n69450 , n69451 , n69452 , n69453 , n69454 , 
 n69455 , n69456 , n69457 , n69458 , n69459 , n69460 , n69461 , n69462 , n69463 , n69464 , 
 n69465 , n69466 , n69467 , n69468 , n69469 , n69470 , n69471 , n69472 , n69473 , n69474 , 
 n69475 , n69476 , n69477 , n69478 , n69479 , n69480 , n69481 , n69482 , n69483 , n69484 , 
 n69485 , n69486 , n69487 , n69488 , n69489 , n69490 , n69491 , n69492 , n69493 , n69494 , 
 n69495 , n69496 , n69497 , n69498 , n69499 , n69500 , n69501 , n69502 , n69503 , n69504 , 
 n69505 , n69506 , n69507 , n69508 , n69509 , n69510 , n69511 , n69512 , n69513 , n69514 , 
 n69515 , n69516 , n69517 , n69518 , n69519 , n69520 , n69521 , n69522 , n69523 , n69524 , 
 n69525 , n69526 , n69527 , n69528 , n69529 , n69530 , n69531 , n69532 , n69533 , n69534 , 
 n69535 , n69536 , n69537 , n69538 , n69539 , n69540 , n69541 , n69542 , n69543 , n69544 , 
 n69545 , n69546 , n69547 , n69548 , n69549 , n69550 , n69551 , n69552 , n69553 , n69554 , 
 n69555 , n69556 , n69557 , n69558 , n69559 , n69560 , n69561 , n69562 , n69563 , n69564 , 
 n69565 , n69566 , n69567 , n69568 , n69569 , n69570 , n69571 , n69572 , n69573 , n69574 , 
 n69575 , n69576 , n69577 , n69578 , n69579 , n69580 , n69581 , n69582 , n69583 , n69584 , 
 n69585 , n69586 , n69587 , n69588 , n69589 , n69590 , n69591 , n69592 , n69593 , n69594 , 
 n69595 , n69596 , n69597 , n69598 , n69599 , n69600 , n69601 , n69602 , n69603 , n69604 , 
 n69605 , n69606 , n69607 , n69608 , n69609 , n69610 , n69611 , n69612 , n69613 , n69614 , 
 n69615 , n69616 , n69617 , n69618 , n69619 , n69620 , n69621 , n69622 , n69623 , n69624 , 
 n69625 , n69626 , n69627 , n69628 , n69629 , n69630 , n69631 , n69632 , n69633 , n69634 , 
 n69635 , n69636 , n69637 , n69638 , n69639 , n69640 , n69641 , n69642 , n69643 , n69644 , 
 n69645 , n69646 , n69647 , n69648 , n69649 , n69650 , n69651 , n69652 , n69653 , n69654 , 
 n69655 , n69656 , n69657 , n69658 , n69659 , n69660 , n69661 , n69662 , n69663 , n69664 , 
 n69665 , n69666 , n69667 , n69668 , n69669 , n69670 , n69671 , n69672 , n69673 , n69674 , 
 n69675 , n69676 , n69677 , n69678 , n69679 , n69680 , n69681 , n69682 , n69683 , n69684 , 
 n69685 , n69686 , n69687 , n69688 , n69689 , n69690 , n69691 , n69692 , n69693 , n69694 , 
 n69695 , n69696 , n69697 , n69698 , n69699 , n69700 , n69701 , n69702 , n69703 , n69704 , 
 n69705 , n69706 , n69707 , n69708 , n69709 , n69710 , n69711 , n69712 , n69713 , n69714 , 
 n69715 , n69716 , n69717 , n69718 , n69719 , n69720 , n69721 , n69722 , n69723 , n69724 , 
 n69725 , n69726 , n69727 , n69728 , n69729 , n69730 , n69731 , n69732 , n69733 , n69734 , 
 n69735 , n69736 , n69737 , n69738 , n69739 , n69740 , n69741 , n69742 , n69743 , n69744 , 
 n69745 , n69746 , n69747 , n69748 , n69749 , n69750 , n69751 , n69752 , n69753 , n69754 , 
 n69755 , n69756 , n69757 , n69758 , n69759 , n69760 , n69761 , n69762 , n69763 , n69764 , 
 n69765 , n69766 , n69767 , n69768 , n69769 , n69770 , n69771 , n69772 , n69773 , n69774 , 
 n69775 , n69776 , n69777 , n69778 , n69779 , n69780 , n69781 , n69782 , n69783 , n69784 , 
 n69785 , n69786 , n69787 , n69788 , n69789 , n69790 , n69791 , n69792 , n69793 , n69794 , 
 n69795 , n69796 , n69797 , n69798 , n69799 , n69800 , n69801 , n69802 , n69803 , n69804 , 
 n69805 , n69806 , n69807 , n69808 , n69809 , n69810 , n69811 , n69812 , n69813 , n69814 , 
 n69815 , n69816 , n69817 , n69818 , n69819 , n69820 , n69821 , n69822 , n69823 , n69824 , 
 n69825 , n69826 , n69827 , n69828 , n69829 , n69830 , n69831 , n69832 , n69833 , n69834 , 
 n69835 , n69836 , n69837 , n69838 , n69839 , n69840 , n69841 , n69842 , n69843 , n69844 , 
 n69845 , n69846 , n69847 , n69848 , n69849 , n69850 , n69851 , n69852 , n69853 , n69854 , 
 n69855 , n69856 , n69857 , n69858 , n69859 , n69860 , n69861 , n69862 , n69863 , n69864 , 
 n69865 , n69866 , n69867 , n69868 , n69869 , n69870 , n69871 , n69872 , n69873 , n69874 , 
 n69875 , n69876 , n69877 , n69878 , n69879 , n69880 , n69881 , n69882 , n69883 , n69884 , 
 n69885 , n69886 , n69887 , n69888 , n69889 , n69890 , n69891 , n69892 , n69893 , n69894 , 
 n69895 , n69896 , n69897 , n69898 , n69899 , n69900 , n69901 , n69902 , n69903 , n69904 , 
 n69905 , n69906 , n69907 , n69908 , n69909 , n69910 , n69911 , n69912 , n69913 , n69914 , 
 n69915 , n69916 , n69917 , n69918 , n69919 , n69920 , n69921 , n69922 , n69923 , n69924 , 
 n69925 , n69926 , n69927 , n69928 , n69929 , n69930 , n69931 , n69932 , n69933 , n69934 , 
 n69935 , n69936 , n69937 , n69938 , n69939 , n69940 , n69941 , n69942 , n69943 , n69944 , 
 n69945 , n69946 , n69947 , n69948 , n69949 , n69950 , n69951 , n69952 , n69953 , n69954 , 
 n69955 , n69956 , n69957 , n69958 , n69959 , n69960 , n69961 , n69962 , n69963 , n69964 , 
 n69965 , n69966 , n69967 , n69968 , n69969 , n69970 , n69971 , n69972 , n69973 , n69974 , 
 n69975 , n69976 , n69977 , n69978 , n69979 , n69980 , n69981 , n69982 , n69983 , n69984 , 
 n69985 , n69986 , n69987 , n69988 , n69989 , n69990 , n69991 , n69992 , n69993 , n69994 , 
 n69995 , n69996 , n69997 , n69998 , n69999 , n70000 , n70001 , n70002 , n70003 , n70004 , 
 n70005 , n70006 , n70007 , n70008 , n70009 , n70010 , n70011 , n70012 , n70013 , n70014 , 
 n70015 , n70016 , n70017 , n70018 , n70019 , n70020 , n70021 , n70022 , n70023 , n70024 , 
 n70025 , n70026 , n70027 , n70028 , n70029 , n70030 , n70031 , n70032 , n70033 , n70034 , 
 n70035 , n70036 , n70037 , n70038 , n70039 , n70040 , n70041 , n70042 , n70043 , n70044 , 
 n70045 , n70046 , n70047 , n70048 , n70049 , n70050 , n70051 , n70052 , n70053 , n70054 , 
 n70055 , n70056 , n70057 , n70058 , n70059 , n70060 , n70061 , n70062 , n70063 , n70064 , 
 n70065 , n70066 , n70067 , n70068 , n70069 , n70070 , n70071 , n70072 , n70073 , n70074 , 
 n70075 , n70076 , n70077 , n70078 , n70079 , n70080 , n70081 , n70082 , n70083 , n70084 , 
 n70085 , n70086 , n70087 , n70088 , n70089 , n70090 , n70091 , n70092 , n70093 , n70094 , 
 n70095 , n70096 , n70097 , n70098 , n70099 , n70100 , n70101 , n70102 , n70103 , n70104 , 
 n70105 , n70106 , n70107 , n70108 , n70109 , n70110 , n70111 , n70112 , n70113 , n70114 , 
 n70115 , n70116 , n70117 , n70118 , n70119 , n70120 , n70121 , n70122 , n70123 , n70124 , 
 n70125 , n70126 , n70127 , n70128 , n70129 , n70130 , n70131 , n70132 , n70133 , n70134 , 
 n70135 , n70136 , n70137 , n70138 , n70139 , n70140 , n70141 , n70142 , n70143 , n70144 , 
 n70145 , n70146 , n70147 , n70148 , n70149 , n70150 , n70151 , n70152 , n70153 , n70154 , 
 n70155 , n70156 , n70157 , n70158 , n70159 , n70160 , n70161 , n70162 , n70163 , n70164 , 
 n70165 , n70166 , n70167 , n70168 , n70169 , n70170 , n70171 , n70172 , n70173 , n70174 , 
 n70175 , n70176 , n70177 , n70178 , n70179 , n70180 , n70181 , n70182 , n70183 , n70184 , 
 n70185 , n70186 , n70187 , n70188 , n70189 , n70190 , n70191 , n70192 , n70193 , n70194 , 
 n70195 , n70196 , n70197 , n70198 , n70199 , n70200 , n70201 , n70202 , n70203 , n70204 , 
 n70205 , n70206 , n70207 , n70208 , n70209 , n70210 , n70211 , n70212 , n70213 , n70214 , 
 n70215 , n70216 , n70217 , n70218 , n70219 , n70220 , n70221 , n70222 , n70223 , n70224 , 
 n70225 , n70226 , n70227 , n70228 , n70229 , n70230 , n70231 , n70232 , n70233 , n70234 , 
 n70235 , n70236 , n70237 , n70238 , n70239 , n70240 , n70241 , n70242 , n70243 , n70244 , 
 n70245 , n70246 , n70247 , n70248 , n70249 , n70250 , n70251 , n70252 , n70253 , n70254 , 
 n70255 , n70256 , n70257 , n70258 , n70259 , n70260 , n70261 , n70262 , n70263 , n70264 , 
 n70265 , n70266 , n70267 , n70268 , n70269 , n70270 , n70271 , n70272 , n70273 , n70274 , 
 n70275 , n70276 , n70277 , n70278 , n70279 , n70280 , n70281 , n70282 , n70283 , n70284 , 
 n70285 , n70286 , n70287 , n70288 , n70289 , n70290 , n70291 , n70292 , n70293 , n70294 , 
 n70295 , n70296 , n70297 , n70298 , n70299 , n70300 , n70301 , n70302 , n70303 , n70304 , 
 n70305 , n70306 , n70307 , n70308 , n70309 , n70310 , n70311 , n70312 , n70313 , n70314 , 
 n70315 , n70316 , n70317 , n70318 , n70319 , n70320 , n70321 , n70322 , n70323 , n70324 , 
 n70325 , n70326 , n70327 , n70328 , n70329 , n70330 , n70331 , n70332 , n70333 , n70334 , 
 n70335 , n70336 , n70337 , n70338 , n70339 , n70340 , n70341 , n70342 , n70343 , n70344 , 
 n70345 , n70346 , n70347 , n70348 , n70349 , n70350 , n70351 , n70352 , n70353 , n70354 , 
 n70355 , n70356 , n70357 , n70358 , n70359 , n70360 , n70361 , n70362 , n70363 , n70364 , 
 n70365 , n70366 , n70367 , n70368 , n70369 , n70370 , n70371 , n70372 , n70373 , n70374 , 
 n70375 , n70376 , n70377 , n70378 , n70379 , n70380 , n70381 , n70382 , n70383 , n70384 , 
 n70385 , n70386 , n70387 , n70388 , n70389 , n70390 , n70391 , n70392 , n70393 , n70394 , 
 n70395 , n70396 , n70397 , n70398 , n70399 , n70400 , n70401 , n70402 , n70403 , n70404 , 
 n70405 , n70406 , n70407 , n70408 , n70409 , n70410 , n70411 , n70412 , n70413 , n70414 , 
 n70415 , n70416 , n70417 , n70418 , n70419 , n70420 , n70421 , n70422 , n70423 , n70424 , 
 n70425 , n70426 , n70427 , n70428 , n70429 , n70430 , n70431 , n70432 , n70433 , n70434 , 
 n70435 , n70436 , n70437 , n70438 , n70439 , n70440 , n70441 , n70442 , n70443 , n70444 , 
 n70445 , n70446 , n70447 , n70448 , n70449 , n70450 , n70451 , n70452 , n70453 , n70454 , 
 n70455 , n70456 , n70457 , n70458 , n70459 , n70460 , n70461 , n70462 , n70463 , n70464 , 
 n70465 , n70466 , n70467 , n70468 , n70469 , n70470 , n70471 , n70472 , n70473 , n70474 , 
 n70475 , n70476 , n70477 , n70478 , n70479 , n70480 , n70481 , n70482 , n70483 , n70484 , 
 n70485 , n70486 , n70487 , n70488 , n70489 , n70490 , n70491 , n70492 , n70493 , n70494 , 
 n70495 , n70496 , n70497 , n70498 , n70499 , n70500 , n70501 , n70502 , n70503 , n70504 , 
 n70505 , n70506 , n70507 , n70508 , n70509 , n70510 , n70511 , n70512 , n70513 , n70514 , 
 n70515 , n70516 , n70517 , n70518 , n70519 , n70520 , n70521 , n70522 , n70523 , n70524 , 
 n70525 , n70526 , n70527 , n70528 , n70529 , n70530 , n70531 , n70532 , n70533 , n70534 , 
 n70535 , n70536 , n70537 , n70538 , n70539 , n70540 , n70541 , n70542 , n70543 , n70544 , 
 n70545 , n70546 , n70547 , n70548 , n70549 , n70550 , n70551 , n70552 , n70553 , n70554 , 
 n70555 , n70556 , n70557 , n70558 , n70559 , n70560 , n70561 , n70562 , n70563 , n70564 , 
 n70565 , n70566 , n70567 , n70568 , n70569 , n70570 , n70571 , n70572 , n70573 , n70574 , 
 n70575 , n70576 , n70577 , n70578 , n70579 , n70580 , n70581 , n70582 , n70583 , n70584 , 
 n70585 , n70586 , n70587 , n70588 , n70589 , n70590 , n70591 , n70592 , n70593 , n70594 , 
 n70595 , n70596 , n70597 , n70598 , n70599 , n70600 , n70601 , n70602 , n70603 , n70604 , 
 n70605 , n70606 , n70607 , n70608 , n70609 , n70610 , n70611 , n70612 , n70613 , n70614 , 
 n70615 , n70616 , n70617 , n70618 , n70619 , n70620 , n70621 , n70622 , n70623 , n70624 , 
 n70625 , n70626 , n70627 , n70628 , n70629 , n70630 , n70631 , n70632 , n70633 , n70634 , 
 n70635 , n70636 , n70637 , n70638 , n70639 , n70640 , n70641 , n70642 , n70643 , n70644 , 
 n70645 , n70646 , n70647 , n70648 , n70649 , n70650 , n70651 , n70652 , n70653 , n70654 , 
 n70655 , n70656 , n70657 , n70658 , n70659 , n70660 , n70661 , n70662 , n70663 , n70664 , 
 n70665 , n70666 , n70667 , n70668 , n70669 , n70670 , n70671 , n70672 , n70673 , n70674 , 
 n70675 , n70676 , n70677 , n70678 , n70679 , n70680 , n70681 , n70682 , n70683 , n70684 , 
 n70685 , n70686 , n70687 , n70688 , n70689 , n70690 , n70691 , n70692 , n70693 , n70694 , 
 n70695 , n70696 , n70697 , n70698 , n70699 , n70700 , n70701 , n70702 , n70703 , n70704 , 
 n70705 , n70706 , n70707 , n70708 , n70709 , n70710 , n70711 , n70712 , n70713 , n70714 , 
 n70715 , n70716 , n70717 , n70718 , n70719 , n70720 , n70721 , n70722 , n70723 , n70724 , 
 n70725 , n70726 , n70727 , n70728 , n70729 , n70730 , n70731 , n70732 , n70733 , n70734 , 
 n70735 , n70736 , n70737 , n70738 , n70739 , n70740 , n70741 , n70742 , n70743 , n70744 , 
 n70745 , n70746 , n70747 , n70748 , n70749 , n70750 , n70751 , n70752 , n70753 , n70754 , 
 n70755 , n70756 , n70757 , n70758 , n70759 , n70760 , n70761 , n70762 , n70763 , n70764 , 
 n70765 , n70766 , n70767 , n70768 , n70769 , n70770 , n70771 , n70772 , n70773 , n70774 , 
 n70775 , n70776 , n70777 , n70778 , n70779 , n70780 , n70781 , n70782 , n70783 , n70784 , 
 n70785 , n70786 , n70787 , n70788 , n70789 , n70790 , n70791 , n70792 , n70793 , n70794 , 
 n70795 , n70796 , n70797 , n70798 , n70799 , n70800 , n70801 , n70802 , n70803 , n70804 , 
 n70805 , n70806 , n70807 , n70808 , n70809 , n70810 , n70811 , n70812 , n70813 , n70814 , 
 n70815 , n70816 , n70817 , n70818 , n70819 , n70820 , n70821 , n70822 , n70823 , n70824 , 
 n70825 , n70826 , n70827 , n70828 , n70829 , n70830 , n70831 , n70832 , n70833 , n70834 , 
 n70835 , n70836 , n70837 , n70838 , n70839 , n70840 , n70841 , n70842 , n70843 , n70844 , 
 n70845 , n70846 , n70847 , n70848 , n70849 , n70850 , n70851 , n70852 , n70853 , n70854 , 
 n70855 , n70856 , n70857 , n70858 , n70859 , n70860 , n70861 , n70862 , n70863 , n70864 , 
 n70865 , n70866 , n70867 , n70868 , n70869 , n70870 , n70871 , n70872 , n70873 , n70874 , 
 n70875 , n70876 , n70877 , n70878 , n70879 , n70880 , n70881 , n70882 , n70883 , n70884 , 
 n70885 , n70886 , n70887 , n70888 , n70889 , n70890 , n70891 , n70892 , n70893 , n70894 , 
 n70895 , n70896 , n70897 , n70898 , n70899 , n70900 , n70901 , n70902 , n70903 , n70904 , 
 n70905 , n70906 , n70907 , n70908 , n70909 , n70910 , n70911 , n70912 , n70913 , n70914 , 
 n70915 , n70916 , n70917 , n70918 , n70919 , n70920 , n70921 , n70922 , n70923 , n70924 , 
 n70925 , n70926 , n70927 , n70928 , n70929 , n70930 , n70931 , n70932 , n70933 , n70934 , 
 n70935 , n70936 , n70937 , n70938 , n70939 , n70940 , n70941 , n70942 , n70943 , n70944 , 
 n70945 , n70946 , n70947 , n70948 , n70949 , n70950 , n70951 , n70952 , n70953 , n70954 , 
 n70955 , n70956 , n70957 , n70958 , n70959 , n70960 , n70961 , n70962 , n70963 , n70964 , 
 n70965 , n70966 , n70967 , n70968 , n70969 , n70970 , n70971 , n70972 , n70973 , n70974 , 
 n70975 , n70976 , n70977 , n70978 , n70979 , n70980 , n70981 , n70982 , n70983 , n70984 , 
 n70985 , n70986 , n70987 , n70988 , n70989 , n70990 , n70991 , n70992 , n70993 , n70994 , 
 n70995 , n70996 , n70997 , n70998 , n70999 , n71000 , n71001 , n71002 , n71003 , n71004 , 
 n71005 , n71006 , n71007 , n71008 , n71009 , n71010 , n71011 , n71012 , n71013 , n71014 , 
 n71015 , n71016 , n71017 , n71018 , n71019 , n71020 , n71021 , n71022 , n71023 , n71024 , 
 n71025 , n71026 , n71027 , n71028 , n71029 , n71030 , n71031 , n71032 , n71033 , n71034 , 
 n71035 , n71036 , n71037 , n71038 , n71039 , n71040 , n71041 , n71042 , n71043 , n71044 , 
 n71045 , n71046 , n71047 , n71048 , n71049 , n71050 , n71051 , n71052 , n71053 , n71054 , 
 n71055 , n71056 , n71057 , n71058 , n71059 , n71060 , n71061 , n71062 , n71063 , n71064 , 
 n71065 , n71066 , n71067 , n71068 , n71069 , n71070 , n71071 , n71072 , n71073 , n71074 , 
 n71075 , n71076 , n71077 , n71078 , n71079 , n71080 , n71081 , n71082 , n71083 , n71084 , 
 n71085 , n71086 , n71087 , n71088 , n71089 , n71090 , n71091 , n71092 , n71093 , n71094 , 
 n71095 , n71096 , n71097 , n71098 , n71099 , n71100 , n71101 , n71102 , n71103 , n71104 , 
 n71105 , n71106 , n71107 , n71108 , n71109 , n71110 , n71111 , n71112 , n71113 , n71114 , 
 n71115 , n71116 , n71117 , n71118 , n71119 , n71120 , n71121 , n71122 , n71123 , n71124 , 
 n71125 , n71126 , n71127 , n71128 , n71129 , n71130 , n71131 , n71132 , n71133 , n71134 , 
 n71135 , n71136 , n71137 , n71138 , n71139 , n71140 , n71141 , n71142 , n71143 , n71144 , 
 n71145 , n71146 , n71147 , n71148 , n71149 , n71150 , n71151 , n71152 , n71153 , n71154 , 
 n71155 , n71156 , n71157 , n71158 , n71159 , n71160 , n71161 , n71162 , n71163 , n71164 , 
 n71165 , n71166 , n71167 , n71168 , n71169 , n71170 , n71171 , n71172 , n71173 , n71174 , 
 n71175 , n71176 , n71177 , n71178 , n71179 , n71180 , n71181 , n71182 , n71183 , n71184 , 
 n71185 , n71186 , n71187 , n71188 , n71189 , n71190 , n71191 , n71192 , n71193 , n71194 , 
 n71195 , n71196 , n71197 , n71198 , n71199 , n71200 , n71201 , n71202 , n71203 , n71204 , 
 n71205 , n71206 , n71207 , n71208 , n71209 , n71210 , n71211 , n71212 , n71213 , n71214 , 
 n71215 , n71216 , n71217 , n71218 , n71219 , n71220 , n71221 , n71222 , n71223 , n71224 , 
 n71225 , n71226 , n71227 , n71228 , n71229 , n71230 , n71231 , n71232 , n71233 , n71234 , 
 n71235 , n71236 , n71237 , n71238 , n71239 , n71240 , n71241 , n71242 , n71243 , n71244 , 
 n71245 , n71246 , n71247 , n71248 , n71249 , n71250 , n71251 , n71252 , n71253 , n71254 , 
 n71255 , n71256 , n71257 , n71258 , n71259 , n71260 , n71261 , n71262 , n71263 , n71264 , 
 n71265 , n71266 , n71267 , n71268 , n71269 , n71270 , n71271 , n71272 , n71273 , n71274 , 
 n71275 , n71276 , n71277 , n71278 , n71279 , n71280 , n71281 , n71282 , n71283 , n71284 , 
 n71285 , n71286 , n71287 , n71288 , n71289 , n71290 , n71291 , n71292 , n71293 , n71294 , 
 n71295 , n71296 , n71297 , n71298 , n71299 , n71300 , n71301 , n71302 , n71303 , n71304 , 
 n71305 , n71306 , n71307 , n71308 , n71309 , n71310 , n71311 , n71312 , n71313 , n71314 , 
 n71315 , n71316 , n71317 , n71318 , n71319 , n71320 , n71321 , n71322 , n71323 , n71324 , 
 n71325 , n71326 , n71327 , n71328 , n71329 , n71330 , n71331 , n71332 , n71333 , n71334 , 
 n71335 , n71336 , n71337 , n71338 , n71339 , n71340 , n71341 , n71342 , n71343 , n71344 , 
 n71345 , n71346 , n71347 , n71348 , n71349 , n71350 , n71351 , n71352 , n71353 , n71354 , 
 n71355 , n71356 , n71357 , n71358 , n71359 , n71360 , n71361 , n71362 , n71363 , n71364 , 
 n71365 , n71366 , n71367 , n71368 , n71369 , n71370 , n71371 , n71372 , n71373 , n71374 , 
 n71375 , n71376 , n71377 , n71378 , n71379 , n71380 , n71381 , n71382 , n71383 , n71384 , 
 n71385 , n71386 , n71387 , n71388 , n71389 , n71390 , n71391 , n71392 , n71393 , n71394 , 
 n71395 , n71396 , n71397 , n71398 , n71399 , n71400 , n71401 , n71402 , n71403 , n71404 , 
 n71405 , n71406 , n71407 , n71408 , n71409 , n71410 , n71411 , n71412 , n71413 , n71414 , 
 n71415 , n71416 , n71417 , n71418 , n71419 , n71420 , n71421 , n71422 , n71423 , n71424 , 
 n71425 , n71426 , n71427 , n71428 , n71429 , n71430 , n71431 , n71432 , n71433 , n71434 , 
 n71435 , n71436 , n71437 , n71438 , n71439 , n71440 , n71441 , n71442 , n71443 , n71444 , 
 n71445 , n71446 , n71447 , n71448 , n71449 , n71450 , n71451 , n71452 , n71453 , n71454 , 
 n71455 , n71456 , n71457 , n71458 , n71459 , n71460 , n71461 , n71462 , n71463 , n71464 , 
 n71465 , n71466 , n71467 , n71468 , n71469 , n71470 , n71471 , n71472 , n71473 , n71474 , 
 n71475 , n71476 , n71477 , n71478 , n71479 , n71480 , n71481 , n71482 , n71483 , n71484 , 
 n71485 , n71486 , n71487 , n71488 , n71489 , n71490 , n71491 , n71492 , n71493 , n71494 , 
 n71495 , n71496 , n71497 , n71498 , n71499 , n71500 , n71501 , n71502 , n71503 , n71504 , 
 n71505 , n71506 , n71507 , n71508 , n71509 , n71510 , n71511 , n71512 , n71513 , n71514 , 
 n71515 , n71516 , n71517 , n71518 , n71519 , n71520 , n71521 , n71522 , n71523 , n71524 , 
 n71525 , n71526 , n71527 , n71528 , n71529 , n71530 , n71531 , n71532 , n71533 , n71534 , 
 n71535 , n71536 , n71537 , n71538 , n71539 , n71540 , n71541 , n71542 , n71543 , n71544 , 
 n71545 , n71546 , n71547 , n71548 , n71549 , n71550 , n71551 , n71552 , n71553 , n71554 , 
 n71555 , n71556 , n71557 , n71558 , n71559 , n71560 , n71561 , n71562 , n71563 , n71564 , 
 n71565 , n71566 , n71567 , n71568 , n71569 , n71570 , n71571 , n71572 , n71573 , n71574 , 
 n71575 , n71576 , n71577 , n71578 , n71579 , n71580 , n71581 , n71582 , n71583 , n71584 , 
 n71585 , n71586 , n71587 , n71588 , n71589 , n71590 , n71591 , n71592 , n71593 , n71594 , 
 n71595 , n71596 , n71597 , n71598 , n71599 , n71600 , n71601 , n71602 , n71603 , n71604 , 
 n71605 , n71606 , n71607 , n71608 , n71609 , n71610 , n71611 , n71612 , n71613 , n71614 , 
 n71615 , n71616 , n71617 , n71618 , n71619 , n71620 , n71621 , n71622 , n71623 , n71624 , 
 n71625 , n71626 , n71627 , n71628 , n71629 , n71630 , n71631 , n71632 , n71633 , n71634 , 
 n71635 , n71636 , n71637 , n71638 , n71639 , n71640 , n71641 , n71642 , n71643 , n71644 , 
 n71645 , n71646 , n71647 , n71648 , n71649 , n71650 , n71651 , n71652 , n71653 , n71654 , 
 n71655 , n71656 , n71657 , n71658 , n71659 , n71660 , n71661 , n71662 , n71663 , n71664 , 
 n71665 , n71666 , n71667 , n71668 , n71669 , n71670 , n71671 , n71672 , n71673 , n71674 , 
 n71675 , n71676 , n71677 , n71678 , n71679 , n71680 , n71681 , n71682 , n71683 , n71684 , 
 n71685 , n71686 , n71687 , n71688 , n71689 , n71690 , n71691 , n71692 , n71693 , n71694 , 
 n71695 , n71696 , n71697 , n71698 , n71699 , n71700 , n71701 , n71702 , n71703 , n71704 , 
 n71705 , n71706 , n71707 , n71708 , n71709 , n71710 , n71711 , n71712 , n71713 , n71714 , 
 n71715 , n71716 , n71717 , n71718 , n71719 , n71720 , n71721 , n71722 , n71723 , n71724 , 
 n71725 , n71726 , n71727 , n71728 , n71729 , n71730 , n71731 , n71732 , n71733 , n71734 , 
 n71735 , n71736 , n71737 , n71738 , n71739 , n71740 , n71741 , n71742 , n71743 , n71744 , 
 n71745 , n71746 , n71747 , n71748 , n71749 , n71750 , n71751 , n71752 , n71753 , n71754 , 
 n71755 , n71756 , n71757 , n71758 , n71759 , n71760 , n71761 , n71762 , n71763 , n71764 , 
 n71765 , n71766 , n71767 , n71768 , n71769 , n71770 , n71771 , n71772 , n71773 , n71774 , 
 n71775 , n71776 , n71777 , n71778 , n71779 , n71780 , n71781 , n71782 , n71783 , n71784 , 
 n71785 , n71786 , n71787 , n71788 , n71789 , n71790 , n71791 , n71792 , n71793 , n71794 , 
 n71795 , n71796 , n71797 , n71798 , n71799 , n71800 , n71801 , n71802 , n71803 , n71804 , 
 n71805 , n71806 , n71807 , n71808 , n71809 , n71810 , n71811 , n71812 , n71813 , n71814 , 
 n71815 , n71816 , n71817 , n71818 , n71819 , n71820 , n71821 , n71822 , n71823 , n71824 , 
 n71825 , n71826 , n71827 , n71828 , n71829 , n71830 , n71831 , n71832 , n71833 , n71834 , 
 n71835 , n71836 , n71837 , n71838 , n71839 , n71840 , n71841 , n71842 , n71843 , n71844 , 
 n71845 , n71846 , n71847 , n71848 , n71849 , n71850 , n71851 , n71852 , n71853 , n71854 , 
 n71855 , n71856 , n71857 , n71858 , n71859 , n71860 , n71861 , n71862 , n71863 , n71864 , 
 n71865 , n71866 , n71867 , n71868 , n71869 , n71870 , n71871 , n71872 , n71873 , n71874 , 
 n71875 , n71876 , n71877 , n71878 , n71879 , n71880 , n71881 , n71882 , n71883 , n71884 , 
 n71885 , n71886 , n71887 , n71888 , n71889 , n71890 , n71891 , n71892 , n71893 , n71894 , 
 n71895 , n71896 , n71897 , n71898 , n71899 , n71900 , n71901 , n71902 , n71903 , n71904 , 
 n71905 , n71906 , n71907 , n71908 , n71909 , n71910 , n71911 , n71912 , n71913 , n71914 , 
 n71915 , n71916 , n71917 , n71918 , n71919 , n71920 , n71921 , n71922 , n71923 , n71924 , 
 n71925 , n71926 , n71927 , n71928 , n71929 , n71930 , n71931 , n71932 , n71933 , n71934 , 
 n71935 , n71936 , n71937 , n71938 , n71939 , n71940 , n71941 , n71942 , n71943 , n71944 , 
 n71945 , n71946 , n71947 , n71948 , n71949 , n71950 , n71951 , n71952 , n71953 , n71954 , 
 n71955 , n71956 , n71957 , n71958 , n71959 , n71960 , n71961 , n71962 , n71963 , n71964 , 
 n71965 , n71966 , n71967 , n71968 , n71969 , n71970 , n71971 , n71972 , n71973 , n71974 , 
 n71975 , n71976 , n71977 , n71978 , n71979 , n71980 , n71981 , n71982 , n71983 , n71984 , 
 n71985 , n71986 , n71987 , n71988 , n71989 , n71990 , n71991 , n71992 , n71993 , n71994 , 
 n71995 , n71996 , n71997 , n71998 , n71999 , n72000 , n72001 , n72002 , n72003 , n72004 , 
 n72005 , n72006 , n72007 , n72008 , n72009 , n72010 , n72011 , n72012 , n72013 , n72014 , 
 n72015 , n72016 , n72017 , n72018 , n72019 , n72020 , n72021 , n72022 , n72023 , n72024 , 
 n72025 , n72026 , n72027 , n72028 , n72029 , n72030 , n72031 , n72032 , n72033 , n72034 , 
 n72035 , n72036 , n72037 , n72038 , n72039 , n72040 , n72041 , n72042 , n72043 , n72044 , 
 n72045 , n72046 , n72047 , n72048 , n72049 , n72050 , n72051 , n72052 , n72053 , n72054 , 
 n72055 , n72056 , n72057 , n72058 , n72059 , n72060 , n72061 , n72062 , n72063 , n72064 , 
 n72065 , n72066 , n72067 , n72068 , n72069 , n72070 , n72071 , n72072 , n72073 , n72074 , 
 n72075 , n72076 , n72077 , n72078 , n72079 , n72080 , n72081 , n72082 , n72083 , n72084 , 
 n72085 , n72086 , n72087 , n72088 , n72089 , n72090 , n72091 , n72092 , n72093 , n72094 , 
 n72095 , n72096 , n72097 , n72098 , n72099 , n72100 , n72101 , n72102 , n72103 , n72104 , 
 n72105 , n72106 , n72107 , n72108 , n72109 , n72110 , n72111 , n72112 , n72113 , n72114 , 
 n72115 , n72116 , n72117 , n72118 , n72119 , n72120 , n72121 , n72122 , n72123 , n72124 , 
 n72125 , n72126 , n72127 , n72128 , n72129 , n72130 , n72131 , n72132 , n72133 , n72134 , 
 n72135 , n72136 , n72137 , n72138 , n72139 , n72140 , n72141 , n72142 , n72143 , n72144 , 
 n72145 , n72146 , n72147 , n72148 , n72149 , n72150 , n72151 , n72152 , n72153 , n72154 , 
 n72155 , n72156 , n72157 , n72158 , n72159 , n72160 , n72161 , n72162 , n72163 , n72164 , 
 n72165 , n72166 , n72167 , n72168 , n72169 , n72170 , n72171 , n72172 , n72173 , n72174 , 
 n72175 , n72176 , n72177 , n72178 , n72179 , n72180 , n72181 , n72182 , n72183 , n72184 , 
 n72185 , n72186 , n72187 , n72188 , n72189 , n72190 , n72191 , n72192 , n72193 , n72194 , 
 n72195 , n72196 , n72197 , n72198 , n72199 , n72200 , n72201 , n72202 , n72203 , n72204 , 
 n72205 , n72206 , n72207 , n72208 , n72209 , n72210 , n72211 , n72212 , n72213 , n72214 , 
 n72215 , n72216 , n72217 , n72218 , n72219 , n72220 , n72221 , n72222 , n72223 , n72224 , 
 n72225 , n72226 , n72227 , n72228 , n72229 , n72230 , n72231 , n72232 , n72233 , n72234 , 
 n72235 , n72236 , n72237 , n72238 , n72239 , n72240 , n72241 , n72242 , n72243 , n72244 , 
 n72245 , n72246 , n72247 , n72248 , n72249 , n72250 , n72251 , n72252 , n72253 , n72254 , 
 n72255 , n72256 , n72257 , n72258 , n72259 , n72260 , n72261 , n72262 , n72263 , n72264 , 
 n72265 , n72266 , n72267 , n72268 , n72269 , n72270 , n72271 , n72272 , n72273 , n72274 , 
 n72275 , n72276 , n72277 , n72278 , n72279 , n72280 , n72281 , n72282 , n72283 , n72284 , 
 n72285 , n72286 , n72287 , n72288 , n72289 , n72290 , n72291 , n72292 , n72293 , n72294 , 
 n72295 , n72296 , n72297 , n72298 , n72299 , n72300 , n72301 , n72302 , n72303 , n72304 , 
 n72305 , n72306 , n72307 , n72308 , n72309 , n72310 , n72311 , n72312 , n72313 , n72314 , 
 n72315 , n72316 , n72317 , n72318 , n72319 , n72320 , n72321 , n72322 , n72323 , n72324 , 
 n72325 , n72326 , n72327 , n72328 , n72329 , n72330 , n72331 , n72332 , n72333 , n72334 , 
 n72335 , n72336 , n72337 , n72338 , n72339 , n72340 , n72341 , n72342 , n72343 , n72344 , 
 n72345 , n72346 , n72347 , n72348 , n72349 , n72350 , n72351 , n72352 , n72353 , n72354 , 
 n72355 , n72356 , n72357 , n72358 , n72359 , n72360 , n72361 , n72362 , n72363 , n72364 , 
 n72365 , n72366 , n72367 , n72368 , n72369 , n72370 , n72371 , n72372 , n72373 , n72374 , 
 n72375 , n72376 , n72377 , n72378 , n72379 , n72380 , n72381 , n72382 , n72383 , n72384 , 
 n72385 , n72386 , n72387 , n72388 , n72389 , n72390 , n72391 , n72392 , n72393 , n72394 , 
 n72395 , n72396 , n72397 , n72398 , n72399 , n72400 , n72401 , n72402 , n72403 , n72404 , 
 n72405 , n72406 , n72407 , n72408 , n72409 , n72410 , n72411 , n72412 , n72413 , n72414 , 
 n72415 , n72416 , n72417 , n72418 , n72419 , n72420 , n72421 , n72422 , n72423 , n72424 , 
 n72425 , n72426 , n72427 , n72428 , n72429 , n72430 , n72431 , n72432 , n72433 , n72434 , 
 n72435 , n72436 , n72437 , n72438 , n72439 , n72440 , n72441 , n72442 , n72443 , n72444 , 
 n72445 , n72446 , n72447 , n72448 , n72449 , n72450 , n72451 , n72452 , n72453 , n72454 , 
 n72455 , n72456 , n72457 , n72458 , n72459 , n72460 , n72461 , n72462 , n72463 , n72464 , 
 n72465 , n72466 , n72467 , n72468 , n72469 , n72470 , n72471 , n72472 , n72473 , n72474 , 
 n72475 , n72476 , n72477 , n72478 , n72479 , n72480 , n72481 , n72482 , n72483 , n72484 , 
 n72485 , n72486 , n72487 , n72488 , n72489 , n72490 , n72491 , n72492 , n72493 , n72494 , 
 n72495 , n72496 , n72497 , n72498 , n72499 , n72500 , n72501 , n72502 , n72503 , n72504 , 
 n72505 , n72506 , n72507 , n72508 , n72509 , n72510 , n72511 , n72512 , n72513 , n72514 , 
 n72515 , n72516 , n72517 , n72518 , n72519 , n72520 , n72521 , n72522 , n72523 , n72524 , 
 n72525 , n72526 , n72527 , n72528 , n72529 , n72530 , n72531 , n72532 , n72533 , n72534 , 
 n72535 , n72536 , n72537 , n72538 , n72539 , n72540 , n72541 , n72542 , n72543 , n72544 , 
 n72545 , n72546 , n72547 , n72548 , n72549 , n72550 , n72551 , n72552 , n72553 , n72554 , 
 n72555 , n72556 , n72557 , n72558 , n72559 , n72560 , n72561 , n72562 , n72563 , n72564 , 
 n72565 , n72566 , n72567 , n72568 , n72569 , n72570 , n72571 , n72572 , n72573 , n72574 , 
 n72575 , n72576 , n72577 , n72578 , n72579 , n72580 , n72581 , n72582 , n72583 , n72584 , 
 n72585 , n72586 , n72587 , n72588 , n72589 , n72590 , n72591 , n72592 , n72593 , n72594 , 
 n72595 , n72596 , n72597 , n72598 , n72599 , n72600 , n72601 , n72602 , n72603 , n72604 , 
 n72605 , n72606 , n72607 , n72608 , n72609 , n72610 , n72611 , n72612 , n72613 , n72614 , 
 n72615 , n72616 , n72617 , n72618 , n72619 , n72620 , n72621 , n72622 , n72623 , n72624 , 
 n72625 , n72626 , n72627 , n72628 , n72629 , n72630 , n72631 , n72632 , n72633 , n72634 , 
 n72635 , n72636 , n72637 , n72638 , n72639 , n72640 , n72641 , n72642 , n72643 , n72644 , 
 n72645 , n72646 , n72647 , n72648 , n72649 , n72650 , n72651 , n72652 , n72653 , n72654 , 
 n72655 , n72656 , n72657 , n72658 , n72659 , n72660 , n72661 , n72662 , n72663 , n72664 , 
 n72665 , n72666 , n72667 , n72668 , n72669 , n72670 , n72671 , n72672 , n72673 , n72674 , 
 n72675 , n72676 , n72677 , n72678 , n72679 , n72680 , n72681 , n72682 , n72683 , n72684 , 
 n72685 , n72686 , n72687 , n72688 , n72689 , n72690 , n72691 , n72692 , n72693 , n72694 , 
 n72695 , n72696 , n72697 , n72698 , n72699 , n72700 , n72701 , n72702 , n72703 , n72704 , 
 n72705 , n72706 , n72707 , n72708 , n72709 , n72710 , n72711 , n72712 , n72713 , n72714 , 
 n72715 , n72716 , n72717 , n72718 , n72719 , n72720 , n72721 , n72722 , n72723 , n72724 , 
 n72725 , n72726 , n72727 , n72728 , n72729 , n72730 , n72731 , n72732 , n72733 , n72734 , 
 n72735 , n72736 , n72737 , n72738 , n72739 , n72740 , n72741 , n72742 , n72743 , n72744 , 
 n72745 , n72746 , n72747 , n72748 , n72749 , n72750 , n72751 , n72752 , n72753 , n72754 , 
 n72755 , n72756 , n72757 , n72758 , n72759 , n72760 , n72761 , n72762 , n72763 , n72764 , 
 n72765 , n72766 , n72767 , n72768 , n72769 , n72770 , n72771 , n72772 , n72773 , n72774 , 
 n72775 , n72776 , n72777 , n72778 , n72779 , n72780 , n72781 , n72782 , n72783 , n72784 , 
 n72785 , n72786 , n72787 , n72788 , n72789 , n72790 , n72791 , n72792 , n72793 , n72794 , 
 n72795 , n72796 , n72797 , n72798 , n72799 , n72800 , n72801 , n72802 , n72803 , n72804 , 
 n72805 , n72806 , n72807 , n72808 , n72809 , n72810 , n72811 , n72812 , n72813 , n72814 , 
 n72815 , n72816 , n72817 , n72818 , n72819 , n72820 , n72821 , n72822 , n72823 , n72824 , 
 n72825 , n72826 , n72827 , n72828 , n72829 , n72830 , n72831 , n72832 , n72833 , n72834 , 
 n72835 , n72836 , n72837 , n72838 , n72839 , n72840 , n72841 , n72842 , n72843 , n72844 , 
 n72845 , n72846 , n72847 , n72848 , n72849 , n72850 , n72851 , n72852 , n72853 , n72854 , 
 n72855 , n72856 , n72857 , n72858 , n72859 , n72860 , n72861 , n72862 , n72863 , n72864 , 
 n72865 , n72866 , n72867 , n72868 , n72869 , n72870 , n72871 , n72872 , n72873 , n72874 , 
 n72875 , n72876 , n72877 , n72878 , n72879 , n72880 , n72881 , n72882 , n72883 , n72884 , 
 n72885 , n72886 , n72887 , n72888 , n72889 , n72890 , n72891 , n72892 , n72893 , n72894 , 
 n72895 , n72896 , n72897 , n72898 , n72899 , n72900 , n72901 , n72902 , n72903 , n72904 , 
 n72905 , n72906 , n72907 , n72908 , n72909 , n72910 , n72911 , n72912 , n72913 , n72914 , 
 n72915 , n72916 , n72917 , n72918 , n72919 , n72920 , n72921 , n72922 , n72923 , n72924 , 
 n72925 , n72926 , n72927 , n72928 , n72929 , n72930 , n72931 , n72932 , n72933 , n72934 , 
 n72935 , n72936 , n72937 , n72938 , n72939 , n72940 , n72941 , n72942 , n72943 , n72944 , 
 n72945 , n72946 , n72947 , n72948 , n72949 , n72950 , n72951 , n72952 , n72953 , n72954 , 
 n72955 , n72956 , n72957 , n72958 , n72959 , n72960 , n72961 , n72962 , n72963 , n72964 , 
 n72965 , n72966 , n72967 , n72968 , n72969 , n72970 , n72971 , n72972 , n72973 , n72974 , 
 n72975 , n72976 , n72977 , n72978 , n72979 , n72980 , n72981 , n72982 , n72983 , n72984 , 
 n72985 , n72986 , n72987 , n72988 , n72989 , n72990 , n72991 , n72992 , n72993 , n72994 , 
 n72995 , n72996 , n72997 , n72998 , n72999 , n73000 , n73001 , n73002 , n73003 , n73004 , 
 n73005 , n73006 , n73007 , n73008 , n73009 , n73010 , n73011 , n73012 , n73013 , n73014 , 
 n73015 , n73016 , n73017 , n73018 , n73019 , n73020 , n73021 , n73022 , n73023 , n73024 , 
 n73025 , n73026 , n73027 , n73028 , n73029 , n73030 , n73031 , n73032 , n73033 , n73034 , 
 n73035 , n73036 , n73037 , n73038 , n73039 , n73040 , n73041 , n73042 , n73043 , n73044 , 
 n73045 , n73046 , n73047 , n73048 , n73049 , n73050 , n73051 , n73052 , n73053 , n73054 , 
 n73055 , n73056 , n73057 , n73058 , n73059 , n73060 , n73061 , n73062 , n73063 , n73064 , 
 n73065 , n73066 , n73067 , n73068 , n73069 , n73070 , n73071 , n73072 , n73073 , n73074 , 
 n73075 , n73076 , n73077 , n73078 , n73079 , n73080 , n73081 , n73082 , n73083 , n73084 , 
 n73085 , n73086 , n73087 , n73088 , n73089 , n73090 , n73091 , n73092 , n73093 , n73094 , 
 n73095 , n73096 , n73097 , n73098 , n73099 , n73100 , n73101 , n73102 , n73103 , n73104 , 
 n73105 , n73106 , n73107 , n73108 , n73109 , n73110 , n73111 , n73112 , n73113 , n73114 , 
 n73115 , n73116 , n73117 , n73118 , n73119 , n73120 , n73121 , n73122 , n73123 , n73124 , 
 n73125 , n73126 , n73127 , n73128 , n73129 , n73130 , n73131 , n73132 , n73133 , n73134 , 
 n73135 , n73136 , n73137 , n73138 , n73139 , n73140 , n73141 , n73142 , n73143 , n73144 , 
 n73145 , n73146 , n73147 , n73148 , n73149 , n73150 , n73151 , n73152 , n73153 , n73154 , 
 n73155 , n73156 , n73157 , n73158 , n73159 , n73160 , n73161 , n73162 , n73163 , n73164 , 
 n73165 , n73166 , n73167 , n73168 , n73169 , n73170 , n73171 , n73172 , n73173 , n73174 , 
 n73175 , n73176 , n73177 , n73178 , n73179 , n73180 , n73181 , n73182 , n73183 , n73184 , 
 n73185 , n73186 , n73187 , n73188 , n73189 , n73190 , n73191 , n73192 , n73193 , n73194 , 
 n73195 , n73196 , n73197 , n73198 , n73199 , n73200 , n73201 , n73202 , n73203 , n73204 , 
 n73205 , n73206 , n73207 , n73208 , n73209 , n73210 , n73211 , n73212 , n73213 , n73214 , 
 n73215 , n73216 , n73217 , n73218 , n73219 , n73220 , n73221 , n73222 , n73223 , n73224 , 
 n73225 , n73226 , n73227 , n73228 , n73229 , n73230 , n73231 , n73232 , n73233 , n73234 , 
 n73235 , n73236 , n73237 , n73238 , n73239 , n73240 , n73241 , n73242 , n73243 , n73244 , 
 n73245 , n73246 , n73247 , n73248 , n73249 , n73250 , n73251 , n73252 , n73253 , n73254 , 
 n73255 , n73256 , n73257 , n73258 , n73259 , n73260 , n73261 , n73262 , n73263 , n73264 , 
 n73265 , n73266 , n73267 , n73268 , n73269 , n73270 , n73271 , n73272 , n73273 , n73274 , 
 n73275 , n73276 , n73277 , n73278 , n73279 , n73280 , n73281 , n73282 , n73283 , n73284 , 
 n73285 , n73286 , n73287 , n73288 , n73289 , n73290 , n73291 , n73292 , n73293 , n73294 , 
 n73295 , n73296 , n73297 , n73298 , n73299 , n73300 , n73301 , n73302 , n73303 , n73304 , 
 n73305 , n73306 , n73307 , n73308 , n73309 , n73310 , n73311 , n73312 , n73313 , n73314 , 
 n73315 , n73316 , n73317 , n73318 , n73319 , n73320 , n73321 , n73322 , n73323 , n73324 , 
 n73325 , n73326 , n73327 , n73328 , n73329 , n73330 , n73331 , n73332 , n73333 , n73334 , 
 n73335 , n73336 , n73337 , n73338 , n73339 , n73340 , n73341 , n73342 , n73343 , n73344 , 
 n73345 , n73346 , n73347 , n73348 , n73349 , n73350 , n73351 , n73352 , n73353 , n73354 , 
 n73355 , n73356 , n73357 , n73358 , n73359 , n73360 , n73361 , n73362 , n73363 , n73364 , 
 n73365 , n73366 , n73367 , n73368 , n73369 , n73370 , n73371 , n73372 , n73373 , n73374 , 
 n73375 , n73376 , n73377 , n73378 , n73379 , n73380 , n73381 , n73382 , n73383 , n73384 , 
 n73385 , n73386 , n73387 , n73388 , n73389 , n73390 , n73391 , n73392 , n73393 , n73394 , 
 n73395 , n73396 , n73397 , n73398 , n73399 , n73400 , n73401 , n73402 , n73403 , n73404 , 
 n73405 , n73406 , n73407 , n73408 , n73409 , n73410 , n73411 , n73412 , n73413 , n73414 , 
 n73415 , n73416 , n73417 , n73418 , n73419 , n73420 , n73421 , n73422 , n73423 , n73424 , 
 n73425 , n73426 , n73427 , n73428 , n73429 , n73430 , n73431 , n73432 , n73433 , n73434 , 
 n73435 , n73436 , n73437 , n73438 , n73439 , n73440 , n73441 , n73442 , n73443 , n73444 , 
 n73445 , n73446 , n73447 , n73448 , n73449 , n73450 , n73451 , n73452 , n73453 , n73454 , 
 n73455 , n73456 , n73457 , n73458 , n73459 , n73460 , n73461 , n73462 , n73463 , n73464 , 
 n73465 , n73466 , n73467 , n73468 , n73469 , n73470 , n73471 , n73472 , n73473 , n73474 , 
 n73475 , n73476 , n73477 , n73478 , n73479 , n73480 , n73481 , n73482 , n73483 , n73484 , 
 n73485 , n73486 , n73487 , n73488 , n73489 , n73490 , n73491 , n73492 , n73493 , n73494 , 
 n73495 , n73496 , n73497 , n73498 , n73499 , n73500 , n73501 , n73502 , n73503 , n73504 , 
 n73505 , n73506 , n73507 , n73508 , n73509 , n73510 , n73511 , n73512 , n73513 , n73514 , 
 n73515 , n73516 , n73517 , n73518 , n73519 , n73520 , n73521 , n73522 , n73523 , n73524 , 
 n73525 , n73526 , n73527 , n73528 , n73529 , n73530 , n73531 , n73532 , n73533 , n73534 , 
 n73535 , n73536 , n73537 , n73538 , n73539 , n73540 , n73541 , n73542 , n73543 , n73544 , 
 n73545 , n73546 , n73547 , n73548 , n73549 , n73550 , n73551 , n73552 , n73553 , n73554 , 
 n73555 , n73556 , n73557 , n73558 , n73559 , n73560 , n73561 , n73562 , n73563 , n73564 , 
 n73565 , n73566 , n73567 , n73568 , n73569 , n73570 , n73571 , n73572 , n73573 , n73574 , 
 n73575 , n73576 , n73577 , n73578 , n73579 , n73580 , n73581 , n73582 , n73583 , n73584 , 
 n73585 , n73586 , n73587 , n73588 , n73589 , n73590 , n73591 , n73592 , n73593 , n73594 , 
 n73595 , n73596 , n73597 , n73598 , n73599 , n73600 , n73601 , n73602 , n73603 , n73604 , 
 n73605 , n73606 , n73607 , n73608 , n73609 , n73610 , n73611 , n73612 , n73613 , n73614 , 
 n73615 , n73616 , n73617 , n73618 , n73619 , n73620 , n73621 , n73622 , n73623 , n73624 , 
 n73625 , n73626 , n73627 , n73628 , n73629 , n73630 , n73631 , n73632 , n73633 , n73634 , 
 n73635 , n73636 , n73637 , n73638 , n73639 , n73640 , n73641 , n73642 , n73643 , n73644 , 
 n73645 , n73646 , n73647 , n73648 , n73649 , n73650 , n73651 , n73652 , n73653 , n73654 , 
 n73655 , n73656 , n73657 , n73658 , n73659 , n73660 , n73661 , n73662 , n73663 , n73664 , 
 n73665 , n73666 , n73667 , n73668 , n73669 , n73670 , n73671 , n73672 , n73673 , n73674 , 
 n73675 , n73676 , n73677 , n73678 , n73679 , n73680 , n73681 , n73682 , n73683 , n73684 , 
 n73685 , n73686 , n73687 , n73688 , n73689 , n73690 , n73691 , n73692 , n73693 , n73694 , 
 n73695 , n73696 , n73697 , n73698 , n73699 , n73700 , n73701 , n73702 , n73703 , n73704 , 
 n73705 , n73706 , n73707 , n73708 , n73709 , n73710 , n73711 , n73712 , n73713 , n73714 , 
 n73715 , n73716 , n73717 , n73718 , n73719 , n73720 , n73721 , n73722 , n73723 , n73724 , 
 n73725 , n73726 , n73727 , n73728 , n73729 , n73730 , n73731 , n73732 , n73733 , n73734 , 
 n73735 , n73736 , n73737 , n73738 , n73739 , n73740 , n73741 , n73742 , n73743 , n73744 , 
 n73745 , n73746 , n73747 , n73748 , n73749 , n73750 , n73751 , n73752 , n73753 , n73754 , 
 n73755 , n73756 , n73757 , n73758 , n73759 , n73760 , n73761 , n73762 , n73763 , n73764 , 
 n73765 , n73766 , n73767 , n73768 , n73769 , n73770 , n73771 , n73772 , n73773 , n73774 , 
 n73775 , n73776 , n73777 , n73778 , n73779 , n73780 , n73781 , n73782 , n73783 , n73784 , 
 n73785 , n73786 , n73787 , n73788 , n73789 , n73790 , n73791 , n73792 , n73793 , n73794 , 
 n73795 , n73796 , n73797 , n73798 , n73799 , n73800 , n73801 , n73802 , n73803 , n73804 , 
 n73805 , n73806 , n73807 , n73808 , n73809 , n73810 , n73811 , n73812 , n73813 , n73814 , 
 n73815 , n73816 , n73817 , n73818 , n73819 , n73820 , n73821 , n73822 , n73823 , n73824 , 
 n73825 , n73826 , n73827 , n73828 , n73829 , n73830 , n73831 , n73832 , n73833 , n73834 , 
 n73835 , n73836 , n73837 , n73838 , n73839 , n73840 , n73841 , n73842 , n73843 , n73844 , 
 n73845 , n73846 , n73847 , n73848 , n73849 , n73850 , n73851 , n73852 , n73853 , n73854 , 
 n73855 , n73856 , n73857 , n73858 , n73859 , n73860 , n73861 , n73862 , n73863 , n73864 , 
 n73865 , n73866 , n73867 , n73868 , n73869 , n73870 , n73871 , n73872 , n73873 , n73874 , 
 n73875 , n73876 , n73877 , n73878 , n73879 , n73880 , n73881 , n73882 , n73883 , n73884 , 
 n73885 , n73886 , n73887 , n73888 , n73889 , n73890 , n73891 , n73892 , n73893 , n73894 , 
 n73895 , n73896 , n73897 , n73898 , n73899 , n73900 , n73901 , n73902 , n73903 , n73904 , 
 n73905 , n73906 , n73907 , n73908 , n73909 , n73910 , n73911 , n73912 , n73913 , n73914 , 
 n73915 , n73916 , n73917 , n73918 , n73919 , n73920 , n73921 , n73922 , n73923 , n73924 , 
 n73925 , n73926 , n73927 , n73928 , n73929 , n73930 , n73931 , n73932 , n73933 , n73934 , 
 n73935 , n73936 , n73937 , n73938 , n73939 , n73940 , n73941 , n73942 , n73943 , n73944 , 
 n73945 , n73946 , n73947 , n73948 , n73949 , n73950 , n73951 , n73952 , n73953 , n73954 , 
 n73955 , n73956 , n73957 , n73958 , n73959 , n73960 , n73961 , n73962 , n73963 , n73964 , 
 n73965 , n73966 , n73967 , n73968 , n73969 , n73970 , n73971 , n73972 , n73973 , n73974 , 
 n73975 , n73976 , n73977 , n73978 , n73979 , n73980 , n73981 , n73982 , n73983 , n73984 , 
 n73985 , n73986 , n73987 , n73988 , n73989 , n73990 , n73991 , n73992 , n73993 , n73994 , 
 n73995 , n73996 , n73997 , n73998 , n73999 , n74000 , n74001 , n74002 , n74003 , n74004 , 
 n74005 , n74006 , n74007 , n74008 , n74009 , n74010 , n74011 , n74012 , n74013 , n74014 , 
 n74015 , n74016 , n74017 , n74018 , n74019 , n74020 , n74021 , n74022 , n74023 , n74024 , 
 n74025 , n74026 , n74027 , n74028 , n74029 , n74030 , n74031 , n74032 , n74033 , n74034 , 
 n74035 , n74036 , n74037 , n74038 , n74039 , n74040 , n74041 , n74042 , n74043 , n74044 , 
 n74045 , n74046 , n74047 , n74048 , n74049 , n74050 , n74051 , n74052 , n74053 , n74054 , 
 n74055 , n74056 , n74057 , n74058 , n74059 , n74060 , n74061 , n74062 , n74063 , n74064 , 
 n74065 , n74066 , n74067 , n74068 , n74069 , n74070 , n74071 , n74072 , n74073 , n74074 , 
 n74075 , n74076 , n74077 , n74078 , n74079 , n74080 , n74081 , n74082 , n74083 , n74084 , 
 n74085 , n74086 , n74087 , n74088 , n74089 , n74090 , n74091 , n74092 , n74093 , n74094 , 
 n74095 , n74096 , n74097 , n74098 , n74099 , n74100 , n74101 , n74102 , n74103 , n74104 , 
 n74105 , n74106 , n74107 , n74108 , n74109 , n74110 , n74111 , n74112 , n74113 , n74114 , 
 n74115 , n74116 , n74117 , n74118 , n74119 , n74120 , n74121 , n74122 , n74123 , n74124 , 
 n74125 , n74126 , n74127 , n74128 , n74129 , n74130 , n74131 , n74132 , n74133 , n74134 , 
 n74135 , n74136 , n74137 , n74138 , n74139 , n74140 , n74141 , n74142 , n74143 , n74144 , 
 n74145 , n74146 , n74147 , n74148 , n74149 , n74150 , n74151 , n74152 , n74153 , n74154 , 
 n74155 , n74156 , n74157 , n74158 , n74159 , n74160 , n74161 , n74162 , n74163 , n74164 , 
 n74165 , n74166 , n74167 , n74168 , n74169 , n74170 , n74171 , n74172 , n74173 , n74174 , 
 n74175 , n74176 , n74177 , n74178 , n74179 , n74180 , n74181 , n74182 , n74183 , n74184 , 
 n74185 , n74186 , n74187 , n74188 , n74189 , n74190 , n74191 , n74192 , n74193 , n74194 , 
 n74195 , n74196 , n74197 , n74198 , n74199 , n74200 , n74201 , n74202 , n74203 , n74204 , 
 n74205 , n74206 , n74207 , n74208 , n74209 , n74210 , n74211 , n74212 , n74213 , n74214 , 
 n74215 , n74216 , n74217 , n74218 , n74219 , n74220 , n74221 , n74222 , n74223 , n74224 , 
 n74225 , n74226 , n74227 , n74228 , n74229 , n74230 , n74231 , n74232 , n74233 , n74234 , 
 n74235 , n74236 , n74237 , n74238 , n74239 , n74240 , n74241 , n74242 , n74243 , n74244 , 
 n74245 , n74246 , n74247 , n74248 , n74249 , n74250 , n74251 , n74252 , n74253 , n74254 , 
 n74255 , n74256 , n74257 , n74258 , n74259 , n74260 , n74261 , n74262 , n74263 , n74264 , 
 n74265 , n74266 , n74267 , n74268 , n74269 , n74270 , n74271 , n74272 , n74273 , n74274 , 
 n74275 , n74276 , n74277 , n74278 , n74279 , n74280 , n74281 , n74282 , n74283 , n74284 , 
 n74285 , n74286 , n74287 , n74288 , n74289 , n74290 , n74291 , n74292 , n74293 , n74294 , 
 n74295 , n74296 , n74297 , n74298 , n74299 , n74300 , n74301 , n74302 , n74303 , n74304 , 
 n74305 , n74306 , n74307 , n74308 , n74309 , n74310 , n74311 , n74312 , n74313 , n74314 , 
 n74315 , n74316 , n74317 , n74318 , n74319 , n74320 , n74321 , n74322 , n74323 , n74324 , 
 n74325 , n74326 , n74327 , n74328 , n74329 , n74330 , n74331 , n74332 , n74333 , n74334 , 
 n74335 , n74336 , n74337 , n74338 , n74339 , n74340 , n74341 , n74342 , n74343 , n74344 , 
 n74345 , n74346 , n74347 , n74348 , n74349 , n74350 , n74351 , n74352 , n74353 , n74354 , 
 n74355 , n74356 , n74357 , n74358 , n74359 , n74360 , n74361 , n74362 , n74363 , n74364 , 
 n74365 , n74366 , n74367 , n74368 , n74369 , n74370 , n74371 , n74372 , n74373 , n74374 , 
 n74375 , n74376 , n74377 , n74378 , n74379 , n74380 , n74381 , n74382 , n74383 , n74384 , 
 n74385 , n74386 , n74387 , n74388 , n74389 , n74390 , n74391 , n74392 , n74393 , n74394 , 
 n74395 , n74396 , n74397 , n74398 , n74399 , n74400 , n74401 , n74402 , n74403 , n74404 , 
 n74405 , n74406 , n74407 , n74408 , n74409 , n74410 , n74411 , n74412 , n74413 , n74414 , 
 n74415 , n74416 , n74417 , n74418 , n74419 , n74420 , n74421 , n74422 , n74423 , n74424 , 
 n74425 , n74426 , n74427 , n74428 , n74429 , n74430 , n74431 , n74432 , n74433 , n74434 , 
 n74435 , n74436 , n74437 , n74438 , n74439 , n74440 , n74441 , n74442 , n74443 , n74444 , 
 n74445 , n74446 , n74447 , n74448 , n74449 , n74450 , n74451 , n74452 , n74453 , n74454 , 
 n74455 , n74456 , n74457 , n74458 , n74459 , n74460 , n74461 , n74462 , n74463 , n74464 , 
 n74465 , n74466 , n74467 , n74468 , n74469 , n74470 , n74471 , n74472 , n74473 , n74474 , 
 n74475 , n74476 , n74477 , n74478 , n74479 , n74480 , n74481 , n74482 , n74483 , n74484 , 
 n74485 , n74486 , n74487 , n74488 , n74489 , n74490 , n74491 , n74492 , n74493 , n74494 , 
 n74495 , n74496 , n74497 , n74498 , n74499 , n74500 , n74501 , n74502 , n74503 , n74504 , 
 n74505 , n74506 , n74507 , n74508 , n74509 , n74510 , n74511 , n74512 , n74513 , n74514 , 
 n74515 , n74516 , n74517 , n74518 , n74519 , n74520 , n74521 , n74522 , n74523 , n74524 , 
 n74525 , n74526 , n74527 , n74528 , n74529 , n74530 , n74531 , n74532 , n74533 , n74534 , 
 n74535 , n74536 , n74537 , n74538 , n74539 , n74540 , n74541 , n74542 , n74543 , n74544 , 
 n74545 , n74546 , n74547 , n74548 , n74549 , n74550 , n74551 , n74552 , n74553 , n74554 , 
 n74555 , n74556 , n74557 , n74558 , n74559 , n74560 , n74561 , n74562 , n74563 , n74564 , 
 n74565 , n74566 , n74567 , n74568 , n74569 , n74570 , n74571 , n74572 , n74573 , n74574 , 
 n74575 , n74576 , n74577 , n74578 , n74579 , n74580 , n74581 , n74582 , n74583 , n74584 , 
 n74585 , n74586 , n74587 , n74588 , n74589 , n74590 , n74591 , n74592 , n74593 , n74594 , 
 n74595 , n74596 , n74597 , n74598 , n74599 , n74600 , n74601 , n74602 , n74603 , n74604 , 
 n74605 , n74606 , n74607 , n74608 , n74609 , n74610 , n74611 , n74612 , n74613 , n74614 , 
 n74615 , n74616 , n74617 , n74618 , n74619 , n74620 , n74621 , n74622 , n74623 , n74624 , 
 n74625 , n74626 , n74627 , n74628 , n74629 , n74630 , n74631 , n74632 , n74633 , n74634 , 
 n74635 , n74636 , n74637 , n74638 , n74639 , n74640 , n74641 , n74642 , n74643 , n74644 , 
 n74645 , n74646 , n74647 , n74648 , n74649 , n74650 , n74651 , n74652 , n74653 , n74654 , 
 n74655 , n74656 , n74657 , n74658 , n74659 , n74660 , n74661 , n74662 , n74663 , n74664 , 
 n74665 , n74666 , n74667 , n74668 , n74669 , n74670 , n74671 , n74672 , n74673 , n74674 , 
 n74675 , n74676 , n74677 , n74678 , n74679 , n74680 , n74681 , n74682 , n74683 , n74684 , 
 n74685 , n74686 , n74687 , n74688 , n74689 , n74690 , n74691 , n74692 , n74693 , n74694 , 
 n74695 , n74696 , n74697 , n74698 , n74699 , n74700 , n74701 , n74702 , n74703 , n74704 , 
 n74705 , n74706 , n74707 , n74708 , n74709 , n74710 , n74711 , n74712 , n74713 , n74714 , 
 n74715 , n74716 , n74717 , n74718 , n74719 , n74720 , n74721 , n74722 , n74723 , n74724 , 
 n74725 , n74726 , n74727 , n74728 , n74729 , n74730 , n74731 , n74732 , n74733 , n74734 , 
 n74735 , n74736 , n74737 , n74738 , n74739 , n74740 , n74741 , n74742 , n74743 , n74744 , 
 n74745 , n74746 , n74747 , n74748 , n74749 , n74750 , n74751 , n74752 , n74753 , n74754 , 
 n74755 , n74756 , n74757 , n74758 , n74759 , n74760 , n74761 , n74762 , n74763 , n74764 , 
 n74765 , n74766 , n74767 , n74768 , n74769 , n74770 , n74771 , n74772 , n74773 , n74774 , 
 n74775 , n74776 , n74777 , n74778 , n74779 , n74780 , n74781 , n74782 , n74783 , n74784 , 
 n74785 , n74786 , n74787 , n74788 , n74789 , n74790 , n74791 , n74792 , n74793 , n74794 , 
 n74795 , n74796 , n74797 , n74798 , n74799 , n74800 , n74801 , n74802 , n74803 , n74804 , 
 n74805 , n74806 , n74807 , n74808 , n74809 , n74810 , n74811 , n74812 , n74813 , n74814 , 
 n74815 , n74816 , n74817 , n74818 , n74819 , n74820 , n74821 , n74822 , n74823 , n74824 , 
 n74825 , n74826 , n74827 , n74828 , n74829 , n74830 , n74831 , n74832 , n74833 , n74834 , 
 n74835 , n74836 , n74837 , n74838 , n74839 , n74840 , n74841 , n74842 , n74843 , n74844 , 
 n74845 , n74846 , n74847 , n74848 , n74849 , n74850 , n74851 , n74852 , n74853 , n74854 , 
 n74855 , n74856 , n74857 , n74858 , n74859 , n74860 , n74861 , n74862 , n74863 , n74864 , 
 n74865 , n74866 , n74867 , n74868 , n74869 , n74870 , n74871 , n74872 , n74873 , n74874 , 
 n74875 , n74876 , n74877 , n74878 , n74879 , n74880 , n74881 , n74882 , n74883 , n74884 , 
 n74885 , n74886 , n74887 , n74888 , n74889 , n74890 , n74891 , n74892 , n74893 , n74894 , 
 n74895 , n74896 , n74897 , n74898 , n74899 , n74900 , n74901 , n74902 , n74903 , n74904 , 
 n74905 , n74906 , n74907 , n74908 , n74909 , n74910 , n74911 , n74912 , n74913 , n74914 , 
 n74915 , n74916 , n74917 , n74918 , n74919 , n74920 , n74921 , n74922 , n74923 , n74924 , 
 n74925 , n74926 , n74927 , n74928 , n74929 , n74930 , n74931 , n74932 , n74933 , n74934 , 
 n74935 , n74936 , n74937 , n74938 , n74939 , n74940 , n74941 , n74942 , n74943 , n74944 , 
 n74945 , n74946 , n74947 , n74948 , n74949 , n74950 , n74951 , n74952 , n74953 , n74954 , 
 n74955 , n74956 , n74957 , n74958 , n74959 , n74960 , n74961 , n74962 , n74963 , n74964 , 
 n74965 , n74966 , n74967 , n74968 , n74969 , n74970 , n74971 , n74972 , n74973 , n74974 , 
 n74975 , n74976 , n74977 , n74978 , n74979 , n74980 , n74981 , n74982 , n74983 , n74984 , 
 n74985 , n74986 , n74987 , n74988 , n74989 , n74990 , n74991 , n74992 , n74993 , n74994 , 
 n74995 , n74996 , n74997 , n74998 , n74999 , n75000 , n75001 , n75002 , n75003 , n75004 , 
 n75005 , n75006 , n75007 , n75008 , n75009 , n75010 , n75011 , n75012 , n75013 , n75014 , 
 n75015 , n75016 , n75017 , n75018 , n75019 , n75020 , n75021 , n75022 , n75023 , n75024 , 
 n75025 , n75026 , n75027 , n75028 , n75029 , n75030 , n75031 , n75032 , n75033 , n75034 , 
 n75035 , n75036 , n75037 , n75038 , n75039 , n75040 , n75041 , n75042 , n75043 , n75044 , 
 n75045 , n75046 , n75047 , n75048 , n75049 , n75050 , n75051 , n75052 , n75053 , n75054 , 
 n75055 , n75056 , n75057 , n75058 , n75059 , n75060 , n75061 , n75062 , n75063 , n75064 , 
 n75065 , n75066 , n75067 , n75068 , n75069 , n75070 , n75071 , n75072 , n75073 , n75074 , 
 n75075 , n75076 , n75077 , n75078 , n75079 , n75080 , n75081 , n75082 , n75083 , n75084 , 
 n75085 , n75086 , n75087 , n75088 , n75089 , n75090 , n75091 , n75092 , n75093 , n75094 , 
 n75095 , n75096 , n75097 , n75098 , n75099 , n75100 , n75101 , n75102 , n75103 , n75104 , 
 n75105 , n75106 , n75107 , n75108 , n75109 , n75110 , n75111 , n75112 , n75113 , n75114 , 
 n75115 , n75116 , n75117 , n75118 , n75119 , n75120 , n75121 , n75122 , n75123 , n75124 , 
 n75125 , n75126 , n75127 , n75128 , n75129 , n75130 , n75131 , n75132 , n75133 , n75134 , 
 n75135 , n75136 , n75137 , n75138 , n75139 , n75140 , n75141 , n75142 , n75143 , n75144 , 
 n75145 , n75146 , n75147 , n75148 , n75149 , n75150 , n75151 , n75152 , n75153 , n75154 , 
 n75155 , n75156 , n75157 , n75158 , n75159 , n75160 , n75161 , n75162 , n75163 , n75164 , 
 n75165 , n75166 , n75167 , n75168 , n75169 , n75170 , n75171 , n75172 , n75173 , n75174 , 
 n75175 , n75176 , n75177 , n75178 , n75179 , n75180 , n75181 , n75182 , n75183 , n75184 , 
 n75185 , n75186 , n75187 , n75188 , n75189 , n75190 , n75191 , n75192 , n75193 , n75194 , 
 n75195 , n75196 , n75197 , n75198 , n75199 , n75200 , n75201 , n75202 , n75203 , n75204 , 
 n75205 , n75206 , n75207 , n75208 , n75209 , n75210 , n75211 , n75212 , n75213 , n75214 , 
 n75215 , n75216 , n75217 , n75218 , n75219 , n75220 , n75221 , n75222 , n75223 , n75224 , 
 n75225 , n75226 , n75227 , n75228 , n75229 , n75230 , n75231 , n75232 , n75233 , n75234 , 
 n75235 , n75236 , n75237 , n75238 , n75239 , n75240 , n75241 , n75242 , n75243 , n75244 , 
 n75245 , n75246 , n75247 , n75248 , n75249 , n75250 , n75251 , n75252 , n75253 , n75254 , 
 n75255 , n75256 , n75257 , n75258 , n75259 , n75260 , n75261 , n75262 , n75263 , n75264 , 
 n75265 , n75266 , n75267 , n75268 , n75269 , n75270 , n75271 , n75272 , n75273 , n75274 , 
 n75275 , n75276 , n75277 , n75278 , n75279 , n75280 , n75281 , n75282 , n75283 , n75284 , 
 n75285 , n75286 , n75287 , n75288 , n75289 , n75290 , n75291 , n75292 , n75293 , n75294 , 
 n75295 , n75296 , n75297 , n75298 , n75299 , n75300 , n75301 , n75302 , n75303 , n75304 , 
 n75305 , n75306 , n75307 , n75308 , n75309 , n75310 , n75311 , n75312 , n75313 , n75314 , 
 n75315 , n75316 , n75317 , n75318 , n75319 , n75320 , n75321 , n75322 , n75323 , n75324 , 
 n75325 , n75326 , n75327 , n75328 , n75329 , n75330 , n75331 , n75332 , n75333 , n75334 , 
 n75335 , n75336 , n75337 , n75338 , n75339 , n75340 , n75341 , n75342 , n75343 , n75344 , 
 n75345 , n75346 , n75347 , n75348 , n75349 , n75350 , n75351 , n75352 , n75353 , n75354 , 
 n75355 , n75356 , n75357 , n75358 , n75359 , n75360 , n75361 , n75362 , n75363 , n75364 , 
 n75365 , n75366 , n75367 , n75368 , n75369 , n75370 , n75371 , n75372 , n75373 , n75374 , 
 n75375 , n75376 , n75377 , n75378 , n75379 , n75380 , n75381 , n75382 , n75383 , n75384 , 
 n75385 , n75386 , n75387 , n75388 , n75389 , n75390 , n75391 , n75392 , n75393 , n75394 , 
 n75395 , n75396 , n75397 , n75398 , n75399 , n75400 , n75401 , n75402 , n75403 , n75404 , 
 n75405 , n75406 , n75407 , n75408 , n75409 , n75410 , n75411 , n75412 , n75413 , n75414 , 
 n75415 , n75416 , n75417 , n75418 , n75419 , n75420 , n75421 , n75422 , n75423 , n75424 , 
 n75425 , n75426 , n75427 , n75428 , n75429 , n75430 , n75431 , n75432 , n75433 , n75434 , 
 n75435 , n75436 , n75437 , n75438 , n75439 , n75440 , n75441 , n75442 , n75443 , n75444 , 
 n75445 , n75446 , n75447 , n75448 , n75449 , n75450 , n75451 , n75452 , n75453 , n75454 , 
 n75455 , n75456 , n75457 , n75458 , n75459 , n75460 , n75461 , n75462 , n75463 , n75464 , 
 n75465 , n75466 , n75467 , n75468 , n75469 , n75470 , n75471 , n75472 , n75473 , n75474 , 
 n75475 , n75476 , n75477 , n75478 , n75479 , n75480 , n75481 , n75482 , n75483 , n75484 , 
 n75485 , n75486 , n75487 , n75488 , n75489 , n75490 , n75491 , n75492 , n75493 , n75494 , 
 n75495 , n75496 , n75497 , n75498 , n75499 , n75500 , n75501 , n75502 , n75503 , n75504 , 
 n75505 , n75506 , n75507 , n75508 , n75509 , n75510 , n75511 , n75512 , n75513 , n75514 , 
 n75515 , n75516 , n75517 , n75518 , n75519 , n75520 , n75521 , n75522 , n75523 , n75524 , 
 n75525 , n75526 , n75527 , n75528 , n75529 , n75530 , n75531 , n75532 , n75533 , n75534 , 
 n75535 , n75536 , n75537 , n75538 , n75539 , n75540 , n75541 , n75542 , n75543 , n75544 , 
 n75545 , n75546 , n75547 , n75548 , n75549 , n75550 , n75551 , n75552 , n75553 , n75554 , 
 n75555 , n75556 , n75557 , n75558 , n75559 , n75560 , n75561 , n75562 , n75563 , n75564 , 
 n75565 , n75566 , n75567 , n75568 , n75569 , n75570 , n75571 , n75572 , n75573 , n75574 , 
 n75575 , n75576 , n75577 , n75578 , n75579 , n75580 , n75581 , n75582 , n75583 , n75584 , 
 n75585 , n75586 , n75587 , n75588 , n75589 , n75590 , n75591 , n75592 , n75593 , n75594 , 
 n75595 , n75596 , n75597 , n75598 , n75599 , n75600 , n75601 , n75602 , n75603 , n75604 , 
 n75605 , n75606 , n75607 , n75608 , n75609 , n75610 , n75611 , n75612 , n75613 , n75614 , 
 n75615 , n75616 , n75617 , n75618 , n75619 , n75620 , n75621 , n75622 , n75623 , n75624 , 
 n75625 , n75626 , n75627 , n75628 , n75629 , n75630 , n75631 , n75632 , n75633 , n75634 , 
 n75635 , n75636 , n75637 , n75638 , n75639 , n75640 , n75641 , n75642 , n75643 , n75644 , 
 n75645 , n75646 , n75647 , n75648 , n75649 , n75650 , n75651 , n75652 , n75653 , n75654 , 
 n75655 , n75656 , n75657 , n75658 , n75659 , n75660 , n75661 , n75662 , n75663 , n75664 , 
 n75665 , n75666 , n75667 , n75668 , n75669 , n75670 , n75671 , n75672 , n75673 , n75674 , 
 n75675 , n75676 , n75677 , n75678 , n75679 , n75680 , n75681 , n75682 , n75683 , n75684 , 
 n75685 , n75686 , n75687 , n75688 , n75689 , n75690 , n75691 , n75692 , n75693 , n75694 , 
 n75695 , n75696 , n75697 , n75698 , n75699 , n75700 , n75701 , n75702 , n75703 , n75704 , 
 n75705 , n75706 , n75707 , n75708 , n75709 , n75710 , n75711 , n75712 , n75713 , n75714 , 
 n75715 , n75716 , n75717 , n75718 , n75719 , n75720 , n75721 , n75722 , n75723 , n75724 , 
 n75725 , n75726 , n75727 , n75728 , n75729 , n75730 , n75731 , n75732 , n75733 , n75734 , 
 n75735 , n75736 , n75737 , n75738 , n75739 , n75740 , n75741 , n75742 , n75743 , n75744 , 
 n75745 , n75746 , n75747 , n75748 , n75749 , n75750 , n75751 , n75752 , n75753 , n75754 , 
 n75755 , n75756 , n75757 , n75758 , n75759 , n75760 , n75761 , n75762 , n75763 , n75764 , 
 n75765 , n75766 , n75767 , n75768 , n75769 , n75770 , n75771 , n75772 , n75773 , n75774 , 
 n75775 , n75776 , n75777 , n75778 , n75779 , n75780 , n75781 , n75782 , n75783 , n75784 , 
 n75785 , n75786 , n75787 , n75788 , n75789 , n75790 , n75791 , n75792 , n75793 , n75794 , 
 n75795 , n75796 , n75797 , n75798 , n75799 , n75800 , n75801 , n75802 , n75803 , n75804 , 
 n75805 , n75806 , n75807 , n75808 , n75809 , n75810 , n75811 , n75812 , n75813 , n75814 , 
 n75815 , n75816 , n75817 , n75818 , n75819 , n75820 , n75821 , n75822 , n75823 , n75824 , 
 n75825 , n75826 , n75827 , n75828 , n75829 , n75830 , n75831 , n75832 , n75833 , n75834 , 
 n75835 , n75836 , n75837 , n75838 , n75839 , n75840 , n75841 , n75842 , n75843 , n75844 , 
 n75845 , n75846 , n75847 , n75848 , n75849 , n75850 , n75851 , n75852 , n75853 , n75854 , 
 n75855 , n75856 , n75857 , n75858 , n75859 , n75860 , n75861 , n75862 , n75863 , n75864 , 
 n75865 , n75866 , n75867 , n75868 , n75869 , n75870 , n75871 , n75872 , n75873 , n75874 , 
 n75875 , n75876 , n75877 , n75878 , n75879 , n75880 , n75881 , n75882 , n75883 , n75884 , 
 n75885 , n75886 , n75887 , n75888 , n75889 , n75890 , n75891 , n75892 , n75893 , n75894 , 
 n75895 , n75896 , n75897 , n75898 , n75899 , n75900 , n75901 , n75902 , n75903 , n75904 , 
 n75905 , n75906 , n75907 , n75908 , n75909 , n75910 , n75911 , n75912 , n75913 , n75914 , 
 n75915 , n75916 , n75917 , n75918 , n75919 , n75920 , n75921 , n75922 , n75923 , n75924 , 
 n75925 , n75926 , n75927 , n75928 , n75929 , n75930 , n75931 , n75932 , n75933 , n75934 , 
 n75935 , n75936 , n75937 , n75938 , n75939 , n75940 , n75941 , n75942 , n75943 , n75944 , 
 n75945 , n75946 , n75947 , n75948 , n75949 , n75950 , n75951 , n75952 , n75953 , n75954 , 
 n75955 , n75956 , n75957 , n75958 , n75959 , n75960 , n75961 , n75962 , n75963 , n75964 , 
 n75965 , n75966 , n75967 , n75968 , n75969 , n75970 , n75971 , n75972 , n75973 , n75974 , 
 n75975 , n75976 , n75977 , n75978 , n75979 , n75980 , n75981 , n75982 , n75983 , n75984 , 
 n75985 , n75986 , n75987 , n75988 , n75989 , n75990 , n75991 , n75992 , n75993 , n75994 , 
 n75995 , n75996 , n75997 , n75998 , n75999 , n76000 , n76001 , n76002 , n76003 , n76004 , 
 n76005 , n76006 , n76007 , n76008 , n76009 , n76010 , n76011 , n76012 , n76013 , n76014 , 
 n76015 , n76016 , n76017 , n76018 , n76019 , n76020 , n76021 , n76022 , n76023 , n76024 , 
 n76025 , n76026 , n76027 , n76028 , n76029 , n76030 , n76031 , n76032 , n76033 , n76034 , 
 n76035 , n76036 , n76037 , n76038 , n76039 , n76040 , n76041 , n76042 , n76043 , n76044 , 
 n76045 , n76046 , n76047 , n76048 , n76049 , n76050 , n76051 , n76052 , n76053 , n76054 , 
 n76055 , n76056 , n76057 , n76058 , n76059 , n76060 , n76061 , n76062 , n76063 , n76064 , 
 n76065 , n76066 , n76067 , n76068 , n76069 , n76070 , n76071 , n76072 , n76073 , n76074 , 
 n76075 , n76076 , n76077 , n76078 , n76079 , n76080 , n76081 , n76082 , n76083 , n76084 , 
 n76085 , n76086 , n76087 , n76088 , n76089 , n76090 , n76091 , n76092 , n76093 , n76094 , 
 n76095 , n76096 , n76097 , n76098 , n76099 , n76100 , n76101 , n76102 , n76103 , n76104 , 
 n76105 , n76106 , n76107 , n76108 , n76109 , n76110 , n76111 , n76112 , n76113 , n76114 , 
 n76115 , n76116 , n76117 , n76118 , n76119 , n76120 , n76121 , n76122 , n76123 , n76124 , 
 n76125 , n76126 , n76127 , n76128 , n76129 , n76130 , n76131 , n76132 , n76133 , n76134 , 
 n76135 , n76136 , n76137 , n76138 , n76139 , n76140 , n76141 , n76142 , n76143 , n76144 , 
 n76145 , n76146 , n76147 , n76148 , n76149 , n76150 , n76151 , n76152 , n76153 , n76154 , 
 n76155 , n76156 , n76157 , n76158 , n76159 , n76160 , n76161 , n76162 , n76163 , n76164 , 
 n76165 , n76166 , n76167 , n76168 , n76169 , n76170 , n76171 , n76172 , n76173 , n76174 , 
 n76175 , n76176 , n76177 , n76178 , n76179 , n76180 , n76181 , n76182 , n76183 , n76184 , 
 n76185 , n76186 , n76187 , n76188 , n76189 , n76190 , n76191 , n76192 , n76193 , n76194 , 
 n76195 , n76196 , n76197 , n76198 , n76199 , n76200 , n76201 , n76202 , n76203 , n76204 , 
 n76205 , n76206 , n76207 , n76208 , n76209 , n76210 , n76211 , n76212 , n76213 , n76214 , 
 n76215 , n76216 , n76217 , n76218 , n76219 , n76220 , n76221 , n76222 , n76223 , n76224 , 
 n76225 , n76226 , n76227 , n76228 , n76229 , n76230 , n76231 , n76232 , n76233 , n76234 , 
 n76235 , n76236 , n76237 , n76238 , n76239 , n76240 , n76241 , n76242 , n76243 , n76244 , 
 n76245 , n76246 , n76247 , n76248 , n76249 , n76250 , n76251 , n76252 , n76253 , n76254 , 
 n76255 , n76256 , n76257 , n76258 , n76259 , n76260 , n76261 , n76262 , n76263 , n76264 , 
 n76265 , n76266 , n76267 , n76268 , n76269 , n76270 , n76271 , n76272 , n76273 , n76274 , 
 n76275 , n76276 , n76277 , n76278 , n76279 , n76280 , n76281 , n76282 , n76283 , n76284 , 
 n76285 , n76286 , n76287 , n76288 , n76289 , n76290 , n76291 , n76292 , n76293 , n76294 , 
 n76295 , n76296 , n76297 , n76298 , n76299 , n76300 , n76301 , n76302 , n76303 , n76304 , 
 n76305 , n76306 , n76307 , n76308 , n76309 , n76310 , n76311 , n76312 , n76313 , n76314 , 
 n76315 , n76316 , n76317 , n76318 , n76319 , n76320 , n76321 , n76322 , n76323 , n76324 , 
 n76325 , n76326 , n76327 , n76328 , n76329 , n76330 , n76331 , n76332 , n76333 , n76334 , 
 n76335 , n76336 , n76337 , n76338 , n76339 , n76340 , n76341 , n76342 , n76343 , n76344 , 
 n76345 , n76346 , n76347 , n76348 , n76349 , n76350 , n76351 , n76352 , n76353 , n76354 , 
 n76355 , n76356 , n76357 , n76358 , n76359 , n76360 , n76361 , n76362 , n76363 , n76364 , 
 n76365 , n76366 , n76367 , n76368 , n76369 , n76370 , n76371 , n76372 , n76373 , n76374 , 
 n76375 , n76376 , n76377 , n76378 , n76379 , n76380 , n76381 , n76382 , n76383 , n76384 , 
 n76385 , n76386 , n76387 , n76388 , n76389 , n76390 , n76391 , n76392 , n76393 , n76394 , 
 n76395 , n76396 , n76397 , n76398 , n76399 , n76400 , n76401 , n76402 , n76403 , n76404 , 
 n76405 , n76406 , n76407 , n76408 , n76409 , n76410 , n76411 , n76412 , n76413 , n76414 , 
 n76415 , n76416 , n76417 , n76418 , n76419 , n76420 , n76421 , n76422 , n76423 , n76424 , 
 n76425 , n76426 , n76427 , n76428 , n76429 , n76430 , n76431 , n76432 , n76433 , n76434 , 
 n76435 , n76436 , n76437 , n76438 , n76439 , n76440 , n76441 , n76442 , n76443 , n76444 , 
 n76445 , n76446 , n76447 , n76448 , n76449 , n76450 , n76451 , n76452 , n76453 , n76454 , 
 n76455 , n76456 , n76457 , n76458 , n76459 , n76460 , n76461 , n76462 , n76463 , n76464 , 
 n76465 , n76466 , n76467 , n76468 , n76469 , n76470 , n76471 , n76472 , n76473 , n76474 , 
 n76475 , n76476 , n76477 , n76478 , n76479 , n76480 , n76481 , n76482 , n76483 , n76484 , 
 n76485 , n76486 , n76487 , n76488 , n76489 , n76490 , n76491 , n76492 , n76493 , n76494 , 
 n76495 , n76496 , n76497 , n76498 , n76499 , n76500 , n76501 , n76502 , n76503 , n76504 , 
 n76505 , n76506 , n76507 , n76508 , n76509 , n76510 , n76511 , n76512 , n76513 , n76514 , 
 n76515 , n76516 , n76517 , n76518 , n76519 , n76520 , n76521 , n76522 , n76523 , n76524 , 
 n76525 , n76526 , n76527 , n76528 , n76529 , n76530 , n76531 , n76532 , n76533 , n76534 , 
 n76535 , n76536 , n76537 , n76538 , n76539 , n76540 , n76541 , n76542 , n76543 , n76544 , 
 n76545 , n76546 , n76547 , n76548 , n76549 , n76550 , n76551 , n76552 , n76553 , n76554 , 
 n76555 , n76556 , n76557 , n76558 , n76559 , n76560 , n76561 , n76562 , n76563 , n76564 , 
 n76565 , n76566 , n76567 , n76568 , n76569 , n76570 , n76571 , n76572 , n76573 , n76574 , 
 n76575 , n76576 , n76577 , n76578 , n76579 , n76580 , n76581 , n76582 , n76583 , n76584 , 
 n76585 , n76586 , n76587 , n76588 , n76589 , n76590 , n76591 , n76592 , n76593 , n76594 , 
 n76595 , n76596 , n76597 , n76598 , n76599 , n76600 , n76601 , n76602 , n76603 , n76604 , 
 n76605 , n76606 , n76607 , n76608 , n76609 , n76610 , n76611 , n76612 , n76613 , n76614 , 
 n76615 , n76616 , n76617 , n76618 , n76619 , n76620 , n76621 , n76622 , n76623 , n76624 , 
 n76625 , n76626 , n76627 , n76628 , n76629 , n76630 , n76631 , n76632 , n76633 , n76634 , 
 n76635 , n76636 , n76637 , n76638 , n76639 , n76640 , n76641 , n76642 , n76643 , n76644 , 
 n76645 , n76646 , n76647 , n76648 , n76649 , n76650 , n76651 , n76652 , n76653 , n76654 , 
 n76655 , n76656 , n76657 , n76658 , n76659 , n76660 , n76661 , n76662 , n76663 , n76664 , 
 n76665 , n76666 , n76667 , n76668 , n76669 , n76670 , n76671 , n76672 , n76673 , n76674 , 
 n76675 , n76676 , n76677 , n76678 , n76679 , n76680 , n76681 , n76682 , n76683 , n76684 , 
 n76685 , n76686 , n76687 , n76688 , n76689 , n76690 , n76691 , n76692 , n76693 , n76694 , 
 n76695 , n76696 , n76697 , n76698 , n76699 , n76700 , n76701 , n76702 , n76703 , n76704 , 
 n76705 , n76706 , n76707 , n76708 , n76709 , n76710 , n76711 , n76712 , n76713 , n76714 , 
 n76715 , n76716 , n76717 , n76718 , n76719 , n76720 , n76721 , n76722 , n76723 , n76724 , 
 n76725 , n76726 , n76727 , n76728 , n76729 , n76730 , n76731 , n76732 , n76733 , n76734 , 
 n76735 , n76736 , n76737 , n76738 , n76739 , n76740 , n76741 , n76742 , n76743 , n76744 , 
 n76745 , n76746 , n76747 , n76748 , n76749 , n76750 , n76751 , n76752 , n76753 , n76754 , 
 n76755 , n76756 , n76757 , n76758 , n76759 , n76760 , n76761 , n76762 , n76763 , n76764 , 
 n76765 , n76766 , n76767 , n76768 , n76769 , n76770 , n76771 , n76772 , n76773 , n76774 , 
 n76775 , n76776 , n76777 , n76778 , n76779 , n76780 , n76781 , n76782 , n76783 , n76784 , 
 n76785 , n76786 , n76787 , n76788 , n76789 , n76790 , n76791 , n76792 , n76793 , n76794 , 
 n76795 , n76796 , n76797 , n76798 , n76799 , n76800 , n76801 , n76802 , n76803 , n76804 , 
 n76805 , n76806 , n76807 , n76808 , n76809 , n76810 , n76811 , n76812 , n76813 , n76814 , 
 n76815 , n76816 , n76817 , n76818 , n76819 , n76820 , n76821 , n76822 , n76823 , n76824 , 
 n76825 , n76826 , n76827 , n76828 , n76829 , n76830 , n76831 , n76832 , n76833 , n76834 , 
 n76835 , n76836 , n76837 , n76838 , n76839 , n76840 , n76841 , n76842 , n76843 , n76844 , 
 n76845 , n76846 , n76847 , n76848 , n76849 , n76850 , n76851 , n76852 , n76853 , n76854 , 
 n76855 , n76856 , n76857 , n76858 , n76859 , n76860 , n76861 , n76862 , n76863 , n76864 , 
 n76865 , n76866 , n76867 , n76868 , n76869 , n76870 , n76871 , n76872 , n76873 , n76874 , 
 n76875 , n76876 , n76877 , n76878 , n76879 , n76880 , n76881 , n76882 , n76883 , n76884 , 
 n76885 , n76886 , n76887 , n76888 , n76889 , n76890 , n76891 , n76892 , n76893 , n76894 , 
 n76895 , n76896 , n76897 , n76898 , n76899 , n76900 , n76901 , n76902 , n76903 , n76904 , 
 n76905 , n76906 , n76907 , n76908 , n76909 , n76910 , n76911 , n76912 , n76913 , n76914 , 
 n76915 , n76916 , n76917 , n76918 , n76919 , n76920 , n76921 , n76922 , n76923 , n76924 , 
 n76925 , n76926 , n76927 , n76928 , n76929 , n76930 , n76931 , n76932 , n76933 , n76934 , 
 n76935 , n76936 , n76937 , n76938 , n76939 , n76940 , n76941 , n76942 , n76943 , n76944 , 
 n76945 , n76946 , n76947 , n76948 , n76949 , n76950 , n76951 , n76952 , n76953 , n76954 , 
 n76955 , n76956 , n76957 , n76958 , n76959 , n76960 , n76961 , n76962 , n76963 , n76964 , 
 n76965 , n76966 , n76967 , n76968 , n76969 , n76970 , n76971 , n76972 , n76973 , n76974 , 
 n76975 , n76976 , n76977 , n76978 , n76979 , n76980 , n76981 , n76982 , n76983 , n76984 , 
 n76985 , n76986 , n76987 , n76988 , n76989 , n76990 , n76991 , n76992 , n76993 , n76994 , 
 n76995 , n76996 , n76997 , n76998 , n76999 , n77000 , n77001 , n77002 , n77003 , n77004 , 
 n77005 , n77006 , n77007 , n77008 , n77009 , n77010 , n77011 , n77012 , n77013 , n77014 , 
 n77015 , n77016 , n77017 , n77018 , n77019 , n77020 , n77021 , n77022 , n77023 , n77024 , 
 n77025 , n77026 , n77027 , n77028 , n77029 , n77030 , n77031 , n77032 , n77033 , n77034 , 
 n77035 , n77036 , n77037 , n77038 , n77039 , n77040 , n77041 , n77042 , n77043 , n77044 , 
 n77045 , n77046 , n77047 , n77048 , n77049 , n77050 , n77051 , n77052 , n77053 , n77054 , 
 n77055 , n77056 , n77057 , n77058 , n77059 , n77060 , n77061 , n77062 , n77063 , n77064 , 
 n77065 , n77066 , n77067 , n77068 , n77069 , n77070 , n77071 , n77072 , n77073 , n77074 , 
 n77075 , n77076 , n77077 , n77078 , n77079 , n77080 , n77081 , n77082 , n77083 , n77084 , 
 n77085 , n77086 , n77087 , n77088 , n77089 , n77090 , n77091 , n77092 , n77093 , n77094 , 
 n77095 , n77096 , n77097 , n77098 , n77099 , n77100 , n77101 , n77102 , n77103 , n77104 , 
 n77105 , n77106 , n77107 , n77108 , n77109 , n77110 , n77111 , n77112 , n77113 , n77114 , 
 n77115 , n77116 , n77117 , n77118 , n77119 , n77120 , n77121 , n77122 , n77123 , n77124 , 
 n77125 , n77126 , n77127 , n77128 , n77129 , n77130 , n77131 , n77132 , n77133 , n77134 , 
 n77135 , n77136 , n77137 , n77138 , n77139 , n77140 , n77141 , n77142 , n77143 , n77144 , 
 n77145 , n77146 , n77147 , n77148 , n77149 , n77150 , n77151 , n77152 , n77153 , n77154 , 
 n77155 , n77156 , n77157 , n77158 , n77159 , n77160 , n77161 , n77162 , n77163 , n77164 , 
 n77165 , n77166 , n77167 , n77168 , n77169 , n77170 , n77171 , n77172 , n77173 , n77174 , 
 n77175 , n77176 , n77177 , n77178 , n77179 , n77180 , n77181 , n77182 , n77183 , n77184 , 
 n77185 , n77186 , n77187 , n77188 , n77189 , n77190 , n77191 , n77192 , n77193 , n77194 , 
 n77195 , n77196 , n77197 , n77198 , n77199 , n77200 , n77201 , n77202 , n77203 , n77204 , 
 n77205 , n77206 , n77207 , n77208 , n77209 , n77210 , n77211 , n77212 , n77213 , n77214 , 
 n77215 , n77216 , n77217 , n77218 , n77219 , n77220 , n77221 , n77222 , n77223 , n77224 , 
 n77225 , n77226 , n77227 , n77228 , n77229 , n77230 , n77231 , n77232 , n77233 , n77234 , 
 n77235 , n77236 , n77237 , n77238 , n77239 , n77240 , n77241 , n77242 , n77243 , n77244 , 
 n77245 , n77246 , n77247 , n77248 , n77249 , n77250 , n77251 , n77252 , n77253 , n77254 , 
 n77255 , n77256 , n77257 , n77258 , n77259 , n77260 , n77261 , n77262 , n77263 , n77264 , 
 n77265 , n77266 , n77267 , n77268 , n77269 , n77270 , n77271 , n77272 , n77273 , n77274 , 
 n77275 , n77276 , n77277 , n77278 , n77279 , n77280 , n77281 , n77282 , n77283 , n77284 , 
 n77285 , n77286 , n77287 , n77288 , n77289 , n77290 , n77291 , n77292 , n77293 , n77294 , 
 n77295 , n77296 , n77297 , n77298 , n77299 , n77300 , n77301 , n77302 , n77303 , n77304 , 
 n77305 , n77306 , n77307 , n77308 , n77309 , n77310 , n77311 , n77312 , n77313 , n77314 , 
 n77315 , n77316 , n77317 , n77318 , n77319 , n77320 , n77321 , n77322 , n77323 , n77324 , 
 n77325 , n77326 , n77327 , n77328 , n77329 , n77330 , n77331 , n77332 , n77333 , n77334 , 
 n77335 , n77336 , n77337 , n77338 , n77339 , n77340 , n77341 , n77342 , n77343 , n77344 , 
 n77345 , n77346 , n77347 , n77348 , n77349 , n77350 , n77351 , n77352 , n77353 , n77354 , 
 n77355 , n77356 , n77357 , n77358 , n77359 , n77360 , n77361 , n77362 , n77363 , n77364 , 
 n77365 , n77366 , n77367 , n77368 , n77369 , n77370 , n77371 , n77372 , n77373 , n77374 , 
 n77375 , n77376 , n77377 , n77378 , n77379 , n77380 , n77381 , n77382 , n77383 , n77384 , 
 n77385 , n77386 , n77387 , n77388 , n77389 , n77390 , n77391 , n77392 , n77393 , n77394 , 
 n77395 , n77396 , n77397 , n77398 , n77399 , n77400 , n77401 , n77402 , n77403 , n77404 , 
 n77405 , n77406 , n77407 , n77408 , n77409 , n77410 , n77411 , n77412 , n77413 , n77414 , 
 n77415 , n77416 , n77417 , n77418 , n77419 , n77420 , n77421 , n77422 , n77423 , n77424 , 
 n77425 , n77426 , n77427 , n77428 , n77429 , n77430 , n77431 , n77432 , n77433 , n77434 , 
 n77435 , n77436 , n77437 , n77438 , n77439 , n77440 , n77441 , n77442 , n77443 , n77444 , 
 n77445 , n77446 , n77447 , n77448 , n77449 , n77450 , n77451 , n77452 , n77453 , n77454 , 
 n77455 , n77456 , n77457 , n77458 , n77459 , n77460 , n77461 , n77462 , n77463 , n77464 , 
 n77465 , n77466 , n77467 , n77468 , n77469 , n77470 , n77471 , n77472 , n77473 , n77474 , 
 n77475 , n77476 , n77477 , n77478 , n77479 , n77480 , n77481 , n77482 , n77483 , n77484 , 
 n77485 , n77486 , n77487 , n77488 , n77489 , n77490 , n77491 , n77492 , n77493 , n77494 , 
 n77495 , n77496 , n77497 , n77498 , n77499 , n77500 , n77501 , n77502 , n77503 , n77504 , 
 n77505 , n77506 , n77507 , n77508 , n77509 , n77510 , n77511 , n77512 , n77513 , n77514 , 
 n77515 , n77516 , n77517 , n77518 , n77519 , n77520 , n77521 , n77522 , n77523 , n77524 , 
 n77525 , n77526 , n77527 , n77528 , n77529 , n77530 , n77531 , n77532 , n77533 , n77534 , 
 n77535 , n77536 , n77537 , n77538 , n77539 , n77540 , n77541 , n77542 , n77543 , n77544 , 
 n77545 , n77546 , n77547 , n77548 , n77549 , n77550 , n77551 , n77552 , n77553 , n77554 , 
 n77555 , n77556 , n77557 , n77558 , n77559 , n77560 , n77561 , n77562 , n77563 , n77564 , 
 n77565 , n77566 , n77567 , n77568 , n77569 , n77570 , n77571 , n77572 , n77573 , n77574 , 
 n77575 , n77576 , n77577 , n77578 , n77579 , n77580 , n77581 , n77582 , n77583 , n77584 , 
 n77585 , n77586 , n77587 , n77588 , n77589 , n77590 , n77591 , n77592 , n77593 , n77594 , 
 n77595 , n77596 , n77597 , n77598 , n77599 , n77600 , n77601 , n77602 , n77603 , n77604 , 
 n77605 , n77606 , n77607 , n77608 , n77609 , n77610 , n77611 , n77612 , n77613 , n77614 , 
 n77615 , n77616 , n77617 , n77618 , n77619 , n77620 , n77621 , n77622 , n77623 , n77624 , 
 n77625 , n77626 , n77627 , n77628 , n77629 , n77630 , n77631 , n77632 , n77633 , n77634 , 
 n77635 , n77636 , n77637 , n77638 , n77639 , n77640 , n77641 , n77642 , n77643 , n77644 , 
 n77645 , n77646 , n77647 , n77648 , n77649 , n77650 , n77651 , n77652 , n77653 , n77654 , 
 n77655 , n77656 , n77657 , n77658 , n77659 , n77660 , n77661 , n77662 , n77663 , n77664 , 
 n77665 , n77666 , n77667 , n77668 , n77669 , n77670 , n77671 , n77672 , n77673 , n77674 , 
 n77675 , n77676 , n77677 , n77678 , n77679 , n77680 , n77681 , n77682 , n77683 , n77684 , 
 n77685 , n77686 , n77687 , n77688 , n77689 , n77690 , n77691 , n77692 , n77693 , n77694 , 
 n77695 , n77696 , n77697 , n77698 , n77699 , n77700 , n77701 , n77702 , n77703 , n77704 , 
 n77705 , n77706 , n77707 , n77708 , n77709 , n77710 , n77711 , n77712 , n77713 , n77714 , 
 n77715 , n77716 , n77717 , n77718 , n77719 , n77720 , n77721 , n77722 , n77723 , n77724 , 
 n77725 , n77726 , n77727 , n77728 , n77729 , n77730 , n77731 , n77732 , n77733 , n77734 , 
 n77735 , n77736 , n77737 , n77738 , n77739 , n77740 , n77741 , n77742 , n77743 , n77744 , 
 n77745 , n77746 , n77747 , n77748 , n77749 , n77750 , n77751 , n77752 , n77753 , n77754 , 
 n77755 , n77756 , n77757 , n77758 , n77759 , n77760 , n77761 , n77762 , n77763 , n77764 , 
 n77765 , n77766 , n77767 , n77768 , n77769 , n77770 , n77771 , n77772 , n77773 , n77774 , 
 n77775 , n77776 , n77777 , n77778 , n77779 , n77780 , n77781 , n77782 , n77783 , n77784 , 
 n77785 , n77786 , n77787 , n77788 , n77789 , n77790 , n77791 , n77792 , n77793 , n77794 , 
 n77795 , n77796 , n77797 , n77798 , n77799 , n77800 , n77801 , n77802 , n77803 , n77804 , 
 n77805 , n77806 , n77807 , n77808 , n77809 , n77810 , n77811 , n77812 , n77813 , n77814 , 
 n77815 , n77816 , n77817 , n77818 , n77819 , n77820 , n77821 , n77822 , n77823 , n77824 , 
 n77825 , n77826 , n77827 , n77828 , n77829 , n77830 , n77831 , n77832 , n77833 , n77834 , 
 n77835 , n77836 , n77837 , n77838 , n77839 , n77840 , n77841 , n77842 , n77843 , n77844 , 
 n77845 , n77846 , n77847 , n77848 , n77849 , n77850 , n77851 , n77852 , n77853 , n77854 , 
 n77855 , n77856 , n77857 , n77858 , n77859 , n77860 , n77861 , n77862 , n77863 , n77864 , 
 n77865 , n77866 , n77867 , n77868 , n77869 , n77870 , n77871 , n77872 , n77873 , n77874 , 
 n77875 , n77876 , n77877 , n77878 , n77879 , n77880 , n77881 , n77882 , n77883 , n77884 , 
 n77885 , n77886 , n77887 , n77888 , n77889 , n77890 , n77891 , n77892 , n77893 , n77894 , 
 n77895 , n77896 , n77897 , n77898 , n77899 , n77900 , n77901 , n77902 , n77903 , n77904 , 
 n77905 , n77906 , n77907 , n77908 , n77909 , n77910 , n77911 , n77912 , n77913 , n77914 , 
 n77915 , n77916 , n77917 , n77918 , n77919 , n77920 , n77921 , n77922 , n77923 , n77924 , 
 n77925 , n77926 , n77927 , n77928 , n77929 , n77930 , n77931 , n77932 , n77933 , n77934 , 
 n77935 , n77936 , n77937 , n77938 , n77939 , n77940 , n77941 , n77942 , n77943 , n77944 , 
 n77945 , n77946 , n77947 , n77948 , n77949 , n77950 , n77951 , n77952 , n77953 , n77954 , 
 n77955 , n77956 , n77957 , n77958 , n77959 , n77960 , n77961 , n77962 , n77963 , n77964 , 
 n77965 , n77966 , n77967 , n77968 , n77969 , n77970 , n77971 , n77972 , n77973 , n77974 , 
 n77975 , n77976 , n77977 , n77978 , n77979 , n77980 , n77981 , n77982 , n77983 , n77984 , 
 n77985 , n77986 , n77987 , n77988 , n77989 , n77990 , n77991 , n77992 , n77993 , n77994 , 
 n77995 , n77996 , n77997 , n77998 , n77999 , n78000 , n78001 , n78002 , n78003 , n78004 , 
 n78005 , n78006 , n78007 , n78008 , n78009 , n78010 , n78011 , n78012 , n78013 , n78014 , 
 n78015 , n78016 , n78017 , n78018 , n78019 , n78020 , n78021 , n78022 , n78023 , n78024 , 
 n78025 , n78026 , n78027 , n78028 , n78029 , n78030 , n78031 , n78032 , n78033 , n78034 , 
 n78035 , n78036 , n78037 , n78038 , n78039 , n78040 , n78041 , n78042 , n78043 , n78044 , 
 n78045 , n78046 , n78047 , n78048 , n78049 , n78050 , n78051 , n78052 , n78053 , n78054 , 
 n78055 , n78056 , n78057 , n78058 , n78059 , n78060 , n78061 , n78062 , n78063 , n78064 , 
 n78065 , n78066 , n78067 , n78068 , n78069 , n78070 , n78071 , n78072 , n78073 , n78074 , 
 n78075 , n78076 , n78077 , n78078 , n78079 , n78080 , n78081 , n78082 , n78083 , n78084 , 
 n78085 , n78086 , n78087 , n78088 , n78089 , n78090 , n78091 , n78092 , n78093 , n78094 , 
 n78095 , n78096 , n78097 , n78098 , n78099 , n78100 , n78101 , n78102 , n78103 , n78104 , 
 n78105 , n78106 , n78107 , n78108 , n78109 , n78110 , n78111 , n78112 , n78113 , n78114 , 
 n78115 , n78116 , n78117 , n78118 , n78119 , n78120 , n78121 , n78122 , n78123 , n78124 , 
 n78125 , n78126 , n78127 , n78128 , n78129 , n78130 , n78131 , n78132 , n78133 , n78134 , 
 n78135 , n78136 , n78137 , n78138 , n78139 , n78140 , n78141 , n78142 , n78143 , n78144 , 
 n78145 , n78146 , n78147 , n78148 , n78149 , n78150 , n78151 , n78152 , n78153 , n78154 , 
 n78155 , n78156 , n78157 , n78158 , n78159 , n78160 , n78161 , n78162 , n78163 , n78164 , 
 n78165 , n78166 , n78167 , n78168 , n78169 , n78170 , n78171 , n78172 , n78173 , n78174 , 
 n78175 , n78176 , n78177 , n78178 , n78179 , n78180 , n78181 , n78182 , n78183 , n78184 , 
 n78185 , n78186 , n78187 , n78188 , n78189 , n78190 , n78191 , n78192 , n78193 , n78194 , 
 n78195 , n78196 , n78197 , n78198 , n78199 , n78200 , n78201 , n78202 , n78203 , n78204 , 
 n78205 , n78206 , n78207 , n78208 , n78209 , n78210 , n78211 , n78212 , n78213 , n78214 , 
 n78215 , n78216 , n78217 , n78218 , n78219 , n78220 , n78221 , n78222 , n78223 , n78224 , 
 n78225 , n78226 , n78227 , n78228 , n78229 , n78230 , n78231 , n78232 , n78233 , n78234 , 
 n78235 , n78236 , n78237 , n78238 , n78239 , n78240 , n78241 , n78242 , n78243 , n78244 , 
 n78245 , n78246 , n78247 , n78248 , n78249 , n78250 , n78251 , n78252 , n78253 , n78254 , 
 n78255 , n78256 , n78257 , n78258 , n78259 , n78260 , n78261 , n78262 , n78263 , n78264 , 
 n78265 , n78266 , n78267 , n78268 , n78269 , n78270 , n78271 , n78272 , n78273 , n78274 , 
 n78275 , n78276 , n78277 , n78278 , n78279 , n78280 , n78281 , n78282 , n78283 , n78284 , 
 n78285 , n78286 , n78287 , n78288 , n78289 , n78290 , n78291 , n78292 , n78293 , n78294 , 
 n78295 , n78296 , n78297 , n78298 , n78299 , n78300 , n78301 , n78302 , n78303 , n78304 , 
 n78305 , n78306 , n78307 , n78308 , n78309 , n78310 , n78311 , n78312 , n78313 , n78314 , 
 n78315 , n78316 , n78317 , n78318 , n78319 , n78320 , n78321 , n78322 , n78323 , n78324 , 
 n78325 , n78326 , n78327 , n78328 , n78329 , n78330 , n78331 , n78332 , n78333 , n78334 , 
 n78335 , n78336 , n78337 , n78338 , n78339 , n78340 , n78341 , n78342 , n78343 , n78344 , 
 n78345 , n78346 , n78347 , n78348 , n78349 , n78350 , n78351 , n78352 , n78353 , n78354 , 
 n78355 , n78356 , n78357 , n78358 , n78359 , n78360 , n78361 , n78362 , n78363 , n78364 , 
 n78365 , n78366 , n78367 , n78368 , n78369 , n78370 , n78371 , n78372 , n78373 , n78374 , 
 n78375 , n78376 , n78377 , n78378 , n78379 , n78380 , n78381 , n78382 , n78383 , n78384 , 
 n78385 , n78386 , n78387 , n78388 , n78389 , n78390 , n78391 , n78392 , n78393 , n78394 , 
 n78395 , n78396 , n78397 , n78398 , n78399 , n78400 , n78401 , n78402 , n78403 , n78404 , 
 n78405 , n78406 , n78407 , n78408 , n78409 , n78410 , n78411 , n78412 , n78413 , n78414 , 
 n78415 , n78416 , n78417 , n78418 , n78419 , n78420 , n78421 , n78422 , n78423 , n78424 , 
 n78425 , n78426 , n78427 , n78428 , n78429 , n78430 , n78431 , n78432 , n78433 , n78434 , 
 n78435 , n78436 , n78437 , n78438 , n78439 , n78440 , n78441 , n78442 , n78443 , n78444 , 
 n78445 , n78446 , n78447 , n78448 , n78449 , n78450 , n78451 , n78452 , n78453 , n78454 , 
 n78455 , n78456 , n78457 , n78458 , n78459 , n78460 , n78461 , n78462 , n78463 , n78464 , 
 n78465 , n78466 , n78467 , n78468 , n78469 , n78470 , n78471 , n78472 , n78473 , n78474 , 
 n78475 , n78476 , n78477 , n78478 , n78479 , n78480 , n78481 , n78482 , n78483 , n78484 , 
 n78485 , n78486 , n78487 , n78488 , n78489 , n78490 , n78491 , n78492 , n78493 , n78494 , 
 n78495 , n78496 , n78497 , n78498 , n78499 , n78500 , n78501 , n78502 , n78503 , n78504 , 
 n78505 , n78506 , n78507 , n78508 , n78509 , n78510 , n78511 , n78512 , n78513 , n78514 , 
 n78515 , n78516 , n78517 , n78518 , n78519 , n78520 , n78521 , n78522 , n78523 , n78524 , 
 n78525 , n78526 , n78527 , n78528 , n78529 , n78530 , n78531 , n78532 , n78533 , n78534 , 
 n78535 , n78536 , n78537 , n78538 , n78539 , n78540 , n78541 , n78542 , n78543 , n78544 , 
 n78545 , n78546 , n78547 , n78548 , n78549 , n78550 , n78551 , n78552 , n78553 , n78554 , 
 n78555 , n78556 , n78557 , n78558 , n78559 , n78560 , n78561 , n78562 , n78563 , n78564 , 
 n78565 , n78566 , n78567 , n78568 , n78569 , n78570 , n78571 , n78572 , n78573 , n78574 , 
 n78575 , n78576 , n78577 , n78578 , n78579 , n78580 , n78581 , n78582 , n78583 , n78584 , 
 n78585 , n78586 , n78587 , n78588 , n78589 , n78590 , n78591 , n78592 , n78593 , n78594 , 
 n78595 , n78596 , n78597 , n78598 , n78599 , n78600 , n78601 , n78602 , n78603 , n78604 , 
 n78605 , n78606 , n78607 , n78608 , n78609 , n78610 , n78611 , n78612 , n78613 , n78614 , 
 n78615 , n78616 , n78617 , n78618 , n78619 , n78620 , n78621 , n78622 , n78623 , n78624 , 
 n78625 , n78626 , n78627 , n78628 , n78629 , n78630 , n78631 , n78632 , n78633 , n78634 , 
 n78635 , n78636 , n78637 , n78638 , n78639 , n78640 , n78641 , n78642 , n78643 , n78644 , 
 n78645 , n78646 , n78647 , n78648 , n78649 , n78650 , n78651 , n78652 , n78653 , n78654 , 
 n78655 , n78656 , n78657 , n78658 , n78659 , n78660 , n78661 , n78662 , n78663 , n78664 , 
 n78665 , n78666 , n78667 , n78668 , n78669 , n78670 , n78671 , n78672 , n78673 , n78674 , 
 n78675 , n78676 , n78677 , n78678 , n78679 , n78680 , n78681 , n78682 , n78683 , n78684 , 
 n78685 , n78686 , n78687 , n78688 , n78689 , n78690 , n78691 , n78692 , n78693 , n78694 , 
 n78695 , n78696 , n78697 , n78698 , n78699 , n78700 , n78701 , n78702 , n78703 , n78704 , 
 n78705 , n78706 , n78707 , n78708 , n78709 , n78710 , n78711 , n78712 , n78713 , n78714 , 
 n78715 , n78716 , n78717 , n78718 , n78719 , n78720 , n78721 , n78722 , n78723 , n78724 , 
 n78725 , n78726 , n78727 , n78728 , n78729 , n78730 , n78731 , n78732 , n78733 , n78734 , 
 n78735 , n78736 , n78737 , n78738 , n78739 , n78740 , n78741 , n78742 , n78743 , n78744 , 
 n78745 , n78746 , n78747 , n78748 , n78749 , n78750 , n78751 , n78752 , n78753 , n78754 , 
 n78755 , n78756 , n78757 , n78758 , n78759 , n78760 , n78761 , n78762 , n78763 , n78764 , 
 n78765 , n78766 , n78767 , n78768 , n78769 , n78770 , n78771 , n78772 , n78773 , n78774 , 
 n78775 , n78776 , n78777 , n78778 , n78779 , n78780 , n78781 , n78782 , n78783 , n78784 , 
 n78785 , n78786 , n78787 , n78788 , n78789 , n78790 , n78791 , n78792 , n78793 , n78794 , 
 n78795 , n78796 , n78797 , n78798 , n78799 , n78800 , n78801 , n78802 , n78803 , n78804 , 
 n78805 , n78806 , n78807 , n78808 , n78809 , n78810 , n78811 , n78812 , n78813 , n78814 , 
 n78815 , n78816 , n78817 , n78818 , n78819 , n78820 , n78821 , n78822 , n78823 , n78824 , 
 n78825 , n78826 , n78827 , n78828 , n78829 , n78830 , n78831 , n78832 , n78833 , n78834 , 
 n78835 , n78836 , n78837 , n78838 , n78839 , n78840 , n78841 , n78842 , n78843 , n78844 , 
 n78845 , n78846 , n78847 , n78848 , n78849 , n78850 , n78851 , n78852 , n78853 , n78854 , 
 n78855 , n78856 , n78857 , n78858 , n78859 , n78860 , n78861 , n78862 , n78863 , n78864 , 
 n78865 , n78866 , n78867 , n78868 , n78869 , n78870 , n78871 , n78872 , n78873 , n78874 , 
 n78875 , n78876 , n78877 , n78878 , n78879 , n78880 , n78881 , n78882 , n78883 , n78884 , 
 n78885 , n78886 , n78887 , n78888 , n78889 , n78890 , n78891 , n78892 , n78893 , n78894 , 
 n78895 , n78896 , n78897 , n78898 , n78899 , n78900 , n78901 , n78902 , n78903 , n78904 , 
 n78905 , n78906 , n78907 , n78908 , n78909 , n78910 , n78911 , n78912 , n78913 , n78914 , 
 n78915 , n78916 , n78917 , n78918 , n78919 , n78920 , n78921 , n78922 , n78923 , n78924 , 
 n78925 , n78926 , n78927 , n78928 , n78929 , n78930 , n78931 , n78932 , n78933 , n78934 , 
 n78935 , n78936 , n78937 , n78938 , n78939 , n78940 , n78941 , n78942 , n78943 , n78944 , 
 n78945 , n78946 , n78947 , n78948 , n78949 , n78950 , n78951 , n78952 , n78953 , n78954 , 
 n78955 , n78956 , n78957 , n78958 , n78959 , n78960 , n78961 , n78962 , n78963 , n78964 , 
 n78965 , n78966 , n78967 , n78968 , n78969 , n78970 , n78971 , n78972 , n78973 , n78974 , 
 n78975 , n78976 , n78977 , n78978 , n78979 , n78980 , n78981 , n78982 , n78983 , n78984 , 
 n78985 , n78986 , n78987 , n78988 , n78989 , n78990 , n78991 , n78992 , n78993 , n78994 , 
 n78995 , n78996 , n78997 , n78998 , n78999 , n79000 , n79001 , n79002 , n79003 , n79004 , 
 n79005 , n79006 , n79007 , n79008 , n79009 , n79010 , n79011 , n79012 , n79013 , n79014 , 
 n79015 , n79016 , n79017 , n79018 , n79019 , n79020 , n79021 , n79022 , n79023 , n79024 , 
 n79025 , n79026 , n79027 , n79028 , n79029 , n79030 , n79031 , n79032 , n79033 , n79034 , 
 n79035 , n79036 , n79037 , n79038 , n79039 , n79040 , n79041 , n79042 , n79043 , n79044 , 
 n79045 , n79046 , n79047 , n79048 , n79049 , n79050 , n79051 , n79052 , n79053 , n79054 , 
 n79055 , n79056 , n79057 , n79058 , n79059 , n79060 , n79061 , n79062 , n79063 , n79064 , 
 n79065 , n79066 , n79067 , n79068 , n79069 , n79070 , n79071 , n79072 , n79073 , n79074 , 
 n79075 , n79076 , n79077 , n79078 , n79079 , n79080 , n79081 , n79082 , n79083 , n79084 , 
 n79085 , n79086 , n79087 , n79088 , n79089 , n79090 , n79091 , n79092 , n79093 , n79094 , 
 n79095 , n79096 , n79097 , n79098 , n79099 , n79100 , n79101 , n79102 , n79103 , n79104 , 
 n79105 , n79106 , n79107 , n79108 , n79109 , n79110 , n79111 , n79112 , n79113 , n79114 , 
 n79115 , n79116 , n79117 , n79118 , n79119 , n79120 , n79121 , n79122 , n79123 , n79124 , 
 n79125 , n79126 , n79127 , n79128 , n79129 , n79130 , n79131 , n79132 , n79133 , n79134 , 
 n79135 , n79136 , n79137 , n79138 , n79139 , n79140 , n79141 , n79142 , n79143 , n79144 , 
 n79145 , n79146 , n79147 , n79148 , n79149 , n79150 , n79151 , n79152 , n79153 , n79154 , 
 n79155 , n79156 , n79157 , n79158 , n79159 , n79160 , n79161 , n79162 , n79163 , n79164 , 
 n79165 , n79166 , n79167 , n79168 , n79169 , n79170 , n79171 , n79172 , n79173 , n79174 , 
 n79175 , n79176 , n79177 , n79178 , n79179 , n79180 , n79181 , n79182 , n79183 , n79184 , 
 n79185 , n79186 , n79187 , n79188 , n79189 , n79190 , n79191 , n79192 , n79193 , n79194 , 
 n79195 , n79196 , n79197 , n79198 , n79199 , n79200 , n79201 , n79202 , n79203 , n79204 , 
 n79205 , n79206 , n79207 , n79208 , n79209 , n79210 , n79211 , n79212 , n79213 , n79214 , 
 n79215 , n79216 , n79217 , n79218 , n79219 , n79220 , n79221 , n79222 , n79223 , n79224 , 
 n79225 , n79226 , n79227 , n79228 , n79229 , n79230 , n79231 , n79232 , n79233 , n79234 , 
 n79235 , n79236 , n79237 , n79238 , n79239 , n79240 , n79241 , n79242 , n79243 , n79244 , 
 n79245 , n79246 , n79247 , n79248 , n79249 , n79250 , n79251 , n79252 , n79253 , n79254 , 
 n79255 , n79256 , n79257 , n79258 , n79259 , n79260 , n79261 , n79262 , n79263 , n79264 , 
 n79265 , n79266 , n79267 , n79268 , n79269 , n79270 , n79271 , n79272 , n79273 , n79274 , 
 n79275 , n79276 , n79277 , n79278 , n79279 , n79280 , n79281 , n79282 , n79283 , n79284 , 
 n79285 , n79286 , n79287 , n79288 , n79289 , n79290 , n79291 , n79292 , n79293 , n79294 , 
 n79295 , n79296 , n79297 , n79298 , n79299 , n79300 , n79301 , n79302 , n79303 , n79304 , 
 n79305 , n79306 , n79307 , n79308 , n79309 , n79310 , n79311 , n79312 , n79313 , n79314 , 
 n79315 , n79316 , n79317 , n79318 , n79319 , n79320 , n79321 , n79322 , n79323 , n79324 , 
 n79325 , n79326 , n79327 , n79328 , n79329 , n79330 , n79331 , n79332 , n79333 , n79334 , 
 n79335 , n79336 , n79337 , n79338 , n79339 , n79340 , n79341 , n79342 , n79343 , n79344 , 
 n79345 , n79346 , n79347 , n79348 , n79349 , n79350 , n79351 , n79352 , n79353 , n79354 , 
 n79355 , n79356 , n79357 , n79358 , n79359 , n79360 , n79361 , n79362 , n79363 , n79364 , 
 n79365 , n79366 , n79367 , n79368 , n79369 , n79370 , n79371 , n79372 , n79373 , n79374 , 
 n79375 , n79376 , n79377 , n79378 , n79379 , n79380 , n79381 , n79382 , n79383 , n79384 , 
 n79385 , n79386 , n79387 , n79388 , n79389 , n79390 , n79391 , n79392 , n79393 , n79394 , 
 n79395 , n79396 , n79397 , n79398 , n79399 , n79400 , n79401 , n79402 , n79403 , n79404 , 
 n79405 , n79406 , n79407 , n79408 , n79409 , n79410 , n79411 , n79412 , n79413 , n79414 , 
 n79415 , n79416 , n79417 , n79418 , n79419 , n79420 , n79421 , n79422 , n79423 , n79424 , 
 n79425 , n79426 , n79427 , n79428 , n79429 , n79430 , n79431 , n79432 , n79433 , n79434 , 
 n79435 , n79436 , n79437 , n79438 , n79439 , n79440 , n79441 , n79442 , n79443 , n79444 , 
 n79445 , n79446 , n79447 , n79448 , n79449 , n79450 , n79451 , n79452 , n79453 , n79454 , 
 n79455 , n79456 , n79457 , n79458 , n79459 , n79460 , n79461 , n79462 , n79463 , n79464 , 
 n79465 , n79466 , n79467 , n79468 , n79469 , n79470 , n79471 , n79472 , n79473 , n79474 , 
 n79475 , n79476 , n79477 , n79478 , n79479 , n79480 , n79481 , n79482 , n79483 , n79484 , 
 n79485 , n79486 , n79487 , n79488 , n79489 , n79490 , n79491 , n79492 , n79493 , n79494 , 
 n79495 , n79496 , n79497 , n79498 , n79499 , n79500 , n79501 , n79502 , n79503 , n79504 , 
 n79505 , n79506 , n79507 , n79508 , n79509 , n79510 , n79511 , n79512 , n79513 , n79514 , 
 n79515 , n79516 , n79517 , n79518 , n79519 , n79520 , n79521 , n79522 , n79523 , n79524 , 
 n79525 , n79526 , n79527 , n79528 , n79529 , n79530 , n79531 , n79532 , n79533 , n79534 , 
 n79535 , n79536 , n79537 , n79538 , n79539 , n79540 , n79541 , n79542 , n79543 , n79544 , 
 n79545 , n79546 , n79547 , n79548 , n79549 , n79550 , n79551 , n79552 , n79553 , n79554 , 
 n79555 , n79556 , n79557 , n79558 , n79559 , n79560 , n79561 , n79562 , n79563 , n79564 , 
 n79565 , n79566 , n79567 , n79568 , n79569 , n79570 , n79571 , n79572 , n79573 , n79574 , 
 n79575 , n79576 , n79577 , n79578 , n79579 , n79580 , n79581 , n79582 , n79583 , n79584 , 
 n79585 , n79586 , n79587 , n79588 , n79589 , n79590 , n79591 , n79592 , n79593 , n79594 , 
 n79595 , n79596 , n79597 , n79598 , n79599 , n79600 , n79601 , n79602 , n79603 , n79604 , 
 n79605 , n79606 , n79607 , n79608 , n79609 , n79610 , n79611 , n79612 , n79613 , n79614 , 
 n79615 , n79616 , n79617 , n79618 , n79619 , n79620 , n79621 , n79622 , n79623 , n79624 , 
 n79625 , n79626 , n79627 , n79628 , n79629 , n79630 , n79631 , n79632 , n79633 , n79634 , 
 n79635 , n79636 , n79637 , n79638 , n79639 , n79640 , n79641 , n79642 , n79643 , n79644 , 
 n79645 , n79646 , n79647 , n79648 , n79649 , n79650 , n79651 , n79652 , n79653 , n79654 , 
 n79655 , n79656 , n79657 , n79658 , n79659 , n79660 , n79661 , n79662 , n79663 , n79664 , 
 n79665 , n79666 , n79667 , n79668 , n79669 , n79670 , n79671 , n79672 , n79673 , n79674 , 
 n79675 , n79676 , n79677 , n79678 , n79679 , n79680 , n79681 , n79682 , n79683 , n79684 , 
 n79685 , n79686 , n79687 , n79688 , n79689 , n79690 , n79691 , n79692 , n79693 , n79694 , 
 n79695 , n79696 , n79697 , n79698 , n79699 , n79700 , n79701 , n79702 , n79703 , n79704 , 
 n79705 , n79706 , n79707 , n79708 , n79709 , n79710 , n79711 , n79712 , n79713 , n79714 , 
 n79715 , n79716 , n79717 , n79718 , n79719 , n79720 , n79721 , n79722 , n79723 , n79724 , 
 n79725 , n79726 , n79727 , n79728 , n79729 , n79730 , n79731 , n79732 , n79733 , n79734 , 
 n79735 , n79736 , n79737 , n79738 , n79739 , n79740 , n79741 , n79742 , n79743 , n79744 , 
 n79745 , n79746 , n79747 , n79748 , n79749 , n79750 , n79751 , n79752 , n79753 , n79754 , 
 n79755 , n79756 , n79757 , n79758 , n79759 , n79760 , n79761 , n79762 , n79763 , n79764 , 
 n79765 , n79766 , n79767 , n79768 , n79769 , n79770 , n79771 , n79772 , n79773 , n79774 , 
 n79775 , n79776 , n79777 , n79778 , n79779 , n79780 , n79781 , n79782 , n79783 , n79784 , 
 n79785 , n79786 , n79787 , n79788 , n79789 , n79790 , n79791 , n79792 , n79793 , n79794 , 
 n79795 , n79796 , n79797 , n79798 , n79799 , n79800 , n79801 , n79802 , n79803 , n79804 , 
 n79805 , n79806 , n79807 , n79808 , n79809 , n79810 , n79811 , n79812 , n79813 , n79814 , 
 n79815 , n79816 , n79817 , n79818 , n79819 , n79820 , n79821 , n79822 , n79823 , n79824 , 
 n79825 , n79826 , n79827 , n79828 , n79829 , n79830 , n79831 , n79832 , n79833 , n79834 , 
 n79835 , n79836 , n79837 , n79838 , n79839 , n79840 , n79841 , n79842 , n79843 , n79844 , 
 n79845 , n79846 , n79847 , n79848 , n79849 , n79850 , n79851 , n79852 , n79853 , n79854 , 
 n79855 , n79856 , n79857 , n79858 , n79859 , n79860 , n79861 , n79862 , n79863 , n79864 , 
 n79865 , n79866 , n79867 , n79868 , n79869 , n79870 , n79871 , n79872 , n79873 , n79874 , 
 n79875 , n79876 , n79877 , n79878 , n79879 , n79880 , n79881 , n79882 , n79883 , n79884 , 
 n79885 , n79886 , n79887 , n79888 , n79889 , n79890 , n79891 , n79892 , n79893 , n79894 , 
 n79895 , n79896 , n79897 , n79898 , n79899 , n79900 , n79901 , n79902 , n79903 , n79904 , 
 n79905 , n79906 , n79907 , n79908 , n79909 , n79910 , n79911 , n79912 , n79913 , n79914 , 
 n79915 , n79916 , n79917 , n79918 , n79919 , n79920 , n79921 , n79922 , n79923 , n79924 , 
 n79925 , n79926 , n79927 , n79928 , n79929 , n79930 , n79931 , n79932 , n79933 , n79934 , 
 n79935 , n79936 , n79937 , n79938 , n79939 , n79940 , n79941 , n79942 , n79943 , n79944 , 
 n79945 , n79946 , n79947 , n79948 , n79949 , n79950 , n79951 , n79952 , n79953 , n79954 , 
 n79955 , n79956 , n79957 , n79958 , n79959 , n79960 , n79961 , n79962 , n79963 , n79964 , 
 n79965 , n79966 , n79967 , n79968 , n79969 , n79970 , n79971 , n79972 , n79973 , n79974 , 
 n79975 , n79976 , n79977 , n79978 , n79979 , n79980 , n79981 , n79982 , n79983 , n79984 , 
 n79985 , n79986 , n79987 , n79988 , n79989 , n79990 , n79991 , n79992 , n79993 , n79994 , 
 n79995 , n79996 , n79997 , n79998 , n79999 , n80000 , n80001 , n80002 , n80003 , n80004 , 
 n80005 , n80006 , n80007 , n80008 , n80009 , n80010 , n80011 , n80012 , n80013 , n80014 , 
 n80015 , n80016 , n80017 , n80018 , n80019 , n80020 , n80021 , n80022 , n80023 , n80024 , 
 n80025 , n80026 , n80027 , n80028 , n80029 , n80030 , n80031 , n80032 , n80033 , n80034 , 
 n80035 , n80036 , n80037 , n80038 , n80039 , n80040 , n80041 , n80042 , n80043 , n80044 , 
 n80045 , n80046 , n80047 , n80048 , n80049 , n80050 , n80051 , n80052 , n80053 , n80054 , 
 n80055 , n80056 , n80057 , n80058 , n80059 , n80060 , n80061 , n80062 , n80063 , n80064 , 
 n80065 , n80066 , n80067 , n80068 , n80069 , n80070 , n80071 , n80072 , n80073 , n80074 , 
 n80075 , n80076 , n80077 , n80078 , n80079 , n80080 , n80081 , n80082 , n80083 , n80084 , 
 n80085 , n80086 , n80087 , n80088 , n80089 , n80090 , n80091 , n80092 , n80093 , n80094 , 
 n80095 , n80096 , n80097 , n80098 , n80099 , n80100 , n80101 , n80102 , n80103 , n80104 , 
 n80105 , n80106 , n80107 , n80108 , n80109 , n80110 , n80111 , n80112 , n80113 , n80114 , 
 n80115 , n80116 , n80117 , n80118 , n80119 , n80120 , n80121 , n80122 , n80123 , n80124 , 
 n80125 , n80126 , n80127 , n80128 , n80129 , n80130 , n80131 , n80132 , n80133 , n80134 , 
 n80135 , n80136 , n80137 , n80138 , n80139 , n80140 , n80141 , n80142 , n80143 , n80144 , 
 n80145 , n80146 , n80147 , n80148 , n80149 , n80150 , n80151 , n80152 , n80153 , n80154 , 
 n80155 , n80156 , n80157 , n80158 , n80159 , n80160 , n80161 , n80162 , n80163 , n80164 , 
 n80165 , n80166 , n80167 , n80168 , n80169 , n80170 , n80171 , n80172 , n80173 , n80174 , 
 n80175 , n80176 , n80177 , n80178 , n80179 , n80180 , n80181 , n80182 , n80183 , n80184 , 
 n80185 , n80186 , n80187 , n80188 , n80189 , n80190 , n80191 , n80192 , n80193 , n80194 , 
 n80195 , n80196 , n80197 , n80198 , n80199 , n80200 , n80201 , n80202 , n80203 , n80204 , 
 n80205 , n80206 , n80207 , n80208 , n80209 , n80210 , n80211 , n80212 , n80213 , n80214 , 
 n80215 , n80216 , n80217 , n80218 , n80219 , n80220 , n80221 , n80222 , n80223 , n80224 , 
 n80225 , n80226 , n80227 , n80228 , n80229 , n80230 , n80231 , n80232 , n80233 , n80234 , 
 n80235 , n80236 , n80237 , n80238 , n80239 , n80240 , n80241 , n80242 , n80243 , n80244 , 
 n80245 , n80246 , n80247 , n80248 , n80249 , n80250 , n80251 , n80252 , n80253 , n80254 , 
 n80255 , n80256 , n80257 , n80258 , n80259 , n80260 , n80261 , n80262 , n80263 , n80264 , 
 n80265 , n80266 , n80267 , n80268 , n80269 , n80270 , n80271 , n80272 , n80273 , n80274 , 
 n80275 , n80276 , n80277 , n80278 , n80279 , n80280 , n80281 , n80282 , n80283 , n80284 , 
 n80285 , n80286 , n80287 , n80288 , n80289 , n80290 , n80291 , n80292 , n80293 , n80294 , 
 n80295 , n80296 , n80297 , n80298 , n80299 , n80300 , n80301 , n80302 , n80303 , n80304 , 
 n80305 , n80306 , n80307 , n80308 , n80309 , n80310 , n80311 , n80312 , n80313 , n80314 , 
 n80315 , n80316 , n80317 , n80318 , n80319 , n80320 , n80321 , n80322 , n80323 , n80324 , 
 n80325 , n80326 , n80327 , n80328 , n80329 , n80330 , n80331 , n80332 , n80333 , n80334 , 
 n80335 , n80336 , n80337 , n80338 , n80339 , n80340 , n80341 , n80342 , n80343 , n80344 , 
 n80345 , n80346 , n80347 , n80348 , n80349 , n80350 , n80351 , n80352 , n80353 , n80354 , 
 n80355 , n80356 , n80357 , n80358 , n80359 , n80360 , n80361 , n80362 , n80363 , n80364 , 
 n80365 , n80366 , n80367 , n80368 , n80369 , n80370 , n80371 , n80372 , n80373 , n80374 , 
 n80375 , n80376 , n80377 , n80378 , n80379 , n80380 , n80381 , n80382 , n80383 , n80384 , 
 n80385 , n80386 , n80387 , n80388 , n80389 , n80390 , n80391 , n80392 , n80393 , n80394 , 
 n80395 , n80396 , n80397 , n80398 , n80399 , n80400 , n80401 , n80402 , n80403 , n80404 , 
 n80405 , n80406 , n80407 , n80408 , n80409 , n80410 , n80411 , n80412 , n80413 , n80414 , 
 n80415 , n80416 , n80417 , n80418 , n80419 , n80420 , n80421 , n80422 , n80423 , n80424 , 
 n80425 , n80426 , n80427 , n80428 , n80429 , n80430 , n80431 , n80432 , n80433 , n80434 , 
 n80435 , n80436 , n80437 , n80438 , n80439 , n80440 , n80441 , n80442 , n80443 , n80444 , 
 n80445 , n80446 , n80447 , n80448 , n80449 , n80450 , n80451 , n80452 , n80453 , n80454 , 
 n80455 , n80456 , n80457 , n80458 , n80459 , n80460 , n80461 , n80462 , n80463 , n80464 , 
 n80465 , n80466 , n80467 , n80468 , n80469 , n80470 , n80471 , n80472 , n80473 , n80474 , 
 n80475 , n80476 , n80477 , n80478 , n80479 , n80480 , n80481 , n80482 , n80483 , n80484 , 
 n80485 , n80486 , n80487 , n80488 , n80489 , n80490 , n80491 , n80492 , n80493 , n80494 , 
 n80495 , n80496 , n80497 , n80498 , n80499 , n80500 , n80501 , n80502 , n80503 , n80504 , 
 n80505 , n80506 , n80507 , n80508 , n80509 , n80510 , n80511 , n80512 , n80513 , n80514 , 
 n80515 , n80516 , n80517 , n80518 , n80519 , n80520 , n80521 , n80522 , n80523 , n80524 , 
 n80525 , n80526 , n80527 , n80528 , n80529 , n80530 , n80531 , n80532 , n80533 , n80534 , 
 n80535 , n80536 , n80537 , n80538 , n80539 , n80540 , n80541 , n80542 , n80543 , n80544 , 
 n80545 , n80546 , n80547 , n80548 , n80549 , n80550 , n80551 , n80552 , n80553 , n80554 , 
 n80555 , n80556 , n80557 , n80558 , n80559 , n80560 , n80561 , n80562 , n80563 , n80564 , 
 n80565 , n80566 , n80567 , n80568 , n80569 , n80570 , n80571 , n80572 , n80573 , n80574 , 
 n80575 , n80576 , n80577 , n80578 , n80579 , n80580 , n80581 , n80582 , n80583 , n80584 , 
 n80585 , n80586 , n80587 , n80588 , n80589 , n80590 , n80591 , n80592 , n80593 , n80594 , 
 n80595 , n80596 , n80597 , n80598 , n80599 , n80600 , n80601 , n80602 , n80603 , n80604 , 
 n80605 , n80606 , n80607 , n80608 , n80609 , n80610 , n80611 , n80612 , n80613 , n80614 , 
 n80615 , n80616 , n80617 , n80618 , n80619 , n80620 , n80621 , n80622 , n80623 , n80624 , 
 n80625 , n80626 , n80627 , n80628 , n80629 , n80630 , n80631 , n80632 , n80633 , n80634 , 
 n80635 , n80636 , n80637 , n80638 , n80639 , n80640 , n80641 , n80642 , n80643 , n80644 , 
 n80645 , n80646 , n80647 , n80648 , n80649 , n80650 , n80651 , n80652 , n80653 , n80654 , 
 n80655 , n80656 , n80657 , n80658 , n80659 , n80660 , n80661 , n80662 , n80663 , n80664 , 
 n80665 , n80666 , n80667 , n80668 , n80669 , n80670 , n80671 , n80672 , n80673 , n80674 , 
 n80675 , n80676 , n80677 , n80678 , n80679 , n80680 , n80681 , n80682 , n80683 , n80684 , 
 n80685 , n80686 , n80687 , n80688 , n80689 , n80690 , n80691 , n80692 , n80693 , n80694 , 
 n80695 , n80696 , n80697 , n80698 , n80699 , n80700 , n80701 , n80702 , n80703 , n80704 , 
 n80705 , n80706 , n80707 , n80708 , n80709 , n80710 , n80711 , n80712 , n80713 , n80714 , 
 n80715 , n80716 , n80717 , n80718 , n80719 , n80720 , n80721 , n80722 , n80723 , n80724 , 
 n80725 , n80726 , n80727 , n80728 , n80729 , n80730 , n80731 , n80732 , n80733 , n80734 , 
 n80735 , n80736 , n80737 , n80738 , n80739 , n80740 , n80741 , n80742 , n80743 , n80744 , 
 n80745 , n80746 , n80747 , n80748 , n80749 , n80750 , n80751 , n80752 , n80753 , n80754 , 
 n80755 , n80756 , n80757 , n80758 , n80759 , n80760 , n80761 , n80762 , n80763 , n80764 , 
 n80765 , n80766 , n80767 , n80768 , n80769 , n80770 , n80771 , n80772 , n80773 , n80774 , 
 n80775 , n80776 , n80777 , n80778 , n80779 , n80780 , n80781 , n80782 , n80783 , n80784 , 
 n80785 , n80786 , n80787 , n80788 , n80789 , n80790 , n80791 , n80792 , n80793 , n80794 , 
 n80795 , n80796 , n80797 , n80798 , n80799 , n80800 , n80801 , n80802 , n80803 , n80804 , 
 n80805 , n80806 , n80807 , n80808 , n80809 , n80810 , n80811 , n80812 , n80813 , n80814 , 
 n80815 , n80816 , n80817 , n80818 , n80819 , n80820 , n80821 , n80822 , n80823 , n80824 , 
 n80825 , n80826 , n80827 , n80828 , n80829 , n80830 , n80831 , n80832 , n80833 , n80834 , 
 n80835 , n80836 , n80837 , n80838 , n80839 , n80840 , n80841 , n80842 , n80843 , n80844 , 
 n80845 , n80846 , n80847 , n80848 , n80849 , n80850 , n80851 , n80852 , n80853 , n80854 , 
 n80855 , n80856 , n80857 , n80858 , n80859 , n80860 , n80861 , n80862 , n80863 , n80864 , 
 n80865 , n80866 , n80867 , n80868 , n80869 , n80870 , n80871 , n80872 , n80873 , n80874 , 
 n80875 , n80876 , n80877 , n80878 , n80879 , n80880 , n80881 , n80882 , n80883 , n80884 , 
 n80885 , n80886 , n80887 , n80888 , n80889 , n80890 , n80891 , n80892 , n80893 , n80894 , 
 n80895 , n80896 , n80897 , n80898 , n80899 , n80900 , n80901 , n80902 , n80903 , n80904 , 
 n80905 , n80906 , n80907 , n80908 , n80909 , n80910 , n80911 , n80912 , n80913 , n80914 , 
 n80915 , n80916 , n80917 , n80918 , n80919 , n80920 , n80921 , n80922 , n80923 , n80924 , 
 n80925 , n80926 , n80927 , n80928 , n80929 , n80930 , n80931 , n80932 , n80933 , n80934 , 
 n80935 , n80936 , n80937 , n80938 , n80939 , n80940 , n80941 , n80942 , n80943 , n80944 , 
 n80945 , n80946 , n80947 , n80948 , n80949 , n80950 , n80951 , n80952 , n80953 , n80954 , 
 n80955 , n80956 , n80957 , n80958 , n80959 , n80960 , n80961 , n80962 , n80963 , n80964 , 
 n80965 , n80966 , n80967 , n80968 , n80969 , n80970 , n80971 , n80972 , n80973 , n80974 , 
 n80975 , n80976 , n80977 , n80978 , n80979 , n80980 , n80981 , n80982 , n80983 , n80984 , 
 n80985 , n80986 , n80987 , n80988 , n80989 , n80990 , n80991 , n80992 , n80993 , n80994 , 
 n80995 , n80996 , n80997 , n80998 , n80999 , n81000 , n81001 , n81002 , n81003 , n81004 , 
 n81005 , n81006 , n81007 , n81008 , n81009 , n81010 , n81011 , n81012 , n81013 , n81014 , 
 n81015 , n81016 , n81017 , n81018 , n81019 , n81020 , n81021 , n81022 , n81023 , n81024 , 
 n81025 , n81026 , n81027 , n81028 , n81029 , n81030 , n81031 , n81032 , n81033 , n81034 , 
 n81035 , n81036 , n81037 , n81038 , n81039 , n81040 , n81041 , n81042 , n81043 , n81044 , 
 n81045 , n81046 , n81047 , n81048 , n81049 , n81050 , n81051 , n81052 , n81053 , n81054 , 
 n81055 , n81056 , n81057 , n81058 , n81059 , n81060 , n81061 , n81062 , n81063 , n81064 , 
 n81065 , n81066 , n81067 , n81068 , n81069 , n81070 , n81071 , n81072 , n81073 , n81074 , 
 n81075 , n81076 , n81077 , n81078 , n81079 , n81080 , n81081 , n81082 , n81083 , n81084 , 
 n81085 , n81086 , n81087 , n81088 , n81089 , n81090 , n81091 , n81092 , n81093 , n81094 , 
 n81095 , n81096 , n81097 , n81098 , n81099 , n81100 , n81101 , n81102 , n81103 , n81104 , 
 n81105 , n81106 , n81107 , n81108 , n81109 , n81110 , n81111 , n81112 , n81113 , n81114 , 
 n81115 , n81116 , n81117 , n81118 , n81119 , n81120 , n81121 , n81122 , n81123 , n81124 , 
 n81125 , n81126 , n81127 , n81128 , n81129 , n81130 , n81131 , n81132 , n81133 , n81134 , 
 n81135 , n81136 , n81137 , n81138 , n81139 , n81140 , n81141 , n81142 , n81143 , n81144 , 
 n81145 , n81146 , n81147 , n81148 , n81149 , n81150 , n81151 , n81152 , n81153 , n81154 , 
 n81155 , n81156 , n81157 , n81158 , n81159 , n81160 , n81161 , n81162 , n81163 , n81164 , 
 n81165 , n81166 , n81167 , n81168 , n81169 , n81170 , n81171 , n81172 , n81173 , n81174 , 
 n81175 , n81176 , n81177 , n81178 , n81179 , n81180 , n81181 , n81182 , n81183 , n81184 , 
 n81185 , n81186 , n81187 , n81188 , n81189 , n81190 , n81191 , n81192 , n81193 , n81194 , 
 n81195 , n81196 , n81197 , n81198 , n81199 , n81200 , n81201 , n81202 , n81203 , n81204 , 
 n81205 , n81206 , n81207 , n81208 , n81209 , n81210 , n81211 , n81212 , n81213 , n81214 , 
 n81215 , n81216 , n81217 , n81218 , n81219 , n81220 , n81221 , n81222 , n81223 , n81224 , 
 n81225 , n81226 , n81227 , n81228 , n81229 , n81230 , n81231 , n81232 , n81233 , n81234 , 
 n81235 , n81236 , n81237 , n81238 , n81239 , n81240 , n81241 , n81242 , n81243 , n81244 , 
 n81245 , n81246 , n81247 , n81248 , n81249 , n81250 , n81251 , n81252 , n81253 , n81254 , 
 n81255 , n81256 , n81257 , n81258 , n81259 , n81260 , n81261 , n81262 , n81263 , n81264 , 
 n81265 , n81266 , n81267 , n81268 , n81269 , n81270 , n81271 , n81272 , n81273 , n81274 , 
 n81275 , n81276 , n81277 , n81278 , n81279 , n81280 , n81281 , n81282 , n81283 , n81284 , 
 n81285 , n81286 , n81287 , n81288 , n81289 , n81290 , n81291 , n81292 , n81293 , n81294 , 
 n81295 , n81296 , n81297 , n81298 , n81299 , n81300 , n81301 , n81302 , n81303 , n81304 , 
 n81305 , n81306 , n81307 , n81308 , n81309 , n81310 , n81311 , n81312 , n81313 , n81314 , 
 n81315 , n81316 , n81317 , n81318 , n81319 , n81320 , n81321 , n81322 , n81323 , n81324 , 
 n81325 , n81326 , n81327 , n81328 , n81329 , n81330 , n81331 , n81332 , n81333 , n81334 , 
 n81335 , n81336 , n81337 , n81338 , n81339 , n81340 , n81341 , n81342 , n81343 , n81344 , 
 n81345 , n81346 , n81347 , n81348 , n81349 , n81350 , n81351 , n81352 , n81353 , n81354 , 
 n81355 , n81356 , n81357 , n81358 , n81359 , n81360 , n81361 , n81362 , n81363 , n81364 , 
 n81365 , n81366 , n81367 , n81368 , n81369 , n81370 , n81371 , n81372 , n81373 , n81374 , 
 n81375 , n81376 , n81377 , n81378 , n81379 , n81380 , n81381 , n81382 , n81383 , n81384 , 
 n81385 , n81386 , n81387 , n81388 , n81389 , n81390 , n81391 , n81392 , n81393 , n81394 , 
 n81395 , n81396 , n81397 , n81398 , n81399 , n81400 , n81401 , n81402 , n81403 , n81404 , 
 n81405 , n81406 , n81407 , n81408 , n81409 , n81410 , n81411 , n81412 , n81413 , n81414 , 
 n81415 , n81416 , n81417 , n81418 , n81419 , n81420 , n81421 , n81422 , n81423 , n81424 , 
 n81425 , n81426 , n81427 , n81428 , n81429 , n81430 , n81431 , n81432 , n81433 , n81434 , 
 n81435 , n81436 , n81437 , n81438 , n81439 , n81440 , n81441 , n81442 , n81443 , n81444 , 
 n81445 , n81446 , n81447 , n81448 , n81449 , n81450 , n81451 , n81452 , n81453 , n81454 , 
 n81455 , n81456 , n81457 , n81458 , n81459 , n81460 , n81461 , n81462 , n81463 , n81464 , 
 n81465 , n81466 , n81467 , n81468 , n81469 , n81470 , n81471 , n81472 , n81473 , n81474 , 
 n81475 , n81476 , n81477 , n81478 , n81479 , n81480 , n81481 , n81482 , n81483 , n81484 , 
 n81485 , n81486 , n81487 , n81488 , n81489 , n81490 , n81491 , n81492 , n81493 , n81494 , 
 n81495 , n81496 , n81497 , n81498 , n81499 , n81500 , n81501 , n81502 , n81503 , n81504 , 
 n81505 , n81506 , n81507 , n81508 , n81509 , n81510 , n81511 , n81512 , n81513 , n81514 , 
 n81515 , n81516 , n81517 , n81518 , n81519 , n81520 , n81521 , n81522 , n81523 , n81524 , 
 n81525 , n81526 , n81527 , n81528 , n81529 , n81530 , n81531 , n81532 , n81533 , n81534 , 
 n81535 , n81536 , n81537 , n81538 , n81539 , n81540 , n81541 , n81542 , n81543 , n81544 , 
 n81545 , n81546 , n81547 , n81548 , n81549 , n81550 , n81551 , n81552 , n81553 , n81554 , 
 n81555 , n81556 , n81557 , n81558 , n81559 , n81560 , n81561 , n81562 , n81563 , n81564 , 
 n81565 , n81566 , n81567 , n81568 , n81569 , n81570 , n81571 , n81572 , n81573 , n81574 , 
 n81575 , n81576 , n81577 , n81578 , n81579 , n81580 , n81581 , n81582 , n81583 , n81584 , 
 n81585 , n81586 , n81587 , n81588 , n81589 , n81590 , n81591 , n81592 , n81593 , n81594 , 
 n81595 , n81596 , n81597 , n81598 , n81599 , n81600 , n81601 , n81602 , n81603 , n81604 , 
 n81605 , n81606 , n81607 , n81608 , n81609 , n81610 , n81611 , n81612 , n81613 , n81614 , 
 n81615 , n81616 , n81617 , n81618 , n81619 , n81620 , n81621 , n81622 , n81623 , n81624 , 
 n81625 , n81626 , n81627 , n81628 , n81629 , n81630 , n81631 , n81632 , n81633 , n81634 , 
 n81635 , n81636 , n81637 , n81638 , n81639 , n81640 , n81641 , n81642 , n81643 , n81644 , 
 n81645 , n81646 , n81647 , n81648 , n81649 , n81650 , n81651 , n81652 , n81653 , n81654 , 
 n81655 , n81656 , n81657 , n81658 , n81659 , n81660 , n81661 , n81662 , n81663 , n81664 , 
 n81665 , n81666 , n81667 , n81668 , n81669 , n81670 , n81671 , n81672 , n81673 , n81674 , 
 n81675 , n81676 , n81677 , n81678 , n81679 , n81680 , n81681 , n81682 , n81683 , n81684 , 
 n81685 , n81686 , n81687 , n81688 , n81689 , n81690 , n81691 , n81692 , n81693 , n81694 , 
 n81695 , n81696 , n81697 , n81698 , n81699 , n81700 , n81701 , n81702 , n81703 , n81704 , 
 n81705 , n81706 , n81707 , n81708 , n81709 , n81710 , n81711 , n81712 , n81713 , n81714 , 
 n81715 , n81716 , n81717 , n81718 , n81719 , n81720 , n81721 , n81722 , n81723 , n81724 , 
 n81725 , n81726 , n81727 , n81728 , n81729 , n81730 , n81731 , n81732 , n81733 , n81734 , 
 n81735 , n81736 , n81737 , n81738 , n81739 , n81740 , n81741 , n81742 , n81743 , n81744 , 
 n81745 , n81746 , n81747 , n81748 , n81749 , n81750 , n81751 , n81752 , n81753 , n81754 , 
 n81755 , n81756 , n81757 , n81758 , n81759 , n81760 , n81761 , n81762 , n81763 , n81764 , 
 n81765 , n81766 , n81767 , n81768 , n81769 , n81770 , n81771 , n81772 , n81773 , n81774 , 
 n81775 , n81776 , n81777 , n81778 , n81779 , n81780 , n81781 , n81782 , n81783 , n81784 , 
 n81785 , n81786 , n81787 , n81788 , n81789 , n81790 , n81791 , n81792 , n81793 , n81794 , 
 n81795 , n81796 , n81797 , n81798 , n81799 , n81800 , n81801 , n81802 , n81803 , n81804 , 
 n81805 , n81806 , n81807 , n81808 , n81809 , n81810 , n81811 , n81812 , n81813 , n81814 , 
 n81815 , n81816 , n81817 , n81818 , n81819 , n81820 , n81821 , n81822 , n81823 , n81824 , 
 n81825 , n81826 , n81827 , n81828 , n81829 , n81830 , n81831 , n81832 , n81833 , n81834 , 
 n81835 , n81836 , n81837 , n81838 , n81839 , n81840 , n81841 , n81842 , n81843 , n81844 , 
 n81845 , n81846 , n81847 , n81848 , n81849 , n81850 , n81851 , n81852 , n81853 , n81854 , 
 n81855 , n81856 , n81857 , n81858 , n81859 , n81860 , n81861 , n81862 , n81863 , n81864 , 
 n81865 , n81866 , n81867 , n81868 , n81869 , n81870 , n81871 , n81872 , n81873 , n81874 , 
 n81875 , n81876 , n81877 , n81878 , n81879 , n81880 , n81881 , n81882 , n81883 , n81884 , 
 n81885 , n81886 , n81887 , n81888 , n81889 , n81890 , n81891 , n81892 , n81893 , n81894 , 
 n81895 , n81896 , n81897 , n81898 , n81899 , n81900 , n81901 , n81902 , n81903 , n81904 , 
 n81905 , n81906 , n81907 , n81908 , n81909 , n81910 , n81911 , n81912 , n81913 , n81914 , 
 n81915 , n81916 , n81917 , n81918 , n81919 , n81920 , n81921 , n81922 , n81923 , n81924 , 
 n81925 , n81926 , n81927 , n81928 , n81929 , n81930 , n81931 , n81932 , n81933 , n81934 , 
 n81935 , n81936 , n81937 , n81938 , n81939 , n81940 , n81941 , n81942 , n81943 , n81944 , 
 n81945 , n81946 , n81947 , n81948 , n81949 , n81950 , n81951 , n81952 , n81953 , n81954 , 
 n81955 , n81956 , n81957 , n81958 , n81959 , n81960 , n81961 , n81962 , n81963 , n81964 , 
 n81965 , n81966 , n81967 , n81968 , n81969 , n81970 , n81971 , n81972 , n81973 , n81974 , 
 n81975 , n81976 , n81977 , n81978 , n81979 , n81980 , n81981 , n81982 , n81983 , n81984 , 
 n81985 , n81986 , n81987 , n81988 , n81989 , n81990 , n81991 , n81992 , n81993 , n81994 , 
 n81995 , n81996 , n81997 , n81998 , n81999 , n82000 , n82001 , n82002 , n82003 , n82004 , 
 n82005 , n82006 , n82007 , n82008 , n82009 , n82010 , n82011 , n82012 , n82013 , n82014 , 
 n82015 , n82016 , n82017 , n82018 , n82019 , n82020 , n82021 , n82022 , n82023 , n82024 , 
 n82025 , n82026 , n82027 , n82028 , n82029 , n82030 , n82031 , n82032 , n82033 , n82034 , 
 n82035 , n82036 , n82037 , n82038 , n82039 , n82040 , n82041 , n82042 , n82043 , n82044 , 
 n82045 , n82046 , n82047 , n82048 , n82049 , n82050 , n82051 , n82052 , n82053 , n82054 , 
 n82055 , n82056 , n82057 , n82058 , n82059 , n82060 , n82061 , n82062 , n82063 , n82064 , 
 n82065 , n82066 , n82067 , n82068 , n82069 , n82070 , n82071 , n82072 , n82073 , n82074 , 
 n82075 , n82076 , n82077 , n82078 , n82079 , n82080 , n82081 , n82082 , n82083 , n82084 , 
 n82085 , n82086 , n82087 , n82088 , n82089 , n82090 , n82091 , n82092 , n82093 , n82094 , 
 n82095 , n82096 , n82097 , n82098 , n82099 , n82100 , n82101 , n82102 , n82103 , n82104 , 
 n82105 , n82106 , n82107 , n82108 , n82109 , n82110 , n82111 , n82112 , n82113 , n82114 , 
 n82115 , n82116 , n82117 , n82118 , n82119 , n82120 , n82121 , n82122 , n82123 , n82124 , 
 n82125 , n82126 , n82127 , n82128 , n82129 , n82130 , n82131 , n82132 , n82133 , n82134 , 
 n82135 , n82136 , n82137 , n82138 , n82139 , n82140 , n82141 , n82142 , n82143 , n82144 , 
 n82145 , n82146 , n82147 , n82148 , n82149 , n82150 , n82151 , n82152 , n82153 , n82154 , 
 n82155 , n82156 , n82157 , n82158 , n82159 , n82160 , n82161 , n82162 , n82163 , n82164 , 
 n82165 , n82166 , n82167 , n82168 , n82169 , n82170 , n82171 , n82172 , n82173 , n82174 , 
 n82175 , n82176 , n82177 , n82178 , n82179 , n82180 , n82181 , n82182 , n82183 , n82184 , 
 n82185 , n82186 , n82187 , n82188 , n82189 , n82190 , n82191 , n82192 , n82193 , n82194 , 
 n82195 , n82196 , n82197 , n82198 , n82199 , n82200 , n82201 , n82202 , n82203 , n82204 , 
 n82205 , n82206 , n82207 , n82208 , n82209 , n82210 , n82211 , n82212 , n82213 , n82214 , 
 n82215 , n82216 , n82217 , n82218 , n82219 , n82220 , n82221 , n82222 , n82223 , n82224 , 
 n82225 , n82226 , n82227 , n82228 , n82229 , n82230 , n82231 , n82232 , n82233 , n82234 , 
 n82235 , n82236 , n82237 , n82238 , n82239 , n82240 , n82241 , n82242 , n82243 , n82244 , 
 n82245 , n82246 , n82247 , n82248 , n82249 , n82250 , n82251 , n82252 , n82253 , n82254 , 
 n82255 , n82256 , n82257 , n82258 , n82259 , n82260 , n82261 , n82262 , n82263 , n82264 , 
 n82265 , n82266 , n82267 , n82268 , n82269 , n82270 , n82271 , n82272 , n82273 , n82274 , 
 n82275 , n82276 , n82277 , n82278 , n82279 , n82280 , n82281 , n82282 , n82283 , n82284 , 
 n82285 , n82286 , n82287 , n82288 , n82289 , n82290 , n82291 , n82292 , n82293 , n82294 , 
 n82295 , n82296 , n82297 , n82298 , n82299 , n82300 , n82301 , n82302 , n82303 , n82304 , 
 n82305 , n82306 , n82307 , n82308 , n82309 , n82310 , n82311 , n82312 , n82313 , n82314 , 
 n82315 , n82316 , n82317 , n82318 , n82319 , n82320 , n82321 , n82322 , n82323 , n82324 , 
 n82325 , n82326 , n82327 , n82328 , n82329 , n82330 , n82331 , n82332 , n82333 , n82334 , 
 n82335 , n82336 , n82337 , n82338 , n82339 , n82340 , n82341 , n82342 , n82343 , n82344 , 
 n82345 , n82346 , n82347 , n82348 , n82349 , n82350 , n82351 , n82352 , n82353 , n82354 , 
 n82355 , n82356 , n82357 , n82358 , n82359 , n82360 , n82361 , n82362 , n82363 , n82364 , 
 n82365 , n82366 , n82367 , n82368 , n82369 , n82370 , n82371 , n82372 , n82373 , n82374 , 
 n82375 , n82376 , n82377 , n82378 , n82379 , n82380 , n82381 , n82382 , n82383 , n82384 , 
 n82385 , n82386 , n82387 , n82388 , n82389 , n82390 , n82391 , n82392 , n82393 , n82394 , 
 n82395 , n82396 , n82397 , n82398 , n82399 , n82400 , n82401 , n82402 , n82403 , n82404 , 
 n82405 , n82406 , n82407 , n82408 , n82409 , n82410 , n82411 , n82412 , n82413 , n82414 , 
 n82415 , n82416 , n82417 , n82418 , n82419 , n82420 , n82421 , n82422 , n82423 , n82424 , 
 n82425 , n82426 , n82427 , n82428 , n82429 , n82430 , n82431 , n82432 , n82433 , n82434 , 
 n82435 , n82436 , n82437 , n82438 , n82439 , n82440 , n82441 , n82442 , n82443 , n82444 , 
 n82445 , n82446 , n82447 , n82448 , n82449 , n82450 , n82451 , n82452 , n82453 , n82454 , 
 n82455 , n82456 , n82457 , n82458 , n82459 , n82460 , n82461 , n82462 , n82463 , n82464 , 
 n82465 , n82466 , n82467 , n82468 , n82469 , n82470 , n82471 , n82472 , n82473 , n82474 , 
 n82475 , n82476 , n82477 , n82478 , n82479 , n82480 , n82481 , n82482 , n82483 , n82484 , 
 n82485 , n82486 , n82487 , n82488 , n82489 , n82490 , n82491 , n82492 , n82493 , n82494 , 
 n82495 , n82496 , n82497 , n82498 , n82499 , n82500 , n82501 , n82502 , n82503 , n82504 , 
 n82505 , n82506 , n82507 , n82508 , n82509 , n82510 , n82511 , n82512 , n82513 , n82514 , 
 n82515 , n82516 , n82517 , n82518 , n82519 , n82520 , n82521 , n82522 , n82523 , n82524 , 
 n82525 , n82526 , n82527 , n82528 , n82529 , n82530 , n82531 , n82532 , n82533 , n82534 , 
 n82535 , n82536 , n82537 , n82538 , n82539 , n82540 , n82541 , n82542 , n82543 , n82544 , 
 n82545 , n82546 , n82547 , n82548 , n82549 , n82550 , n82551 , n82552 , n82553 , n82554 , 
 n82555 , n82556 , n82557 , n82558 , n82559 , n82560 , n82561 , n82562 , n82563 , n82564 , 
 n82565 , n82566 , n82567 , n82568 , n82569 , n82570 , n82571 , n82572 , n82573 , n82574 , 
 n82575 , n82576 , n82577 , n82578 , n82579 , n82580 , n82581 , n82582 , n82583 , n82584 , 
 n82585 , n82586 , n82587 , n82588 , n82589 , n82590 , n82591 , n82592 , n82593 , n82594 , 
 n82595 , n82596 , n82597 , n82598 , n82599 , n82600 , n82601 , n82602 , n82603 , n82604 , 
 n82605 , n82606 , n82607 , n82608 , n82609 , n82610 , n82611 , n82612 , n82613 , n82614 , 
 n82615 , n82616 , n82617 , n82618 , n82619 , n82620 , n82621 , n82622 , n82623 , n82624 , 
 n82625 , n82626 , n82627 , n82628 , n82629 , n82630 , n82631 , n82632 , n82633 , n82634 , 
 n82635 , n82636 , n82637 , n82638 , n82639 , n82640 , n82641 , n82642 , n82643 , n82644 , 
 n82645 , n82646 , n82647 , n82648 , n82649 , n82650 , n82651 , n82652 , n82653 , n82654 , 
 n82655 , n82656 , n82657 , n82658 , n82659 , n82660 , n82661 , n82662 , n82663 , n82664 , 
 n82665 , n82666 , n82667 , n82668 , n82669 , n82670 , n82671 , n82672 , n82673 , n82674 , 
 n82675 , n82676 , n82677 , n82678 , n82679 , n82680 , n82681 , n82682 , n82683 , n82684 , 
 n82685 , n82686 , n82687 , n82688 , n82689 , n82690 , n82691 , n82692 , n82693 , n82694 , 
 n82695 , n82696 , n82697 , n82698 , n82699 , n82700 , n82701 , n82702 , n82703 , n82704 , 
 n82705 , n82706 , n82707 , n82708 , n82709 , n82710 , n82711 , n82712 , n82713 , n82714 , 
 n82715 , n82716 , n82717 , n82718 , n82719 , n82720 , n82721 , n82722 , n82723 , n82724 , 
 n82725 , n82726 , n82727 , n82728 , n82729 , n82730 , n82731 , n82732 , n82733 , n82734 , 
 n82735 , n82736 , n82737 , n82738 , n82739 , n82740 , n82741 , n82742 , n82743 , n82744 , 
 n82745 , n82746 , n82747 , n82748 , n82749 , n82750 , n82751 , n82752 , n82753 , n82754 , 
 n82755 , n82756 , n82757 , n82758 , n82759 , n82760 , n82761 , n82762 , n82763 , n82764 , 
 n82765 , n82766 , n82767 , n82768 , n82769 , n82770 , n82771 , n82772 , n82773 , n82774 , 
 n82775 , n82776 , n82777 , n82778 , n82779 , n82780 , n82781 , n82782 , n82783 , n82784 , 
 n82785 , n82786 , n82787 , n82788 , n82789 , n82790 , n82791 , n82792 , n82793 , n82794 , 
 n82795 , n82796 , n82797 , n82798 , n82799 , n82800 , n82801 , n82802 , n82803 , n82804 , 
 n82805 , n82806 , n82807 , n82808 , n82809 , n82810 , n82811 , n82812 , n82813 , n82814 , 
 n82815 , n82816 , n82817 , n82818 , n82819 , n82820 , n82821 , n82822 , n82823 , n82824 , 
 n82825 , n82826 , n82827 , n82828 , n82829 , n82830 , n82831 , n82832 , n82833 , n82834 , 
 n82835 , n82836 , n82837 , n82838 , n82839 , n82840 , n82841 , n82842 , n82843 , n82844 , 
 n82845 , n82846 , n82847 , n82848 , n82849 , n82850 , n82851 , n82852 , n82853 , n82854 , 
 n82855 , n82856 , n82857 , n82858 , n82859 , n82860 , n82861 , n82862 , n82863 , n82864 , 
 n82865 , n82866 , n82867 , n82868 , n82869 , n82870 , n82871 , n82872 , n82873 , n82874 , 
 n82875 , n82876 , n82877 , n82878 , n82879 , n82880 , n82881 , n82882 , n82883 , n82884 , 
 n82885 , n82886 , n82887 , n82888 , n82889 , n82890 , n82891 , n82892 , n82893 , n82894 , 
 n82895 , n82896 , n82897 , n82898 , n82899 , n82900 , n82901 , n82902 , n82903 , n82904 , 
 n82905 , n82906 , n82907 , n82908 , n82909 , n82910 , n82911 , n82912 , n82913 , n82914 , 
 n82915 , n82916 , n82917 , n82918 , n82919 , n82920 , n82921 , n82922 , n82923 , n82924 , 
 n82925 , n82926 , n82927 , n82928 , n82929 , n82930 , n82931 , n82932 , n82933 , n82934 , 
 n82935 , n82936 , n82937 , n82938 , n82939 , n82940 , n82941 , n82942 , n82943 , n82944 , 
 n82945 , n82946 , n82947 , n82948 , n82949 , n82950 , n82951 , n82952 , n82953 , n82954 , 
 n82955 , n82956 , n82957 , n82958 , n82959 , n82960 , n82961 , n82962 , n82963 , n82964 , 
 n82965 , n82966 , n82967 , n82968 , n82969 , n82970 , n82971 , n82972 , n82973 , n82974 , 
 n82975 , n82976 , n82977 , n82978 , n82979 , n82980 , n82981 , n82982 , n82983 , n82984 , 
 n82985 , n82986 , n82987 , n82988 , n82989 , n82990 , n82991 , n82992 , n82993 , n82994 , 
 n82995 , n82996 , n82997 , n82998 , n82999 , n83000 , n83001 , n83002 , n83003 , n83004 , 
 n83005 , n83006 , n83007 , n83008 , n83009 , n83010 , n83011 , n83012 , n83013 , n83014 , 
 n83015 , n83016 , n83017 , n83018 , n83019 , n83020 , n83021 , n83022 , n83023 , n83024 , 
 n83025 , n83026 , n83027 , n83028 , n83029 , n83030 , n83031 , n83032 , n83033 , n83034 , 
 n83035 , n83036 , n83037 , n83038 , n83039 , n83040 , n83041 , n83042 , n83043 , n83044 , 
 n83045 , n83046 , n83047 , n83048 , n83049 , n83050 , n83051 , n83052 , n83053 , n83054 , 
 n83055 , n83056 , n83057 , n83058 , n83059 , n83060 , n83061 , n83062 , n83063 , n83064 , 
 n83065 , n83066 , n83067 , n83068 , n83069 , n83070 , n83071 , n83072 , n83073 , n83074 , 
 n83075 , n83076 , n83077 , n83078 , n83079 , n83080 , n83081 , n83082 , n83083 , n83084 , 
 n83085 , n83086 , n83087 , n83088 , n83089 , n83090 , n83091 , n83092 , n83093 , n83094 , 
 n83095 , n83096 , n83097 , n83098 , n83099 , n83100 , n83101 , n83102 , n83103 , n83104 , 
 n83105 , n83106 , n83107 , n83108 , n83109 , n83110 , n83111 , n83112 , n83113 , n83114 , 
 n83115 , n83116 , n83117 , n83118 , n83119 , n83120 , n83121 , n83122 , n83123 , n83124 , 
 n83125 , n83126 , n83127 , n83128 , n83129 , n83130 , n83131 , n83132 , n83133 , n83134 , 
 n83135 , n83136 , n83137 , n83138 , n83139 , n83140 , n83141 , n83142 , n83143 , n83144 , 
 n83145 , n83146 , n83147 , n83148 , n83149 , n83150 , n83151 , n83152 , n83153 , n83154 , 
 n83155 , n83156 , n83157 , n83158 , n83159 , n83160 , n83161 , n83162 , n83163 , n83164 , 
 n83165 , n83166 , n83167 , n83168 , n83169 , n83170 , n83171 , n83172 , n83173 , n83174 , 
 n83175 , n83176 , n83177 , n83178 , n83179 , n83180 , n83181 , n83182 , n83183 , n83184 , 
 n83185 , n83186 , n83187 , n83188 , n83189 , n83190 , n83191 , n83192 , n83193 , n83194 , 
 n83195 , n83196 , n83197 , n83198 , n83199 , n83200 , n83201 , n83202 , n83203 , n83204 , 
 n83205 , n83206 , n83207 , n83208 , n83209 , n83210 , n83211 , n83212 , n83213 , n83214 , 
 n83215 , n83216 , n83217 , n83218 , n83219 , n83220 , n83221 , n83222 , n83223 , n83224 , 
 n83225 , n83226 , n83227 , n83228 , n83229 , n83230 , n83231 , n83232 , n83233 , n83234 , 
 n83235 , n83236 , n83237 , n83238 , n83239 , n83240 , n83241 , n83242 , n83243 , n83244 , 
 n83245 , n83246 , n83247 , n83248 , n83249 , n83250 , n83251 , n83252 , n83253 , n83254 , 
 n83255 , n83256 , n83257 , n83258 , n83259 , n83260 , n83261 , n83262 , n83263 , n83264 , 
 n83265 , n83266 , n83267 , n83268 , n83269 , n83270 , n83271 , n83272 , n83273 , n83274 , 
 n83275 , n83276 , n83277 , n83278 , n83279 , n83280 , n83281 , n83282 , n83283 , n83284 , 
 n83285 , n83286 , n83287 , n83288 , n83289 , n83290 , n83291 , n83292 , n83293 , n83294 , 
 n83295 , n83296 , n83297 , n83298 , n83299 , n83300 , n83301 , n83302 , n83303 , n83304 , 
 n83305 , n83306 , n83307 , n83308 , n83309 , n83310 , n83311 , n83312 , n83313 , n83314 , 
 n83315 , n83316 , n83317 , n83318 , n83319 , n83320 , n83321 , n83322 , n83323 , n83324 , 
 n83325 , n83326 , n83327 , n83328 , n83329 , n83330 , n83331 , n83332 , n83333 , n83334 , 
 n83335 , n83336 , n83337 , n83338 , n83339 , n83340 , n83341 , n83342 , n83343 , n83344 , 
 n83345 , n83346 , n83347 , n83348 , n83349 , n83350 , n83351 , n83352 , n83353 , n83354 , 
 n83355 , n83356 , n83357 , n83358 , n83359 , n83360 , n83361 , n83362 , n83363 , n83364 , 
 n83365 , n83366 , n83367 , n83368 , n83369 , n83370 , n83371 , n83372 , n83373 , n83374 , 
 n83375 , n83376 , n83377 , n83378 , n83379 , n83380 , n83381 , n83382 , n83383 , n83384 , 
 n83385 , n83386 , n83387 , n83388 , n83389 , n83390 , n83391 , n83392 , n83393 , n83394 , 
 n83395 , n83396 , n83397 , n83398 , n83399 , n83400 , n83401 , n83402 , n83403 , n83404 , 
 n83405 , n83406 , n83407 , n83408 , n83409 , n83410 , n83411 , n83412 , n83413 , n83414 , 
 n83415 , n83416 , n83417 , n83418 , n83419 , n83420 , n83421 , n83422 , n83423 , n83424 , 
 n83425 , n83426 , n83427 , n83428 , n83429 , n83430 , n83431 , n83432 , n83433 , n83434 , 
 n83435 , n83436 , n83437 , n83438 , n83439 , n83440 , n83441 , n83442 , n83443 , n83444 , 
 n83445 , n83446 , n83447 , n83448 , n83449 , n83450 , n83451 , n83452 , n83453 , n83454 , 
 n83455 , n83456 , n83457 , n83458 , n83459 , n83460 , n83461 , n83462 , n83463 , n83464 , 
 n83465 , n83466 , n83467 , n83468 , n83469 , n83470 , n83471 , n83472 , n83473 , n83474 , 
 n83475 , n83476 , n83477 , n83478 , n83479 , n83480 , n83481 , n83482 , n83483 , n83484 , 
 n83485 , n83486 , n83487 , n83488 , n83489 , n83490 , n83491 , n83492 , n83493 , n83494 , 
 n83495 , n83496 , n83497 , n83498 , n83499 , n83500 , n83501 , n83502 , n83503 , n83504 , 
 n83505 , n83506 , n83507 , n83508 , n83509 , n83510 , n83511 , n83512 , n83513 , n83514 , 
 n83515 , n83516 , n83517 , n83518 , n83519 , n83520 , n83521 , n83522 , n83523 , n83524 , 
 n83525 , n83526 , n83527 , n83528 , n83529 , n83530 , n83531 , n83532 , n83533 , n83534 , 
 n83535 , n83536 , n83537 , n83538 , n83539 , n83540 , n83541 , n83542 , n83543 , n83544 , 
 n83545 , n83546 , n83547 , n83548 , n83549 , n83550 , n83551 , n83552 , n83553 , n83554 , 
 n83555 , n83556 , n83557 , n83558 , n83559 , n83560 , n83561 , n83562 , n83563 , n83564 , 
 n83565 , n83566 , n83567 , n83568 , n83569 , n83570 , n83571 , n83572 , n83573 , n83574 , 
 n83575 , n83576 , n83577 , n83578 , n83579 , n83580 , n83581 , n83582 , n83583 , n83584 , 
 n83585 , n83586 , n83587 , n83588 , n83589 , n83590 , n83591 , n83592 , n83593 , n83594 , 
 n83595 , n83596 , n83597 , n83598 , n83599 , n83600 , n83601 , n83602 , n83603 , n83604 , 
 n83605 , n83606 , n83607 , n83608 , n83609 , n83610 , n83611 , n83612 , n83613 , n83614 , 
 n83615 , n83616 , n83617 , n83618 , n83619 , n83620 , n83621 , n83622 , n83623 , n83624 , 
 n83625 , n83626 , n83627 , n83628 , n83629 , n83630 , n83631 , n83632 , n83633 , n83634 , 
 n83635 , n83636 , n83637 , n83638 , n83639 , n83640 , n83641 , n83642 , n83643 , n83644 , 
 n83645 , n83646 , n83647 , n83648 , n83649 , n83650 , n83651 , n83652 , n83653 , n83654 , 
 n83655 , n83656 , n83657 , n83658 , n83659 , n83660 , n83661 , n83662 , n83663 , n83664 , 
 n83665 , n83666 , n83667 , n83668 , n83669 , n83670 , n83671 , n83672 , n83673 , n83674 , 
 n83675 , n83676 , n83677 , n83678 , n83679 , n83680 , n83681 , n83682 , n83683 , n83684 , 
 n83685 , n83686 , n83687 , n83688 , n83689 , n83690 , n83691 , n83692 , n83693 , n83694 , 
 n83695 , n83696 , n83697 , n83698 , n83699 , n83700 , n83701 , n83702 , n83703 , n83704 , 
 n83705 , n83706 , n83707 , n83708 , n83709 , n83710 , n83711 , n83712 , n83713 , n83714 , 
 n83715 , n83716 , n83717 , n83718 , n83719 , n83720 , n83721 , n83722 , n83723 , n83724 , 
 n83725 , n83726 , n83727 , n83728 , n83729 , n83730 , n83731 , n83732 , n83733 , n83734 , 
 n83735 , n83736 , n83737 , n83738 , n83739 , n83740 , n83741 , n83742 , n83743 , n83744 , 
 n83745 , n83746 , n83747 , n83748 , n83749 , n83750 , n83751 , n83752 , n83753 , n83754 , 
 n83755 , n83756 , n83757 , n83758 , n83759 , n83760 , n83761 , n83762 , n83763 , n83764 , 
 n83765 , n83766 , n83767 , n83768 , n83769 , n83770 , n83771 , n83772 , n83773 , n83774 , 
 n83775 , n83776 , n83777 , n83778 , n83779 , n83780 , n83781 , n83782 , n83783 , n83784 , 
 n83785 , n83786 , n83787 , n83788 , n83789 , n83790 , n83791 , n83792 , n83793 , n83794 , 
 n83795 , n83796 , n83797 , n83798 , n83799 , n83800 , n83801 , n83802 , n83803 , n83804 , 
 n83805 , n83806 , n83807 , n83808 , n83809 , n83810 , n83811 , n83812 , n83813 , n83814 , 
 n83815 , n83816 , n83817 , n83818 , n83819 , n83820 , n83821 , n83822 , n83823 , n83824 , 
 n83825 , n83826 , n83827 , n83828 , n83829 , n83830 , n83831 , n83832 , n83833 , n83834 , 
 n83835 , n83836 , n83837 , n83838 , n83839 , n83840 , n83841 , n83842 , n83843 , n83844 , 
 n83845 , n83846 , n83847 , n83848 , n83849 , n83850 , n83851 , n83852 , n83853 , n83854 , 
 n83855 , n83856 , n83857 , n83858 , n83859 , n83860 , n83861 , n83862 , n83863 , n83864 , 
 n83865 , n83866 , n83867 , n83868 , n83869 , n83870 , n83871 , n83872 , n83873 , n83874 , 
 n83875 , n83876 , n83877 , n83878 , n83879 , n83880 , n83881 , n83882 , n83883 , n83884 , 
 n83885 , n83886 , n83887 , n83888 , n83889 , n83890 , n83891 , n83892 , n83893 , n83894 , 
 n83895 , n83896 , n83897 , n83898 , n83899 , n83900 , n83901 , n83902 , n83903 , n83904 , 
 n83905 , n83906 , n83907 , n83908 , n83909 , n83910 , n83911 , n83912 , n83913 , n83914 , 
 n83915 , n83916 , n83917 , n83918 , n83919 , n83920 , n83921 , n83922 , n83923 , n83924 , 
 n83925 , n83926 , n83927 , n83928 , n83929 , n83930 , n83931 , n83932 , n83933 , n83934 , 
 n83935 , n83936 , n83937 , n83938 , n83939 , n83940 , n83941 , n83942 , n83943 , n83944 , 
 n83945 , n83946 , n83947 , n83948 , n83949 , n83950 , n83951 , n83952 , n83953 , n83954 , 
 n83955 , n83956 , n83957 , n83958 , n83959 , n83960 , n83961 , n83962 , n83963 , n83964 , 
 n83965 , n83966 , n83967 , n83968 , n83969 , n83970 , n83971 , n83972 , n83973 , n83974 , 
 n83975 , n83976 , n83977 , n83978 , n83979 , n83980 , n83981 , n83982 , n83983 , n83984 , 
 n83985 , n83986 , n83987 , n83988 , n83989 , n83990 , n83991 , n83992 , n83993 , n83994 , 
 n83995 , n83996 , n83997 , n83998 , n83999 , n84000 , n84001 , n84002 , n84003 , n84004 , 
 n84005 , n84006 , n84007 , n84008 , n84009 , n84010 , n84011 , n84012 , n84013 , n84014 , 
 n84015 , n84016 , n84017 , n84018 , n84019 , n84020 , n84021 , n84022 , n84023 , n84024 , 
 n84025 , n84026 , n84027 , n84028 , n84029 , n84030 , n84031 , n84032 , n84033 , n84034 , 
 n84035 , n84036 , n84037 , n84038 , n84039 , n84040 , n84041 , n84042 , n84043 , n84044 , 
 n84045 , n84046 , n84047 , n84048 , n84049 , n84050 , n84051 , n84052 , n84053 , n84054 , 
 n84055 , n84056 , n84057 , n84058 , n84059 , n84060 , n84061 , n84062 , n84063 , n84064 , 
 n84065 , n84066 , n84067 , n84068 , n84069 , n84070 , n84071 , n84072 , n84073 , n84074 , 
 n84075 , n84076 , n84077 , n84078 , n84079 , n84080 , n84081 , n84082 , n84083 , n84084 , 
 n84085 , n84086 , n84087 , n84088 , n84089 , n84090 , n84091 , n84092 , n84093 , n84094 , 
 n84095 , n84096 , n84097 , n84098 , n84099 , n84100 , n84101 , n84102 , n84103 , n84104 , 
 n84105 , n84106 , n84107 , n84108 , n84109 , n84110 , n84111 , n84112 , n84113 , n84114 , 
 n84115 , n84116 , n84117 , n84118 , n84119 , n84120 , n84121 , n84122 , n84123 , n84124 , 
 n84125 , n84126 , n84127 , n84128 , n84129 , n84130 , n84131 , n84132 , n84133 , n84134 , 
 n84135 , n84136 , n84137 , n84138 , n84139 , n84140 , n84141 , n84142 , n84143 , n84144 , 
 n84145 , n84146 , n84147 , n84148 , n84149 , n84150 , n84151 , n84152 , n84153 , n84154 , 
 n84155 , n84156 , n84157 , n84158 , n84159 , n84160 , n84161 , n84162 , n84163 , n84164 , 
 n84165 , n84166 , n84167 , n84168 , n84169 , n84170 , n84171 , n84172 , n84173 , n84174 , 
 n84175 , n84176 , n84177 , n84178 , n84179 , n84180 , n84181 , n84182 , n84183 , n84184 , 
 n84185 , n84186 , n84187 , n84188 , n84189 , n84190 , n84191 , n84192 , n84193 , n84194 , 
 n84195 , n84196 , n84197 , n84198 , n84199 , n84200 , n84201 , n84202 , n84203 , n84204 , 
 n84205 , n84206 , n84207 , n84208 , n84209 , n84210 , n84211 , n84212 , n84213 , n84214 , 
 n84215 , n84216 , n84217 , n84218 , n84219 , n84220 , n84221 , n84222 , n84223 , n84224 , 
 n84225 , n84226 , n84227 , n84228 , n84229 , n84230 , n84231 , n84232 , n84233 , n84234 , 
 n84235 , n84236 , n84237 , n84238 , n84239 , n84240 , n84241 , n84242 , n84243 , n84244 , 
 n84245 , n84246 , n84247 , n84248 , n84249 , n84250 , n84251 , n84252 , n84253 , n84254 , 
 n84255 , n84256 , n84257 , n84258 , n84259 , n84260 , n84261 , n84262 , n84263 , n84264 , 
 n84265 , n84266 , n84267 , n84268 , n84269 , n84270 , n84271 , n84272 , n84273 , n84274 , 
 n84275 , n84276 , n84277 , n84278 , n84279 , n84280 , n84281 , n84282 , n84283 , n84284 , 
 n84285 , n84286 , n84287 , n84288 , n84289 , n84290 , n84291 , n84292 , n84293 , n84294 , 
 n84295 , n84296 , n84297 , n84298 , n84299 , n84300 , n84301 , n84302 , n84303 , n84304 , 
 n84305 , n84306 , n84307 , n84308 , n84309 , n84310 , n84311 , n84312 , n84313 , n84314 , 
 n84315 , n84316 , n84317 , n84318 , n84319 , n84320 , n84321 , n84322 , n84323 , n84324 , 
 n84325 , n84326 , n84327 , n84328 , n84329 , n84330 , n84331 , n84332 , n84333 , n84334 , 
 n84335 , n84336 , n84337 , n84338 , n84339 , n84340 , n84341 , n84342 , n84343 , n84344 , 
 n84345 , n84346 , n84347 , n84348 , n84349 , n84350 , n84351 , n84352 , n84353 , n84354 , 
 n84355 , n84356 , n84357 , n84358 , n84359 , n84360 , n84361 , n84362 , n84363 , n84364 , 
 n84365 , n84366 , n84367 , n84368 , n84369 , n84370 , n84371 , n84372 , n84373 , n84374 , 
 n84375 , n84376 , n84377 , n84378 , n84379 , n84380 , n84381 , n84382 , n84383 , n84384 , 
 n84385 , n84386 , n84387 , n84388 , n84389 , n84390 , n84391 , n84392 , n84393 , n84394 , 
 n84395 , n84396 , n84397 , n84398 , n84399 , n84400 , n84401 , n84402 , n84403 , n84404 , 
 n84405 , n84406 , n84407 , n84408 , n84409 , n84410 , n84411 , n84412 , n84413 , n84414 , 
 n84415 , n84416 , n84417 , n84418 , n84419 , n84420 , n84421 , n84422 , n84423 , n84424 , 
 n84425 , n84426 , n84427 , n84428 , n84429 , n84430 , n84431 , n84432 , n84433 , n84434 , 
 n84435 , n84436 , n84437 , n84438 , n84439 , n84440 , n84441 , n84442 , n84443 , n84444 , 
 n84445 , n84446 , n84447 , n84448 , n84449 , n84450 , n84451 , n84452 , n84453 , n84454 , 
 n84455 , n84456 , n84457 , n84458 , n84459 , n84460 , n84461 , n84462 , n84463 , n84464 , 
 n84465 , n84466 , n84467 , n84468 , n84469 , n84470 , n84471 , n84472 , n84473 , n84474 , 
 n84475 , n84476 , n84477 , n84478 , n84479 , n84480 , n84481 , n84482 , n84483 , n84484 , 
 n84485 , n84486 , n84487 , n84488 , n84489 , n84490 , n84491 , n84492 , n84493 , n84494 , 
 n84495 , n84496 , n84497 , n84498 , n84499 , n84500 , n84501 , n84502 , n84503 , n84504 , 
 n84505 , n84506 , n84507 , n84508 , n84509 , n84510 , n84511 , n84512 , n84513 , n84514 , 
 n84515 , n84516 , n84517 , n84518 , n84519 , n84520 , n84521 , n84522 , n84523 , n84524 , 
 n84525 , n84526 , n84527 , n84528 , n84529 , n84530 , n84531 , n84532 , n84533 , n84534 , 
 n84535 , n84536 , n84537 , n84538 , n84539 , n84540 , n84541 , n84542 , n84543 , n84544 , 
 n84545 , n84546 , n84547 , n84548 , n84549 , n84550 , n84551 , n84552 , n84553 , n84554 , 
 n84555 , n84556 , n84557 , n84558 , n84559 , n84560 , n84561 , n84562 , n84563 , n84564 , 
 n84565 , n84566 , n84567 , n84568 , n84569 , n84570 , n84571 , n84572 , n84573 , n84574 , 
 n84575 , n84576 , n84577 , n84578 , n84579 , n84580 , n84581 , n84582 , n84583 , n84584 , 
 n84585 , n84586 , n84587 , n84588 , n84589 , n84590 , n84591 , n84592 , n84593 , n84594 , 
 n84595 , n84596 , n84597 , n84598 , n84599 , n84600 , n84601 , n84602 , n84603 , n84604 , 
 n84605 , n84606 , n84607 , n84608 , n84609 , n84610 , n84611 , n84612 , n84613 , n84614 , 
 n84615 , n84616 , n84617 , n84618 , n84619 , n84620 , n84621 , n84622 , n84623 , n84624 , 
 n84625 , n84626 , n84627 , n84628 , n84629 , n84630 , n84631 , n84632 , n84633 , n84634 , 
 n84635 , n84636 , n84637 , n84638 , n84639 , n84640 , n84641 , n84642 , n84643 , n84644 , 
 n84645 , n84646 , n84647 , n84648 , n84649 , n84650 , n84651 , n84652 , n84653 , n84654 , 
 n84655 , n84656 , n84657 , n84658 , n84659 , n84660 , n84661 , n84662 , n84663 , n84664 , 
 n84665 , n84666 , n84667 , n84668 , n84669 , n84670 , n84671 , n84672 , n84673 , n84674 , 
 n84675 , n84676 , n84677 , n84678 , n84679 , n84680 , n84681 , n84682 , n84683 , n84684 , 
 n84685 , n84686 , n84687 , n84688 , n84689 , n84690 , n84691 , n84692 , n84693 , n84694 , 
 n84695 , n84696 , n84697 , n84698 , n84699 , n84700 , n84701 , n84702 , n84703 , n84704 , 
 n84705 , n84706 , n84707 , n84708 , n84709 , n84710 , n84711 , n84712 , n84713 , n84714 , 
 n84715 , n84716 , n84717 , n84718 , n84719 , n84720 , n84721 , n84722 , n84723 , n84724 , 
 n84725 , n84726 , n84727 , n84728 , n84729 , n84730 , n84731 , n84732 , n84733 , n84734 , 
 n84735 , n84736 , n84737 , n84738 , n84739 , n84740 , n84741 , n84742 , n84743 , n84744 , 
 n84745 , n84746 , n84747 , n84748 , n84749 , n84750 , n84751 , n84752 , n84753 , n84754 , 
 n84755 , n84756 , n84757 , n84758 , n84759 , n84760 , n84761 , n84762 , n84763 , n84764 , 
 n84765 , n84766 , n84767 , n84768 , n84769 , n84770 , n84771 , n84772 , n84773 , n84774 , 
 n84775 , n84776 , n84777 , n84778 , n84779 , n84780 , n84781 , n84782 , n84783 , n84784 , 
 n84785 , n84786 , n84787 , n84788 , n84789 , n84790 , n84791 , n84792 , n84793 , n84794 , 
 n84795 , n84796 , n84797 , n84798 , n84799 , n84800 , n84801 , n84802 , n84803 , n84804 , 
 n84805 , n84806 , n84807 , n84808 , n84809 , n84810 , n84811 , n84812 , n84813 , n84814 , 
 n84815 , n84816 , n84817 , n84818 , n84819 , n84820 , n84821 , n84822 , n84823 , n84824 , 
 n84825 , n84826 , n84827 , n84828 , n84829 , n84830 , n84831 , n84832 , n84833 , n84834 , 
 n84835 , n84836 , n84837 , n84838 , n84839 , n84840 , n84841 , n84842 , n84843 , n84844 , 
 n84845 , n84846 , n84847 , n84848 , n84849 , n84850 , n84851 , n84852 , n84853 , n84854 , 
 n84855 , n84856 , n84857 , n84858 , n84859 , n84860 , n84861 , n84862 , n84863 , n84864 , 
 n84865 , n84866 , n84867 , n84868 , n84869 , n84870 , n84871 , n84872 , n84873 , n84874 , 
 n84875 , n84876 , n84877 , n84878 , n84879 , n84880 , n84881 , n84882 , n84883 , n84884 , 
 n84885 , n84886 , n84887 , n84888 , n84889 , n84890 , n84891 , n84892 , n84893 , n84894 , 
 n84895 , n84896 , n84897 , n84898 , n84899 , n84900 , n84901 , n84902 , n84903 , n84904 , 
 n84905 , n84906 , n84907 , n84908 , n84909 , n84910 , n84911 , n84912 , n84913 , n84914 , 
 n84915 , n84916 , n84917 , n84918 , n84919 , n84920 , n84921 , n84922 , n84923 , n84924 , 
 n84925 , n84926 , n84927 , n84928 , n84929 , n84930 , n84931 , n84932 , n84933 , n84934 , 
 n84935 , n84936 , n84937 , n84938 , n84939 , n84940 , n84941 , n84942 , n84943 , n84944 , 
 n84945 , n84946 , n84947 , n84948 , n84949 , n84950 , n84951 , n84952 , n84953 , n84954 , 
 n84955 , n84956 , n84957 , n84958 , n84959 , n84960 , n84961 , n84962 , n84963 , n84964 , 
 n84965 , n84966 , n84967 , n84968 , n84969 , n84970 , n84971 , n84972 , n84973 , n84974 , 
 n84975 , n84976 , n84977 , n84978 , n84979 , n84980 , n84981 , n84982 , n84983 , n84984 , 
 n84985 , n84986 , n84987 , n84988 , n84989 , n84990 , n84991 , n84992 , n84993 , n84994 , 
 n84995 , n84996 , n84997 , n84998 , n84999 , n85000 , n85001 , n85002 , n85003 , n85004 , 
 n85005 , n85006 , n85007 , n85008 , n85009 , n85010 , n85011 , n85012 , n85013 , n85014 , 
 n85015 , n85016 , n85017 , n85018 , n85019 , n85020 , n85021 , n85022 , n85023 , n85024 , 
 n85025 , n85026 , n85027 , n85028 , n85029 , n85030 , n85031 , n85032 , n85033 , n85034 , 
 n85035 , n85036 , n85037 , n85038 , n85039 , n85040 , n85041 , n85042 , n85043 , n85044 , 
 n85045 , n85046 , n85047 , n85048 , n85049 , n85050 , n85051 , n85052 , n85053 , n85054 , 
 n85055 , n85056 , n85057 , n85058 , n85059 , n85060 , n85061 , n85062 , n85063 , n85064 , 
 n85065 , n85066 , n85067 , n85068 , n85069 , n85070 , n85071 , n85072 , n85073 , n85074 , 
 n85075 , n85076 , n85077 , n85078 , n85079 , n85080 , n85081 , n85082 , n85083 , n85084 , 
 n85085 , n85086 , n85087 , n85088 , n85089 , n85090 , n85091 , n85092 , n85093 , n85094 , 
 n85095 , n85096 , n85097 , n85098 , n85099 , n85100 , n85101 , n85102 , n85103 , n85104 , 
 n85105 , n85106 , n85107 , n85108 , n85109 , n85110 , n85111 , n85112 , n85113 , n85114 , 
 n85115 , n85116 , n85117 , n85118 , n85119 , n85120 , n85121 , n85122 , n85123 , n85124 , 
 n85125 , n85126 , n85127 , n85128 , n85129 , n85130 , n85131 , n85132 , n85133 , n85134 , 
 n85135 , n85136 , n85137 , n85138 , n85139 , n85140 , n85141 , n85142 , n85143 , n85144 , 
 n85145 , n85146 , n85147 , n85148 , n85149 , n85150 , n85151 , n85152 , n85153 , n85154 , 
 n85155 , n85156 , n85157 , n85158 , n85159 , n85160 , n85161 , n85162 , n85163 , n85164 , 
 n85165 , n85166 , n85167 , n85168 , n85169 , n85170 , n85171 , n85172 , n85173 , n85174 , 
 n85175 , n85176 , n85177 , n85178 , n85179 , n85180 , n85181 , n85182 , n85183 , n85184 , 
 n85185 , n85186 , n85187 , n85188 , n85189 , n85190 , n85191 , n85192 , n85193 , n85194 , 
 n85195 , n85196 , n85197 , n85198 , n85199 , n85200 , n85201 , n85202 , n85203 , n85204 , 
 n85205 , n85206 , n85207 , n85208 , n85209 , n85210 , n85211 , n85212 , n85213 , n85214 , 
 n85215 , n85216 , n85217 , n85218 , n85219 , n85220 , n85221 , n85222 , n85223 , n85224 , 
 n85225 , n85226 , n85227 , n85228 , n85229 , n85230 , n85231 , n85232 , n85233 , n85234 , 
 n85235 , n85236 , n85237 , n85238 , n85239 , n85240 , n85241 , n85242 , n85243 , n85244 , 
 n85245 , n85246 , n85247 , n85248 , n85249 , n85250 , n85251 , n85252 , n85253 , n85254 , 
 n85255 , n85256 , n85257 , n85258 , n85259 , n85260 , n85261 , n85262 , n85263 , n85264 , 
 n85265 , n85266 , n85267 , n85268 , n85269 , n85270 , n85271 , n85272 , n85273 , n85274 , 
 n85275 , n85276 , n85277 , n85278 , n85279 , n85280 , n85281 , n85282 , n85283 , n85284 , 
 n85285 , n85286 , n85287 , n85288 , n85289 , n85290 , n85291 , n85292 , n85293 , n85294 , 
 n85295 , n85296 , n85297 , n85298 , n85299 , n85300 , n85301 , n85302 , n85303 , n85304 , 
 n85305 , n85306 , n85307 , n85308 , n85309 , n85310 , n85311 , n85312 , n85313 , n85314 , 
 n85315 , n85316 , n85317 , n85318 , n85319 , n85320 , n85321 , n85322 , n85323 , n85324 , 
 n85325 , n85326 , n85327 , n85328 , n85329 , n85330 , n85331 , n85332 , n85333 , n85334 , 
 n85335 , n85336 , n85337 , n85338 , n85339 , n85340 , n85341 , n85342 , n85343 , n85344 , 
 n85345 , n85346 , n85347 , n85348 , n85349 , n85350 , n85351 , n85352 , n85353 , n85354 , 
 n85355 , n85356 , n85357 , n85358 , n85359 , n85360 , n85361 , n85362 , n85363 , n85364 , 
 n85365 , n85366 , n85367 , n85368 , n85369 , n85370 , n85371 , n85372 , n85373 , n85374 , 
 n85375 , n85376 , n85377 , n85378 , n85379 , n85380 , n85381 , n85382 , n85383 , n85384 , 
 n85385 , n85386 , n85387 , n85388 , n85389 , n85390 , n85391 , n85392 , n85393 , n85394 , 
 n85395 , n85396 , n85397 , n85398 , n85399 , n85400 , n85401 , n85402 , n85403 , n85404 , 
 n85405 , n85406 , n85407 , n85408 , n85409 , n85410 , n85411 , n85412 , n85413 , n85414 , 
 n85415 , n85416 , n85417 , n85418 , n85419 , n85420 , n85421 , n85422 , n85423 , n85424 , 
 n85425 , n85426 , n85427 , n85428 , n85429 , n85430 , n85431 , n85432 , n85433 , n85434 , 
 n85435 , n85436 , n85437 , n85438 , n85439 , n85440 , n85441 , n85442 , n85443 , n85444 , 
 n85445 , n85446 , n85447 , n85448 , n85449 , n85450 , n85451 , n85452 , n85453 , n85454 , 
 n85455 , n85456 , n85457 , n85458 , n85459 , n85460 , n85461 , n85462 , n85463 , n85464 , 
 n85465 , n85466 , n85467 , n85468 , n85469 , n85470 , n85471 , n85472 , n85473 , n85474 , 
 n85475 , n85476 , n85477 , n85478 , n85479 , n85480 , n85481 , n85482 , n85483 , n85484 , 
 n85485 , n85486 , n85487 , n85488 , n85489 , n85490 , n85491 , n85492 , n85493 , n85494 , 
 n85495 , n85496 , n85497 , n85498 , n85499 , n85500 , n85501 , n85502 , n85503 , n85504 , 
 n85505 , n85506 , n85507 , n85508 , n85509 , n85510 , n85511 , n85512 , n85513 , n85514 , 
 n85515 , n85516 , n85517 , n85518 , n85519 , n85520 , n85521 , n85522 , n85523 , n85524 , 
 n85525 , n85526 , n85527 , n85528 , n85529 , n85530 , n85531 , n85532 , n85533 , n85534 , 
 n85535 , n85536 , n85537 , n85538 , n85539 , n85540 , n85541 , n85542 , n85543 , n85544 , 
 n85545 , n85546 , n85547 , n85548 , n85549 , n85550 , n85551 , n85552 , n85553 , n85554 , 
 n85555 , n85556 , n85557 , n85558 , n85559 , n85560 , n85561 , n85562 , n85563 , n85564 , 
 n85565 , n85566 , n85567 , n85568 , n85569 , n85570 , n85571 , n85572 , n85573 , n85574 , 
 n85575 , n85576 , n85577 , n85578 , n85579 , n85580 , n85581 , n85582 , n85583 , n85584 , 
 n85585 , n85586 , n85587 , n85588 , n85589 , n85590 , n85591 , n85592 , n85593 , n85594 , 
 n85595 , n85596 , n85597 , n85598 , n85599 , n85600 , n85601 , n85602 , n85603 , n85604 , 
 n85605 , n85606 , n85607 , n85608 , n85609 , n85610 , n85611 , n85612 , n85613 , n85614 , 
 n85615 , n85616 , n85617 , n85618 , n85619 , n85620 , n85621 , n85622 , n85623 , n85624 , 
 n85625 , n85626 , n85627 , n85628 , n85629 , n85630 , n85631 , n85632 , n85633 , n85634 , 
 n85635 , n85636 , n85637 , n85638 , n85639 , n85640 , n85641 , n85642 , n85643 , n85644 , 
 n85645 , n85646 , n85647 , n85648 , n85649 , n85650 , n85651 , n85652 , n85653 , n85654 , 
 n85655 , n85656 , n85657 , n85658 , n85659 , n85660 , n85661 , n85662 , n85663 , n85664 , 
 n85665 , n85666 , n85667 , n85668 , n85669 , n85670 , n85671 , n85672 , n85673 , n85674 , 
 n85675 , n85676 , n85677 , n85678 , n85679 , n85680 , n85681 , n85682 , n85683 , n85684 , 
 n85685 , n85686 , n85687 , n85688 , n85689 , n85690 , n85691 , n85692 , n85693 , n85694 , 
 n85695 , n85696 , n85697 , n85698 , n85699 , n85700 , n85701 , n85702 , n85703 , n85704 , 
 n85705 , n85706 , n85707 , n85708 , n85709 , n85710 , n85711 , n85712 , n85713 , n85714 , 
 n85715 , n85716 , n85717 , n85718 , n85719 , n85720 , n85721 , n85722 , n85723 , n85724 , 
 n85725 , n85726 , n85727 , n85728 , n85729 , n85730 , n85731 , n85732 , n85733 , n85734 , 
 n85735 , n85736 , n85737 , n85738 , n85739 , n85740 , n85741 , n85742 , n85743 , n85744 , 
 n85745 , n85746 , n85747 , n85748 , n85749 , n85750 , n85751 , n85752 , n85753 , n85754 , 
 n85755 , n85756 , n85757 , n85758 , n85759 , n85760 , n85761 , n85762 , n85763 , n85764 , 
 n85765 , n85766 , n85767 , n85768 , n85769 , n85770 , n85771 , n85772 , n85773 , n85774 , 
 n85775 , n85776 , n85777 , n85778 , n85779 , n85780 , n85781 , n85782 , n85783 , n85784 , 
 n85785 , n85786 , n85787 , n85788 , n85789 , n85790 , n85791 , n85792 , n85793 , n85794 , 
 n85795 , n85796 , n85797 , n85798 , n85799 , n85800 , n85801 , n85802 , n85803 , n85804 , 
 n85805 , n85806 , n85807 , n85808 , n85809 , n85810 , n85811 , n85812 , n85813 , n85814 , 
 n85815 , n85816 , n85817 , n85818 , n85819 , n85820 , n85821 , n85822 , n85823 , n85824 , 
 n85825 , n85826 , n85827 , n85828 , n85829 , n85830 , n85831 , n85832 , n85833 , n85834 , 
 n85835 , n85836 , n85837 , n85838 , n85839 , n85840 , n85841 , n85842 , n85843 , n85844 , 
 n85845 , n85846 , n85847 , n85848 , n85849 , n85850 , n85851 , n85852 , n85853 , n85854 , 
 n85855 , n85856 , n85857 , n85858 , n85859 , n85860 , n85861 , n85862 , n85863 , n85864 , 
 n85865 , n85866 , n85867 , n85868 , n85869 , n85870 , n85871 , n85872 , n85873 , n85874 , 
 n85875 , n85876 , n85877 , n85878 , n85879 , n85880 , n85881 , n85882 , n85883 , n85884 , 
 n85885 , n85886 , n85887 , n85888 , n85889 , n85890 , n85891 , n85892 , n85893 , n85894 , 
 n85895 , n85896 , n85897 , n85898 , n85899 , n85900 , n85901 , n85902 , n85903 , n85904 , 
 n85905 , n85906 , n85907 , n85908 , n85909 , n85910 , n85911 , n85912 , n85913 , n85914 , 
 n85915 , n85916 , n85917 , n85918 , n85919 , n85920 , n85921 , n85922 , n85923 , n85924 , 
 n85925 , n85926 , n85927 , n85928 , n85929 , n85930 , n85931 , n85932 , n85933 , n85934 , 
 n85935 , n85936 , n85937 , n85938 , n85939 , n85940 , n85941 , n85942 , n85943 , n85944 , 
 n85945 , n85946 , n85947 , n85948 , n85949 , n85950 , n85951 , n85952 , n85953 , n85954 , 
 n85955 , n85956 , n85957 , n85958 , n85959 , n85960 , n85961 , n85962 , n85963 , n85964 , 
 n85965 , n85966 , n85967 , n85968 , n85969 , n85970 , n85971 , n85972 , n85973 , n85974 , 
 n85975 , n85976 , n85977 , n85978 , n85979 , n85980 , n85981 , n85982 , n85983 , n85984 , 
 n85985 , n85986 , n85987 , n85988 , n85989 , n85990 , n85991 , n85992 , n85993 , n85994 , 
 n85995 , n85996 , n85997 , n85998 , n85999 , n86000 , n86001 , n86002 , n86003 , n86004 , 
 n86005 , n86006 , n86007 , n86008 , n86009 , n86010 , n86011 , n86012 , n86013 , n86014 , 
 n86015 , n86016 , n86017 , n86018 , n86019 , n86020 , n86021 , n86022 , n86023 , n86024 , 
 n86025 , n86026 , n86027 , n86028 , n86029 , n86030 , n86031 , n86032 , n86033 , n86034 , 
 n86035 , n86036 , n86037 , n86038 , n86039 , n86040 , n86041 , n86042 , n86043 , n86044 , 
 n86045 , n86046 , n86047 , n86048 , n86049 , n86050 , n86051 , n86052 , n86053 , n86054 , 
 n86055 , n86056 , n86057 , n86058 , n86059 , n86060 , n86061 , n86062 , n86063 , n86064 , 
 n86065 , n86066 , n86067 , n86068 , n86069 , n86070 , n86071 , n86072 , n86073 , n86074 , 
 n86075 , n86076 , n86077 , n86078 , n86079 , n86080 , n86081 , n86082 , n86083 , n86084 , 
 n86085 , n86086 , n86087 , n86088 , n86089 , n86090 , n86091 , n86092 , n86093 , n86094 , 
 n86095 , n86096 , n86097 , n86098 , n86099 , n86100 , n86101 , n86102 , n86103 , n86104 , 
 n86105 , n86106 , n86107 , n86108 , n86109 , n86110 , n86111 , n86112 , n86113 , n86114 , 
 n86115 , n86116 , n86117 , n86118 , n86119 , n86120 , n86121 , n86122 , n86123 , n86124 , 
 n86125 , n86126 , n86127 , n86128 , n86129 , n86130 , n86131 , n86132 , n86133 , n86134 , 
 n86135 , n86136 , n86137 , n86138 , n86139 , n86140 , n86141 , n86142 , n86143 , n86144 , 
 n86145 , n86146 , n86147 , n86148 , n86149 , n86150 , n86151 , n86152 , n86153 , n86154 , 
 n86155 , n86156 , n86157 , n86158 , n86159 , n86160 , n86161 , n86162 , n86163 , n86164 , 
 n86165 , n86166 , n86167 , n86168 , n86169 , n86170 , n86171 , n86172 , n86173 , n86174 , 
 n86175 , n86176 , n86177 , n86178 , n86179 , n86180 , n86181 , n86182 , n86183 , n86184 , 
 n86185 , n86186 , n86187 , n86188 , n86189 , n86190 , n86191 , n86192 , n86193 , n86194 , 
 n86195 , n86196 , n86197 , n86198 , n86199 , n86200 , n86201 , n86202 , n86203 , n86204 , 
 n86205 , n86206 , n86207 , n86208 , n86209 , n86210 , n86211 , n86212 , n86213 , n86214 , 
 n86215 , n86216 , n86217 , n86218 , n86219 , n86220 , n86221 , n86222 , n86223 , n86224 , 
 n86225 , n86226 , n86227 , n86228 , n86229 , n86230 , n86231 , n86232 , n86233 , n86234 , 
 n86235 , n86236 , n86237 , n86238 , n86239 , n86240 , n86241 , n86242 , n86243 , n86244 , 
 n86245 , n86246 , n86247 , n86248 , n86249 , n86250 , n86251 , n86252 , n86253 , n86254 , 
 n86255 , n86256 , n86257 , n86258 , n86259 , n86260 , n86261 , n86262 , n86263 , n86264 , 
 n86265 , n86266 , n86267 , n86268 , n86269 , n86270 , n86271 , n86272 , n86273 , n86274 , 
 n86275 , n86276 , n86277 , n86278 , n86279 , n86280 , n86281 , n86282 , n86283 , n86284 , 
 n86285 , n86286 , n86287 , n86288 , n86289 , n86290 , n86291 , n86292 , n86293 , n86294 , 
 n86295 , n86296 , n86297 , n86298 , n86299 , n86300 , n86301 , n86302 , n86303 , n86304 , 
 n86305 , n86306 , n86307 , n86308 , n86309 , n86310 , n86311 , n86312 , n86313 , n86314 , 
 n86315 , n86316 , n86317 , n86318 , n86319 , n86320 , n86321 , n86322 , n86323 , n86324 , 
 n86325 , n86326 , n86327 , n86328 , n86329 , n86330 , n86331 , n86332 , n86333 , n86334 , 
 n86335 , n86336 , n86337 , n86338 , n86339 , n86340 , n86341 , n86342 , n86343 , n86344 , 
 n86345 , n86346 , n86347 , n86348 , n86349 , n86350 , n86351 , n86352 , n86353 , n86354 , 
 n86355 , n86356 , n86357 , n86358 , n86359 , n86360 , n86361 , n86362 , n86363 , n86364 , 
 n86365 , n86366 , n86367 , n86368 , n86369 , n86370 , n86371 , n86372 , n86373 , n86374 , 
 n86375 , n86376 , n86377 , n86378 , n86379 , n86380 , n86381 , n86382 , n86383 , n86384 , 
 n86385 , n86386 , n86387 , n86388 , n86389 , n86390 , n86391 , n86392 , n86393 , n86394 , 
 n86395 , n86396 , n86397 , n86398 , n86399 , n86400 , n86401 , n86402 , n86403 , n86404 , 
 n86405 , n86406 , n86407 , n86408 , n86409 , n86410 , n86411 , n86412 , n86413 , n86414 , 
 n86415 , n86416 , n86417 , n86418 , n86419 , n86420 , n86421 , n86422 , n86423 , n86424 , 
 n86425 , n86426 , n86427 , n86428 , n86429 , n86430 , n86431 , n86432 , n86433 , n86434 , 
 n86435 , n86436 , n86437 , n86438 , n86439 , n86440 , n86441 , n86442 , n86443 , n86444 , 
 n86445 , n86446 , n86447 , n86448 , n86449 , n86450 , n86451 , n86452 , n86453 , n86454 , 
 n86455 , n86456 , n86457 , n86458 , n86459 , n86460 , n86461 , n86462 , n86463 , n86464 , 
 n86465 , n86466 , n86467 , n86468 , n86469 , n86470 , n86471 , n86472 , n86473 , n86474 , 
 n86475 , n86476 , n86477 , n86478 , n86479 , n86480 , n86481 , n86482 , n86483 , n86484 , 
 n86485 , n86486 , n86487 , n86488 , n86489 , n86490 , n86491 , n86492 , n86493 , n86494 , 
 n86495 , n86496 , n86497 , n86498 , n86499 , n86500 , n86501 , n86502 , n86503 , n86504 , 
 n86505 , n86506 , n86507 , n86508 , n86509 , n86510 , n86511 , n86512 , n86513 , n86514 , 
 n86515 , n86516 , n86517 , n86518 , n86519 , n86520 , n86521 , n86522 , n86523 , n86524 , 
 n86525 , n86526 , n86527 , n86528 , n86529 , n86530 , n86531 , n86532 , n86533 , n86534 , 
 n86535 , n86536 , n86537 , n86538 , n86539 , n86540 , n86541 , n86542 , n86543 , n86544 , 
 n86545 , n86546 , n86547 , n86548 , n86549 , n86550 , n86551 , n86552 , n86553 , n86554 , 
 n86555 , n86556 , n86557 , n86558 , n86559 , n86560 , n86561 , n86562 , n86563 , n86564 , 
 n86565 , n86566 , n86567 , n86568 , n86569 , n86570 , n86571 , n86572 , n86573 , n86574 , 
 n86575 , n86576 , n86577 , n86578 , n86579 , n86580 , n86581 , n86582 , n86583 , n86584 , 
 n86585 , n86586 , n86587 , n86588 , n86589 , n86590 , n86591 , n86592 , n86593 , n86594 , 
 n86595 , n86596 , n86597 , n86598 , n86599 , n86600 , n86601 , n86602 , n86603 , n86604 , 
 n86605 , n86606 , n86607 , n86608 , n86609 , n86610 , n86611 , n86612 , n86613 , n86614 , 
 n86615 , n86616 , n86617 , n86618 , n86619 , n86620 , n86621 , n86622 , n86623 , n86624 , 
 n86625 , n86626 , n86627 , n86628 , n86629 , n86630 , n86631 , n86632 , n86633 , n86634 , 
 n86635 , n86636 , n86637 , n86638 , n86639 , n86640 , n86641 , n86642 , n86643 , n86644 , 
 n86645 , n86646 , n86647 , n86648 , n86649 , n86650 , n86651 , n86652 , n86653 , n86654 , 
 n86655 , n86656 , n86657 , n86658 , n86659 , n86660 , n86661 , n86662 , n86663 , n86664 , 
 n86665 , n86666 , n86667 , n86668 , n86669 , n86670 , n86671 , n86672 , n86673 , n86674 , 
 n86675 , n86676 , n86677 , n86678 , n86679 , n86680 , n86681 , n86682 , n86683 , n86684 , 
 n86685 , n86686 , n86687 , n86688 , n86689 , n86690 , n86691 , n86692 , n86693 , n86694 , 
 n86695 , n86696 , n86697 , n86698 , n86699 , n86700 , n86701 , n86702 , n86703 , n86704 , 
 n86705 , n86706 , n86707 , n86708 , n86709 , n86710 , n86711 , n86712 , n86713 , n86714 , 
 n86715 , n86716 , n86717 , n86718 , n86719 , n86720 , n86721 , n86722 , n86723 , n86724 , 
 n86725 , n86726 , n86727 , n86728 , n86729 , n86730 , n86731 , n86732 , n86733 , n86734 , 
 n86735 , n86736 , n86737 , n86738 , n86739 , n86740 , n86741 , n86742 , n86743 , n86744 , 
 n86745 , n86746 , n86747 , n86748 , n86749 , n86750 , n86751 , n86752 , n86753 , n86754 , 
 n86755 , n86756 , n86757 , n86758 , n86759 , n86760 , n86761 , n86762 , n86763 , n86764 , 
 n86765 , n86766 , n86767 , n86768 , n86769 , n86770 , n86771 , n86772 , n86773 , n86774 , 
 n86775 , n86776 , n86777 , n86778 , n86779 , n86780 , n86781 , n86782 , n86783 , n86784 , 
 n86785 , n86786 , n86787 , n86788 , n86789 , n86790 , n86791 , n86792 , n86793 , n86794 , 
 n86795 , n86796 , n86797 , n86798 , n86799 , n86800 , n86801 , n86802 , n86803 , n86804 , 
 n86805 , n86806 , n86807 , n86808 , n86809 , n86810 , n86811 , n86812 , n86813 , n86814 , 
 n86815 , n86816 , n86817 , n86818 , n86819 , n86820 , n86821 , n86822 , n86823 , n86824 , 
 n86825 , n86826 , n86827 , n86828 , n86829 , n86830 , n86831 , n86832 , n86833 , n86834 , 
 n86835 , n86836 , n86837 , n86838 , n86839 , n86840 , n86841 , n86842 , n86843 , n86844 , 
 n86845 , n86846 , n86847 , n86848 , n86849 , n86850 , n86851 , n86852 , n86853 , n86854 , 
 n86855 , n86856 , n86857 , n86858 , n86859 , n86860 , n86861 , n86862 , n86863 , n86864 , 
 n86865 , n86866 , n86867 , n86868 , n86869 , n86870 , n86871 , n86872 , n86873 , n86874 , 
 n86875 , n86876 , n86877 , n86878 , n86879 , n86880 , n86881 , n86882 , n86883 , n86884 , 
 n86885 , n86886 , n86887 , n86888 , n86889 , n86890 , n86891 , n86892 , n86893 , n86894 , 
 n86895 , n86896 , n86897 , n86898 , n86899 , n86900 , n86901 , n86902 , n86903 , n86904 , 
 n86905 , n86906 , n86907 , n86908 , n86909 , n86910 , n86911 , n86912 , n86913 , n86914 , 
 n86915 , n86916 , n86917 , n86918 , n86919 , n86920 , n86921 , n86922 , n86923 , n86924 , 
 n86925 , n86926 , n86927 , n86928 , n86929 , n86930 , n86931 , n86932 , n86933 , n86934 , 
 n86935 , n86936 , n86937 , n86938 , n86939 , n86940 , n86941 , n86942 , n86943 , n86944 , 
 n86945 , n86946 , n86947 , n86948 , n86949 , n86950 , n86951 , n86952 , n86953 , n86954 , 
 n86955 , n86956 , n86957 , n86958 , n86959 , n86960 , n86961 , n86962 , n86963 , n86964 , 
 n86965 , n86966 , n86967 , n86968 , n86969 , n86970 , n86971 , n86972 , n86973 , n86974 , 
 n86975 , n86976 , n86977 , n86978 , n86979 , n86980 , n86981 , n86982 , n86983 , n86984 , 
 n86985 , n86986 , n86987 , n86988 , n86989 , n86990 , n86991 , n86992 , n86993 , n86994 , 
 n86995 , n86996 , n86997 , n86998 , n86999 , n87000 , n87001 , n87002 , n87003 , n87004 , 
 n87005 , n87006 , n87007 , n87008 , n87009 , n87010 , n87011 , n87012 , n87013 , n87014 , 
 n87015 , n87016 , n87017 , n87018 , n87019 , n87020 , n87021 , n87022 , n87023 , n87024 , 
 n87025 , n87026 , n87027 , n87028 , n87029 , n87030 , n87031 , n87032 , n87033 , n87034 , 
 n87035 , n87036 , n87037 , n87038 , n87039 , n87040 , n87041 , n87042 , n87043 , n87044 , 
 n87045 , n87046 , n87047 , n87048 , n87049 , n87050 , n87051 , n87052 , n87053 , n87054 , 
 n87055 , n87056 , n87057 , n87058 , n87059 , n87060 , n87061 , n87062 , n87063 , n87064 , 
 n87065 , n87066 , n87067 , n87068 , n87069 , n87070 , n87071 , n87072 , n87073 , n87074 , 
 n87075 , n87076 , n87077 , n87078 , n87079 , n87080 , n87081 , n87082 , n87083 , n87084 , 
 n87085 , n87086 , n87087 , n87088 , n87089 , n87090 , n87091 , n87092 , n87093 , n87094 , 
 n87095 , n87096 , n87097 , n87098 , n87099 , n87100 , n87101 , n87102 , n87103 , n87104 , 
 n87105 , n87106 , n87107 , n87108 , n87109 , n87110 , n87111 , n87112 , n87113 , n87114 , 
 n87115 , n87116 , n87117 , n87118 , n87119 , n87120 , n87121 , n87122 , n87123 , n87124 , 
 n87125 , n87126 , n87127 , n87128 , n87129 , n87130 , n87131 , n87132 , n87133 , n87134 , 
 n87135 , n87136 , n87137 , n87138 , n87139 , n87140 , n87141 , n87142 , n87143 , n87144 , 
 n87145 , n87146 , n87147 , n87148 , n87149 , n87150 , n87151 , n87152 , n87153 , n87154 , 
 n87155 , n87156 , n87157 , n87158 , n87159 , n87160 , n87161 , n87162 , n87163 , n87164 , 
 n87165 , n87166 , n87167 , n87168 , n87169 , n87170 , n87171 , n87172 , n87173 , n87174 , 
 n87175 , n87176 , n87177 , n87178 , n87179 , n87180 , n87181 , n87182 , n87183 , n87184 , 
 n87185 , n87186 , n87187 , n87188 , n87189 , n87190 , n87191 , n87192 , n87193 , n87194 , 
 n87195 , n87196 , n87197 , n87198 , n87199 , n87200 , n87201 , n87202 , n87203 , n87204 , 
 n87205 , n87206 , n87207 , n87208 , n87209 , n87210 , n87211 , n87212 , n87213 , n87214 , 
 n87215 , n87216 , n87217 , n87218 , n87219 , n87220 , n87221 , n87222 , n87223 , n87224 , 
 n87225 , n87226 , n87227 , n87228 , n87229 , n87230 , n87231 , n87232 , n87233 , n87234 , 
 n87235 , n87236 , n87237 , n87238 , n87239 , n87240 , n87241 , n87242 , n87243 , n87244 , 
 n87245 , n87246 , n87247 , n87248 , n87249 , n87250 , n87251 , n87252 , n87253 , n87254 , 
 n87255 , n87256 , n87257 , n87258 , n87259 , n87260 , n87261 , n87262 , n87263 , n87264 , 
 n87265 , n87266 , n87267 , n87268 , n87269 , n87270 , n87271 , n87272 , n87273 , n87274 , 
 n87275 , n87276 , n87277 , n87278 , n87279 , n87280 , n87281 , n87282 , n87283 , n87284 , 
 n87285 , n87286 , n87287 , n87288 , n87289 , n87290 , n87291 , n87292 , n87293 , n87294 , 
 n87295 , n87296 , n87297 , n87298 , n87299 , n87300 , n87301 , n87302 , n87303 , n87304 , 
 n87305 , n87306 , n87307 , n87308 , n87309 , n87310 , n87311 , n87312 , n87313 , n87314 , 
 n87315 , n87316 , n87317 , n87318 , n87319 , n87320 , n87321 , n87322 , n87323 , n87324 , 
 n87325 , n87326 , n87327 , n87328 , n87329 , n87330 , n87331 , n87332 , n87333 , n87334 , 
 n87335 , n87336 , n87337 , n87338 , n87339 , n87340 , n87341 , n87342 , n87343 , n87344 , 
 n87345 , n87346 , n87347 , n87348 , n87349 , n87350 , n87351 , n87352 , n87353 , n87354 , 
 n87355 , n87356 , n87357 , n87358 , n87359 , n87360 , n87361 , n87362 , n87363 , n87364 , 
 n87365 , n87366 , n87367 , n87368 , n87369 , n87370 , n87371 , n87372 , n87373 , n87374 , 
 n87375 , n87376 , n87377 , n87378 , n87379 , n87380 , n87381 , n87382 , n87383 , n87384 , 
 n87385 , n87386 , n87387 , n87388 , n87389 , n87390 , n87391 , n87392 , n87393 , n87394 , 
 n87395 , n87396 , n87397 , n87398 , n87399 , n87400 , n87401 , n87402 , n87403 , n87404 , 
 n87405 , n87406 , n87407 , n87408 , n87409 , n87410 , n87411 , n87412 , n87413 , n87414 , 
 n87415 , n87416 , n87417 , n87418 , n87419 , n87420 , n87421 , n87422 , n87423 , n87424 , 
 n87425 , n87426 , n87427 , n87428 , n87429 , n87430 , n87431 , n87432 , n87433 , n87434 , 
 n87435 , n87436 , n87437 , n87438 , n87439 , n87440 , n87441 , n87442 , n87443 , n87444 , 
 n87445 , n87446 , n87447 , n87448 , n87449 , n87450 , n87451 , n87452 , n87453 , n87454 , 
 n87455 , n87456 , n87457 , n87458 , n87459 , n87460 , n87461 , n87462 , n87463 , n87464 , 
 n87465 , n87466 , n87467 , n87468 , n87469 , n87470 , n87471 , n87472 , n87473 , n87474 , 
 n87475 , n87476 , n87477 , n87478 , n87479 , n87480 , n87481 , n87482 , n87483 , n87484 , 
 n87485 , n87486 , n87487 , n87488 , n87489 , n87490 , n87491 , n87492 , n87493 , n87494 , 
 n87495 , n87496 , n87497 , n87498 , n87499 , n87500 , n87501 , n87502 , n87503 , n87504 , 
 n87505 , n87506 , n87507 , n87508 , n87509 , n87510 , n87511 , n87512 , n87513 , n87514 , 
 n87515 , n87516 , n87517 , n87518 , n87519 , n87520 , n87521 , n87522 , n87523 , n87524 , 
 n87525 , n87526 , n87527 , n87528 , n87529 , n87530 , n87531 , n87532 , n87533 , n87534 , 
 n87535 , n87536 , n87537 , n87538 , n87539 , n87540 , n87541 , n87542 , n87543 , n87544 , 
 n87545 , n87546 , n87547 , n87548 , n87549 , n87550 , n87551 , n87552 , n87553 , n87554 , 
 n87555 , n87556 , n87557 , n87558 , n87559 , n87560 , n87561 , n87562 , n87563 , n87564 , 
 n87565 , n87566 , n87567 , n87568 , n87569 , n87570 , n87571 , n87572 , n87573 , n87574 , 
 n87575 , n87576 , n87577 , n87578 , n87579 , n87580 , n87581 , n87582 , n87583 , n87584 , 
 n87585 , n87586 , n87587 , n87588 , n87589 , n87590 ;
buf ( n544 , n0 );
buf ( n545 , n1 );
buf ( n546 , n2 );
buf ( n547 , n3 );
buf ( n548 , n4 );
buf ( n549 , n5 );
buf ( n550 , n6 );
buf ( n551 , n7 );
buf ( n552 , n8 );
buf ( n553 , n9 );
buf ( n554 , n10 );
buf ( n555 , n11 );
buf ( n556 , n12 );
buf ( n557 , n13 );
buf ( n558 , n14 );
buf ( n559 , n15 );
buf ( n560 , n16 );
buf ( n561 , n17 );
buf ( n562 , n18 );
buf ( n563 , n19 );
buf ( n564 , n20 );
buf ( n565 , n21 );
buf ( n566 , n22 );
buf ( n567 , n23 );
buf ( n568 , n24 );
buf ( n569 , n25 );
buf ( n570 , n26 );
buf ( n571 , n27 );
buf ( n572 , n28 );
buf ( n573 , n29 );
buf ( n574 , n30 );
buf ( n575 , n31 );
buf ( n576 , n32 );
buf ( n577 , n33 );
buf ( n578 , n34 );
buf ( n579 , n35 );
buf ( n580 , n36 );
buf ( n581 , n37 );
buf ( n582 , n38 );
buf ( n583 , n39 );
buf ( n584 , n40 );
buf ( n585 , n41 );
buf ( n586 , n42 );
buf ( n587 , n43 );
buf ( n588 , n44 );
buf ( n589 , n45 );
buf ( n590 , n46 );
buf ( n591 , n47 );
buf ( n592 , n48 );
buf ( n593 , n49 );
buf ( n594 , n50 );
buf ( n595 , n51 );
buf ( n596 , n52 );
buf ( n597 , n53 );
buf ( n598 , n54 );
buf ( n599 , n55 );
buf ( n600 , n56 );
buf ( n601 , n57 );
buf ( n602 , n58 );
buf ( n603 , n59 );
buf ( n604 , n60 );
buf ( n605 , n61 );
buf ( n606 , n62 );
buf ( n607 , n63 );
buf ( n608 , n64 );
buf ( n609 , n65 );
buf ( n610 , n66 );
buf ( n611 , n67 );
buf ( n612 , n68 );
buf ( n613 , n69 );
buf ( n614 , n70 );
buf ( n615 , n71 );
buf ( n616 , n72 );
buf ( n617 , n73 );
buf ( n618 , n74 );
buf ( n619 , n75 );
buf ( n620 , n76 );
buf ( n621 , n77 );
buf ( n622 , n78 );
buf ( n623 , n79 );
buf ( n80 , n624 );
buf ( n81 , n625 );
buf ( n82 , n626 );
buf ( n83 , n627 );
buf ( n84 , n628 );
buf ( n85 , n629 );
buf ( n86 , n630 );
buf ( n87 , n631 );
buf ( n88 , n632 );
buf ( n89 , n633 );
buf ( n90 , n634 );
buf ( n91 , n635 );
buf ( n92 , n636 );
buf ( n93 , n637 );
buf ( n94 , n638 );
buf ( n95 , n639 );
buf ( n96 , n640 );
buf ( n97 , n641 );
buf ( n98 , n642 );
buf ( n99 , n643 );
buf ( n100 , n644 );
buf ( n101 , n645 );
buf ( n102 , n646 );
buf ( n103 , n647 );
buf ( n104 , n648 );
buf ( n105 , n649 );
buf ( n106 , n650 );
buf ( n107 , n651 );
buf ( n108 , n652 );
buf ( n109 , n653 );
buf ( n110 , n654 );
buf ( n111 , n655 );
buf ( n112 , n656 );
buf ( n113 , n657 );
buf ( n114 , n658 );
buf ( n115 , n659 );
buf ( n116 , n660 );
buf ( n117 , n661 );
buf ( n118 , n662 );
buf ( n119 , n663 );
buf ( n120 , n664 );
buf ( n121 , n665 );
buf ( n122 , n666 );
buf ( n123 , n667 );
buf ( n124 , n668 );
buf ( n125 , n669 );
buf ( n126 , n670 );
buf ( n127 , n671 );
buf ( n128 , n672 );
buf ( n129 , n673 );
buf ( n130 , n674 );
buf ( n131 , n675 );
buf ( n132 , n676 );
buf ( n133 , n677 );
buf ( n134 , n678 );
buf ( n135 , n679 );
buf ( n136 , n680 );
buf ( n137 , n681 );
buf ( n138 , n682 );
buf ( n139 , n683 );
buf ( n140 , n684 );
buf ( n141 , n685 );
buf ( n142 , n686 );
buf ( n143 , n687 );
buf ( n144 , n688 );
buf ( n145 , n689 );
buf ( n146 , n690 );
buf ( n147 , n691 );
buf ( n148 , n692 );
buf ( n149 , n693 );
buf ( n150 , n694 );
buf ( n151 , n695 );
buf ( n152 , n696 );
buf ( n153 , n697 );
buf ( n154 , n698 );
buf ( n155 , n699 );
buf ( n156 , n700 );
buf ( n157 , n701 );
buf ( n158 , n702 );
buf ( n159 , n703 );
buf ( n160 , n704 );
buf ( n161 , n705 );
buf ( n162 , n706 );
buf ( n163 , n707 );
buf ( n164 , n708 );
buf ( n165 , n709 );
buf ( n166 , n710 );
buf ( n167 , n711 );
buf ( n168 , n712 );
buf ( n169 , n713 );
buf ( n170 , n714 );
buf ( n171 , n715 );
buf ( n172 , n716 );
buf ( n173 , n717 );
buf ( n174 , n718 );
buf ( n175 , n719 );
buf ( n176 , n720 );
buf ( n177 , n721 );
buf ( n178 , n722 );
buf ( n179 , n723 );
buf ( n180 , n724 );
buf ( n181 , n725 );
buf ( n182 , n726 );
buf ( n183 , n727 );
buf ( n184 , n728 );
buf ( n185 , n729 );
buf ( n186 , n730 );
buf ( n187 , n731 );
buf ( n188 , n732 );
buf ( n189 , n733 );
buf ( n190 , n734 );
buf ( n191 , n735 );
buf ( n192 , n736 );
buf ( n193 , n737 );
buf ( n194 , n738 );
buf ( n195 , n739 );
buf ( n196 , n740 );
buf ( n197 , n741 );
buf ( n198 , n742 );
buf ( n199 , n743 );
buf ( n200 , n744 );
buf ( n201 , n745 );
buf ( n202 , n746 );
buf ( n203 , n747 );
buf ( n204 , n748 );
buf ( n205 , n749 );
buf ( n206 , n750 );
buf ( n207 , n751 );
buf ( n208 , n752 );
buf ( n209 , n753 );
buf ( n210 , n754 );
buf ( n211 , n755 );
buf ( n212 , n756 );
buf ( n213 , n757 );
buf ( n214 , n758 );
buf ( n215 , n759 );
buf ( n216 , n760 );
buf ( n217 , n761 );
buf ( n218 , n762 );
buf ( n219 , n763 );
buf ( n220 , n764 );
buf ( n221 , n765 );
buf ( n222 , n766 );
buf ( n223 , n767 );
buf ( n224 , n768 );
buf ( n225 , n769 );
buf ( n226 , n770 );
buf ( n227 , n771 );
buf ( n228 , n772 );
buf ( n229 , n773 );
buf ( n230 , n774 );
buf ( n231 , n775 );
buf ( n232 , n776 );
buf ( n233 , n777 );
buf ( n234 , n778 );
buf ( n235 , n779 );
buf ( n236 , n780 );
buf ( n237 , n781 );
buf ( n238 , n782 );
buf ( n239 , n783 );
buf ( n240 , n784 );
buf ( n241 , n785 );
buf ( n242 , n786 );
buf ( n243 , n787 );
buf ( n244 , n788 );
buf ( n245 , n789 );
buf ( n246 , n790 );
buf ( n247 , n791 );
buf ( n248 , n792 );
buf ( n249 , n793 );
buf ( n250 , n794 );
buf ( n251 , n795 );
buf ( n252 , n796 );
buf ( n253 , n797 );
buf ( n254 , n798 );
buf ( n255 , n799 );
buf ( n256 , n800 );
buf ( n257 , n801 );
buf ( n258 , n802 );
buf ( n259 , n803 );
buf ( n260 , n804 );
buf ( n261 , n805 );
buf ( n262 , n806 );
buf ( n263 , n807 );
buf ( n264 , n808 );
buf ( n265 , n809 );
buf ( n266 , n810 );
buf ( n267 , n811 );
buf ( n268 , n812 );
buf ( n269 , n813 );
buf ( n270 , n814 );
buf ( n271 , n815 );
buf ( n624 , n87528 );
buf ( n625 , n87530 );
buf ( n626 , n87532 );
buf ( n627 , n87534 );
buf ( n628 , n87536 );
buf ( n629 , n87538 );
buf ( n630 , n87540 );
buf ( n631 , n87542 );
buf ( n632 , n87544 );
buf ( n633 , n87546 );
buf ( n634 , n87548 );
buf ( n635 , n87550 );
buf ( n636 , n87552 );
buf ( n637 , n87554 );
buf ( n638 , n87556 );
buf ( n639 , n87558 );
buf ( n640 , n87560 );
buf ( n641 , n87562 );
buf ( n642 , n87564 );
buf ( n643 , n87566 );
buf ( n644 , n87568 );
buf ( n645 , n87570 );
buf ( n646 , n87572 );
buf ( n647 , n87574 );
buf ( n648 , n87576 );
buf ( n649 , n87578 );
buf ( n650 , n87580 );
buf ( n651 , n87582 );
buf ( n652 , n87584 );
buf ( n653 , n87586 );
buf ( n654 , n87588 );
buf ( n655 , n87590 );
buf ( n656 , n85579 );
buf ( n657 , n85581 );
buf ( n658 , n85583 );
buf ( n659 , n85585 );
buf ( n660 , n85587 );
buf ( n661 , n85589 );
buf ( n662 , n85591 );
buf ( n663 , n85593 );
buf ( n664 , n85595 );
buf ( n665 , n85597 );
buf ( n666 , n85599 );
buf ( n667 , n85601 );
buf ( n668 , n85603 );
buf ( n669 , n85605 );
buf ( n670 , n85607 );
buf ( n671 , n85609 );
buf ( n672 , n85611 );
buf ( n673 , n85613 );
buf ( n674 , n85615 );
buf ( n675 , n85617 );
buf ( n676 , n85619 );
buf ( n677 , n85621 );
buf ( n678 , n85623 );
buf ( n679 , n85625 );
buf ( n680 , n85627 );
buf ( n681 , n85629 );
buf ( n682 , n85631 );
buf ( n683 , n85633 );
buf ( n684 , n85635 );
buf ( n685 , n85637 );
buf ( n686 , n85639 );
buf ( n687 , n85641 );
buf ( n688 , n83568 );
buf ( n689 , n83570 );
buf ( n690 , n83572 );
buf ( n691 , n83574 );
buf ( n692 , n83576 );
buf ( n693 , n83578 );
buf ( n694 , n83580 );
buf ( n695 , n83582 );
buf ( n696 , n83584 );
buf ( n697 , n83586 );
buf ( n698 , n83588 );
buf ( n699 , n83590 );
buf ( n700 , n83592 );
buf ( n701 , n83594 );
buf ( n702 , n83596 );
buf ( n703 , n83598 );
buf ( n704 , n83600 );
buf ( n705 , n83602 );
buf ( n706 , n83604 );
buf ( n707 , n83606 );
buf ( n708 , n83608 );
buf ( n709 , n83610 );
buf ( n710 , n83612 );
buf ( n711 , n83614 );
buf ( n712 , n83616 );
buf ( n713 , n83618 );
buf ( n714 , n83620 );
buf ( n715 , n83622 );
buf ( n716 , n83624 );
buf ( n717 , n83626 );
buf ( n718 , n83628 );
buf ( n719 , n83630 );
buf ( n720 , n83632 );
buf ( n721 , n83634 );
buf ( n722 , n83636 );
buf ( n723 , n83638 );
buf ( n724 , n83640 );
buf ( n725 , n83642 );
buf ( n726 , n83644 );
buf ( n727 , n83646 );
buf ( n728 , n83648 );
buf ( n729 , n83650 );
buf ( n730 , n83652 );
buf ( n731 , n83654 );
buf ( n732 , n83656 );
buf ( n733 , n83658 );
buf ( n734 , n83660 );
buf ( n735 , n83662 );
buf ( n736 , n83664 );
buf ( n737 , n83666 );
buf ( n738 , n83668 );
buf ( n739 , n83670 );
buf ( n740 , n83672 );
buf ( n741 , n83674 );
buf ( n742 , n83676 );
buf ( n743 , n83678 );
buf ( n744 , n83680 );
buf ( n745 , n83682 );
buf ( n746 , n83684 );
buf ( n747 , n83686 );
buf ( n748 , n83688 );
buf ( n749 , n83690 );
buf ( n750 , n83692 );
buf ( n751 , n83694 );
buf ( n752 , n83696 );
buf ( n753 , n83698 );
buf ( n754 , n83700 );
buf ( n755 , n83702 );
buf ( n756 , n83704 );
buf ( n757 , n83706 );
buf ( n758 , n83708 );
buf ( n759 , n83710 );
buf ( n760 , n83712 );
buf ( n761 , n83714 );
buf ( n762 , n83716 );
buf ( n763 , n83718 );
buf ( n764 , n83720 );
buf ( n765 , n83722 );
buf ( n766 , n83724 );
buf ( n767 , n83727 );
buf ( n768 , n83730 );
buf ( n769 , n83733 );
buf ( n770 , n83736 );
buf ( n771 , n83739 );
buf ( n772 , n83742 );
buf ( n773 , n83745 );
buf ( n774 , n83748 );
buf ( n775 , n83751 );
buf ( n776 , n83754 );
buf ( n777 , n83757 );
buf ( n778 , n83760 );
buf ( n779 , n83763 );
buf ( n780 , n83766 );
buf ( n781 , n83769 );
buf ( n782 , n83772 );
buf ( n783 , n83775 );
buf ( n784 , n83778 );
buf ( n785 , n83781 );
buf ( n786 , n83784 );
buf ( n787 , n83787 );
buf ( n788 , n83790 );
buf ( n789 , n83793 );
buf ( n790 , n83796 );
buf ( n791 , n83799 );
buf ( n792 , n83802 );
buf ( n793 , n83805 );
buf ( n794 , n83808 );
buf ( n795 , n83811 );
buf ( n796 , n83814 );
buf ( n797 , n83817 );
buf ( n798 , n83820 );
buf ( n799 , n83823 );
buf ( n800 , n83826 );
buf ( n801 , n83829 );
buf ( n802 , n83832 );
buf ( n803 , n83835 );
buf ( n804 , n83838 );
buf ( n805 , n83841 );
buf ( n806 , n83844 );
buf ( n807 , n83847 );
buf ( n808 , n83850 );
buf ( n809 , n83853 );
buf ( n810 , n83856 );
buf ( n811 , n83859 );
buf ( n812 , n83862 );
buf ( n813 , n83865 );
buf ( n814 , n83868 );
buf ( n815 , n83870 );
buf ( n816 , n592 );
buf ( n817 , n593 );
buf ( n818 , n594 );
buf ( n819 , n595 );
buf ( n820 , n596 );
buf ( n821 , n597 );
buf ( n822 , n598 );
buf ( n823 , n599 );
buf ( n824 , n600 );
buf ( n825 , n601 );
buf ( n826 , n602 );
buf ( n827 , n603 );
buf ( n828 , n604 );
buf ( n829 , n605 );
buf ( n830 , n606 );
buf ( n831 , n607 );
buf ( n832 , n562 );
buf ( n833 , n832 );
buf ( n834 , n563 );
buf ( n835 , n834 );
buf ( n836 , n564 );
buf ( n837 , n836 );
and ( n838 , n835 , n837 );
not ( n839 , n838 );
and ( n840 , n833 , n839 );
not ( n841 , n840 );
buf ( n842 , n545 );
buf ( n843 , n842 );
buf ( n844 , n560 );
buf ( n845 , n844 );
buf ( n846 , n561 );
buf ( n847 , n846 );
xor ( n848 , n845 , n847 );
xor ( n849 , n847 , n833 );
not ( n850 , n849 );
and ( n851 , n848 , n850 );
and ( n852 , n843 , n851 );
buf ( n853 , n544 );
buf ( n854 , n853 );
and ( n855 , n854 , n849 );
nor ( n856 , n852 , n855 );
and ( n857 , n847 , n833 );
not ( n858 , n857 );
and ( n859 , n845 , n858 );
xnor ( n860 , n856 , n859 );
and ( n861 , n841 , n860 );
buf ( n862 , n546 );
buf ( n863 , n862 );
and ( n864 , n863 , n845 );
and ( n865 , n860 , n864 );
and ( n866 , n841 , n864 );
or ( n867 , n861 , n865 , n866 );
and ( n868 , n854 , n851 );
not ( n869 , n868 );
xnor ( n870 , n869 , n859 );
and ( n871 , n867 , n870 );
and ( n872 , n843 , n845 );
not ( n873 , n872 );
and ( n874 , n870 , n873 );
and ( n875 , n867 , n873 );
or ( n876 , n871 , n874 , n875 );
buf ( n877 , n544 );
buf ( n878 , n877 );
buf ( n879 , n578 );
buf ( n880 , n879 );
buf ( n881 , n579 );
buf ( n882 , n881 );
xor ( n883 , n880 , n882 );
buf ( n884 , n580 );
buf ( n885 , n884 );
xor ( n886 , n882 , n885 );
not ( n887 , n886 );
and ( n888 , n883 , n887 );
and ( n889 , n878 , n888 );
not ( n890 , n889 );
and ( n891 , n882 , n885 );
not ( n892 , n891 );
and ( n893 , n880 , n892 );
xnor ( n894 , n890 , n893 );
not ( n895 , n894 );
buf ( n896 , n546 );
buf ( n897 , n896 );
buf ( n898 , n576 );
buf ( n899 , n898 );
buf ( n900 , n577 );
buf ( n901 , n900 );
xor ( n902 , n899 , n901 );
xor ( n903 , n901 , n880 );
not ( n904 , n903 );
and ( n905 , n902 , n904 );
and ( n906 , n897 , n905 );
buf ( n907 , n545 );
buf ( n908 , n907 );
and ( n909 , n908 , n903 );
nor ( n910 , n906 , n909 );
and ( n911 , n901 , n880 );
not ( n912 , n911 );
and ( n913 , n899 , n912 );
xnor ( n914 , n910 , n913 );
and ( n915 , n895 , n914 );
buf ( n916 , n547 );
buf ( n917 , n916 );
and ( n918 , n917 , n899 );
and ( n919 , n914 , n918 );
and ( n920 , n895 , n918 );
or ( n921 , n915 , n919 , n920 );
buf ( n922 , n894 );
and ( n923 , n921 , n922 );
not ( n924 , n893 );
and ( n925 , n908 , n905 );
and ( n926 , n878 , n903 );
nor ( n927 , n925 , n926 );
xnor ( n928 , n927 , n913 );
xor ( n929 , n924 , n928 );
and ( n930 , n897 , n899 );
xor ( n931 , n929 , n930 );
and ( n932 , n922 , n931 );
and ( n933 , n921 , n931 );
or ( n934 , n923 , n932 , n933 );
xor ( n935 , n867 , n870 );
xor ( n936 , n935 , n873 );
and ( n937 , n934 , n936 );
and ( n938 , n924 , n928 );
and ( n939 , n928 , n930 );
and ( n940 , n924 , n930 );
or ( n941 , n938 , n939 , n940 );
and ( n942 , n878 , n905 );
not ( n943 , n942 );
xnor ( n944 , n943 , n913 );
xor ( n945 , n941 , n944 );
and ( n946 , n908 , n899 );
not ( n947 , n946 );
xor ( n948 , n945 , n947 );
and ( n949 , n936 , n948 );
and ( n950 , n934 , n948 );
or ( n951 , n937 , n949 , n950 );
xor ( n952 , n876 , n951 );
and ( n953 , n941 , n944 );
and ( n954 , n944 , n947 );
and ( n955 , n941 , n947 );
or ( n956 , n953 , n954 , n955 );
buf ( n957 , n946 );
not ( n958 , n913 );
xor ( n959 , n957 , n958 );
and ( n960 , n878 , n899 );
xor ( n961 , n959 , n960 );
xor ( n962 , n956 , n961 );
buf ( n963 , n872 );
not ( n964 , n859 );
xor ( n965 , n963 , n964 );
and ( n966 , n854 , n845 );
xor ( n967 , n965 , n966 );
xor ( n968 , n962 , n967 );
xor ( n969 , n952 , n968 );
xor ( n970 , n833 , n835 );
xor ( n971 , n835 , n837 );
not ( n972 , n971 );
and ( n973 , n970 , n972 );
and ( n974 , n854 , n973 );
not ( n975 , n974 );
xnor ( n976 , n975 , n840 );
not ( n977 , n976 );
and ( n978 , n863 , n851 );
and ( n979 , n843 , n849 );
nor ( n980 , n978 , n979 );
xnor ( n981 , n980 , n859 );
and ( n982 , n977 , n981 );
buf ( n983 , n547 );
buf ( n984 , n983 );
and ( n985 , n984 , n845 );
and ( n986 , n981 , n985 );
and ( n987 , n977 , n985 );
or ( n988 , n982 , n986 , n987 );
buf ( n989 , n976 );
and ( n990 , n988 , n989 );
xor ( n991 , n841 , n860 );
xor ( n992 , n991 , n864 );
and ( n993 , n989 , n992 );
and ( n994 , n988 , n992 );
or ( n995 , n990 , n993 , n994 );
buf ( n996 , n581 );
buf ( n997 , n996 );
buf ( n998 , n582 );
buf ( n999 , n998 );
and ( n1000 , n997 , n999 );
not ( n1001 , n1000 );
and ( n1002 , n885 , n1001 );
not ( n1003 , n1002 );
and ( n1004 , n908 , n888 );
and ( n1005 , n878 , n886 );
nor ( n1006 , n1004 , n1005 );
xnor ( n1007 , n1006 , n893 );
and ( n1008 , n1003 , n1007 );
buf ( n1009 , n548 );
buf ( n1010 , n1009 );
and ( n1011 , n1010 , n899 );
and ( n1012 , n1007 , n1011 );
and ( n1013 , n1003 , n1011 );
or ( n1014 , n1008 , n1012 , n1013 );
and ( n1015 , n897 , n888 );
and ( n1016 , n908 , n886 );
nor ( n1017 , n1015 , n1016 );
xnor ( n1018 , n1017 , n893 );
and ( n1019 , n1010 , n905 );
and ( n1020 , n917 , n903 );
nor ( n1021 , n1019 , n1020 );
xnor ( n1022 , n1021 , n913 );
and ( n1023 , n1018 , n1022 );
buf ( n1024 , n549 );
buf ( n1025 , n1024 );
and ( n1026 , n1025 , n899 );
and ( n1027 , n1022 , n1026 );
and ( n1028 , n1018 , n1026 );
or ( n1029 , n1023 , n1027 , n1028 );
xor ( n1030 , n885 , n997 );
xor ( n1031 , n997 , n999 );
not ( n1032 , n1031 );
and ( n1033 , n1030 , n1032 );
and ( n1034 , n878 , n1033 );
not ( n1035 , n1034 );
xnor ( n1036 , n1035 , n1002 );
buf ( n1037 , n1036 );
and ( n1038 , n1029 , n1037 );
and ( n1039 , n917 , n905 );
and ( n1040 , n897 , n903 );
nor ( n1041 , n1039 , n1040 );
xnor ( n1042 , n1041 , n913 );
and ( n1043 , n1037 , n1042 );
and ( n1044 , n1029 , n1042 );
or ( n1045 , n1038 , n1043 , n1044 );
and ( n1046 , n1014 , n1045 );
xor ( n1047 , n895 , n914 );
xor ( n1048 , n1047 , n918 );
and ( n1049 , n1045 , n1048 );
and ( n1050 , n1014 , n1048 );
or ( n1051 , n1046 , n1049 , n1050 );
xor ( n1052 , n988 , n989 );
xor ( n1053 , n1052 , n992 );
and ( n1054 , n1051 , n1053 );
xor ( n1055 , n921 , n922 );
xor ( n1056 , n1055 , n931 );
and ( n1057 , n1053 , n1056 );
and ( n1058 , n1051 , n1056 );
or ( n1059 , n1054 , n1057 , n1058 );
and ( n1060 , n995 , n1059 );
xor ( n1061 , n934 , n936 );
xor ( n1062 , n1061 , n948 );
and ( n1063 , n1059 , n1062 );
and ( n1064 , n995 , n1062 );
or ( n1065 , n1060 , n1063 , n1064 );
xor ( n1066 , n969 , n1065 );
xor ( n1067 , n995 , n1059 );
xor ( n1068 , n1067 , n1062 );
buf ( n1069 , n565 );
buf ( n1070 , n1069 );
buf ( n1071 , n566 );
buf ( n1072 , n1071 );
and ( n1073 , n1070 , n1072 );
not ( n1074 , n1073 );
and ( n1075 , n837 , n1074 );
not ( n1076 , n1075 );
and ( n1077 , n843 , n973 );
and ( n1078 , n854 , n971 );
nor ( n1079 , n1077 , n1078 );
xnor ( n1080 , n1079 , n840 );
and ( n1081 , n1076 , n1080 );
buf ( n1082 , n548 );
buf ( n1083 , n1082 );
and ( n1084 , n1083 , n845 );
and ( n1085 , n1080 , n1084 );
and ( n1086 , n1076 , n1084 );
or ( n1087 , n1081 , n1085 , n1086 );
and ( n1088 , n863 , n973 );
and ( n1089 , n843 , n971 );
nor ( n1090 , n1088 , n1089 );
xnor ( n1091 , n1090 , n840 );
and ( n1092 , n1083 , n851 );
and ( n1093 , n984 , n849 );
nor ( n1094 , n1092 , n1093 );
xnor ( n1095 , n1094 , n859 );
and ( n1096 , n1091 , n1095 );
buf ( n1097 , n549 );
buf ( n1098 , n1097 );
and ( n1099 , n1098 , n845 );
and ( n1100 , n1095 , n1099 );
and ( n1101 , n1091 , n1099 );
or ( n1102 , n1096 , n1100 , n1101 );
xor ( n1103 , n837 , n1070 );
xor ( n1104 , n1070 , n1072 );
not ( n1105 , n1104 );
and ( n1106 , n1103 , n1105 );
and ( n1107 , n854 , n1106 );
not ( n1108 , n1107 );
xnor ( n1109 , n1108 , n1075 );
buf ( n1110 , n1109 );
and ( n1111 , n1102 , n1110 );
and ( n1112 , n984 , n851 );
and ( n1113 , n863 , n849 );
nor ( n1114 , n1112 , n1113 );
xnor ( n1115 , n1114 , n859 );
and ( n1116 , n1110 , n1115 );
and ( n1117 , n1102 , n1115 );
or ( n1118 , n1111 , n1116 , n1117 );
and ( n1119 , n1087 , n1118 );
xor ( n1120 , n977 , n981 );
xor ( n1121 , n1120 , n985 );
and ( n1122 , n1118 , n1121 );
and ( n1123 , n1087 , n1121 );
or ( n1124 , n1119 , n1122 , n1123 );
buf ( n1125 , n583 );
buf ( n1126 , n1125 );
buf ( n1127 , n584 );
buf ( n1128 , n1127 );
and ( n1129 , n1126 , n1128 );
not ( n1130 , n1129 );
and ( n1131 , n999 , n1130 );
not ( n1132 , n1131 );
and ( n1133 , n908 , n1033 );
and ( n1134 , n878 , n1031 );
nor ( n1135 , n1133 , n1134 );
xnor ( n1136 , n1135 , n1002 );
and ( n1137 , n1132 , n1136 );
and ( n1138 , n1025 , n905 );
and ( n1139 , n1010 , n903 );
nor ( n1140 , n1138 , n1139 );
xnor ( n1141 , n1140 , n913 );
and ( n1142 , n1136 , n1141 );
and ( n1143 , n1132 , n1141 );
or ( n1144 , n1137 , n1142 , n1143 );
not ( n1145 , n1036 );
and ( n1146 , n1144 , n1145 );
xor ( n1147 , n1018 , n1022 );
xor ( n1148 , n1147 , n1026 );
and ( n1149 , n1145 , n1148 );
and ( n1150 , n1144 , n1148 );
or ( n1151 , n1146 , n1149 , n1150 );
xor ( n1152 , n1003 , n1007 );
xor ( n1153 , n1152 , n1011 );
and ( n1154 , n1151 , n1153 );
xor ( n1155 , n1029 , n1037 );
xor ( n1156 , n1155 , n1042 );
and ( n1157 , n1153 , n1156 );
and ( n1158 , n1151 , n1156 );
or ( n1159 , n1154 , n1157 , n1158 );
xor ( n1160 , n1014 , n1045 );
xor ( n1161 , n1160 , n1048 );
and ( n1162 , n1159 , n1161 );
xor ( n1163 , n1087 , n1118 );
xor ( n1164 , n1163 , n1121 );
and ( n1165 , n1161 , n1164 );
and ( n1166 , n1159 , n1164 );
or ( n1167 , n1162 , n1165 , n1166 );
and ( n1168 , n1124 , n1167 );
xor ( n1169 , n1051 , n1053 );
xor ( n1170 , n1169 , n1056 );
and ( n1171 , n1167 , n1170 );
and ( n1172 , n1124 , n1170 );
or ( n1173 , n1168 , n1171 , n1172 );
and ( n1174 , n1068 , n1173 );
xor ( n1175 , n1068 , n1173 );
xor ( n1176 , n1124 , n1167 );
xor ( n1177 , n1176 , n1170 );
buf ( n1178 , n567 );
buf ( n1179 , n1178 );
buf ( n1180 , n568 );
buf ( n1181 , n1180 );
and ( n1182 , n1179 , n1181 );
not ( n1183 , n1182 );
and ( n1184 , n1072 , n1183 );
not ( n1185 , n1184 );
and ( n1186 , n843 , n1106 );
and ( n1187 , n854 , n1104 );
nor ( n1188 , n1186 , n1187 );
xnor ( n1189 , n1188 , n1075 );
and ( n1190 , n1185 , n1189 );
and ( n1191 , n1098 , n851 );
and ( n1192 , n1083 , n849 );
nor ( n1193 , n1191 , n1192 );
xnor ( n1194 , n1193 , n859 );
and ( n1195 , n1189 , n1194 );
and ( n1196 , n1185 , n1194 );
or ( n1197 , n1190 , n1195 , n1196 );
not ( n1198 , n1109 );
and ( n1199 , n1197 , n1198 );
xor ( n1200 , n1091 , n1095 );
xor ( n1201 , n1200 , n1099 );
and ( n1202 , n1198 , n1201 );
and ( n1203 , n1197 , n1201 );
or ( n1204 , n1199 , n1202 , n1203 );
xor ( n1205 , n1076 , n1080 );
xor ( n1206 , n1205 , n1084 );
and ( n1207 , n1204 , n1206 );
xor ( n1208 , n1102 , n1110 );
xor ( n1209 , n1208 , n1115 );
and ( n1210 , n1206 , n1209 );
and ( n1211 , n1204 , n1209 );
or ( n1212 , n1207 , n1210 , n1211 );
and ( n1213 , n897 , n1033 );
and ( n1214 , n908 , n1031 );
nor ( n1215 , n1213 , n1214 );
xnor ( n1216 , n1215 , n1002 );
buf ( n1217 , n1216 );
and ( n1218 , n917 , n888 );
and ( n1219 , n897 , n886 );
nor ( n1220 , n1218 , n1219 );
xnor ( n1221 , n1220 , n893 );
and ( n1222 , n1217 , n1221 );
buf ( n1223 , n550 );
buf ( n1224 , n1223 );
and ( n1225 , n1224 , n899 );
and ( n1226 , n1221 , n1225 );
and ( n1227 , n1217 , n1225 );
or ( n1228 , n1222 , n1226 , n1227 );
xor ( n1229 , n999 , n1126 );
xor ( n1230 , n1126 , n1128 );
not ( n1231 , n1230 );
and ( n1232 , n1229 , n1231 );
and ( n1233 , n878 , n1232 );
not ( n1234 , n1233 );
xnor ( n1235 , n1234 , n1131 );
and ( n1236 , n1224 , n905 );
and ( n1237 , n1025 , n903 );
nor ( n1238 , n1236 , n1237 );
xnor ( n1239 , n1238 , n913 );
and ( n1240 , n1235 , n1239 );
buf ( n1241 , n551 );
buf ( n1242 , n1241 );
and ( n1243 , n1242 , n899 );
and ( n1244 , n1239 , n1243 );
and ( n1245 , n1235 , n1243 );
or ( n1246 , n1240 , n1244 , n1245 );
xor ( n1247 , n1132 , n1136 );
xor ( n1248 , n1247 , n1141 );
and ( n1249 , n1246 , n1248 );
xor ( n1250 , n1217 , n1221 );
xor ( n1251 , n1250 , n1225 );
and ( n1252 , n1248 , n1251 );
and ( n1253 , n1246 , n1251 );
or ( n1254 , n1249 , n1252 , n1253 );
and ( n1255 , n1228 , n1254 );
xor ( n1256 , n1144 , n1145 );
xor ( n1257 , n1256 , n1148 );
and ( n1258 , n1254 , n1257 );
and ( n1259 , n1228 , n1257 );
or ( n1260 , n1255 , n1258 , n1259 );
xor ( n1261 , n1204 , n1206 );
xor ( n1262 , n1261 , n1209 );
and ( n1263 , n1260 , n1262 );
xor ( n1264 , n1151 , n1153 );
xor ( n1265 , n1264 , n1156 );
and ( n1266 , n1262 , n1265 );
and ( n1267 , n1260 , n1265 );
or ( n1268 , n1263 , n1266 , n1267 );
and ( n1269 , n1212 , n1268 );
xor ( n1270 , n1159 , n1161 );
xor ( n1271 , n1270 , n1164 );
and ( n1272 , n1268 , n1271 );
and ( n1273 , n1212 , n1271 );
or ( n1274 , n1269 , n1272 , n1273 );
and ( n1275 , n1177 , n1274 );
xor ( n1276 , n1177 , n1274 );
xor ( n1277 , n1212 , n1268 );
xor ( n1278 , n1277 , n1271 );
and ( n1279 , n863 , n1106 );
and ( n1280 , n843 , n1104 );
nor ( n1281 , n1279 , n1280 );
xnor ( n1282 , n1281 , n1075 );
buf ( n1283 , n1282 );
and ( n1284 , n984 , n973 );
and ( n1285 , n863 , n971 );
nor ( n1286 , n1284 , n1285 );
xnor ( n1287 , n1286 , n840 );
and ( n1288 , n1283 , n1287 );
buf ( n1289 , n550 );
buf ( n1290 , n1289 );
and ( n1291 , n1290 , n845 );
and ( n1292 , n1287 , n1291 );
and ( n1293 , n1283 , n1291 );
or ( n1294 , n1288 , n1292 , n1293 );
xor ( n1295 , n1072 , n1179 );
xor ( n1296 , n1179 , n1181 );
not ( n1297 , n1296 );
and ( n1298 , n1295 , n1297 );
and ( n1299 , n854 , n1298 );
not ( n1300 , n1299 );
xnor ( n1301 , n1300 , n1184 );
and ( n1302 , n1290 , n851 );
and ( n1303 , n1098 , n849 );
nor ( n1304 , n1302 , n1303 );
xnor ( n1305 , n1304 , n859 );
and ( n1306 , n1301 , n1305 );
buf ( n1307 , n551 );
buf ( n1308 , n1307 );
and ( n1309 , n1308 , n845 );
and ( n1310 , n1305 , n1309 );
and ( n1311 , n1301 , n1309 );
or ( n1312 , n1306 , n1310 , n1311 );
xor ( n1313 , n1185 , n1189 );
xor ( n1314 , n1313 , n1194 );
and ( n1315 , n1312 , n1314 );
xor ( n1316 , n1283 , n1287 );
xor ( n1317 , n1316 , n1291 );
and ( n1318 , n1314 , n1317 );
and ( n1319 , n1312 , n1317 );
or ( n1320 , n1315 , n1318 , n1319 );
and ( n1321 , n1294 , n1320 );
xor ( n1322 , n1197 , n1198 );
xor ( n1323 , n1322 , n1201 );
and ( n1324 , n1320 , n1323 );
and ( n1325 , n1294 , n1323 );
or ( n1326 , n1321 , n1324 , n1325 );
and ( n1327 , n917 , n1033 );
and ( n1328 , n897 , n1031 );
nor ( n1329 , n1327 , n1328 );
xnor ( n1330 , n1329 , n1002 );
and ( n1331 , n1242 , n905 );
and ( n1332 , n1224 , n903 );
nor ( n1333 , n1331 , n1332 );
xnor ( n1334 , n1333 , n913 );
and ( n1335 , n1330 , n1334 );
buf ( n1336 , n552 );
buf ( n1337 , n1336 );
and ( n1338 , n1337 , n899 );
and ( n1339 , n1334 , n1338 );
and ( n1340 , n1330 , n1338 );
or ( n1341 , n1335 , n1339 , n1340 );
not ( n1342 , n1216 );
and ( n1343 , n1341 , n1342 );
and ( n1344 , n1010 , n888 );
and ( n1345 , n917 , n886 );
nor ( n1346 , n1344 , n1345 );
xnor ( n1347 , n1346 , n893 );
and ( n1348 , n1342 , n1347 );
and ( n1349 , n1341 , n1347 );
or ( n1350 , n1343 , n1348 , n1349 );
buf ( n1351 , n585 );
buf ( n1352 , n1351 );
buf ( n1353 , n586 );
buf ( n1354 , n1353 );
and ( n1355 , n1352 , n1354 );
not ( n1356 , n1355 );
and ( n1357 , n1128 , n1356 );
not ( n1358 , n1357 );
and ( n1359 , n908 , n1232 );
and ( n1360 , n878 , n1230 );
nor ( n1361 , n1359 , n1360 );
xnor ( n1362 , n1361 , n1131 );
and ( n1363 , n1358 , n1362 );
and ( n1364 , n1025 , n888 );
and ( n1365 , n1010 , n886 );
nor ( n1366 , n1364 , n1365 );
xnor ( n1367 , n1366 , n893 );
and ( n1368 , n1362 , n1367 );
and ( n1369 , n1358 , n1367 );
or ( n1370 , n1363 , n1368 , n1369 );
xor ( n1371 , n1235 , n1239 );
xor ( n1372 , n1371 , n1243 );
and ( n1373 , n1370 , n1372 );
xor ( n1374 , n1341 , n1342 );
xor ( n1375 , n1374 , n1347 );
and ( n1376 , n1372 , n1375 );
and ( n1377 , n1370 , n1375 );
or ( n1378 , n1373 , n1376 , n1377 );
and ( n1379 , n1350 , n1378 );
xor ( n1380 , n1246 , n1248 );
xor ( n1381 , n1380 , n1251 );
and ( n1382 , n1378 , n1381 );
and ( n1383 , n1350 , n1381 );
or ( n1384 , n1379 , n1382 , n1383 );
xor ( n1385 , n1294 , n1320 );
xor ( n1386 , n1385 , n1323 );
and ( n1387 , n1384 , n1386 );
xor ( n1388 , n1228 , n1254 );
xor ( n1389 , n1388 , n1257 );
and ( n1390 , n1386 , n1389 );
and ( n1391 , n1384 , n1389 );
or ( n1392 , n1387 , n1390 , n1391 );
and ( n1393 , n1326 , n1392 );
xor ( n1394 , n1260 , n1262 );
xor ( n1395 , n1394 , n1265 );
and ( n1396 , n1392 , n1395 );
and ( n1397 , n1326 , n1395 );
or ( n1398 , n1393 , n1396 , n1397 );
and ( n1399 , n1278 , n1398 );
xor ( n1400 , n1278 , n1398 );
xor ( n1401 , n1326 , n1392 );
xor ( n1402 , n1401 , n1395 );
and ( n1403 , n984 , n1106 );
and ( n1404 , n863 , n1104 );
nor ( n1405 , n1403 , n1404 );
xnor ( n1406 , n1405 , n1075 );
and ( n1407 , n1308 , n851 );
and ( n1408 , n1290 , n849 );
nor ( n1409 , n1407 , n1408 );
xnor ( n1410 , n1409 , n859 );
and ( n1411 , n1406 , n1410 );
buf ( n1412 , n552 );
buf ( n1413 , n1412 );
and ( n1414 , n1413 , n845 );
and ( n1415 , n1410 , n1414 );
and ( n1416 , n1406 , n1414 );
or ( n1417 , n1411 , n1415 , n1416 );
not ( n1418 , n1282 );
and ( n1419 , n1417 , n1418 );
and ( n1420 , n1083 , n973 );
and ( n1421 , n984 , n971 );
nor ( n1422 , n1420 , n1421 );
xnor ( n1423 , n1422 , n840 );
and ( n1424 , n1418 , n1423 );
and ( n1425 , n1417 , n1423 );
or ( n1426 , n1419 , n1424 , n1425 );
buf ( n1427 , n569 );
buf ( n1428 , n1427 );
buf ( n1429 , n570 );
buf ( n1430 , n1429 );
and ( n1431 , n1428 , n1430 );
not ( n1432 , n1431 );
and ( n1433 , n1181 , n1432 );
not ( n1434 , n1433 );
and ( n1435 , n843 , n1298 );
and ( n1436 , n854 , n1296 );
nor ( n1437 , n1435 , n1436 );
xnor ( n1438 , n1437 , n1184 );
and ( n1439 , n1434 , n1438 );
and ( n1440 , n1098 , n973 );
and ( n1441 , n1083 , n971 );
nor ( n1442 , n1440 , n1441 );
xnor ( n1443 , n1442 , n840 );
and ( n1444 , n1438 , n1443 );
and ( n1445 , n1434 , n1443 );
or ( n1446 , n1439 , n1444 , n1445 );
xor ( n1447 , n1301 , n1305 );
xor ( n1448 , n1447 , n1309 );
and ( n1449 , n1446 , n1448 );
xor ( n1450 , n1417 , n1418 );
xor ( n1451 , n1450 , n1423 );
and ( n1452 , n1448 , n1451 );
and ( n1453 , n1446 , n1451 );
or ( n1454 , n1449 , n1452 , n1453 );
and ( n1455 , n1426 , n1454 );
xor ( n1456 , n1312 , n1314 );
xor ( n1457 , n1456 , n1317 );
and ( n1458 , n1454 , n1457 );
and ( n1459 , n1426 , n1457 );
or ( n1460 , n1455 , n1458 , n1459 );
xor ( n1461 , n1128 , n1352 );
xor ( n1462 , n1352 , n1354 );
not ( n1463 , n1462 );
and ( n1464 , n1461 , n1463 );
and ( n1465 , n878 , n1464 );
not ( n1466 , n1465 );
xnor ( n1467 , n1466 , n1357 );
and ( n1468 , n1224 , n888 );
and ( n1469 , n1025 , n886 );
nor ( n1470 , n1468 , n1469 );
xnor ( n1471 , n1470 , n893 );
and ( n1472 , n1467 , n1471 );
and ( n1473 , n1337 , n905 );
and ( n1474 , n1242 , n903 );
nor ( n1475 , n1473 , n1474 );
xnor ( n1476 , n1475 , n913 );
and ( n1477 , n1471 , n1476 );
and ( n1478 , n1467 , n1476 );
or ( n1479 , n1472 , n1477 , n1478 );
and ( n1480 , n897 , n1232 );
and ( n1481 , n908 , n1230 );
nor ( n1482 , n1480 , n1481 );
xnor ( n1483 , n1482 , n1131 );
buf ( n1484 , n1483 );
and ( n1485 , n1479 , n1484 );
xor ( n1486 , n1330 , n1334 );
xor ( n1487 , n1486 , n1338 );
and ( n1488 , n1484 , n1487 );
and ( n1489 , n1479 , n1487 );
or ( n1490 , n1485 , n1488 , n1489 );
not ( n1491 , n1483 );
and ( n1492 , n1010 , n1033 );
and ( n1493 , n917 , n1031 );
nor ( n1494 , n1492 , n1493 );
xnor ( n1495 , n1494 , n1002 );
and ( n1496 , n1491 , n1495 );
buf ( n1497 , n553 );
buf ( n1498 , n1497 );
and ( n1499 , n1498 , n899 );
and ( n1500 , n1495 , n1499 );
and ( n1501 , n1491 , n1499 );
or ( n1502 , n1496 , n1500 , n1501 );
xor ( n1503 , n1358 , n1362 );
xor ( n1504 , n1503 , n1367 );
and ( n1505 , n1502 , n1504 );
xor ( n1506 , n1479 , n1484 );
xor ( n1507 , n1506 , n1487 );
and ( n1508 , n1504 , n1507 );
and ( n1509 , n1502 , n1507 );
or ( n1510 , n1505 , n1508 , n1509 );
and ( n1511 , n1490 , n1510 );
xor ( n1512 , n1370 , n1372 );
xor ( n1513 , n1512 , n1375 );
and ( n1514 , n1510 , n1513 );
and ( n1515 , n1490 , n1513 );
or ( n1516 , n1511 , n1514 , n1515 );
xor ( n1517 , n1350 , n1378 );
xor ( n1518 , n1517 , n1381 );
and ( n1519 , n1516 , n1518 );
xor ( n1520 , n1426 , n1454 );
xor ( n1521 , n1520 , n1457 );
and ( n1522 , n1518 , n1521 );
and ( n1523 , n1516 , n1521 );
or ( n1524 , n1519 , n1522 , n1523 );
and ( n1525 , n1460 , n1524 );
xor ( n1526 , n1384 , n1386 );
xor ( n1527 , n1526 , n1389 );
and ( n1528 , n1524 , n1527 );
and ( n1529 , n1460 , n1527 );
or ( n1530 , n1525 , n1528 , n1529 );
and ( n1531 , n1402 , n1530 );
xor ( n1532 , n1402 , n1530 );
xor ( n1533 , n1460 , n1524 );
xor ( n1534 , n1533 , n1527 );
xor ( n1535 , n1181 , n1428 );
xor ( n1536 , n1428 , n1430 );
not ( n1537 , n1536 );
and ( n1538 , n1535 , n1537 );
and ( n1539 , n854 , n1538 );
not ( n1540 , n1539 );
xnor ( n1541 , n1540 , n1433 );
and ( n1542 , n1290 , n973 );
and ( n1543 , n1098 , n971 );
nor ( n1544 , n1542 , n1543 );
xnor ( n1545 , n1544 , n840 );
and ( n1546 , n1541 , n1545 );
and ( n1547 , n1413 , n851 );
and ( n1548 , n1308 , n849 );
nor ( n1549 , n1547 , n1548 );
xnor ( n1550 , n1549 , n859 );
and ( n1551 , n1545 , n1550 );
and ( n1552 , n1541 , n1550 );
or ( n1553 , n1546 , n1551 , n1552 );
and ( n1554 , n863 , n1298 );
and ( n1555 , n843 , n1296 );
nor ( n1556 , n1554 , n1555 );
xnor ( n1557 , n1556 , n1184 );
buf ( n1558 , n1557 );
and ( n1559 , n1553 , n1558 );
xor ( n1560 , n1406 , n1410 );
xor ( n1561 , n1560 , n1414 );
and ( n1562 , n1558 , n1561 );
and ( n1563 , n1553 , n1561 );
or ( n1564 , n1559 , n1562 , n1563 );
not ( n1565 , n1557 );
and ( n1566 , n1083 , n1106 );
and ( n1567 , n984 , n1104 );
nor ( n1568 , n1566 , n1567 );
xnor ( n1569 , n1568 , n1075 );
and ( n1570 , n1565 , n1569 );
buf ( n1571 , n553 );
buf ( n1572 , n1571 );
and ( n1573 , n1572 , n845 );
and ( n1574 , n1569 , n1573 );
and ( n1575 , n1565 , n1573 );
or ( n1576 , n1570 , n1574 , n1575 );
xor ( n1577 , n1434 , n1438 );
xor ( n1578 , n1577 , n1443 );
and ( n1579 , n1576 , n1578 );
xor ( n1580 , n1553 , n1558 );
xor ( n1581 , n1580 , n1561 );
and ( n1582 , n1578 , n1581 );
and ( n1583 , n1576 , n1581 );
or ( n1584 , n1579 , n1582 , n1583 );
and ( n1585 , n1564 , n1584 );
xor ( n1586 , n1446 , n1448 );
xor ( n1587 , n1586 , n1451 );
and ( n1588 , n1584 , n1587 );
and ( n1589 , n1564 , n1587 );
or ( n1590 , n1585 , n1588 , n1589 );
buf ( n1591 , n571 );
buf ( n1592 , n1591 );
buf ( n1593 , n572 );
buf ( n1594 , n1593 );
and ( n1595 , n1592 , n1594 );
not ( n1596 , n1595 );
and ( n1597 , n1430 , n1596 );
not ( n1598 , n1597 );
and ( n1599 , n843 , n1538 );
and ( n1600 , n854 , n1536 );
nor ( n1601 , n1599 , n1600 );
xnor ( n1602 , n1601 , n1433 );
and ( n1603 , n1598 , n1602 );
and ( n1604 , n1098 , n1106 );
and ( n1605 , n1083 , n1104 );
nor ( n1606 , n1604 , n1605 );
xnor ( n1607 , n1606 , n1075 );
and ( n1608 , n1602 , n1607 );
and ( n1609 , n1598 , n1607 );
or ( n1610 , n1603 , n1608 , n1609 );
and ( n1611 , n984 , n1298 );
and ( n1612 , n863 , n1296 );
nor ( n1613 , n1611 , n1612 );
xnor ( n1614 , n1613 , n1184 );
and ( n1615 , n1308 , n973 );
and ( n1616 , n1290 , n971 );
nor ( n1617 , n1615 , n1616 );
xnor ( n1618 , n1617 , n840 );
and ( n1619 , n1614 , n1618 );
and ( n1620 , n1572 , n851 );
and ( n1621 , n1413 , n849 );
nor ( n1622 , n1620 , n1621 );
xnor ( n1623 , n1622 , n859 );
and ( n1624 , n1618 , n1623 );
and ( n1625 , n1614 , n1623 );
or ( n1626 , n1619 , n1624 , n1625 );
and ( n1627 , n1610 , n1626 );
xor ( n1628 , n1541 , n1545 );
xor ( n1629 , n1628 , n1550 );
and ( n1630 , n1626 , n1629 );
and ( n1631 , n1610 , n1629 );
or ( n1632 , n1627 , n1630 , n1631 );
and ( n1633 , n863 , n1538 );
and ( n1634 , n843 , n1536 );
nor ( n1635 , n1633 , n1634 );
xnor ( n1636 , n1635 , n1433 );
and ( n1637 , n1290 , n1106 );
and ( n1638 , n1098 , n1104 );
nor ( n1639 , n1637 , n1638 );
xnor ( n1640 , n1639 , n1075 );
and ( n1641 , n1636 , n1640 );
and ( n1642 , n1413 , n973 );
and ( n1643 , n1308 , n971 );
nor ( n1644 , n1642 , n1643 );
xnor ( n1645 , n1644 , n840 );
and ( n1646 , n1640 , n1645 );
and ( n1647 , n1636 , n1645 );
or ( n1648 , n1641 , n1646 , n1647 );
xor ( n1649 , n1430 , n1592 );
xor ( n1650 , n1592 , n1594 );
not ( n1651 , n1650 );
and ( n1652 , n1649 , n1651 );
and ( n1653 , n854 , n1652 );
not ( n1654 , n1653 );
xnor ( n1655 , n1654 , n1597 );
buf ( n1656 , n1655 );
and ( n1657 , n1648 , n1656 );
buf ( n1658 , n554 );
buf ( n1659 , n1658 );
and ( n1660 , n1659 , n845 );
and ( n1661 , n1656 , n1660 );
and ( n1662 , n1648 , n1660 );
or ( n1663 , n1657 , n1661 , n1662 );
and ( n1664 , n1083 , n1298 );
and ( n1665 , n984 , n1296 );
nor ( n1666 , n1664 , n1665 );
xnor ( n1667 , n1666 , n1184 );
and ( n1668 , n1659 , n851 );
and ( n1669 , n1572 , n849 );
nor ( n1670 , n1668 , n1669 );
xnor ( n1671 , n1670 , n859 );
and ( n1672 , n1667 , n1671 );
buf ( n1673 , n555 );
buf ( n1674 , n1673 );
and ( n1675 , n1674 , n845 );
and ( n1676 , n1671 , n1675 );
and ( n1677 , n1667 , n1675 );
or ( n1678 , n1672 , n1676 , n1677 );
xor ( n1679 , n1598 , n1602 );
xor ( n1680 , n1679 , n1607 );
and ( n1681 , n1678 , n1680 );
xor ( n1682 , n1614 , n1618 );
xor ( n1683 , n1682 , n1623 );
and ( n1684 , n1680 , n1683 );
and ( n1685 , n1678 , n1683 );
or ( n1686 , n1681 , n1684 , n1685 );
and ( n1687 , n1663 , n1686 );
xor ( n1688 , n1565 , n1569 );
xor ( n1689 , n1688 , n1573 );
and ( n1690 , n1686 , n1689 );
and ( n1691 , n1663 , n1689 );
or ( n1692 , n1687 , n1690 , n1691 );
and ( n1693 , n1632 , n1692 );
xor ( n1694 , n1576 , n1578 );
xor ( n1695 , n1694 , n1581 );
and ( n1696 , n1692 , n1695 );
and ( n1697 , n1632 , n1695 );
or ( n1698 , n1693 , n1696 , n1697 );
buf ( n1699 , n587 );
buf ( n1700 , n1699 );
buf ( n1701 , n588 );
buf ( n1702 , n1701 );
and ( n1703 , n1700 , n1702 );
not ( n1704 , n1703 );
and ( n1705 , n1354 , n1704 );
not ( n1706 , n1705 );
and ( n1707 , n908 , n1464 );
and ( n1708 , n878 , n1462 );
nor ( n1709 , n1707 , n1708 );
xnor ( n1710 , n1709 , n1357 );
and ( n1711 , n1706 , n1710 );
and ( n1712 , n1025 , n1033 );
and ( n1713 , n1010 , n1031 );
nor ( n1714 , n1712 , n1713 );
xnor ( n1715 , n1714 , n1002 );
and ( n1716 , n1710 , n1715 );
and ( n1717 , n1706 , n1715 );
or ( n1718 , n1711 , n1716 , n1717 );
and ( n1719 , n917 , n1232 );
and ( n1720 , n897 , n1230 );
nor ( n1721 , n1719 , n1720 );
xnor ( n1722 , n1721 , n1131 );
and ( n1723 , n1242 , n888 );
and ( n1724 , n1224 , n886 );
nor ( n1725 , n1723 , n1724 );
xnor ( n1726 , n1725 , n893 );
and ( n1727 , n1722 , n1726 );
and ( n1728 , n1498 , n905 );
and ( n1729 , n1337 , n903 );
nor ( n1730 , n1728 , n1729 );
xnor ( n1731 , n1730 , n913 );
and ( n1732 , n1726 , n1731 );
and ( n1733 , n1722 , n1731 );
or ( n1734 , n1727 , n1732 , n1733 );
and ( n1735 , n1718 , n1734 );
xor ( n1736 , n1467 , n1471 );
xor ( n1737 , n1736 , n1476 );
and ( n1738 , n1734 , n1737 );
and ( n1739 , n1718 , n1737 );
or ( n1740 , n1735 , n1738 , n1739 );
and ( n1741 , n897 , n1464 );
and ( n1742 , n908 , n1462 );
nor ( n1743 , n1741 , n1742 );
xnor ( n1744 , n1743 , n1357 );
and ( n1745 , n1224 , n1033 );
and ( n1746 , n1025 , n1031 );
nor ( n1747 , n1745 , n1746 );
xnor ( n1748 , n1747 , n1002 );
and ( n1749 , n1744 , n1748 );
and ( n1750 , n1337 , n888 );
and ( n1751 , n1242 , n886 );
nor ( n1752 , n1750 , n1751 );
xnor ( n1753 , n1752 , n893 );
and ( n1754 , n1748 , n1753 );
and ( n1755 , n1744 , n1753 );
or ( n1756 , n1749 , n1754 , n1755 );
xor ( n1757 , n1354 , n1700 );
xor ( n1758 , n1700 , n1702 );
not ( n1759 , n1758 );
and ( n1760 , n1757 , n1759 );
and ( n1761 , n878 , n1760 );
not ( n1762 , n1761 );
xnor ( n1763 , n1762 , n1705 );
buf ( n1764 , n1763 );
and ( n1765 , n1756 , n1764 );
buf ( n1766 , n554 );
buf ( n1767 , n1766 );
and ( n1768 , n1767 , n899 );
and ( n1769 , n1764 , n1768 );
and ( n1770 , n1756 , n1768 );
or ( n1771 , n1765 , n1769 , n1770 );
and ( n1772 , n1010 , n1232 );
and ( n1773 , n917 , n1230 );
nor ( n1774 , n1772 , n1773 );
xnor ( n1775 , n1774 , n1131 );
and ( n1776 , n1767 , n905 );
and ( n1777 , n1498 , n903 );
nor ( n1778 , n1776 , n1777 );
xnor ( n1779 , n1778 , n913 );
and ( n1780 , n1775 , n1779 );
buf ( n1781 , n555 );
buf ( n1782 , n1781 );
and ( n1783 , n1782 , n899 );
and ( n1784 , n1779 , n1783 );
and ( n1785 , n1775 , n1783 );
or ( n1786 , n1780 , n1784 , n1785 );
xor ( n1787 , n1706 , n1710 );
xor ( n1788 , n1787 , n1715 );
and ( n1789 , n1786 , n1788 );
xor ( n1790 , n1722 , n1726 );
xor ( n1791 , n1790 , n1731 );
and ( n1792 , n1788 , n1791 );
and ( n1793 , n1786 , n1791 );
or ( n1794 , n1789 , n1792 , n1793 );
and ( n1795 , n1771 , n1794 );
xor ( n1796 , n1491 , n1495 );
xor ( n1797 , n1796 , n1499 );
and ( n1798 , n1794 , n1797 );
and ( n1799 , n1771 , n1797 );
or ( n1800 , n1795 , n1798 , n1799 );
and ( n1801 , n1740 , n1800 );
xor ( n1802 , n1502 , n1504 );
xor ( n1803 , n1802 , n1507 );
and ( n1804 , n1800 , n1803 );
and ( n1805 , n1740 , n1803 );
or ( n1806 , n1801 , n1804 , n1805 );
and ( n1807 , n1698 , n1806 );
xor ( n1808 , n1490 , n1510 );
xor ( n1809 , n1808 , n1513 );
and ( n1810 , n1806 , n1809 );
and ( n1811 , n1698 , n1809 );
or ( n1812 , n1807 , n1810 , n1811 );
and ( n1813 , n1590 , n1812 );
xor ( n1814 , n1516 , n1518 );
xor ( n1815 , n1814 , n1521 );
and ( n1816 , n1812 , n1815 );
and ( n1817 , n1590 , n1815 );
or ( n1818 , n1813 , n1816 , n1817 );
and ( n1819 , n1534 , n1818 );
xor ( n1820 , n1534 , n1818 );
xor ( n1821 , n1590 , n1812 );
xor ( n1822 , n1821 , n1815 );
and ( n1823 , n984 , n1538 );
and ( n1824 , n863 , n1536 );
nor ( n1825 , n1823 , n1824 );
xnor ( n1826 , n1825 , n1433 );
and ( n1827 , n1308 , n1106 );
and ( n1828 , n1290 , n1104 );
nor ( n1829 , n1827 , n1828 );
xnor ( n1830 , n1829 , n1075 );
and ( n1831 , n1826 , n1830 );
buf ( n1832 , n556 );
buf ( n1833 , n1832 );
and ( n1834 , n1833 , n845 );
and ( n1835 , n1830 , n1834 );
and ( n1836 , n1826 , n1834 );
or ( n1837 , n1831 , n1835 , n1836 );
buf ( n1838 , n573 );
buf ( n1839 , n1838 );
buf ( n1840 , n574 );
buf ( n1841 , n1840 );
and ( n1842 , n1839 , n1841 );
not ( n1843 , n1842 );
and ( n1844 , n1594 , n1843 );
not ( n1845 , n1844 );
and ( n1846 , n843 , n1652 );
and ( n1847 , n854 , n1650 );
nor ( n1848 , n1846 , n1847 );
xnor ( n1849 , n1848 , n1597 );
and ( n1850 , n1845 , n1849 );
and ( n1851 , n1098 , n1298 );
and ( n1852 , n1083 , n1296 );
nor ( n1853 , n1851 , n1852 );
xnor ( n1854 , n1853 , n1184 );
and ( n1855 , n1849 , n1854 );
and ( n1856 , n1845 , n1854 );
or ( n1857 , n1850 , n1855 , n1856 );
and ( n1858 , n1837 , n1857 );
not ( n1859 , n1655 );
and ( n1860 , n1857 , n1859 );
and ( n1861 , n1837 , n1859 );
or ( n1862 , n1858 , n1860 , n1861 );
xor ( n1863 , n1594 , n1839 );
xor ( n1864 , n1839 , n1841 );
not ( n1865 , n1864 );
and ( n1866 , n1863 , n1865 );
and ( n1867 , n854 , n1866 );
not ( n1868 , n1867 );
xnor ( n1869 , n1868 , n1844 );
buf ( n1870 , n1869 );
and ( n1871 , n1572 , n973 );
and ( n1872 , n1413 , n971 );
nor ( n1873 , n1871 , n1872 );
xnor ( n1874 , n1873 , n840 );
and ( n1875 , n1870 , n1874 );
and ( n1876 , n1674 , n851 );
and ( n1877 , n1659 , n849 );
nor ( n1878 , n1876 , n1877 );
xnor ( n1879 , n1878 , n859 );
and ( n1880 , n1874 , n1879 );
and ( n1881 , n1870 , n1879 );
or ( n1882 , n1875 , n1880 , n1881 );
xor ( n1883 , n1667 , n1671 );
xor ( n1884 , n1883 , n1675 );
and ( n1885 , n1882 , n1884 );
xor ( n1886 , n1636 , n1640 );
xor ( n1887 , n1886 , n1645 );
and ( n1888 , n1884 , n1887 );
and ( n1889 , n1882 , n1887 );
or ( n1890 , n1885 , n1888 , n1889 );
and ( n1891 , n1862 , n1890 );
xor ( n1892 , n1648 , n1656 );
xor ( n1893 , n1892 , n1660 );
and ( n1894 , n1890 , n1893 );
and ( n1895 , n1862 , n1893 );
or ( n1896 , n1891 , n1894 , n1895 );
xor ( n1897 , n1610 , n1626 );
xor ( n1898 , n1897 , n1629 );
and ( n1899 , n1896 , n1898 );
xor ( n1900 , n1663 , n1686 );
xor ( n1901 , n1900 , n1689 );
and ( n1902 , n1898 , n1901 );
and ( n1903 , n1896 , n1901 );
or ( n1904 , n1899 , n1902 , n1903 );
and ( n1905 , n917 , n1464 );
and ( n1906 , n897 , n1462 );
nor ( n1907 , n1905 , n1906 );
xnor ( n1908 , n1907 , n1357 );
and ( n1909 , n1242 , n1033 );
and ( n1910 , n1224 , n1031 );
nor ( n1911 , n1909 , n1910 );
xnor ( n1912 , n1911 , n1002 );
and ( n1913 , n1908 , n1912 );
buf ( n1914 , n556 );
buf ( n1915 , n1914 );
and ( n1916 , n1915 , n899 );
and ( n1917 , n1912 , n1916 );
and ( n1918 , n1908 , n1916 );
or ( n1919 , n1913 , n1917 , n1918 );
buf ( n1920 , n589 );
buf ( n1921 , n1920 );
buf ( n1922 , n590 );
buf ( n1923 , n1922 );
and ( n1924 , n1921 , n1923 );
not ( n1925 , n1924 );
and ( n1926 , n1702 , n1925 );
not ( n1927 , n1926 );
and ( n1928 , n908 , n1760 );
and ( n1929 , n878 , n1758 );
nor ( n1930 , n1928 , n1929 );
xnor ( n1931 , n1930 , n1705 );
and ( n1932 , n1927 , n1931 );
and ( n1933 , n1025 , n1232 );
and ( n1934 , n1010 , n1230 );
nor ( n1935 , n1933 , n1934 );
xnor ( n1936 , n1935 , n1131 );
and ( n1937 , n1931 , n1936 );
and ( n1938 , n1927 , n1936 );
or ( n1939 , n1932 , n1937 , n1938 );
and ( n1940 , n1919 , n1939 );
not ( n1941 , n1763 );
and ( n1942 , n1939 , n1941 );
and ( n1943 , n1919 , n1941 );
or ( n1944 , n1940 , n1942 , n1943 );
xor ( n1945 , n1702 , n1921 );
xor ( n1946 , n1921 , n1923 );
not ( n1947 , n1946 );
and ( n1948 , n1945 , n1947 );
and ( n1949 , n878 , n1948 );
not ( n1950 , n1949 );
xnor ( n1951 , n1950 , n1926 );
buf ( n1952 , n1951 );
and ( n1953 , n1498 , n888 );
and ( n1954 , n1337 , n886 );
nor ( n1955 , n1953 , n1954 );
xnor ( n1956 , n1955 , n893 );
and ( n1957 , n1952 , n1956 );
and ( n1958 , n1782 , n905 );
and ( n1959 , n1767 , n903 );
nor ( n1960 , n1958 , n1959 );
xnor ( n1961 , n1960 , n913 );
and ( n1962 , n1956 , n1961 );
and ( n1963 , n1952 , n1961 );
or ( n1964 , n1957 , n1962 , n1963 );
xor ( n1965 , n1775 , n1779 );
xor ( n1966 , n1965 , n1783 );
and ( n1967 , n1964 , n1966 );
xor ( n1968 , n1744 , n1748 );
xor ( n1969 , n1968 , n1753 );
and ( n1970 , n1966 , n1969 );
and ( n1971 , n1964 , n1969 );
or ( n1972 , n1967 , n1970 , n1971 );
and ( n1973 , n1944 , n1972 );
xor ( n1974 , n1756 , n1764 );
xor ( n1975 , n1974 , n1768 );
and ( n1976 , n1972 , n1975 );
and ( n1977 , n1944 , n1975 );
or ( n1978 , n1973 , n1976 , n1977 );
xor ( n1979 , n1718 , n1734 );
xor ( n1980 , n1979 , n1737 );
and ( n1981 , n1978 , n1980 );
xor ( n1982 , n1771 , n1794 );
xor ( n1983 , n1982 , n1797 );
and ( n1984 , n1980 , n1983 );
and ( n1985 , n1978 , n1983 );
or ( n1986 , n1981 , n1984 , n1985 );
and ( n1987 , n1904 , n1986 );
xor ( n1988 , n1740 , n1800 );
xor ( n1989 , n1988 , n1803 );
and ( n1990 , n1986 , n1989 );
and ( n1991 , n1904 , n1989 );
or ( n1992 , n1987 , n1990 , n1991 );
xor ( n1993 , n1564 , n1584 );
xor ( n1994 , n1993 , n1587 );
and ( n1995 , n1992 , n1994 );
xor ( n1996 , n1698 , n1806 );
xor ( n1997 , n1996 , n1809 );
and ( n1998 , n1994 , n1997 );
and ( n1999 , n1992 , n1997 );
or ( n2000 , n1995 , n1998 , n1999 );
and ( n2001 , n1822 , n2000 );
xor ( n2002 , n1822 , n2000 );
xor ( n2003 , n1992 , n1994 );
xor ( n2004 , n2003 , n1997 );
and ( n2005 , n863 , n1652 );
and ( n2006 , n843 , n1650 );
nor ( n2007 , n2005 , n2006 );
xnor ( n2008 , n2007 , n1597 );
and ( n2009 , n1290 , n1298 );
and ( n2010 , n1098 , n1296 );
nor ( n2011 , n2009 , n2010 );
xnor ( n2012 , n2011 , n1184 );
and ( n2013 , n2008 , n2012 );
buf ( n2014 , n557 );
buf ( n2015 , n2014 );
and ( n2016 , n2015 , n845 );
and ( n2017 , n2012 , n2016 );
and ( n2018 , n2008 , n2016 );
or ( n2019 , n2013 , n2017 , n2018 );
and ( n2020 , n1083 , n1538 );
and ( n2021 , n984 , n1536 );
nor ( n2022 , n2020 , n2021 );
xnor ( n2023 , n2022 , n1433 );
and ( n2024 , n1413 , n1106 );
and ( n2025 , n1308 , n1104 );
nor ( n2026 , n2024 , n2025 );
xnor ( n2027 , n2026 , n1075 );
and ( n2028 , n2023 , n2027 );
and ( n2029 , n1659 , n973 );
and ( n2030 , n1572 , n971 );
nor ( n2031 , n2029 , n2030 );
xnor ( n2032 , n2031 , n840 );
and ( n2033 , n2027 , n2032 );
and ( n2034 , n2023 , n2032 );
or ( n2035 , n2028 , n2033 , n2034 );
and ( n2036 , n2019 , n2035 );
xor ( n2037 , n1845 , n1849 );
xor ( n2038 , n2037 , n1854 );
and ( n2039 , n2035 , n2038 );
and ( n2040 , n2019 , n2038 );
or ( n2041 , n2036 , n2039 , n2040 );
xor ( n2042 , n1837 , n1857 );
xor ( n2043 , n2042 , n1859 );
and ( n2044 , n2041 , n2043 );
xor ( n2045 , n1882 , n1884 );
xor ( n2046 , n2045 , n1887 );
and ( n2047 , n2043 , n2046 );
and ( n2048 , n2041 , n2046 );
or ( n2049 , n2044 , n2047 , n2048 );
xor ( n2050 , n1678 , n1680 );
xor ( n2051 , n2050 , n1683 );
and ( n2052 , n2049 , n2051 );
xor ( n2053 , n1862 , n1890 );
xor ( n2054 , n2053 , n1893 );
and ( n2055 , n2051 , n2054 );
and ( n2056 , n2049 , n2054 );
or ( n2057 , n2052 , n2055 , n2056 );
and ( n2058 , n897 , n1760 );
and ( n2059 , n908 , n1758 );
nor ( n2060 , n2058 , n2059 );
xnor ( n2061 , n2060 , n1705 );
and ( n2062 , n1224 , n1232 );
and ( n2063 , n1025 , n1230 );
nor ( n2064 , n2062 , n2063 );
xnor ( n2065 , n2064 , n1131 );
and ( n2066 , n2061 , n2065 );
buf ( n2067 , n557 );
buf ( n2068 , n2067 );
and ( n2069 , n2068 , n899 );
and ( n2070 , n2065 , n2069 );
and ( n2071 , n2061 , n2069 );
or ( n2072 , n2066 , n2070 , n2071 );
and ( n2073 , n1010 , n1464 );
and ( n2074 , n917 , n1462 );
nor ( n2075 , n2073 , n2074 );
xnor ( n2076 , n2075 , n1357 );
and ( n2077 , n1337 , n1033 );
and ( n2078 , n1242 , n1031 );
nor ( n2079 , n2077 , n2078 );
xnor ( n2080 , n2079 , n1002 );
and ( n2081 , n2076 , n2080 );
and ( n2082 , n1767 , n888 );
and ( n2083 , n1498 , n886 );
nor ( n2084 , n2082 , n2083 );
xnor ( n2085 , n2084 , n893 );
and ( n2086 , n2080 , n2085 );
and ( n2087 , n2076 , n2085 );
or ( n2088 , n2081 , n2086 , n2087 );
and ( n2089 , n2072 , n2088 );
xor ( n2090 , n1927 , n1931 );
xor ( n2091 , n2090 , n1936 );
and ( n2092 , n2088 , n2091 );
and ( n2093 , n2072 , n2091 );
or ( n2094 , n2089 , n2092 , n2093 );
xor ( n2095 , n1919 , n1939 );
xor ( n2096 , n2095 , n1941 );
and ( n2097 , n2094 , n2096 );
xor ( n2098 , n1964 , n1966 );
xor ( n2099 , n2098 , n1969 );
and ( n2100 , n2096 , n2099 );
and ( n2101 , n2094 , n2099 );
or ( n2102 , n2097 , n2100 , n2101 );
xor ( n2103 , n1786 , n1788 );
xor ( n2104 , n2103 , n1791 );
and ( n2105 , n2102 , n2104 );
xor ( n2106 , n1944 , n1972 );
xor ( n2107 , n2106 , n1975 );
and ( n2108 , n2104 , n2107 );
and ( n2109 , n2102 , n2107 );
or ( n2110 , n2105 , n2108 , n2109 );
and ( n2111 , n2057 , n2110 );
xor ( n2112 , n1978 , n1980 );
xor ( n2113 , n2112 , n1983 );
and ( n2114 , n2110 , n2113 );
and ( n2115 , n2057 , n2113 );
or ( n2116 , n2111 , n2114 , n2115 );
xor ( n2117 , n1632 , n1692 );
xor ( n2118 , n2117 , n1695 );
and ( n2119 , n2116 , n2118 );
xor ( n2120 , n1904 , n1986 );
xor ( n2121 , n2120 , n1989 );
and ( n2122 , n2118 , n2121 );
and ( n2123 , n2116 , n2121 );
or ( n2124 , n2119 , n2122 , n2123 );
and ( n2125 , n2004 , n2124 );
xor ( n2126 , n2004 , n2124 );
xor ( n2127 , n2116 , n2118 );
xor ( n2128 , n2127 , n2121 );
and ( n2129 , n1098 , n1538 );
and ( n2130 , n1083 , n1536 );
nor ( n2131 , n2129 , n2130 );
xnor ( n2132 , n2131 , n1433 );
buf ( n2133 , n2132 );
not ( n2134 , n1869 );
and ( n2135 , n2133 , n2134 );
and ( n2136 , n1833 , n851 );
and ( n2137 , n1674 , n849 );
nor ( n2138 , n2136 , n2137 );
xnor ( n2139 , n2138 , n859 );
and ( n2140 , n2134 , n2139 );
and ( n2141 , n2133 , n2139 );
or ( n2142 , n2135 , n2140 , n2141 );
xor ( n2143 , n1826 , n1830 );
xor ( n2144 , n2143 , n1834 );
and ( n2145 , n2142 , n2144 );
xor ( n2146 , n1870 , n1874 );
xor ( n2147 , n2146 , n1879 );
and ( n2148 , n2144 , n2147 );
and ( n2149 , n2142 , n2147 );
or ( n2150 , n2145 , n2148 , n2149 );
not ( n2151 , n1841 );
and ( n2152 , n2015 , n851 );
and ( n2153 , n1833 , n849 );
nor ( n2154 , n2152 , n2153 );
xnor ( n2155 , n2154 , n859 );
and ( n2156 , n2151 , n2155 );
buf ( n2157 , n558 );
buf ( n2158 , n2157 );
and ( n2159 , n2158 , n845 );
and ( n2160 , n2155 , n2159 );
and ( n2161 , n2151 , n2159 );
or ( n2162 , n2156 , n2160 , n2161 );
and ( n2163 , n843 , n1866 );
and ( n2164 , n854 , n1864 );
nor ( n2165 , n2163 , n2164 );
xnor ( n2166 , n2165 , n1844 );
and ( n2167 , n984 , n1652 );
and ( n2168 , n863 , n1650 );
nor ( n2169 , n2167 , n2168 );
xnor ( n2170 , n2169 , n1597 );
and ( n2171 , n2166 , n2170 );
and ( n2172 , n1308 , n1298 );
and ( n2173 , n1290 , n1296 );
nor ( n2174 , n2172 , n2173 );
xnor ( n2175 , n2174 , n1184 );
and ( n2176 , n2170 , n2175 );
and ( n2177 , n2166 , n2175 );
or ( n2178 , n2171 , n2176 , n2177 );
and ( n2179 , n2162 , n2178 );
xor ( n2180 , n2023 , n2027 );
xor ( n2181 , n2180 , n2032 );
and ( n2182 , n2178 , n2181 );
and ( n2183 , n2162 , n2181 );
or ( n2184 , n2179 , n2182 , n2183 );
buf ( n2185 , n575 );
buf ( n2186 , n2185 );
xor ( n2187 , n1841 , n2186 );
not ( n2188 , n2186 );
and ( n2189 , n2187 , n2188 );
and ( n2190 , n854 , n2189 );
not ( n2191 , n2190 );
xnor ( n2192 , n2191 , n1841 );
and ( n2193 , n863 , n1866 );
and ( n2194 , n843 , n1864 );
nor ( n2195 , n2193 , n2194 );
xnor ( n2196 , n2195 , n1844 );
and ( n2197 , n2192 , n2196 );
buf ( n2198 , n559 );
buf ( n2199 , n2198 );
and ( n2200 , n2199 , n845 );
and ( n2201 , n2196 , n2200 );
and ( n2202 , n2192 , n2200 );
or ( n2203 , n2197 , n2201 , n2202 );
and ( n2204 , n1083 , n1652 );
and ( n2205 , n984 , n1650 );
nor ( n2206 , n2204 , n2205 );
xnor ( n2207 , n2206 , n1597 );
and ( n2208 , n1659 , n1106 );
and ( n2209 , n1572 , n1104 );
nor ( n2210 , n2208 , n2209 );
xnor ( n2211 , n2210 , n1075 );
and ( n2212 , n2207 , n2211 );
and ( n2213 , n1833 , n973 );
and ( n2214 , n1674 , n971 );
nor ( n2215 , n2213 , n2214 );
xnor ( n2216 , n2215 , n840 );
and ( n2217 , n2211 , n2216 );
and ( n2218 , n2207 , n2216 );
or ( n2219 , n2212 , n2217 , n2218 );
and ( n2220 , n2203 , n2219 );
and ( n2221 , n1290 , n1538 );
and ( n2222 , n1098 , n1536 );
nor ( n2223 , n2221 , n2222 );
xnor ( n2224 , n2223 , n1433 );
and ( n2225 , n1413 , n1298 );
and ( n2226 , n1308 , n1296 );
nor ( n2227 , n2225 , n2226 );
xnor ( n2228 , n2227 , n1184 );
and ( n2229 , n2224 , n2228 );
and ( n2230 , n2158 , n851 );
and ( n2231 , n2015 , n849 );
nor ( n2232 , n2230 , n2231 );
xnor ( n2233 , n2232 , n859 );
and ( n2234 , n2228 , n2233 );
and ( n2235 , n2224 , n2233 );
or ( n2236 , n2229 , n2234 , n2235 );
and ( n2237 , n2219 , n2236 );
and ( n2238 , n2203 , n2236 );
or ( n2239 , n2220 , n2237 , n2238 );
xor ( n2240 , n2008 , n2012 );
xor ( n2241 , n2240 , n2016 );
and ( n2242 , n2239 , n2241 );
xor ( n2243 , n2133 , n2134 );
xor ( n2244 , n2243 , n2139 );
and ( n2245 , n2241 , n2244 );
and ( n2246 , n2239 , n2244 );
or ( n2247 , n2242 , n2245 , n2246 );
and ( n2248 , n2184 , n2247 );
xor ( n2249 , n2019 , n2035 );
xor ( n2250 , n2249 , n2038 );
and ( n2251 , n2247 , n2250 );
and ( n2252 , n2184 , n2250 );
or ( n2253 , n2248 , n2251 , n2252 );
and ( n2254 , n2150 , n2253 );
xor ( n2255 , n2041 , n2043 );
xor ( n2256 , n2255 , n2046 );
and ( n2257 , n2253 , n2256 );
and ( n2258 , n2150 , n2256 );
or ( n2259 , n2254 , n2257 , n2258 );
and ( n2260 , n1025 , n1464 );
and ( n2261 , n1010 , n1462 );
nor ( n2262 , n2260 , n2261 );
xnor ( n2263 , n2262 , n1357 );
buf ( n2264 , n2263 );
not ( n2265 , n1951 );
and ( n2266 , n2264 , n2265 );
and ( n2267 , n1915 , n905 );
and ( n2268 , n1782 , n903 );
nor ( n2269 , n2267 , n2268 );
xnor ( n2270 , n2269 , n913 );
and ( n2271 , n2265 , n2270 );
and ( n2272 , n2264 , n2270 );
or ( n2273 , n2266 , n2271 , n2272 );
xor ( n2274 , n1908 , n1912 );
xor ( n2275 , n2274 , n1916 );
and ( n2276 , n2273 , n2275 );
xor ( n2277 , n1952 , n1956 );
xor ( n2278 , n2277 , n1961 );
and ( n2279 , n2275 , n2278 );
and ( n2280 , n2273 , n2278 );
or ( n2281 , n2276 , n2279 , n2280 );
not ( n2282 , n1923 );
and ( n2283 , n2068 , n905 );
and ( n2284 , n1915 , n903 );
nor ( n2285 , n2283 , n2284 );
xnor ( n2286 , n2285 , n913 );
and ( n2287 , n2282 , n2286 );
buf ( n2288 , n558 );
buf ( n2289 , n2288 );
and ( n2290 , n2289 , n899 );
and ( n2291 , n2286 , n2290 );
and ( n2292 , n2282 , n2290 );
or ( n2293 , n2287 , n2291 , n2292 );
and ( n2294 , n908 , n1948 );
and ( n2295 , n878 , n1946 );
nor ( n2296 , n2294 , n2295 );
xnor ( n2297 , n2296 , n1926 );
and ( n2298 , n917 , n1760 );
and ( n2299 , n897 , n1758 );
nor ( n2300 , n2298 , n2299 );
xnor ( n2301 , n2300 , n1705 );
and ( n2302 , n2297 , n2301 );
and ( n2303 , n1242 , n1232 );
and ( n2304 , n1224 , n1230 );
nor ( n2305 , n2303 , n2304 );
xnor ( n2306 , n2305 , n1131 );
and ( n2307 , n2301 , n2306 );
and ( n2308 , n2297 , n2306 );
or ( n2309 , n2302 , n2307 , n2308 );
and ( n2310 , n2293 , n2309 );
xor ( n2311 , n2076 , n2080 );
xor ( n2312 , n2311 , n2085 );
and ( n2313 , n2309 , n2312 );
and ( n2314 , n2293 , n2312 );
or ( n2315 , n2310 , n2313 , n2314 );
and ( n2316 , n1010 , n1760 );
and ( n2317 , n917 , n1758 );
nor ( n2318 , n2316 , n2317 );
xnor ( n2319 , n2318 , n1705 );
and ( n2320 , n1767 , n1033 );
and ( n2321 , n1498 , n1031 );
nor ( n2322 , n2320 , n2321 );
xnor ( n2323 , n2322 , n1002 );
and ( n2324 , n2319 , n2323 );
and ( n2325 , n1915 , n888 );
and ( n2326 , n1782 , n886 );
nor ( n2327 , n2325 , n2326 );
xnor ( n2328 , n2327 , n893 );
and ( n2329 , n2323 , n2328 );
and ( n2330 , n2319 , n2328 );
or ( n2331 , n2324 , n2329 , n2330 );
buf ( n2332 , n591 );
buf ( n2333 , n2332 );
xor ( n2334 , n1923 , n2333 );
not ( n2335 , n2333 );
and ( n2336 , n2334 , n2335 );
and ( n2337 , n878 , n2336 );
not ( n2338 , n2337 );
xnor ( n2339 , n2338 , n1923 );
and ( n2340 , n897 , n1948 );
and ( n2341 , n908 , n1946 );
nor ( n2342 , n2340 , n2341 );
xnor ( n2343 , n2342 , n1926 );
and ( n2344 , n2339 , n2343 );
buf ( n2345 , n559 );
buf ( n2346 , n2345 );
and ( n2347 , n2346 , n899 );
and ( n2348 , n2343 , n2347 );
and ( n2349 , n2339 , n2347 );
or ( n2350 , n2344 , n2348 , n2349 );
and ( n2351 , n2331 , n2350 );
and ( n2352 , n1224 , n1464 );
and ( n2353 , n1025 , n1462 );
nor ( n2354 , n2352 , n2353 );
xnor ( n2355 , n2354 , n1357 );
and ( n2356 , n1337 , n1232 );
and ( n2357 , n1242 , n1230 );
nor ( n2358 , n2356 , n2357 );
xnor ( n2359 , n2358 , n1131 );
and ( n2360 , n2355 , n2359 );
and ( n2361 , n2289 , n905 );
and ( n2362 , n2068 , n903 );
nor ( n2363 , n2361 , n2362 );
xnor ( n2364 , n2363 , n913 );
and ( n2365 , n2359 , n2364 );
and ( n2366 , n2355 , n2364 );
or ( n2367 , n2360 , n2365 , n2366 );
and ( n2368 , n2350 , n2367 );
and ( n2369 , n2331 , n2367 );
or ( n2370 , n2351 , n2368 , n2369 );
xor ( n2371 , n2061 , n2065 );
xor ( n2372 , n2371 , n2069 );
and ( n2373 , n2370 , n2372 );
xor ( n2374 , n2264 , n2265 );
xor ( n2375 , n2374 , n2270 );
and ( n2376 , n2372 , n2375 );
and ( n2377 , n2370 , n2375 );
or ( n2378 , n2373 , n2376 , n2377 );
and ( n2379 , n2315 , n2378 );
xor ( n2380 , n2072 , n2088 );
xor ( n2381 , n2380 , n2091 );
and ( n2382 , n2378 , n2381 );
and ( n2383 , n2315 , n2381 );
or ( n2384 , n2379 , n2382 , n2383 );
and ( n2385 , n2281 , n2384 );
xor ( n2386 , n2094 , n2096 );
xor ( n2387 , n2386 , n2099 );
and ( n2388 , n2384 , n2387 );
and ( n2389 , n2281 , n2387 );
or ( n2390 , n2385 , n2388 , n2389 );
and ( n2391 , n2259 , n2390 );
xor ( n2392 , n2102 , n2104 );
xor ( n2393 , n2392 , n2107 );
and ( n2394 , n2390 , n2393 );
and ( n2395 , n2259 , n2393 );
or ( n2396 , n2391 , n2394 , n2395 );
xor ( n2397 , n1896 , n1898 );
xor ( n2398 , n2397 , n1901 );
and ( n2399 , n2396 , n2398 );
xor ( n2400 , n2057 , n2110 );
xor ( n2401 , n2400 , n2113 );
and ( n2402 , n2398 , n2401 );
and ( n2403 , n2396 , n2401 );
or ( n2404 , n2399 , n2402 , n2403 );
and ( n2405 , n2128 , n2404 );
xor ( n2406 , n2128 , n2404 );
xor ( n2407 , n2396 , n2398 );
xor ( n2408 , n2407 , n2401 );
not ( n2409 , n2132 );
and ( n2410 , n1572 , n1106 );
and ( n2411 , n1413 , n1104 );
nor ( n2412 , n2410 , n2411 );
xnor ( n2413 , n2412 , n1075 );
and ( n2414 , n2409 , n2413 );
and ( n2415 , n1674 , n973 );
and ( n2416 , n1659 , n971 );
nor ( n2417 , n2415 , n2416 );
xnor ( n2418 , n2417 , n840 );
and ( n2419 , n2413 , n2418 );
and ( n2420 , n2409 , n2418 );
or ( n2421 , n2414 , n2419 , n2420 );
and ( n2422 , n1098 , n1652 );
and ( n2423 , n1083 , n1650 );
nor ( n2424 , n2422 , n2423 );
xnor ( n2425 , n2424 , n1597 );
and ( n2426 , n1572 , n1298 );
and ( n2427 , n1413 , n1296 );
nor ( n2428 , n2426 , n2427 );
xnor ( n2429 , n2428 , n1184 );
and ( n2430 , n2425 , n2429 );
and ( n2431 , n1674 , n1106 );
and ( n2432 , n1659 , n1104 );
nor ( n2433 , n2431 , n2432 );
xnor ( n2434 , n2433 , n1075 );
and ( n2435 , n2429 , n2434 );
and ( n2436 , n2425 , n2434 );
or ( n2437 , n2430 , n2435 , n2436 );
and ( n2438 , n984 , n1866 );
and ( n2439 , n863 , n1864 );
nor ( n2440 , n2438 , n2439 );
xnor ( n2441 , n2440 , n1844 );
and ( n2442 , n1308 , n1538 );
and ( n2443 , n1290 , n1536 );
nor ( n2444 , n2442 , n2443 );
xnor ( n2445 , n2444 , n1433 );
and ( n2446 , n2441 , n2445 );
and ( n2447 , n2199 , n851 );
and ( n2448 , n2158 , n849 );
nor ( n2449 , n2447 , n2448 );
xnor ( n2450 , n2449 , n859 );
and ( n2451 , n2445 , n2450 );
and ( n2452 , n2441 , n2450 );
or ( n2453 , n2446 , n2451 , n2452 );
and ( n2454 , n2437 , n2453 );
and ( n2455 , n843 , n2189 );
and ( n2456 , n854 , n2186 );
nor ( n2457 , n2455 , n2456 );
xnor ( n2458 , n2457 , n1841 );
and ( n2459 , n2199 , n849 );
not ( n2460 , n2459 );
and ( n2461 , n2460 , n859 );
and ( n2462 , n2458 , n2461 );
and ( n2463 , n2453 , n2462 );
and ( n2464 , n2437 , n2462 );
or ( n2465 , n2454 , n2463 , n2464 );
xor ( n2466 , n2151 , n2155 );
xor ( n2467 , n2466 , n2159 );
and ( n2468 , n2465 , n2467 );
xor ( n2469 , n2166 , n2170 );
xor ( n2470 , n2469 , n2175 );
and ( n2471 , n2467 , n2470 );
and ( n2472 , n2465 , n2470 );
or ( n2473 , n2468 , n2471 , n2472 );
and ( n2474 , n2421 , n2473 );
xor ( n2475 , n2162 , n2178 );
xor ( n2476 , n2475 , n2181 );
and ( n2477 , n2473 , n2476 );
and ( n2478 , n2421 , n2476 );
or ( n2479 , n2474 , n2477 , n2478 );
xor ( n2480 , n2142 , n2144 );
xor ( n2481 , n2480 , n2147 );
and ( n2482 , n2479 , n2481 );
xor ( n2483 , n2184 , n2247 );
xor ( n2484 , n2483 , n2250 );
and ( n2485 , n2481 , n2484 );
and ( n2486 , n2479 , n2484 );
or ( n2487 , n2482 , n2485 , n2486 );
not ( n2488 , n2263 );
and ( n2489 , n1498 , n1033 );
and ( n2490 , n1337 , n1031 );
nor ( n2491 , n2489 , n2490 );
xnor ( n2492 , n2491 , n1002 );
and ( n2493 , n2488 , n2492 );
and ( n2494 , n1782 , n888 );
and ( n2495 , n1767 , n886 );
nor ( n2496 , n2494 , n2495 );
xnor ( n2497 , n2496 , n893 );
and ( n2498 , n2492 , n2497 );
and ( n2499 , n2488 , n2497 );
or ( n2500 , n2493 , n2498 , n2499 );
and ( n2501 , n1025 , n1760 );
and ( n2502 , n1010 , n1758 );
nor ( n2503 , n2501 , n2502 );
xnor ( n2504 , n2503 , n1705 );
and ( n2505 , n1498 , n1232 );
and ( n2506 , n1337 , n1230 );
nor ( n2507 , n2505 , n2506 );
xnor ( n2508 , n2507 , n1131 );
and ( n2509 , n2504 , n2508 );
and ( n2510 , n1782 , n1033 );
and ( n2511 , n1767 , n1031 );
nor ( n2512 , n2510 , n2511 );
xnor ( n2513 , n2512 , n1002 );
and ( n2514 , n2508 , n2513 );
and ( n2515 , n2504 , n2513 );
or ( n2516 , n2509 , n2514 , n2515 );
and ( n2517 , n917 , n1948 );
and ( n2518 , n897 , n1946 );
nor ( n2519 , n2517 , n2518 );
xnor ( n2520 , n2519 , n1926 );
and ( n2521 , n1242 , n1464 );
and ( n2522 , n1224 , n1462 );
nor ( n2523 , n2521 , n2522 );
xnor ( n2524 , n2523 , n1357 );
and ( n2525 , n2520 , n2524 );
and ( n2526 , n2346 , n905 );
and ( n2527 , n2289 , n903 );
nor ( n2528 , n2526 , n2527 );
xnor ( n2529 , n2528 , n913 );
and ( n2530 , n2524 , n2529 );
and ( n2531 , n2520 , n2529 );
or ( n2532 , n2525 , n2530 , n2531 );
and ( n2533 , n2516 , n2532 );
and ( n2534 , n908 , n2336 );
and ( n2535 , n878 , n2333 );
nor ( n2536 , n2534 , n2535 );
xnor ( n2537 , n2536 , n1923 );
and ( n2538 , n2346 , n903 );
not ( n2539 , n2538 );
and ( n2540 , n2539 , n913 );
and ( n2541 , n2537 , n2540 );
and ( n2542 , n2532 , n2541 );
and ( n2543 , n2516 , n2541 );
or ( n2544 , n2533 , n2542 , n2543 );
xor ( n2545 , n2282 , n2286 );
xor ( n2546 , n2545 , n2290 );
and ( n2547 , n2544 , n2546 );
xor ( n2548 , n2297 , n2301 );
xor ( n2549 , n2548 , n2306 );
and ( n2550 , n2546 , n2549 );
and ( n2551 , n2544 , n2549 );
or ( n2552 , n2547 , n2550 , n2551 );
and ( n2553 , n2500 , n2552 );
xor ( n2554 , n2293 , n2309 );
xor ( n2555 , n2554 , n2312 );
and ( n2556 , n2552 , n2555 );
and ( n2557 , n2500 , n2555 );
or ( n2558 , n2553 , n2556 , n2557 );
xor ( n2559 , n2273 , n2275 );
xor ( n2560 , n2559 , n2278 );
and ( n2561 , n2558 , n2560 );
xor ( n2562 , n2315 , n2378 );
xor ( n2563 , n2562 , n2381 );
and ( n2564 , n2560 , n2563 );
and ( n2565 , n2558 , n2563 );
or ( n2566 , n2561 , n2564 , n2565 );
and ( n2567 , n2487 , n2566 );
xor ( n2568 , n2281 , n2384 );
xor ( n2569 , n2568 , n2387 );
and ( n2570 , n2566 , n2569 );
and ( n2571 , n2487 , n2569 );
or ( n2572 , n2567 , n2570 , n2571 );
xor ( n2573 , n2049 , n2051 );
xor ( n2574 , n2573 , n2054 );
and ( n2575 , n2572 , n2574 );
xor ( n2576 , n2259 , n2390 );
xor ( n2577 , n2576 , n2393 );
and ( n2578 , n2574 , n2577 );
and ( n2579 , n2572 , n2577 );
or ( n2580 , n2575 , n2578 , n2579 );
and ( n2581 , n2408 , n2580 );
xor ( n2582 , n2408 , n2580 );
xor ( n2583 , n2572 , n2574 );
xor ( n2584 , n2583 , n2577 );
xor ( n2585 , n2192 , n2196 );
xor ( n2586 , n2585 , n2200 );
xor ( n2587 , n2207 , n2211 );
xor ( n2588 , n2587 , n2216 );
and ( n2589 , n2586 , n2588 );
xor ( n2590 , n2224 , n2228 );
xor ( n2591 , n2590 , n2233 );
and ( n2592 , n2588 , n2591 );
and ( n2593 , n2586 , n2591 );
or ( n2594 , n2589 , n2592 , n2593 );
xor ( n2595 , n2203 , n2219 );
xor ( n2596 , n2595 , n2236 );
and ( n2597 , n2594 , n2596 );
xor ( n2598 , n2409 , n2413 );
xor ( n2599 , n2598 , n2418 );
and ( n2600 , n2596 , n2599 );
and ( n2601 , n2594 , n2599 );
or ( n2602 , n2597 , n2600 , n2601 );
xor ( n2603 , n2239 , n2241 );
xor ( n2604 , n2603 , n2244 );
and ( n2605 , n2602 , n2604 );
xor ( n2606 , n2421 , n2473 );
xor ( n2607 , n2606 , n2476 );
and ( n2608 , n2604 , n2607 );
and ( n2609 , n2602 , n2607 );
or ( n2610 , n2605 , n2608 , n2609 );
xor ( n2611 , n2319 , n2323 );
xor ( n2612 , n2611 , n2328 );
xor ( n2613 , n2339 , n2343 );
xor ( n2614 , n2613 , n2347 );
and ( n2615 , n2612 , n2614 );
xor ( n2616 , n2355 , n2359 );
xor ( n2617 , n2616 , n2364 );
and ( n2618 , n2614 , n2617 );
and ( n2619 , n2612 , n2617 );
or ( n2620 , n2615 , n2618 , n2619 );
xor ( n2621 , n2331 , n2350 );
xor ( n2622 , n2621 , n2367 );
and ( n2623 , n2620 , n2622 );
xor ( n2624 , n2488 , n2492 );
xor ( n2625 , n2624 , n2497 );
and ( n2626 , n2622 , n2625 );
and ( n2627 , n2620 , n2625 );
or ( n2628 , n2623 , n2626 , n2627 );
xor ( n2629 , n2370 , n2372 );
xor ( n2630 , n2629 , n2375 );
and ( n2631 , n2628 , n2630 );
xor ( n2632 , n2500 , n2552 );
xor ( n2633 , n2632 , n2555 );
and ( n2634 , n2630 , n2633 );
and ( n2635 , n2628 , n2633 );
or ( n2636 , n2631 , n2634 , n2635 );
and ( n2637 , n2610 , n2636 );
xor ( n2638 , n2558 , n2560 );
xor ( n2639 , n2638 , n2563 );
and ( n2640 , n2636 , n2639 );
and ( n2641 , n2610 , n2639 );
or ( n2642 , n2637 , n2640 , n2641 );
xor ( n2643 , n2150 , n2253 );
xor ( n2644 , n2643 , n2256 );
and ( n2645 , n2642 , n2644 );
xor ( n2646 , n2487 , n2566 );
xor ( n2647 , n2646 , n2569 );
and ( n2648 , n2644 , n2647 );
and ( n2649 , n2642 , n2647 );
or ( n2650 , n2645 , n2648 , n2649 );
and ( n2651 , n2584 , n2650 );
xor ( n2652 , n2584 , n2650 );
xor ( n2653 , n2458 , n2461 );
and ( n2654 , n863 , n2189 );
and ( n2655 , n843 , n2186 );
nor ( n2656 , n2654 , n2655 );
xnor ( n2657 , n2656 , n1841 );
and ( n2658 , n1083 , n1866 );
and ( n2659 , n984 , n1864 );
nor ( n2660 , n2658 , n2659 );
xnor ( n2661 , n2660 , n1844 );
and ( n2662 , n2657 , n2661 );
and ( n2663 , n2661 , n2459 );
and ( n2664 , n2657 , n2459 );
or ( n2665 , n2662 , n2663 , n2664 );
and ( n2666 , n2653 , n2665 );
and ( n2667 , n2015 , n973 );
and ( n2668 , n1833 , n971 );
nor ( n2669 , n2667 , n2668 );
xnor ( n2670 , n2669 , n840 );
and ( n2671 , n2665 , n2670 );
and ( n2672 , n2653 , n2670 );
or ( n2673 , n2666 , n2671 , n2672 );
and ( n2674 , n1290 , n1652 );
and ( n2675 , n1098 , n1650 );
nor ( n2676 , n2674 , n2675 );
xnor ( n2677 , n2676 , n1597 );
and ( n2678 , n1413 , n1538 );
and ( n2679 , n1308 , n1536 );
nor ( n2680 , n2678 , n2679 );
xnor ( n2681 , n2680 , n1433 );
and ( n2682 , n2677 , n2681 );
and ( n2683 , n1659 , n1298 );
and ( n2684 , n1572 , n1296 );
nor ( n2685 , n2683 , n2684 );
xnor ( n2686 , n2685 , n1184 );
and ( n2687 , n2681 , n2686 );
and ( n2688 , n2677 , n2686 );
or ( n2689 , n2682 , n2687 , n2688 );
xor ( n2690 , n2425 , n2429 );
xor ( n2691 , n2690 , n2434 );
and ( n2692 , n2689 , n2691 );
xor ( n2693 , n2441 , n2445 );
xor ( n2694 , n2693 , n2450 );
and ( n2695 , n2691 , n2694 );
and ( n2696 , n2689 , n2694 );
or ( n2697 , n2692 , n2695 , n2696 );
and ( n2698 , n2673 , n2697 );
xor ( n2699 , n2437 , n2453 );
xor ( n2700 , n2699 , n2462 );
and ( n2701 , n2697 , n2700 );
and ( n2702 , n2673 , n2700 );
or ( n2703 , n2698 , n2701 , n2702 );
xor ( n2704 , n2465 , n2467 );
xor ( n2705 , n2704 , n2470 );
and ( n2706 , n2703 , n2705 );
xor ( n2707 , n2594 , n2596 );
xor ( n2708 , n2707 , n2599 );
and ( n2709 , n2705 , n2708 );
and ( n2710 , n2703 , n2708 );
or ( n2711 , n2706 , n2709 , n2710 );
xor ( n2712 , n2537 , n2540 );
and ( n2713 , n897 , n2336 );
and ( n2714 , n908 , n2333 );
nor ( n2715 , n2713 , n2714 );
xnor ( n2716 , n2715 , n1923 );
and ( n2717 , n1010 , n1948 );
and ( n2718 , n917 , n1946 );
nor ( n2719 , n2717 , n2718 );
xnor ( n2720 , n2719 , n1926 );
and ( n2721 , n2716 , n2720 );
and ( n2722 , n2720 , n2538 );
and ( n2723 , n2716 , n2538 );
or ( n2724 , n2721 , n2722 , n2723 );
and ( n2725 , n2712 , n2724 );
and ( n2726 , n2068 , n888 );
and ( n2727 , n1915 , n886 );
nor ( n2728 , n2726 , n2727 );
xnor ( n2729 , n2728 , n893 );
and ( n2730 , n2724 , n2729 );
and ( n2731 , n2712 , n2729 );
or ( n2732 , n2725 , n2730 , n2731 );
and ( n2733 , n1224 , n1760 );
and ( n2734 , n1025 , n1758 );
nor ( n2735 , n2733 , n2734 );
xnor ( n2736 , n2735 , n1705 );
and ( n2737 , n1337 , n1464 );
and ( n2738 , n1242 , n1462 );
nor ( n2739 , n2737 , n2738 );
xnor ( n2740 , n2739 , n1357 );
and ( n2741 , n2736 , n2740 );
and ( n2742 , n1767 , n1232 );
and ( n2743 , n1498 , n1230 );
nor ( n2744 , n2742 , n2743 );
xnor ( n2745 , n2744 , n1131 );
and ( n2746 , n2740 , n2745 );
and ( n2747 , n2736 , n2745 );
or ( n2748 , n2741 , n2746 , n2747 );
xor ( n2749 , n2504 , n2508 );
xor ( n2750 , n2749 , n2513 );
and ( n2751 , n2748 , n2750 );
xor ( n2752 , n2520 , n2524 );
xor ( n2753 , n2752 , n2529 );
and ( n2754 , n2750 , n2753 );
and ( n2755 , n2748 , n2753 );
or ( n2756 , n2751 , n2754 , n2755 );
and ( n2757 , n2732 , n2756 );
xor ( n2758 , n2516 , n2532 );
xor ( n2759 , n2758 , n2541 );
and ( n2760 , n2756 , n2759 );
and ( n2761 , n2732 , n2759 );
or ( n2762 , n2757 , n2760 , n2761 );
xor ( n2763 , n2544 , n2546 );
xor ( n2764 , n2763 , n2549 );
and ( n2765 , n2762 , n2764 );
xor ( n2766 , n2620 , n2622 );
xor ( n2767 , n2766 , n2625 );
and ( n2768 , n2764 , n2767 );
and ( n2769 , n2762 , n2767 );
or ( n2770 , n2765 , n2768 , n2769 );
and ( n2771 , n2711 , n2770 );
xor ( n2772 , n2628 , n2630 );
xor ( n2773 , n2772 , n2633 );
and ( n2774 , n2770 , n2773 );
and ( n2775 , n2711 , n2773 );
or ( n2776 , n2771 , n2774 , n2775 );
xor ( n2777 , n2479 , n2481 );
xor ( n2778 , n2777 , n2484 );
and ( n2779 , n2776 , n2778 );
xor ( n2780 , n2610 , n2636 );
xor ( n2781 , n2780 , n2639 );
and ( n2782 , n2778 , n2781 );
and ( n2783 , n2776 , n2781 );
or ( n2784 , n2779 , n2782 , n2783 );
xor ( n2785 , n2642 , n2644 );
xor ( n2786 , n2785 , n2647 );
and ( n2787 , n2784 , n2786 );
xor ( n2788 , n2784 , n2786 );
xor ( n2789 , n2776 , n2778 );
xor ( n2790 , n2789 , n2781 );
and ( n2791 , n984 , n2189 );
and ( n2792 , n863 , n2186 );
nor ( n2793 , n2791 , n2792 );
xnor ( n2794 , n2793 , n1841 );
and ( n2795 , n2199 , n971 );
not ( n2796 , n2795 );
and ( n2797 , n2796 , n840 );
and ( n2798 , n2794 , n2797 );
and ( n2799 , n1833 , n1106 );
and ( n2800 , n1674 , n1104 );
nor ( n2801 , n2799 , n2800 );
xnor ( n2802 , n2801 , n1075 );
and ( n2803 , n2798 , n2802 );
and ( n2804 , n2158 , n973 );
and ( n2805 , n2015 , n971 );
nor ( n2806 , n2804 , n2805 );
xnor ( n2807 , n2806 , n840 );
and ( n2808 , n2802 , n2807 );
and ( n2809 , n2798 , n2807 );
or ( n2810 , n2803 , n2808 , n2809 );
and ( n2811 , n1308 , n1652 );
and ( n2812 , n1290 , n1650 );
nor ( n2813 , n2811 , n2812 );
xnor ( n2814 , n2813 , n1597 );
and ( n2815 , n2015 , n1106 );
and ( n2816 , n1833 , n1104 );
nor ( n2817 , n2815 , n2816 );
xnor ( n2818 , n2817 , n1075 );
and ( n2819 , n2814 , n2818 );
and ( n2820 , n2199 , n973 );
and ( n2821 , n2158 , n971 );
nor ( n2822 , n2820 , n2821 );
xnor ( n2823 , n2822 , n840 );
and ( n2824 , n2818 , n2823 );
and ( n2825 , n2814 , n2823 );
or ( n2826 , n2819 , n2824 , n2825 );
and ( n2827 , n1098 , n1866 );
and ( n2828 , n1083 , n1864 );
nor ( n2829 , n2827 , n2828 );
xnor ( n2830 , n2829 , n1844 );
and ( n2831 , n1572 , n1538 );
and ( n2832 , n1413 , n1536 );
nor ( n2833 , n2831 , n2832 );
xnor ( n2834 , n2833 , n1433 );
and ( n2835 , n2830 , n2834 );
and ( n2836 , n1674 , n1298 );
and ( n2837 , n1659 , n1296 );
nor ( n2838 , n2836 , n2837 );
xnor ( n2839 , n2838 , n1184 );
and ( n2840 , n2834 , n2839 );
and ( n2841 , n2830 , n2839 );
or ( n2842 , n2835 , n2840 , n2841 );
and ( n2843 , n2826 , n2842 );
xor ( n2844 , n2657 , n2661 );
xor ( n2845 , n2844 , n2459 );
and ( n2846 , n2842 , n2845 );
and ( n2847 , n2826 , n2845 );
or ( n2848 , n2843 , n2846 , n2847 );
and ( n2849 , n2810 , n2848 );
xor ( n2850 , n2653 , n2665 );
xor ( n2851 , n2850 , n2670 );
and ( n2852 , n2848 , n2851 );
and ( n2853 , n2810 , n2851 );
or ( n2854 , n2849 , n2852 , n2853 );
xor ( n2855 , n2586 , n2588 );
xor ( n2856 , n2855 , n2591 );
and ( n2857 , n2854 , n2856 );
xor ( n2858 , n2673 , n2697 );
xor ( n2859 , n2858 , n2700 );
and ( n2860 , n2856 , n2859 );
and ( n2861 , n2854 , n2859 );
or ( n2862 , n2857 , n2860 , n2861 );
and ( n2863 , n917 , n2336 );
and ( n2864 , n897 , n2333 );
nor ( n2865 , n2863 , n2864 );
xnor ( n2866 , n2865 , n1923 );
and ( n2867 , n2346 , n886 );
not ( n2868 , n2867 );
and ( n2869 , n2868 , n893 );
and ( n2870 , n2866 , n2869 );
and ( n2871 , n1915 , n1033 );
and ( n2872 , n1782 , n1031 );
nor ( n2873 , n2871 , n2872 );
xnor ( n2874 , n2873 , n1002 );
and ( n2875 , n2870 , n2874 );
and ( n2876 , n2289 , n888 );
and ( n2877 , n2068 , n886 );
nor ( n2878 , n2876 , n2877 );
xnor ( n2879 , n2878 , n893 );
and ( n2880 , n2874 , n2879 );
and ( n2881 , n2870 , n2879 );
or ( n2882 , n2875 , n2880 , n2881 );
and ( n2883 , n1025 , n1948 );
and ( n2884 , n1010 , n1946 );
nor ( n2885 , n2883 , n2884 );
xnor ( n2886 , n2885 , n1926 );
and ( n2887 , n1498 , n1464 );
and ( n2888 , n1337 , n1462 );
nor ( n2889 , n2887 , n2888 );
xnor ( n2890 , n2889 , n1357 );
and ( n2891 , n2886 , n2890 );
and ( n2892 , n1782 , n1232 );
and ( n2893 , n1767 , n1230 );
nor ( n2894 , n2892 , n2893 );
xnor ( n2895 , n2894 , n1131 );
and ( n2896 , n2890 , n2895 );
and ( n2897 , n2886 , n2895 );
or ( n2898 , n2891 , n2896 , n2897 );
and ( n2899 , n1242 , n1760 );
and ( n2900 , n1224 , n1758 );
nor ( n2901 , n2899 , n2900 );
xnor ( n2902 , n2901 , n1705 );
and ( n2903 , n2068 , n1033 );
and ( n2904 , n1915 , n1031 );
nor ( n2905 , n2903 , n2904 );
xnor ( n2906 , n2905 , n1002 );
and ( n2907 , n2902 , n2906 );
and ( n2908 , n2346 , n888 );
and ( n2909 , n2289 , n886 );
nor ( n2910 , n2908 , n2909 );
xnor ( n2911 , n2910 , n893 );
and ( n2912 , n2906 , n2911 );
and ( n2913 , n2902 , n2911 );
or ( n2914 , n2907 , n2912 , n2913 );
and ( n2915 , n2898 , n2914 );
xor ( n2916 , n2716 , n2720 );
xor ( n2917 , n2916 , n2538 );
and ( n2918 , n2914 , n2917 );
and ( n2919 , n2898 , n2917 );
or ( n2920 , n2915 , n2918 , n2919 );
and ( n2921 , n2882 , n2920 );
xor ( n2922 , n2712 , n2724 );
xor ( n2923 , n2922 , n2729 );
and ( n2924 , n2920 , n2923 );
and ( n2925 , n2882 , n2923 );
or ( n2926 , n2921 , n2924 , n2925 );
xor ( n2927 , n2612 , n2614 );
xor ( n2928 , n2927 , n2617 );
and ( n2929 , n2926 , n2928 );
xor ( n2930 , n2732 , n2756 );
xor ( n2931 , n2930 , n2759 );
and ( n2932 , n2928 , n2931 );
and ( n2933 , n2926 , n2931 );
or ( n2934 , n2929 , n2932 , n2933 );
and ( n2935 , n2862 , n2934 );
xor ( n2936 , n2762 , n2764 );
xor ( n2937 , n2936 , n2767 );
and ( n2938 , n2934 , n2937 );
and ( n2939 , n2862 , n2937 );
or ( n2940 , n2935 , n2938 , n2939 );
xor ( n2941 , n2602 , n2604 );
xor ( n2942 , n2941 , n2607 );
and ( n2943 , n2940 , n2942 );
xor ( n2944 , n2711 , n2770 );
xor ( n2945 , n2944 , n2773 );
and ( n2946 , n2942 , n2945 );
and ( n2947 , n2940 , n2945 );
or ( n2948 , n2943 , n2946 , n2947 );
and ( n2949 , n2790 , n2948 );
xor ( n2950 , n2790 , n2948 );
xor ( n2951 , n2794 , n2797 );
and ( n2952 , n1083 , n2189 );
and ( n2953 , n984 , n2186 );
nor ( n2954 , n2952 , n2953 );
xnor ( n2955 , n2954 , n1841 );
and ( n2956 , n1833 , n1298 );
and ( n2957 , n1674 , n1296 );
nor ( n2958 , n2956 , n2957 );
xnor ( n2959 , n2958 , n1184 );
and ( n2960 , n2955 , n2959 );
and ( n2961 , n2158 , n1106 );
and ( n2962 , n2015 , n1104 );
nor ( n2963 , n2961 , n2962 );
xnor ( n2964 , n2963 , n1075 );
and ( n2965 , n2959 , n2964 );
and ( n2966 , n2955 , n2964 );
or ( n2967 , n2960 , n2965 , n2966 );
and ( n2968 , n2951 , n2967 );
and ( n2969 , n1290 , n1866 );
and ( n2970 , n1098 , n1864 );
nor ( n2971 , n2969 , n2970 );
xnor ( n2972 , n2971 , n1844 );
and ( n2973 , n1659 , n1538 );
and ( n2974 , n1572 , n1536 );
nor ( n2975 , n2973 , n2974 );
xnor ( n2976 , n2975 , n1433 );
and ( n2977 , n2972 , n2976 );
and ( n2978 , n2976 , n2795 );
and ( n2979 , n2972 , n2795 );
or ( n2980 , n2977 , n2978 , n2979 );
and ( n2981 , n2967 , n2980 );
and ( n2982 , n2951 , n2980 );
or ( n2983 , n2968 , n2981 , n2982 );
xor ( n2984 , n2677 , n2681 );
xor ( n2985 , n2984 , n2686 );
and ( n2986 , n2983 , n2985 );
xor ( n2987 , n2798 , n2802 );
xor ( n2988 , n2987 , n2807 );
and ( n2989 , n2985 , n2988 );
and ( n2990 , n2983 , n2988 );
or ( n2991 , n2986 , n2989 , n2990 );
xor ( n2992 , n2689 , n2691 );
xor ( n2993 , n2992 , n2694 );
and ( n2994 , n2991 , n2993 );
xor ( n2995 , n2810 , n2848 );
xor ( n2996 , n2995 , n2851 );
and ( n2997 , n2993 , n2996 );
and ( n2998 , n2991 , n2996 );
or ( n2999 , n2994 , n2997 , n2998 );
xor ( n3000 , n2866 , n2869 );
and ( n3001 , n1224 , n1948 );
and ( n3002 , n1025 , n1946 );
nor ( n3003 , n3001 , n3002 );
xnor ( n3004 , n3003 , n1926 );
and ( n3005 , n1767 , n1464 );
and ( n3006 , n1498 , n1462 );
nor ( n3007 , n3005 , n3006 );
xnor ( n3008 , n3007 , n1357 );
and ( n3009 , n3004 , n3008 );
and ( n3010 , n3008 , n2867 );
and ( n3011 , n3004 , n2867 );
or ( n3012 , n3009 , n3010 , n3011 );
and ( n3013 , n3000 , n3012 );
and ( n3014 , n1010 , n2336 );
and ( n3015 , n917 , n2333 );
nor ( n3016 , n3014 , n3015 );
xnor ( n3017 , n3016 , n1923 );
and ( n3018 , n1915 , n1232 );
and ( n3019 , n1782 , n1230 );
nor ( n3020 , n3018 , n3019 );
xnor ( n3021 , n3020 , n1131 );
and ( n3022 , n3017 , n3021 );
and ( n3023 , n2289 , n1033 );
and ( n3024 , n2068 , n1031 );
nor ( n3025 , n3023 , n3024 );
xnor ( n3026 , n3025 , n1002 );
and ( n3027 , n3021 , n3026 );
and ( n3028 , n3017 , n3026 );
or ( n3029 , n3022 , n3027 , n3028 );
and ( n3030 , n3012 , n3029 );
and ( n3031 , n3000 , n3029 );
or ( n3032 , n3013 , n3030 , n3031 );
xor ( n3033 , n2736 , n2740 );
xor ( n3034 , n3033 , n2745 );
and ( n3035 , n3032 , n3034 );
xor ( n3036 , n2870 , n2874 );
xor ( n3037 , n3036 , n2879 );
and ( n3038 , n3034 , n3037 );
and ( n3039 , n3032 , n3037 );
or ( n3040 , n3035 , n3038 , n3039 );
xor ( n3041 , n2748 , n2750 );
xor ( n3042 , n3041 , n2753 );
and ( n3043 , n3040 , n3042 );
xor ( n3044 , n2882 , n2920 );
xor ( n3045 , n3044 , n2923 );
and ( n3046 , n3042 , n3045 );
and ( n3047 , n3040 , n3045 );
or ( n3048 , n3043 , n3046 , n3047 );
and ( n3049 , n2999 , n3048 );
xor ( n3050 , n2926 , n2928 );
xor ( n3051 , n3050 , n2931 );
and ( n3052 , n3048 , n3051 );
and ( n3053 , n2999 , n3051 );
or ( n3054 , n3049 , n3052 , n3053 );
xor ( n3055 , n2703 , n2705 );
xor ( n3056 , n3055 , n2708 );
and ( n3057 , n3054 , n3056 );
xor ( n3058 , n2862 , n2934 );
xor ( n3059 , n3058 , n2937 );
and ( n3060 , n3056 , n3059 );
and ( n3061 , n3054 , n3059 );
or ( n3062 , n3057 , n3060 , n3061 );
xor ( n3063 , n2940 , n2942 );
xor ( n3064 , n3063 , n2945 );
and ( n3065 , n3062 , n3064 );
xor ( n3066 , n3062 , n3064 );
xor ( n3067 , n3054 , n3056 );
xor ( n3068 , n3067 , n3059 );
and ( n3069 , n1098 , n2189 );
and ( n3070 , n1083 , n2186 );
nor ( n3071 , n3069 , n3070 );
xnor ( n3072 , n3071 , n1841 );
and ( n3073 , n1674 , n1538 );
and ( n3074 , n1659 , n1536 );
nor ( n3075 , n3073 , n3074 );
xnor ( n3076 , n3075 , n1433 );
and ( n3077 , n3072 , n3076 );
and ( n3078 , n2015 , n1298 );
and ( n3079 , n1833 , n1296 );
nor ( n3080 , n3078 , n3079 );
xnor ( n3081 , n3080 , n1184 );
and ( n3082 , n3076 , n3081 );
and ( n3083 , n3072 , n3081 );
or ( n3084 , n3077 , n3082 , n3083 );
and ( n3085 , n1308 , n1866 );
and ( n3086 , n1290 , n1864 );
nor ( n3087 , n3085 , n3086 );
xnor ( n3088 , n3087 , n1844 );
and ( n3089 , n2199 , n1104 );
not ( n3090 , n3089 );
and ( n3091 , n3090 , n1075 );
and ( n3092 , n3088 , n3091 );
and ( n3093 , n3084 , n3092 );
and ( n3094 , n1413 , n1652 );
and ( n3095 , n1308 , n1650 );
nor ( n3096 , n3094 , n3095 );
xnor ( n3097 , n3096 , n1597 );
and ( n3098 , n3092 , n3097 );
and ( n3099 , n3084 , n3097 );
or ( n3100 , n3093 , n3098 , n3099 );
xor ( n3101 , n2814 , n2818 );
xor ( n3102 , n3101 , n2823 );
and ( n3103 , n3100 , n3102 );
xor ( n3104 , n2830 , n2834 );
xor ( n3105 , n3104 , n2839 );
and ( n3106 , n3102 , n3105 );
and ( n3107 , n3100 , n3105 );
or ( n3108 , n3103 , n3106 , n3107 );
xor ( n3109 , n2826 , n2842 );
xor ( n3110 , n3109 , n2845 );
and ( n3111 , n3108 , n3110 );
xor ( n3112 , n2983 , n2985 );
xor ( n3113 , n3112 , n2988 );
and ( n3114 , n3110 , n3113 );
and ( n3115 , n3108 , n3113 );
or ( n3116 , n3111 , n3114 , n3115 );
and ( n3117 , n1025 , n2336 );
and ( n3118 , n1010 , n2333 );
nor ( n3119 , n3117 , n3118 );
xnor ( n3120 , n3119 , n1923 );
and ( n3121 , n1782 , n1464 );
and ( n3122 , n1767 , n1462 );
nor ( n3123 , n3121 , n3122 );
xnor ( n3124 , n3123 , n1357 );
and ( n3125 , n3120 , n3124 );
and ( n3126 , n2068 , n1232 );
and ( n3127 , n1915 , n1230 );
nor ( n3128 , n3126 , n3127 );
xnor ( n3129 , n3128 , n1131 );
and ( n3130 , n3124 , n3129 );
and ( n3131 , n3120 , n3129 );
or ( n3132 , n3125 , n3130 , n3131 );
and ( n3133 , n1242 , n1948 );
and ( n3134 , n1224 , n1946 );
nor ( n3135 , n3133 , n3134 );
xnor ( n3136 , n3135 , n1926 );
and ( n3137 , n2346 , n1031 );
not ( n3138 , n3137 );
and ( n3139 , n3138 , n1002 );
and ( n3140 , n3136 , n3139 );
and ( n3141 , n3132 , n3140 );
and ( n3142 , n1337 , n1760 );
and ( n3143 , n1242 , n1758 );
nor ( n3144 , n3142 , n3143 );
xnor ( n3145 , n3144 , n1705 );
and ( n3146 , n3140 , n3145 );
and ( n3147 , n3132 , n3145 );
or ( n3148 , n3141 , n3146 , n3147 );
xor ( n3149 , n2886 , n2890 );
xor ( n3150 , n3149 , n2895 );
and ( n3151 , n3148 , n3150 );
xor ( n3152 , n2902 , n2906 );
xor ( n3153 , n3152 , n2911 );
and ( n3154 , n3150 , n3153 );
and ( n3155 , n3148 , n3153 );
or ( n3156 , n3151 , n3154 , n3155 );
xor ( n3157 , n2898 , n2914 );
xor ( n3158 , n3157 , n2917 );
and ( n3159 , n3156 , n3158 );
xor ( n3160 , n3032 , n3034 );
xor ( n3161 , n3160 , n3037 );
and ( n3162 , n3158 , n3161 );
and ( n3163 , n3156 , n3161 );
or ( n3164 , n3159 , n3162 , n3163 );
and ( n3165 , n3116 , n3164 );
xor ( n3166 , n3040 , n3042 );
xor ( n3167 , n3166 , n3045 );
and ( n3168 , n3164 , n3167 );
and ( n3169 , n3116 , n3167 );
or ( n3170 , n3165 , n3168 , n3169 );
xor ( n3171 , n2854 , n2856 );
xor ( n3172 , n3171 , n2859 );
and ( n3173 , n3170 , n3172 );
xor ( n3174 , n2999 , n3048 );
xor ( n3175 , n3174 , n3051 );
and ( n3176 , n3172 , n3175 );
and ( n3177 , n3170 , n3175 );
or ( n3178 , n3173 , n3176 , n3177 );
and ( n3179 , n3068 , n3178 );
xor ( n3180 , n3068 , n3178 );
xor ( n3181 , n3170 , n3172 );
xor ( n3182 , n3181 , n3175 );
xor ( n3183 , n3088 , n3091 );
and ( n3184 , n1572 , n1652 );
and ( n3185 , n1413 , n1650 );
nor ( n3186 , n3184 , n3185 );
xnor ( n3187 , n3186 , n1597 );
and ( n3188 , n3183 , n3187 );
and ( n3189 , n2199 , n1106 );
and ( n3190 , n2158 , n1104 );
nor ( n3191 , n3189 , n3190 );
xnor ( n3192 , n3191 , n1075 );
and ( n3193 , n3187 , n3192 );
and ( n3194 , n3183 , n3192 );
or ( n3195 , n3188 , n3193 , n3194 );
xor ( n3196 , n2955 , n2959 );
xor ( n3197 , n3196 , n2964 );
and ( n3198 , n3195 , n3197 );
xor ( n3199 , n2972 , n2976 );
xor ( n3200 , n3199 , n2795 );
and ( n3201 , n3197 , n3200 );
and ( n3202 , n3195 , n3200 );
or ( n3203 , n3198 , n3201 , n3202 );
xor ( n3204 , n2951 , n2967 );
xor ( n3205 , n3204 , n2980 );
and ( n3206 , n3203 , n3205 );
xor ( n3207 , n3100 , n3102 );
xor ( n3208 , n3207 , n3105 );
and ( n3209 , n3205 , n3208 );
and ( n3210 , n3203 , n3208 );
or ( n3211 , n3206 , n3209 , n3210 );
xor ( n3212 , n3136 , n3139 );
and ( n3213 , n1498 , n1760 );
and ( n3214 , n1337 , n1758 );
nor ( n3215 , n3213 , n3214 );
xnor ( n3216 , n3215 , n1705 );
and ( n3217 , n3212 , n3216 );
and ( n3218 , n2346 , n1033 );
and ( n3219 , n2289 , n1031 );
nor ( n3220 , n3218 , n3219 );
xnor ( n3221 , n3220 , n1002 );
and ( n3222 , n3216 , n3221 );
and ( n3223 , n3212 , n3221 );
or ( n3224 , n3217 , n3222 , n3223 );
xor ( n3225 , n3004 , n3008 );
xor ( n3226 , n3225 , n2867 );
and ( n3227 , n3224 , n3226 );
xor ( n3228 , n3017 , n3021 );
xor ( n3229 , n3228 , n3026 );
and ( n3230 , n3226 , n3229 );
and ( n3231 , n3224 , n3229 );
or ( n3232 , n3227 , n3230 , n3231 );
xor ( n3233 , n3000 , n3012 );
xor ( n3234 , n3233 , n3029 );
and ( n3235 , n3232 , n3234 );
xor ( n3236 , n3148 , n3150 );
xor ( n3237 , n3236 , n3153 );
and ( n3238 , n3234 , n3237 );
and ( n3239 , n3232 , n3237 );
or ( n3240 , n3235 , n3238 , n3239 );
and ( n3241 , n3211 , n3240 );
xor ( n3242 , n3156 , n3158 );
xor ( n3243 , n3242 , n3161 );
and ( n3244 , n3240 , n3243 );
and ( n3245 , n3211 , n3243 );
or ( n3246 , n3241 , n3244 , n3245 );
xor ( n3247 , n2991 , n2993 );
xor ( n3248 , n3247 , n2996 );
and ( n3249 , n3246 , n3248 );
xor ( n3250 , n3116 , n3164 );
xor ( n3251 , n3250 , n3167 );
and ( n3252 , n3248 , n3251 );
and ( n3253 , n3246 , n3251 );
or ( n3254 , n3249 , n3252 , n3253 );
and ( n3255 , n3182 , n3254 );
xor ( n3256 , n3182 , n3254 );
xor ( n3257 , n3246 , n3248 );
xor ( n3258 , n3257 , n3251 );
and ( n3259 , n1224 , n2336 );
and ( n3260 , n1025 , n2333 );
nor ( n3261 , n3259 , n3260 );
xnor ( n3262 , n3261 , n1923 );
and ( n3263 , n1767 , n1760 );
and ( n3264 , n1498 , n1758 );
nor ( n3265 , n3263 , n3264 );
xnor ( n3266 , n3265 , n1705 );
and ( n3267 , n3262 , n3266 );
and ( n3268 , n2289 , n1232 );
and ( n3269 , n2068 , n1230 );
nor ( n3270 , n3268 , n3269 );
xnor ( n3271 , n3270 , n1131 );
and ( n3272 , n3266 , n3271 );
and ( n3273 , n3262 , n3271 );
or ( n3274 , n3267 , n3272 , n3273 );
and ( n3275 , n1337 , n1948 );
and ( n3276 , n1242 , n1946 );
nor ( n3277 , n3275 , n3276 );
xnor ( n3278 , n3277 , n1926 );
and ( n3279 , n1915 , n1464 );
and ( n3280 , n1782 , n1462 );
nor ( n3281 , n3279 , n3280 );
xnor ( n3282 , n3281 , n1357 );
and ( n3283 , n3278 , n3282 );
and ( n3284 , n3282 , n3137 );
and ( n3285 , n3278 , n3137 );
or ( n3286 , n3283 , n3284 , n3285 );
and ( n3287 , n3274 , n3286 );
xor ( n3288 , n3120 , n3124 );
xor ( n3289 , n3288 , n3129 );
and ( n3290 , n3286 , n3289 );
and ( n3291 , n3274 , n3289 );
or ( n3292 , n3287 , n3290 , n3291 );
xor ( n3293 , n3132 , n3140 );
xor ( n3294 , n3293 , n3145 );
and ( n3295 , n3292 , n3294 );
xor ( n3296 , n3224 , n3226 );
xor ( n3297 , n3296 , n3229 );
and ( n3298 , n3294 , n3297 );
and ( n3299 , n3292 , n3297 );
or ( n3300 , n3295 , n3298 , n3299 );
and ( n3301 , n1290 , n2189 );
and ( n3302 , n1098 , n2186 );
nor ( n3303 , n3301 , n3302 );
xnor ( n3304 , n3303 , n1841 );
and ( n3305 , n1659 , n1652 );
and ( n3306 , n1572 , n1650 );
nor ( n3307 , n3305 , n3306 );
xnor ( n3308 , n3307 , n1597 );
and ( n3309 , n3304 , n3308 );
and ( n3310 , n2158 , n1298 );
and ( n3311 , n2015 , n1296 );
nor ( n3312 , n3310 , n3311 );
xnor ( n3313 , n3312 , n1184 );
and ( n3314 , n3308 , n3313 );
and ( n3315 , n3304 , n3313 );
or ( n3316 , n3309 , n3314 , n3315 );
and ( n3317 , n1413 , n1866 );
and ( n3318 , n1308 , n1864 );
nor ( n3319 , n3317 , n3318 );
xnor ( n3320 , n3319 , n1844 );
and ( n3321 , n1833 , n1538 );
and ( n3322 , n1674 , n1536 );
nor ( n3323 , n3321 , n3322 );
xnor ( n3324 , n3323 , n1433 );
and ( n3325 , n3320 , n3324 );
and ( n3326 , n3324 , n3089 );
and ( n3327 , n3320 , n3089 );
or ( n3328 , n3325 , n3326 , n3327 );
and ( n3329 , n3316 , n3328 );
xor ( n3330 , n3072 , n3076 );
xor ( n3331 , n3330 , n3081 );
and ( n3332 , n3328 , n3331 );
and ( n3333 , n3316 , n3331 );
or ( n3334 , n3329 , n3332 , n3333 );
xor ( n3335 , n3084 , n3092 );
xor ( n3336 , n3335 , n3097 );
and ( n3337 , n3334 , n3336 );
xor ( n3338 , n3195 , n3197 );
xor ( n3339 , n3338 , n3200 );
and ( n3340 , n3336 , n3339 );
and ( n3341 , n3334 , n3339 );
or ( n3342 , n3337 , n3340 , n3341 );
and ( n3343 , n3300 , n3342 );
xor ( n3344 , n3232 , n3234 );
xor ( n3345 , n3344 , n3237 );
and ( n3346 , n3342 , n3345 );
and ( n3347 , n3300 , n3345 );
or ( n3348 , n3343 , n3346 , n3347 );
xor ( n3349 , n3108 , n3110 );
xor ( n3350 , n3349 , n3113 );
and ( n3351 , n3348 , n3350 );
xor ( n3352 , n3211 , n3240 );
xor ( n3353 , n3352 , n3243 );
and ( n3354 , n3350 , n3353 );
and ( n3355 , n3348 , n3353 );
or ( n3356 , n3351 , n3354 , n3355 );
and ( n3357 , n3258 , n3356 );
xor ( n3358 , n3258 , n3356 );
xor ( n3359 , n3348 , n3350 );
xor ( n3360 , n3359 , n3353 );
and ( n3361 , n1308 , n2189 );
and ( n3362 , n1290 , n2186 );
nor ( n3363 , n3361 , n3362 );
xnor ( n3364 , n3363 , n1841 );
and ( n3365 , n2015 , n1538 );
and ( n3366 , n1833 , n1536 );
nor ( n3367 , n3365 , n3366 );
xnor ( n3368 , n3367 , n1433 );
and ( n3369 , n3364 , n3368 );
and ( n3370 , n2199 , n1298 );
and ( n3371 , n2158 , n1296 );
nor ( n3372 , n3370 , n3371 );
xnor ( n3373 , n3372 , n1184 );
and ( n3374 , n3368 , n3373 );
and ( n3375 , n3364 , n3373 );
or ( n3376 , n3369 , n3374 , n3375 );
and ( n3377 , n1572 , n1866 );
and ( n3378 , n1413 , n1864 );
nor ( n3379 , n3377 , n3378 );
xnor ( n3380 , n3379 , n1844 );
and ( n3381 , n2199 , n1296 );
not ( n3382 , n3381 );
and ( n3383 , n3382 , n1184 );
and ( n3384 , n3380 , n3383 );
and ( n3385 , n3376 , n3384 );
xor ( n3386 , n3320 , n3324 );
xor ( n3387 , n3386 , n3089 );
and ( n3388 , n3384 , n3387 );
and ( n3389 , n3376 , n3387 );
or ( n3390 , n3385 , n3388 , n3389 );
xor ( n3391 , n3183 , n3187 );
xor ( n3392 , n3391 , n3192 );
and ( n3393 , n3390 , n3392 );
xor ( n3394 , n3316 , n3328 );
xor ( n3395 , n3394 , n3331 );
and ( n3396 , n3392 , n3395 );
and ( n3397 , n3390 , n3395 );
or ( n3398 , n3393 , n3396 , n3397 );
and ( n3399 , n1242 , n2336 );
and ( n3400 , n1224 , n2333 );
nor ( n3401 , n3399 , n3400 );
xnor ( n3402 , n3401 , n1923 );
and ( n3403 , n2068 , n1464 );
and ( n3404 , n1915 , n1462 );
nor ( n3405 , n3403 , n3404 );
xnor ( n3406 , n3405 , n1357 );
and ( n3407 , n3402 , n3406 );
and ( n3408 , n2346 , n1232 );
and ( n3409 , n2289 , n1230 );
nor ( n3410 , n3408 , n3409 );
xnor ( n3411 , n3410 , n1131 );
and ( n3412 , n3406 , n3411 );
and ( n3413 , n3402 , n3411 );
or ( n3414 , n3407 , n3412 , n3413 );
and ( n3415 , n1498 , n1948 );
and ( n3416 , n1337 , n1946 );
nor ( n3417 , n3415 , n3416 );
xnor ( n3418 , n3417 , n1926 );
and ( n3419 , n2346 , n1230 );
not ( n3420 , n3419 );
and ( n3421 , n3420 , n1131 );
and ( n3422 , n3418 , n3421 );
and ( n3423 , n3414 , n3422 );
xor ( n3424 , n3278 , n3282 );
xor ( n3425 , n3424 , n3137 );
and ( n3426 , n3422 , n3425 );
and ( n3427 , n3414 , n3425 );
or ( n3428 , n3423 , n3426 , n3427 );
xor ( n3429 , n3212 , n3216 );
xor ( n3430 , n3429 , n3221 );
and ( n3431 , n3428 , n3430 );
xor ( n3432 , n3274 , n3286 );
xor ( n3433 , n3432 , n3289 );
and ( n3434 , n3430 , n3433 );
and ( n3435 , n3428 , n3433 );
or ( n3436 , n3431 , n3434 , n3435 );
and ( n3437 , n3398 , n3436 );
xor ( n3438 , n3292 , n3294 );
xor ( n3439 , n3438 , n3297 );
and ( n3440 , n3436 , n3439 );
and ( n3441 , n3398 , n3439 );
or ( n3442 , n3437 , n3440 , n3441 );
xor ( n3443 , n3203 , n3205 );
xor ( n3444 , n3443 , n3208 );
and ( n3445 , n3442 , n3444 );
xor ( n3446 , n3300 , n3342 );
xor ( n3447 , n3446 , n3345 );
and ( n3448 , n3444 , n3447 );
and ( n3449 , n3442 , n3447 );
or ( n3450 , n3445 , n3448 , n3449 );
and ( n3451 , n3360 , n3450 );
xor ( n3452 , n3360 , n3450 );
xor ( n3453 , n3442 , n3444 );
xor ( n3454 , n3453 , n3447 );
xor ( n3455 , n3380 , n3383 );
and ( n3456 , n1413 , n2189 );
and ( n3457 , n1308 , n2186 );
nor ( n3458 , n3456 , n3457 );
xnor ( n3459 , n3458 , n1841 );
and ( n3460 , n2158 , n1538 );
and ( n3461 , n2015 , n1536 );
nor ( n3462 , n3460 , n3461 );
xnor ( n3463 , n3462 , n1433 );
and ( n3464 , n3459 , n3463 );
and ( n3465 , n3463 , n3381 );
and ( n3466 , n3459 , n3381 );
or ( n3467 , n3464 , n3465 , n3466 );
and ( n3468 , n3455 , n3467 );
and ( n3469 , n1674 , n1652 );
and ( n3470 , n1659 , n1650 );
nor ( n3471 , n3469 , n3470 );
xnor ( n3472 , n3471 , n1597 );
and ( n3473 , n3467 , n3472 );
and ( n3474 , n3455 , n3472 );
or ( n3475 , n3468 , n3473 , n3474 );
xor ( n3476 , n3304 , n3308 );
xor ( n3477 , n3476 , n3313 );
and ( n3478 , n3475 , n3477 );
xor ( n3479 , n3376 , n3384 );
xor ( n3480 , n3479 , n3387 );
and ( n3481 , n3477 , n3480 );
and ( n3482 , n3475 , n3480 );
or ( n3483 , n3478 , n3481 , n3482 );
xor ( n3484 , n3418 , n3421 );
and ( n3485 , n1337 , n2336 );
and ( n3486 , n1242 , n2333 );
nor ( n3487 , n3485 , n3486 );
xnor ( n3488 , n3487 , n1923 );
and ( n3489 , n2289 , n1464 );
and ( n3490 , n2068 , n1462 );
nor ( n3491 , n3489 , n3490 );
xnor ( n3492 , n3491 , n1357 );
and ( n3493 , n3488 , n3492 );
and ( n3494 , n3492 , n3419 );
and ( n3495 , n3488 , n3419 );
or ( n3496 , n3493 , n3494 , n3495 );
and ( n3497 , n3484 , n3496 );
and ( n3498 , n1782 , n1760 );
and ( n3499 , n1767 , n1758 );
nor ( n3500 , n3498 , n3499 );
xnor ( n3501 , n3500 , n1705 );
and ( n3502 , n3496 , n3501 );
and ( n3503 , n3484 , n3501 );
or ( n3504 , n3497 , n3502 , n3503 );
xor ( n3505 , n3262 , n3266 );
xor ( n3506 , n3505 , n3271 );
and ( n3507 , n3504 , n3506 );
xor ( n3508 , n3414 , n3422 );
xor ( n3509 , n3508 , n3425 );
and ( n3510 , n3506 , n3509 );
and ( n3511 , n3504 , n3509 );
or ( n3512 , n3507 , n3510 , n3511 );
and ( n3513 , n3483 , n3512 );
xor ( n3514 , n3428 , n3430 );
xor ( n3515 , n3514 , n3433 );
and ( n3516 , n3512 , n3515 );
and ( n3517 , n3483 , n3515 );
or ( n3518 , n3513 , n3516 , n3517 );
xor ( n3519 , n3334 , n3336 );
xor ( n3520 , n3519 , n3339 );
and ( n3521 , n3518 , n3520 );
xor ( n3522 , n3398 , n3436 );
xor ( n3523 , n3522 , n3439 );
and ( n3524 , n3520 , n3523 );
and ( n3525 , n3518 , n3523 );
or ( n3526 , n3521 , n3524 , n3525 );
and ( n3527 , n3454 , n3526 );
xor ( n3528 , n3454 , n3526 );
and ( n3529 , n1572 , n2189 );
and ( n3530 , n1413 , n2186 );
nor ( n3531 , n3529 , n3530 );
xnor ( n3532 , n3531 , n1841 );
and ( n3533 , n2199 , n1536 );
not ( n3534 , n3533 );
and ( n3535 , n3534 , n1433 );
and ( n3536 , n3532 , n3535 );
and ( n3537 , n1659 , n1866 );
and ( n3538 , n1572 , n1864 );
nor ( n3539 , n3537 , n3538 );
xnor ( n3540 , n3539 , n1844 );
and ( n3541 , n3536 , n3540 );
and ( n3542 , n1833 , n1652 );
and ( n3543 , n1674 , n1650 );
nor ( n3544 , n3542 , n3543 );
xnor ( n3545 , n3544 , n1597 );
and ( n3546 , n3540 , n3545 );
and ( n3547 , n3536 , n3545 );
or ( n3548 , n3541 , n3546 , n3547 );
xor ( n3549 , n3364 , n3368 );
xor ( n3550 , n3549 , n3373 );
and ( n3551 , n3548 , n3550 );
xor ( n3552 , n3455 , n3467 );
xor ( n3553 , n3552 , n3472 );
and ( n3554 , n3550 , n3553 );
and ( n3555 , n3548 , n3553 );
or ( n3556 , n3551 , n3554 , n3555 );
and ( n3557 , n1498 , n2336 );
and ( n3558 , n1337 , n2333 );
nor ( n3559 , n3557 , n3558 );
xnor ( n3560 , n3559 , n1923 );
and ( n3561 , n2346 , n1462 );
not ( n3562 , n3561 );
and ( n3563 , n3562 , n1357 );
and ( n3564 , n3560 , n3563 );
and ( n3565 , n1767 , n1948 );
and ( n3566 , n1498 , n1946 );
nor ( n3567 , n3565 , n3566 );
xnor ( n3568 , n3567 , n1926 );
and ( n3569 , n3564 , n3568 );
and ( n3570 , n1915 , n1760 );
and ( n3571 , n1782 , n1758 );
nor ( n3572 , n3570 , n3571 );
xnor ( n3573 , n3572 , n1705 );
and ( n3574 , n3568 , n3573 );
and ( n3575 , n3564 , n3573 );
or ( n3576 , n3569 , n3574 , n3575 );
xor ( n3577 , n3402 , n3406 );
xor ( n3578 , n3577 , n3411 );
and ( n3579 , n3576 , n3578 );
xor ( n3580 , n3484 , n3496 );
xor ( n3581 , n3580 , n3501 );
and ( n3582 , n3578 , n3581 );
and ( n3583 , n3576 , n3581 );
or ( n3584 , n3579 , n3582 , n3583 );
and ( n3585 , n3556 , n3584 );
xor ( n3586 , n3504 , n3506 );
xor ( n3587 , n3586 , n3509 );
and ( n3588 , n3584 , n3587 );
and ( n3589 , n3556 , n3587 );
or ( n3590 , n3585 , n3588 , n3589 );
xor ( n3591 , n3390 , n3392 );
xor ( n3592 , n3591 , n3395 );
and ( n3593 , n3590 , n3592 );
xor ( n3594 , n3483 , n3512 );
xor ( n3595 , n3594 , n3515 );
and ( n3596 , n3592 , n3595 );
and ( n3597 , n3590 , n3595 );
or ( n3598 , n3593 , n3596 , n3597 );
xor ( n3599 , n3518 , n3520 );
xor ( n3600 , n3599 , n3523 );
and ( n3601 , n3598 , n3600 );
xor ( n3602 , n3598 , n3600 );
xor ( n3603 , n3590 , n3592 );
xor ( n3604 , n3603 , n3595 );
and ( n3605 , n1674 , n1866 );
and ( n3606 , n1659 , n1864 );
nor ( n3607 , n3605 , n3606 );
xnor ( n3608 , n3607 , n1844 );
and ( n3609 , n2015 , n1652 );
and ( n3610 , n1833 , n1650 );
nor ( n3611 , n3609 , n3610 );
xnor ( n3612 , n3611 , n1597 );
and ( n3613 , n3608 , n3612 );
and ( n3614 , n2199 , n1538 );
and ( n3615 , n2158 , n1536 );
nor ( n3616 , n3614 , n3615 );
xnor ( n3617 , n3616 , n1433 );
and ( n3618 , n3612 , n3617 );
and ( n3619 , n3608 , n3617 );
or ( n3620 , n3613 , n3618 , n3619 );
xor ( n3621 , n3459 , n3463 );
xor ( n3622 , n3621 , n3381 );
and ( n3623 , n3620 , n3622 );
xor ( n3624 , n3536 , n3540 );
xor ( n3625 , n3624 , n3545 );
and ( n3626 , n3622 , n3625 );
and ( n3627 , n3620 , n3625 );
or ( n3628 , n3623 , n3626 , n3627 );
and ( n3629 , n1782 , n1948 );
and ( n3630 , n1767 , n1946 );
nor ( n3631 , n3629 , n3630 );
xnor ( n3632 , n3631 , n1926 );
and ( n3633 , n2068 , n1760 );
and ( n3634 , n1915 , n1758 );
nor ( n3635 , n3633 , n3634 );
xnor ( n3636 , n3635 , n1705 );
and ( n3637 , n3632 , n3636 );
and ( n3638 , n2346 , n1464 );
and ( n3639 , n2289 , n1462 );
nor ( n3640 , n3638 , n3639 );
xnor ( n3641 , n3640 , n1357 );
and ( n3642 , n3636 , n3641 );
and ( n3643 , n3632 , n3641 );
or ( n3644 , n3637 , n3642 , n3643 );
xor ( n3645 , n3488 , n3492 );
xor ( n3646 , n3645 , n3419 );
and ( n3647 , n3644 , n3646 );
xor ( n3648 , n3564 , n3568 );
xor ( n3649 , n3648 , n3573 );
and ( n3650 , n3646 , n3649 );
and ( n3651 , n3644 , n3649 );
or ( n3652 , n3647 , n3650 , n3651 );
and ( n3653 , n3628 , n3652 );
xor ( n3654 , n3576 , n3578 );
xor ( n3655 , n3654 , n3581 );
and ( n3656 , n3652 , n3655 );
and ( n3657 , n3628 , n3655 );
or ( n3658 , n3653 , n3656 , n3657 );
xor ( n3659 , n3475 , n3477 );
xor ( n3660 , n3659 , n3480 );
and ( n3661 , n3658 , n3660 );
xor ( n3662 , n3556 , n3584 );
xor ( n3663 , n3662 , n3587 );
and ( n3664 , n3660 , n3663 );
and ( n3665 , n3658 , n3663 );
or ( n3666 , n3661 , n3664 , n3665 );
and ( n3667 , n3604 , n3666 );
xor ( n3668 , n3604 , n3666 );
xor ( n3669 , n3658 , n3660 );
xor ( n3670 , n3669 , n3663 );
xor ( n3671 , n3532 , n3535 );
and ( n3672 , n1659 , n2189 );
and ( n3673 , n1572 , n2186 );
nor ( n3674 , n3672 , n3673 );
xnor ( n3675 , n3674 , n1841 );
and ( n3676 , n1833 , n1866 );
and ( n3677 , n1674 , n1864 );
nor ( n3678 , n3676 , n3677 );
xnor ( n3679 , n3678 , n1844 );
and ( n3680 , n3675 , n3679 );
and ( n3681 , n3679 , n3533 );
and ( n3682 , n3675 , n3533 );
or ( n3683 , n3680 , n3681 , n3682 );
and ( n3684 , n3671 , n3683 );
xor ( n3685 , n3608 , n3612 );
xor ( n3686 , n3685 , n3617 );
and ( n3687 , n3683 , n3686 );
and ( n3688 , n3671 , n3686 );
or ( n3689 , n3684 , n3687 , n3688 );
xor ( n3690 , n3560 , n3563 );
and ( n3691 , n1767 , n2336 );
and ( n3692 , n1498 , n2333 );
nor ( n3693 , n3691 , n3692 );
xnor ( n3694 , n3693 , n1923 );
and ( n3695 , n1915 , n1948 );
and ( n3696 , n1782 , n1946 );
nor ( n3697 , n3695 , n3696 );
xnor ( n3698 , n3697 , n1926 );
and ( n3699 , n3694 , n3698 );
and ( n3700 , n3698 , n3561 );
and ( n3701 , n3694 , n3561 );
or ( n3702 , n3699 , n3700 , n3701 );
and ( n3703 , n3690 , n3702 );
xor ( n3704 , n3632 , n3636 );
xor ( n3705 , n3704 , n3641 );
and ( n3706 , n3702 , n3705 );
and ( n3707 , n3690 , n3705 );
or ( n3708 , n3703 , n3706 , n3707 );
and ( n3709 , n3689 , n3708 );
xor ( n3710 , n3644 , n3646 );
xor ( n3711 , n3710 , n3649 );
and ( n3712 , n3708 , n3711 );
and ( n3713 , n3689 , n3711 );
or ( n3714 , n3709 , n3712 , n3713 );
xor ( n3715 , n3548 , n3550 );
xor ( n3716 , n3715 , n3553 );
and ( n3717 , n3714 , n3716 );
xor ( n3718 , n3628 , n3652 );
xor ( n3719 , n3718 , n3655 );
and ( n3720 , n3716 , n3719 );
and ( n3721 , n3714 , n3719 );
or ( n3722 , n3717 , n3720 , n3721 );
and ( n3723 , n3670 , n3722 );
xor ( n3724 , n3670 , n3722 );
xor ( n3725 , n3714 , n3716 );
xor ( n3726 , n3725 , n3719 );
and ( n3727 , n1674 , n2189 );
and ( n3728 , n1659 , n2186 );
nor ( n3729 , n3727 , n3728 );
xnor ( n3730 , n3729 , n1841 );
and ( n3731 , n2199 , n1650 );
not ( n3732 , n3731 );
and ( n3733 , n3732 , n1597 );
and ( n3734 , n3730 , n3733 );
and ( n3735 , n2158 , n1652 );
and ( n3736 , n2015 , n1650 );
nor ( n3737 , n3735 , n3736 );
xnor ( n3738 , n3737 , n1597 );
and ( n3739 , n3734 , n3738 );
xor ( n3740 , n3675 , n3679 );
xor ( n3741 , n3740 , n3533 );
and ( n3742 , n3738 , n3741 );
and ( n3743 , n3734 , n3741 );
or ( n3744 , n3739 , n3742 , n3743 );
and ( n3745 , n1782 , n2336 );
and ( n3746 , n1767 , n2333 );
nor ( n3747 , n3745 , n3746 );
xnor ( n3748 , n3747 , n1923 );
and ( n3749 , n2346 , n1758 );
not ( n3750 , n3749 );
and ( n3751 , n3750 , n1705 );
and ( n3752 , n3748 , n3751 );
and ( n3753 , n2289 , n1760 );
and ( n3754 , n2068 , n1758 );
nor ( n3755 , n3753 , n3754 );
xnor ( n3756 , n3755 , n1705 );
and ( n3757 , n3752 , n3756 );
xor ( n3758 , n3694 , n3698 );
xor ( n3759 , n3758 , n3561 );
and ( n3760 , n3756 , n3759 );
and ( n3761 , n3752 , n3759 );
or ( n3762 , n3757 , n3760 , n3761 );
and ( n3763 , n3744 , n3762 );
xor ( n3764 , n3690 , n3702 );
xor ( n3765 , n3764 , n3705 );
and ( n3766 , n3762 , n3765 );
and ( n3767 , n3744 , n3765 );
or ( n3768 , n3763 , n3766 , n3767 );
xor ( n3769 , n3620 , n3622 );
xor ( n3770 , n3769 , n3625 );
and ( n3771 , n3768 , n3770 );
xor ( n3772 , n3689 , n3708 );
xor ( n3773 , n3772 , n3711 );
and ( n3774 , n3770 , n3773 );
and ( n3775 , n3768 , n3773 );
or ( n3776 , n3771 , n3774 , n3775 );
and ( n3777 , n3726 , n3776 );
xor ( n3778 , n3726 , n3776 );
xor ( n3779 , n3730 , n3733 );
and ( n3780 , n2015 , n1866 );
and ( n3781 , n1833 , n1864 );
nor ( n3782 , n3780 , n3781 );
xnor ( n3783 , n3782 , n1844 );
and ( n3784 , n3779 , n3783 );
and ( n3785 , n2199 , n1652 );
and ( n3786 , n2158 , n1650 );
nor ( n3787 , n3785 , n3786 );
xnor ( n3788 , n3787 , n1597 );
and ( n3789 , n3783 , n3788 );
and ( n3790 , n3779 , n3788 );
or ( n3791 , n3784 , n3789 , n3790 );
xor ( n3792 , n3748 , n3751 );
and ( n3793 , n2068 , n1948 );
and ( n3794 , n1915 , n1946 );
nor ( n3795 , n3793 , n3794 );
xnor ( n3796 , n3795 , n1926 );
and ( n3797 , n3792 , n3796 );
and ( n3798 , n2346 , n1760 );
and ( n3799 , n2289 , n1758 );
nor ( n3800 , n3798 , n3799 );
xnor ( n3801 , n3800 , n1705 );
and ( n3802 , n3796 , n3801 );
and ( n3803 , n3792 , n3801 );
or ( n3804 , n3797 , n3802 , n3803 );
and ( n3805 , n3791 , n3804 );
xor ( n3806 , n3752 , n3756 );
xor ( n3807 , n3806 , n3759 );
and ( n3808 , n3804 , n3807 );
and ( n3809 , n3791 , n3807 );
or ( n3810 , n3805 , n3808 , n3809 );
xor ( n3811 , n3671 , n3683 );
xor ( n3812 , n3811 , n3686 );
and ( n3813 , n3810 , n3812 );
xor ( n3814 , n3744 , n3762 );
xor ( n3815 , n3814 , n3765 );
and ( n3816 , n3812 , n3815 );
and ( n3817 , n3810 , n3815 );
or ( n3818 , n3813 , n3816 , n3817 );
xor ( n3819 , n3768 , n3770 );
xor ( n3820 , n3819 , n3773 );
and ( n3821 , n3818 , n3820 );
xor ( n3822 , n3818 , n3820 );
xor ( n3823 , n3810 , n3812 );
xor ( n3824 , n3823 , n3815 );
and ( n3825 , n1833 , n2189 );
and ( n3826 , n1674 , n2186 );
nor ( n3827 , n3825 , n3826 );
xnor ( n3828 , n3827 , n1841 );
and ( n3829 , n2158 , n1866 );
and ( n3830 , n2015 , n1864 );
nor ( n3831 , n3829 , n3830 );
xnor ( n3832 , n3831 , n1844 );
and ( n3833 , n3828 , n3832 );
and ( n3834 , n3832 , n3731 );
and ( n3835 , n3828 , n3731 );
or ( n3836 , n3833 , n3834 , n3835 );
and ( n3837 , n1915 , n2336 );
and ( n3838 , n1782 , n2333 );
nor ( n3839 , n3837 , n3838 );
xnor ( n3840 , n3839 , n1923 );
and ( n3841 , n2289 , n1948 );
and ( n3842 , n2068 , n1946 );
nor ( n3843 , n3841 , n3842 );
xnor ( n3844 , n3843 , n1926 );
and ( n3845 , n3840 , n3844 );
and ( n3846 , n3844 , n3749 );
and ( n3847 , n3840 , n3749 );
or ( n3848 , n3845 , n3846 , n3847 );
and ( n3849 , n3836 , n3848 );
xor ( n3850 , n3792 , n3796 );
xor ( n3851 , n3850 , n3801 );
and ( n3852 , n3848 , n3851 );
and ( n3853 , n3836 , n3851 );
or ( n3854 , n3849 , n3852 , n3853 );
xor ( n3855 , n3734 , n3738 );
xor ( n3856 , n3855 , n3741 );
and ( n3857 , n3854 , n3856 );
xor ( n3858 , n3791 , n3804 );
xor ( n3859 , n3858 , n3807 );
and ( n3860 , n3856 , n3859 );
and ( n3861 , n3854 , n3859 );
or ( n3862 , n3857 , n3860 , n3861 );
and ( n3863 , n3824 , n3862 );
xor ( n3864 , n3824 , n3862 );
xor ( n3865 , n3854 , n3856 );
xor ( n3866 , n3865 , n3859 );
and ( n3867 , n2068 , n2336 );
and ( n3868 , n1915 , n2333 );
nor ( n3869 , n3867 , n3868 );
xnor ( n3870 , n3869 , n1923 );
and ( n3871 , n2346 , n1946 );
not ( n3872 , n3871 );
and ( n3873 , n3872 , n1926 );
and ( n3874 , n3870 , n3873 );
and ( n3875 , n2015 , n2189 );
and ( n3876 , n1833 , n2186 );
nor ( n3877 , n3875 , n3876 );
xnor ( n3878 , n3877 , n1841 );
and ( n3879 , n2199 , n1864 );
not ( n3880 , n3879 );
and ( n3881 , n3880 , n1844 );
and ( n3882 , n3878 , n3881 );
and ( n3883 , n3874 , n3882 );
xor ( n3884 , n3840 , n3844 );
xor ( n3885 , n3884 , n3749 );
and ( n3886 , n3882 , n3885 );
and ( n3887 , n3874 , n3885 );
or ( n3888 , n3883 , n3886 , n3887 );
xor ( n3889 , n3779 , n3783 );
xor ( n3890 , n3889 , n3788 );
and ( n3891 , n3888 , n3890 );
xor ( n3892 , n3836 , n3848 );
xor ( n3893 , n3892 , n3851 );
and ( n3894 , n3890 , n3893 );
and ( n3895 , n3888 , n3893 );
or ( n3896 , n3891 , n3894 , n3895 );
and ( n3897 , n3866 , n3896 );
xor ( n3898 , n3866 , n3896 );
xor ( n3899 , n3870 , n3873 );
and ( n3900 , n2199 , n1866 );
and ( n3901 , n2158 , n1864 );
nor ( n3902 , n3900 , n3901 );
xnor ( n3903 , n3902 , n1844 );
and ( n3904 , n3899 , n3903 );
and ( n3905 , n2346 , n1948 );
and ( n3906 , n2289 , n1946 );
nor ( n3907 , n3905 , n3906 );
xnor ( n3908 , n3907 , n1926 );
and ( n3909 , n3903 , n3908 );
and ( n3910 , n3899 , n3908 );
or ( n3911 , n3904 , n3909 , n3910 );
xor ( n3912 , n3828 , n3832 );
xor ( n3913 , n3912 , n3731 );
and ( n3914 , n3911 , n3913 );
xor ( n3915 , n3874 , n3882 );
xor ( n3916 , n3915 , n3885 );
and ( n3917 , n3913 , n3916 );
and ( n3918 , n3911 , n3916 );
or ( n3919 , n3914 , n3917 , n3918 );
xor ( n3920 , n3888 , n3890 );
xor ( n3921 , n3920 , n3893 );
and ( n3922 , n3919 , n3921 );
xor ( n3923 , n3919 , n3921 );
xor ( n3924 , n3911 , n3913 );
xor ( n3925 , n3924 , n3916 );
xor ( n3926 , n3878 , n3881 );
and ( n3927 , n2289 , n2336 );
and ( n3928 , n2068 , n2333 );
nor ( n3929 , n3927 , n3928 );
xnor ( n3930 , n3929 , n1923 );
and ( n3931 , n3879 , n3930 );
and ( n3932 , n3926 , n3931 );
xor ( n3933 , n3899 , n3903 );
xor ( n3934 , n3933 , n3908 );
and ( n3935 , n3931 , n3934 );
and ( n3936 , n3926 , n3934 );
or ( n3937 , n3932 , n3935 , n3936 );
and ( n3938 , n3925 , n3937 );
xor ( n3939 , n3925 , n3937 );
xor ( n3940 , n3879 , n3930 );
and ( n3941 , n2158 , n2189 );
and ( n3942 , n2015 , n2186 );
nor ( n3943 , n3941 , n3942 );
xnor ( n3944 , n3943 , n1841 );
and ( n3945 , n3940 , n3944 );
and ( n3946 , n3944 , n3871 );
and ( n3947 , n3940 , n3871 );
or ( n3948 , n3945 , n3946 , n3947 );
xor ( n3949 , n3926 , n3931 );
xor ( n3950 , n3949 , n3934 );
and ( n3951 , n3948 , n3950 );
xor ( n3952 , n3948 , n3950 );
and ( n3953 , n2199 , n2186 );
not ( n3954 , n3953 );
and ( n3955 , n3954 , n1841 );
and ( n3956 , n2346 , n2333 );
not ( n3957 , n3956 );
and ( n3958 , n3957 , n1923 );
and ( n3959 , n3955 , n3958 );
and ( n3960 , n2346 , n2336 );
and ( n3961 , n2289 , n2333 );
nor ( n3962 , n3960 , n3961 );
xnor ( n3963 , n3962 , n1923 );
and ( n3964 , n3958 , n3963 );
and ( n3965 , n3955 , n3963 );
or ( n3966 , n3959 , n3964 , n3965 );
xor ( n3967 , n3940 , n3944 );
xor ( n3968 , n3967 , n3871 );
and ( n3969 , n3966 , n3968 );
xor ( n3970 , n3966 , n3968 );
and ( n3971 , n2199 , n2189 );
and ( n3972 , n2158 , n2186 );
nor ( n3973 , n3971 , n3972 );
xnor ( n3974 , n3973 , n1841 );
xor ( n3975 , n3955 , n3958 );
xor ( n3976 , n3975 , n3963 );
and ( n3977 , n3974 , n3976 );
xor ( n3978 , n3974 , n3976 );
and ( n3979 , n3953 , n3956 );
and ( n3980 , n3978 , n3979 );
or ( n3981 , n3977 , n3980 );
and ( n3982 , n3970 , n3981 );
or ( n3983 , n3969 , n3982 );
and ( n3984 , n3952 , n3983 );
or ( n3985 , n3951 , n3984 );
and ( n3986 , n3939 , n3985 );
or ( n3987 , n3938 , n3986 );
and ( n3988 , n3923 , n3987 );
or ( n3989 , n3922 , n3988 );
and ( n3990 , n3898 , n3989 );
or ( n3991 , n3897 , n3990 );
and ( n3992 , n3864 , n3991 );
or ( n3993 , n3863 , n3992 );
and ( n3994 , n3822 , n3993 );
or ( n3995 , n3821 , n3994 );
and ( n3996 , n3778 , n3995 );
or ( n3997 , n3777 , n3996 );
and ( n3998 , n3724 , n3997 );
or ( n3999 , n3723 , n3998 );
and ( n4000 , n3668 , n3999 );
or ( n4001 , n3667 , n4000 );
and ( n4002 , n3602 , n4001 );
or ( n4003 , n3601 , n4002 );
and ( n4004 , n3528 , n4003 );
or ( n4005 , n3527 , n4004 );
and ( n4006 , n3452 , n4005 );
or ( n4007 , n3451 , n4006 );
and ( n4008 , n3358 , n4007 );
or ( n4009 , n3357 , n4008 );
and ( n4010 , n3256 , n4009 );
or ( n4011 , n3255 , n4010 );
and ( n4012 , n3180 , n4011 );
or ( n4013 , n3179 , n4012 );
and ( n4014 , n3066 , n4013 );
or ( n4015 , n3065 , n4014 );
and ( n4016 , n2950 , n4015 );
or ( n4017 , n2949 , n4016 );
and ( n4018 , n2788 , n4017 );
or ( n4019 , n2787 , n4018 );
and ( n4020 , n2652 , n4019 );
or ( n4021 , n2651 , n4020 );
and ( n4022 , n2582 , n4021 );
or ( n4023 , n2581 , n4022 );
and ( n4024 , n2406 , n4023 );
or ( n4025 , n2405 , n4024 );
and ( n4026 , n2126 , n4025 );
or ( n4027 , n2125 , n4026 );
and ( n4028 , n2002 , n4027 );
or ( n4029 , n2001 , n4028 );
and ( n4030 , n1820 , n4029 );
or ( n4031 , n1819 , n4030 );
and ( n4032 , n1532 , n4031 );
or ( n4033 , n1531 , n4032 );
and ( n4034 , n1400 , n4033 );
or ( n4035 , n1399 , n4034 );
and ( n4036 , n1276 , n4035 );
or ( n4037 , n1275 , n4036 );
and ( n4038 , n1175 , n4037 );
or ( n4039 , n1174 , n4038 );
xor ( n4040 , n1066 , n4039 );
buf ( n4041 , n4040 );
buf ( n4042 , n4041 );
buf ( n4043 , n560 );
buf ( n4044 , n576 );
and ( n4045 , n4043 , n4044 );
buf ( n4046 , n561 );
buf ( n4047 , n577 );
and ( n4048 , n4046 , n4047 );
buf ( n4049 , n562 );
buf ( n4050 , n578 );
and ( n4051 , n4049 , n4050 );
buf ( n4052 , n563 );
buf ( n4053 , n579 );
and ( n4054 , n4052 , n4053 );
buf ( n4055 , n564 );
buf ( n4056 , n580 );
and ( n4057 , n4055 , n4056 );
buf ( n4058 , n565 );
buf ( n4059 , n581 );
and ( n4060 , n4058 , n4059 );
buf ( n4061 , n566 );
buf ( n4062 , n582 );
and ( n4063 , n4061 , n4062 );
buf ( n4064 , n567 );
buf ( n4065 , n583 );
and ( n4066 , n4064 , n4065 );
buf ( n4067 , n568 );
buf ( n4068 , n584 );
and ( n4069 , n4067 , n4068 );
buf ( n4070 , n569 );
buf ( n4071 , n585 );
and ( n4072 , n4070 , n4071 );
buf ( n4073 , n570 );
buf ( n4074 , n586 );
and ( n4075 , n4073 , n4074 );
buf ( n4076 , n571 );
buf ( n4077 , n587 );
and ( n4078 , n4076 , n4077 );
buf ( n4079 , n572 );
buf ( n4080 , n588 );
and ( n4081 , n4079 , n4080 );
buf ( n4082 , n573 );
buf ( n4083 , n589 );
and ( n4084 , n4082 , n4083 );
buf ( n4085 , n574 );
buf ( n4086 , n590 );
and ( n4087 , n4085 , n4086 );
buf ( n4088 , n575 );
buf ( n4089 , n591 );
and ( n4090 , n4088 , n4089 );
and ( n4091 , n4086 , n4090 );
and ( n4092 , n4085 , n4090 );
or ( n4093 , n4087 , n4091 , n4092 );
and ( n4094 , n4083 , n4093 );
and ( n4095 , n4082 , n4093 );
or ( n4096 , n4084 , n4094 , n4095 );
and ( n4097 , n4080 , n4096 );
and ( n4098 , n4079 , n4096 );
or ( n4099 , n4081 , n4097 , n4098 );
and ( n4100 , n4077 , n4099 );
and ( n4101 , n4076 , n4099 );
or ( n4102 , n4078 , n4100 , n4101 );
and ( n4103 , n4074 , n4102 );
and ( n4104 , n4073 , n4102 );
or ( n4105 , n4075 , n4103 , n4104 );
and ( n4106 , n4071 , n4105 );
and ( n4107 , n4070 , n4105 );
or ( n4108 , n4072 , n4106 , n4107 );
and ( n4109 , n4068 , n4108 );
and ( n4110 , n4067 , n4108 );
or ( n4111 , n4069 , n4109 , n4110 );
and ( n4112 , n4065 , n4111 );
and ( n4113 , n4064 , n4111 );
or ( n4114 , n4066 , n4112 , n4113 );
and ( n4115 , n4062 , n4114 );
and ( n4116 , n4061 , n4114 );
or ( n4117 , n4063 , n4115 , n4116 );
and ( n4118 , n4059 , n4117 );
and ( n4119 , n4058 , n4117 );
or ( n4120 , n4060 , n4118 , n4119 );
and ( n4121 , n4056 , n4120 );
and ( n4122 , n4055 , n4120 );
or ( n4123 , n4057 , n4121 , n4122 );
and ( n4124 , n4053 , n4123 );
and ( n4125 , n4052 , n4123 );
or ( n4126 , n4054 , n4124 , n4125 );
and ( n4127 , n4050 , n4126 );
and ( n4128 , n4049 , n4126 );
or ( n4129 , n4051 , n4127 , n4128 );
and ( n4130 , n4047 , n4129 );
and ( n4131 , n4046 , n4129 );
or ( n4132 , n4048 , n4130 , n4131 );
and ( n4133 , n4044 , n4132 );
and ( n4134 , n4043 , n4132 );
or ( n4135 , n4045 , n4133 , n4134 );
buf ( n4136 , n4135 );
buf ( n4137 , n4136 );
buf ( n4138 , n4137 );
buf ( n4139 , n546 );
buf ( n4140 , n4139 );
buf ( n4141 , n547 );
buf ( n4142 , n4141 );
xor ( n4143 , n4140 , n4142 );
buf ( n4144 , n548 );
buf ( n4145 , n4144 );
xor ( n4146 , n4142 , n4145 );
not ( n4147 , n4146 );
and ( n4148 , n4143 , n4147 );
and ( n4149 , n4138 , n4148 );
not ( n4150 , n4149 );
and ( n4151 , n4142 , n4145 );
not ( n4152 , n4151 );
and ( n4153 , n4140 , n4152 );
xnor ( n4154 , n4150 , n4153 );
buf ( n4155 , n4154 );
not ( n4156 , n4153 );
and ( n4157 , n4155 , n4156 );
xor ( n4158 , n4043 , n4044 );
xor ( n4159 , n4158 , n4132 );
buf ( n4160 , n4159 );
buf ( n4161 , n4160 );
buf ( n4162 , n4161 );
buf ( n4163 , n544 );
buf ( n4164 , n4163 );
buf ( n4165 , n545 );
buf ( n4166 , n4165 );
xor ( n4167 , n4164 , n4166 );
xor ( n4168 , n4166 , n4140 );
not ( n4169 , n4168 );
and ( n4170 , n4167 , n4169 );
and ( n4171 , n4162 , n4170 );
and ( n4172 , n4138 , n4168 );
nor ( n4173 , n4171 , n4172 );
and ( n4174 , n4166 , n4140 );
not ( n4175 , n4174 );
and ( n4176 , n4164 , n4175 );
xnor ( n4177 , n4173 , n4176 );
and ( n4178 , n4156 , n4177 );
and ( n4179 , n4155 , n4177 );
or ( n4180 , n4157 , n4178 , n4179 );
and ( n4181 , n4138 , n4170 );
not ( n4182 , n4181 );
xnor ( n4183 , n4182 , n4176 );
xor ( n4184 , n4180 , n4183 );
and ( n4185 , n4162 , n4164 );
xor ( n4186 , n4184 , n4185 );
not ( n4187 , n4154 );
xor ( n4188 , n4046 , n4047 );
xor ( n4189 , n4188 , n4129 );
buf ( n4190 , n4189 );
buf ( n4191 , n4190 );
buf ( n4192 , n4191 );
and ( n4193 , n4192 , n4170 );
and ( n4194 , n4162 , n4168 );
nor ( n4195 , n4193 , n4194 );
xnor ( n4196 , n4195 , n4176 );
and ( n4197 , n4187 , n4196 );
xor ( n4198 , n4049 , n4050 );
xor ( n4199 , n4198 , n4126 );
buf ( n4200 , n4199 );
buf ( n4201 , n4200 );
buf ( n4202 , n4201 );
and ( n4203 , n4202 , n4164 );
and ( n4204 , n4196 , n4203 );
and ( n4205 , n4187 , n4203 );
or ( n4206 , n4197 , n4204 , n4205 );
and ( n4207 , n4192 , n4164 );
and ( n4208 , n4206 , n4207 );
xor ( n4209 , n4155 , n4156 );
xor ( n4210 , n4209 , n4177 );
and ( n4211 , n4207 , n4210 );
and ( n4212 , n4206 , n4210 );
or ( n4213 , n4208 , n4211 , n4212 );
xor ( n4214 , n4186 , n4213 );
xor ( n4215 , n4206 , n4207 );
xor ( n4216 , n4215 , n4210 );
buf ( n4217 , n549 );
buf ( n4218 , n4217 );
buf ( n4219 , n550 );
buf ( n4220 , n4219 );
and ( n4221 , n4218 , n4220 );
not ( n4222 , n4221 );
and ( n4223 , n4145 , n4222 );
not ( n4224 , n4223 );
and ( n4225 , n4162 , n4148 );
and ( n4226 , n4138 , n4146 );
nor ( n4227 , n4225 , n4226 );
xnor ( n4228 , n4227 , n4153 );
and ( n4229 , n4224 , n4228 );
xor ( n4230 , n4052 , n4053 );
xor ( n4231 , n4230 , n4123 );
buf ( n4232 , n4231 );
buf ( n4233 , n4232 );
buf ( n4234 , n4233 );
and ( n4235 , n4234 , n4164 );
and ( n4236 , n4228 , n4235 );
and ( n4237 , n4224 , n4235 );
or ( n4238 , n4229 , n4236 , n4237 );
xor ( n4239 , n4145 , n4218 );
xor ( n4240 , n4218 , n4220 );
not ( n4241 , n4240 );
and ( n4242 , n4239 , n4241 );
and ( n4243 , n4138 , n4242 );
not ( n4244 , n4243 );
xnor ( n4245 , n4244 , n4223 );
not ( n4246 , n4245 );
and ( n4247 , n4192 , n4148 );
and ( n4248 , n4162 , n4146 );
nor ( n4249 , n4247 , n4248 );
xnor ( n4250 , n4249 , n4153 );
and ( n4251 , n4246 , n4250 );
xor ( n4252 , n4055 , n4056 );
xor ( n4253 , n4252 , n4120 );
buf ( n4254 , n4253 );
buf ( n4255 , n4254 );
buf ( n4256 , n4255 );
and ( n4257 , n4256 , n4164 );
and ( n4258 , n4250 , n4257 );
and ( n4259 , n4246 , n4257 );
or ( n4260 , n4251 , n4258 , n4259 );
buf ( n4261 , n4245 );
and ( n4262 , n4260 , n4261 );
and ( n4263 , n4202 , n4170 );
and ( n4264 , n4192 , n4168 );
nor ( n4265 , n4263 , n4264 );
xnor ( n4266 , n4265 , n4176 );
and ( n4267 , n4261 , n4266 );
and ( n4268 , n4260 , n4266 );
or ( n4269 , n4262 , n4267 , n4268 );
and ( n4270 , n4238 , n4269 );
xor ( n4271 , n4187 , n4196 );
xor ( n4272 , n4271 , n4203 );
and ( n4273 , n4269 , n4272 );
and ( n4274 , n4238 , n4272 );
or ( n4275 , n4270 , n4273 , n4274 );
and ( n4276 , n4216 , n4275 );
xor ( n4277 , n4238 , n4269 );
xor ( n4278 , n4277 , n4272 );
buf ( n4279 , n551 );
buf ( n4280 , n4279 );
buf ( n4281 , n552 );
buf ( n4282 , n4281 );
and ( n4283 , n4280 , n4282 );
not ( n4284 , n4283 );
and ( n4285 , n4220 , n4284 );
not ( n4286 , n4285 );
and ( n4287 , n4162 , n4242 );
and ( n4288 , n4138 , n4240 );
nor ( n4289 , n4287 , n4288 );
xnor ( n4290 , n4289 , n4223 );
and ( n4291 , n4286 , n4290 );
and ( n4292 , n4256 , n4170 );
and ( n4293 , n4234 , n4168 );
nor ( n4294 , n4292 , n4293 );
xnor ( n4295 , n4294 , n4176 );
and ( n4296 , n4290 , n4295 );
and ( n4297 , n4286 , n4295 );
or ( n4298 , n4291 , n4296 , n4297 );
xor ( n4299 , n4220 , n4280 );
xor ( n4300 , n4280 , n4282 );
not ( n4301 , n4300 );
and ( n4302 , n4299 , n4301 );
and ( n4303 , n4138 , n4302 );
not ( n4304 , n4303 );
xnor ( n4305 , n4304 , n4285 );
buf ( n4306 , n4305 );
and ( n4307 , n4202 , n4148 );
and ( n4308 , n4192 , n4146 );
nor ( n4309 , n4307 , n4308 );
xnor ( n4310 , n4309 , n4153 );
and ( n4311 , n4306 , n4310 );
xor ( n4312 , n4058 , n4059 );
xor ( n4313 , n4312 , n4117 );
buf ( n4314 , n4313 );
buf ( n4315 , n4314 );
buf ( n4316 , n4315 );
and ( n4317 , n4316 , n4164 );
and ( n4318 , n4310 , n4317 );
and ( n4319 , n4306 , n4317 );
or ( n4320 , n4311 , n4318 , n4319 );
and ( n4321 , n4298 , n4320 );
and ( n4322 , n4234 , n4170 );
and ( n4323 , n4202 , n4168 );
nor ( n4324 , n4322 , n4323 );
xnor ( n4325 , n4324 , n4176 );
and ( n4326 , n4320 , n4325 );
and ( n4327 , n4298 , n4325 );
or ( n4328 , n4321 , n4326 , n4327 );
xor ( n4329 , n4224 , n4228 );
xor ( n4330 , n4329 , n4235 );
and ( n4331 , n4328 , n4330 );
xor ( n4332 , n4260 , n4261 );
xor ( n4333 , n4332 , n4266 );
and ( n4334 , n4330 , n4333 );
and ( n4335 , n4328 , n4333 );
or ( n4336 , n4331 , n4334 , n4335 );
and ( n4337 , n4278 , n4336 );
xor ( n4338 , n4328 , n4330 );
xor ( n4339 , n4338 , n4333 );
not ( n4340 , n4305 );
and ( n4341 , n4192 , n4242 );
and ( n4342 , n4162 , n4240 );
nor ( n4343 , n4341 , n4342 );
xnor ( n4344 , n4343 , n4223 );
and ( n4345 , n4340 , n4344 );
and ( n4346 , n4316 , n4170 );
and ( n4347 , n4256 , n4168 );
nor ( n4348 , n4346 , n4347 );
xnor ( n4349 , n4348 , n4176 );
and ( n4350 , n4344 , n4349 );
and ( n4351 , n4340 , n4349 );
or ( n4352 , n4345 , n4350 , n4351 );
xor ( n4353 , n4286 , n4290 );
xor ( n4354 , n4353 , n4295 );
and ( n4355 , n4352 , n4354 );
xor ( n4356 , n4306 , n4310 );
xor ( n4357 , n4356 , n4317 );
and ( n4358 , n4354 , n4357 );
and ( n4359 , n4352 , n4357 );
or ( n4360 , n4355 , n4358 , n4359 );
xor ( n4361 , n4298 , n4320 );
xor ( n4362 , n4361 , n4325 );
and ( n4363 , n4360 , n4362 );
xor ( n4364 , n4246 , n4250 );
xor ( n4365 , n4364 , n4257 );
and ( n4366 , n4362 , n4365 );
and ( n4367 , n4360 , n4365 );
or ( n4368 , n4363 , n4366 , n4367 );
and ( n4369 , n4339 , n4368 );
xor ( n4370 , n4360 , n4362 );
xor ( n4371 , n4370 , n4365 );
and ( n4372 , n4202 , n4242 );
and ( n4373 , n4192 , n4240 );
nor ( n4374 , n4372 , n4373 );
xnor ( n4375 , n4374 , n4223 );
and ( n4376 , n4256 , n4148 );
and ( n4377 , n4234 , n4146 );
nor ( n4378 , n4376 , n4377 );
xnor ( n4379 , n4378 , n4153 );
and ( n4380 , n4375 , n4379 );
xor ( n4381 , n4061 , n4062 );
xor ( n4382 , n4381 , n4114 );
buf ( n4383 , n4382 );
buf ( n4384 , n4383 );
buf ( n4385 , n4384 );
and ( n4386 , n4385 , n4170 );
and ( n4387 , n4316 , n4168 );
nor ( n4388 , n4386 , n4387 );
xnor ( n4389 , n4388 , n4176 );
and ( n4390 , n4379 , n4389 );
and ( n4391 , n4375 , n4389 );
or ( n4392 , n4380 , n4390 , n4391 );
and ( n4393 , n4234 , n4148 );
and ( n4394 , n4202 , n4146 );
nor ( n4395 , n4393 , n4394 );
xnor ( n4396 , n4395 , n4153 );
and ( n4397 , n4392 , n4396 );
and ( n4398 , n4385 , n4164 );
and ( n4399 , n4396 , n4398 );
and ( n4400 , n4392 , n4398 );
or ( n4401 , n4397 , n4399 , n4400 );
buf ( n4402 , n553 );
buf ( n4403 , n4402 );
buf ( n4404 , n554 );
buf ( n4405 , n4404 );
and ( n4406 , n4403 , n4405 );
not ( n4407 , n4406 );
and ( n4408 , n4282 , n4407 );
not ( n4409 , n4408 );
and ( n4410 , n4162 , n4302 );
and ( n4411 , n4138 , n4300 );
nor ( n4412 , n4410 , n4411 );
xnor ( n4413 , n4412 , n4285 );
and ( n4414 , n4409 , n4413 );
xor ( n4415 , n4064 , n4065 );
xor ( n4416 , n4415 , n4111 );
buf ( n4417 , n4416 );
buf ( n4418 , n4417 );
buf ( n4419 , n4418 );
and ( n4420 , n4419 , n4164 );
and ( n4421 , n4413 , n4420 );
and ( n4422 , n4409 , n4420 );
or ( n4423 , n4414 , n4421 , n4422 );
and ( n4424 , n4192 , n4302 );
and ( n4425 , n4162 , n4300 );
nor ( n4426 , n4424 , n4425 );
xnor ( n4427 , n4426 , n4285 );
and ( n4428 , n4316 , n4148 );
and ( n4429 , n4256 , n4146 );
nor ( n4430 , n4428 , n4429 );
xnor ( n4431 , n4430 , n4153 );
and ( n4432 , n4427 , n4431 );
xor ( n4433 , n4067 , n4068 );
xor ( n4434 , n4433 , n4108 );
buf ( n4435 , n4434 );
buf ( n4436 , n4435 );
buf ( n4437 , n4436 );
and ( n4438 , n4437 , n4164 );
and ( n4439 , n4431 , n4438 );
and ( n4440 , n4427 , n4438 );
or ( n4441 , n4432 , n4439 , n4440 );
xor ( n4442 , n4282 , n4403 );
xor ( n4443 , n4403 , n4405 );
not ( n4444 , n4443 );
and ( n4445 , n4442 , n4444 );
and ( n4446 , n4138 , n4445 );
not ( n4447 , n4446 );
xnor ( n4448 , n4447 , n4408 );
not ( n4449 , n4448 );
and ( n4450 , n4234 , n4242 );
and ( n4451 , n4202 , n4240 );
nor ( n4452 , n4450 , n4451 );
xnor ( n4453 , n4452 , n4223 );
and ( n4454 , n4449 , n4453 );
and ( n4455 , n4419 , n4170 );
and ( n4456 , n4385 , n4168 );
nor ( n4457 , n4455 , n4456 );
xnor ( n4458 , n4457 , n4176 );
and ( n4459 , n4453 , n4458 );
and ( n4460 , n4449 , n4458 );
or ( n4461 , n4454 , n4459 , n4460 );
and ( n4462 , n4441 , n4461 );
buf ( n4463 , n4448 );
and ( n4464 , n4461 , n4463 );
and ( n4465 , n4441 , n4463 );
or ( n4466 , n4462 , n4464 , n4465 );
and ( n4467 , n4423 , n4466 );
xor ( n4468 , n4340 , n4344 );
xor ( n4469 , n4468 , n4349 );
and ( n4470 , n4466 , n4469 );
and ( n4471 , n4423 , n4469 );
or ( n4472 , n4467 , n4470 , n4471 );
and ( n4473 , n4401 , n4472 );
xor ( n4474 , n4352 , n4354 );
xor ( n4475 , n4474 , n4357 );
and ( n4476 , n4472 , n4475 );
and ( n4477 , n4401 , n4475 );
or ( n4478 , n4473 , n4476 , n4477 );
and ( n4479 , n4371 , n4478 );
xor ( n4480 , n4401 , n4472 );
xor ( n4481 , n4480 , n4475 );
xor ( n4482 , n4409 , n4413 );
xor ( n4483 , n4482 , n4420 );
xor ( n4484 , n4375 , n4379 );
xor ( n4485 , n4484 , n4389 );
and ( n4486 , n4483 , n4485 );
xor ( n4487 , n4441 , n4461 );
xor ( n4488 , n4487 , n4463 );
and ( n4489 , n4485 , n4488 );
and ( n4490 , n4483 , n4488 );
or ( n4491 , n4486 , n4489 , n4490 );
xor ( n4492 , n4392 , n4396 );
xor ( n4493 , n4492 , n4398 );
and ( n4494 , n4491 , n4493 );
xor ( n4495 , n4423 , n4466 );
xor ( n4496 , n4495 , n4469 );
and ( n4497 , n4493 , n4496 );
and ( n4498 , n4491 , n4496 );
or ( n4499 , n4494 , n4497 , n4498 );
and ( n4500 , n4481 , n4499 );
xor ( n4501 , n4491 , n4493 );
xor ( n4502 , n4501 , n4496 );
xor ( n4503 , n4483 , n4485 );
xor ( n4504 , n4503 , n4488 );
and ( n4505 , n4192 , n4445 );
and ( n4506 , n4162 , n4443 );
nor ( n4507 , n4505 , n4506 );
xnor ( n4508 , n4507 , n4408 );
xor ( n4509 , n4070 , n4071 );
xor ( n4510 , n4509 , n4105 );
buf ( n4511 , n4510 );
buf ( n4512 , n4511 );
buf ( n4513 , n4512 );
and ( n4514 , n4513 , n4170 );
and ( n4515 , n4437 , n4168 );
nor ( n4516 , n4514 , n4515 );
xnor ( n4517 , n4516 , n4176 );
and ( n4518 , n4508 , n4517 );
xor ( n4519 , n4073 , n4074 );
xor ( n4520 , n4519 , n4102 );
buf ( n4521 , n4520 );
buf ( n4522 , n4521 );
buf ( n4523 , n4522 );
and ( n4524 , n4523 , n4164 );
and ( n4525 , n4517 , n4524 );
and ( n4526 , n4508 , n4524 );
or ( n4527 , n4518 , n4525 , n4526 );
and ( n4528 , n4202 , n4302 );
and ( n4529 , n4192 , n4300 );
nor ( n4530 , n4528 , n4529 );
xnor ( n4531 , n4530 , n4285 );
and ( n4532 , n4527 , n4531 );
and ( n4533 , n4385 , n4148 );
and ( n4534 , n4316 , n4146 );
nor ( n4535 , n4533 , n4534 );
xnor ( n4536 , n4535 , n4153 );
and ( n4537 , n4531 , n4536 );
and ( n4538 , n4527 , n4536 );
or ( n4539 , n4532 , n4537 , n4538 );
xor ( n4540 , n4427 , n4431 );
xor ( n4541 , n4540 , n4438 );
and ( n4542 , n4539 , n4541 );
and ( n4543 , n4504 , n4542 );
xor ( n4544 , n4449 , n4453 );
xor ( n4545 , n4544 , n4458 );
buf ( n4546 , n555 );
buf ( n4547 , n4546 );
buf ( n4548 , n556 );
buf ( n4549 , n4548 );
and ( n4550 , n4547 , n4549 );
not ( n4551 , n4550 );
and ( n4552 , n4405 , n4551 );
not ( n4553 , n4552 );
and ( n4554 , n4437 , n4170 );
and ( n4555 , n4419 , n4168 );
nor ( n4556 , n4554 , n4555 );
xnor ( n4557 , n4556 , n4176 );
and ( n4558 , n4553 , n4557 );
and ( n4559 , n4513 , n4164 );
and ( n4560 , n4557 , n4559 );
and ( n4561 , n4553 , n4559 );
or ( n4562 , n4558 , n4560 , n4561 );
and ( n4563 , n4545 , n4562 );
and ( n4564 , n4162 , n4445 );
and ( n4565 , n4138 , n4443 );
nor ( n4566 , n4564 , n4565 );
xnor ( n4567 , n4566 , n4408 );
and ( n4568 , n4256 , n4242 );
and ( n4569 , n4234 , n4240 );
nor ( n4570 , n4568 , n4569 );
xnor ( n4571 , n4570 , n4223 );
and ( n4572 , n4567 , n4571 );
xor ( n4573 , n4553 , n4557 );
xor ( n4574 , n4573 , n4559 );
and ( n4575 , n4571 , n4574 );
and ( n4576 , n4567 , n4574 );
or ( n4577 , n4572 , n4575 , n4576 );
and ( n4578 , n4562 , n4577 );
and ( n4579 , n4545 , n4577 );
or ( n4580 , n4563 , n4578 , n4579 );
and ( n4581 , n4542 , n4580 );
and ( n4582 , n4504 , n4580 );
or ( n4583 , n4543 , n4581 , n4582 );
and ( n4584 , n4502 , n4583 );
xor ( n4585 , n4539 , n4541 );
and ( n4586 , n4234 , n4302 );
and ( n4587 , n4202 , n4300 );
nor ( n4588 , n4586 , n4587 );
xnor ( n4589 , n4588 , n4285 );
and ( n4590 , n4316 , n4242 );
and ( n4591 , n4256 , n4240 );
nor ( n4592 , n4590 , n4591 );
xnor ( n4593 , n4592 , n4223 );
and ( n4594 , n4589 , n4593 );
and ( n4595 , n4419 , n4148 );
and ( n4596 , n4385 , n4146 );
nor ( n4597 , n4595 , n4596 );
xnor ( n4598 , n4597 , n4153 );
and ( n4599 , n4593 , n4598 );
and ( n4600 , n4589 , n4598 );
or ( n4601 , n4594 , n4599 , n4600 );
xor ( n4602 , n4405 , n4547 );
xor ( n4603 , n4547 , n4549 );
not ( n4604 , n4603 );
and ( n4605 , n4602 , n4604 );
and ( n4606 , n4162 , n4605 );
and ( n4607 , n4138 , n4603 );
nor ( n4608 , n4606 , n4607 );
xnor ( n4609 , n4608 , n4552 );
and ( n4610 , n4202 , n4445 );
and ( n4611 , n4192 , n4443 );
nor ( n4612 , n4610 , n4611 );
xnor ( n4613 , n4612 , n4408 );
and ( n4614 , n4609 , n4613 );
and ( n4615 , n4385 , n4242 );
and ( n4616 , n4316 , n4240 );
nor ( n4617 , n4615 , n4616 );
xnor ( n4618 , n4617 , n4223 );
and ( n4619 , n4613 , n4618 );
and ( n4620 , n4609 , n4618 );
or ( n4621 , n4614 , n4619 , n4620 );
xor ( n4622 , n4508 , n4517 );
xor ( n4623 , n4622 , n4524 );
and ( n4624 , n4621 , n4623 );
and ( n4625 , n4601 , n4624 );
xor ( n4626 , n4567 , n4571 );
xor ( n4627 , n4626 , n4574 );
and ( n4628 , n4624 , n4627 );
and ( n4629 , n4601 , n4627 );
or ( n4630 , n4625 , n4628 , n4629 );
and ( n4631 , n4585 , n4630 );
xor ( n4632 , n4545 , n4562 );
xor ( n4633 , n4632 , n4577 );
and ( n4634 , n4630 , n4633 );
and ( n4635 , n4585 , n4633 );
or ( n4636 , n4631 , n4634 , n4635 );
xor ( n4637 , n4504 , n4542 );
xor ( n4638 , n4637 , n4580 );
and ( n4639 , n4636 , n4638 );
xor ( n4640 , n4585 , n4630 );
xor ( n4641 , n4640 , n4633 );
and ( n4642 , n4256 , n4302 );
and ( n4643 , n4234 , n4300 );
nor ( n4644 , n4642 , n4643 );
xnor ( n4645 , n4644 , n4285 );
and ( n4646 , n4437 , n4148 );
and ( n4647 , n4419 , n4146 );
nor ( n4648 , n4646 , n4647 );
xnor ( n4649 , n4648 , n4153 );
and ( n4650 , n4645 , n4649 );
and ( n4651 , n4523 , n4170 );
and ( n4652 , n4513 , n4168 );
nor ( n4653 , n4651 , n4652 );
xnor ( n4654 , n4653 , n4176 );
and ( n4655 , n4649 , n4654 );
and ( n4656 , n4645 , n4654 );
or ( n4657 , n4650 , n4655 , n4656 );
xor ( n4658 , n4079 , n4080 );
xor ( n4659 , n4658 , n4096 );
buf ( n4660 , n4659 );
buf ( n4661 , n4660 );
buf ( n4662 , n4661 );
and ( n4663 , n4662 , n4164 );
buf ( n4664 , n4663 );
buf ( n4665 , n557 );
buf ( n4666 , n4665 );
buf ( n4667 , n558 );
buf ( n4668 , n4667 );
and ( n4669 , n4666 , n4668 );
not ( n4670 , n4669 );
and ( n4671 , n4549 , n4670 );
not ( n4672 , n4671 );
and ( n4673 , n4664 , n4672 );
xor ( n4674 , n4076 , n4077 );
xor ( n4675 , n4674 , n4099 );
buf ( n4676 , n4675 );
buf ( n4677 , n4676 );
buf ( n4678 , n4677 );
and ( n4679 , n4678 , n4164 );
and ( n4680 , n4672 , n4679 );
and ( n4681 , n4664 , n4679 );
or ( n4682 , n4673 , n4680 , n4681 );
and ( n4683 , n4657 , n4682 );
and ( n4684 , n4138 , n4605 );
not ( n4685 , n4684 );
xnor ( n4686 , n4685 , n4552 );
not ( n4687 , n4686 );
and ( n4688 , n4682 , n4687 );
and ( n4689 , n4657 , n4687 );
or ( n4690 , n4683 , n4688 , n4689 );
xor ( n4691 , n4527 , n4531 );
xor ( n4692 , n4691 , n4536 );
and ( n4693 , n4690 , n4692 );
and ( n4694 , n4641 , n4693 );
xor ( n4695 , n4601 , n4624 );
xor ( n4696 , n4695 , n4627 );
buf ( n4697 , n4686 );
and ( n4698 , n4696 , n4697 );
xor ( n4699 , n4690 , n4692 );
and ( n4700 , n4697 , n4699 );
and ( n4701 , n4696 , n4699 );
or ( n4702 , n4698 , n4700 , n4701 );
and ( n4703 , n4693 , n4702 );
and ( n4704 , n4641 , n4702 );
or ( n4705 , n4694 , n4703 , n4704 );
and ( n4706 , n4638 , n4705 );
and ( n4707 , n4636 , n4705 );
or ( n4708 , n4639 , n4706 , n4707 );
and ( n4709 , n4583 , n4708 );
and ( n4710 , n4502 , n4708 );
or ( n4711 , n4584 , n4709 , n4710 );
and ( n4712 , n4499 , n4711 );
and ( n4713 , n4481 , n4711 );
or ( n4714 , n4500 , n4712 , n4713 );
and ( n4715 , n4478 , n4714 );
and ( n4716 , n4371 , n4714 );
or ( n4717 , n4479 , n4715 , n4716 );
and ( n4718 , n4368 , n4717 );
and ( n4719 , n4339 , n4717 );
or ( n4720 , n4369 , n4718 , n4719 );
and ( n4721 , n4336 , n4720 );
and ( n4722 , n4278 , n4720 );
or ( n4723 , n4337 , n4721 , n4722 );
and ( n4724 , n4275 , n4723 );
and ( n4725 , n4216 , n4723 );
or ( n4726 , n4276 , n4724 , n4725 );
xor ( n4727 , n4214 , n4726 );
not ( n4728 , n4727 );
xor ( n4729 , n4216 , n4275 );
xor ( n4730 , n4729 , n4723 );
xor ( n4731 , n4278 , n4336 );
xor ( n4732 , n4731 , n4720 );
xor ( n4733 , n4339 , n4368 );
xor ( n4734 , n4733 , n4717 );
xor ( n4735 , n4371 , n4478 );
xor ( n4736 , n4735 , n4714 );
xor ( n4737 , n4481 , n4499 );
xor ( n4738 , n4737 , n4711 );
xor ( n4739 , n4502 , n4583 );
xor ( n4740 , n4739 , n4708 );
xor ( n4741 , n4636 , n4638 );
xor ( n4742 , n4741 , n4705 );
and ( n4743 , n4316 , n4302 );
and ( n4744 , n4256 , n4300 );
nor ( n4745 , n4743 , n4744 );
xnor ( n4746 , n4745 , n4285 );
and ( n4747 , n4513 , n4148 );
and ( n4748 , n4437 , n4146 );
nor ( n4749 , n4747 , n4748 );
xnor ( n4750 , n4749 , n4153 );
and ( n4751 , n4746 , n4750 );
and ( n4752 , n4678 , n4170 );
and ( n4753 , n4523 , n4168 );
nor ( n4754 , n4752 , n4753 );
xnor ( n4755 , n4754 , n4176 );
and ( n4756 , n4750 , n4755 );
and ( n4757 , n4746 , n4755 );
or ( n4758 , n4751 , n4756 , n4757 );
and ( n4759 , n4192 , n4605 );
and ( n4760 , n4162 , n4603 );
nor ( n4761 , n4759 , n4760 );
xnor ( n4762 , n4761 , n4552 );
and ( n4763 , n4234 , n4445 );
and ( n4764 , n4202 , n4443 );
nor ( n4765 , n4763 , n4764 );
xnor ( n4766 , n4765 , n4408 );
and ( n4767 , n4762 , n4766 );
and ( n4768 , n4419 , n4242 );
and ( n4769 , n4385 , n4240 );
nor ( n4770 , n4768 , n4769 );
xnor ( n4771 , n4770 , n4223 );
and ( n4772 , n4766 , n4771 );
and ( n4773 , n4762 , n4771 );
or ( n4774 , n4767 , n4772 , n4773 );
and ( n4775 , n4758 , n4774 );
xor ( n4776 , n4609 , n4613 );
xor ( n4777 , n4776 , n4618 );
and ( n4778 , n4774 , n4777 );
and ( n4779 , n4758 , n4777 );
or ( n4780 , n4775 , n4778 , n4779 );
not ( n4781 , n4668 );
xor ( n4782 , n4082 , n4083 );
xor ( n4783 , n4782 , n4093 );
buf ( n4784 , n4783 );
buf ( n4785 , n4784 );
buf ( n4786 , n4785 );
and ( n4787 , n4786 , n4164 );
or ( n4788 , n4781 , n4787 );
xor ( n4789 , n4549 , n4666 );
xor ( n4790 , n4666 , n4668 );
not ( n4791 , n4790 );
and ( n4792 , n4789 , n4791 );
and ( n4793 , n4138 , n4792 );
not ( n4794 , n4793 );
xnor ( n4795 , n4794 , n4671 );
and ( n4796 , n4788 , n4795 );
not ( n4797 , n4663 );
and ( n4798 , n4795 , n4797 );
and ( n4799 , n4788 , n4797 );
or ( n4800 , n4796 , n4798 , n4799 );
xor ( n4801 , n4645 , n4649 );
xor ( n4802 , n4801 , n4654 );
and ( n4803 , n4800 , n4802 );
xor ( n4804 , n4664 , n4672 );
xor ( n4805 , n4804 , n4679 );
and ( n4806 , n4802 , n4805 );
and ( n4807 , n4800 , n4805 );
or ( n4808 , n4803 , n4806 , n4807 );
and ( n4809 , n4780 , n4808 );
xor ( n4810 , n4657 , n4682 );
xor ( n4811 , n4810 , n4687 );
and ( n4812 , n4808 , n4811 );
and ( n4813 , n4780 , n4811 );
or ( n4814 , n4809 , n4812 , n4813 );
xor ( n4815 , n4589 , n4593 );
xor ( n4816 , n4815 , n4598 );
xor ( n4817 , n4621 , n4623 );
and ( n4818 , n4816 , n4817 );
xor ( n4819 , n4780 , n4808 );
xor ( n4820 , n4819 , n4811 );
and ( n4821 , n4817 , n4820 );
and ( n4822 , n4816 , n4820 );
or ( n4823 , n4818 , n4821 , n4822 );
and ( n4824 , n4814 , n4823 );
xor ( n4825 , n4696 , n4697 );
xor ( n4826 , n4825 , n4699 );
and ( n4827 , n4823 , n4826 );
and ( n4828 , n4814 , n4826 );
or ( n4829 , n4824 , n4827 , n4828 );
xor ( n4830 , n4641 , n4693 );
xor ( n4831 , n4830 , n4702 );
and ( n4832 , n4829 , n4831 );
xor ( n4833 , n4829 , n4831 );
and ( n4834 , n4256 , n4445 );
and ( n4835 , n4234 , n4443 );
nor ( n4836 , n4834 , n4835 );
xnor ( n4837 , n4836 , n4408 );
and ( n4838 , n4437 , n4242 );
and ( n4839 , n4419 , n4240 );
nor ( n4840 , n4838 , n4839 );
xnor ( n4841 , n4840 , n4223 );
and ( n4842 , n4837 , n4841 );
and ( n4843 , n4523 , n4148 );
and ( n4844 , n4513 , n4146 );
nor ( n4845 , n4843 , n4844 );
xnor ( n4846 , n4845 , n4153 );
and ( n4847 , n4841 , n4846 );
and ( n4848 , n4837 , n4846 );
or ( n4849 , n4842 , n4847 , n4848 );
xor ( n4850 , n4746 , n4750 );
xor ( n4851 , n4850 , n4755 );
and ( n4852 , n4849 , n4851 );
xor ( n4853 , n4762 , n4766 );
xor ( n4854 , n4853 , n4771 );
and ( n4855 , n4851 , n4854 );
and ( n4856 , n4849 , n4854 );
or ( n4857 , n4852 , n4855 , n4856 );
and ( n4858 , n4162 , n4792 );
and ( n4859 , n4138 , n4790 );
nor ( n4860 , n4858 , n4859 );
xnor ( n4861 , n4860 , n4671 );
and ( n4862 , n4202 , n4605 );
and ( n4863 , n4192 , n4603 );
nor ( n4864 , n4862 , n4863 );
xnor ( n4865 , n4864 , n4552 );
and ( n4866 , n4861 , n4865 );
and ( n4867 , n4385 , n4302 );
and ( n4868 , n4316 , n4300 );
nor ( n4869 , n4867 , n4868 );
xnor ( n4870 , n4869 , n4285 );
and ( n4871 , n4865 , n4870 );
and ( n4872 , n4861 , n4870 );
or ( n4873 , n4866 , n4871 , n4872 );
and ( n4874 , n4662 , n4170 );
and ( n4875 , n4678 , n4168 );
nor ( n4876 , n4874 , n4875 );
xnor ( n4877 , n4876 , n4176 );
xnor ( n4878 , n4781 , n4787 );
and ( n4879 , n4877 , n4878 );
and ( n4880 , n4873 , n4879 );
xor ( n4881 , n4788 , n4795 );
xor ( n4882 , n4881 , n4797 );
and ( n4883 , n4879 , n4882 );
and ( n4884 , n4873 , n4882 );
or ( n4885 , n4880 , n4883 , n4884 );
and ( n4886 , n4857 , n4885 );
xor ( n4887 , n4800 , n4802 );
xor ( n4888 , n4887 , n4805 );
and ( n4889 , n4885 , n4888 );
and ( n4890 , n4857 , n4888 );
or ( n4891 , n4886 , n4889 , n4890 );
and ( n4892 , n4316 , n4445 );
and ( n4893 , n4256 , n4443 );
nor ( n4894 , n4892 , n4893 );
xnor ( n4895 , n4894 , n4408 );
and ( n4896 , n4513 , n4242 );
and ( n4897 , n4437 , n4240 );
nor ( n4898 , n4896 , n4897 );
xnor ( n4899 , n4898 , n4223 );
and ( n4900 , n4895 , n4899 );
and ( n4901 , n4678 , n4148 );
and ( n4902 , n4523 , n4146 );
nor ( n4903 , n4901 , n4902 );
xnor ( n4904 , n4903 , n4153 );
and ( n4905 , n4899 , n4904 );
and ( n4906 , n4895 , n4904 );
or ( n4907 , n4900 , n4905 , n4906 );
and ( n4908 , n4662 , n4148 );
and ( n4909 , n4678 , n4146 );
nor ( n4910 , n4908 , n4909 );
xnor ( n4911 , n4910 , n4153 );
xor ( n4912 , n4085 , n4086 );
xor ( n4913 , n4912 , n4090 );
buf ( n4914 , n4913 );
buf ( n4915 , n4914 );
buf ( n4916 , n4915 );
and ( n4917 , n4916 , n4170 );
and ( n4918 , n4786 , n4168 );
nor ( n4919 , n4917 , n4918 );
xnor ( n4920 , n4919 , n4176 );
and ( n4921 , n4911 , n4920 );
xor ( n4922 , n4088 , n4089 );
buf ( n4923 , n4922 );
buf ( n4924 , n4923 );
buf ( n4925 , n4924 );
and ( n4926 , n4925 , n4164 );
and ( n4927 , n4920 , n4926 );
and ( n4928 , n4911 , n4926 );
or ( n4929 , n4921 , n4927 , n4928 );
and ( n4930 , n4192 , n4792 );
and ( n4931 , n4162 , n4790 );
nor ( n4932 , n4930 , n4931 );
xnor ( n4933 , n4932 , n4671 );
and ( n4934 , n4929 , n4933 );
and ( n4935 , n4419 , n4302 );
and ( n4936 , n4385 , n4300 );
nor ( n4937 , n4935 , n4936 );
xnor ( n4938 , n4937 , n4285 );
and ( n4939 , n4933 , n4938 );
and ( n4940 , n4929 , n4938 );
or ( n4941 , n4934 , n4939 , n4940 );
and ( n4942 , n4907 , n4941 );
xor ( n4943 , n4861 , n4865 );
xor ( n4944 , n4943 , n4870 );
and ( n4945 , n4941 , n4944 );
and ( n4946 , n4907 , n4944 );
or ( n4947 , n4942 , n4945 , n4946 );
xor ( n4948 , n4877 , n4878 );
buf ( n4949 , n559 );
buf ( n4950 , n4949 );
xor ( n4951 , n4668 , n4950 );
not ( n4952 , n4950 );
and ( n4953 , n4951 , n4952 );
and ( n4954 , n4138 , n4953 );
not ( n4955 , n4954 );
xnor ( n4956 , n4955 , n4668 );
and ( n4957 , n4786 , n4170 );
and ( n4958 , n4662 , n4168 );
nor ( n4959 , n4957 , n4958 );
xnor ( n4960 , n4959 , n4176 );
and ( n4961 , n4956 , n4960 );
and ( n4962 , n4916 , n4164 );
and ( n4963 , n4960 , n4962 );
and ( n4964 , n4956 , n4962 );
or ( n4965 , n4961 , n4963 , n4964 );
and ( n4966 , n4948 , n4965 );
xor ( n4967 , n4837 , n4841 );
xor ( n4968 , n4967 , n4846 );
and ( n4969 , n4965 , n4968 );
and ( n4970 , n4948 , n4968 );
or ( n4971 , n4966 , n4969 , n4970 );
and ( n4972 , n4947 , n4971 );
xor ( n4973 , n4873 , n4879 );
xor ( n4974 , n4973 , n4882 );
and ( n4975 , n4971 , n4974 );
and ( n4976 , n4947 , n4974 );
or ( n4977 , n4972 , n4975 , n4976 );
xor ( n4978 , n4758 , n4774 );
xor ( n4979 , n4978 , n4777 );
and ( n4980 , n4977 , n4979 );
xor ( n4981 , n4857 , n4885 );
xor ( n4982 , n4981 , n4888 );
and ( n4983 , n4979 , n4982 );
and ( n4984 , n4977 , n4982 );
or ( n4985 , n4980 , n4983 , n4984 );
and ( n4986 , n4891 , n4985 );
xor ( n4987 , n4816 , n4817 );
xor ( n4988 , n4987 , n4820 );
and ( n4989 , n4985 , n4988 );
and ( n4990 , n4891 , n4988 );
or ( n4991 , n4986 , n4989 , n4990 );
xor ( n4992 , n4814 , n4823 );
xor ( n4993 , n4992 , n4826 );
and ( n4994 , n4991 , n4993 );
xor ( n4995 , n4991 , n4993 );
xor ( n4996 , n4891 , n4985 );
xor ( n4997 , n4996 , n4988 );
and ( n4998 , n4162 , n4953 );
and ( n4999 , n4138 , n4950 );
nor ( n5000 , n4998 , n4999 );
xnor ( n5001 , n5000 , n4668 );
and ( n5002 , n4202 , n4792 );
and ( n5003 , n4192 , n4790 );
nor ( n5004 , n5002 , n5003 );
xnor ( n5005 , n5004 , n4671 );
and ( n5006 , n5001 , n5005 );
and ( n5007 , n4385 , n4445 );
and ( n5008 , n4316 , n4443 );
nor ( n5009 , n5007 , n5008 );
xnor ( n5010 , n5009 , n4408 );
and ( n5011 , n5005 , n5010 );
and ( n5012 , n5001 , n5010 );
or ( n5013 , n5006 , n5011 , n5012 );
xor ( n5014 , n4895 , n4899 );
xor ( n5015 , n5014 , n4904 );
and ( n5016 , n5013 , n5015 );
xor ( n5017 , n4929 , n4933 );
xor ( n5018 , n5017 , n4938 );
and ( n5019 , n5015 , n5018 );
and ( n5020 , n5013 , n5018 );
or ( n5021 , n5016 , n5019 , n5020 );
and ( n5022 , n4925 , n4168 );
not ( n5023 , n5022 );
and ( n5024 , n5023 , n4176 );
and ( n5025 , n4925 , n4170 );
and ( n5026 , n4916 , n4168 );
nor ( n5027 , n5025 , n5026 );
xnor ( n5028 , n5027 , n4176 );
and ( n5029 , n5024 , n5028 );
and ( n5030 , n4437 , n4302 );
and ( n5031 , n4419 , n4300 );
nor ( n5032 , n5030 , n5031 );
xnor ( n5033 , n5032 , n4285 );
and ( n5034 , n5029 , n5033 );
and ( n5035 , n4523 , n4242 );
and ( n5036 , n4513 , n4240 );
nor ( n5037 , n5035 , n5036 );
xnor ( n5038 , n5037 , n4223 );
and ( n5039 , n5033 , n5038 );
and ( n5040 , n5029 , n5038 );
or ( n5041 , n5034 , n5039 , n5040 );
and ( n5042 , n4234 , n4605 );
and ( n5043 , n4202 , n4603 );
nor ( n5044 , n5042 , n5043 );
xnor ( n5045 , n5044 , n4552 );
and ( n5046 , n5041 , n5045 );
xor ( n5047 , n4956 , n4960 );
xor ( n5048 , n5047 , n4962 );
and ( n5049 , n5045 , n5048 );
and ( n5050 , n5041 , n5048 );
or ( n5051 , n5046 , n5049 , n5050 );
and ( n5052 , n5021 , n5051 );
xor ( n5053 , n4948 , n4965 );
xor ( n5054 , n5053 , n4968 );
and ( n5055 , n5051 , n5054 );
and ( n5056 , n5021 , n5054 );
or ( n5057 , n5052 , n5055 , n5056 );
xor ( n5058 , n4849 , n4851 );
xor ( n5059 , n5058 , n4854 );
and ( n5060 , n5057 , n5059 );
xor ( n5061 , n4947 , n4971 );
xor ( n5062 , n5061 , n4974 );
and ( n5063 , n5059 , n5062 );
and ( n5064 , n5057 , n5062 );
or ( n5065 , n5060 , n5063 , n5064 );
xor ( n5066 , n4977 , n4979 );
xor ( n5067 , n5066 , n4982 );
and ( n5068 , n5065 , n5067 );
xor ( n5069 , n5057 , n5059 );
xor ( n5070 , n5069 , n5062 );
xor ( n5071 , n5024 , n5028 );
and ( n5072 , n4678 , n4242 );
and ( n5073 , n4523 , n4240 );
nor ( n5074 , n5072 , n5073 );
xnor ( n5075 , n5074 , n4223 );
and ( n5076 , n5071 , n5075 );
and ( n5077 , n4786 , n4148 );
and ( n5078 , n4662 , n4146 );
nor ( n5079 , n5077 , n5078 );
xnor ( n5080 , n5079 , n4153 );
and ( n5081 , n5075 , n5080 );
and ( n5082 , n5071 , n5080 );
or ( n5083 , n5076 , n5081 , n5082 );
and ( n5084 , n4256 , n4605 );
and ( n5085 , n4234 , n4603 );
nor ( n5086 , n5084 , n5085 );
xnor ( n5087 , n5086 , n4552 );
and ( n5088 , n5083 , n5087 );
xor ( n5089 , n4911 , n4920 );
xor ( n5090 , n5089 , n4926 );
and ( n5091 , n5087 , n5090 );
and ( n5092 , n5083 , n5090 );
or ( n5093 , n5088 , n5091 , n5092 );
and ( n5094 , n4192 , n4953 );
and ( n5095 , n4162 , n4950 );
nor ( n5096 , n5094 , n5095 );
xnor ( n5097 , n5096 , n4668 );
and ( n5098 , n4419 , n4445 );
and ( n5099 , n4385 , n4443 );
nor ( n5100 , n5098 , n5099 );
xnor ( n5101 , n5100 , n4408 );
and ( n5102 , n5097 , n5101 );
and ( n5103 , n4513 , n4302 );
and ( n5104 , n4437 , n4300 );
nor ( n5105 , n5103 , n5104 );
xnor ( n5106 , n5105 , n4285 );
and ( n5107 , n5101 , n5106 );
and ( n5108 , n5097 , n5106 );
or ( n5109 , n5102 , n5107 , n5108 );
and ( n5110 , n4925 , n4146 );
not ( n5111 , n5110 );
and ( n5112 , n5111 , n4153 );
and ( n5113 , n4925 , n4148 );
and ( n5114 , n4916 , n4146 );
nor ( n5115 , n5113 , n5114 );
xnor ( n5116 , n5115 , n4153 );
and ( n5117 , n5112 , n5116 );
and ( n5118 , n4916 , n4148 );
and ( n5119 , n4786 , n4146 );
nor ( n5120 , n5118 , n5119 );
xnor ( n5121 , n5120 , n4153 );
and ( n5122 , n5117 , n5121 );
and ( n5123 , n5121 , n5022 );
and ( n5124 , n5117 , n5022 );
or ( n5125 , n5122 , n5123 , n5124 );
and ( n5126 , n4234 , n4792 );
and ( n5127 , n4202 , n4790 );
nor ( n5128 , n5126 , n5127 );
xnor ( n5129 , n5128 , n4671 );
and ( n5130 , n5125 , n5129 );
and ( n5131 , n4316 , n4605 );
and ( n5132 , n4256 , n4603 );
nor ( n5133 , n5131 , n5132 );
xnor ( n5134 , n5133 , n4552 );
and ( n5135 , n5129 , n5134 );
and ( n5136 , n5125 , n5134 );
or ( n5137 , n5130 , n5135 , n5136 );
and ( n5138 , n5109 , n5137 );
xor ( n5139 , n5029 , n5033 );
xor ( n5140 , n5139 , n5038 );
and ( n5141 , n5137 , n5140 );
and ( n5142 , n5109 , n5140 );
or ( n5143 , n5138 , n5141 , n5142 );
and ( n5144 , n5093 , n5143 );
xor ( n5145 , n5041 , n5045 );
xor ( n5146 , n5145 , n5048 );
and ( n5147 , n5143 , n5146 );
and ( n5148 , n5093 , n5146 );
or ( n5149 , n5144 , n5147 , n5148 );
xor ( n5150 , n4907 , n4941 );
xor ( n5151 , n5150 , n4944 );
and ( n5152 , n5149 , n5151 );
xor ( n5153 , n5021 , n5051 );
xor ( n5154 , n5153 , n5054 );
and ( n5155 , n5151 , n5154 );
and ( n5156 , n5149 , n5154 );
or ( n5157 , n5152 , n5155 , n5156 );
and ( n5158 , n5070 , n5157 );
xor ( n5159 , n5149 , n5151 );
xor ( n5160 , n5159 , n5154 );
and ( n5161 , n4437 , n4445 );
and ( n5162 , n4419 , n4443 );
nor ( n5163 , n5161 , n5162 );
xnor ( n5164 , n5163 , n4408 );
and ( n5165 , n4523 , n4302 );
and ( n5166 , n4513 , n4300 );
nor ( n5167 , n5165 , n5166 );
xnor ( n5168 , n5167 , n4285 );
and ( n5169 , n5164 , n5168 );
and ( n5170 , n4662 , n4242 );
and ( n5171 , n4678 , n4240 );
nor ( n5172 , n5170 , n5171 );
xnor ( n5173 , n5172 , n4223 );
and ( n5174 , n5168 , n5173 );
and ( n5175 , n5164 , n5173 );
or ( n5176 , n5169 , n5174 , n5175 );
and ( n5177 , n4202 , n4953 );
and ( n5178 , n4192 , n4950 );
nor ( n5179 , n5177 , n5178 );
xnor ( n5180 , n5179 , n4668 );
and ( n5181 , n4256 , n4792 );
and ( n5182 , n4234 , n4790 );
nor ( n5183 , n5181 , n5182 );
xnor ( n5184 , n5183 , n4671 );
and ( n5185 , n5180 , n5184 );
xor ( n5186 , n5117 , n5121 );
xor ( n5187 , n5186 , n5022 );
and ( n5188 , n5184 , n5187 );
and ( n5189 , n5180 , n5187 );
or ( n5190 , n5185 , n5188 , n5189 );
and ( n5191 , n5176 , n5190 );
xor ( n5192 , n5071 , n5075 );
xor ( n5193 , n5192 , n5080 );
and ( n5194 , n5190 , n5193 );
and ( n5195 , n5176 , n5193 );
or ( n5196 , n5191 , n5194 , n5195 );
xor ( n5197 , n5001 , n5005 );
xor ( n5198 , n5197 , n5010 );
and ( n5199 , n5196 , n5198 );
xor ( n5200 , n5083 , n5087 );
xor ( n5201 , n5200 , n5090 );
and ( n5202 , n5198 , n5201 );
and ( n5203 , n5196 , n5201 );
or ( n5204 , n5199 , n5202 , n5203 );
xor ( n5205 , n5013 , n5015 );
xor ( n5206 , n5205 , n5018 );
and ( n5207 , n5204 , n5206 );
xor ( n5208 , n5093 , n5143 );
xor ( n5209 , n5208 , n5146 );
and ( n5210 , n5206 , n5209 );
and ( n5211 , n5204 , n5209 );
or ( n5212 , n5207 , n5210 , n5211 );
and ( n5213 , n5160 , n5212 );
xor ( n5214 , n5204 , n5206 );
xor ( n5215 , n5214 , n5209 );
xor ( n5216 , n5097 , n5101 );
xor ( n5217 , n5216 , n5106 );
xor ( n5218 , n5125 , n5129 );
xor ( n5219 , n5218 , n5134 );
and ( n5220 , n5217 , n5219 );
xor ( n5221 , n5176 , n5190 );
xor ( n5222 , n5221 , n5193 );
and ( n5223 , n5219 , n5222 );
and ( n5224 , n5217 , n5222 );
or ( n5225 , n5220 , n5223 , n5224 );
xor ( n5226 , n5109 , n5137 );
xor ( n5227 , n5226 , n5140 );
and ( n5228 , n5225 , n5227 );
xor ( n5229 , n5196 , n5198 );
xor ( n5230 , n5229 , n5201 );
and ( n5231 , n5227 , n5230 );
and ( n5232 , n5225 , n5230 );
or ( n5233 , n5228 , n5231 , n5232 );
and ( n5234 , n5215 , n5233 );
xor ( n5235 , n5225 , n5227 );
xor ( n5236 , n5235 , n5230 );
xor ( n5237 , n5112 , n5116 );
and ( n5238 , n4678 , n4302 );
and ( n5239 , n4523 , n4300 );
nor ( n5240 , n5238 , n5239 );
xnor ( n5241 , n5240 , n4285 );
and ( n5242 , n5237 , n5241 );
and ( n5243 , n4786 , n4242 );
and ( n5244 , n4662 , n4240 );
nor ( n5245 , n5243 , n5244 );
xnor ( n5246 , n5245 , n4223 );
and ( n5247 , n5241 , n5246 );
and ( n5248 , n5237 , n5246 );
or ( n5249 , n5242 , n5247 , n5248 );
and ( n5250 , n4385 , n4605 );
and ( n5251 , n4316 , n4603 );
nor ( n5252 , n5250 , n5251 );
xnor ( n5253 , n5252 , n4552 );
and ( n5254 , n5249 , n5253 );
xor ( n5255 , n5164 , n5168 );
xor ( n5256 , n5255 , n5173 );
and ( n5257 , n5253 , n5256 );
and ( n5258 , n5249 , n5256 );
or ( n5259 , n5254 , n5257 , n5258 );
and ( n5260 , n4925 , n4240 );
not ( n5261 , n5260 );
and ( n5262 , n5261 , n4223 );
and ( n5263 , n4925 , n4242 );
and ( n5264 , n4916 , n4240 );
nor ( n5265 , n5263 , n5264 );
xnor ( n5266 , n5265 , n4223 );
and ( n5267 , n5262 , n5266 );
and ( n5268 , n4916 , n4242 );
and ( n5269 , n4786 , n4240 );
nor ( n5270 , n5268 , n5269 );
xnor ( n5271 , n5270 , n4223 );
and ( n5272 , n5267 , n5271 );
and ( n5273 , n5271 , n5110 );
and ( n5274 , n5267 , n5110 );
or ( n5275 , n5272 , n5273 , n5274 );
and ( n5276 , n4316 , n4792 );
and ( n5277 , n4256 , n4790 );
nor ( n5278 , n5276 , n5277 );
xnor ( n5279 , n5278 , n4671 );
and ( n5280 , n5275 , n5279 );
and ( n5281 , n4513 , n4445 );
and ( n5282 , n4437 , n4443 );
nor ( n5283 , n5281 , n5282 );
xnor ( n5284 , n5283 , n4408 );
and ( n5285 , n5279 , n5284 );
and ( n5286 , n5275 , n5284 );
or ( n5287 , n5280 , n5285 , n5286 );
xor ( n5288 , n5180 , n5184 );
xor ( n5289 , n5288 , n5187 );
and ( n5290 , n5287 , n5289 );
and ( n5291 , n5259 , n5290 );
xor ( n5292 , n5217 , n5219 );
xor ( n5293 , n5292 , n5222 );
and ( n5294 , n5290 , n5293 );
and ( n5295 , n5259 , n5293 );
or ( n5296 , n5291 , n5294 , n5295 );
and ( n5297 , n5236 , n5296 );
and ( n5298 , n4234 , n4953 );
and ( n5299 , n4202 , n4950 );
nor ( n5300 , n5298 , n5299 );
xnor ( n5301 , n5300 , n4668 );
and ( n5302 , n4419 , n4605 );
and ( n5303 , n4385 , n4603 );
nor ( n5304 , n5302 , n5303 );
xnor ( n5305 , n5304 , n4552 );
and ( n5306 , n5301 , n5305 );
and ( n5307 , n4437 , n4605 );
and ( n5308 , n4419 , n4603 );
nor ( n5309 , n5307 , n5308 );
xnor ( n5310 , n5309 , n4552 );
and ( n5311 , n4523 , n4445 );
and ( n5312 , n4513 , n4443 );
nor ( n5313 , n5311 , n5312 );
xnor ( n5314 , n5313 , n4408 );
and ( n5315 , n5310 , n5314 );
and ( n5316 , n4662 , n4302 );
and ( n5317 , n4678 , n4300 );
nor ( n5318 , n5316 , n5317 );
xnor ( n5319 , n5318 , n4285 );
and ( n5320 , n5314 , n5319 );
and ( n5321 , n5310 , n5319 );
or ( n5322 , n5315 , n5320 , n5321 );
and ( n5323 , n5305 , n5322 );
and ( n5324 , n5301 , n5322 );
or ( n5325 , n5306 , n5323 , n5324 );
xor ( n5326 , n5249 , n5253 );
xor ( n5327 , n5326 , n5256 );
and ( n5328 , n5325 , n5327 );
xor ( n5329 , n5287 , n5289 );
and ( n5330 , n5327 , n5329 );
and ( n5331 , n5325 , n5329 );
or ( n5332 , n5328 , n5330 , n5331 );
xor ( n5333 , n5237 , n5241 );
xor ( n5334 , n5333 , n5246 );
xor ( n5335 , n5301 , n5305 );
xor ( n5336 , n5335 , n5322 );
and ( n5337 , n5334 , n5336 );
xor ( n5338 , n5275 , n5279 );
xor ( n5339 , n5338 , n5284 );
and ( n5340 , n5336 , n5339 );
and ( n5341 , n5334 , n5339 );
or ( n5342 , n5337 , n5340 , n5341 );
and ( n5343 , n4662 , n4445 );
and ( n5344 , n4678 , n4443 );
nor ( n5345 , n5343 , n5344 );
xnor ( n5346 , n5345 , n4408 );
and ( n5347 , n4916 , n4302 );
and ( n5348 , n4786 , n4300 );
nor ( n5349 , n5347 , n5348 );
xnor ( n5350 , n5349 , n4285 );
and ( n5351 , n5346 , n5350 );
and ( n5352 , n5350 , n5260 );
and ( n5353 , n5346 , n5260 );
or ( n5354 , n5351 , n5352 , n5353 );
and ( n5355 , n4419 , n4792 );
and ( n5356 , n4385 , n4790 );
nor ( n5357 , n5355 , n5356 );
xnor ( n5358 , n5357 , n4671 );
and ( n5359 , n5354 , n5358 );
and ( n5360 , n4513 , n4605 );
and ( n5361 , n4437 , n4603 );
nor ( n5362 , n5360 , n5361 );
xnor ( n5363 , n5362 , n4552 );
and ( n5364 , n5358 , n5363 );
and ( n5365 , n5354 , n5363 );
or ( n5366 , n5359 , n5364 , n5365 );
xor ( n5367 , n5262 , n5266 );
and ( n5368 , n4678 , n4445 );
and ( n5369 , n4523 , n4443 );
nor ( n5370 , n5368 , n5369 );
xnor ( n5371 , n5370 , n4408 );
and ( n5372 , n5367 , n5371 );
and ( n5373 , n4786 , n4302 );
and ( n5374 , n4662 , n4300 );
nor ( n5375 , n5373 , n5374 );
xnor ( n5376 , n5375 , n4285 );
and ( n5377 , n5371 , n5376 );
and ( n5378 , n5367 , n5376 );
or ( n5379 , n5372 , n5377 , n5378 );
and ( n5380 , n5366 , n5379 );
xor ( n5381 , n5310 , n5314 );
xor ( n5382 , n5381 , n5319 );
and ( n5383 , n5379 , n5382 );
and ( n5384 , n5366 , n5382 );
or ( n5385 , n5380 , n5383 , n5384 );
and ( n5386 , n4385 , n4792 );
and ( n5387 , n4316 , n4790 );
nor ( n5388 , n5386 , n5387 );
xnor ( n5389 , n5388 , n4671 );
xor ( n5390 , n5267 , n5271 );
xor ( n5391 , n5390 , n5110 );
and ( n5392 , n5389 , n5391 );
and ( n5393 , n5385 , n5392 );
and ( n5394 , n4256 , n4953 );
and ( n5395 , n4234 , n4950 );
nor ( n5396 , n5394 , n5395 );
xnor ( n5397 , n5396 , n4668 );
xor ( n5398 , n5366 , n5379 );
xor ( n5399 , n5398 , n5382 );
and ( n5400 , n5397 , n5399 );
xor ( n5401 , n5389 , n5391 );
and ( n5402 , n5399 , n5401 );
and ( n5403 , n5397 , n5401 );
or ( n5404 , n5400 , n5402 , n5403 );
and ( n5405 , n5392 , n5404 );
and ( n5406 , n5385 , n5404 );
or ( n5407 , n5393 , n5405 , n5406 );
and ( n5408 , n5342 , n5407 );
xor ( n5409 , n5325 , n5327 );
xor ( n5410 , n5409 , n5329 );
and ( n5411 , n5407 , n5410 );
and ( n5412 , n5342 , n5410 );
or ( n5413 , n5408 , n5411 , n5412 );
and ( n5414 , n5332 , n5413 );
xor ( n5415 , n5259 , n5290 );
xor ( n5416 , n5415 , n5293 );
and ( n5417 , n5413 , n5416 );
and ( n5418 , n5332 , n5416 );
or ( n5419 , n5414 , n5417 , n5418 );
and ( n5420 , n5296 , n5419 );
and ( n5421 , n5236 , n5419 );
or ( n5422 , n5297 , n5420 , n5421 );
and ( n5423 , n5233 , n5422 );
and ( n5424 , n5215 , n5422 );
or ( n5425 , n5234 , n5423 , n5424 );
and ( n5426 , n5212 , n5425 );
and ( n5427 , n5160 , n5425 );
or ( n5428 , n5213 , n5426 , n5427 );
and ( n5429 , n5157 , n5428 );
and ( n5430 , n5070 , n5428 );
or ( n5431 , n5158 , n5429 , n5430 );
and ( n5432 , n5067 , n5431 );
and ( n5433 , n5065 , n5431 );
or ( n5434 , n5068 , n5432 , n5433 );
and ( n5435 , n4997 , n5434 );
xor ( n5436 , n4997 , n5434 );
xor ( n5437 , n5065 , n5067 );
xor ( n5438 , n5437 , n5431 );
xor ( n5439 , n5070 , n5157 );
xor ( n5440 , n5439 , n5428 );
xor ( n5441 , n5160 , n5212 );
xor ( n5442 , n5441 , n5425 );
xor ( n5443 , n5215 , n5233 );
xor ( n5444 , n5443 , n5422 );
xor ( n5445 , n5236 , n5296 );
xor ( n5446 , n5445 , n5419 );
xor ( n5447 , n5332 , n5413 );
xor ( n5448 , n5447 , n5416 );
xor ( n5449 , n5334 , n5336 );
xor ( n5450 , n5449 , n5339 );
and ( n5451 , n4925 , n4300 );
not ( n5452 , n5451 );
and ( n5453 , n5452 , n4285 );
and ( n5454 , n4925 , n4302 );
and ( n5455 , n4916 , n4300 );
nor ( n5456 , n5454 , n5455 );
xnor ( n5457 , n5456 , n4285 );
and ( n5458 , n5453 , n5457 );
and ( n5459 , n4437 , n4792 );
and ( n5460 , n4419 , n4790 );
nor ( n5461 , n5459 , n5460 );
xnor ( n5462 , n5461 , n4671 );
and ( n5463 , n5458 , n5462 );
and ( n5464 , n4523 , n4605 );
and ( n5465 , n4513 , n4603 );
nor ( n5466 , n5464 , n5465 );
xnor ( n5467 , n5466 , n4552 );
and ( n5468 , n5462 , n5467 );
and ( n5469 , n5458 , n5467 );
or ( n5470 , n5463 , n5468 , n5469 );
and ( n5471 , n4316 , n4953 );
and ( n5472 , n4256 , n4950 );
nor ( n5473 , n5471 , n5472 );
xnor ( n5474 , n5473 , n4668 );
and ( n5475 , n5470 , n5474 );
xor ( n5476 , n5367 , n5371 );
xor ( n5477 , n5476 , n5376 );
and ( n5478 , n5474 , n5477 );
and ( n5479 , n5470 , n5477 );
or ( n5480 , n5475 , n5478 , n5479 );
xor ( n5481 , n5453 , n5457 );
and ( n5482 , n4513 , n4792 );
and ( n5483 , n4437 , n4790 );
nor ( n5484 , n5482 , n5483 );
xnor ( n5485 , n5484 , n4671 );
and ( n5486 , n5481 , n5485 );
and ( n5487 , n4786 , n4445 );
and ( n5488 , n4662 , n4443 );
nor ( n5489 , n5487 , n5488 );
xnor ( n5490 , n5489 , n4408 );
and ( n5491 , n5485 , n5490 );
and ( n5492 , n5481 , n5490 );
or ( n5493 , n5486 , n5491 , n5492 );
and ( n5494 , n4385 , n4953 );
and ( n5495 , n4316 , n4950 );
nor ( n5496 , n5494 , n5495 );
xnor ( n5497 , n5496 , n4668 );
and ( n5498 , n5493 , n5497 );
xor ( n5499 , n5346 , n5350 );
xor ( n5500 , n5499 , n5260 );
and ( n5501 , n5497 , n5500 );
and ( n5502 , n5493 , n5500 );
or ( n5503 , n5498 , n5501 , n5502 );
xor ( n5504 , n5354 , n5358 );
xor ( n5505 , n5504 , n5363 );
and ( n5506 , n5503 , n5505 );
xor ( n5507 , n5470 , n5474 );
xor ( n5508 , n5507 , n5477 );
and ( n5509 , n5505 , n5508 );
and ( n5510 , n5503 , n5508 );
or ( n5511 , n5506 , n5509 , n5510 );
and ( n5512 , n5480 , n5511 );
xor ( n5513 , n5397 , n5399 );
xor ( n5514 , n5513 , n5401 );
and ( n5515 , n5511 , n5514 );
and ( n5516 , n5480 , n5514 );
or ( n5517 , n5512 , n5515 , n5516 );
and ( n5518 , n5450 , n5517 );
xor ( n5519 , n5385 , n5392 );
xor ( n5520 , n5519 , n5404 );
and ( n5521 , n5517 , n5520 );
and ( n5522 , n5450 , n5520 );
or ( n5523 , n5518 , n5521 , n5522 );
xor ( n5524 , n5342 , n5407 );
xor ( n5525 , n5524 , n5410 );
and ( n5526 , n5523 , n5525 );
xor ( n5527 , n5523 , n5525 );
xor ( n5528 , n5450 , n5517 );
xor ( n5529 , n5528 , n5520 );
xor ( n5530 , n5480 , n5511 );
xor ( n5531 , n5530 , n5514 );
xor ( n5532 , n5503 , n5505 );
xor ( n5533 , n5532 , n5508 );
and ( n5534 , n4662 , n4605 );
and ( n5535 , n4678 , n4603 );
nor ( n5536 , n5534 , n5535 );
xnor ( n5537 , n5536 , n4552 );
and ( n5538 , n4916 , n4445 );
and ( n5539 , n4786 , n4443 );
nor ( n5540 , n5538 , n5539 );
xnor ( n5541 , n5540 , n4408 );
and ( n5542 , n5537 , n5541 );
and ( n5543 , n5541 , n5451 );
and ( n5544 , n5537 , n5451 );
or ( n5545 , n5542 , n5543 , n5544 );
and ( n5546 , n4419 , n4953 );
and ( n5547 , n4385 , n4950 );
nor ( n5548 , n5546 , n5547 );
xnor ( n5549 , n5548 , n4668 );
and ( n5550 , n5545 , n5549 );
and ( n5551 , n4678 , n4605 );
and ( n5552 , n4523 , n4603 );
nor ( n5553 , n5551 , n5552 );
xnor ( n5554 , n5553 , n4552 );
and ( n5555 , n5549 , n5554 );
and ( n5556 , n5545 , n5554 );
or ( n5557 , n5550 , n5555 , n5556 );
xor ( n5558 , n5458 , n5462 );
xor ( n5559 , n5558 , n5467 );
and ( n5560 , n5557 , n5559 );
xor ( n5561 , n5493 , n5497 );
xor ( n5562 , n5561 , n5500 );
and ( n5563 , n5559 , n5562 );
and ( n5564 , n5557 , n5562 );
or ( n5565 , n5560 , n5563 , n5564 );
and ( n5566 , n5533 , n5565 );
xor ( n5567 , n5533 , n5565 );
and ( n5568 , n4925 , n4443 );
not ( n5569 , n5568 );
and ( n5570 , n5569 , n4408 );
and ( n5571 , n4925 , n4445 );
and ( n5572 , n4916 , n4443 );
nor ( n5573 , n5571 , n5572 );
xnor ( n5574 , n5573 , n4408 );
and ( n5575 , n5570 , n5574 );
and ( n5576 , n4437 , n4953 );
and ( n5577 , n4419 , n4950 );
nor ( n5578 , n5576 , n5577 );
xnor ( n5579 , n5578 , n4668 );
and ( n5580 , n5575 , n5579 );
and ( n5581 , n4523 , n4792 );
and ( n5582 , n4513 , n4790 );
nor ( n5583 , n5581 , n5582 );
xnor ( n5584 , n5583 , n4671 );
and ( n5585 , n5579 , n5584 );
and ( n5586 , n5575 , n5584 );
or ( n5587 , n5580 , n5585 , n5586 );
xor ( n5588 , n5545 , n5549 );
xor ( n5589 , n5588 , n5554 );
and ( n5590 , n5587 , n5589 );
xor ( n5591 , n5481 , n5485 );
xor ( n5592 , n5591 , n5490 );
and ( n5593 , n5589 , n5592 );
and ( n5594 , n5587 , n5592 );
or ( n5595 , n5590 , n5593 , n5594 );
xor ( n5596 , n5557 , n5559 );
xor ( n5597 , n5596 , n5562 );
and ( n5598 , n5595 , n5597 );
xor ( n5599 , n5595 , n5597 );
xor ( n5600 , n5587 , n5589 );
xor ( n5601 , n5600 , n5592 );
xor ( n5602 , n5570 , n5574 );
and ( n5603 , n4678 , n4792 );
and ( n5604 , n4523 , n4790 );
nor ( n5605 , n5603 , n5604 );
xnor ( n5606 , n5605 , n4671 );
and ( n5607 , n5602 , n5606 );
and ( n5608 , n4786 , n4605 );
and ( n5609 , n4662 , n4603 );
nor ( n5610 , n5608 , n5609 );
xnor ( n5611 , n5610 , n4552 );
and ( n5612 , n5606 , n5611 );
and ( n5613 , n5602 , n5611 );
or ( n5614 , n5607 , n5612 , n5613 );
xor ( n5615 , n5537 , n5541 );
xor ( n5616 , n5615 , n5451 );
and ( n5617 , n5614 , n5616 );
xor ( n5618 , n5575 , n5579 );
xor ( n5619 , n5618 , n5584 );
and ( n5620 , n5616 , n5619 );
and ( n5621 , n5614 , n5619 );
or ( n5622 , n5617 , n5620 , n5621 );
and ( n5623 , n5601 , n5622 );
xor ( n5624 , n5601 , n5622 );
xor ( n5625 , n5614 , n5616 );
xor ( n5626 , n5625 , n5619 );
and ( n5627 , n4925 , n4603 );
not ( n5628 , n5627 );
and ( n5629 , n5628 , n4552 );
and ( n5630 , n4925 , n4605 );
and ( n5631 , n4916 , n4603 );
nor ( n5632 , n5630 , n5631 );
xnor ( n5633 , n5632 , n4552 );
and ( n5634 , n5629 , n5633 );
and ( n5635 , n4916 , n4605 );
and ( n5636 , n4786 , n4603 );
nor ( n5637 , n5635 , n5636 );
xnor ( n5638 , n5637 , n4552 );
and ( n5639 , n5634 , n5638 );
and ( n5640 , n5638 , n5568 );
and ( n5641 , n5634 , n5568 );
or ( n5642 , n5639 , n5640 , n5641 );
and ( n5643 , n4513 , n4953 );
and ( n5644 , n4437 , n4950 );
nor ( n5645 , n5643 , n5644 );
xnor ( n5646 , n5645 , n4668 );
and ( n5647 , n5642 , n5646 );
xor ( n5648 , n5602 , n5606 );
xor ( n5649 , n5648 , n5611 );
and ( n5650 , n5646 , n5649 );
and ( n5651 , n5642 , n5649 );
or ( n5652 , n5647 , n5650 , n5651 );
and ( n5653 , n5626 , n5652 );
xor ( n5654 , n5626 , n5652 );
xor ( n5655 , n5642 , n5646 );
xor ( n5656 , n5655 , n5649 );
and ( n5657 , n4523 , n4953 );
and ( n5658 , n4513 , n4950 );
nor ( n5659 , n5657 , n5658 );
xnor ( n5660 , n5659 , n4668 );
and ( n5661 , n4662 , n4792 );
and ( n5662 , n4678 , n4790 );
nor ( n5663 , n5661 , n5662 );
xnor ( n5664 , n5663 , n4671 );
and ( n5665 , n5660 , n5664 );
xor ( n5666 , n5634 , n5638 );
xor ( n5667 , n5666 , n5568 );
and ( n5668 , n5664 , n5667 );
and ( n5669 , n5660 , n5667 );
or ( n5670 , n5665 , n5668 , n5669 );
and ( n5671 , n5656 , n5670 );
xor ( n5672 , n5656 , n5670 );
xor ( n5673 , n5629 , n5633 );
and ( n5674 , n4678 , n4953 );
and ( n5675 , n4523 , n4950 );
nor ( n5676 , n5674 , n5675 );
xnor ( n5677 , n5676 , n4668 );
and ( n5678 , n5673 , n5677 );
and ( n5679 , n4786 , n4792 );
and ( n5680 , n4662 , n4790 );
nor ( n5681 , n5679 , n5680 );
xnor ( n5682 , n5681 , n4671 );
and ( n5683 , n5677 , n5682 );
and ( n5684 , n5673 , n5682 );
or ( n5685 , n5678 , n5683 , n5684 );
xor ( n5686 , n5660 , n5664 );
xor ( n5687 , n5686 , n5667 );
and ( n5688 , n5685 , n5687 );
xor ( n5689 , n5685 , n5687 );
xor ( n5690 , n5673 , n5677 );
xor ( n5691 , n5690 , n5682 );
and ( n5692 , n4925 , n4790 );
not ( n5693 , n5692 );
and ( n5694 , n5693 , n4671 );
and ( n5695 , n4925 , n4792 );
and ( n5696 , n4916 , n4790 );
nor ( n5697 , n5695 , n5696 );
xnor ( n5698 , n5697 , n4671 );
and ( n5699 , n5694 , n5698 );
and ( n5700 , n4916 , n4792 );
and ( n5701 , n4786 , n4790 );
nor ( n5702 , n5700 , n5701 );
xnor ( n5703 , n5702 , n4671 );
and ( n5704 , n5699 , n5703 );
and ( n5705 , n5703 , n5627 );
and ( n5706 , n5699 , n5627 );
or ( n5707 , n5704 , n5705 , n5706 );
and ( n5708 , n5691 , n5707 );
xor ( n5709 , n5691 , n5707 );
and ( n5710 , n4662 , n4953 );
and ( n5711 , n4678 , n4950 );
nor ( n5712 , n5710 , n5711 );
xnor ( n5713 , n5712 , n4668 );
xor ( n5714 , n5699 , n5703 );
xor ( n5715 , n5714 , n5627 );
and ( n5716 , n5713 , n5715 );
xor ( n5717 , n5713 , n5715 );
and ( n5718 , n4786 , n4953 );
and ( n5719 , n4662 , n4950 );
nor ( n5720 , n5718 , n5719 );
xnor ( n5721 , n5720 , n4668 );
xor ( n5722 , n5694 , n5698 );
and ( n5723 , n5721 , n5722 );
xor ( n5724 , n5721 , n5722 );
and ( n5725 , n4916 , n4953 );
and ( n5726 , n4786 , n4950 );
nor ( n5727 , n5725 , n5726 );
xnor ( n5728 , n5727 , n4668 );
and ( n5729 , n5728 , n5692 );
xor ( n5730 , n5728 , n5692 );
and ( n5731 , n4925 , n4953 );
and ( n5732 , n4916 , n4950 );
nor ( n5733 , n5731 , n5732 );
xnor ( n5734 , n5733 , n4668 );
and ( n5735 , n4925 , n4950 );
not ( n5736 , n5735 );
and ( n5737 , n5736 , n4668 );
and ( n5738 , n5734 , n5737 );
and ( n5739 , n5730 , n5738 );
or ( n5740 , n5729 , n5739 );
and ( n5741 , n5724 , n5740 );
or ( n5742 , n5723 , n5741 );
and ( n5743 , n5717 , n5742 );
or ( n5744 , n5716 , n5743 );
and ( n5745 , n5709 , n5744 );
or ( n5746 , n5708 , n5745 );
and ( n5747 , n5689 , n5746 );
or ( n5748 , n5688 , n5747 );
and ( n5749 , n5672 , n5748 );
or ( n5750 , n5671 , n5749 );
and ( n5751 , n5654 , n5750 );
or ( n5752 , n5653 , n5751 );
and ( n5753 , n5624 , n5752 );
or ( n5754 , n5623 , n5753 );
and ( n5755 , n5599 , n5754 );
or ( n5756 , n5598 , n5755 );
and ( n5757 , n5567 , n5756 );
or ( n5758 , n5566 , n5757 );
and ( n5759 , n5531 , n5758 );
and ( n5760 , n5529 , n5759 );
and ( n5761 , n5527 , n5760 );
or ( n5762 , n5526 , n5761 );
and ( n5763 , n5448 , n5762 );
and ( n5764 , n5446 , n5763 );
and ( n5765 , n5444 , n5764 );
and ( n5766 , n5442 , n5765 );
and ( n5767 , n5440 , n5766 );
and ( n5768 , n5438 , n5767 );
and ( n5769 , n5436 , n5768 );
or ( n5770 , n5435 , n5769 );
and ( n5771 , n4995 , n5770 );
or ( n5772 , n4994 , n5771 );
and ( n5773 , n4833 , n5772 );
or ( n5774 , n4832 , n5773 );
and ( n5775 , n4742 , n5774 );
and ( n5776 , n4740 , n5775 );
and ( n5777 , n4738 , n5776 );
and ( n5778 , n4736 , n5777 );
and ( n5779 , n4734 , n5778 );
and ( n5780 , n4732 , n5779 );
and ( n5781 , n4730 , n5780 );
xor ( n5782 , n4728 , n5781 );
buf ( n5783 , n5782 );
buf ( n5784 , n5783 );
not ( n5785 , n5784 );
and ( n5786 , n4042 , n5785 );
xor ( n5787 , n1175 , n4037 );
buf ( n5788 , n5787 );
buf ( n5789 , n5788 );
xor ( n5790 , n4730 , n5780 );
buf ( n5791 , n5790 );
buf ( n5792 , n5791 );
not ( n5793 , n5792 );
and ( n5794 , n5789 , n5793 );
xor ( n5795 , n1276 , n4035 );
buf ( n5796 , n5795 );
buf ( n5797 , n5796 );
xor ( n5798 , n4732 , n5779 );
buf ( n5799 , n5798 );
buf ( n5800 , n5799 );
not ( n5801 , n5800 );
and ( n5802 , n5797 , n5801 );
xor ( n5803 , n1400 , n4033 );
buf ( n5804 , n5803 );
buf ( n5805 , n5804 );
xor ( n5806 , n4734 , n5778 );
buf ( n5807 , n5806 );
buf ( n5808 , n5807 );
not ( n5809 , n5808 );
and ( n5810 , n5805 , n5809 );
xor ( n5811 , n1532 , n4031 );
buf ( n5812 , n5811 );
buf ( n5813 , n5812 );
xor ( n5814 , n4736 , n5777 );
buf ( n5815 , n5814 );
buf ( n5816 , n5815 );
not ( n5817 , n5816 );
and ( n5818 , n5813 , n5817 );
xor ( n5819 , n1820 , n4029 );
buf ( n5820 , n5819 );
buf ( n5821 , n5820 );
xor ( n5822 , n4738 , n5776 );
buf ( n5823 , n5822 );
buf ( n5824 , n5823 );
not ( n5825 , n5824 );
and ( n5826 , n5821 , n5825 );
xor ( n5827 , n2002 , n4027 );
buf ( n5828 , n5827 );
buf ( n5829 , n5828 );
xor ( n5830 , n4740 , n5775 );
buf ( n5831 , n5830 );
buf ( n5832 , n5831 );
not ( n5833 , n5832 );
and ( n5834 , n5829 , n5833 );
xor ( n5835 , n2126 , n4025 );
buf ( n5836 , n5835 );
buf ( n5837 , n5836 );
xor ( n5838 , n4742 , n5774 );
buf ( n5839 , n5838 );
buf ( n5840 , n5839 );
not ( n5841 , n5840 );
and ( n5842 , n5837 , n5841 );
xor ( n5843 , n2406 , n4023 );
buf ( n5844 , n5843 );
buf ( n5845 , n5844 );
xor ( n5846 , n4833 , n5772 );
buf ( n5847 , n5846 );
buf ( n5848 , n5847 );
not ( n5849 , n5848 );
and ( n5850 , n5845 , n5849 );
xor ( n5851 , n2582 , n4021 );
buf ( n5852 , n5851 );
buf ( n5853 , n5852 );
xor ( n5854 , n4995 , n5770 );
buf ( n5855 , n5854 );
buf ( n5856 , n5855 );
not ( n5857 , n5856 );
and ( n5858 , n5853 , n5857 );
xor ( n5859 , n2652 , n4019 );
buf ( n5860 , n5859 );
buf ( n5861 , n5860 );
xor ( n5862 , n5436 , n5768 );
buf ( n5863 , n5862 );
buf ( n5864 , n5863 );
not ( n5865 , n5864 );
and ( n5866 , n5861 , n5865 );
xor ( n5867 , n2788 , n4017 );
buf ( n5868 , n5867 );
buf ( n5869 , n5868 );
xor ( n5870 , n5438 , n5767 );
buf ( n5871 , n5870 );
buf ( n5872 , n5871 );
not ( n5873 , n5872 );
and ( n5874 , n5869 , n5873 );
xor ( n5875 , n2950 , n4015 );
buf ( n5876 , n5875 );
buf ( n5877 , n5876 );
xor ( n5878 , n5440 , n5766 );
buf ( n5879 , n5878 );
buf ( n5880 , n5879 );
not ( n5881 , n5880 );
and ( n5882 , n5877 , n5881 );
xor ( n5883 , n3066 , n4013 );
buf ( n5884 , n5883 );
buf ( n5885 , n5884 );
xor ( n5886 , n5442 , n5765 );
buf ( n5887 , n5886 );
buf ( n5888 , n5887 );
not ( n5889 , n5888 );
and ( n5890 , n5885 , n5889 );
xor ( n5891 , n3180 , n4011 );
buf ( n5892 , n5891 );
buf ( n5893 , n5892 );
xor ( n5894 , n5444 , n5764 );
buf ( n5895 , n5894 );
buf ( n5896 , n5895 );
not ( n5897 , n5896 );
and ( n5898 , n5893 , n5897 );
xor ( n5899 , n3256 , n4009 );
buf ( n5900 , n5899 );
buf ( n5901 , n5900 );
xor ( n5902 , n5446 , n5763 );
buf ( n5903 , n5902 );
buf ( n5904 , n5903 );
not ( n5905 , n5904 );
and ( n5906 , n5901 , n5905 );
xor ( n5907 , n3358 , n4007 );
buf ( n5908 , n5907 );
buf ( n5909 , n5908 );
xor ( n5910 , n5448 , n5762 );
buf ( n5911 , n5910 );
buf ( n5912 , n5911 );
not ( n5913 , n5912 );
and ( n5914 , n5909 , n5913 );
xor ( n5915 , n3452 , n4005 );
buf ( n5916 , n5915 );
buf ( n5917 , n5916 );
xor ( n5918 , n5527 , n5760 );
buf ( n5919 , n5918 );
buf ( n5920 , n5919 );
not ( n5921 , n5920 );
and ( n5922 , n5917 , n5921 );
xor ( n5923 , n3528 , n4003 );
buf ( n5924 , n5923 );
buf ( n5925 , n5924 );
xor ( n5926 , n5529 , n5759 );
buf ( n5927 , n5926 );
buf ( n5928 , n5927 );
not ( n5929 , n5928 );
and ( n5930 , n5925 , n5929 );
xor ( n5931 , n3602 , n4001 );
buf ( n5932 , n5931 );
buf ( n5933 , n5932 );
xor ( n5934 , n5531 , n5758 );
buf ( n5935 , n5934 );
buf ( n5936 , n5935 );
not ( n5937 , n5936 );
and ( n5938 , n5933 , n5937 );
xor ( n5939 , n3668 , n3999 );
buf ( n5940 , n5939 );
buf ( n5941 , n5940 );
xor ( n5942 , n5567 , n5756 );
buf ( n5943 , n5942 );
buf ( n5944 , n5943 );
not ( n5945 , n5944 );
and ( n5946 , n5941 , n5945 );
xor ( n5947 , n3724 , n3997 );
buf ( n5948 , n5947 );
buf ( n5949 , n5948 );
xor ( n5950 , n5599 , n5754 );
buf ( n5951 , n5950 );
buf ( n5952 , n5951 );
not ( n5953 , n5952 );
and ( n5954 , n5949 , n5953 );
xor ( n5955 , n3778 , n3995 );
buf ( n5956 , n5955 );
buf ( n5957 , n5956 );
xor ( n5958 , n5624 , n5752 );
buf ( n5959 , n5958 );
buf ( n5960 , n5959 );
not ( n5961 , n5960 );
and ( n5962 , n5957 , n5961 );
xor ( n5963 , n3822 , n3993 );
buf ( n5964 , n5963 );
buf ( n5965 , n5964 );
xor ( n5966 , n5654 , n5750 );
buf ( n5967 , n5966 );
buf ( n5968 , n5967 );
not ( n5969 , n5968 );
and ( n5970 , n5965 , n5969 );
xor ( n5971 , n3864 , n3991 );
buf ( n5972 , n5971 );
buf ( n5973 , n5972 );
xor ( n5974 , n5672 , n5748 );
buf ( n5975 , n5974 );
buf ( n5976 , n5975 );
not ( n5977 , n5976 );
and ( n5978 , n5973 , n5977 );
xor ( n5979 , n3898 , n3989 );
buf ( n5980 , n5979 );
buf ( n5981 , n5980 );
xor ( n5982 , n5689 , n5746 );
buf ( n5983 , n5982 );
buf ( n5984 , n5983 );
not ( n5985 , n5984 );
and ( n5986 , n5981 , n5985 );
xor ( n5987 , n3923 , n3987 );
buf ( n5988 , n5987 );
buf ( n5989 , n5988 );
xor ( n5990 , n5709 , n5744 );
buf ( n5991 , n5990 );
buf ( n5992 , n5991 );
not ( n5993 , n5992 );
and ( n5994 , n5989 , n5993 );
xor ( n5995 , n3939 , n3985 );
buf ( n5996 , n5995 );
buf ( n5997 , n5996 );
xor ( n5998 , n5717 , n5742 );
buf ( n5999 , n5998 );
buf ( n6000 , n5999 );
not ( n6001 , n6000 );
and ( n6002 , n5997 , n6001 );
xor ( n6003 , n3952 , n3983 );
buf ( n6004 , n6003 );
buf ( n6005 , n6004 );
xor ( n6006 , n5724 , n5740 );
buf ( n6007 , n6006 );
buf ( n6008 , n6007 );
not ( n6009 , n6008 );
and ( n6010 , n6005 , n6009 );
xor ( n6011 , n3970 , n3981 );
buf ( n6012 , n6011 );
buf ( n6013 , n6012 );
xor ( n6014 , n5730 , n5738 );
buf ( n6015 , n6014 );
buf ( n6016 , n6015 );
not ( n6017 , n6016 );
and ( n6018 , n6013 , n6017 );
xor ( n6019 , n3978 , n3979 );
buf ( n6020 , n6019 );
buf ( n6021 , n6020 );
xor ( n6022 , n5734 , n5737 );
buf ( n6023 , n6022 );
buf ( n6024 , n6023 );
not ( n6025 , n6024 );
and ( n6026 , n6021 , n6025 );
buf ( n6027 , n6025 );
buf ( n6028 , n6021 );
or ( n6029 , n6026 , n6027 , n6028 );
and ( n6030 , n6017 , n6029 );
and ( n6031 , n6013 , n6029 );
or ( n6032 , n6018 , n6030 , n6031 );
and ( n6033 , n6009 , n6032 );
and ( n6034 , n6005 , n6032 );
or ( n6035 , n6010 , n6033 , n6034 );
and ( n6036 , n6001 , n6035 );
and ( n6037 , n5997 , n6035 );
or ( n6038 , n6002 , n6036 , n6037 );
and ( n6039 , n5993 , n6038 );
and ( n6040 , n5989 , n6038 );
or ( n6041 , n5994 , n6039 , n6040 );
and ( n6042 , n5985 , n6041 );
and ( n6043 , n5981 , n6041 );
or ( n6044 , n5986 , n6042 , n6043 );
and ( n6045 , n5977 , n6044 );
and ( n6046 , n5973 , n6044 );
or ( n6047 , n5978 , n6045 , n6046 );
and ( n6048 , n5969 , n6047 );
and ( n6049 , n5965 , n6047 );
or ( n6050 , n5970 , n6048 , n6049 );
and ( n6051 , n5961 , n6050 );
and ( n6052 , n5957 , n6050 );
or ( n6053 , n5962 , n6051 , n6052 );
and ( n6054 , n5953 , n6053 );
and ( n6055 , n5949 , n6053 );
or ( n6056 , n5954 , n6054 , n6055 );
and ( n6057 , n5945 , n6056 );
and ( n6058 , n5941 , n6056 );
or ( n6059 , n5946 , n6057 , n6058 );
and ( n6060 , n5937 , n6059 );
and ( n6061 , n5933 , n6059 );
or ( n6062 , n5938 , n6060 , n6061 );
and ( n6063 , n5929 , n6062 );
and ( n6064 , n5925 , n6062 );
or ( n6065 , n5930 , n6063 , n6064 );
and ( n6066 , n5921 , n6065 );
and ( n6067 , n5917 , n6065 );
or ( n6068 , n5922 , n6066 , n6067 );
and ( n6069 , n5913 , n6068 );
and ( n6070 , n5909 , n6068 );
or ( n6071 , n5914 , n6069 , n6070 );
and ( n6072 , n5905 , n6071 );
and ( n6073 , n5901 , n6071 );
or ( n6074 , n5906 , n6072 , n6073 );
and ( n6075 , n5897 , n6074 );
and ( n6076 , n5893 , n6074 );
or ( n6077 , n5898 , n6075 , n6076 );
and ( n6078 , n5889 , n6077 );
and ( n6079 , n5885 , n6077 );
or ( n6080 , n5890 , n6078 , n6079 );
and ( n6081 , n5881 , n6080 );
and ( n6082 , n5877 , n6080 );
or ( n6083 , n5882 , n6081 , n6082 );
and ( n6084 , n5873 , n6083 );
and ( n6085 , n5869 , n6083 );
or ( n6086 , n5874 , n6084 , n6085 );
and ( n6087 , n5865 , n6086 );
and ( n6088 , n5861 , n6086 );
or ( n6089 , n5866 , n6087 , n6088 );
and ( n6090 , n5857 , n6089 );
and ( n6091 , n5853 , n6089 );
or ( n6092 , n5858 , n6090 , n6091 );
and ( n6093 , n5849 , n6092 );
and ( n6094 , n5845 , n6092 );
or ( n6095 , n5850 , n6093 , n6094 );
and ( n6096 , n5841 , n6095 );
and ( n6097 , n5837 , n6095 );
or ( n6098 , n5842 , n6096 , n6097 );
and ( n6099 , n5833 , n6098 );
and ( n6100 , n5829 , n6098 );
or ( n6101 , n5834 , n6099 , n6100 );
and ( n6102 , n5825 , n6101 );
and ( n6103 , n5821 , n6101 );
or ( n6104 , n5826 , n6102 , n6103 );
and ( n6105 , n5817 , n6104 );
and ( n6106 , n5813 , n6104 );
or ( n6107 , n5818 , n6105 , n6106 );
and ( n6108 , n5809 , n6107 );
and ( n6109 , n5805 , n6107 );
or ( n6110 , n5810 , n6108 , n6109 );
and ( n6111 , n5801 , n6110 );
and ( n6112 , n5797 , n6110 );
or ( n6113 , n5802 , n6111 , n6112 );
and ( n6114 , n5793 , n6113 );
and ( n6115 , n5789 , n6113 );
or ( n6116 , n5794 , n6114 , n6115 );
and ( n6117 , n5785 , n6116 );
and ( n6118 , n4042 , n6116 );
or ( n6119 , n5786 , n6117 , n6118 );
not ( n6120 , n6119 );
buf ( n6121 , n6120 );
buf ( n6122 , n6121 );
buf ( n6123 , n6120 );
buf ( n6124 , n6123 );
buf ( n6125 , n6120 );
buf ( n6126 , n6125 );
buf ( n6127 , n6120 );
buf ( n6128 , n6127 );
buf ( n6129 , n6120 );
buf ( n6130 , n6129 );
buf ( n6131 , n6120 );
buf ( n6132 , n6131 );
buf ( n6133 , n6120 );
buf ( n6134 , n6133 );
buf ( n6135 , n6120 );
buf ( n6136 , n6135 );
buf ( n6137 , n6120 );
buf ( n6138 , n6137 );
buf ( n6139 , n6120 );
buf ( n6140 , n6139 );
buf ( n6141 , n6120 );
buf ( n6142 , n6141 );
buf ( n6143 , n6120 );
buf ( n6144 , n6143 );
buf ( n6145 , n6120 );
buf ( n6146 , n6145 );
buf ( n6147 , n6120 );
buf ( n6148 , n6147 );
buf ( n6149 , n6120 );
buf ( n6150 , n6149 );
buf ( n6151 , n6120 );
buf ( n6152 , n6151 );
buf ( n6153 , n6120 );
buf ( n6154 , n6153 );
buf ( n6155 , n6120 );
buf ( n6156 , n6155 );
buf ( n6157 , n6120 );
buf ( n6158 , n6157 );
buf ( n6159 , n6120 );
buf ( n6160 , n6159 );
buf ( n6161 , n6120 );
buf ( n6162 , n6161 );
buf ( n6163 , n6120 );
buf ( n6164 , n6163 );
buf ( n6165 , n6120 );
buf ( n6166 , n6165 );
buf ( n6167 , n6120 );
buf ( n6168 , n6167 );
buf ( n6169 , n6120 );
buf ( n6170 , n6169 );
buf ( n6171 , n6120 );
buf ( n6172 , n6171 );
buf ( n6173 , n6120 );
buf ( n6174 , n6173 );
buf ( n6175 , n6120 );
buf ( n6176 , n6175 );
buf ( n6177 , n6120 );
buf ( n6178 , n6177 );
buf ( n6179 , n6120 );
buf ( n6180 , n6179 );
buf ( n6181 , n6120 );
buf ( n6182 , n6181 );
buf ( n6183 , n6120 );
buf ( n6184 , n6183 );
buf ( n6185 , n6120 );
buf ( n6186 , n6185 );
buf ( n6187 , n6120 );
buf ( n6188 , n6187 );
buf ( n6189 , n6120 );
buf ( n6190 , n6189 );
buf ( n6191 , n6120 );
buf ( n6192 , n6191 );
buf ( n6193 , n6120 );
buf ( n6194 , n6193 );
buf ( n6195 , n6120 );
buf ( n6196 , n6195 );
buf ( n6197 , n6120 );
buf ( n6198 , n6197 );
buf ( n6199 , n6120 );
buf ( n6200 , n6199 );
buf ( n6201 , n6120 );
buf ( n6202 , n6201 );
buf ( n6203 , n6120 );
buf ( n6204 , n6203 );
buf ( n6205 , n6120 );
buf ( n6206 , n6205 );
buf ( n6207 , n6120 );
buf ( n6208 , n6207 );
buf ( n6209 , n6120 );
buf ( n6210 , n6209 );
buf ( n6211 , n6120 );
buf ( n6212 , n6211 );
buf ( n6213 , n6120 );
buf ( n6214 , n6213 );
buf ( n6215 , n6120 );
buf ( n6216 , n6215 );
buf ( n6217 , n6120 );
buf ( n6218 , n6217 );
buf ( n6219 , n6120 );
buf ( n6220 , n6219 );
buf ( n6221 , n6120 );
buf ( n6222 , n6221 );
buf ( n6223 , n6120 );
buf ( n6224 , n6223 );
buf ( n6225 , n6120 );
buf ( n6226 , n6225 );
buf ( n6227 , n6120 );
buf ( n6228 , n6227 );
buf ( n6229 , n6120 );
buf ( n6230 , n6229 );
buf ( n6231 , n6120 );
buf ( n6232 , n6231 );
buf ( n6233 , n6120 );
buf ( n6234 , n6233 );
buf ( n6235 , n6120 );
buf ( n6236 , n6235 );
buf ( n6237 , n6120 );
buf ( n6238 , n6237 );
buf ( n6239 , n6120 );
buf ( n6240 , n6239 );
buf ( n6241 , n6120 );
buf ( n6242 , n6241 );
buf ( n6243 , n6120 );
buf ( n6244 , n6243 );
buf ( n6245 , n6120 );
buf ( n6246 , n6245 );
buf ( n6247 , n6120 );
buf ( n6248 , n6247 );
buf ( n6249 , n6120 );
buf ( n6250 , n6249 );
buf ( n6251 , n6120 );
buf ( n6252 , n6251 );
buf ( n6253 , n6120 );
buf ( n6254 , n6253 );
buf ( n6255 , n6120 );
buf ( n6256 , n6255 );
buf ( n6257 , n6120 );
buf ( n6258 , n6257 );
buf ( n6259 , n6120 );
buf ( n6260 , n6259 );
buf ( n6261 , n6120 );
buf ( n6262 , n6261 );
buf ( n6263 , n6120 );
buf ( n6264 , n6263 );
buf ( n6265 , n6120 );
buf ( n6266 , n6265 );
buf ( n6267 , n6120 );
buf ( n6268 , n6267 );
buf ( n6269 , n6120 );
buf ( n6270 , n6269 );
buf ( n6271 , n6120 );
buf ( n6272 , n6271 );
buf ( n6273 , n6120 );
buf ( n6274 , n6273 );
buf ( n6275 , n6120 );
buf ( n6276 , n6275 );
buf ( n6277 , n6120 );
buf ( n6278 , n6277 );
buf ( n6279 , n6120 );
buf ( n6280 , n6279 );
buf ( n6281 , n6120 );
buf ( n6282 , n6281 );
buf ( n6283 , n6120 );
buf ( n6284 , n6283 );
buf ( n6285 , n6120 );
buf ( n6286 , n6285 );
buf ( n6287 , n6120 );
buf ( n6288 , n6287 );
buf ( n6289 , n6120 );
buf ( n6290 , n6289 );
buf ( n6291 , n6120 );
buf ( n6292 , n6291 );
buf ( n6293 , n6120 );
buf ( n6294 , n6293 );
buf ( n6295 , n6120 );
buf ( n6296 , n6295 );
buf ( n6297 , n6120 );
buf ( n6298 , n6297 );
buf ( n6299 , n6120 );
buf ( n6300 , n6299 );
buf ( n6301 , n6120 );
buf ( n6302 , n6301 );
buf ( n6303 , n6120 );
buf ( n6304 , n6303 );
buf ( n6305 , n6120 );
buf ( n6306 , n6305 );
buf ( n6307 , n6120 );
buf ( n6308 , n6307 );
buf ( n6309 , n6120 );
buf ( n6310 , n6309 );
xor ( n6311 , n4042 , n5785 );
xor ( n6312 , n6311 , n6116 );
buf ( n6313 , n6312 );
buf ( n6314 , n6313 );
xor ( n6315 , n5789 , n5793 );
xor ( n6316 , n6315 , n6113 );
buf ( n6317 , n6316 );
buf ( n6318 , n6317 );
xor ( n6319 , n5797 , n5801 );
xor ( n6320 , n6319 , n6110 );
buf ( n6321 , n6320 );
buf ( n6322 , n6321 );
xor ( n6323 , n5805 , n5809 );
xor ( n6324 , n6323 , n6107 );
buf ( n6325 , n6324 );
buf ( n6326 , n6325 );
xor ( n6327 , n5813 , n5817 );
xor ( n6328 , n6327 , n6104 );
buf ( n6329 , n6328 );
buf ( n6330 , n6329 );
xor ( n6331 , n5821 , n5825 );
xor ( n6332 , n6331 , n6101 );
buf ( n6333 , n6332 );
buf ( n6334 , n6333 );
xor ( n6335 , n5829 , n5833 );
xor ( n6336 , n6335 , n6098 );
buf ( n6337 , n6336 );
buf ( n6338 , n6337 );
xor ( n6339 , n5837 , n5841 );
xor ( n6340 , n6339 , n6095 );
buf ( n6341 , n6340 );
buf ( n6342 , n6341 );
xor ( n6343 , n5845 , n5849 );
xor ( n6344 , n6343 , n6092 );
buf ( n6345 , n6344 );
buf ( n6346 , n6345 );
xor ( n6347 , n5853 , n5857 );
xor ( n6348 , n6347 , n6089 );
buf ( n6349 , n6348 );
buf ( n6350 , n6349 );
xor ( n6351 , n5861 , n5865 );
xor ( n6352 , n6351 , n6086 );
buf ( n6353 , n6352 );
buf ( n6354 , n6353 );
xor ( n6355 , n5869 , n5873 );
xor ( n6356 , n6355 , n6083 );
buf ( n6357 , n6356 );
buf ( n6358 , n6357 );
xor ( n6359 , n5877 , n5881 );
xor ( n6360 , n6359 , n6080 );
buf ( n6361 , n6360 );
buf ( n6362 , n6361 );
xor ( n6363 , n5885 , n5889 );
xor ( n6364 , n6363 , n6077 );
buf ( n6365 , n6364 );
buf ( n6366 , n6365 );
xor ( n6367 , n5893 , n5897 );
xor ( n6368 , n6367 , n6074 );
buf ( n6369 , n6368 );
buf ( n6370 , n6369 );
xor ( n6371 , n5901 , n5905 );
xor ( n6372 , n6371 , n6071 );
buf ( n6373 , n6372 );
buf ( n6374 , n6373 );
xor ( n6375 , n5909 , n5913 );
xor ( n6376 , n6375 , n6068 );
buf ( n6377 , n6376 );
buf ( n6378 , n6377 );
buf ( n6379 , n576 );
and ( n6380 , n6378 , n6379 );
xor ( n6381 , n5917 , n5921 );
xor ( n6382 , n6381 , n6065 );
buf ( n6383 , n6382 );
buf ( n6384 , n6383 );
buf ( n6385 , n577 );
and ( n6386 , n6384 , n6385 );
xor ( n6387 , n5925 , n5929 );
xor ( n6388 , n6387 , n6062 );
buf ( n6389 , n6388 );
buf ( n6390 , n6389 );
buf ( n6391 , n578 );
and ( n6392 , n6390 , n6391 );
xor ( n6393 , n5933 , n5937 );
xor ( n6394 , n6393 , n6059 );
buf ( n6395 , n6394 );
buf ( n6396 , n6395 );
buf ( n6397 , n579 );
and ( n6398 , n6396 , n6397 );
xor ( n6399 , n5941 , n5945 );
xor ( n6400 , n6399 , n6056 );
buf ( n6401 , n6400 );
buf ( n6402 , n6401 );
buf ( n6403 , n580 );
and ( n6404 , n6402 , n6403 );
xor ( n6405 , n5949 , n5953 );
xor ( n6406 , n6405 , n6053 );
buf ( n6407 , n6406 );
buf ( n6408 , n6407 );
buf ( n6409 , n581 );
and ( n6410 , n6408 , n6409 );
xor ( n6411 , n5957 , n5961 );
xor ( n6412 , n6411 , n6050 );
buf ( n6413 , n6412 );
buf ( n6414 , n6413 );
buf ( n6415 , n582 );
and ( n6416 , n6414 , n6415 );
xor ( n6417 , n5965 , n5969 );
xor ( n6418 , n6417 , n6047 );
buf ( n6419 , n6418 );
buf ( n6420 , n6419 );
buf ( n6421 , n583 );
and ( n6422 , n6420 , n6421 );
xor ( n6423 , n5973 , n5977 );
xor ( n6424 , n6423 , n6044 );
buf ( n6425 , n6424 );
buf ( n6426 , n6425 );
buf ( n6427 , n584 );
and ( n6428 , n6426 , n6427 );
xor ( n6429 , n5981 , n5985 );
xor ( n6430 , n6429 , n6041 );
buf ( n6431 , n6430 );
buf ( n6432 , n6431 );
buf ( n6433 , n585 );
and ( n6434 , n6432 , n6433 );
xor ( n6435 , n5989 , n5993 );
xor ( n6436 , n6435 , n6038 );
buf ( n6437 , n6436 );
buf ( n6438 , n6437 );
buf ( n6439 , n586 );
and ( n6440 , n6438 , n6439 );
xor ( n6441 , n5997 , n6001 );
xor ( n6442 , n6441 , n6035 );
buf ( n6443 , n6442 );
buf ( n6444 , n6443 );
buf ( n6445 , n587 );
and ( n6446 , n6444 , n6445 );
xor ( n6447 , n6005 , n6009 );
xor ( n6448 , n6447 , n6032 );
buf ( n6449 , n6448 );
buf ( n6450 , n6449 );
buf ( n6451 , n588 );
and ( n6452 , n6450 , n6451 );
xor ( n6453 , n6013 , n6017 );
xor ( n6454 , n6453 , n6029 );
buf ( n6455 , n6454 );
buf ( n6456 , n6455 );
buf ( n6457 , n589 );
and ( n6458 , n6456 , n6457 );
xor ( n6459 , n6021 , n6025 );
not ( n6460 , n6459 );
buf ( n6461 , n6460 );
buf ( n6462 , n6461 );
buf ( n6463 , n590 );
and ( n6464 , n6462 , n6463 );
buf ( n6465 , n6464 );
and ( n6466 , n6457 , n6465 );
and ( n6467 , n6456 , n6465 );
or ( n6468 , n6458 , n6466 , n6467 );
and ( n6469 , n6451 , n6468 );
and ( n6470 , n6450 , n6468 );
or ( n6471 , n6452 , n6469 , n6470 );
and ( n6472 , n6445 , n6471 );
and ( n6473 , n6444 , n6471 );
or ( n6474 , n6446 , n6472 , n6473 );
and ( n6475 , n6439 , n6474 );
and ( n6476 , n6438 , n6474 );
or ( n6477 , n6440 , n6475 , n6476 );
and ( n6478 , n6433 , n6477 );
and ( n6479 , n6432 , n6477 );
or ( n6480 , n6434 , n6478 , n6479 );
and ( n6481 , n6427 , n6480 );
and ( n6482 , n6426 , n6480 );
or ( n6483 , n6428 , n6481 , n6482 );
and ( n6484 , n6421 , n6483 );
and ( n6485 , n6420 , n6483 );
or ( n6486 , n6422 , n6484 , n6485 );
and ( n6487 , n6415 , n6486 );
and ( n6488 , n6414 , n6486 );
or ( n6489 , n6416 , n6487 , n6488 );
and ( n6490 , n6409 , n6489 );
and ( n6491 , n6408 , n6489 );
or ( n6492 , n6410 , n6490 , n6491 );
and ( n6493 , n6403 , n6492 );
and ( n6494 , n6402 , n6492 );
or ( n6495 , n6404 , n6493 , n6494 );
and ( n6496 , n6397 , n6495 );
and ( n6497 , n6396 , n6495 );
or ( n6498 , n6398 , n6496 , n6497 );
and ( n6499 , n6391 , n6498 );
and ( n6500 , n6390 , n6498 );
or ( n6501 , n6392 , n6499 , n6500 );
and ( n6502 , n6385 , n6501 );
and ( n6503 , n6384 , n6501 );
or ( n6504 , n6386 , n6502 , n6503 );
and ( n6505 , n6379 , n6504 );
and ( n6506 , n6378 , n6504 );
or ( n6507 , n6380 , n6505 , n6506 );
and ( n6508 , n6374 , n6507 );
and ( n6509 , n6370 , n6508 );
and ( n6510 , n6366 , n6509 );
and ( n6511 , n6362 , n6510 );
and ( n6512 , n6358 , n6511 );
and ( n6513 , n6354 , n6512 );
and ( n6514 , n6350 , n6513 );
and ( n6515 , n6346 , n6514 );
and ( n6516 , n6342 , n6515 );
and ( n6517 , n6338 , n6516 );
and ( n6518 , n6334 , n6517 );
and ( n6519 , n6330 , n6518 );
and ( n6520 , n6326 , n6519 );
and ( n6521 , n6322 , n6520 );
and ( n6522 , n6318 , n6521 );
and ( n6523 , n6314 , n6522 );
and ( n6524 , n6310 , n6523 );
and ( n6525 , n6308 , n6524 );
and ( n6526 , n6306 , n6525 );
and ( n6527 , n6304 , n6526 );
and ( n6528 , n6302 , n6527 );
and ( n6529 , n6300 , n6528 );
and ( n6530 , n6298 , n6529 );
and ( n6531 , n6296 , n6530 );
and ( n6532 , n6294 , n6531 );
and ( n6533 , n6292 , n6532 );
and ( n6534 , n6290 , n6533 );
and ( n6535 , n6288 , n6534 );
and ( n6536 , n6286 , n6535 );
and ( n6537 , n6284 , n6536 );
and ( n6538 , n6282 , n6537 );
and ( n6539 , n6280 , n6538 );
and ( n6540 , n6278 , n6539 );
and ( n6541 , n6276 , n6540 );
and ( n6542 , n6274 , n6541 );
and ( n6543 , n6272 , n6542 );
and ( n6544 , n6270 , n6543 );
and ( n6545 , n6268 , n6544 );
and ( n6546 , n6266 , n6545 );
and ( n6547 , n6264 , n6546 );
and ( n6548 , n6262 , n6547 );
and ( n6549 , n6260 , n6548 );
and ( n6550 , n6258 , n6549 );
and ( n6551 , n6256 , n6550 );
and ( n6552 , n6254 , n6551 );
and ( n6553 , n6252 , n6552 );
and ( n6554 , n6250 , n6553 );
and ( n6555 , n6248 , n6554 );
and ( n6556 , n6246 , n6555 );
and ( n6557 , n6244 , n6556 );
and ( n6558 , n6242 , n6557 );
and ( n6559 , n6240 , n6558 );
and ( n6560 , n6238 , n6559 );
and ( n6561 , n6236 , n6560 );
and ( n6562 , n6234 , n6561 );
and ( n6563 , n6232 , n6562 );
and ( n6564 , n6230 , n6563 );
and ( n6565 , n6228 , n6564 );
and ( n6566 , n6226 , n6565 );
and ( n6567 , n6224 , n6566 );
and ( n6568 , n6222 , n6567 );
and ( n6569 , n6220 , n6568 );
and ( n6570 , n6218 , n6569 );
and ( n6571 , n6216 , n6570 );
and ( n6572 , n6214 , n6571 );
and ( n6573 , n6212 , n6572 );
and ( n6574 , n6210 , n6573 );
and ( n6575 , n6208 , n6574 );
and ( n6576 , n6206 , n6575 );
and ( n6577 , n6204 , n6576 );
and ( n6578 , n6202 , n6577 );
and ( n6579 , n6200 , n6578 );
and ( n6580 , n6198 , n6579 );
and ( n6581 , n6196 , n6580 );
and ( n6582 , n6194 , n6581 );
and ( n6583 , n6192 , n6582 );
and ( n6584 , n6190 , n6583 );
and ( n6585 , n6188 , n6584 );
and ( n6586 , n6186 , n6585 );
and ( n6587 , n6184 , n6586 );
and ( n6588 , n6182 , n6587 );
and ( n6589 , n6180 , n6588 );
and ( n6590 , n6178 , n6589 );
and ( n6591 , n6176 , n6590 );
and ( n6592 , n6174 , n6591 );
and ( n6593 , n6172 , n6592 );
and ( n6594 , n6170 , n6593 );
and ( n6595 , n6168 , n6594 );
and ( n6596 , n6166 , n6595 );
and ( n6597 , n6164 , n6596 );
and ( n6598 , n6162 , n6597 );
and ( n6599 , n6160 , n6598 );
and ( n6600 , n6158 , n6599 );
and ( n6601 , n6156 , n6600 );
and ( n6602 , n6154 , n6601 );
and ( n6603 , n6152 , n6602 );
and ( n6604 , n6150 , n6603 );
and ( n6605 , n6148 , n6604 );
and ( n6606 , n6146 , n6605 );
and ( n6607 , n6144 , n6606 );
and ( n6608 , n6142 , n6607 );
and ( n6609 , n6140 , n6608 );
and ( n6610 , n6138 , n6609 );
and ( n6611 , n6136 , n6610 );
and ( n6612 , n6134 , n6611 );
and ( n6613 , n6132 , n6612 );
and ( n6614 , n6130 , n6613 );
and ( n6615 , n6128 , n6614 );
and ( n6616 , n6126 , n6615 );
and ( n6617 , n6124 , n6616 );
xor ( n6618 , n6122 , n6617 );
buf ( n6619 , n6618 );
buf ( n6620 , n6619 );
xor ( n6621 , n6124 , n6616 );
buf ( n6622 , n6621 );
buf ( n6623 , n6622 );
xor ( n6624 , n6126 , n6615 );
buf ( n6625 , n6624 );
buf ( n6626 , n6625 );
xor ( n6627 , n6128 , n6614 );
buf ( n6628 , n6627 );
buf ( n6629 , n6628 );
xor ( n6630 , n6130 , n6613 );
buf ( n6631 , n6630 );
buf ( n6632 , n6631 );
xor ( n6633 , n6132 , n6612 );
buf ( n6634 , n6633 );
buf ( n6635 , n6634 );
xor ( n6636 , n6134 , n6611 );
buf ( n6637 , n6636 );
buf ( n6638 , n6637 );
xor ( n6639 , n6136 , n6610 );
buf ( n6640 , n6639 );
buf ( n6641 , n6640 );
xor ( n6642 , n6138 , n6609 );
buf ( n6643 , n6642 );
buf ( n6644 , n6643 );
xor ( n6645 , n6140 , n6608 );
buf ( n6646 , n6645 );
buf ( n6647 , n6646 );
xor ( n6648 , n6142 , n6607 );
buf ( n6649 , n6648 );
buf ( n6650 , n6649 );
xor ( n6651 , n6144 , n6606 );
buf ( n6652 , n6651 );
buf ( n6653 , n6652 );
xor ( n6654 , n6146 , n6605 );
buf ( n6655 , n6654 );
buf ( n6656 , n6655 );
xor ( n6657 , n6148 , n6604 );
buf ( n6658 , n6657 );
buf ( n6659 , n6658 );
xor ( n6660 , n6150 , n6603 );
buf ( n6661 , n6660 );
buf ( n6662 , n6661 );
xor ( n6663 , n6152 , n6602 );
buf ( n6664 , n6663 );
buf ( n6665 , n6664 );
xor ( n6666 , n6154 , n6601 );
buf ( n6667 , n6666 );
buf ( n6668 , n6667 );
xor ( n6669 , n6156 , n6600 );
buf ( n6670 , n6669 );
buf ( n6671 , n6670 );
xor ( n6672 , n6158 , n6599 );
buf ( n6673 , n6672 );
buf ( n6674 , n6673 );
xor ( n6675 , n6160 , n6598 );
buf ( n6676 , n6675 );
buf ( n6677 , n6676 );
xor ( n6678 , n6162 , n6597 );
buf ( n6679 , n6678 );
buf ( n6680 , n6679 );
xor ( n6681 , n6164 , n6596 );
buf ( n6682 , n6681 );
buf ( n6683 , n6682 );
xor ( n6684 , n6166 , n6595 );
buf ( n6685 , n6684 );
buf ( n6686 , n6685 );
xor ( n6687 , n6168 , n6594 );
buf ( n6688 , n6687 );
buf ( n6689 , n6688 );
xor ( n6690 , n6170 , n6593 );
buf ( n6691 , n6690 );
buf ( n6692 , n6691 );
xor ( n6693 , n6172 , n6592 );
buf ( n6694 , n6693 );
buf ( n6695 , n6694 );
xor ( n6696 , n6174 , n6591 );
buf ( n6697 , n6696 );
buf ( n6698 , n6697 );
xor ( n6699 , n6176 , n6590 );
buf ( n6700 , n6699 );
buf ( n6701 , n6700 );
xor ( n6702 , n6178 , n6589 );
buf ( n6703 , n6702 );
buf ( n6704 , n6703 );
xor ( n6705 , n6180 , n6588 );
buf ( n6706 , n6705 );
buf ( n6707 , n6706 );
xor ( n6708 , n6182 , n6587 );
buf ( n6709 , n6708 );
buf ( n6710 , n6709 );
xor ( n6711 , n6184 , n6586 );
buf ( n6712 , n6711 );
buf ( n6713 , n6712 );
xor ( n6714 , n6186 , n6585 );
buf ( n6715 , n6714 );
buf ( n6716 , n6715 );
xor ( n6717 , n6188 , n6584 );
buf ( n6718 , n6717 );
buf ( n6719 , n6718 );
xor ( n6720 , n6190 , n6583 );
buf ( n6721 , n6720 );
buf ( n6722 , n6721 );
xor ( n6723 , n6192 , n6582 );
buf ( n6724 , n6723 );
buf ( n6725 , n6724 );
xor ( n6726 , n6194 , n6581 );
buf ( n6727 , n6726 );
buf ( n6728 , n6727 );
xor ( n6729 , n6196 , n6580 );
buf ( n6730 , n6729 );
buf ( n6731 , n6730 );
xor ( n6732 , n6198 , n6579 );
buf ( n6733 , n6732 );
buf ( n6734 , n6733 );
xor ( n6735 , n6200 , n6578 );
buf ( n6736 , n6735 );
buf ( n6737 , n6736 );
xor ( n6738 , n6202 , n6577 );
buf ( n6739 , n6738 );
buf ( n6740 , n6739 );
xor ( n6741 , n6204 , n6576 );
buf ( n6742 , n6741 );
buf ( n6743 , n6742 );
xor ( n6744 , n6206 , n6575 );
buf ( n6745 , n6744 );
buf ( n6746 , n6745 );
xor ( n6747 , n6208 , n6574 );
buf ( n6748 , n6747 );
buf ( n6749 , n6748 );
xor ( n6750 , n6210 , n6573 );
buf ( n6751 , n6750 );
buf ( n6752 , n6751 );
xor ( n6753 , n6212 , n6572 );
buf ( n6754 , n6753 );
buf ( n6755 , n6754 );
xor ( n6756 , n6214 , n6571 );
buf ( n6757 , n6756 );
buf ( n6758 , n6757 );
xor ( n6759 , n6216 , n6570 );
buf ( n6760 , n6759 );
buf ( n6761 , n6760 );
xor ( n6762 , n6218 , n6569 );
buf ( n6763 , n6762 );
buf ( n6764 , n6763 );
xor ( n6765 , n6220 , n6568 );
buf ( n6766 , n6765 );
buf ( n6767 , n6766 );
xor ( n6768 , n6222 , n6567 );
buf ( n6769 , n6768 );
buf ( n6770 , n6769 );
xor ( n6771 , n6224 , n6566 );
buf ( n6772 , n6771 );
buf ( n6773 , n6772 );
xor ( n6774 , n6226 , n6565 );
buf ( n6775 , n6774 );
buf ( n6776 , n6775 );
xor ( n6777 , n6228 , n6564 );
buf ( n6778 , n6777 );
buf ( n6779 , n6778 );
xor ( n6780 , n6230 , n6563 );
buf ( n6781 , n6780 );
buf ( n6782 , n6781 );
xor ( n6783 , n6232 , n6562 );
buf ( n6784 , n6783 );
buf ( n6785 , n6784 );
xor ( n6786 , n6234 , n6561 );
buf ( n6787 , n6786 );
buf ( n6788 , n6787 );
xor ( n6789 , n6236 , n6560 );
buf ( n6790 , n6789 );
buf ( n6791 , n6790 );
xor ( n6792 , n6238 , n6559 );
buf ( n6793 , n6792 );
buf ( n6794 , n6793 );
xor ( n6795 , n6240 , n6558 );
buf ( n6796 , n6795 );
buf ( n6797 , n6796 );
xor ( n6798 , n6242 , n6557 );
buf ( n6799 , n6798 );
buf ( n6800 , n6799 );
xor ( n6801 , n6244 , n6556 );
buf ( n6802 , n6801 );
buf ( n6803 , n6802 );
xor ( n6804 , n6246 , n6555 );
buf ( n6805 , n6804 );
buf ( n6806 , n6805 );
xor ( n6807 , n6248 , n6554 );
buf ( n6808 , n6807 );
buf ( n6809 , n6808 );
xor ( n6810 , n6250 , n6553 );
buf ( n6811 , n6810 );
buf ( n6812 , n6811 );
xor ( n6813 , n6252 , n6552 );
buf ( n6814 , n6813 );
buf ( n6815 , n6814 );
xor ( n6816 , n6254 , n6551 );
buf ( n6817 , n6816 );
buf ( n6818 , n6817 );
xor ( n6819 , n6256 , n6550 );
buf ( n6820 , n6819 );
buf ( n6821 , n6820 );
xor ( n6822 , n6258 , n6549 );
buf ( n6823 , n6822 );
buf ( n6824 , n6823 );
xor ( n6825 , n6260 , n6548 );
buf ( n6826 , n6825 );
buf ( n6827 , n6826 );
xor ( n6828 , n6262 , n6547 );
buf ( n6829 , n6828 );
buf ( n6830 , n6829 );
xor ( n6831 , n6264 , n6546 );
buf ( n6832 , n6831 );
buf ( n6833 , n6832 );
xor ( n6834 , n6266 , n6545 );
buf ( n6835 , n6834 );
buf ( n6836 , n6835 );
xor ( n6837 , n6268 , n6544 );
buf ( n6838 , n6837 );
buf ( n6839 , n6838 );
xor ( n6840 , n6270 , n6543 );
buf ( n6841 , n6840 );
buf ( n6842 , n6841 );
xor ( n6843 , n6272 , n6542 );
buf ( n6844 , n6843 );
buf ( n6845 , n6844 );
xor ( n6846 , n6274 , n6541 );
buf ( n6847 , n6846 );
buf ( n6848 , n6847 );
xor ( n6849 , n6276 , n6540 );
buf ( n6850 , n6849 );
buf ( n6851 , n6850 );
xor ( n6852 , n6278 , n6539 );
buf ( n6853 , n6852 );
buf ( n6854 , n6853 );
xor ( n6855 , n6280 , n6538 );
buf ( n6856 , n6855 );
buf ( n6857 , n6856 );
xor ( n6858 , n6282 , n6537 );
buf ( n6859 , n6858 );
buf ( n6860 , n6859 );
xor ( n6861 , n6284 , n6536 );
buf ( n6862 , n6861 );
buf ( n6863 , n6862 );
xor ( n6864 , n6286 , n6535 );
buf ( n6865 , n6864 );
buf ( n6866 , n6865 );
xor ( n6867 , n6288 , n6534 );
buf ( n6868 , n6867 );
buf ( n6869 , n6868 );
xor ( n6870 , n6290 , n6533 );
buf ( n6871 , n6870 );
buf ( n6872 , n6871 );
xor ( n6873 , n6292 , n6532 );
buf ( n6874 , n6873 );
buf ( n6875 , n6874 );
xor ( n6876 , n6294 , n6531 );
buf ( n6877 , n6876 );
buf ( n6878 , n6877 );
xor ( n6879 , n6296 , n6530 );
buf ( n6880 , n6879 );
buf ( n6881 , n6880 );
xor ( n6882 , n6298 , n6529 );
buf ( n6883 , n6882 );
buf ( n6884 , n6883 );
xor ( n6885 , n6300 , n6528 );
buf ( n6886 , n6885 );
buf ( n6887 , n6886 );
xor ( n6888 , n6302 , n6527 );
buf ( n6889 , n6888 );
buf ( n6890 , n6889 );
xor ( n6891 , n6304 , n6526 );
buf ( n6892 , n6891 );
buf ( n6893 , n6892 );
xor ( n6894 , n6306 , n6525 );
buf ( n6895 , n6894 );
buf ( n6896 , n6895 );
xor ( n6897 , n6308 , n6524 );
buf ( n6898 , n6897 );
buf ( n6899 , n6898 );
xor ( n6900 , n6310 , n6523 );
buf ( n6901 , n6900 );
buf ( n6902 , n6901 );
xor ( n6903 , n6314 , n6522 );
buf ( n6904 , n6903 );
buf ( n6905 , n6904 );
xor ( n6906 , n6318 , n6521 );
buf ( n6907 , n6906 );
buf ( n6908 , n6907 );
xor ( n6909 , n6322 , n6520 );
buf ( n6910 , n6909 );
buf ( n6911 , n6910 );
xor ( n6912 , n6326 , n6519 );
buf ( n6913 , n6912 );
buf ( n6914 , n6913 );
xor ( n6915 , n6330 , n6518 );
buf ( n6916 , n6915 );
buf ( n6917 , n6916 );
xor ( n6918 , n6334 , n6517 );
buf ( n6919 , n6918 );
buf ( n6920 , n6919 );
xor ( n6921 , n6338 , n6516 );
buf ( n6922 , n6921 );
buf ( n6923 , n6922 );
xor ( n6924 , n6342 , n6515 );
buf ( n6925 , n6924 );
buf ( n6926 , n6925 );
xor ( n6927 , n6346 , n6514 );
buf ( n6928 , n6927 );
buf ( n6929 , n6928 );
xor ( n6930 , n6350 , n6513 );
buf ( n6931 , n6930 );
buf ( n6932 , n6931 );
xor ( n6933 , n6354 , n6512 );
buf ( n6934 , n6933 );
buf ( n6935 , n6934 );
xor ( n6936 , n6358 , n6511 );
buf ( n6937 , n6936 );
buf ( n6938 , n6937 );
xor ( n6939 , n6362 , n6510 );
buf ( n6940 , n6939 );
buf ( n6941 , n6940 );
xor ( n6942 , n6366 , n6509 );
buf ( n6943 , n6942 );
buf ( n6944 , n6943 );
xor ( n6945 , n6370 , n6508 );
buf ( n6946 , n6945 );
buf ( n6947 , n6946 );
xor ( n6948 , n6374 , n6507 );
buf ( n6949 , n6948 );
buf ( n6950 , n6949 );
xor ( n6951 , n6378 , n6379 );
xor ( n6952 , n6951 , n6504 );
buf ( n6953 , n6952 );
buf ( n6954 , n6953 );
xor ( n6955 , n6384 , n6385 );
xor ( n6956 , n6955 , n6501 );
buf ( n6957 , n6956 );
buf ( n6958 , n6957 );
xor ( n6959 , n6390 , n6391 );
xor ( n6960 , n6959 , n6498 );
buf ( n6961 , n6960 );
buf ( n6962 , n6961 );
xor ( n6963 , n6396 , n6397 );
xor ( n6964 , n6963 , n6495 );
buf ( n6965 , n6964 );
buf ( n6966 , n6965 );
xor ( n6967 , n6402 , n6403 );
xor ( n6968 , n6967 , n6492 );
buf ( n6969 , n6968 );
buf ( n6970 , n6969 );
xor ( n6971 , n6408 , n6409 );
xor ( n6972 , n6971 , n6489 );
buf ( n6973 , n6972 );
buf ( n6974 , n6973 );
xor ( n6975 , n6414 , n6415 );
xor ( n6976 , n6975 , n6486 );
buf ( n6977 , n6976 );
buf ( n6978 , n6977 );
xor ( n6979 , n6420 , n6421 );
xor ( n6980 , n6979 , n6483 );
buf ( n6981 , n6980 );
buf ( n6982 , n6981 );
xor ( n6983 , n6426 , n6427 );
xor ( n6984 , n6983 , n6480 );
buf ( n6985 , n6984 );
buf ( n6986 , n6985 );
xor ( n6987 , n6432 , n6433 );
xor ( n6988 , n6987 , n6477 );
buf ( n6989 , n6988 );
buf ( n6990 , n6989 );
xor ( n6991 , n6438 , n6439 );
xor ( n6992 , n6991 , n6474 );
buf ( n6993 , n6992 );
buf ( n6994 , n6993 );
xor ( n6995 , n6444 , n6445 );
xor ( n6996 , n6995 , n6471 );
buf ( n6997 , n6996 );
buf ( n6998 , n6997 );
xor ( n6999 , n6450 , n6451 );
xor ( n7000 , n6999 , n6468 );
buf ( n7001 , n7000 );
buf ( n7002 , n7001 );
xor ( n7003 , n6456 , n6457 );
xor ( n7004 , n7003 , n6465 );
buf ( n7005 , n7004 );
buf ( n7006 , n7005 );
xor ( n7007 , n6462 , n6463 );
buf ( n7008 , n7007 );
buf ( n7009 , n7008 );
buf ( n7010 , n7009 );
buf ( n7011 , n591 );
buf ( n7012 , n7011 );
buf ( n7013 , n7012 );
buf ( n7014 , n7013 );
and ( n7015 , n816 , n7010 );
and ( n7016 , n816 , n7014 );
and ( n7017 , n817 , n7010 );
and ( n7018 , n7016 , n7017 );
xor ( n7019 , n7016 , n7017 );
and ( n7020 , n817 , n7014 );
and ( n7021 , n818 , n7010 );
and ( n7022 , n7020 , n7021 );
xor ( n7023 , n7020 , n7021 );
and ( n7024 , n818 , n7014 );
and ( n7025 , n819 , n7010 );
and ( n7026 , n7024 , n7025 );
xor ( n7027 , n7024 , n7025 );
and ( n7028 , n819 , n7014 );
and ( n7029 , n820 , n7010 );
and ( n7030 , n7028 , n7029 );
xor ( n7031 , n7028 , n7029 );
and ( n7032 , n820 , n7014 );
and ( n7033 , n821 , n7010 );
and ( n7034 , n7032 , n7033 );
xor ( n7035 , n7032 , n7033 );
and ( n7036 , n821 , n7014 );
and ( n7037 , n822 , n7010 );
and ( n7038 , n7036 , n7037 );
xor ( n7039 , n7036 , n7037 );
and ( n7040 , n822 , n7014 );
and ( n7041 , n823 , n7010 );
and ( n7042 , n7040 , n7041 );
xor ( n7043 , n7040 , n7041 );
and ( n7044 , n823 , n7014 );
and ( n7045 , n824 , n7010 );
and ( n7046 , n7044 , n7045 );
xor ( n7047 , n7044 , n7045 );
and ( n7048 , n824 , n7014 );
and ( n7049 , n825 , n7010 );
and ( n7050 , n7048 , n7049 );
xor ( n7051 , n7048 , n7049 );
and ( n7052 , n825 , n7014 );
and ( n7053 , n826 , n7010 );
and ( n7054 , n7052 , n7053 );
xor ( n7055 , n7052 , n7053 );
and ( n7056 , n826 , n7014 );
and ( n7057 , n827 , n7010 );
and ( n7058 , n7056 , n7057 );
xor ( n7059 , n7056 , n7057 );
and ( n7060 , n827 , n7014 );
and ( n7061 , n828 , n7010 );
and ( n7062 , n7060 , n7061 );
xor ( n7063 , n7060 , n7061 );
and ( n7064 , n828 , n7014 );
and ( n7065 , n829 , n7010 );
and ( n7066 , n7064 , n7065 );
xor ( n7067 , n7064 , n7065 );
and ( n7068 , n829 , n7014 );
and ( n7069 , n830 , n7010 );
and ( n7070 , n7068 , n7069 );
xor ( n7071 , n7068 , n7069 );
and ( n7072 , n830 , n7014 );
and ( n7073 , n831 , n7010 );
and ( n7074 , n7072 , n7073 );
and ( n7075 , n7071 , n7074 );
or ( n7076 , n7070 , n7075 );
and ( n7077 , n7067 , n7076 );
or ( n7078 , n7066 , n7077 );
and ( n7079 , n7063 , n7078 );
or ( n7080 , n7062 , n7079 );
and ( n7081 , n7059 , n7080 );
or ( n7082 , n7058 , n7081 );
and ( n7083 , n7055 , n7082 );
or ( n7084 , n7054 , n7083 );
and ( n7085 , n7051 , n7084 );
or ( n7086 , n7050 , n7085 );
and ( n7087 , n7047 , n7086 );
or ( n7088 , n7046 , n7087 );
and ( n7089 , n7043 , n7088 );
or ( n7090 , n7042 , n7089 );
and ( n7091 , n7039 , n7090 );
or ( n7092 , n7038 , n7091 );
and ( n7093 , n7035 , n7092 );
or ( n7094 , n7034 , n7093 );
and ( n7095 , n7031 , n7094 );
or ( n7096 , n7030 , n7095 );
and ( n7097 , n7027 , n7096 );
or ( n7098 , n7026 , n7097 );
and ( n7099 , n7023 , n7098 );
or ( n7100 , n7022 , n7099 );
and ( n7101 , n7019 , n7100 );
or ( n7102 , n7018 , n7101 );
and ( n7103 , n7015 , n7102 );
and ( n7104 , n816 , n7006 );
and ( n7105 , n7103 , n7104 );
xor ( n7106 , n7103 , n7104 );
xor ( n7107 , n7015 , n7102 );
and ( n7108 , n817 , n7006 );
and ( n7109 , n7107 , n7108 );
xor ( n7110 , n7107 , n7108 );
xor ( n7111 , n7019 , n7100 );
and ( n7112 , n818 , n7006 );
and ( n7113 , n7111 , n7112 );
xor ( n7114 , n7111 , n7112 );
xor ( n7115 , n7023 , n7098 );
and ( n7116 , n819 , n7006 );
and ( n7117 , n7115 , n7116 );
xor ( n7118 , n7115 , n7116 );
xor ( n7119 , n7027 , n7096 );
and ( n7120 , n820 , n7006 );
and ( n7121 , n7119 , n7120 );
xor ( n7122 , n7119 , n7120 );
xor ( n7123 , n7031 , n7094 );
and ( n7124 , n821 , n7006 );
and ( n7125 , n7123 , n7124 );
xor ( n7126 , n7123 , n7124 );
xor ( n7127 , n7035 , n7092 );
and ( n7128 , n822 , n7006 );
and ( n7129 , n7127 , n7128 );
xor ( n7130 , n7127 , n7128 );
xor ( n7131 , n7039 , n7090 );
and ( n7132 , n823 , n7006 );
and ( n7133 , n7131 , n7132 );
xor ( n7134 , n7131 , n7132 );
xor ( n7135 , n7043 , n7088 );
and ( n7136 , n824 , n7006 );
and ( n7137 , n7135 , n7136 );
xor ( n7138 , n7135 , n7136 );
xor ( n7139 , n7047 , n7086 );
and ( n7140 , n825 , n7006 );
and ( n7141 , n7139 , n7140 );
xor ( n7142 , n7139 , n7140 );
xor ( n7143 , n7051 , n7084 );
and ( n7144 , n826 , n7006 );
and ( n7145 , n7143 , n7144 );
xor ( n7146 , n7143 , n7144 );
xor ( n7147 , n7055 , n7082 );
and ( n7148 , n827 , n7006 );
and ( n7149 , n7147 , n7148 );
xor ( n7150 , n7147 , n7148 );
xor ( n7151 , n7059 , n7080 );
and ( n7152 , n828 , n7006 );
and ( n7153 , n7151 , n7152 );
xor ( n7154 , n7151 , n7152 );
xor ( n7155 , n7063 , n7078 );
and ( n7156 , n829 , n7006 );
and ( n7157 , n7155 , n7156 );
xor ( n7158 , n7155 , n7156 );
xor ( n7159 , n7067 , n7076 );
and ( n7160 , n830 , n7006 );
and ( n7161 , n7159 , n7160 );
xor ( n7162 , n7159 , n7160 );
xor ( n7163 , n7071 , n7074 );
and ( n7164 , n831 , n7006 );
and ( n7165 , n7163 , n7164 );
and ( n7166 , n7162 , n7165 );
or ( n7167 , n7161 , n7166 );
and ( n7168 , n7158 , n7167 );
or ( n7169 , n7157 , n7168 );
and ( n7170 , n7154 , n7169 );
or ( n7171 , n7153 , n7170 );
and ( n7172 , n7150 , n7171 );
or ( n7173 , n7149 , n7172 );
and ( n7174 , n7146 , n7173 );
or ( n7175 , n7145 , n7174 );
and ( n7176 , n7142 , n7175 );
or ( n7177 , n7141 , n7176 );
and ( n7178 , n7138 , n7177 );
or ( n7179 , n7137 , n7178 );
and ( n7180 , n7134 , n7179 );
or ( n7181 , n7133 , n7180 );
and ( n7182 , n7130 , n7181 );
or ( n7183 , n7129 , n7182 );
and ( n7184 , n7126 , n7183 );
or ( n7185 , n7125 , n7184 );
and ( n7186 , n7122 , n7185 );
or ( n7187 , n7121 , n7186 );
and ( n7188 , n7118 , n7187 );
or ( n7189 , n7117 , n7188 );
and ( n7190 , n7114 , n7189 );
or ( n7191 , n7113 , n7190 );
and ( n7192 , n7110 , n7191 );
or ( n7193 , n7109 , n7192 );
and ( n7194 , n7106 , n7193 );
or ( n7195 , n7105 , n7194 );
and ( n7196 , n816 , n7002 );
and ( n7197 , n7195 , n7196 );
xor ( n7198 , n7195 , n7196 );
xor ( n7199 , n7106 , n7193 );
and ( n7200 , n817 , n7002 );
and ( n7201 , n7199 , n7200 );
xor ( n7202 , n7199 , n7200 );
xor ( n7203 , n7110 , n7191 );
and ( n7204 , n818 , n7002 );
and ( n7205 , n7203 , n7204 );
xor ( n7206 , n7203 , n7204 );
xor ( n7207 , n7114 , n7189 );
and ( n7208 , n819 , n7002 );
and ( n7209 , n7207 , n7208 );
xor ( n7210 , n7207 , n7208 );
xor ( n7211 , n7118 , n7187 );
and ( n7212 , n820 , n7002 );
and ( n7213 , n7211 , n7212 );
xor ( n7214 , n7211 , n7212 );
xor ( n7215 , n7122 , n7185 );
and ( n7216 , n821 , n7002 );
and ( n7217 , n7215 , n7216 );
xor ( n7218 , n7215 , n7216 );
xor ( n7219 , n7126 , n7183 );
and ( n7220 , n822 , n7002 );
and ( n7221 , n7219 , n7220 );
xor ( n7222 , n7219 , n7220 );
xor ( n7223 , n7130 , n7181 );
and ( n7224 , n823 , n7002 );
and ( n7225 , n7223 , n7224 );
xor ( n7226 , n7223 , n7224 );
xor ( n7227 , n7134 , n7179 );
and ( n7228 , n824 , n7002 );
and ( n7229 , n7227 , n7228 );
xor ( n7230 , n7227 , n7228 );
xor ( n7231 , n7138 , n7177 );
and ( n7232 , n825 , n7002 );
and ( n7233 , n7231 , n7232 );
xor ( n7234 , n7231 , n7232 );
xor ( n7235 , n7142 , n7175 );
and ( n7236 , n826 , n7002 );
and ( n7237 , n7235 , n7236 );
xor ( n7238 , n7235 , n7236 );
xor ( n7239 , n7146 , n7173 );
and ( n7240 , n827 , n7002 );
and ( n7241 , n7239 , n7240 );
xor ( n7242 , n7239 , n7240 );
xor ( n7243 , n7150 , n7171 );
and ( n7244 , n828 , n7002 );
and ( n7245 , n7243 , n7244 );
xor ( n7246 , n7243 , n7244 );
xor ( n7247 , n7154 , n7169 );
and ( n7248 , n829 , n7002 );
and ( n7249 , n7247 , n7248 );
xor ( n7250 , n7247 , n7248 );
xor ( n7251 , n7158 , n7167 );
and ( n7252 , n830 , n7002 );
and ( n7253 , n7251 , n7252 );
xor ( n7254 , n7251 , n7252 );
xor ( n7255 , n7162 , n7165 );
and ( n7256 , n831 , n7002 );
and ( n7257 , n7255 , n7256 );
and ( n7258 , n7254 , n7257 );
or ( n7259 , n7253 , n7258 );
and ( n7260 , n7250 , n7259 );
or ( n7261 , n7249 , n7260 );
and ( n7262 , n7246 , n7261 );
or ( n7263 , n7245 , n7262 );
and ( n7264 , n7242 , n7263 );
or ( n7265 , n7241 , n7264 );
and ( n7266 , n7238 , n7265 );
or ( n7267 , n7237 , n7266 );
and ( n7268 , n7234 , n7267 );
or ( n7269 , n7233 , n7268 );
and ( n7270 , n7230 , n7269 );
or ( n7271 , n7229 , n7270 );
and ( n7272 , n7226 , n7271 );
or ( n7273 , n7225 , n7272 );
and ( n7274 , n7222 , n7273 );
or ( n7275 , n7221 , n7274 );
and ( n7276 , n7218 , n7275 );
or ( n7277 , n7217 , n7276 );
and ( n7278 , n7214 , n7277 );
or ( n7279 , n7213 , n7278 );
and ( n7280 , n7210 , n7279 );
or ( n7281 , n7209 , n7280 );
and ( n7282 , n7206 , n7281 );
or ( n7283 , n7205 , n7282 );
and ( n7284 , n7202 , n7283 );
or ( n7285 , n7201 , n7284 );
and ( n7286 , n7198 , n7285 );
or ( n7287 , n7197 , n7286 );
and ( n7288 , n816 , n6998 );
and ( n7289 , n7287 , n7288 );
xor ( n7290 , n7287 , n7288 );
xor ( n7291 , n7198 , n7285 );
and ( n7292 , n817 , n6998 );
and ( n7293 , n7291 , n7292 );
xor ( n7294 , n7291 , n7292 );
xor ( n7295 , n7202 , n7283 );
and ( n7296 , n818 , n6998 );
and ( n7297 , n7295 , n7296 );
xor ( n7298 , n7295 , n7296 );
xor ( n7299 , n7206 , n7281 );
and ( n7300 , n819 , n6998 );
and ( n7301 , n7299 , n7300 );
xor ( n7302 , n7299 , n7300 );
xor ( n7303 , n7210 , n7279 );
and ( n7304 , n820 , n6998 );
and ( n7305 , n7303 , n7304 );
xor ( n7306 , n7303 , n7304 );
xor ( n7307 , n7214 , n7277 );
and ( n7308 , n821 , n6998 );
and ( n7309 , n7307 , n7308 );
xor ( n7310 , n7307 , n7308 );
xor ( n7311 , n7218 , n7275 );
and ( n7312 , n822 , n6998 );
and ( n7313 , n7311 , n7312 );
xor ( n7314 , n7311 , n7312 );
xor ( n7315 , n7222 , n7273 );
and ( n7316 , n823 , n6998 );
and ( n7317 , n7315 , n7316 );
xor ( n7318 , n7315 , n7316 );
xor ( n7319 , n7226 , n7271 );
and ( n7320 , n824 , n6998 );
and ( n7321 , n7319 , n7320 );
xor ( n7322 , n7319 , n7320 );
xor ( n7323 , n7230 , n7269 );
and ( n7324 , n825 , n6998 );
and ( n7325 , n7323 , n7324 );
xor ( n7326 , n7323 , n7324 );
xor ( n7327 , n7234 , n7267 );
and ( n7328 , n826 , n6998 );
and ( n7329 , n7327 , n7328 );
xor ( n7330 , n7327 , n7328 );
xor ( n7331 , n7238 , n7265 );
and ( n7332 , n827 , n6998 );
and ( n7333 , n7331 , n7332 );
xor ( n7334 , n7331 , n7332 );
xor ( n7335 , n7242 , n7263 );
and ( n7336 , n828 , n6998 );
and ( n7337 , n7335 , n7336 );
xor ( n7338 , n7335 , n7336 );
xor ( n7339 , n7246 , n7261 );
and ( n7340 , n829 , n6998 );
and ( n7341 , n7339 , n7340 );
xor ( n7342 , n7339 , n7340 );
xor ( n7343 , n7250 , n7259 );
and ( n7344 , n830 , n6998 );
and ( n7345 , n7343 , n7344 );
xor ( n7346 , n7343 , n7344 );
xor ( n7347 , n7254 , n7257 );
and ( n7348 , n831 , n6998 );
and ( n7349 , n7347 , n7348 );
and ( n7350 , n7346 , n7349 );
or ( n7351 , n7345 , n7350 );
and ( n7352 , n7342 , n7351 );
or ( n7353 , n7341 , n7352 );
and ( n7354 , n7338 , n7353 );
or ( n7355 , n7337 , n7354 );
and ( n7356 , n7334 , n7355 );
or ( n7357 , n7333 , n7356 );
and ( n7358 , n7330 , n7357 );
or ( n7359 , n7329 , n7358 );
and ( n7360 , n7326 , n7359 );
or ( n7361 , n7325 , n7360 );
and ( n7362 , n7322 , n7361 );
or ( n7363 , n7321 , n7362 );
and ( n7364 , n7318 , n7363 );
or ( n7365 , n7317 , n7364 );
and ( n7366 , n7314 , n7365 );
or ( n7367 , n7313 , n7366 );
and ( n7368 , n7310 , n7367 );
or ( n7369 , n7309 , n7368 );
and ( n7370 , n7306 , n7369 );
or ( n7371 , n7305 , n7370 );
and ( n7372 , n7302 , n7371 );
or ( n7373 , n7301 , n7372 );
and ( n7374 , n7298 , n7373 );
or ( n7375 , n7297 , n7374 );
and ( n7376 , n7294 , n7375 );
or ( n7377 , n7293 , n7376 );
and ( n7378 , n7290 , n7377 );
or ( n7379 , n7289 , n7378 );
and ( n7380 , n816 , n6994 );
and ( n7381 , n7379 , n7380 );
xor ( n7382 , n7379 , n7380 );
xor ( n7383 , n7290 , n7377 );
and ( n7384 , n817 , n6994 );
and ( n7385 , n7383 , n7384 );
xor ( n7386 , n7383 , n7384 );
xor ( n7387 , n7294 , n7375 );
and ( n7388 , n818 , n6994 );
and ( n7389 , n7387 , n7388 );
xor ( n7390 , n7387 , n7388 );
xor ( n7391 , n7298 , n7373 );
and ( n7392 , n819 , n6994 );
and ( n7393 , n7391 , n7392 );
xor ( n7394 , n7391 , n7392 );
xor ( n7395 , n7302 , n7371 );
and ( n7396 , n820 , n6994 );
and ( n7397 , n7395 , n7396 );
xor ( n7398 , n7395 , n7396 );
xor ( n7399 , n7306 , n7369 );
and ( n7400 , n821 , n6994 );
and ( n7401 , n7399 , n7400 );
xor ( n7402 , n7399 , n7400 );
xor ( n7403 , n7310 , n7367 );
and ( n7404 , n822 , n6994 );
and ( n7405 , n7403 , n7404 );
xor ( n7406 , n7403 , n7404 );
xor ( n7407 , n7314 , n7365 );
and ( n7408 , n823 , n6994 );
and ( n7409 , n7407 , n7408 );
xor ( n7410 , n7407 , n7408 );
xor ( n7411 , n7318 , n7363 );
and ( n7412 , n824 , n6994 );
and ( n7413 , n7411 , n7412 );
xor ( n7414 , n7411 , n7412 );
xor ( n7415 , n7322 , n7361 );
and ( n7416 , n825 , n6994 );
and ( n7417 , n7415 , n7416 );
xor ( n7418 , n7415 , n7416 );
xor ( n7419 , n7326 , n7359 );
and ( n7420 , n826 , n6994 );
and ( n7421 , n7419 , n7420 );
xor ( n7422 , n7419 , n7420 );
xor ( n7423 , n7330 , n7357 );
and ( n7424 , n827 , n6994 );
and ( n7425 , n7423 , n7424 );
xor ( n7426 , n7423 , n7424 );
xor ( n7427 , n7334 , n7355 );
and ( n7428 , n828 , n6994 );
and ( n7429 , n7427 , n7428 );
xor ( n7430 , n7427 , n7428 );
xor ( n7431 , n7338 , n7353 );
and ( n7432 , n829 , n6994 );
and ( n7433 , n7431 , n7432 );
xor ( n7434 , n7431 , n7432 );
xor ( n7435 , n7342 , n7351 );
and ( n7436 , n830 , n6994 );
and ( n7437 , n7435 , n7436 );
xor ( n7438 , n7435 , n7436 );
xor ( n7439 , n7346 , n7349 );
and ( n7440 , n831 , n6994 );
and ( n7441 , n7439 , n7440 );
and ( n7442 , n7438 , n7441 );
or ( n7443 , n7437 , n7442 );
and ( n7444 , n7434 , n7443 );
or ( n7445 , n7433 , n7444 );
and ( n7446 , n7430 , n7445 );
or ( n7447 , n7429 , n7446 );
and ( n7448 , n7426 , n7447 );
or ( n7449 , n7425 , n7448 );
and ( n7450 , n7422 , n7449 );
or ( n7451 , n7421 , n7450 );
and ( n7452 , n7418 , n7451 );
or ( n7453 , n7417 , n7452 );
and ( n7454 , n7414 , n7453 );
or ( n7455 , n7413 , n7454 );
and ( n7456 , n7410 , n7455 );
or ( n7457 , n7409 , n7456 );
and ( n7458 , n7406 , n7457 );
or ( n7459 , n7405 , n7458 );
and ( n7460 , n7402 , n7459 );
or ( n7461 , n7401 , n7460 );
and ( n7462 , n7398 , n7461 );
or ( n7463 , n7397 , n7462 );
and ( n7464 , n7394 , n7463 );
or ( n7465 , n7393 , n7464 );
and ( n7466 , n7390 , n7465 );
or ( n7467 , n7389 , n7466 );
and ( n7468 , n7386 , n7467 );
or ( n7469 , n7385 , n7468 );
and ( n7470 , n7382 , n7469 );
or ( n7471 , n7381 , n7470 );
and ( n7472 , n816 , n6990 );
and ( n7473 , n7471 , n7472 );
xor ( n7474 , n7471 , n7472 );
xor ( n7475 , n7382 , n7469 );
and ( n7476 , n817 , n6990 );
and ( n7477 , n7475 , n7476 );
xor ( n7478 , n7475 , n7476 );
xor ( n7479 , n7386 , n7467 );
and ( n7480 , n818 , n6990 );
and ( n7481 , n7479 , n7480 );
xor ( n7482 , n7479 , n7480 );
xor ( n7483 , n7390 , n7465 );
and ( n7484 , n819 , n6990 );
and ( n7485 , n7483 , n7484 );
xor ( n7486 , n7483 , n7484 );
xor ( n7487 , n7394 , n7463 );
and ( n7488 , n820 , n6990 );
and ( n7489 , n7487 , n7488 );
xor ( n7490 , n7487 , n7488 );
xor ( n7491 , n7398 , n7461 );
and ( n7492 , n821 , n6990 );
and ( n7493 , n7491 , n7492 );
xor ( n7494 , n7491 , n7492 );
xor ( n7495 , n7402 , n7459 );
and ( n7496 , n822 , n6990 );
and ( n7497 , n7495 , n7496 );
xor ( n7498 , n7495 , n7496 );
xor ( n7499 , n7406 , n7457 );
and ( n7500 , n823 , n6990 );
and ( n7501 , n7499 , n7500 );
xor ( n7502 , n7499 , n7500 );
xor ( n7503 , n7410 , n7455 );
and ( n7504 , n824 , n6990 );
and ( n7505 , n7503 , n7504 );
xor ( n7506 , n7503 , n7504 );
xor ( n7507 , n7414 , n7453 );
and ( n7508 , n825 , n6990 );
and ( n7509 , n7507 , n7508 );
xor ( n7510 , n7507 , n7508 );
xor ( n7511 , n7418 , n7451 );
and ( n7512 , n826 , n6990 );
and ( n7513 , n7511 , n7512 );
xor ( n7514 , n7511 , n7512 );
xor ( n7515 , n7422 , n7449 );
and ( n7516 , n827 , n6990 );
and ( n7517 , n7515 , n7516 );
xor ( n7518 , n7515 , n7516 );
xor ( n7519 , n7426 , n7447 );
and ( n7520 , n828 , n6990 );
and ( n7521 , n7519 , n7520 );
xor ( n7522 , n7519 , n7520 );
xor ( n7523 , n7430 , n7445 );
and ( n7524 , n829 , n6990 );
and ( n7525 , n7523 , n7524 );
xor ( n7526 , n7523 , n7524 );
xor ( n7527 , n7434 , n7443 );
and ( n7528 , n830 , n6990 );
and ( n7529 , n7527 , n7528 );
xor ( n7530 , n7527 , n7528 );
xor ( n7531 , n7438 , n7441 );
and ( n7532 , n831 , n6990 );
and ( n7533 , n7531 , n7532 );
and ( n7534 , n7530 , n7533 );
or ( n7535 , n7529 , n7534 );
and ( n7536 , n7526 , n7535 );
or ( n7537 , n7525 , n7536 );
and ( n7538 , n7522 , n7537 );
or ( n7539 , n7521 , n7538 );
and ( n7540 , n7518 , n7539 );
or ( n7541 , n7517 , n7540 );
and ( n7542 , n7514 , n7541 );
or ( n7543 , n7513 , n7542 );
and ( n7544 , n7510 , n7543 );
or ( n7545 , n7509 , n7544 );
and ( n7546 , n7506 , n7545 );
or ( n7547 , n7505 , n7546 );
and ( n7548 , n7502 , n7547 );
or ( n7549 , n7501 , n7548 );
and ( n7550 , n7498 , n7549 );
or ( n7551 , n7497 , n7550 );
and ( n7552 , n7494 , n7551 );
or ( n7553 , n7493 , n7552 );
and ( n7554 , n7490 , n7553 );
or ( n7555 , n7489 , n7554 );
and ( n7556 , n7486 , n7555 );
or ( n7557 , n7485 , n7556 );
and ( n7558 , n7482 , n7557 );
or ( n7559 , n7481 , n7558 );
and ( n7560 , n7478 , n7559 );
or ( n7561 , n7477 , n7560 );
and ( n7562 , n7474 , n7561 );
or ( n7563 , n7473 , n7562 );
and ( n7564 , n816 , n6986 );
and ( n7565 , n7563 , n7564 );
xor ( n7566 , n7563 , n7564 );
xor ( n7567 , n7474 , n7561 );
and ( n7568 , n817 , n6986 );
and ( n7569 , n7567 , n7568 );
xor ( n7570 , n7567 , n7568 );
xor ( n7571 , n7478 , n7559 );
and ( n7572 , n818 , n6986 );
and ( n7573 , n7571 , n7572 );
xor ( n7574 , n7571 , n7572 );
xor ( n7575 , n7482 , n7557 );
and ( n7576 , n819 , n6986 );
and ( n7577 , n7575 , n7576 );
xor ( n7578 , n7575 , n7576 );
xor ( n7579 , n7486 , n7555 );
and ( n7580 , n820 , n6986 );
and ( n7581 , n7579 , n7580 );
xor ( n7582 , n7579 , n7580 );
xor ( n7583 , n7490 , n7553 );
and ( n7584 , n821 , n6986 );
and ( n7585 , n7583 , n7584 );
xor ( n7586 , n7583 , n7584 );
xor ( n7587 , n7494 , n7551 );
and ( n7588 , n822 , n6986 );
and ( n7589 , n7587 , n7588 );
xor ( n7590 , n7587 , n7588 );
xor ( n7591 , n7498 , n7549 );
and ( n7592 , n823 , n6986 );
and ( n7593 , n7591 , n7592 );
xor ( n7594 , n7591 , n7592 );
xor ( n7595 , n7502 , n7547 );
and ( n7596 , n824 , n6986 );
and ( n7597 , n7595 , n7596 );
xor ( n7598 , n7595 , n7596 );
xor ( n7599 , n7506 , n7545 );
and ( n7600 , n825 , n6986 );
and ( n7601 , n7599 , n7600 );
xor ( n7602 , n7599 , n7600 );
xor ( n7603 , n7510 , n7543 );
and ( n7604 , n826 , n6986 );
and ( n7605 , n7603 , n7604 );
xor ( n7606 , n7603 , n7604 );
xor ( n7607 , n7514 , n7541 );
and ( n7608 , n827 , n6986 );
and ( n7609 , n7607 , n7608 );
xor ( n7610 , n7607 , n7608 );
xor ( n7611 , n7518 , n7539 );
and ( n7612 , n828 , n6986 );
and ( n7613 , n7611 , n7612 );
xor ( n7614 , n7611 , n7612 );
xor ( n7615 , n7522 , n7537 );
and ( n7616 , n829 , n6986 );
and ( n7617 , n7615 , n7616 );
xor ( n7618 , n7615 , n7616 );
xor ( n7619 , n7526 , n7535 );
and ( n7620 , n830 , n6986 );
and ( n7621 , n7619 , n7620 );
xor ( n7622 , n7619 , n7620 );
xor ( n7623 , n7530 , n7533 );
and ( n7624 , n831 , n6986 );
and ( n7625 , n7623 , n7624 );
and ( n7626 , n7622 , n7625 );
or ( n7627 , n7621 , n7626 );
and ( n7628 , n7618 , n7627 );
or ( n7629 , n7617 , n7628 );
and ( n7630 , n7614 , n7629 );
or ( n7631 , n7613 , n7630 );
and ( n7632 , n7610 , n7631 );
or ( n7633 , n7609 , n7632 );
and ( n7634 , n7606 , n7633 );
or ( n7635 , n7605 , n7634 );
and ( n7636 , n7602 , n7635 );
or ( n7637 , n7601 , n7636 );
and ( n7638 , n7598 , n7637 );
or ( n7639 , n7597 , n7638 );
and ( n7640 , n7594 , n7639 );
or ( n7641 , n7593 , n7640 );
and ( n7642 , n7590 , n7641 );
or ( n7643 , n7589 , n7642 );
and ( n7644 , n7586 , n7643 );
or ( n7645 , n7585 , n7644 );
and ( n7646 , n7582 , n7645 );
or ( n7647 , n7581 , n7646 );
and ( n7648 , n7578 , n7647 );
or ( n7649 , n7577 , n7648 );
and ( n7650 , n7574 , n7649 );
or ( n7651 , n7573 , n7650 );
and ( n7652 , n7570 , n7651 );
or ( n7653 , n7569 , n7652 );
and ( n7654 , n7566 , n7653 );
or ( n7655 , n7565 , n7654 );
and ( n7656 , n816 , n6982 );
and ( n7657 , n7655 , n7656 );
xor ( n7658 , n7655 , n7656 );
xor ( n7659 , n7566 , n7653 );
and ( n7660 , n817 , n6982 );
and ( n7661 , n7659 , n7660 );
xor ( n7662 , n7659 , n7660 );
xor ( n7663 , n7570 , n7651 );
and ( n7664 , n818 , n6982 );
and ( n7665 , n7663 , n7664 );
xor ( n7666 , n7663 , n7664 );
xor ( n7667 , n7574 , n7649 );
and ( n7668 , n819 , n6982 );
and ( n7669 , n7667 , n7668 );
xor ( n7670 , n7667 , n7668 );
xor ( n7671 , n7578 , n7647 );
and ( n7672 , n820 , n6982 );
and ( n7673 , n7671 , n7672 );
xor ( n7674 , n7671 , n7672 );
xor ( n7675 , n7582 , n7645 );
and ( n7676 , n821 , n6982 );
and ( n7677 , n7675 , n7676 );
xor ( n7678 , n7675 , n7676 );
xor ( n7679 , n7586 , n7643 );
and ( n7680 , n822 , n6982 );
and ( n7681 , n7679 , n7680 );
xor ( n7682 , n7679 , n7680 );
xor ( n7683 , n7590 , n7641 );
and ( n7684 , n823 , n6982 );
and ( n7685 , n7683 , n7684 );
xor ( n7686 , n7683 , n7684 );
xor ( n7687 , n7594 , n7639 );
and ( n7688 , n824 , n6982 );
and ( n7689 , n7687 , n7688 );
xor ( n7690 , n7687 , n7688 );
xor ( n7691 , n7598 , n7637 );
and ( n7692 , n825 , n6982 );
and ( n7693 , n7691 , n7692 );
xor ( n7694 , n7691 , n7692 );
xor ( n7695 , n7602 , n7635 );
and ( n7696 , n826 , n6982 );
and ( n7697 , n7695 , n7696 );
xor ( n7698 , n7695 , n7696 );
xor ( n7699 , n7606 , n7633 );
and ( n7700 , n827 , n6982 );
and ( n7701 , n7699 , n7700 );
xor ( n7702 , n7699 , n7700 );
xor ( n7703 , n7610 , n7631 );
and ( n7704 , n828 , n6982 );
and ( n7705 , n7703 , n7704 );
xor ( n7706 , n7703 , n7704 );
xor ( n7707 , n7614 , n7629 );
and ( n7708 , n829 , n6982 );
and ( n7709 , n7707 , n7708 );
xor ( n7710 , n7707 , n7708 );
xor ( n7711 , n7618 , n7627 );
and ( n7712 , n830 , n6982 );
and ( n7713 , n7711 , n7712 );
xor ( n7714 , n7711 , n7712 );
xor ( n7715 , n7622 , n7625 );
and ( n7716 , n831 , n6982 );
and ( n7717 , n7715 , n7716 );
and ( n7718 , n7714 , n7717 );
or ( n7719 , n7713 , n7718 );
and ( n7720 , n7710 , n7719 );
or ( n7721 , n7709 , n7720 );
and ( n7722 , n7706 , n7721 );
or ( n7723 , n7705 , n7722 );
and ( n7724 , n7702 , n7723 );
or ( n7725 , n7701 , n7724 );
and ( n7726 , n7698 , n7725 );
or ( n7727 , n7697 , n7726 );
and ( n7728 , n7694 , n7727 );
or ( n7729 , n7693 , n7728 );
and ( n7730 , n7690 , n7729 );
or ( n7731 , n7689 , n7730 );
and ( n7732 , n7686 , n7731 );
or ( n7733 , n7685 , n7732 );
and ( n7734 , n7682 , n7733 );
or ( n7735 , n7681 , n7734 );
and ( n7736 , n7678 , n7735 );
or ( n7737 , n7677 , n7736 );
and ( n7738 , n7674 , n7737 );
or ( n7739 , n7673 , n7738 );
and ( n7740 , n7670 , n7739 );
or ( n7741 , n7669 , n7740 );
and ( n7742 , n7666 , n7741 );
or ( n7743 , n7665 , n7742 );
and ( n7744 , n7662 , n7743 );
or ( n7745 , n7661 , n7744 );
and ( n7746 , n7658 , n7745 );
or ( n7747 , n7657 , n7746 );
and ( n7748 , n816 , n6978 );
and ( n7749 , n7747 , n7748 );
xor ( n7750 , n7747 , n7748 );
xor ( n7751 , n7658 , n7745 );
and ( n7752 , n817 , n6978 );
and ( n7753 , n7751 , n7752 );
xor ( n7754 , n7751 , n7752 );
xor ( n7755 , n7662 , n7743 );
and ( n7756 , n818 , n6978 );
and ( n7757 , n7755 , n7756 );
xor ( n7758 , n7755 , n7756 );
xor ( n7759 , n7666 , n7741 );
and ( n7760 , n819 , n6978 );
and ( n7761 , n7759 , n7760 );
xor ( n7762 , n7759 , n7760 );
xor ( n7763 , n7670 , n7739 );
and ( n7764 , n820 , n6978 );
and ( n7765 , n7763 , n7764 );
xor ( n7766 , n7763 , n7764 );
xor ( n7767 , n7674 , n7737 );
and ( n7768 , n821 , n6978 );
and ( n7769 , n7767 , n7768 );
xor ( n7770 , n7767 , n7768 );
xor ( n7771 , n7678 , n7735 );
and ( n7772 , n822 , n6978 );
and ( n7773 , n7771 , n7772 );
xor ( n7774 , n7771 , n7772 );
xor ( n7775 , n7682 , n7733 );
and ( n7776 , n823 , n6978 );
and ( n7777 , n7775 , n7776 );
xor ( n7778 , n7775 , n7776 );
xor ( n7779 , n7686 , n7731 );
and ( n7780 , n824 , n6978 );
and ( n7781 , n7779 , n7780 );
xor ( n7782 , n7779 , n7780 );
xor ( n7783 , n7690 , n7729 );
and ( n7784 , n825 , n6978 );
and ( n7785 , n7783 , n7784 );
xor ( n7786 , n7783 , n7784 );
xor ( n7787 , n7694 , n7727 );
and ( n7788 , n826 , n6978 );
and ( n7789 , n7787 , n7788 );
xor ( n7790 , n7787 , n7788 );
xor ( n7791 , n7698 , n7725 );
and ( n7792 , n827 , n6978 );
and ( n7793 , n7791 , n7792 );
xor ( n7794 , n7791 , n7792 );
xor ( n7795 , n7702 , n7723 );
and ( n7796 , n828 , n6978 );
and ( n7797 , n7795 , n7796 );
xor ( n7798 , n7795 , n7796 );
xor ( n7799 , n7706 , n7721 );
and ( n7800 , n829 , n6978 );
and ( n7801 , n7799 , n7800 );
xor ( n7802 , n7799 , n7800 );
xor ( n7803 , n7710 , n7719 );
and ( n7804 , n830 , n6978 );
and ( n7805 , n7803 , n7804 );
xor ( n7806 , n7803 , n7804 );
xor ( n7807 , n7714 , n7717 );
and ( n7808 , n831 , n6978 );
and ( n7809 , n7807 , n7808 );
and ( n7810 , n7806 , n7809 );
or ( n7811 , n7805 , n7810 );
and ( n7812 , n7802 , n7811 );
or ( n7813 , n7801 , n7812 );
and ( n7814 , n7798 , n7813 );
or ( n7815 , n7797 , n7814 );
and ( n7816 , n7794 , n7815 );
or ( n7817 , n7793 , n7816 );
and ( n7818 , n7790 , n7817 );
or ( n7819 , n7789 , n7818 );
and ( n7820 , n7786 , n7819 );
or ( n7821 , n7785 , n7820 );
and ( n7822 , n7782 , n7821 );
or ( n7823 , n7781 , n7822 );
and ( n7824 , n7778 , n7823 );
or ( n7825 , n7777 , n7824 );
and ( n7826 , n7774 , n7825 );
or ( n7827 , n7773 , n7826 );
and ( n7828 , n7770 , n7827 );
or ( n7829 , n7769 , n7828 );
and ( n7830 , n7766 , n7829 );
or ( n7831 , n7765 , n7830 );
and ( n7832 , n7762 , n7831 );
or ( n7833 , n7761 , n7832 );
and ( n7834 , n7758 , n7833 );
or ( n7835 , n7757 , n7834 );
and ( n7836 , n7754 , n7835 );
or ( n7837 , n7753 , n7836 );
and ( n7838 , n7750 , n7837 );
or ( n7839 , n7749 , n7838 );
and ( n7840 , n816 , n6974 );
and ( n7841 , n7839 , n7840 );
xor ( n7842 , n7839 , n7840 );
xor ( n7843 , n7750 , n7837 );
and ( n7844 , n817 , n6974 );
and ( n7845 , n7843 , n7844 );
xor ( n7846 , n7843 , n7844 );
xor ( n7847 , n7754 , n7835 );
and ( n7848 , n818 , n6974 );
and ( n7849 , n7847 , n7848 );
xor ( n7850 , n7847 , n7848 );
xor ( n7851 , n7758 , n7833 );
and ( n7852 , n819 , n6974 );
and ( n7853 , n7851 , n7852 );
xor ( n7854 , n7851 , n7852 );
xor ( n7855 , n7762 , n7831 );
and ( n7856 , n820 , n6974 );
and ( n7857 , n7855 , n7856 );
xor ( n7858 , n7855 , n7856 );
xor ( n7859 , n7766 , n7829 );
and ( n7860 , n821 , n6974 );
and ( n7861 , n7859 , n7860 );
xor ( n7862 , n7859 , n7860 );
xor ( n7863 , n7770 , n7827 );
and ( n7864 , n822 , n6974 );
and ( n7865 , n7863 , n7864 );
xor ( n7866 , n7863 , n7864 );
xor ( n7867 , n7774 , n7825 );
and ( n7868 , n823 , n6974 );
and ( n7869 , n7867 , n7868 );
xor ( n7870 , n7867 , n7868 );
xor ( n7871 , n7778 , n7823 );
and ( n7872 , n824 , n6974 );
and ( n7873 , n7871 , n7872 );
xor ( n7874 , n7871 , n7872 );
xor ( n7875 , n7782 , n7821 );
and ( n7876 , n825 , n6974 );
and ( n7877 , n7875 , n7876 );
xor ( n7878 , n7875 , n7876 );
xor ( n7879 , n7786 , n7819 );
and ( n7880 , n826 , n6974 );
and ( n7881 , n7879 , n7880 );
xor ( n7882 , n7879 , n7880 );
xor ( n7883 , n7790 , n7817 );
and ( n7884 , n827 , n6974 );
and ( n7885 , n7883 , n7884 );
xor ( n7886 , n7883 , n7884 );
xor ( n7887 , n7794 , n7815 );
and ( n7888 , n828 , n6974 );
and ( n7889 , n7887 , n7888 );
xor ( n7890 , n7887 , n7888 );
xor ( n7891 , n7798 , n7813 );
and ( n7892 , n829 , n6974 );
and ( n7893 , n7891 , n7892 );
xor ( n7894 , n7891 , n7892 );
xor ( n7895 , n7802 , n7811 );
and ( n7896 , n830 , n6974 );
and ( n7897 , n7895 , n7896 );
xor ( n7898 , n7895 , n7896 );
xor ( n7899 , n7806 , n7809 );
and ( n7900 , n831 , n6974 );
and ( n7901 , n7899 , n7900 );
and ( n7902 , n7898 , n7901 );
or ( n7903 , n7897 , n7902 );
and ( n7904 , n7894 , n7903 );
or ( n7905 , n7893 , n7904 );
and ( n7906 , n7890 , n7905 );
or ( n7907 , n7889 , n7906 );
and ( n7908 , n7886 , n7907 );
or ( n7909 , n7885 , n7908 );
and ( n7910 , n7882 , n7909 );
or ( n7911 , n7881 , n7910 );
and ( n7912 , n7878 , n7911 );
or ( n7913 , n7877 , n7912 );
and ( n7914 , n7874 , n7913 );
or ( n7915 , n7873 , n7914 );
and ( n7916 , n7870 , n7915 );
or ( n7917 , n7869 , n7916 );
and ( n7918 , n7866 , n7917 );
or ( n7919 , n7865 , n7918 );
and ( n7920 , n7862 , n7919 );
or ( n7921 , n7861 , n7920 );
and ( n7922 , n7858 , n7921 );
or ( n7923 , n7857 , n7922 );
and ( n7924 , n7854 , n7923 );
or ( n7925 , n7853 , n7924 );
and ( n7926 , n7850 , n7925 );
or ( n7927 , n7849 , n7926 );
and ( n7928 , n7846 , n7927 );
or ( n7929 , n7845 , n7928 );
and ( n7930 , n7842 , n7929 );
or ( n7931 , n7841 , n7930 );
and ( n7932 , n816 , n6970 );
and ( n7933 , n7931 , n7932 );
xor ( n7934 , n7931 , n7932 );
xor ( n7935 , n7842 , n7929 );
and ( n7936 , n817 , n6970 );
and ( n7937 , n7935 , n7936 );
xor ( n7938 , n7935 , n7936 );
xor ( n7939 , n7846 , n7927 );
and ( n7940 , n818 , n6970 );
and ( n7941 , n7939 , n7940 );
xor ( n7942 , n7939 , n7940 );
xor ( n7943 , n7850 , n7925 );
and ( n7944 , n819 , n6970 );
and ( n7945 , n7943 , n7944 );
xor ( n7946 , n7943 , n7944 );
xor ( n7947 , n7854 , n7923 );
and ( n7948 , n820 , n6970 );
and ( n7949 , n7947 , n7948 );
xor ( n7950 , n7947 , n7948 );
xor ( n7951 , n7858 , n7921 );
and ( n7952 , n821 , n6970 );
and ( n7953 , n7951 , n7952 );
xor ( n7954 , n7951 , n7952 );
xor ( n7955 , n7862 , n7919 );
and ( n7956 , n822 , n6970 );
and ( n7957 , n7955 , n7956 );
xor ( n7958 , n7955 , n7956 );
xor ( n7959 , n7866 , n7917 );
and ( n7960 , n823 , n6970 );
and ( n7961 , n7959 , n7960 );
xor ( n7962 , n7959 , n7960 );
xor ( n7963 , n7870 , n7915 );
and ( n7964 , n824 , n6970 );
and ( n7965 , n7963 , n7964 );
xor ( n7966 , n7963 , n7964 );
xor ( n7967 , n7874 , n7913 );
and ( n7968 , n825 , n6970 );
and ( n7969 , n7967 , n7968 );
xor ( n7970 , n7967 , n7968 );
xor ( n7971 , n7878 , n7911 );
and ( n7972 , n826 , n6970 );
and ( n7973 , n7971 , n7972 );
xor ( n7974 , n7971 , n7972 );
xor ( n7975 , n7882 , n7909 );
and ( n7976 , n827 , n6970 );
and ( n7977 , n7975 , n7976 );
xor ( n7978 , n7975 , n7976 );
xor ( n7979 , n7886 , n7907 );
and ( n7980 , n828 , n6970 );
and ( n7981 , n7979 , n7980 );
xor ( n7982 , n7979 , n7980 );
xor ( n7983 , n7890 , n7905 );
and ( n7984 , n829 , n6970 );
and ( n7985 , n7983 , n7984 );
xor ( n7986 , n7983 , n7984 );
xor ( n7987 , n7894 , n7903 );
and ( n7988 , n830 , n6970 );
and ( n7989 , n7987 , n7988 );
xor ( n7990 , n7987 , n7988 );
xor ( n7991 , n7898 , n7901 );
and ( n7992 , n831 , n6970 );
and ( n7993 , n7991 , n7992 );
and ( n7994 , n7990 , n7993 );
or ( n7995 , n7989 , n7994 );
and ( n7996 , n7986 , n7995 );
or ( n7997 , n7985 , n7996 );
and ( n7998 , n7982 , n7997 );
or ( n7999 , n7981 , n7998 );
and ( n8000 , n7978 , n7999 );
or ( n8001 , n7977 , n8000 );
and ( n8002 , n7974 , n8001 );
or ( n8003 , n7973 , n8002 );
and ( n8004 , n7970 , n8003 );
or ( n8005 , n7969 , n8004 );
and ( n8006 , n7966 , n8005 );
or ( n8007 , n7965 , n8006 );
and ( n8008 , n7962 , n8007 );
or ( n8009 , n7961 , n8008 );
and ( n8010 , n7958 , n8009 );
or ( n8011 , n7957 , n8010 );
and ( n8012 , n7954 , n8011 );
or ( n8013 , n7953 , n8012 );
and ( n8014 , n7950 , n8013 );
or ( n8015 , n7949 , n8014 );
and ( n8016 , n7946 , n8015 );
or ( n8017 , n7945 , n8016 );
and ( n8018 , n7942 , n8017 );
or ( n8019 , n7941 , n8018 );
and ( n8020 , n7938 , n8019 );
or ( n8021 , n7937 , n8020 );
and ( n8022 , n7934 , n8021 );
or ( n8023 , n7933 , n8022 );
and ( n8024 , n816 , n6966 );
and ( n8025 , n8023 , n8024 );
xor ( n8026 , n8023 , n8024 );
xor ( n8027 , n7934 , n8021 );
and ( n8028 , n817 , n6966 );
and ( n8029 , n8027 , n8028 );
xor ( n8030 , n8027 , n8028 );
xor ( n8031 , n7938 , n8019 );
and ( n8032 , n818 , n6966 );
and ( n8033 , n8031 , n8032 );
xor ( n8034 , n8031 , n8032 );
xor ( n8035 , n7942 , n8017 );
and ( n8036 , n819 , n6966 );
and ( n8037 , n8035 , n8036 );
xor ( n8038 , n8035 , n8036 );
xor ( n8039 , n7946 , n8015 );
and ( n8040 , n820 , n6966 );
and ( n8041 , n8039 , n8040 );
xor ( n8042 , n8039 , n8040 );
xor ( n8043 , n7950 , n8013 );
and ( n8044 , n821 , n6966 );
and ( n8045 , n8043 , n8044 );
xor ( n8046 , n8043 , n8044 );
xor ( n8047 , n7954 , n8011 );
and ( n8048 , n822 , n6966 );
and ( n8049 , n8047 , n8048 );
xor ( n8050 , n8047 , n8048 );
xor ( n8051 , n7958 , n8009 );
and ( n8052 , n823 , n6966 );
and ( n8053 , n8051 , n8052 );
xor ( n8054 , n8051 , n8052 );
xor ( n8055 , n7962 , n8007 );
and ( n8056 , n824 , n6966 );
and ( n8057 , n8055 , n8056 );
xor ( n8058 , n8055 , n8056 );
xor ( n8059 , n7966 , n8005 );
and ( n8060 , n825 , n6966 );
and ( n8061 , n8059 , n8060 );
xor ( n8062 , n8059 , n8060 );
xor ( n8063 , n7970 , n8003 );
and ( n8064 , n826 , n6966 );
and ( n8065 , n8063 , n8064 );
xor ( n8066 , n8063 , n8064 );
xor ( n8067 , n7974 , n8001 );
and ( n8068 , n827 , n6966 );
and ( n8069 , n8067 , n8068 );
xor ( n8070 , n8067 , n8068 );
xor ( n8071 , n7978 , n7999 );
and ( n8072 , n828 , n6966 );
and ( n8073 , n8071 , n8072 );
xor ( n8074 , n8071 , n8072 );
xor ( n8075 , n7982 , n7997 );
and ( n8076 , n829 , n6966 );
and ( n8077 , n8075 , n8076 );
xor ( n8078 , n8075 , n8076 );
xor ( n8079 , n7986 , n7995 );
and ( n8080 , n830 , n6966 );
and ( n8081 , n8079 , n8080 );
xor ( n8082 , n8079 , n8080 );
xor ( n8083 , n7990 , n7993 );
and ( n8084 , n831 , n6966 );
and ( n8085 , n8083 , n8084 );
and ( n8086 , n8082 , n8085 );
or ( n8087 , n8081 , n8086 );
and ( n8088 , n8078 , n8087 );
or ( n8089 , n8077 , n8088 );
and ( n8090 , n8074 , n8089 );
or ( n8091 , n8073 , n8090 );
and ( n8092 , n8070 , n8091 );
or ( n8093 , n8069 , n8092 );
and ( n8094 , n8066 , n8093 );
or ( n8095 , n8065 , n8094 );
and ( n8096 , n8062 , n8095 );
or ( n8097 , n8061 , n8096 );
and ( n8098 , n8058 , n8097 );
or ( n8099 , n8057 , n8098 );
and ( n8100 , n8054 , n8099 );
or ( n8101 , n8053 , n8100 );
and ( n8102 , n8050 , n8101 );
or ( n8103 , n8049 , n8102 );
and ( n8104 , n8046 , n8103 );
or ( n8105 , n8045 , n8104 );
and ( n8106 , n8042 , n8105 );
or ( n8107 , n8041 , n8106 );
and ( n8108 , n8038 , n8107 );
or ( n8109 , n8037 , n8108 );
and ( n8110 , n8034 , n8109 );
or ( n8111 , n8033 , n8110 );
and ( n8112 , n8030 , n8111 );
or ( n8113 , n8029 , n8112 );
and ( n8114 , n8026 , n8113 );
or ( n8115 , n8025 , n8114 );
and ( n8116 , n816 , n6962 );
and ( n8117 , n8115 , n8116 );
xor ( n8118 , n8115 , n8116 );
xor ( n8119 , n8026 , n8113 );
and ( n8120 , n817 , n6962 );
and ( n8121 , n8119 , n8120 );
xor ( n8122 , n8119 , n8120 );
xor ( n8123 , n8030 , n8111 );
and ( n8124 , n818 , n6962 );
and ( n8125 , n8123 , n8124 );
xor ( n8126 , n8123 , n8124 );
xor ( n8127 , n8034 , n8109 );
and ( n8128 , n819 , n6962 );
and ( n8129 , n8127 , n8128 );
xor ( n8130 , n8127 , n8128 );
xor ( n8131 , n8038 , n8107 );
and ( n8132 , n820 , n6962 );
and ( n8133 , n8131 , n8132 );
xor ( n8134 , n8131 , n8132 );
xor ( n8135 , n8042 , n8105 );
and ( n8136 , n821 , n6962 );
and ( n8137 , n8135 , n8136 );
xor ( n8138 , n8135 , n8136 );
xor ( n8139 , n8046 , n8103 );
and ( n8140 , n822 , n6962 );
and ( n8141 , n8139 , n8140 );
xor ( n8142 , n8139 , n8140 );
xor ( n8143 , n8050 , n8101 );
and ( n8144 , n823 , n6962 );
and ( n8145 , n8143 , n8144 );
xor ( n8146 , n8143 , n8144 );
xor ( n8147 , n8054 , n8099 );
and ( n8148 , n824 , n6962 );
and ( n8149 , n8147 , n8148 );
xor ( n8150 , n8147 , n8148 );
xor ( n8151 , n8058 , n8097 );
and ( n8152 , n825 , n6962 );
and ( n8153 , n8151 , n8152 );
xor ( n8154 , n8151 , n8152 );
xor ( n8155 , n8062 , n8095 );
and ( n8156 , n826 , n6962 );
and ( n8157 , n8155 , n8156 );
xor ( n8158 , n8155 , n8156 );
xor ( n8159 , n8066 , n8093 );
and ( n8160 , n827 , n6962 );
and ( n8161 , n8159 , n8160 );
xor ( n8162 , n8159 , n8160 );
xor ( n8163 , n8070 , n8091 );
and ( n8164 , n828 , n6962 );
and ( n8165 , n8163 , n8164 );
xor ( n8166 , n8163 , n8164 );
xor ( n8167 , n8074 , n8089 );
and ( n8168 , n829 , n6962 );
and ( n8169 , n8167 , n8168 );
xor ( n8170 , n8167 , n8168 );
xor ( n8171 , n8078 , n8087 );
and ( n8172 , n830 , n6962 );
and ( n8173 , n8171 , n8172 );
xor ( n8174 , n8171 , n8172 );
xor ( n8175 , n8082 , n8085 );
and ( n8176 , n831 , n6962 );
and ( n8177 , n8175 , n8176 );
and ( n8178 , n8174 , n8177 );
or ( n8179 , n8173 , n8178 );
and ( n8180 , n8170 , n8179 );
or ( n8181 , n8169 , n8180 );
and ( n8182 , n8166 , n8181 );
or ( n8183 , n8165 , n8182 );
and ( n8184 , n8162 , n8183 );
or ( n8185 , n8161 , n8184 );
and ( n8186 , n8158 , n8185 );
or ( n8187 , n8157 , n8186 );
and ( n8188 , n8154 , n8187 );
or ( n8189 , n8153 , n8188 );
and ( n8190 , n8150 , n8189 );
or ( n8191 , n8149 , n8190 );
and ( n8192 , n8146 , n8191 );
or ( n8193 , n8145 , n8192 );
and ( n8194 , n8142 , n8193 );
or ( n8195 , n8141 , n8194 );
and ( n8196 , n8138 , n8195 );
or ( n8197 , n8137 , n8196 );
and ( n8198 , n8134 , n8197 );
or ( n8199 , n8133 , n8198 );
and ( n8200 , n8130 , n8199 );
or ( n8201 , n8129 , n8200 );
and ( n8202 , n8126 , n8201 );
or ( n8203 , n8125 , n8202 );
and ( n8204 , n8122 , n8203 );
or ( n8205 , n8121 , n8204 );
and ( n8206 , n8118 , n8205 );
or ( n8207 , n8117 , n8206 );
and ( n8208 , n816 , n6958 );
and ( n8209 , n8207 , n8208 );
xor ( n8210 , n8207 , n8208 );
xor ( n8211 , n8118 , n8205 );
and ( n8212 , n817 , n6958 );
and ( n8213 , n8211 , n8212 );
xor ( n8214 , n8211 , n8212 );
xor ( n8215 , n8122 , n8203 );
and ( n8216 , n818 , n6958 );
and ( n8217 , n8215 , n8216 );
xor ( n8218 , n8215 , n8216 );
xor ( n8219 , n8126 , n8201 );
and ( n8220 , n819 , n6958 );
and ( n8221 , n8219 , n8220 );
xor ( n8222 , n8219 , n8220 );
xor ( n8223 , n8130 , n8199 );
and ( n8224 , n820 , n6958 );
and ( n8225 , n8223 , n8224 );
xor ( n8226 , n8223 , n8224 );
xor ( n8227 , n8134 , n8197 );
and ( n8228 , n821 , n6958 );
and ( n8229 , n8227 , n8228 );
xor ( n8230 , n8227 , n8228 );
xor ( n8231 , n8138 , n8195 );
and ( n8232 , n822 , n6958 );
and ( n8233 , n8231 , n8232 );
xor ( n8234 , n8231 , n8232 );
xor ( n8235 , n8142 , n8193 );
and ( n8236 , n823 , n6958 );
and ( n8237 , n8235 , n8236 );
xor ( n8238 , n8235 , n8236 );
xor ( n8239 , n8146 , n8191 );
and ( n8240 , n824 , n6958 );
and ( n8241 , n8239 , n8240 );
xor ( n8242 , n8239 , n8240 );
xor ( n8243 , n8150 , n8189 );
and ( n8244 , n825 , n6958 );
and ( n8245 , n8243 , n8244 );
xor ( n8246 , n8243 , n8244 );
xor ( n8247 , n8154 , n8187 );
and ( n8248 , n826 , n6958 );
and ( n8249 , n8247 , n8248 );
xor ( n8250 , n8247 , n8248 );
xor ( n8251 , n8158 , n8185 );
and ( n8252 , n827 , n6958 );
and ( n8253 , n8251 , n8252 );
xor ( n8254 , n8251 , n8252 );
xor ( n8255 , n8162 , n8183 );
and ( n8256 , n828 , n6958 );
and ( n8257 , n8255 , n8256 );
xor ( n8258 , n8255 , n8256 );
xor ( n8259 , n8166 , n8181 );
and ( n8260 , n829 , n6958 );
and ( n8261 , n8259 , n8260 );
xor ( n8262 , n8259 , n8260 );
xor ( n8263 , n8170 , n8179 );
and ( n8264 , n830 , n6958 );
and ( n8265 , n8263 , n8264 );
xor ( n8266 , n8263 , n8264 );
xor ( n8267 , n8174 , n8177 );
and ( n8268 , n831 , n6958 );
and ( n8269 , n8267 , n8268 );
and ( n8270 , n8266 , n8269 );
or ( n8271 , n8265 , n8270 );
and ( n8272 , n8262 , n8271 );
or ( n8273 , n8261 , n8272 );
and ( n8274 , n8258 , n8273 );
or ( n8275 , n8257 , n8274 );
and ( n8276 , n8254 , n8275 );
or ( n8277 , n8253 , n8276 );
and ( n8278 , n8250 , n8277 );
or ( n8279 , n8249 , n8278 );
and ( n8280 , n8246 , n8279 );
or ( n8281 , n8245 , n8280 );
and ( n8282 , n8242 , n8281 );
or ( n8283 , n8241 , n8282 );
and ( n8284 , n8238 , n8283 );
or ( n8285 , n8237 , n8284 );
and ( n8286 , n8234 , n8285 );
or ( n8287 , n8233 , n8286 );
and ( n8288 , n8230 , n8287 );
or ( n8289 , n8229 , n8288 );
and ( n8290 , n8226 , n8289 );
or ( n8291 , n8225 , n8290 );
and ( n8292 , n8222 , n8291 );
or ( n8293 , n8221 , n8292 );
and ( n8294 , n8218 , n8293 );
or ( n8295 , n8217 , n8294 );
and ( n8296 , n8214 , n8295 );
or ( n8297 , n8213 , n8296 );
and ( n8298 , n8210 , n8297 );
or ( n8299 , n8209 , n8298 );
and ( n8300 , n816 , n6954 );
and ( n8301 , n8299 , n8300 );
xor ( n8302 , n8299 , n8300 );
xor ( n8303 , n8210 , n8297 );
and ( n8304 , n817 , n6954 );
and ( n8305 , n8303 , n8304 );
xor ( n8306 , n8303 , n8304 );
xor ( n8307 , n8214 , n8295 );
and ( n8308 , n818 , n6954 );
and ( n8309 , n8307 , n8308 );
xor ( n8310 , n8307 , n8308 );
xor ( n8311 , n8218 , n8293 );
and ( n8312 , n819 , n6954 );
and ( n8313 , n8311 , n8312 );
xor ( n8314 , n8311 , n8312 );
xor ( n8315 , n8222 , n8291 );
and ( n8316 , n820 , n6954 );
and ( n8317 , n8315 , n8316 );
xor ( n8318 , n8315 , n8316 );
xor ( n8319 , n8226 , n8289 );
and ( n8320 , n821 , n6954 );
and ( n8321 , n8319 , n8320 );
xor ( n8322 , n8319 , n8320 );
xor ( n8323 , n8230 , n8287 );
and ( n8324 , n822 , n6954 );
and ( n8325 , n8323 , n8324 );
xor ( n8326 , n8323 , n8324 );
xor ( n8327 , n8234 , n8285 );
and ( n8328 , n823 , n6954 );
and ( n8329 , n8327 , n8328 );
xor ( n8330 , n8327 , n8328 );
xor ( n8331 , n8238 , n8283 );
and ( n8332 , n824 , n6954 );
and ( n8333 , n8331 , n8332 );
xor ( n8334 , n8331 , n8332 );
xor ( n8335 , n8242 , n8281 );
and ( n8336 , n825 , n6954 );
and ( n8337 , n8335 , n8336 );
xor ( n8338 , n8335 , n8336 );
xor ( n8339 , n8246 , n8279 );
and ( n8340 , n826 , n6954 );
and ( n8341 , n8339 , n8340 );
xor ( n8342 , n8339 , n8340 );
xor ( n8343 , n8250 , n8277 );
and ( n8344 , n827 , n6954 );
and ( n8345 , n8343 , n8344 );
xor ( n8346 , n8343 , n8344 );
xor ( n8347 , n8254 , n8275 );
and ( n8348 , n828 , n6954 );
and ( n8349 , n8347 , n8348 );
xor ( n8350 , n8347 , n8348 );
xor ( n8351 , n8258 , n8273 );
and ( n8352 , n829 , n6954 );
and ( n8353 , n8351 , n8352 );
xor ( n8354 , n8351 , n8352 );
xor ( n8355 , n8262 , n8271 );
and ( n8356 , n830 , n6954 );
and ( n8357 , n8355 , n8356 );
xor ( n8358 , n8355 , n8356 );
xor ( n8359 , n8266 , n8269 );
and ( n8360 , n831 , n6954 );
and ( n8361 , n8359 , n8360 );
and ( n8362 , n8358 , n8361 );
or ( n8363 , n8357 , n8362 );
and ( n8364 , n8354 , n8363 );
or ( n8365 , n8353 , n8364 );
and ( n8366 , n8350 , n8365 );
or ( n8367 , n8349 , n8366 );
and ( n8368 , n8346 , n8367 );
or ( n8369 , n8345 , n8368 );
and ( n8370 , n8342 , n8369 );
or ( n8371 , n8341 , n8370 );
and ( n8372 , n8338 , n8371 );
or ( n8373 , n8337 , n8372 );
and ( n8374 , n8334 , n8373 );
or ( n8375 , n8333 , n8374 );
and ( n8376 , n8330 , n8375 );
or ( n8377 , n8329 , n8376 );
and ( n8378 , n8326 , n8377 );
or ( n8379 , n8325 , n8378 );
and ( n8380 , n8322 , n8379 );
or ( n8381 , n8321 , n8380 );
and ( n8382 , n8318 , n8381 );
or ( n8383 , n8317 , n8382 );
and ( n8384 , n8314 , n8383 );
or ( n8385 , n8313 , n8384 );
and ( n8386 , n8310 , n8385 );
or ( n8387 , n8309 , n8386 );
and ( n8388 , n8306 , n8387 );
or ( n8389 , n8305 , n8388 );
and ( n8390 , n8302 , n8389 );
or ( n8391 , n8301 , n8390 );
and ( n8392 , n816 , n6950 );
and ( n8393 , n8391 , n8392 );
xor ( n8394 , n8391 , n8392 );
xor ( n8395 , n8302 , n8389 );
and ( n8396 , n817 , n6950 );
and ( n8397 , n8395 , n8396 );
xor ( n8398 , n8395 , n8396 );
xor ( n8399 , n8306 , n8387 );
and ( n8400 , n818 , n6950 );
and ( n8401 , n8399 , n8400 );
xor ( n8402 , n8399 , n8400 );
xor ( n8403 , n8310 , n8385 );
and ( n8404 , n819 , n6950 );
and ( n8405 , n8403 , n8404 );
xor ( n8406 , n8403 , n8404 );
xor ( n8407 , n8314 , n8383 );
and ( n8408 , n820 , n6950 );
and ( n8409 , n8407 , n8408 );
xor ( n8410 , n8407 , n8408 );
xor ( n8411 , n8318 , n8381 );
and ( n8412 , n821 , n6950 );
and ( n8413 , n8411 , n8412 );
xor ( n8414 , n8411 , n8412 );
xor ( n8415 , n8322 , n8379 );
and ( n8416 , n822 , n6950 );
and ( n8417 , n8415 , n8416 );
xor ( n8418 , n8415 , n8416 );
xor ( n8419 , n8326 , n8377 );
and ( n8420 , n823 , n6950 );
and ( n8421 , n8419 , n8420 );
xor ( n8422 , n8419 , n8420 );
xor ( n8423 , n8330 , n8375 );
and ( n8424 , n824 , n6950 );
and ( n8425 , n8423 , n8424 );
xor ( n8426 , n8423 , n8424 );
xor ( n8427 , n8334 , n8373 );
and ( n8428 , n825 , n6950 );
and ( n8429 , n8427 , n8428 );
xor ( n8430 , n8427 , n8428 );
xor ( n8431 , n8338 , n8371 );
and ( n8432 , n826 , n6950 );
and ( n8433 , n8431 , n8432 );
xor ( n8434 , n8431 , n8432 );
xor ( n8435 , n8342 , n8369 );
and ( n8436 , n827 , n6950 );
and ( n8437 , n8435 , n8436 );
xor ( n8438 , n8435 , n8436 );
xor ( n8439 , n8346 , n8367 );
and ( n8440 , n828 , n6950 );
and ( n8441 , n8439 , n8440 );
xor ( n8442 , n8439 , n8440 );
xor ( n8443 , n8350 , n8365 );
and ( n8444 , n829 , n6950 );
and ( n8445 , n8443 , n8444 );
xor ( n8446 , n8443 , n8444 );
xor ( n8447 , n8354 , n8363 );
and ( n8448 , n830 , n6950 );
and ( n8449 , n8447 , n8448 );
xor ( n8450 , n8447 , n8448 );
xor ( n8451 , n8358 , n8361 );
and ( n8452 , n831 , n6950 );
and ( n8453 , n8451 , n8452 );
and ( n8454 , n8450 , n8453 );
or ( n8455 , n8449 , n8454 );
and ( n8456 , n8446 , n8455 );
or ( n8457 , n8445 , n8456 );
and ( n8458 , n8442 , n8457 );
or ( n8459 , n8441 , n8458 );
and ( n8460 , n8438 , n8459 );
or ( n8461 , n8437 , n8460 );
and ( n8462 , n8434 , n8461 );
or ( n8463 , n8433 , n8462 );
and ( n8464 , n8430 , n8463 );
or ( n8465 , n8429 , n8464 );
and ( n8466 , n8426 , n8465 );
or ( n8467 , n8425 , n8466 );
and ( n8468 , n8422 , n8467 );
or ( n8469 , n8421 , n8468 );
and ( n8470 , n8418 , n8469 );
or ( n8471 , n8417 , n8470 );
and ( n8472 , n8414 , n8471 );
or ( n8473 , n8413 , n8472 );
and ( n8474 , n8410 , n8473 );
or ( n8475 , n8409 , n8474 );
and ( n8476 , n8406 , n8475 );
or ( n8477 , n8405 , n8476 );
and ( n8478 , n8402 , n8477 );
or ( n8479 , n8401 , n8478 );
and ( n8480 , n8398 , n8479 );
or ( n8481 , n8397 , n8480 );
and ( n8482 , n8394 , n8481 );
or ( n8483 , n8393 , n8482 );
and ( n8484 , n816 , n6947 );
and ( n8485 , n8483 , n8484 );
xor ( n8486 , n8483 , n8484 );
xor ( n8487 , n8394 , n8481 );
and ( n8488 , n817 , n6947 );
and ( n8489 , n8487 , n8488 );
xor ( n8490 , n8487 , n8488 );
xor ( n8491 , n8398 , n8479 );
and ( n8492 , n818 , n6947 );
and ( n8493 , n8491 , n8492 );
xor ( n8494 , n8491 , n8492 );
xor ( n8495 , n8402 , n8477 );
and ( n8496 , n819 , n6947 );
and ( n8497 , n8495 , n8496 );
xor ( n8498 , n8495 , n8496 );
xor ( n8499 , n8406 , n8475 );
and ( n8500 , n820 , n6947 );
and ( n8501 , n8499 , n8500 );
xor ( n8502 , n8499 , n8500 );
xor ( n8503 , n8410 , n8473 );
and ( n8504 , n821 , n6947 );
and ( n8505 , n8503 , n8504 );
xor ( n8506 , n8503 , n8504 );
xor ( n8507 , n8414 , n8471 );
and ( n8508 , n822 , n6947 );
and ( n8509 , n8507 , n8508 );
xor ( n8510 , n8507 , n8508 );
xor ( n8511 , n8418 , n8469 );
and ( n8512 , n823 , n6947 );
and ( n8513 , n8511 , n8512 );
xor ( n8514 , n8511 , n8512 );
xor ( n8515 , n8422 , n8467 );
and ( n8516 , n824 , n6947 );
and ( n8517 , n8515 , n8516 );
xor ( n8518 , n8515 , n8516 );
xor ( n8519 , n8426 , n8465 );
and ( n8520 , n825 , n6947 );
and ( n8521 , n8519 , n8520 );
xor ( n8522 , n8519 , n8520 );
xor ( n8523 , n8430 , n8463 );
and ( n8524 , n826 , n6947 );
and ( n8525 , n8523 , n8524 );
xor ( n8526 , n8523 , n8524 );
xor ( n8527 , n8434 , n8461 );
and ( n8528 , n827 , n6947 );
and ( n8529 , n8527 , n8528 );
xor ( n8530 , n8527 , n8528 );
xor ( n8531 , n8438 , n8459 );
and ( n8532 , n828 , n6947 );
and ( n8533 , n8531 , n8532 );
xor ( n8534 , n8531 , n8532 );
xor ( n8535 , n8442 , n8457 );
and ( n8536 , n829 , n6947 );
and ( n8537 , n8535 , n8536 );
xor ( n8538 , n8535 , n8536 );
xor ( n8539 , n8446 , n8455 );
and ( n8540 , n830 , n6947 );
and ( n8541 , n8539 , n8540 );
xor ( n8542 , n8539 , n8540 );
xor ( n8543 , n8450 , n8453 );
and ( n8544 , n831 , n6947 );
and ( n8545 , n8543 , n8544 );
and ( n8546 , n8542 , n8545 );
or ( n8547 , n8541 , n8546 );
and ( n8548 , n8538 , n8547 );
or ( n8549 , n8537 , n8548 );
and ( n8550 , n8534 , n8549 );
or ( n8551 , n8533 , n8550 );
and ( n8552 , n8530 , n8551 );
or ( n8553 , n8529 , n8552 );
and ( n8554 , n8526 , n8553 );
or ( n8555 , n8525 , n8554 );
and ( n8556 , n8522 , n8555 );
or ( n8557 , n8521 , n8556 );
and ( n8558 , n8518 , n8557 );
or ( n8559 , n8517 , n8558 );
and ( n8560 , n8514 , n8559 );
or ( n8561 , n8513 , n8560 );
and ( n8562 , n8510 , n8561 );
or ( n8563 , n8509 , n8562 );
and ( n8564 , n8506 , n8563 );
or ( n8565 , n8505 , n8564 );
and ( n8566 , n8502 , n8565 );
or ( n8567 , n8501 , n8566 );
and ( n8568 , n8498 , n8567 );
or ( n8569 , n8497 , n8568 );
and ( n8570 , n8494 , n8569 );
or ( n8571 , n8493 , n8570 );
and ( n8572 , n8490 , n8571 );
or ( n8573 , n8489 , n8572 );
and ( n8574 , n8486 , n8573 );
or ( n8575 , n8485 , n8574 );
and ( n8576 , n816 , n6944 );
and ( n8577 , n8575 , n8576 );
xor ( n8578 , n8575 , n8576 );
xor ( n8579 , n8486 , n8573 );
and ( n8580 , n817 , n6944 );
and ( n8581 , n8579 , n8580 );
xor ( n8582 , n8579 , n8580 );
xor ( n8583 , n8490 , n8571 );
and ( n8584 , n818 , n6944 );
and ( n8585 , n8583 , n8584 );
xor ( n8586 , n8583 , n8584 );
xor ( n8587 , n8494 , n8569 );
and ( n8588 , n819 , n6944 );
and ( n8589 , n8587 , n8588 );
xor ( n8590 , n8587 , n8588 );
xor ( n8591 , n8498 , n8567 );
and ( n8592 , n820 , n6944 );
and ( n8593 , n8591 , n8592 );
xor ( n8594 , n8591 , n8592 );
xor ( n8595 , n8502 , n8565 );
and ( n8596 , n821 , n6944 );
and ( n8597 , n8595 , n8596 );
xor ( n8598 , n8595 , n8596 );
xor ( n8599 , n8506 , n8563 );
and ( n8600 , n822 , n6944 );
and ( n8601 , n8599 , n8600 );
xor ( n8602 , n8599 , n8600 );
xor ( n8603 , n8510 , n8561 );
and ( n8604 , n823 , n6944 );
and ( n8605 , n8603 , n8604 );
xor ( n8606 , n8603 , n8604 );
xor ( n8607 , n8514 , n8559 );
and ( n8608 , n824 , n6944 );
and ( n8609 , n8607 , n8608 );
xor ( n8610 , n8607 , n8608 );
xor ( n8611 , n8518 , n8557 );
and ( n8612 , n825 , n6944 );
and ( n8613 , n8611 , n8612 );
xor ( n8614 , n8611 , n8612 );
xor ( n8615 , n8522 , n8555 );
and ( n8616 , n826 , n6944 );
and ( n8617 , n8615 , n8616 );
xor ( n8618 , n8615 , n8616 );
xor ( n8619 , n8526 , n8553 );
and ( n8620 , n827 , n6944 );
and ( n8621 , n8619 , n8620 );
xor ( n8622 , n8619 , n8620 );
xor ( n8623 , n8530 , n8551 );
and ( n8624 , n828 , n6944 );
and ( n8625 , n8623 , n8624 );
xor ( n8626 , n8623 , n8624 );
xor ( n8627 , n8534 , n8549 );
and ( n8628 , n829 , n6944 );
and ( n8629 , n8627 , n8628 );
xor ( n8630 , n8627 , n8628 );
xor ( n8631 , n8538 , n8547 );
and ( n8632 , n830 , n6944 );
and ( n8633 , n8631 , n8632 );
xor ( n8634 , n8631 , n8632 );
xor ( n8635 , n8542 , n8545 );
and ( n8636 , n831 , n6944 );
and ( n8637 , n8635 , n8636 );
and ( n8638 , n8634 , n8637 );
or ( n8639 , n8633 , n8638 );
and ( n8640 , n8630 , n8639 );
or ( n8641 , n8629 , n8640 );
and ( n8642 , n8626 , n8641 );
or ( n8643 , n8625 , n8642 );
and ( n8644 , n8622 , n8643 );
or ( n8645 , n8621 , n8644 );
and ( n8646 , n8618 , n8645 );
or ( n8647 , n8617 , n8646 );
and ( n8648 , n8614 , n8647 );
or ( n8649 , n8613 , n8648 );
and ( n8650 , n8610 , n8649 );
or ( n8651 , n8609 , n8650 );
and ( n8652 , n8606 , n8651 );
or ( n8653 , n8605 , n8652 );
and ( n8654 , n8602 , n8653 );
or ( n8655 , n8601 , n8654 );
and ( n8656 , n8598 , n8655 );
or ( n8657 , n8597 , n8656 );
and ( n8658 , n8594 , n8657 );
or ( n8659 , n8593 , n8658 );
and ( n8660 , n8590 , n8659 );
or ( n8661 , n8589 , n8660 );
and ( n8662 , n8586 , n8661 );
or ( n8663 , n8585 , n8662 );
and ( n8664 , n8582 , n8663 );
or ( n8665 , n8581 , n8664 );
and ( n8666 , n8578 , n8665 );
or ( n8667 , n8577 , n8666 );
and ( n8668 , n816 , n6941 );
and ( n8669 , n8667 , n8668 );
xor ( n8670 , n8667 , n8668 );
xor ( n8671 , n8578 , n8665 );
and ( n8672 , n817 , n6941 );
and ( n8673 , n8671 , n8672 );
xor ( n8674 , n8671 , n8672 );
xor ( n8675 , n8582 , n8663 );
and ( n8676 , n818 , n6941 );
and ( n8677 , n8675 , n8676 );
xor ( n8678 , n8675 , n8676 );
xor ( n8679 , n8586 , n8661 );
and ( n8680 , n819 , n6941 );
and ( n8681 , n8679 , n8680 );
xor ( n8682 , n8679 , n8680 );
xor ( n8683 , n8590 , n8659 );
and ( n8684 , n820 , n6941 );
and ( n8685 , n8683 , n8684 );
xor ( n8686 , n8683 , n8684 );
xor ( n8687 , n8594 , n8657 );
and ( n8688 , n821 , n6941 );
and ( n8689 , n8687 , n8688 );
xor ( n8690 , n8687 , n8688 );
xor ( n8691 , n8598 , n8655 );
and ( n8692 , n822 , n6941 );
and ( n8693 , n8691 , n8692 );
xor ( n8694 , n8691 , n8692 );
xor ( n8695 , n8602 , n8653 );
and ( n8696 , n823 , n6941 );
and ( n8697 , n8695 , n8696 );
xor ( n8698 , n8695 , n8696 );
xor ( n8699 , n8606 , n8651 );
and ( n8700 , n824 , n6941 );
and ( n8701 , n8699 , n8700 );
xor ( n8702 , n8699 , n8700 );
xor ( n8703 , n8610 , n8649 );
and ( n8704 , n825 , n6941 );
and ( n8705 , n8703 , n8704 );
xor ( n8706 , n8703 , n8704 );
xor ( n8707 , n8614 , n8647 );
and ( n8708 , n826 , n6941 );
and ( n8709 , n8707 , n8708 );
xor ( n8710 , n8707 , n8708 );
xor ( n8711 , n8618 , n8645 );
and ( n8712 , n827 , n6941 );
and ( n8713 , n8711 , n8712 );
xor ( n8714 , n8711 , n8712 );
xor ( n8715 , n8622 , n8643 );
and ( n8716 , n828 , n6941 );
and ( n8717 , n8715 , n8716 );
xor ( n8718 , n8715 , n8716 );
xor ( n8719 , n8626 , n8641 );
and ( n8720 , n829 , n6941 );
and ( n8721 , n8719 , n8720 );
xor ( n8722 , n8719 , n8720 );
xor ( n8723 , n8630 , n8639 );
and ( n8724 , n830 , n6941 );
and ( n8725 , n8723 , n8724 );
xor ( n8726 , n8723 , n8724 );
xor ( n8727 , n8634 , n8637 );
and ( n8728 , n831 , n6941 );
and ( n8729 , n8727 , n8728 );
and ( n8730 , n8726 , n8729 );
or ( n8731 , n8725 , n8730 );
and ( n8732 , n8722 , n8731 );
or ( n8733 , n8721 , n8732 );
and ( n8734 , n8718 , n8733 );
or ( n8735 , n8717 , n8734 );
and ( n8736 , n8714 , n8735 );
or ( n8737 , n8713 , n8736 );
and ( n8738 , n8710 , n8737 );
or ( n8739 , n8709 , n8738 );
and ( n8740 , n8706 , n8739 );
or ( n8741 , n8705 , n8740 );
and ( n8742 , n8702 , n8741 );
or ( n8743 , n8701 , n8742 );
and ( n8744 , n8698 , n8743 );
or ( n8745 , n8697 , n8744 );
and ( n8746 , n8694 , n8745 );
or ( n8747 , n8693 , n8746 );
and ( n8748 , n8690 , n8747 );
or ( n8749 , n8689 , n8748 );
and ( n8750 , n8686 , n8749 );
or ( n8751 , n8685 , n8750 );
and ( n8752 , n8682 , n8751 );
or ( n8753 , n8681 , n8752 );
and ( n8754 , n8678 , n8753 );
or ( n8755 , n8677 , n8754 );
and ( n8756 , n8674 , n8755 );
or ( n8757 , n8673 , n8756 );
and ( n8758 , n8670 , n8757 );
or ( n8759 , n8669 , n8758 );
and ( n8760 , n816 , n6938 );
and ( n8761 , n8759 , n8760 );
xor ( n8762 , n8759 , n8760 );
xor ( n8763 , n8670 , n8757 );
and ( n8764 , n817 , n6938 );
and ( n8765 , n8763 , n8764 );
xor ( n8766 , n8763 , n8764 );
xor ( n8767 , n8674 , n8755 );
and ( n8768 , n818 , n6938 );
and ( n8769 , n8767 , n8768 );
xor ( n8770 , n8767 , n8768 );
xor ( n8771 , n8678 , n8753 );
and ( n8772 , n819 , n6938 );
and ( n8773 , n8771 , n8772 );
xor ( n8774 , n8771 , n8772 );
xor ( n8775 , n8682 , n8751 );
and ( n8776 , n820 , n6938 );
and ( n8777 , n8775 , n8776 );
xor ( n8778 , n8775 , n8776 );
xor ( n8779 , n8686 , n8749 );
and ( n8780 , n821 , n6938 );
and ( n8781 , n8779 , n8780 );
xor ( n8782 , n8779 , n8780 );
xor ( n8783 , n8690 , n8747 );
and ( n8784 , n822 , n6938 );
and ( n8785 , n8783 , n8784 );
xor ( n8786 , n8783 , n8784 );
xor ( n8787 , n8694 , n8745 );
and ( n8788 , n823 , n6938 );
and ( n8789 , n8787 , n8788 );
xor ( n8790 , n8787 , n8788 );
xor ( n8791 , n8698 , n8743 );
and ( n8792 , n824 , n6938 );
and ( n8793 , n8791 , n8792 );
xor ( n8794 , n8791 , n8792 );
xor ( n8795 , n8702 , n8741 );
and ( n8796 , n825 , n6938 );
and ( n8797 , n8795 , n8796 );
xor ( n8798 , n8795 , n8796 );
xor ( n8799 , n8706 , n8739 );
and ( n8800 , n826 , n6938 );
and ( n8801 , n8799 , n8800 );
xor ( n8802 , n8799 , n8800 );
xor ( n8803 , n8710 , n8737 );
and ( n8804 , n827 , n6938 );
and ( n8805 , n8803 , n8804 );
xor ( n8806 , n8803 , n8804 );
xor ( n8807 , n8714 , n8735 );
and ( n8808 , n828 , n6938 );
and ( n8809 , n8807 , n8808 );
xor ( n8810 , n8807 , n8808 );
xor ( n8811 , n8718 , n8733 );
and ( n8812 , n829 , n6938 );
and ( n8813 , n8811 , n8812 );
xor ( n8814 , n8811 , n8812 );
xor ( n8815 , n8722 , n8731 );
and ( n8816 , n830 , n6938 );
and ( n8817 , n8815 , n8816 );
xor ( n8818 , n8815 , n8816 );
xor ( n8819 , n8726 , n8729 );
and ( n8820 , n831 , n6938 );
and ( n8821 , n8819 , n8820 );
and ( n8822 , n8818 , n8821 );
or ( n8823 , n8817 , n8822 );
and ( n8824 , n8814 , n8823 );
or ( n8825 , n8813 , n8824 );
and ( n8826 , n8810 , n8825 );
or ( n8827 , n8809 , n8826 );
and ( n8828 , n8806 , n8827 );
or ( n8829 , n8805 , n8828 );
and ( n8830 , n8802 , n8829 );
or ( n8831 , n8801 , n8830 );
and ( n8832 , n8798 , n8831 );
or ( n8833 , n8797 , n8832 );
and ( n8834 , n8794 , n8833 );
or ( n8835 , n8793 , n8834 );
and ( n8836 , n8790 , n8835 );
or ( n8837 , n8789 , n8836 );
and ( n8838 , n8786 , n8837 );
or ( n8839 , n8785 , n8838 );
and ( n8840 , n8782 , n8839 );
or ( n8841 , n8781 , n8840 );
and ( n8842 , n8778 , n8841 );
or ( n8843 , n8777 , n8842 );
and ( n8844 , n8774 , n8843 );
or ( n8845 , n8773 , n8844 );
and ( n8846 , n8770 , n8845 );
or ( n8847 , n8769 , n8846 );
and ( n8848 , n8766 , n8847 );
or ( n8849 , n8765 , n8848 );
and ( n8850 , n8762 , n8849 );
or ( n8851 , n8761 , n8850 );
and ( n8852 , n816 , n6935 );
and ( n8853 , n8851 , n8852 );
xor ( n8854 , n8851 , n8852 );
xor ( n8855 , n8762 , n8849 );
and ( n8856 , n817 , n6935 );
and ( n8857 , n8855 , n8856 );
xor ( n8858 , n8855 , n8856 );
xor ( n8859 , n8766 , n8847 );
and ( n8860 , n818 , n6935 );
and ( n8861 , n8859 , n8860 );
xor ( n8862 , n8859 , n8860 );
xor ( n8863 , n8770 , n8845 );
and ( n8864 , n819 , n6935 );
and ( n8865 , n8863 , n8864 );
xor ( n8866 , n8863 , n8864 );
xor ( n8867 , n8774 , n8843 );
and ( n8868 , n820 , n6935 );
and ( n8869 , n8867 , n8868 );
xor ( n8870 , n8867 , n8868 );
xor ( n8871 , n8778 , n8841 );
and ( n8872 , n821 , n6935 );
and ( n8873 , n8871 , n8872 );
xor ( n8874 , n8871 , n8872 );
xor ( n8875 , n8782 , n8839 );
and ( n8876 , n822 , n6935 );
and ( n8877 , n8875 , n8876 );
xor ( n8878 , n8875 , n8876 );
xor ( n8879 , n8786 , n8837 );
and ( n8880 , n823 , n6935 );
and ( n8881 , n8879 , n8880 );
xor ( n8882 , n8879 , n8880 );
xor ( n8883 , n8790 , n8835 );
and ( n8884 , n824 , n6935 );
and ( n8885 , n8883 , n8884 );
xor ( n8886 , n8883 , n8884 );
xor ( n8887 , n8794 , n8833 );
and ( n8888 , n825 , n6935 );
and ( n8889 , n8887 , n8888 );
xor ( n8890 , n8887 , n8888 );
xor ( n8891 , n8798 , n8831 );
and ( n8892 , n826 , n6935 );
and ( n8893 , n8891 , n8892 );
xor ( n8894 , n8891 , n8892 );
xor ( n8895 , n8802 , n8829 );
and ( n8896 , n827 , n6935 );
and ( n8897 , n8895 , n8896 );
xor ( n8898 , n8895 , n8896 );
xor ( n8899 , n8806 , n8827 );
and ( n8900 , n828 , n6935 );
and ( n8901 , n8899 , n8900 );
xor ( n8902 , n8899 , n8900 );
xor ( n8903 , n8810 , n8825 );
and ( n8904 , n829 , n6935 );
and ( n8905 , n8903 , n8904 );
xor ( n8906 , n8903 , n8904 );
xor ( n8907 , n8814 , n8823 );
and ( n8908 , n830 , n6935 );
and ( n8909 , n8907 , n8908 );
xor ( n8910 , n8907 , n8908 );
xor ( n8911 , n8818 , n8821 );
and ( n8912 , n831 , n6935 );
and ( n8913 , n8911 , n8912 );
and ( n8914 , n8910 , n8913 );
or ( n8915 , n8909 , n8914 );
and ( n8916 , n8906 , n8915 );
or ( n8917 , n8905 , n8916 );
and ( n8918 , n8902 , n8917 );
or ( n8919 , n8901 , n8918 );
and ( n8920 , n8898 , n8919 );
or ( n8921 , n8897 , n8920 );
and ( n8922 , n8894 , n8921 );
or ( n8923 , n8893 , n8922 );
and ( n8924 , n8890 , n8923 );
or ( n8925 , n8889 , n8924 );
and ( n8926 , n8886 , n8925 );
or ( n8927 , n8885 , n8926 );
and ( n8928 , n8882 , n8927 );
or ( n8929 , n8881 , n8928 );
and ( n8930 , n8878 , n8929 );
or ( n8931 , n8877 , n8930 );
and ( n8932 , n8874 , n8931 );
or ( n8933 , n8873 , n8932 );
and ( n8934 , n8870 , n8933 );
or ( n8935 , n8869 , n8934 );
and ( n8936 , n8866 , n8935 );
or ( n8937 , n8865 , n8936 );
and ( n8938 , n8862 , n8937 );
or ( n8939 , n8861 , n8938 );
and ( n8940 , n8858 , n8939 );
or ( n8941 , n8857 , n8940 );
and ( n8942 , n8854 , n8941 );
or ( n8943 , n8853 , n8942 );
and ( n8944 , n816 , n6932 );
and ( n8945 , n8943 , n8944 );
xor ( n8946 , n8943 , n8944 );
xor ( n8947 , n8854 , n8941 );
and ( n8948 , n817 , n6932 );
and ( n8949 , n8947 , n8948 );
xor ( n8950 , n8947 , n8948 );
xor ( n8951 , n8858 , n8939 );
and ( n8952 , n818 , n6932 );
and ( n8953 , n8951 , n8952 );
xor ( n8954 , n8951 , n8952 );
xor ( n8955 , n8862 , n8937 );
and ( n8956 , n819 , n6932 );
and ( n8957 , n8955 , n8956 );
xor ( n8958 , n8955 , n8956 );
xor ( n8959 , n8866 , n8935 );
and ( n8960 , n820 , n6932 );
and ( n8961 , n8959 , n8960 );
xor ( n8962 , n8959 , n8960 );
xor ( n8963 , n8870 , n8933 );
and ( n8964 , n821 , n6932 );
and ( n8965 , n8963 , n8964 );
xor ( n8966 , n8963 , n8964 );
xor ( n8967 , n8874 , n8931 );
and ( n8968 , n822 , n6932 );
and ( n8969 , n8967 , n8968 );
xor ( n8970 , n8967 , n8968 );
xor ( n8971 , n8878 , n8929 );
and ( n8972 , n823 , n6932 );
and ( n8973 , n8971 , n8972 );
xor ( n8974 , n8971 , n8972 );
xor ( n8975 , n8882 , n8927 );
and ( n8976 , n824 , n6932 );
and ( n8977 , n8975 , n8976 );
xor ( n8978 , n8975 , n8976 );
xor ( n8979 , n8886 , n8925 );
and ( n8980 , n825 , n6932 );
and ( n8981 , n8979 , n8980 );
xor ( n8982 , n8979 , n8980 );
xor ( n8983 , n8890 , n8923 );
and ( n8984 , n826 , n6932 );
and ( n8985 , n8983 , n8984 );
xor ( n8986 , n8983 , n8984 );
xor ( n8987 , n8894 , n8921 );
and ( n8988 , n827 , n6932 );
and ( n8989 , n8987 , n8988 );
xor ( n8990 , n8987 , n8988 );
xor ( n8991 , n8898 , n8919 );
and ( n8992 , n828 , n6932 );
and ( n8993 , n8991 , n8992 );
xor ( n8994 , n8991 , n8992 );
xor ( n8995 , n8902 , n8917 );
and ( n8996 , n829 , n6932 );
and ( n8997 , n8995 , n8996 );
xor ( n8998 , n8995 , n8996 );
xor ( n8999 , n8906 , n8915 );
and ( n9000 , n830 , n6932 );
and ( n9001 , n8999 , n9000 );
xor ( n9002 , n8999 , n9000 );
xor ( n9003 , n8910 , n8913 );
and ( n9004 , n831 , n6932 );
and ( n9005 , n9003 , n9004 );
and ( n9006 , n9002 , n9005 );
or ( n9007 , n9001 , n9006 );
and ( n9008 , n8998 , n9007 );
or ( n9009 , n8997 , n9008 );
and ( n9010 , n8994 , n9009 );
or ( n9011 , n8993 , n9010 );
and ( n9012 , n8990 , n9011 );
or ( n9013 , n8989 , n9012 );
and ( n9014 , n8986 , n9013 );
or ( n9015 , n8985 , n9014 );
and ( n9016 , n8982 , n9015 );
or ( n9017 , n8981 , n9016 );
and ( n9018 , n8978 , n9017 );
or ( n9019 , n8977 , n9018 );
and ( n9020 , n8974 , n9019 );
or ( n9021 , n8973 , n9020 );
and ( n9022 , n8970 , n9021 );
or ( n9023 , n8969 , n9022 );
and ( n9024 , n8966 , n9023 );
or ( n9025 , n8965 , n9024 );
and ( n9026 , n8962 , n9025 );
or ( n9027 , n8961 , n9026 );
and ( n9028 , n8958 , n9027 );
or ( n9029 , n8957 , n9028 );
and ( n9030 , n8954 , n9029 );
or ( n9031 , n8953 , n9030 );
and ( n9032 , n8950 , n9031 );
or ( n9033 , n8949 , n9032 );
and ( n9034 , n8946 , n9033 );
or ( n9035 , n8945 , n9034 );
and ( n9036 , n816 , n6929 );
and ( n9037 , n9035 , n9036 );
xor ( n9038 , n9035 , n9036 );
xor ( n9039 , n8946 , n9033 );
and ( n9040 , n817 , n6929 );
and ( n9041 , n9039 , n9040 );
xor ( n9042 , n9039 , n9040 );
xor ( n9043 , n8950 , n9031 );
and ( n9044 , n818 , n6929 );
and ( n9045 , n9043 , n9044 );
xor ( n9046 , n9043 , n9044 );
xor ( n9047 , n8954 , n9029 );
and ( n9048 , n819 , n6929 );
and ( n9049 , n9047 , n9048 );
xor ( n9050 , n9047 , n9048 );
xor ( n9051 , n8958 , n9027 );
and ( n9052 , n820 , n6929 );
and ( n9053 , n9051 , n9052 );
xor ( n9054 , n9051 , n9052 );
xor ( n9055 , n8962 , n9025 );
and ( n9056 , n821 , n6929 );
and ( n9057 , n9055 , n9056 );
xor ( n9058 , n9055 , n9056 );
xor ( n9059 , n8966 , n9023 );
and ( n9060 , n822 , n6929 );
and ( n9061 , n9059 , n9060 );
xor ( n9062 , n9059 , n9060 );
xor ( n9063 , n8970 , n9021 );
and ( n9064 , n823 , n6929 );
and ( n9065 , n9063 , n9064 );
xor ( n9066 , n9063 , n9064 );
xor ( n9067 , n8974 , n9019 );
and ( n9068 , n824 , n6929 );
and ( n9069 , n9067 , n9068 );
xor ( n9070 , n9067 , n9068 );
xor ( n9071 , n8978 , n9017 );
and ( n9072 , n825 , n6929 );
and ( n9073 , n9071 , n9072 );
xor ( n9074 , n9071 , n9072 );
xor ( n9075 , n8982 , n9015 );
and ( n9076 , n826 , n6929 );
and ( n9077 , n9075 , n9076 );
xor ( n9078 , n9075 , n9076 );
xor ( n9079 , n8986 , n9013 );
and ( n9080 , n827 , n6929 );
and ( n9081 , n9079 , n9080 );
xor ( n9082 , n9079 , n9080 );
xor ( n9083 , n8990 , n9011 );
and ( n9084 , n828 , n6929 );
and ( n9085 , n9083 , n9084 );
xor ( n9086 , n9083 , n9084 );
xor ( n9087 , n8994 , n9009 );
and ( n9088 , n829 , n6929 );
and ( n9089 , n9087 , n9088 );
xor ( n9090 , n9087 , n9088 );
xor ( n9091 , n8998 , n9007 );
and ( n9092 , n830 , n6929 );
and ( n9093 , n9091 , n9092 );
xor ( n9094 , n9091 , n9092 );
xor ( n9095 , n9002 , n9005 );
and ( n9096 , n831 , n6929 );
and ( n9097 , n9095 , n9096 );
and ( n9098 , n9094 , n9097 );
or ( n9099 , n9093 , n9098 );
and ( n9100 , n9090 , n9099 );
or ( n9101 , n9089 , n9100 );
and ( n9102 , n9086 , n9101 );
or ( n9103 , n9085 , n9102 );
and ( n9104 , n9082 , n9103 );
or ( n9105 , n9081 , n9104 );
and ( n9106 , n9078 , n9105 );
or ( n9107 , n9077 , n9106 );
and ( n9108 , n9074 , n9107 );
or ( n9109 , n9073 , n9108 );
and ( n9110 , n9070 , n9109 );
or ( n9111 , n9069 , n9110 );
and ( n9112 , n9066 , n9111 );
or ( n9113 , n9065 , n9112 );
and ( n9114 , n9062 , n9113 );
or ( n9115 , n9061 , n9114 );
and ( n9116 , n9058 , n9115 );
or ( n9117 , n9057 , n9116 );
and ( n9118 , n9054 , n9117 );
or ( n9119 , n9053 , n9118 );
and ( n9120 , n9050 , n9119 );
or ( n9121 , n9049 , n9120 );
and ( n9122 , n9046 , n9121 );
or ( n9123 , n9045 , n9122 );
and ( n9124 , n9042 , n9123 );
or ( n9125 , n9041 , n9124 );
and ( n9126 , n9038 , n9125 );
or ( n9127 , n9037 , n9126 );
and ( n9128 , n816 , n6926 );
and ( n9129 , n9127 , n9128 );
xor ( n9130 , n9127 , n9128 );
xor ( n9131 , n9038 , n9125 );
and ( n9132 , n817 , n6926 );
and ( n9133 , n9131 , n9132 );
xor ( n9134 , n9131 , n9132 );
xor ( n9135 , n9042 , n9123 );
and ( n9136 , n818 , n6926 );
and ( n9137 , n9135 , n9136 );
xor ( n9138 , n9135 , n9136 );
xor ( n9139 , n9046 , n9121 );
and ( n9140 , n819 , n6926 );
and ( n9141 , n9139 , n9140 );
xor ( n9142 , n9139 , n9140 );
xor ( n9143 , n9050 , n9119 );
and ( n9144 , n820 , n6926 );
and ( n9145 , n9143 , n9144 );
xor ( n9146 , n9143 , n9144 );
xor ( n9147 , n9054 , n9117 );
and ( n9148 , n821 , n6926 );
and ( n9149 , n9147 , n9148 );
xor ( n9150 , n9147 , n9148 );
xor ( n9151 , n9058 , n9115 );
and ( n9152 , n822 , n6926 );
and ( n9153 , n9151 , n9152 );
xor ( n9154 , n9151 , n9152 );
xor ( n9155 , n9062 , n9113 );
and ( n9156 , n823 , n6926 );
and ( n9157 , n9155 , n9156 );
xor ( n9158 , n9155 , n9156 );
xor ( n9159 , n9066 , n9111 );
and ( n9160 , n824 , n6926 );
and ( n9161 , n9159 , n9160 );
xor ( n9162 , n9159 , n9160 );
xor ( n9163 , n9070 , n9109 );
and ( n9164 , n825 , n6926 );
and ( n9165 , n9163 , n9164 );
xor ( n9166 , n9163 , n9164 );
xor ( n9167 , n9074 , n9107 );
and ( n9168 , n826 , n6926 );
and ( n9169 , n9167 , n9168 );
xor ( n9170 , n9167 , n9168 );
xor ( n9171 , n9078 , n9105 );
and ( n9172 , n827 , n6926 );
and ( n9173 , n9171 , n9172 );
xor ( n9174 , n9171 , n9172 );
xor ( n9175 , n9082 , n9103 );
and ( n9176 , n828 , n6926 );
and ( n9177 , n9175 , n9176 );
xor ( n9178 , n9175 , n9176 );
xor ( n9179 , n9086 , n9101 );
and ( n9180 , n829 , n6926 );
and ( n9181 , n9179 , n9180 );
xor ( n9182 , n9179 , n9180 );
xor ( n9183 , n9090 , n9099 );
and ( n9184 , n830 , n6926 );
and ( n9185 , n9183 , n9184 );
xor ( n9186 , n9183 , n9184 );
xor ( n9187 , n9094 , n9097 );
and ( n9188 , n831 , n6926 );
and ( n9189 , n9187 , n9188 );
and ( n9190 , n9186 , n9189 );
or ( n9191 , n9185 , n9190 );
and ( n9192 , n9182 , n9191 );
or ( n9193 , n9181 , n9192 );
and ( n9194 , n9178 , n9193 );
or ( n9195 , n9177 , n9194 );
and ( n9196 , n9174 , n9195 );
or ( n9197 , n9173 , n9196 );
and ( n9198 , n9170 , n9197 );
or ( n9199 , n9169 , n9198 );
and ( n9200 , n9166 , n9199 );
or ( n9201 , n9165 , n9200 );
and ( n9202 , n9162 , n9201 );
or ( n9203 , n9161 , n9202 );
and ( n9204 , n9158 , n9203 );
or ( n9205 , n9157 , n9204 );
and ( n9206 , n9154 , n9205 );
or ( n9207 , n9153 , n9206 );
and ( n9208 , n9150 , n9207 );
or ( n9209 , n9149 , n9208 );
and ( n9210 , n9146 , n9209 );
or ( n9211 , n9145 , n9210 );
and ( n9212 , n9142 , n9211 );
or ( n9213 , n9141 , n9212 );
and ( n9214 , n9138 , n9213 );
or ( n9215 , n9137 , n9214 );
and ( n9216 , n9134 , n9215 );
or ( n9217 , n9133 , n9216 );
and ( n9218 , n9130 , n9217 );
or ( n9219 , n9129 , n9218 );
and ( n9220 , n816 , n6923 );
and ( n9221 , n9219 , n9220 );
xor ( n9222 , n9219 , n9220 );
xor ( n9223 , n9130 , n9217 );
and ( n9224 , n817 , n6923 );
and ( n9225 , n9223 , n9224 );
xor ( n9226 , n9223 , n9224 );
xor ( n9227 , n9134 , n9215 );
and ( n9228 , n818 , n6923 );
and ( n9229 , n9227 , n9228 );
xor ( n9230 , n9227 , n9228 );
xor ( n9231 , n9138 , n9213 );
and ( n9232 , n819 , n6923 );
and ( n9233 , n9231 , n9232 );
xor ( n9234 , n9231 , n9232 );
xor ( n9235 , n9142 , n9211 );
and ( n9236 , n820 , n6923 );
and ( n9237 , n9235 , n9236 );
xor ( n9238 , n9235 , n9236 );
xor ( n9239 , n9146 , n9209 );
and ( n9240 , n821 , n6923 );
and ( n9241 , n9239 , n9240 );
xor ( n9242 , n9239 , n9240 );
xor ( n9243 , n9150 , n9207 );
and ( n9244 , n822 , n6923 );
and ( n9245 , n9243 , n9244 );
xor ( n9246 , n9243 , n9244 );
xor ( n9247 , n9154 , n9205 );
and ( n9248 , n823 , n6923 );
and ( n9249 , n9247 , n9248 );
xor ( n9250 , n9247 , n9248 );
xor ( n9251 , n9158 , n9203 );
and ( n9252 , n824 , n6923 );
and ( n9253 , n9251 , n9252 );
xor ( n9254 , n9251 , n9252 );
xor ( n9255 , n9162 , n9201 );
and ( n9256 , n825 , n6923 );
and ( n9257 , n9255 , n9256 );
xor ( n9258 , n9255 , n9256 );
xor ( n9259 , n9166 , n9199 );
and ( n9260 , n826 , n6923 );
and ( n9261 , n9259 , n9260 );
xor ( n9262 , n9259 , n9260 );
xor ( n9263 , n9170 , n9197 );
and ( n9264 , n827 , n6923 );
and ( n9265 , n9263 , n9264 );
xor ( n9266 , n9263 , n9264 );
xor ( n9267 , n9174 , n9195 );
and ( n9268 , n828 , n6923 );
and ( n9269 , n9267 , n9268 );
xor ( n9270 , n9267 , n9268 );
xor ( n9271 , n9178 , n9193 );
and ( n9272 , n829 , n6923 );
and ( n9273 , n9271 , n9272 );
xor ( n9274 , n9271 , n9272 );
xor ( n9275 , n9182 , n9191 );
and ( n9276 , n830 , n6923 );
and ( n9277 , n9275 , n9276 );
xor ( n9278 , n9275 , n9276 );
xor ( n9279 , n9186 , n9189 );
and ( n9280 , n831 , n6923 );
and ( n9281 , n9279 , n9280 );
and ( n9282 , n9278 , n9281 );
or ( n9283 , n9277 , n9282 );
and ( n9284 , n9274 , n9283 );
or ( n9285 , n9273 , n9284 );
and ( n9286 , n9270 , n9285 );
or ( n9287 , n9269 , n9286 );
and ( n9288 , n9266 , n9287 );
or ( n9289 , n9265 , n9288 );
and ( n9290 , n9262 , n9289 );
or ( n9291 , n9261 , n9290 );
and ( n9292 , n9258 , n9291 );
or ( n9293 , n9257 , n9292 );
and ( n9294 , n9254 , n9293 );
or ( n9295 , n9253 , n9294 );
and ( n9296 , n9250 , n9295 );
or ( n9297 , n9249 , n9296 );
and ( n9298 , n9246 , n9297 );
or ( n9299 , n9245 , n9298 );
and ( n9300 , n9242 , n9299 );
or ( n9301 , n9241 , n9300 );
and ( n9302 , n9238 , n9301 );
or ( n9303 , n9237 , n9302 );
and ( n9304 , n9234 , n9303 );
or ( n9305 , n9233 , n9304 );
and ( n9306 , n9230 , n9305 );
or ( n9307 , n9229 , n9306 );
and ( n9308 , n9226 , n9307 );
or ( n9309 , n9225 , n9308 );
and ( n9310 , n9222 , n9309 );
or ( n9311 , n9221 , n9310 );
and ( n9312 , n816 , n6920 );
and ( n9313 , n9311 , n9312 );
xor ( n9314 , n9311 , n9312 );
xor ( n9315 , n9222 , n9309 );
and ( n9316 , n817 , n6920 );
and ( n9317 , n9315 , n9316 );
xor ( n9318 , n9315 , n9316 );
xor ( n9319 , n9226 , n9307 );
and ( n9320 , n818 , n6920 );
and ( n9321 , n9319 , n9320 );
xor ( n9322 , n9319 , n9320 );
xor ( n9323 , n9230 , n9305 );
and ( n9324 , n819 , n6920 );
and ( n9325 , n9323 , n9324 );
xor ( n9326 , n9323 , n9324 );
xor ( n9327 , n9234 , n9303 );
and ( n9328 , n820 , n6920 );
and ( n9329 , n9327 , n9328 );
xor ( n9330 , n9327 , n9328 );
xor ( n9331 , n9238 , n9301 );
and ( n9332 , n821 , n6920 );
and ( n9333 , n9331 , n9332 );
xor ( n9334 , n9331 , n9332 );
xor ( n9335 , n9242 , n9299 );
and ( n9336 , n822 , n6920 );
and ( n9337 , n9335 , n9336 );
xor ( n9338 , n9335 , n9336 );
xor ( n9339 , n9246 , n9297 );
and ( n9340 , n823 , n6920 );
and ( n9341 , n9339 , n9340 );
xor ( n9342 , n9339 , n9340 );
xor ( n9343 , n9250 , n9295 );
and ( n9344 , n824 , n6920 );
and ( n9345 , n9343 , n9344 );
xor ( n9346 , n9343 , n9344 );
xor ( n9347 , n9254 , n9293 );
and ( n9348 , n825 , n6920 );
and ( n9349 , n9347 , n9348 );
xor ( n9350 , n9347 , n9348 );
xor ( n9351 , n9258 , n9291 );
and ( n9352 , n826 , n6920 );
and ( n9353 , n9351 , n9352 );
xor ( n9354 , n9351 , n9352 );
xor ( n9355 , n9262 , n9289 );
and ( n9356 , n827 , n6920 );
and ( n9357 , n9355 , n9356 );
xor ( n9358 , n9355 , n9356 );
xor ( n9359 , n9266 , n9287 );
and ( n9360 , n828 , n6920 );
and ( n9361 , n9359 , n9360 );
xor ( n9362 , n9359 , n9360 );
xor ( n9363 , n9270 , n9285 );
and ( n9364 , n829 , n6920 );
and ( n9365 , n9363 , n9364 );
xor ( n9366 , n9363 , n9364 );
xor ( n9367 , n9274 , n9283 );
and ( n9368 , n830 , n6920 );
and ( n9369 , n9367 , n9368 );
xor ( n9370 , n9367 , n9368 );
xor ( n9371 , n9278 , n9281 );
and ( n9372 , n831 , n6920 );
and ( n9373 , n9371 , n9372 );
and ( n9374 , n9370 , n9373 );
or ( n9375 , n9369 , n9374 );
and ( n9376 , n9366 , n9375 );
or ( n9377 , n9365 , n9376 );
and ( n9378 , n9362 , n9377 );
or ( n9379 , n9361 , n9378 );
and ( n9380 , n9358 , n9379 );
or ( n9381 , n9357 , n9380 );
and ( n9382 , n9354 , n9381 );
or ( n9383 , n9353 , n9382 );
and ( n9384 , n9350 , n9383 );
or ( n9385 , n9349 , n9384 );
and ( n9386 , n9346 , n9385 );
or ( n9387 , n9345 , n9386 );
and ( n9388 , n9342 , n9387 );
or ( n9389 , n9341 , n9388 );
and ( n9390 , n9338 , n9389 );
or ( n9391 , n9337 , n9390 );
and ( n9392 , n9334 , n9391 );
or ( n9393 , n9333 , n9392 );
and ( n9394 , n9330 , n9393 );
or ( n9395 , n9329 , n9394 );
and ( n9396 , n9326 , n9395 );
or ( n9397 , n9325 , n9396 );
and ( n9398 , n9322 , n9397 );
or ( n9399 , n9321 , n9398 );
and ( n9400 , n9318 , n9399 );
or ( n9401 , n9317 , n9400 );
and ( n9402 , n9314 , n9401 );
or ( n9403 , n9313 , n9402 );
and ( n9404 , n816 , n6917 );
and ( n9405 , n9403 , n9404 );
xor ( n9406 , n9403 , n9404 );
xor ( n9407 , n9314 , n9401 );
and ( n9408 , n817 , n6917 );
and ( n9409 , n9407 , n9408 );
xor ( n9410 , n9407 , n9408 );
xor ( n9411 , n9318 , n9399 );
and ( n9412 , n818 , n6917 );
and ( n9413 , n9411 , n9412 );
xor ( n9414 , n9411 , n9412 );
xor ( n9415 , n9322 , n9397 );
and ( n9416 , n819 , n6917 );
and ( n9417 , n9415 , n9416 );
xor ( n9418 , n9415 , n9416 );
xor ( n9419 , n9326 , n9395 );
and ( n9420 , n820 , n6917 );
and ( n9421 , n9419 , n9420 );
xor ( n9422 , n9419 , n9420 );
xor ( n9423 , n9330 , n9393 );
and ( n9424 , n821 , n6917 );
and ( n9425 , n9423 , n9424 );
xor ( n9426 , n9423 , n9424 );
xor ( n9427 , n9334 , n9391 );
and ( n9428 , n822 , n6917 );
and ( n9429 , n9427 , n9428 );
xor ( n9430 , n9427 , n9428 );
xor ( n9431 , n9338 , n9389 );
and ( n9432 , n823 , n6917 );
and ( n9433 , n9431 , n9432 );
xor ( n9434 , n9431 , n9432 );
xor ( n9435 , n9342 , n9387 );
and ( n9436 , n824 , n6917 );
and ( n9437 , n9435 , n9436 );
xor ( n9438 , n9435 , n9436 );
xor ( n9439 , n9346 , n9385 );
and ( n9440 , n825 , n6917 );
and ( n9441 , n9439 , n9440 );
xor ( n9442 , n9439 , n9440 );
xor ( n9443 , n9350 , n9383 );
and ( n9444 , n826 , n6917 );
and ( n9445 , n9443 , n9444 );
xor ( n9446 , n9443 , n9444 );
xor ( n9447 , n9354 , n9381 );
and ( n9448 , n827 , n6917 );
and ( n9449 , n9447 , n9448 );
xor ( n9450 , n9447 , n9448 );
xor ( n9451 , n9358 , n9379 );
and ( n9452 , n828 , n6917 );
and ( n9453 , n9451 , n9452 );
xor ( n9454 , n9451 , n9452 );
xor ( n9455 , n9362 , n9377 );
and ( n9456 , n829 , n6917 );
and ( n9457 , n9455 , n9456 );
xor ( n9458 , n9455 , n9456 );
xor ( n9459 , n9366 , n9375 );
and ( n9460 , n830 , n6917 );
and ( n9461 , n9459 , n9460 );
xor ( n9462 , n9459 , n9460 );
xor ( n9463 , n9370 , n9373 );
and ( n9464 , n831 , n6917 );
and ( n9465 , n9463 , n9464 );
and ( n9466 , n9462 , n9465 );
or ( n9467 , n9461 , n9466 );
and ( n9468 , n9458 , n9467 );
or ( n9469 , n9457 , n9468 );
and ( n9470 , n9454 , n9469 );
or ( n9471 , n9453 , n9470 );
and ( n9472 , n9450 , n9471 );
or ( n9473 , n9449 , n9472 );
and ( n9474 , n9446 , n9473 );
or ( n9475 , n9445 , n9474 );
and ( n9476 , n9442 , n9475 );
or ( n9477 , n9441 , n9476 );
and ( n9478 , n9438 , n9477 );
or ( n9479 , n9437 , n9478 );
and ( n9480 , n9434 , n9479 );
or ( n9481 , n9433 , n9480 );
and ( n9482 , n9430 , n9481 );
or ( n9483 , n9429 , n9482 );
and ( n9484 , n9426 , n9483 );
or ( n9485 , n9425 , n9484 );
and ( n9486 , n9422 , n9485 );
or ( n9487 , n9421 , n9486 );
and ( n9488 , n9418 , n9487 );
or ( n9489 , n9417 , n9488 );
and ( n9490 , n9414 , n9489 );
or ( n9491 , n9413 , n9490 );
and ( n9492 , n9410 , n9491 );
or ( n9493 , n9409 , n9492 );
and ( n9494 , n9406 , n9493 );
or ( n9495 , n9405 , n9494 );
and ( n9496 , n816 , n6914 );
and ( n9497 , n9495 , n9496 );
xor ( n9498 , n9495 , n9496 );
xor ( n9499 , n9406 , n9493 );
and ( n9500 , n817 , n6914 );
and ( n9501 , n9499 , n9500 );
xor ( n9502 , n9499 , n9500 );
xor ( n9503 , n9410 , n9491 );
and ( n9504 , n818 , n6914 );
and ( n9505 , n9503 , n9504 );
xor ( n9506 , n9503 , n9504 );
xor ( n9507 , n9414 , n9489 );
and ( n9508 , n819 , n6914 );
and ( n9509 , n9507 , n9508 );
xor ( n9510 , n9507 , n9508 );
xor ( n9511 , n9418 , n9487 );
and ( n9512 , n820 , n6914 );
and ( n9513 , n9511 , n9512 );
xor ( n9514 , n9511 , n9512 );
xor ( n9515 , n9422 , n9485 );
and ( n9516 , n821 , n6914 );
and ( n9517 , n9515 , n9516 );
xor ( n9518 , n9515 , n9516 );
xor ( n9519 , n9426 , n9483 );
and ( n9520 , n822 , n6914 );
and ( n9521 , n9519 , n9520 );
xor ( n9522 , n9519 , n9520 );
xor ( n9523 , n9430 , n9481 );
and ( n9524 , n823 , n6914 );
and ( n9525 , n9523 , n9524 );
xor ( n9526 , n9523 , n9524 );
xor ( n9527 , n9434 , n9479 );
and ( n9528 , n824 , n6914 );
and ( n9529 , n9527 , n9528 );
xor ( n9530 , n9527 , n9528 );
xor ( n9531 , n9438 , n9477 );
and ( n9532 , n825 , n6914 );
and ( n9533 , n9531 , n9532 );
xor ( n9534 , n9531 , n9532 );
xor ( n9535 , n9442 , n9475 );
and ( n9536 , n826 , n6914 );
and ( n9537 , n9535 , n9536 );
xor ( n9538 , n9535 , n9536 );
xor ( n9539 , n9446 , n9473 );
and ( n9540 , n827 , n6914 );
and ( n9541 , n9539 , n9540 );
xor ( n9542 , n9539 , n9540 );
xor ( n9543 , n9450 , n9471 );
and ( n9544 , n828 , n6914 );
and ( n9545 , n9543 , n9544 );
xor ( n9546 , n9543 , n9544 );
xor ( n9547 , n9454 , n9469 );
and ( n9548 , n829 , n6914 );
and ( n9549 , n9547 , n9548 );
xor ( n9550 , n9547 , n9548 );
xor ( n9551 , n9458 , n9467 );
and ( n9552 , n830 , n6914 );
and ( n9553 , n9551 , n9552 );
xor ( n9554 , n9551 , n9552 );
xor ( n9555 , n9462 , n9465 );
and ( n9556 , n831 , n6914 );
and ( n9557 , n9555 , n9556 );
and ( n9558 , n9554 , n9557 );
or ( n9559 , n9553 , n9558 );
and ( n9560 , n9550 , n9559 );
or ( n9561 , n9549 , n9560 );
and ( n9562 , n9546 , n9561 );
or ( n9563 , n9545 , n9562 );
and ( n9564 , n9542 , n9563 );
or ( n9565 , n9541 , n9564 );
and ( n9566 , n9538 , n9565 );
or ( n9567 , n9537 , n9566 );
and ( n9568 , n9534 , n9567 );
or ( n9569 , n9533 , n9568 );
and ( n9570 , n9530 , n9569 );
or ( n9571 , n9529 , n9570 );
and ( n9572 , n9526 , n9571 );
or ( n9573 , n9525 , n9572 );
and ( n9574 , n9522 , n9573 );
or ( n9575 , n9521 , n9574 );
and ( n9576 , n9518 , n9575 );
or ( n9577 , n9517 , n9576 );
and ( n9578 , n9514 , n9577 );
or ( n9579 , n9513 , n9578 );
and ( n9580 , n9510 , n9579 );
or ( n9581 , n9509 , n9580 );
and ( n9582 , n9506 , n9581 );
or ( n9583 , n9505 , n9582 );
and ( n9584 , n9502 , n9583 );
or ( n9585 , n9501 , n9584 );
and ( n9586 , n9498 , n9585 );
or ( n9587 , n9497 , n9586 );
and ( n9588 , n816 , n6911 );
and ( n9589 , n9587 , n9588 );
xor ( n9590 , n9587 , n9588 );
xor ( n9591 , n9498 , n9585 );
and ( n9592 , n817 , n6911 );
and ( n9593 , n9591 , n9592 );
xor ( n9594 , n9591 , n9592 );
xor ( n9595 , n9502 , n9583 );
and ( n9596 , n818 , n6911 );
and ( n9597 , n9595 , n9596 );
xor ( n9598 , n9595 , n9596 );
xor ( n9599 , n9506 , n9581 );
and ( n9600 , n819 , n6911 );
and ( n9601 , n9599 , n9600 );
xor ( n9602 , n9599 , n9600 );
xor ( n9603 , n9510 , n9579 );
and ( n9604 , n820 , n6911 );
and ( n9605 , n9603 , n9604 );
xor ( n9606 , n9603 , n9604 );
xor ( n9607 , n9514 , n9577 );
and ( n9608 , n821 , n6911 );
and ( n9609 , n9607 , n9608 );
xor ( n9610 , n9607 , n9608 );
xor ( n9611 , n9518 , n9575 );
and ( n9612 , n822 , n6911 );
and ( n9613 , n9611 , n9612 );
xor ( n9614 , n9611 , n9612 );
xor ( n9615 , n9522 , n9573 );
and ( n9616 , n823 , n6911 );
and ( n9617 , n9615 , n9616 );
xor ( n9618 , n9615 , n9616 );
xor ( n9619 , n9526 , n9571 );
and ( n9620 , n824 , n6911 );
and ( n9621 , n9619 , n9620 );
xor ( n9622 , n9619 , n9620 );
xor ( n9623 , n9530 , n9569 );
and ( n9624 , n825 , n6911 );
and ( n9625 , n9623 , n9624 );
xor ( n9626 , n9623 , n9624 );
xor ( n9627 , n9534 , n9567 );
and ( n9628 , n826 , n6911 );
and ( n9629 , n9627 , n9628 );
xor ( n9630 , n9627 , n9628 );
xor ( n9631 , n9538 , n9565 );
and ( n9632 , n827 , n6911 );
and ( n9633 , n9631 , n9632 );
xor ( n9634 , n9631 , n9632 );
xor ( n9635 , n9542 , n9563 );
and ( n9636 , n828 , n6911 );
and ( n9637 , n9635 , n9636 );
xor ( n9638 , n9635 , n9636 );
xor ( n9639 , n9546 , n9561 );
and ( n9640 , n829 , n6911 );
and ( n9641 , n9639 , n9640 );
xor ( n9642 , n9639 , n9640 );
xor ( n9643 , n9550 , n9559 );
and ( n9644 , n830 , n6911 );
and ( n9645 , n9643 , n9644 );
xor ( n9646 , n9643 , n9644 );
xor ( n9647 , n9554 , n9557 );
and ( n9648 , n831 , n6911 );
and ( n9649 , n9647 , n9648 );
and ( n9650 , n9646 , n9649 );
or ( n9651 , n9645 , n9650 );
and ( n9652 , n9642 , n9651 );
or ( n9653 , n9641 , n9652 );
and ( n9654 , n9638 , n9653 );
or ( n9655 , n9637 , n9654 );
and ( n9656 , n9634 , n9655 );
or ( n9657 , n9633 , n9656 );
and ( n9658 , n9630 , n9657 );
or ( n9659 , n9629 , n9658 );
and ( n9660 , n9626 , n9659 );
or ( n9661 , n9625 , n9660 );
and ( n9662 , n9622 , n9661 );
or ( n9663 , n9621 , n9662 );
and ( n9664 , n9618 , n9663 );
or ( n9665 , n9617 , n9664 );
and ( n9666 , n9614 , n9665 );
or ( n9667 , n9613 , n9666 );
and ( n9668 , n9610 , n9667 );
or ( n9669 , n9609 , n9668 );
and ( n9670 , n9606 , n9669 );
or ( n9671 , n9605 , n9670 );
and ( n9672 , n9602 , n9671 );
or ( n9673 , n9601 , n9672 );
and ( n9674 , n9598 , n9673 );
or ( n9675 , n9597 , n9674 );
and ( n9676 , n9594 , n9675 );
or ( n9677 , n9593 , n9676 );
and ( n9678 , n9590 , n9677 );
or ( n9679 , n9589 , n9678 );
and ( n9680 , n816 , n6908 );
and ( n9681 , n9679 , n9680 );
xor ( n9682 , n9679 , n9680 );
xor ( n9683 , n9590 , n9677 );
and ( n9684 , n817 , n6908 );
and ( n9685 , n9683 , n9684 );
xor ( n9686 , n9683 , n9684 );
xor ( n9687 , n9594 , n9675 );
and ( n9688 , n818 , n6908 );
and ( n9689 , n9687 , n9688 );
xor ( n9690 , n9687 , n9688 );
xor ( n9691 , n9598 , n9673 );
and ( n9692 , n819 , n6908 );
and ( n9693 , n9691 , n9692 );
xor ( n9694 , n9691 , n9692 );
xor ( n9695 , n9602 , n9671 );
and ( n9696 , n820 , n6908 );
and ( n9697 , n9695 , n9696 );
xor ( n9698 , n9695 , n9696 );
xor ( n9699 , n9606 , n9669 );
and ( n9700 , n821 , n6908 );
and ( n9701 , n9699 , n9700 );
xor ( n9702 , n9699 , n9700 );
xor ( n9703 , n9610 , n9667 );
and ( n9704 , n822 , n6908 );
and ( n9705 , n9703 , n9704 );
xor ( n9706 , n9703 , n9704 );
xor ( n9707 , n9614 , n9665 );
and ( n9708 , n823 , n6908 );
and ( n9709 , n9707 , n9708 );
xor ( n9710 , n9707 , n9708 );
xor ( n9711 , n9618 , n9663 );
and ( n9712 , n824 , n6908 );
and ( n9713 , n9711 , n9712 );
xor ( n9714 , n9711 , n9712 );
xor ( n9715 , n9622 , n9661 );
and ( n9716 , n825 , n6908 );
and ( n9717 , n9715 , n9716 );
xor ( n9718 , n9715 , n9716 );
xor ( n9719 , n9626 , n9659 );
and ( n9720 , n826 , n6908 );
and ( n9721 , n9719 , n9720 );
xor ( n9722 , n9719 , n9720 );
xor ( n9723 , n9630 , n9657 );
and ( n9724 , n827 , n6908 );
and ( n9725 , n9723 , n9724 );
xor ( n9726 , n9723 , n9724 );
xor ( n9727 , n9634 , n9655 );
and ( n9728 , n828 , n6908 );
and ( n9729 , n9727 , n9728 );
xor ( n9730 , n9727 , n9728 );
xor ( n9731 , n9638 , n9653 );
and ( n9732 , n829 , n6908 );
and ( n9733 , n9731 , n9732 );
xor ( n9734 , n9731 , n9732 );
xor ( n9735 , n9642 , n9651 );
and ( n9736 , n830 , n6908 );
and ( n9737 , n9735 , n9736 );
xor ( n9738 , n9735 , n9736 );
xor ( n9739 , n9646 , n9649 );
and ( n9740 , n831 , n6908 );
and ( n9741 , n9739 , n9740 );
and ( n9742 , n9738 , n9741 );
or ( n9743 , n9737 , n9742 );
and ( n9744 , n9734 , n9743 );
or ( n9745 , n9733 , n9744 );
and ( n9746 , n9730 , n9745 );
or ( n9747 , n9729 , n9746 );
and ( n9748 , n9726 , n9747 );
or ( n9749 , n9725 , n9748 );
and ( n9750 , n9722 , n9749 );
or ( n9751 , n9721 , n9750 );
and ( n9752 , n9718 , n9751 );
or ( n9753 , n9717 , n9752 );
and ( n9754 , n9714 , n9753 );
or ( n9755 , n9713 , n9754 );
and ( n9756 , n9710 , n9755 );
or ( n9757 , n9709 , n9756 );
and ( n9758 , n9706 , n9757 );
or ( n9759 , n9705 , n9758 );
and ( n9760 , n9702 , n9759 );
or ( n9761 , n9701 , n9760 );
and ( n9762 , n9698 , n9761 );
or ( n9763 , n9697 , n9762 );
and ( n9764 , n9694 , n9763 );
or ( n9765 , n9693 , n9764 );
and ( n9766 , n9690 , n9765 );
or ( n9767 , n9689 , n9766 );
and ( n9768 , n9686 , n9767 );
or ( n9769 , n9685 , n9768 );
and ( n9770 , n9682 , n9769 );
or ( n9771 , n9681 , n9770 );
and ( n9772 , n816 , n6905 );
and ( n9773 , n9771 , n9772 );
xor ( n9774 , n9771 , n9772 );
xor ( n9775 , n9682 , n9769 );
and ( n9776 , n817 , n6905 );
and ( n9777 , n9775 , n9776 );
xor ( n9778 , n9775 , n9776 );
xor ( n9779 , n9686 , n9767 );
and ( n9780 , n818 , n6905 );
and ( n9781 , n9779 , n9780 );
xor ( n9782 , n9779 , n9780 );
xor ( n9783 , n9690 , n9765 );
and ( n9784 , n819 , n6905 );
and ( n9785 , n9783 , n9784 );
xor ( n9786 , n9783 , n9784 );
xor ( n9787 , n9694 , n9763 );
and ( n9788 , n820 , n6905 );
and ( n9789 , n9787 , n9788 );
xor ( n9790 , n9787 , n9788 );
xor ( n9791 , n9698 , n9761 );
and ( n9792 , n821 , n6905 );
and ( n9793 , n9791 , n9792 );
xor ( n9794 , n9791 , n9792 );
xor ( n9795 , n9702 , n9759 );
and ( n9796 , n822 , n6905 );
and ( n9797 , n9795 , n9796 );
xor ( n9798 , n9795 , n9796 );
xor ( n9799 , n9706 , n9757 );
and ( n9800 , n823 , n6905 );
and ( n9801 , n9799 , n9800 );
xor ( n9802 , n9799 , n9800 );
xor ( n9803 , n9710 , n9755 );
and ( n9804 , n824 , n6905 );
and ( n9805 , n9803 , n9804 );
xor ( n9806 , n9803 , n9804 );
xor ( n9807 , n9714 , n9753 );
and ( n9808 , n825 , n6905 );
and ( n9809 , n9807 , n9808 );
xor ( n9810 , n9807 , n9808 );
xor ( n9811 , n9718 , n9751 );
and ( n9812 , n826 , n6905 );
and ( n9813 , n9811 , n9812 );
xor ( n9814 , n9811 , n9812 );
xor ( n9815 , n9722 , n9749 );
and ( n9816 , n827 , n6905 );
and ( n9817 , n9815 , n9816 );
xor ( n9818 , n9815 , n9816 );
xor ( n9819 , n9726 , n9747 );
and ( n9820 , n828 , n6905 );
and ( n9821 , n9819 , n9820 );
xor ( n9822 , n9819 , n9820 );
xor ( n9823 , n9730 , n9745 );
and ( n9824 , n829 , n6905 );
and ( n9825 , n9823 , n9824 );
xor ( n9826 , n9823 , n9824 );
xor ( n9827 , n9734 , n9743 );
and ( n9828 , n830 , n6905 );
and ( n9829 , n9827 , n9828 );
xor ( n9830 , n9827 , n9828 );
xor ( n9831 , n9738 , n9741 );
and ( n9832 , n831 , n6905 );
and ( n9833 , n9831 , n9832 );
and ( n9834 , n9830 , n9833 );
or ( n9835 , n9829 , n9834 );
and ( n9836 , n9826 , n9835 );
or ( n9837 , n9825 , n9836 );
and ( n9838 , n9822 , n9837 );
or ( n9839 , n9821 , n9838 );
and ( n9840 , n9818 , n9839 );
or ( n9841 , n9817 , n9840 );
and ( n9842 , n9814 , n9841 );
or ( n9843 , n9813 , n9842 );
and ( n9844 , n9810 , n9843 );
or ( n9845 , n9809 , n9844 );
and ( n9846 , n9806 , n9845 );
or ( n9847 , n9805 , n9846 );
and ( n9848 , n9802 , n9847 );
or ( n9849 , n9801 , n9848 );
and ( n9850 , n9798 , n9849 );
or ( n9851 , n9797 , n9850 );
and ( n9852 , n9794 , n9851 );
or ( n9853 , n9793 , n9852 );
and ( n9854 , n9790 , n9853 );
or ( n9855 , n9789 , n9854 );
and ( n9856 , n9786 , n9855 );
or ( n9857 , n9785 , n9856 );
and ( n9858 , n9782 , n9857 );
or ( n9859 , n9781 , n9858 );
and ( n9860 , n9778 , n9859 );
or ( n9861 , n9777 , n9860 );
and ( n9862 , n9774 , n9861 );
or ( n9863 , n9773 , n9862 );
and ( n9864 , n816 , n6902 );
and ( n9865 , n9863 , n9864 );
xor ( n9866 , n9863 , n9864 );
xor ( n9867 , n9774 , n9861 );
and ( n9868 , n817 , n6902 );
and ( n9869 , n9867 , n9868 );
xor ( n9870 , n9867 , n9868 );
xor ( n9871 , n9778 , n9859 );
and ( n9872 , n818 , n6902 );
and ( n9873 , n9871 , n9872 );
xor ( n9874 , n9871 , n9872 );
xor ( n9875 , n9782 , n9857 );
and ( n9876 , n819 , n6902 );
and ( n9877 , n9875 , n9876 );
xor ( n9878 , n9875 , n9876 );
xor ( n9879 , n9786 , n9855 );
and ( n9880 , n820 , n6902 );
and ( n9881 , n9879 , n9880 );
xor ( n9882 , n9879 , n9880 );
xor ( n9883 , n9790 , n9853 );
and ( n9884 , n821 , n6902 );
and ( n9885 , n9883 , n9884 );
xor ( n9886 , n9883 , n9884 );
xor ( n9887 , n9794 , n9851 );
and ( n9888 , n822 , n6902 );
and ( n9889 , n9887 , n9888 );
xor ( n9890 , n9887 , n9888 );
xor ( n9891 , n9798 , n9849 );
and ( n9892 , n823 , n6902 );
and ( n9893 , n9891 , n9892 );
xor ( n9894 , n9891 , n9892 );
xor ( n9895 , n9802 , n9847 );
and ( n9896 , n824 , n6902 );
and ( n9897 , n9895 , n9896 );
xor ( n9898 , n9895 , n9896 );
xor ( n9899 , n9806 , n9845 );
and ( n9900 , n825 , n6902 );
and ( n9901 , n9899 , n9900 );
xor ( n9902 , n9899 , n9900 );
xor ( n9903 , n9810 , n9843 );
and ( n9904 , n826 , n6902 );
and ( n9905 , n9903 , n9904 );
xor ( n9906 , n9903 , n9904 );
xor ( n9907 , n9814 , n9841 );
and ( n9908 , n827 , n6902 );
and ( n9909 , n9907 , n9908 );
xor ( n9910 , n9907 , n9908 );
xor ( n9911 , n9818 , n9839 );
and ( n9912 , n828 , n6902 );
and ( n9913 , n9911 , n9912 );
xor ( n9914 , n9911 , n9912 );
xor ( n9915 , n9822 , n9837 );
and ( n9916 , n829 , n6902 );
and ( n9917 , n9915 , n9916 );
xor ( n9918 , n9915 , n9916 );
xor ( n9919 , n9826 , n9835 );
and ( n9920 , n830 , n6902 );
and ( n9921 , n9919 , n9920 );
xor ( n9922 , n9919 , n9920 );
xor ( n9923 , n9830 , n9833 );
and ( n9924 , n831 , n6902 );
and ( n9925 , n9923 , n9924 );
and ( n9926 , n9922 , n9925 );
or ( n9927 , n9921 , n9926 );
and ( n9928 , n9918 , n9927 );
or ( n9929 , n9917 , n9928 );
and ( n9930 , n9914 , n9929 );
or ( n9931 , n9913 , n9930 );
and ( n9932 , n9910 , n9931 );
or ( n9933 , n9909 , n9932 );
and ( n9934 , n9906 , n9933 );
or ( n9935 , n9905 , n9934 );
and ( n9936 , n9902 , n9935 );
or ( n9937 , n9901 , n9936 );
and ( n9938 , n9898 , n9937 );
or ( n9939 , n9897 , n9938 );
and ( n9940 , n9894 , n9939 );
or ( n9941 , n9893 , n9940 );
and ( n9942 , n9890 , n9941 );
or ( n9943 , n9889 , n9942 );
and ( n9944 , n9886 , n9943 );
or ( n9945 , n9885 , n9944 );
and ( n9946 , n9882 , n9945 );
or ( n9947 , n9881 , n9946 );
and ( n9948 , n9878 , n9947 );
or ( n9949 , n9877 , n9948 );
and ( n9950 , n9874 , n9949 );
or ( n9951 , n9873 , n9950 );
and ( n9952 , n9870 , n9951 );
or ( n9953 , n9869 , n9952 );
and ( n9954 , n9866 , n9953 );
or ( n9955 , n9865 , n9954 );
and ( n9956 , n816 , n6899 );
and ( n9957 , n9955 , n9956 );
xor ( n9958 , n9955 , n9956 );
xor ( n9959 , n9866 , n9953 );
and ( n9960 , n817 , n6899 );
and ( n9961 , n9959 , n9960 );
xor ( n9962 , n9959 , n9960 );
xor ( n9963 , n9870 , n9951 );
and ( n9964 , n818 , n6899 );
and ( n9965 , n9963 , n9964 );
xor ( n9966 , n9963 , n9964 );
xor ( n9967 , n9874 , n9949 );
and ( n9968 , n819 , n6899 );
and ( n9969 , n9967 , n9968 );
xor ( n9970 , n9967 , n9968 );
xor ( n9971 , n9878 , n9947 );
and ( n9972 , n820 , n6899 );
and ( n9973 , n9971 , n9972 );
xor ( n9974 , n9971 , n9972 );
xor ( n9975 , n9882 , n9945 );
and ( n9976 , n821 , n6899 );
and ( n9977 , n9975 , n9976 );
xor ( n9978 , n9975 , n9976 );
xor ( n9979 , n9886 , n9943 );
and ( n9980 , n822 , n6899 );
and ( n9981 , n9979 , n9980 );
xor ( n9982 , n9979 , n9980 );
xor ( n9983 , n9890 , n9941 );
and ( n9984 , n823 , n6899 );
and ( n9985 , n9983 , n9984 );
xor ( n9986 , n9983 , n9984 );
xor ( n9987 , n9894 , n9939 );
and ( n9988 , n824 , n6899 );
and ( n9989 , n9987 , n9988 );
xor ( n9990 , n9987 , n9988 );
xor ( n9991 , n9898 , n9937 );
and ( n9992 , n825 , n6899 );
and ( n9993 , n9991 , n9992 );
xor ( n9994 , n9991 , n9992 );
xor ( n9995 , n9902 , n9935 );
and ( n9996 , n826 , n6899 );
and ( n9997 , n9995 , n9996 );
xor ( n9998 , n9995 , n9996 );
xor ( n9999 , n9906 , n9933 );
and ( n10000 , n827 , n6899 );
and ( n10001 , n9999 , n10000 );
xor ( n10002 , n9999 , n10000 );
xor ( n10003 , n9910 , n9931 );
and ( n10004 , n828 , n6899 );
and ( n10005 , n10003 , n10004 );
xor ( n10006 , n10003 , n10004 );
xor ( n10007 , n9914 , n9929 );
and ( n10008 , n829 , n6899 );
and ( n10009 , n10007 , n10008 );
xor ( n10010 , n10007 , n10008 );
xor ( n10011 , n9918 , n9927 );
and ( n10012 , n830 , n6899 );
and ( n10013 , n10011 , n10012 );
xor ( n10014 , n10011 , n10012 );
xor ( n10015 , n9922 , n9925 );
and ( n10016 , n831 , n6899 );
and ( n10017 , n10015 , n10016 );
and ( n10018 , n10014 , n10017 );
or ( n10019 , n10013 , n10018 );
and ( n10020 , n10010 , n10019 );
or ( n10021 , n10009 , n10020 );
and ( n10022 , n10006 , n10021 );
or ( n10023 , n10005 , n10022 );
and ( n10024 , n10002 , n10023 );
or ( n10025 , n10001 , n10024 );
and ( n10026 , n9998 , n10025 );
or ( n10027 , n9997 , n10026 );
and ( n10028 , n9994 , n10027 );
or ( n10029 , n9993 , n10028 );
and ( n10030 , n9990 , n10029 );
or ( n10031 , n9989 , n10030 );
and ( n10032 , n9986 , n10031 );
or ( n10033 , n9985 , n10032 );
and ( n10034 , n9982 , n10033 );
or ( n10035 , n9981 , n10034 );
and ( n10036 , n9978 , n10035 );
or ( n10037 , n9977 , n10036 );
and ( n10038 , n9974 , n10037 );
or ( n10039 , n9973 , n10038 );
and ( n10040 , n9970 , n10039 );
or ( n10041 , n9969 , n10040 );
and ( n10042 , n9966 , n10041 );
or ( n10043 , n9965 , n10042 );
and ( n10044 , n9962 , n10043 );
or ( n10045 , n9961 , n10044 );
and ( n10046 , n9958 , n10045 );
or ( n10047 , n9957 , n10046 );
and ( n10048 , n816 , n6896 );
and ( n10049 , n10047 , n10048 );
xor ( n10050 , n10047 , n10048 );
xor ( n10051 , n9958 , n10045 );
and ( n10052 , n817 , n6896 );
and ( n10053 , n10051 , n10052 );
xor ( n10054 , n10051 , n10052 );
xor ( n10055 , n9962 , n10043 );
and ( n10056 , n818 , n6896 );
and ( n10057 , n10055 , n10056 );
xor ( n10058 , n10055 , n10056 );
xor ( n10059 , n9966 , n10041 );
and ( n10060 , n819 , n6896 );
and ( n10061 , n10059 , n10060 );
xor ( n10062 , n10059 , n10060 );
xor ( n10063 , n9970 , n10039 );
and ( n10064 , n820 , n6896 );
and ( n10065 , n10063 , n10064 );
xor ( n10066 , n10063 , n10064 );
xor ( n10067 , n9974 , n10037 );
and ( n10068 , n821 , n6896 );
and ( n10069 , n10067 , n10068 );
xor ( n10070 , n10067 , n10068 );
xor ( n10071 , n9978 , n10035 );
and ( n10072 , n822 , n6896 );
and ( n10073 , n10071 , n10072 );
xor ( n10074 , n10071 , n10072 );
xor ( n10075 , n9982 , n10033 );
and ( n10076 , n823 , n6896 );
and ( n10077 , n10075 , n10076 );
xor ( n10078 , n10075 , n10076 );
xor ( n10079 , n9986 , n10031 );
and ( n10080 , n824 , n6896 );
and ( n10081 , n10079 , n10080 );
xor ( n10082 , n10079 , n10080 );
xor ( n10083 , n9990 , n10029 );
and ( n10084 , n825 , n6896 );
and ( n10085 , n10083 , n10084 );
xor ( n10086 , n10083 , n10084 );
xor ( n10087 , n9994 , n10027 );
and ( n10088 , n826 , n6896 );
and ( n10089 , n10087 , n10088 );
xor ( n10090 , n10087 , n10088 );
xor ( n10091 , n9998 , n10025 );
and ( n10092 , n827 , n6896 );
and ( n10093 , n10091 , n10092 );
xor ( n10094 , n10091 , n10092 );
xor ( n10095 , n10002 , n10023 );
and ( n10096 , n828 , n6896 );
and ( n10097 , n10095 , n10096 );
xor ( n10098 , n10095 , n10096 );
xor ( n10099 , n10006 , n10021 );
and ( n10100 , n829 , n6896 );
and ( n10101 , n10099 , n10100 );
xor ( n10102 , n10099 , n10100 );
xor ( n10103 , n10010 , n10019 );
and ( n10104 , n830 , n6896 );
and ( n10105 , n10103 , n10104 );
xor ( n10106 , n10103 , n10104 );
xor ( n10107 , n10014 , n10017 );
and ( n10108 , n831 , n6896 );
and ( n10109 , n10107 , n10108 );
and ( n10110 , n10106 , n10109 );
or ( n10111 , n10105 , n10110 );
and ( n10112 , n10102 , n10111 );
or ( n10113 , n10101 , n10112 );
and ( n10114 , n10098 , n10113 );
or ( n10115 , n10097 , n10114 );
and ( n10116 , n10094 , n10115 );
or ( n10117 , n10093 , n10116 );
and ( n10118 , n10090 , n10117 );
or ( n10119 , n10089 , n10118 );
and ( n10120 , n10086 , n10119 );
or ( n10121 , n10085 , n10120 );
and ( n10122 , n10082 , n10121 );
or ( n10123 , n10081 , n10122 );
and ( n10124 , n10078 , n10123 );
or ( n10125 , n10077 , n10124 );
and ( n10126 , n10074 , n10125 );
or ( n10127 , n10073 , n10126 );
and ( n10128 , n10070 , n10127 );
or ( n10129 , n10069 , n10128 );
and ( n10130 , n10066 , n10129 );
or ( n10131 , n10065 , n10130 );
and ( n10132 , n10062 , n10131 );
or ( n10133 , n10061 , n10132 );
and ( n10134 , n10058 , n10133 );
or ( n10135 , n10057 , n10134 );
and ( n10136 , n10054 , n10135 );
or ( n10137 , n10053 , n10136 );
and ( n10138 , n10050 , n10137 );
or ( n10139 , n10049 , n10138 );
and ( n10140 , n816 , n6893 );
and ( n10141 , n10139 , n10140 );
xor ( n10142 , n10139 , n10140 );
xor ( n10143 , n10050 , n10137 );
and ( n10144 , n817 , n6893 );
and ( n10145 , n10143 , n10144 );
xor ( n10146 , n10143 , n10144 );
xor ( n10147 , n10054 , n10135 );
and ( n10148 , n818 , n6893 );
and ( n10149 , n10147 , n10148 );
xor ( n10150 , n10147 , n10148 );
xor ( n10151 , n10058 , n10133 );
and ( n10152 , n819 , n6893 );
and ( n10153 , n10151 , n10152 );
xor ( n10154 , n10151 , n10152 );
xor ( n10155 , n10062 , n10131 );
and ( n10156 , n820 , n6893 );
and ( n10157 , n10155 , n10156 );
xor ( n10158 , n10155 , n10156 );
xor ( n10159 , n10066 , n10129 );
and ( n10160 , n821 , n6893 );
and ( n10161 , n10159 , n10160 );
xor ( n10162 , n10159 , n10160 );
xor ( n10163 , n10070 , n10127 );
and ( n10164 , n822 , n6893 );
and ( n10165 , n10163 , n10164 );
xor ( n10166 , n10163 , n10164 );
xor ( n10167 , n10074 , n10125 );
and ( n10168 , n823 , n6893 );
and ( n10169 , n10167 , n10168 );
xor ( n10170 , n10167 , n10168 );
xor ( n10171 , n10078 , n10123 );
and ( n10172 , n824 , n6893 );
and ( n10173 , n10171 , n10172 );
xor ( n10174 , n10171 , n10172 );
xor ( n10175 , n10082 , n10121 );
and ( n10176 , n825 , n6893 );
and ( n10177 , n10175 , n10176 );
xor ( n10178 , n10175 , n10176 );
xor ( n10179 , n10086 , n10119 );
and ( n10180 , n826 , n6893 );
and ( n10181 , n10179 , n10180 );
xor ( n10182 , n10179 , n10180 );
xor ( n10183 , n10090 , n10117 );
and ( n10184 , n827 , n6893 );
and ( n10185 , n10183 , n10184 );
xor ( n10186 , n10183 , n10184 );
xor ( n10187 , n10094 , n10115 );
and ( n10188 , n828 , n6893 );
and ( n10189 , n10187 , n10188 );
xor ( n10190 , n10187 , n10188 );
xor ( n10191 , n10098 , n10113 );
and ( n10192 , n829 , n6893 );
and ( n10193 , n10191 , n10192 );
xor ( n10194 , n10191 , n10192 );
xor ( n10195 , n10102 , n10111 );
and ( n10196 , n830 , n6893 );
and ( n10197 , n10195 , n10196 );
xor ( n10198 , n10195 , n10196 );
xor ( n10199 , n10106 , n10109 );
and ( n10200 , n831 , n6893 );
and ( n10201 , n10199 , n10200 );
and ( n10202 , n10198 , n10201 );
or ( n10203 , n10197 , n10202 );
and ( n10204 , n10194 , n10203 );
or ( n10205 , n10193 , n10204 );
and ( n10206 , n10190 , n10205 );
or ( n10207 , n10189 , n10206 );
and ( n10208 , n10186 , n10207 );
or ( n10209 , n10185 , n10208 );
and ( n10210 , n10182 , n10209 );
or ( n10211 , n10181 , n10210 );
and ( n10212 , n10178 , n10211 );
or ( n10213 , n10177 , n10212 );
and ( n10214 , n10174 , n10213 );
or ( n10215 , n10173 , n10214 );
and ( n10216 , n10170 , n10215 );
or ( n10217 , n10169 , n10216 );
and ( n10218 , n10166 , n10217 );
or ( n10219 , n10165 , n10218 );
and ( n10220 , n10162 , n10219 );
or ( n10221 , n10161 , n10220 );
and ( n10222 , n10158 , n10221 );
or ( n10223 , n10157 , n10222 );
and ( n10224 , n10154 , n10223 );
or ( n10225 , n10153 , n10224 );
and ( n10226 , n10150 , n10225 );
or ( n10227 , n10149 , n10226 );
and ( n10228 , n10146 , n10227 );
or ( n10229 , n10145 , n10228 );
and ( n10230 , n10142 , n10229 );
or ( n10231 , n10141 , n10230 );
and ( n10232 , n816 , n6890 );
and ( n10233 , n10231 , n10232 );
xor ( n10234 , n10231 , n10232 );
xor ( n10235 , n10142 , n10229 );
and ( n10236 , n817 , n6890 );
and ( n10237 , n10235 , n10236 );
xor ( n10238 , n10235 , n10236 );
xor ( n10239 , n10146 , n10227 );
and ( n10240 , n818 , n6890 );
and ( n10241 , n10239 , n10240 );
xor ( n10242 , n10239 , n10240 );
xor ( n10243 , n10150 , n10225 );
and ( n10244 , n819 , n6890 );
and ( n10245 , n10243 , n10244 );
xor ( n10246 , n10243 , n10244 );
xor ( n10247 , n10154 , n10223 );
and ( n10248 , n820 , n6890 );
and ( n10249 , n10247 , n10248 );
xor ( n10250 , n10247 , n10248 );
xor ( n10251 , n10158 , n10221 );
and ( n10252 , n821 , n6890 );
and ( n10253 , n10251 , n10252 );
xor ( n10254 , n10251 , n10252 );
xor ( n10255 , n10162 , n10219 );
and ( n10256 , n822 , n6890 );
and ( n10257 , n10255 , n10256 );
xor ( n10258 , n10255 , n10256 );
xor ( n10259 , n10166 , n10217 );
and ( n10260 , n823 , n6890 );
and ( n10261 , n10259 , n10260 );
xor ( n10262 , n10259 , n10260 );
xor ( n10263 , n10170 , n10215 );
and ( n10264 , n824 , n6890 );
and ( n10265 , n10263 , n10264 );
xor ( n10266 , n10263 , n10264 );
xor ( n10267 , n10174 , n10213 );
and ( n10268 , n825 , n6890 );
and ( n10269 , n10267 , n10268 );
xor ( n10270 , n10267 , n10268 );
xor ( n10271 , n10178 , n10211 );
and ( n10272 , n826 , n6890 );
and ( n10273 , n10271 , n10272 );
xor ( n10274 , n10271 , n10272 );
xor ( n10275 , n10182 , n10209 );
and ( n10276 , n827 , n6890 );
and ( n10277 , n10275 , n10276 );
xor ( n10278 , n10275 , n10276 );
xor ( n10279 , n10186 , n10207 );
and ( n10280 , n828 , n6890 );
and ( n10281 , n10279 , n10280 );
xor ( n10282 , n10279 , n10280 );
xor ( n10283 , n10190 , n10205 );
and ( n10284 , n829 , n6890 );
and ( n10285 , n10283 , n10284 );
xor ( n10286 , n10283 , n10284 );
xor ( n10287 , n10194 , n10203 );
and ( n10288 , n830 , n6890 );
and ( n10289 , n10287 , n10288 );
xor ( n10290 , n10287 , n10288 );
xor ( n10291 , n10198 , n10201 );
and ( n10292 , n831 , n6890 );
and ( n10293 , n10291 , n10292 );
and ( n10294 , n10290 , n10293 );
or ( n10295 , n10289 , n10294 );
and ( n10296 , n10286 , n10295 );
or ( n10297 , n10285 , n10296 );
and ( n10298 , n10282 , n10297 );
or ( n10299 , n10281 , n10298 );
and ( n10300 , n10278 , n10299 );
or ( n10301 , n10277 , n10300 );
and ( n10302 , n10274 , n10301 );
or ( n10303 , n10273 , n10302 );
and ( n10304 , n10270 , n10303 );
or ( n10305 , n10269 , n10304 );
and ( n10306 , n10266 , n10305 );
or ( n10307 , n10265 , n10306 );
and ( n10308 , n10262 , n10307 );
or ( n10309 , n10261 , n10308 );
and ( n10310 , n10258 , n10309 );
or ( n10311 , n10257 , n10310 );
and ( n10312 , n10254 , n10311 );
or ( n10313 , n10253 , n10312 );
and ( n10314 , n10250 , n10313 );
or ( n10315 , n10249 , n10314 );
and ( n10316 , n10246 , n10315 );
or ( n10317 , n10245 , n10316 );
and ( n10318 , n10242 , n10317 );
or ( n10319 , n10241 , n10318 );
and ( n10320 , n10238 , n10319 );
or ( n10321 , n10237 , n10320 );
and ( n10322 , n10234 , n10321 );
or ( n10323 , n10233 , n10322 );
and ( n10324 , n816 , n6887 );
and ( n10325 , n10323 , n10324 );
xor ( n10326 , n10323 , n10324 );
xor ( n10327 , n10234 , n10321 );
and ( n10328 , n817 , n6887 );
and ( n10329 , n10327 , n10328 );
xor ( n10330 , n10327 , n10328 );
xor ( n10331 , n10238 , n10319 );
and ( n10332 , n818 , n6887 );
and ( n10333 , n10331 , n10332 );
xor ( n10334 , n10331 , n10332 );
xor ( n10335 , n10242 , n10317 );
and ( n10336 , n819 , n6887 );
and ( n10337 , n10335 , n10336 );
xor ( n10338 , n10335 , n10336 );
xor ( n10339 , n10246 , n10315 );
and ( n10340 , n820 , n6887 );
and ( n10341 , n10339 , n10340 );
xor ( n10342 , n10339 , n10340 );
xor ( n10343 , n10250 , n10313 );
and ( n10344 , n821 , n6887 );
and ( n10345 , n10343 , n10344 );
xor ( n10346 , n10343 , n10344 );
xor ( n10347 , n10254 , n10311 );
and ( n10348 , n822 , n6887 );
and ( n10349 , n10347 , n10348 );
xor ( n10350 , n10347 , n10348 );
xor ( n10351 , n10258 , n10309 );
and ( n10352 , n823 , n6887 );
and ( n10353 , n10351 , n10352 );
xor ( n10354 , n10351 , n10352 );
xor ( n10355 , n10262 , n10307 );
and ( n10356 , n824 , n6887 );
and ( n10357 , n10355 , n10356 );
xor ( n10358 , n10355 , n10356 );
xor ( n10359 , n10266 , n10305 );
and ( n10360 , n825 , n6887 );
and ( n10361 , n10359 , n10360 );
xor ( n10362 , n10359 , n10360 );
xor ( n10363 , n10270 , n10303 );
and ( n10364 , n826 , n6887 );
and ( n10365 , n10363 , n10364 );
xor ( n10366 , n10363 , n10364 );
xor ( n10367 , n10274 , n10301 );
and ( n10368 , n827 , n6887 );
and ( n10369 , n10367 , n10368 );
xor ( n10370 , n10367 , n10368 );
xor ( n10371 , n10278 , n10299 );
and ( n10372 , n828 , n6887 );
and ( n10373 , n10371 , n10372 );
xor ( n10374 , n10371 , n10372 );
xor ( n10375 , n10282 , n10297 );
and ( n10376 , n829 , n6887 );
and ( n10377 , n10375 , n10376 );
xor ( n10378 , n10375 , n10376 );
xor ( n10379 , n10286 , n10295 );
and ( n10380 , n830 , n6887 );
and ( n10381 , n10379 , n10380 );
xor ( n10382 , n10379 , n10380 );
xor ( n10383 , n10290 , n10293 );
and ( n10384 , n831 , n6887 );
and ( n10385 , n10383 , n10384 );
and ( n10386 , n10382 , n10385 );
or ( n10387 , n10381 , n10386 );
and ( n10388 , n10378 , n10387 );
or ( n10389 , n10377 , n10388 );
and ( n10390 , n10374 , n10389 );
or ( n10391 , n10373 , n10390 );
and ( n10392 , n10370 , n10391 );
or ( n10393 , n10369 , n10392 );
and ( n10394 , n10366 , n10393 );
or ( n10395 , n10365 , n10394 );
and ( n10396 , n10362 , n10395 );
or ( n10397 , n10361 , n10396 );
and ( n10398 , n10358 , n10397 );
or ( n10399 , n10357 , n10398 );
and ( n10400 , n10354 , n10399 );
or ( n10401 , n10353 , n10400 );
and ( n10402 , n10350 , n10401 );
or ( n10403 , n10349 , n10402 );
and ( n10404 , n10346 , n10403 );
or ( n10405 , n10345 , n10404 );
and ( n10406 , n10342 , n10405 );
or ( n10407 , n10341 , n10406 );
and ( n10408 , n10338 , n10407 );
or ( n10409 , n10337 , n10408 );
and ( n10410 , n10334 , n10409 );
or ( n10411 , n10333 , n10410 );
and ( n10412 , n10330 , n10411 );
or ( n10413 , n10329 , n10412 );
and ( n10414 , n10326 , n10413 );
or ( n10415 , n10325 , n10414 );
and ( n10416 , n816 , n6884 );
and ( n10417 , n10415 , n10416 );
xor ( n10418 , n10415 , n10416 );
xor ( n10419 , n10326 , n10413 );
and ( n10420 , n817 , n6884 );
and ( n10421 , n10419 , n10420 );
xor ( n10422 , n10419 , n10420 );
xor ( n10423 , n10330 , n10411 );
and ( n10424 , n818 , n6884 );
and ( n10425 , n10423 , n10424 );
xor ( n10426 , n10423 , n10424 );
xor ( n10427 , n10334 , n10409 );
and ( n10428 , n819 , n6884 );
and ( n10429 , n10427 , n10428 );
xor ( n10430 , n10427 , n10428 );
xor ( n10431 , n10338 , n10407 );
and ( n10432 , n820 , n6884 );
and ( n10433 , n10431 , n10432 );
xor ( n10434 , n10431 , n10432 );
xor ( n10435 , n10342 , n10405 );
and ( n10436 , n821 , n6884 );
and ( n10437 , n10435 , n10436 );
xor ( n10438 , n10435 , n10436 );
xor ( n10439 , n10346 , n10403 );
and ( n10440 , n822 , n6884 );
and ( n10441 , n10439 , n10440 );
xor ( n10442 , n10439 , n10440 );
xor ( n10443 , n10350 , n10401 );
and ( n10444 , n823 , n6884 );
and ( n10445 , n10443 , n10444 );
xor ( n10446 , n10443 , n10444 );
xor ( n10447 , n10354 , n10399 );
and ( n10448 , n824 , n6884 );
and ( n10449 , n10447 , n10448 );
xor ( n10450 , n10447 , n10448 );
xor ( n10451 , n10358 , n10397 );
and ( n10452 , n825 , n6884 );
and ( n10453 , n10451 , n10452 );
xor ( n10454 , n10451 , n10452 );
xor ( n10455 , n10362 , n10395 );
and ( n10456 , n826 , n6884 );
and ( n10457 , n10455 , n10456 );
xor ( n10458 , n10455 , n10456 );
xor ( n10459 , n10366 , n10393 );
and ( n10460 , n827 , n6884 );
and ( n10461 , n10459 , n10460 );
xor ( n10462 , n10459 , n10460 );
xor ( n10463 , n10370 , n10391 );
and ( n10464 , n828 , n6884 );
and ( n10465 , n10463 , n10464 );
xor ( n10466 , n10463 , n10464 );
xor ( n10467 , n10374 , n10389 );
and ( n10468 , n829 , n6884 );
and ( n10469 , n10467 , n10468 );
xor ( n10470 , n10467 , n10468 );
xor ( n10471 , n10378 , n10387 );
and ( n10472 , n830 , n6884 );
and ( n10473 , n10471 , n10472 );
xor ( n10474 , n10471 , n10472 );
xor ( n10475 , n10382 , n10385 );
and ( n10476 , n831 , n6884 );
and ( n10477 , n10475 , n10476 );
and ( n10478 , n10474 , n10477 );
or ( n10479 , n10473 , n10478 );
and ( n10480 , n10470 , n10479 );
or ( n10481 , n10469 , n10480 );
and ( n10482 , n10466 , n10481 );
or ( n10483 , n10465 , n10482 );
and ( n10484 , n10462 , n10483 );
or ( n10485 , n10461 , n10484 );
and ( n10486 , n10458 , n10485 );
or ( n10487 , n10457 , n10486 );
and ( n10488 , n10454 , n10487 );
or ( n10489 , n10453 , n10488 );
and ( n10490 , n10450 , n10489 );
or ( n10491 , n10449 , n10490 );
and ( n10492 , n10446 , n10491 );
or ( n10493 , n10445 , n10492 );
and ( n10494 , n10442 , n10493 );
or ( n10495 , n10441 , n10494 );
and ( n10496 , n10438 , n10495 );
or ( n10497 , n10437 , n10496 );
and ( n10498 , n10434 , n10497 );
or ( n10499 , n10433 , n10498 );
and ( n10500 , n10430 , n10499 );
or ( n10501 , n10429 , n10500 );
and ( n10502 , n10426 , n10501 );
or ( n10503 , n10425 , n10502 );
and ( n10504 , n10422 , n10503 );
or ( n10505 , n10421 , n10504 );
and ( n10506 , n10418 , n10505 );
or ( n10507 , n10417 , n10506 );
and ( n10508 , n816 , n6881 );
and ( n10509 , n10507 , n10508 );
xor ( n10510 , n10507 , n10508 );
xor ( n10511 , n10418 , n10505 );
and ( n10512 , n817 , n6881 );
and ( n10513 , n10511 , n10512 );
xor ( n10514 , n10511 , n10512 );
xor ( n10515 , n10422 , n10503 );
and ( n10516 , n818 , n6881 );
and ( n10517 , n10515 , n10516 );
xor ( n10518 , n10515 , n10516 );
xor ( n10519 , n10426 , n10501 );
and ( n10520 , n819 , n6881 );
and ( n10521 , n10519 , n10520 );
xor ( n10522 , n10519 , n10520 );
xor ( n10523 , n10430 , n10499 );
and ( n10524 , n820 , n6881 );
and ( n10525 , n10523 , n10524 );
xor ( n10526 , n10523 , n10524 );
xor ( n10527 , n10434 , n10497 );
and ( n10528 , n821 , n6881 );
and ( n10529 , n10527 , n10528 );
xor ( n10530 , n10527 , n10528 );
xor ( n10531 , n10438 , n10495 );
and ( n10532 , n822 , n6881 );
and ( n10533 , n10531 , n10532 );
xor ( n10534 , n10531 , n10532 );
xor ( n10535 , n10442 , n10493 );
and ( n10536 , n823 , n6881 );
and ( n10537 , n10535 , n10536 );
xor ( n10538 , n10535 , n10536 );
xor ( n10539 , n10446 , n10491 );
and ( n10540 , n824 , n6881 );
and ( n10541 , n10539 , n10540 );
xor ( n10542 , n10539 , n10540 );
xor ( n10543 , n10450 , n10489 );
and ( n10544 , n825 , n6881 );
and ( n10545 , n10543 , n10544 );
xor ( n10546 , n10543 , n10544 );
xor ( n10547 , n10454 , n10487 );
and ( n10548 , n826 , n6881 );
and ( n10549 , n10547 , n10548 );
xor ( n10550 , n10547 , n10548 );
xor ( n10551 , n10458 , n10485 );
and ( n10552 , n827 , n6881 );
and ( n10553 , n10551 , n10552 );
xor ( n10554 , n10551 , n10552 );
xor ( n10555 , n10462 , n10483 );
and ( n10556 , n828 , n6881 );
and ( n10557 , n10555 , n10556 );
xor ( n10558 , n10555 , n10556 );
xor ( n10559 , n10466 , n10481 );
and ( n10560 , n829 , n6881 );
and ( n10561 , n10559 , n10560 );
xor ( n10562 , n10559 , n10560 );
xor ( n10563 , n10470 , n10479 );
and ( n10564 , n830 , n6881 );
and ( n10565 , n10563 , n10564 );
xor ( n10566 , n10563 , n10564 );
xor ( n10567 , n10474 , n10477 );
and ( n10568 , n831 , n6881 );
and ( n10569 , n10567 , n10568 );
and ( n10570 , n10566 , n10569 );
or ( n10571 , n10565 , n10570 );
and ( n10572 , n10562 , n10571 );
or ( n10573 , n10561 , n10572 );
and ( n10574 , n10558 , n10573 );
or ( n10575 , n10557 , n10574 );
and ( n10576 , n10554 , n10575 );
or ( n10577 , n10553 , n10576 );
and ( n10578 , n10550 , n10577 );
or ( n10579 , n10549 , n10578 );
and ( n10580 , n10546 , n10579 );
or ( n10581 , n10545 , n10580 );
and ( n10582 , n10542 , n10581 );
or ( n10583 , n10541 , n10582 );
and ( n10584 , n10538 , n10583 );
or ( n10585 , n10537 , n10584 );
and ( n10586 , n10534 , n10585 );
or ( n10587 , n10533 , n10586 );
and ( n10588 , n10530 , n10587 );
or ( n10589 , n10529 , n10588 );
and ( n10590 , n10526 , n10589 );
or ( n10591 , n10525 , n10590 );
and ( n10592 , n10522 , n10591 );
or ( n10593 , n10521 , n10592 );
and ( n10594 , n10518 , n10593 );
or ( n10595 , n10517 , n10594 );
and ( n10596 , n10514 , n10595 );
or ( n10597 , n10513 , n10596 );
and ( n10598 , n10510 , n10597 );
or ( n10599 , n10509 , n10598 );
and ( n10600 , n816 , n6878 );
and ( n10601 , n10599 , n10600 );
xor ( n10602 , n10599 , n10600 );
xor ( n10603 , n10510 , n10597 );
and ( n10604 , n817 , n6878 );
and ( n10605 , n10603 , n10604 );
xor ( n10606 , n10603 , n10604 );
xor ( n10607 , n10514 , n10595 );
and ( n10608 , n818 , n6878 );
and ( n10609 , n10607 , n10608 );
xor ( n10610 , n10607 , n10608 );
xor ( n10611 , n10518 , n10593 );
and ( n10612 , n819 , n6878 );
and ( n10613 , n10611 , n10612 );
xor ( n10614 , n10611 , n10612 );
xor ( n10615 , n10522 , n10591 );
and ( n10616 , n820 , n6878 );
and ( n10617 , n10615 , n10616 );
xor ( n10618 , n10615 , n10616 );
xor ( n10619 , n10526 , n10589 );
and ( n10620 , n821 , n6878 );
and ( n10621 , n10619 , n10620 );
xor ( n10622 , n10619 , n10620 );
xor ( n10623 , n10530 , n10587 );
and ( n10624 , n822 , n6878 );
and ( n10625 , n10623 , n10624 );
xor ( n10626 , n10623 , n10624 );
xor ( n10627 , n10534 , n10585 );
and ( n10628 , n823 , n6878 );
and ( n10629 , n10627 , n10628 );
xor ( n10630 , n10627 , n10628 );
xor ( n10631 , n10538 , n10583 );
and ( n10632 , n824 , n6878 );
and ( n10633 , n10631 , n10632 );
xor ( n10634 , n10631 , n10632 );
xor ( n10635 , n10542 , n10581 );
and ( n10636 , n825 , n6878 );
and ( n10637 , n10635 , n10636 );
xor ( n10638 , n10635 , n10636 );
xor ( n10639 , n10546 , n10579 );
and ( n10640 , n826 , n6878 );
and ( n10641 , n10639 , n10640 );
xor ( n10642 , n10639 , n10640 );
xor ( n10643 , n10550 , n10577 );
and ( n10644 , n827 , n6878 );
and ( n10645 , n10643 , n10644 );
xor ( n10646 , n10643 , n10644 );
xor ( n10647 , n10554 , n10575 );
and ( n10648 , n828 , n6878 );
and ( n10649 , n10647 , n10648 );
xor ( n10650 , n10647 , n10648 );
xor ( n10651 , n10558 , n10573 );
and ( n10652 , n829 , n6878 );
and ( n10653 , n10651 , n10652 );
xor ( n10654 , n10651 , n10652 );
xor ( n10655 , n10562 , n10571 );
and ( n10656 , n830 , n6878 );
and ( n10657 , n10655 , n10656 );
xor ( n10658 , n10655 , n10656 );
xor ( n10659 , n10566 , n10569 );
and ( n10660 , n831 , n6878 );
and ( n10661 , n10659 , n10660 );
and ( n10662 , n10658 , n10661 );
or ( n10663 , n10657 , n10662 );
and ( n10664 , n10654 , n10663 );
or ( n10665 , n10653 , n10664 );
and ( n10666 , n10650 , n10665 );
or ( n10667 , n10649 , n10666 );
and ( n10668 , n10646 , n10667 );
or ( n10669 , n10645 , n10668 );
and ( n10670 , n10642 , n10669 );
or ( n10671 , n10641 , n10670 );
and ( n10672 , n10638 , n10671 );
or ( n10673 , n10637 , n10672 );
and ( n10674 , n10634 , n10673 );
or ( n10675 , n10633 , n10674 );
and ( n10676 , n10630 , n10675 );
or ( n10677 , n10629 , n10676 );
and ( n10678 , n10626 , n10677 );
or ( n10679 , n10625 , n10678 );
and ( n10680 , n10622 , n10679 );
or ( n10681 , n10621 , n10680 );
and ( n10682 , n10618 , n10681 );
or ( n10683 , n10617 , n10682 );
and ( n10684 , n10614 , n10683 );
or ( n10685 , n10613 , n10684 );
and ( n10686 , n10610 , n10685 );
or ( n10687 , n10609 , n10686 );
and ( n10688 , n10606 , n10687 );
or ( n10689 , n10605 , n10688 );
and ( n10690 , n10602 , n10689 );
or ( n10691 , n10601 , n10690 );
and ( n10692 , n816 , n6875 );
and ( n10693 , n10691 , n10692 );
xor ( n10694 , n10691 , n10692 );
xor ( n10695 , n10602 , n10689 );
and ( n10696 , n817 , n6875 );
and ( n10697 , n10695 , n10696 );
xor ( n10698 , n10695 , n10696 );
xor ( n10699 , n10606 , n10687 );
and ( n10700 , n818 , n6875 );
and ( n10701 , n10699 , n10700 );
xor ( n10702 , n10699 , n10700 );
xor ( n10703 , n10610 , n10685 );
and ( n10704 , n819 , n6875 );
and ( n10705 , n10703 , n10704 );
xor ( n10706 , n10703 , n10704 );
xor ( n10707 , n10614 , n10683 );
and ( n10708 , n820 , n6875 );
and ( n10709 , n10707 , n10708 );
xor ( n10710 , n10707 , n10708 );
xor ( n10711 , n10618 , n10681 );
and ( n10712 , n821 , n6875 );
and ( n10713 , n10711 , n10712 );
xor ( n10714 , n10711 , n10712 );
xor ( n10715 , n10622 , n10679 );
and ( n10716 , n822 , n6875 );
and ( n10717 , n10715 , n10716 );
xor ( n10718 , n10715 , n10716 );
xor ( n10719 , n10626 , n10677 );
and ( n10720 , n823 , n6875 );
and ( n10721 , n10719 , n10720 );
xor ( n10722 , n10719 , n10720 );
xor ( n10723 , n10630 , n10675 );
and ( n10724 , n824 , n6875 );
and ( n10725 , n10723 , n10724 );
xor ( n10726 , n10723 , n10724 );
xor ( n10727 , n10634 , n10673 );
and ( n10728 , n825 , n6875 );
and ( n10729 , n10727 , n10728 );
xor ( n10730 , n10727 , n10728 );
xor ( n10731 , n10638 , n10671 );
and ( n10732 , n826 , n6875 );
and ( n10733 , n10731 , n10732 );
xor ( n10734 , n10731 , n10732 );
xor ( n10735 , n10642 , n10669 );
and ( n10736 , n827 , n6875 );
and ( n10737 , n10735 , n10736 );
xor ( n10738 , n10735 , n10736 );
xor ( n10739 , n10646 , n10667 );
and ( n10740 , n828 , n6875 );
and ( n10741 , n10739 , n10740 );
xor ( n10742 , n10739 , n10740 );
xor ( n10743 , n10650 , n10665 );
and ( n10744 , n829 , n6875 );
and ( n10745 , n10743 , n10744 );
xor ( n10746 , n10743 , n10744 );
xor ( n10747 , n10654 , n10663 );
and ( n10748 , n830 , n6875 );
and ( n10749 , n10747 , n10748 );
xor ( n10750 , n10747 , n10748 );
xor ( n10751 , n10658 , n10661 );
and ( n10752 , n831 , n6875 );
and ( n10753 , n10751 , n10752 );
and ( n10754 , n10750 , n10753 );
or ( n10755 , n10749 , n10754 );
and ( n10756 , n10746 , n10755 );
or ( n10757 , n10745 , n10756 );
and ( n10758 , n10742 , n10757 );
or ( n10759 , n10741 , n10758 );
and ( n10760 , n10738 , n10759 );
or ( n10761 , n10737 , n10760 );
and ( n10762 , n10734 , n10761 );
or ( n10763 , n10733 , n10762 );
and ( n10764 , n10730 , n10763 );
or ( n10765 , n10729 , n10764 );
and ( n10766 , n10726 , n10765 );
or ( n10767 , n10725 , n10766 );
and ( n10768 , n10722 , n10767 );
or ( n10769 , n10721 , n10768 );
and ( n10770 , n10718 , n10769 );
or ( n10771 , n10717 , n10770 );
and ( n10772 , n10714 , n10771 );
or ( n10773 , n10713 , n10772 );
and ( n10774 , n10710 , n10773 );
or ( n10775 , n10709 , n10774 );
and ( n10776 , n10706 , n10775 );
or ( n10777 , n10705 , n10776 );
and ( n10778 , n10702 , n10777 );
or ( n10779 , n10701 , n10778 );
and ( n10780 , n10698 , n10779 );
or ( n10781 , n10697 , n10780 );
and ( n10782 , n10694 , n10781 );
or ( n10783 , n10693 , n10782 );
and ( n10784 , n816 , n6872 );
and ( n10785 , n10783 , n10784 );
xor ( n10786 , n10783 , n10784 );
xor ( n10787 , n10694 , n10781 );
and ( n10788 , n817 , n6872 );
and ( n10789 , n10787 , n10788 );
xor ( n10790 , n10787 , n10788 );
xor ( n10791 , n10698 , n10779 );
and ( n10792 , n818 , n6872 );
and ( n10793 , n10791 , n10792 );
xor ( n10794 , n10791 , n10792 );
xor ( n10795 , n10702 , n10777 );
and ( n10796 , n819 , n6872 );
and ( n10797 , n10795 , n10796 );
xor ( n10798 , n10795 , n10796 );
xor ( n10799 , n10706 , n10775 );
and ( n10800 , n820 , n6872 );
and ( n10801 , n10799 , n10800 );
xor ( n10802 , n10799 , n10800 );
xor ( n10803 , n10710 , n10773 );
and ( n10804 , n821 , n6872 );
and ( n10805 , n10803 , n10804 );
xor ( n10806 , n10803 , n10804 );
xor ( n10807 , n10714 , n10771 );
and ( n10808 , n822 , n6872 );
and ( n10809 , n10807 , n10808 );
xor ( n10810 , n10807 , n10808 );
xor ( n10811 , n10718 , n10769 );
and ( n10812 , n823 , n6872 );
and ( n10813 , n10811 , n10812 );
xor ( n10814 , n10811 , n10812 );
xor ( n10815 , n10722 , n10767 );
and ( n10816 , n824 , n6872 );
and ( n10817 , n10815 , n10816 );
xor ( n10818 , n10815 , n10816 );
xor ( n10819 , n10726 , n10765 );
and ( n10820 , n825 , n6872 );
and ( n10821 , n10819 , n10820 );
xor ( n10822 , n10819 , n10820 );
xor ( n10823 , n10730 , n10763 );
and ( n10824 , n826 , n6872 );
and ( n10825 , n10823 , n10824 );
xor ( n10826 , n10823 , n10824 );
xor ( n10827 , n10734 , n10761 );
and ( n10828 , n827 , n6872 );
and ( n10829 , n10827 , n10828 );
xor ( n10830 , n10827 , n10828 );
xor ( n10831 , n10738 , n10759 );
and ( n10832 , n828 , n6872 );
and ( n10833 , n10831 , n10832 );
xor ( n10834 , n10831 , n10832 );
xor ( n10835 , n10742 , n10757 );
and ( n10836 , n829 , n6872 );
and ( n10837 , n10835 , n10836 );
xor ( n10838 , n10835 , n10836 );
xor ( n10839 , n10746 , n10755 );
and ( n10840 , n830 , n6872 );
and ( n10841 , n10839 , n10840 );
xor ( n10842 , n10839 , n10840 );
xor ( n10843 , n10750 , n10753 );
and ( n10844 , n831 , n6872 );
and ( n10845 , n10843 , n10844 );
and ( n10846 , n10842 , n10845 );
or ( n10847 , n10841 , n10846 );
and ( n10848 , n10838 , n10847 );
or ( n10849 , n10837 , n10848 );
and ( n10850 , n10834 , n10849 );
or ( n10851 , n10833 , n10850 );
and ( n10852 , n10830 , n10851 );
or ( n10853 , n10829 , n10852 );
and ( n10854 , n10826 , n10853 );
or ( n10855 , n10825 , n10854 );
and ( n10856 , n10822 , n10855 );
or ( n10857 , n10821 , n10856 );
and ( n10858 , n10818 , n10857 );
or ( n10859 , n10817 , n10858 );
and ( n10860 , n10814 , n10859 );
or ( n10861 , n10813 , n10860 );
and ( n10862 , n10810 , n10861 );
or ( n10863 , n10809 , n10862 );
and ( n10864 , n10806 , n10863 );
or ( n10865 , n10805 , n10864 );
and ( n10866 , n10802 , n10865 );
or ( n10867 , n10801 , n10866 );
and ( n10868 , n10798 , n10867 );
or ( n10869 , n10797 , n10868 );
and ( n10870 , n10794 , n10869 );
or ( n10871 , n10793 , n10870 );
and ( n10872 , n10790 , n10871 );
or ( n10873 , n10789 , n10872 );
and ( n10874 , n10786 , n10873 );
or ( n10875 , n10785 , n10874 );
and ( n10876 , n816 , n6869 );
and ( n10877 , n10875 , n10876 );
xor ( n10878 , n10875 , n10876 );
xor ( n10879 , n10786 , n10873 );
and ( n10880 , n817 , n6869 );
and ( n10881 , n10879 , n10880 );
xor ( n10882 , n10879 , n10880 );
xor ( n10883 , n10790 , n10871 );
and ( n10884 , n818 , n6869 );
and ( n10885 , n10883 , n10884 );
xor ( n10886 , n10883 , n10884 );
xor ( n10887 , n10794 , n10869 );
and ( n10888 , n819 , n6869 );
and ( n10889 , n10887 , n10888 );
xor ( n10890 , n10887 , n10888 );
xor ( n10891 , n10798 , n10867 );
and ( n10892 , n820 , n6869 );
and ( n10893 , n10891 , n10892 );
xor ( n10894 , n10891 , n10892 );
xor ( n10895 , n10802 , n10865 );
and ( n10896 , n821 , n6869 );
and ( n10897 , n10895 , n10896 );
xor ( n10898 , n10895 , n10896 );
xor ( n10899 , n10806 , n10863 );
and ( n10900 , n822 , n6869 );
and ( n10901 , n10899 , n10900 );
xor ( n10902 , n10899 , n10900 );
xor ( n10903 , n10810 , n10861 );
and ( n10904 , n823 , n6869 );
and ( n10905 , n10903 , n10904 );
xor ( n10906 , n10903 , n10904 );
xor ( n10907 , n10814 , n10859 );
and ( n10908 , n824 , n6869 );
and ( n10909 , n10907 , n10908 );
xor ( n10910 , n10907 , n10908 );
xor ( n10911 , n10818 , n10857 );
and ( n10912 , n825 , n6869 );
and ( n10913 , n10911 , n10912 );
xor ( n10914 , n10911 , n10912 );
xor ( n10915 , n10822 , n10855 );
and ( n10916 , n826 , n6869 );
and ( n10917 , n10915 , n10916 );
xor ( n10918 , n10915 , n10916 );
xor ( n10919 , n10826 , n10853 );
and ( n10920 , n827 , n6869 );
and ( n10921 , n10919 , n10920 );
xor ( n10922 , n10919 , n10920 );
xor ( n10923 , n10830 , n10851 );
and ( n10924 , n828 , n6869 );
and ( n10925 , n10923 , n10924 );
xor ( n10926 , n10923 , n10924 );
xor ( n10927 , n10834 , n10849 );
and ( n10928 , n829 , n6869 );
and ( n10929 , n10927 , n10928 );
xor ( n10930 , n10927 , n10928 );
xor ( n10931 , n10838 , n10847 );
and ( n10932 , n830 , n6869 );
and ( n10933 , n10931 , n10932 );
xor ( n10934 , n10931 , n10932 );
xor ( n10935 , n10842 , n10845 );
and ( n10936 , n831 , n6869 );
and ( n10937 , n10935 , n10936 );
and ( n10938 , n10934 , n10937 );
or ( n10939 , n10933 , n10938 );
and ( n10940 , n10930 , n10939 );
or ( n10941 , n10929 , n10940 );
and ( n10942 , n10926 , n10941 );
or ( n10943 , n10925 , n10942 );
and ( n10944 , n10922 , n10943 );
or ( n10945 , n10921 , n10944 );
and ( n10946 , n10918 , n10945 );
or ( n10947 , n10917 , n10946 );
and ( n10948 , n10914 , n10947 );
or ( n10949 , n10913 , n10948 );
and ( n10950 , n10910 , n10949 );
or ( n10951 , n10909 , n10950 );
and ( n10952 , n10906 , n10951 );
or ( n10953 , n10905 , n10952 );
and ( n10954 , n10902 , n10953 );
or ( n10955 , n10901 , n10954 );
and ( n10956 , n10898 , n10955 );
or ( n10957 , n10897 , n10956 );
and ( n10958 , n10894 , n10957 );
or ( n10959 , n10893 , n10958 );
and ( n10960 , n10890 , n10959 );
or ( n10961 , n10889 , n10960 );
and ( n10962 , n10886 , n10961 );
or ( n10963 , n10885 , n10962 );
and ( n10964 , n10882 , n10963 );
or ( n10965 , n10881 , n10964 );
and ( n10966 , n10878 , n10965 );
or ( n10967 , n10877 , n10966 );
and ( n10968 , n816 , n6866 );
and ( n10969 , n10967 , n10968 );
xor ( n10970 , n10967 , n10968 );
xor ( n10971 , n10878 , n10965 );
and ( n10972 , n817 , n6866 );
and ( n10973 , n10971 , n10972 );
xor ( n10974 , n10971 , n10972 );
xor ( n10975 , n10882 , n10963 );
and ( n10976 , n818 , n6866 );
and ( n10977 , n10975 , n10976 );
xor ( n10978 , n10975 , n10976 );
xor ( n10979 , n10886 , n10961 );
and ( n10980 , n819 , n6866 );
and ( n10981 , n10979 , n10980 );
xor ( n10982 , n10979 , n10980 );
xor ( n10983 , n10890 , n10959 );
and ( n10984 , n820 , n6866 );
and ( n10985 , n10983 , n10984 );
xor ( n10986 , n10983 , n10984 );
xor ( n10987 , n10894 , n10957 );
and ( n10988 , n821 , n6866 );
and ( n10989 , n10987 , n10988 );
xor ( n10990 , n10987 , n10988 );
xor ( n10991 , n10898 , n10955 );
and ( n10992 , n822 , n6866 );
and ( n10993 , n10991 , n10992 );
xor ( n10994 , n10991 , n10992 );
xor ( n10995 , n10902 , n10953 );
and ( n10996 , n823 , n6866 );
and ( n10997 , n10995 , n10996 );
xor ( n10998 , n10995 , n10996 );
xor ( n10999 , n10906 , n10951 );
and ( n11000 , n824 , n6866 );
and ( n11001 , n10999 , n11000 );
xor ( n11002 , n10999 , n11000 );
xor ( n11003 , n10910 , n10949 );
and ( n11004 , n825 , n6866 );
and ( n11005 , n11003 , n11004 );
xor ( n11006 , n11003 , n11004 );
xor ( n11007 , n10914 , n10947 );
and ( n11008 , n826 , n6866 );
and ( n11009 , n11007 , n11008 );
xor ( n11010 , n11007 , n11008 );
xor ( n11011 , n10918 , n10945 );
and ( n11012 , n827 , n6866 );
and ( n11013 , n11011 , n11012 );
xor ( n11014 , n11011 , n11012 );
xor ( n11015 , n10922 , n10943 );
and ( n11016 , n828 , n6866 );
and ( n11017 , n11015 , n11016 );
xor ( n11018 , n11015 , n11016 );
xor ( n11019 , n10926 , n10941 );
and ( n11020 , n829 , n6866 );
and ( n11021 , n11019 , n11020 );
xor ( n11022 , n11019 , n11020 );
xor ( n11023 , n10930 , n10939 );
and ( n11024 , n830 , n6866 );
and ( n11025 , n11023 , n11024 );
xor ( n11026 , n11023 , n11024 );
xor ( n11027 , n10934 , n10937 );
and ( n11028 , n831 , n6866 );
and ( n11029 , n11027 , n11028 );
and ( n11030 , n11026 , n11029 );
or ( n11031 , n11025 , n11030 );
and ( n11032 , n11022 , n11031 );
or ( n11033 , n11021 , n11032 );
and ( n11034 , n11018 , n11033 );
or ( n11035 , n11017 , n11034 );
and ( n11036 , n11014 , n11035 );
or ( n11037 , n11013 , n11036 );
and ( n11038 , n11010 , n11037 );
or ( n11039 , n11009 , n11038 );
and ( n11040 , n11006 , n11039 );
or ( n11041 , n11005 , n11040 );
and ( n11042 , n11002 , n11041 );
or ( n11043 , n11001 , n11042 );
and ( n11044 , n10998 , n11043 );
or ( n11045 , n10997 , n11044 );
and ( n11046 , n10994 , n11045 );
or ( n11047 , n10993 , n11046 );
and ( n11048 , n10990 , n11047 );
or ( n11049 , n10989 , n11048 );
and ( n11050 , n10986 , n11049 );
or ( n11051 , n10985 , n11050 );
and ( n11052 , n10982 , n11051 );
or ( n11053 , n10981 , n11052 );
and ( n11054 , n10978 , n11053 );
or ( n11055 , n10977 , n11054 );
and ( n11056 , n10974 , n11055 );
or ( n11057 , n10973 , n11056 );
and ( n11058 , n10970 , n11057 );
or ( n11059 , n10969 , n11058 );
and ( n11060 , n816 , n6863 );
and ( n11061 , n11059 , n11060 );
xor ( n11062 , n11059 , n11060 );
xor ( n11063 , n10970 , n11057 );
and ( n11064 , n817 , n6863 );
and ( n11065 , n11063 , n11064 );
xor ( n11066 , n11063 , n11064 );
xor ( n11067 , n10974 , n11055 );
and ( n11068 , n818 , n6863 );
and ( n11069 , n11067 , n11068 );
xor ( n11070 , n11067 , n11068 );
xor ( n11071 , n10978 , n11053 );
and ( n11072 , n819 , n6863 );
and ( n11073 , n11071 , n11072 );
xor ( n11074 , n11071 , n11072 );
xor ( n11075 , n10982 , n11051 );
and ( n11076 , n820 , n6863 );
and ( n11077 , n11075 , n11076 );
xor ( n11078 , n11075 , n11076 );
xor ( n11079 , n10986 , n11049 );
and ( n11080 , n821 , n6863 );
and ( n11081 , n11079 , n11080 );
xor ( n11082 , n11079 , n11080 );
xor ( n11083 , n10990 , n11047 );
and ( n11084 , n822 , n6863 );
and ( n11085 , n11083 , n11084 );
xor ( n11086 , n11083 , n11084 );
xor ( n11087 , n10994 , n11045 );
and ( n11088 , n823 , n6863 );
and ( n11089 , n11087 , n11088 );
xor ( n11090 , n11087 , n11088 );
xor ( n11091 , n10998 , n11043 );
and ( n11092 , n824 , n6863 );
and ( n11093 , n11091 , n11092 );
xor ( n11094 , n11091 , n11092 );
xor ( n11095 , n11002 , n11041 );
and ( n11096 , n825 , n6863 );
and ( n11097 , n11095 , n11096 );
xor ( n11098 , n11095 , n11096 );
xor ( n11099 , n11006 , n11039 );
and ( n11100 , n826 , n6863 );
and ( n11101 , n11099 , n11100 );
xor ( n11102 , n11099 , n11100 );
xor ( n11103 , n11010 , n11037 );
and ( n11104 , n827 , n6863 );
and ( n11105 , n11103 , n11104 );
xor ( n11106 , n11103 , n11104 );
xor ( n11107 , n11014 , n11035 );
and ( n11108 , n828 , n6863 );
and ( n11109 , n11107 , n11108 );
xor ( n11110 , n11107 , n11108 );
xor ( n11111 , n11018 , n11033 );
and ( n11112 , n829 , n6863 );
and ( n11113 , n11111 , n11112 );
xor ( n11114 , n11111 , n11112 );
xor ( n11115 , n11022 , n11031 );
and ( n11116 , n830 , n6863 );
and ( n11117 , n11115 , n11116 );
xor ( n11118 , n11115 , n11116 );
xor ( n11119 , n11026 , n11029 );
and ( n11120 , n831 , n6863 );
and ( n11121 , n11119 , n11120 );
and ( n11122 , n11118 , n11121 );
or ( n11123 , n11117 , n11122 );
and ( n11124 , n11114 , n11123 );
or ( n11125 , n11113 , n11124 );
and ( n11126 , n11110 , n11125 );
or ( n11127 , n11109 , n11126 );
and ( n11128 , n11106 , n11127 );
or ( n11129 , n11105 , n11128 );
and ( n11130 , n11102 , n11129 );
or ( n11131 , n11101 , n11130 );
and ( n11132 , n11098 , n11131 );
or ( n11133 , n11097 , n11132 );
and ( n11134 , n11094 , n11133 );
or ( n11135 , n11093 , n11134 );
and ( n11136 , n11090 , n11135 );
or ( n11137 , n11089 , n11136 );
and ( n11138 , n11086 , n11137 );
or ( n11139 , n11085 , n11138 );
and ( n11140 , n11082 , n11139 );
or ( n11141 , n11081 , n11140 );
and ( n11142 , n11078 , n11141 );
or ( n11143 , n11077 , n11142 );
and ( n11144 , n11074 , n11143 );
or ( n11145 , n11073 , n11144 );
and ( n11146 , n11070 , n11145 );
or ( n11147 , n11069 , n11146 );
and ( n11148 , n11066 , n11147 );
or ( n11149 , n11065 , n11148 );
and ( n11150 , n11062 , n11149 );
or ( n11151 , n11061 , n11150 );
and ( n11152 , n816 , n6860 );
and ( n11153 , n11151 , n11152 );
xor ( n11154 , n11151 , n11152 );
xor ( n11155 , n11062 , n11149 );
and ( n11156 , n817 , n6860 );
and ( n11157 , n11155 , n11156 );
xor ( n11158 , n11155 , n11156 );
xor ( n11159 , n11066 , n11147 );
and ( n11160 , n818 , n6860 );
and ( n11161 , n11159 , n11160 );
xor ( n11162 , n11159 , n11160 );
xor ( n11163 , n11070 , n11145 );
and ( n11164 , n819 , n6860 );
and ( n11165 , n11163 , n11164 );
xor ( n11166 , n11163 , n11164 );
xor ( n11167 , n11074 , n11143 );
and ( n11168 , n820 , n6860 );
and ( n11169 , n11167 , n11168 );
xor ( n11170 , n11167 , n11168 );
xor ( n11171 , n11078 , n11141 );
and ( n11172 , n821 , n6860 );
and ( n11173 , n11171 , n11172 );
xor ( n11174 , n11171 , n11172 );
xor ( n11175 , n11082 , n11139 );
and ( n11176 , n822 , n6860 );
and ( n11177 , n11175 , n11176 );
xor ( n11178 , n11175 , n11176 );
xor ( n11179 , n11086 , n11137 );
and ( n11180 , n823 , n6860 );
and ( n11181 , n11179 , n11180 );
xor ( n11182 , n11179 , n11180 );
xor ( n11183 , n11090 , n11135 );
and ( n11184 , n824 , n6860 );
and ( n11185 , n11183 , n11184 );
xor ( n11186 , n11183 , n11184 );
xor ( n11187 , n11094 , n11133 );
and ( n11188 , n825 , n6860 );
and ( n11189 , n11187 , n11188 );
xor ( n11190 , n11187 , n11188 );
xor ( n11191 , n11098 , n11131 );
and ( n11192 , n826 , n6860 );
and ( n11193 , n11191 , n11192 );
xor ( n11194 , n11191 , n11192 );
xor ( n11195 , n11102 , n11129 );
and ( n11196 , n827 , n6860 );
and ( n11197 , n11195 , n11196 );
xor ( n11198 , n11195 , n11196 );
xor ( n11199 , n11106 , n11127 );
and ( n11200 , n828 , n6860 );
and ( n11201 , n11199 , n11200 );
xor ( n11202 , n11199 , n11200 );
xor ( n11203 , n11110 , n11125 );
and ( n11204 , n829 , n6860 );
and ( n11205 , n11203 , n11204 );
xor ( n11206 , n11203 , n11204 );
xor ( n11207 , n11114 , n11123 );
and ( n11208 , n830 , n6860 );
and ( n11209 , n11207 , n11208 );
xor ( n11210 , n11207 , n11208 );
xor ( n11211 , n11118 , n11121 );
and ( n11212 , n831 , n6860 );
and ( n11213 , n11211 , n11212 );
and ( n11214 , n11210 , n11213 );
or ( n11215 , n11209 , n11214 );
and ( n11216 , n11206 , n11215 );
or ( n11217 , n11205 , n11216 );
and ( n11218 , n11202 , n11217 );
or ( n11219 , n11201 , n11218 );
and ( n11220 , n11198 , n11219 );
or ( n11221 , n11197 , n11220 );
and ( n11222 , n11194 , n11221 );
or ( n11223 , n11193 , n11222 );
and ( n11224 , n11190 , n11223 );
or ( n11225 , n11189 , n11224 );
and ( n11226 , n11186 , n11225 );
or ( n11227 , n11185 , n11226 );
and ( n11228 , n11182 , n11227 );
or ( n11229 , n11181 , n11228 );
and ( n11230 , n11178 , n11229 );
or ( n11231 , n11177 , n11230 );
and ( n11232 , n11174 , n11231 );
or ( n11233 , n11173 , n11232 );
and ( n11234 , n11170 , n11233 );
or ( n11235 , n11169 , n11234 );
and ( n11236 , n11166 , n11235 );
or ( n11237 , n11165 , n11236 );
and ( n11238 , n11162 , n11237 );
or ( n11239 , n11161 , n11238 );
and ( n11240 , n11158 , n11239 );
or ( n11241 , n11157 , n11240 );
and ( n11242 , n11154 , n11241 );
or ( n11243 , n11153 , n11242 );
and ( n11244 , n816 , n6857 );
and ( n11245 , n11243 , n11244 );
xor ( n11246 , n11243 , n11244 );
xor ( n11247 , n11154 , n11241 );
and ( n11248 , n817 , n6857 );
and ( n11249 , n11247 , n11248 );
xor ( n11250 , n11247 , n11248 );
xor ( n11251 , n11158 , n11239 );
and ( n11252 , n818 , n6857 );
and ( n11253 , n11251 , n11252 );
xor ( n11254 , n11251 , n11252 );
xor ( n11255 , n11162 , n11237 );
and ( n11256 , n819 , n6857 );
and ( n11257 , n11255 , n11256 );
xor ( n11258 , n11255 , n11256 );
xor ( n11259 , n11166 , n11235 );
and ( n11260 , n820 , n6857 );
and ( n11261 , n11259 , n11260 );
xor ( n11262 , n11259 , n11260 );
xor ( n11263 , n11170 , n11233 );
and ( n11264 , n821 , n6857 );
and ( n11265 , n11263 , n11264 );
xor ( n11266 , n11263 , n11264 );
xor ( n11267 , n11174 , n11231 );
and ( n11268 , n822 , n6857 );
and ( n11269 , n11267 , n11268 );
xor ( n11270 , n11267 , n11268 );
xor ( n11271 , n11178 , n11229 );
and ( n11272 , n823 , n6857 );
and ( n11273 , n11271 , n11272 );
xor ( n11274 , n11271 , n11272 );
xor ( n11275 , n11182 , n11227 );
and ( n11276 , n824 , n6857 );
and ( n11277 , n11275 , n11276 );
xor ( n11278 , n11275 , n11276 );
xor ( n11279 , n11186 , n11225 );
and ( n11280 , n825 , n6857 );
and ( n11281 , n11279 , n11280 );
xor ( n11282 , n11279 , n11280 );
xor ( n11283 , n11190 , n11223 );
and ( n11284 , n826 , n6857 );
and ( n11285 , n11283 , n11284 );
xor ( n11286 , n11283 , n11284 );
xor ( n11287 , n11194 , n11221 );
and ( n11288 , n827 , n6857 );
and ( n11289 , n11287 , n11288 );
xor ( n11290 , n11287 , n11288 );
xor ( n11291 , n11198 , n11219 );
and ( n11292 , n828 , n6857 );
and ( n11293 , n11291 , n11292 );
xor ( n11294 , n11291 , n11292 );
xor ( n11295 , n11202 , n11217 );
and ( n11296 , n829 , n6857 );
and ( n11297 , n11295 , n11296 );
xor ( n11298 , n11295 , n11296 );
xor ( n11299 , n11206 , n11215 );
and ( n11300 , n830 , n6857 );
and ( n11301 , n11299 , n11300 );
xor ( n11302 , n11299 , n11300 );
xor ( n11303 , n11210 , n11213 );
and ( n11304 , n831 , n6857 );
and ( n11305 , n11303 , n11304 );
and ( n11306 , n11302 , n11305 );
or ( n11307 , n11301 , n11306 );
and ( n11308 , n11298 , n11307 );
or ( n11309 , n11297 , n11308 );
and ( n11310 , n11294 , n11309 );
or ( n11311 , n11293 , n11310 );
and ( n11312 , n11290 , n11311 );
or ( n11313 , n11289 , n11312 );
and ( n11314 , n11286 , n11313 );
or ( n11315 , n11285 , n11314 );
and ( n11316 , n11282 , n11315 );
or ( n11317 , n11281 , n11316 );
and ( n11318 , n11278 , n11317 );
or ( n11319 , n11277 , n11318 );
and ( n11320 , n11274 , n11319 );
or ( n11321 , n11273 , n11320 );
and ( n11322 , n11270 , n11321 );
or ( n11323 , n11269 , n11322 );
and ( n11324 , n11266 , n11323 );
or ( n11325 , n11265 , n11324 );
and ( n11326 , n11262 , n11325 );
or ( n11327 , n11261 , n11326 );
and ( n11328 , n11258 , n11327 );
or ( n11329 , n11257 , n11328 );
and ( n11330 , n11254 , n11329 );
or ( n11331 , n11253 , n11330 );
and ( n11332 , n11250 , n11331 );
or ( n11333 , n11249 , n11332 );
and ( n11334 , n11246 , n11333 );
or ( n11335 , n11245 , n11334 );
and ( n11336 , n816 , n6854 );
and ( n11337 , n11335 , n11336 );
xor ( n11338 , n11335 , n11336 );
xor ( n11339 , n11246 , n11333 );
and ( n11340 , n817 , n6854 );
and ( n11341 , n11339 , n11340 );
xor ( n11342 , n11339 , n11340 );
xor ( n11343 , n11250 , n11331 );
and ( n11344 , n818 , n6854 );
and ( n11345 , n11343 , n11344 );
xor ( n11346 , n11343 , n11344 );
xor ( n11347 , n11254 , n11329 );
and ( n11348 , n819 , n6854 );
and ( n11349 , n11347 , n11348 );
xor ( n11350 , n11347 , n11348 );
xor ( n11351 , n11258 , n11327 );
and ( n11352 , n820 , n6854 );
and ( n11353 , n11351 , n11352 );
xor ( n11354 , n11351 , n11352 );
xor ( n11355 , n11262 , n11325 );
and ( n11356 , n821 , n6854 );
and ( n11357 , n11355 , n11356 );
xor ( n11358 , n11355 , n11356 );
xor ( n11359 , n11266 , n11323 );
and ( n11360 , n822 , n6854 );
and ( n11361 , n11359 , n11360 );
xor ( n11362 , n11359 , n11360 );
xor ( n11363 , n11270 , n11321 );
and ( n11364 , n823 , n6854 );
and ( n11365 , n11363 , n11364 );
xor ( n11366 , n11363 , n11364 );
xor ( n11367 , n11274 , n11319 );
and ( n11368 , n824 , n6854 );
and ( n11369 , n11367 , n11368 );
xor ( n11370 , n11367 , n11368 );
xor ( n11371 , n11278 , n11317 );
and ( n11372 , n825 , n6854 );
and ( n11373 , n11371 , n11372 );
xor ( n11374 , n11371 , n11372 );
xor ( n11375 , n11282 , n11315 );
and ( n11376 , n826 , n6854 );
and ( n11377 , n11375 , n11376 );
xor ( n11378 , n11375 , n11376 );
xor ( n11379 , n11286 , n11313 );
and ( n11380 , n827 , n6854 );
and ( n11381 , n11379 , n11380 );
xor ( n11382 , n11379 , n11380 );
xor ( n11383 , n11290 , n11311 );
and ( n11384 , n828 , n6854 );
and ( n11385 , n11383 , n11384 );
xor ( n11386 , n11383 , n11384 );
xor ( n11387 , n11294 , n11309 );
and ( n11388 , n829 , n6854 );
and ( n11389 , n11387 , n11388 );
xor ( n11390 , n11387 , n11388 );
xor ( n11391 , n11298 , n11307 );
and ( n11392 , n830 , n6854 );
and ( n11393 , n11391 , n11392 );
xor ( n11394 , n11391 , n11392 );
xor ( n11395 , n11302 , n11305 );
and ( n11396 , n831 , n6854 );
and ( n11397 , n11395 , n11396 );
and ( n11398 , n11394 , n11397 );
or ( n11399 , n11393 , n11398 );
and ( n11400 , n11390 , n11399 );
or ( n11401 , n11389 , n11400 );
and ( n11402 , n11386 , n11401 );
or ( n11403 , n11385 , n11402 );
and ( n11404 , n11382 , n11403 );
or ( n11405 , n11381 , n11404 );
and ( n11406 , n11378 , n11405 );
or ( n11407 , n11377 , n11406 );
and ( n11408 , n11374 , n11407 );
or ( n11409 , n11373 , n11408 );
and ( n11410 , n11370 , n11409 );
or ( n11411 , n11369 , n11410 );
and ( n11412 , n11366 , n11411 );
or ( n11413 , n11365 , n11412 );
and ( n11414 , n11362 , n11413 );
or ( n11415 , n11361 , n11414 );
and ( n11416 , n11358 , n11415 );
or ( n11417 , n11357 , n11416 );
and ( n11418 , n11354 , n11417 );
or ( n11419 , n11353 , n11418 );
and ( n11420 , n11350 , n11419 );
or ( n11421 , n11349 , n11420 );
and ( n11422 , n11346 , n11421 );
or ( n11423 , n11345 , n11422 );
and ( n11424 , n11342 , n11423 );
or ( n11425 , n11341 , n11424 );
and ( n11426 , n11338 , n11425 );
or ( n11427 , n11337 , n11426 );
and ( n11428 , n816 , n6851 );
and ( n11429 , n11427 , n11428 );
xor ( n11430 , n11427 , n11428 );
xor ( n11431 , n11338 , n11425 );
and ( n11432 , n817 , n6851 );
and ( n11433 , n11431 , n11432 );
xor ( n11434 , n11431 , n11432 );
xor ( n11435 , n11342 , n11423 );
and ( n11436 , n818 , n6851 );
and ( n11437 , n11435 , n11436 );
xor ( n11438 , n11435 , n11436 );
xor ( n11439 , n11346 , n11421 );
and ( n11440 , n819 , n6851 );
and ( n11441 , n11439 , n11440 );
xor ( n11442 , n11439 , n11440 );
xor ( n11443 , n11350 , n11419 );
and ( n11444 , n820 , n6851 );
and ( n11445 , n11443 , n11444 );
xor ( n11446 , n11443 , n11444 );
xor ( n11447 , n11354 , n11417 );
and ( n11448 , n821 , n6851 );
and ( n11449 , n11447 , n11448 );
xor ( n11450 , n11447 , n11448 );
xor ( n11451 , n11358 , n11415 );
and ( n11452 , n822 , n6851 );
and ( n11453 , n11451 , n11452 );
xor ( n11454 , n11451 , n11452 );
xor ( n11455 , n11362 , n11413 );
and ( n11456 , n823 , n6851 );
and ( n11457 , n11455 , n11456 );
xor ( n11458 , n11455 , n11456 );
xor ( n11459 , n11366 , n11411 );
and ( n11460 , n824 , n6851 );
and ( n11461 , n11459 , n11460 );
xor ( n11462 , n11459 , n11460 );
xor ( n11463 , n11370 , n11409 );
and ( n11464 , n825 , n6851 );
and ( n11465 , n11463 , n11464 );
xor ( n11466 , n11463 , n11464 );
xor ( n11467 , n11374 , n11407 );
and ( n11468 , n826 , n6851 );
and ( n11469 , n11467 , n11468 );
xor ( n11470 , n11467 , n11468 );
xor ( n11471 , n11378 , n11405 );
and ( n11472 , n827 , n6851 );
and ( n11473 , n11471 , n11472 );
xor ( n11474 , n11471 , n11472 );
xor ( n11475 , n11382 , n11403 );
and ( n11476 , n828 , n6851 );
and ( n11477 , n11475 , n11476 );
xor ( n11478 , n11475 , n11476 );
xor ( n11479 , n11386 , n11401 );
and ( n11480 , n829 , n6851 );
and ( n11481 , n11479 , n11480 );
xor ( n11482 , n11479 , n11480 );
xor ( n11483 , n11390 , n11399 );
and ( n11484 , n830 , n6851 );
and ( n11485 , n11483 , n11484 );
xor ( n11486 , n11483 , n11484 );
xor ( n11487 , n11394 , n11397 );
and ( n11488 , n831 , n6851 );
and ( n11489 , n11487 , n11488 );
and ( n11490 , n11486 , n11489 );
or ( n11491 , n11485 , n11490 );
and ( n11492 , n11482 , n11491 );
or ( n11493 , n11481 , n11492 );
and ( n11494 , n11478 , n11493 );
or ( n11495 , n11477 , n11494 );
and ( n11496 , n11474 , n11495 );
or ( n11497 , n11473 , n11496 );
and ( n11498 , n11470 , n11497 );
or ( n11499 , n11469 , n11498 );
and ( n11500 , n11466 , n11499 );
or ( n11501 , n11465 , n11500 );
and ( n11502 , n11462 , n11501 );
or ( n11503 , n11461 , n11502 );
and ( n11504 , n11458 , n11503 );
or ( n11505 , n11457 , n11504 );
and ( n11506 , n11454 , n11505 );
or ( n11507 , n11453 , n11506 );
and ( n11508 , n11450 , n11507 );
or ( n11509 , n11449 , n11508 );
and ( n11510 , n11446 , n11509 );
or ( n11511 , n11445 , n11510 );
and ( n11512 , n11442 , n11511 );
or ( n11513 , n11441 , n11512 );
and ( n11514 , n11438 , n11513 );
or ( n11515 , n11437 , n11514 );
and ( n11516 , n11434 , n11515 );
or ( n11517 , n11433 , n11516 );
and ( n11518 , n11430 , n11517 );
or ( n11519 , n11429 , n11518 );
and ( n11520 , n816 , n6848 );
and ( n11521 , n11519 , n11520 );
xor ( n11522 , n11519 , n11520 );
xor ( n11523 , n11430 , n11517 );
and ( n11524 , n817 , n6848 );
and ( n11525 , n11523 , n11524 );
xor ( n11526 , n11523 , n11524 );
xor ( n11527 , n11434 , n11515 );
and ( n11528 , n818 , n6848 );
and ( n11529 , n11527 , n11528 );
xor ( n11530 , n11527 , n11528 );
xor ( n11531 , n11438 , n11513 );
and ( n11532 , n819 , n6848 );
and ( n11533 , n11531 , n11532 );
xor ( n11534 , n11531 , n11532 );
xor ( n11535 , n11442 , n11511 );
and ( n11536 , n820 , n6848 );
and ( n11537 , n11535 , n11536 );
xor ( n11538 , n11535 , n11536 );
xor ( n11539 , n11446 , n11509 );
and ( n11540 , n821 , n6848 );
and ( n11541 , n11539 , n11540 );
xor ( n11542 , n11539 , n11540 );
xor ( n11543 , n11450 , n11507 );
and ( n11544 , n822 , n6848 );
and ( n11545 , n11543 , n11544 );
xor ( n11546 , n11543 , n11544 );
xor ( n11547 , n11454 , n11505 );
and ( n11548 , n823 , n6848 );
and ( n11549 , n11547 , n11548 );
xor ( n11550 , n11547 , n11548 );
xor ( n11551 , n11458 , n11503 );
and ( n11552 , n824 , n6848 );
and ( n11553 , n11551 , n11552 );
xor ( n11554 , n11551 , n11552 );
xor ( n11555 , n11462 , n11501 );
and ( n11556 , n825 , n6848 );
and ( n11557 , n11555 , n11556 );
xor ( n11558 , n11555 , n11556 );
xor ( n11559 , n11466 , n11499 );
and ( n11560 , n826 , n6848 );
and ( n11561 , n11559 , n11560 );
xor ( n11562 , n11559 , n11560 );
xor ( n11563 , n11470 , n11497 );
and ( n11564 , n827 , n6848 );
and ( n11565 , n11563 , n11564 );
xor ( n11566 , n11563 , n11564 );
xor ( n11567 , n11474 , n11495 );
and ( n11568 , n828 , n6848 );
and ( n11569 , n11567 , n11568 );
xor ( n11570 , n11567 , n11568 );
xor ( n11571 , n11478 , n11493 );
and ( n11572 , n829 , n6848 );
and ( n11573 , n11571 , n11572 );
xor ( n11574 , n11571 , n11572 );
xor ( n11575 , n11482 , n11491 );
and ( n11576 , n830 , n6848 );
and ( n11577 , n11575 , n11576 );
xor ( n11578 , n11575 , n11576 );
xor ( n11579 , n11486 , n11489 );
and ( n11580 , n831 , n6848 );
and ( n11581 , n11579 , n11580 );
and ( n11582 , n11578 , n11581 );
or ( n11583 , n11577 , n11582 );
and ( n11584 , n11574 , n11583 );
or ( n11585 , n11573 , n11584 );
and ( n11586 , n11570 , n11585 );
or ( n11587 , n11569 , n11586 );
and ( n11588 , n11566 , n11587 );
or ( n11589 , n11565 , n11588 );
and ( n11590 , n11562 , n11589 );
or ( n11591 , n11561 , n11590 );
and ( n11592 , n11558 , n11591 );
or ( n11593 , n11557 , n11592 );
and ( n11594 , n11554 , n11593 );
or ( n11595 , n11553 , n11594 );
and ( n11596 , n11550 , n11595 );
or ( n11597 , n11549 , n11596 );
and ( n11598 , n11546 , n11597 );
or ( n11599 , n11545 , n11598 );
and ( n11600 , n11542 , n11599 );
or ( n11601 , n11541 , n11600 );
and ( n11602 , n11538 , n11601 );
or ( n11603 , n11537 , n11602 );
and ( n11604 , n11534 , n11603 );
or ( n11605 , n11533 , n11604 );
and ( n11606 , n11530 , n11605 );
or ( n11607 , n11529 , n11606 );
and ( n11608 , n11526 , n11607 );
or ( n11609 , n11525 , n11608 );
and ( n11610 , n11522 , n11609 );
or ( n11611 , n11521 , n11610 );
and ( n11612 , n816 , n6845 );
and ( n11613 , n11611 , n11612 );
xor ( n11614 , n11611 , n11612 );
xor ( n11615 , n11522 , n11609 );
and ( n11616 , n817 , n6845 );
and ( n11617 , n11615 , n11616 );
xor ( n11618 , n11615 , n11616 );
xor ( n11619 , n11526 , n11607 );
and ( n11620 , n818 , n6845 );
and ( n11621 , n11619 , n11620 );
xor ( n11622 , n11619 , n11620 );
xor ( n11623 , n11530 , n11605 );
and ( n11624 , n819 , n6845 );
and ( n11625 , n11623 , n11624 );
xor ( n11626 , n11623 , n11624 );
xor ( n11627 , n11534 , n11603 );
and ( n11628 , n820 , n6845 );
and ( n11629 , n11627 , n11628 );
xor ( n11630 , n11627 , n11628 );
xor ( n11631 , n11538 , n11601 );
and ( n11632 , n821 , n6845 );
and ( n11633 , n11631 , n11632 );
xor ( n11634 , n11631 , n11632 );
xor ( n11635 , n11542 , n11599 );
and ( n11636 , n822 , n6845 );
and ( n11637 , n11635 , n11636 );
xor ( n11638 , n11635 , n11636 );
xor ( n11639 , n11546 , n11597 );
and ( n11640 , n823 , n6845 );
and ( n11641 , n11639 , n11640 );
xor ( n11642 , n11639 , n11640 );
xor ( n11643 , n11550 , n11595 );
and ( n11644 , n824 , n6845 );
and ( n11645 , n11643 , n11644 );
xor ( n11646 , n11643 , n11644 );
xor ( n11647 , n11554 , n11593 );
and ( n11648 , n825 , n6845 );
and ( n11649 , n11647 , n11648 );
xor ( n11650 , n11647 , n11648 );
xor ( n11651 , n11558 , n11591 );
and ( n11652 , n826 , n6845 );
and ( n11653 , n11651 , n11652 );
xor ( n11654 , n11651 , n11652 );
xor ( n11655 , n11562 , n11589 );
and ( n11656 , n827 , n6845 );
and ( n11657 , n11655 , n11656 );
xor ( n11658 , n11655 , n11656 );
xor ( n11659 , n11566 , n11587 );
and ( n11660 , n828 , n6845 );
and ( n11661 , n11659 , n11660 );
xor ( n11662 , n11659 , n11660 );
xor ( n11663 , n11570 , n11585 );
and ( n11664 , n829 , n6845 );
and ( n11665 , n11663 , n11664 );
xor ( n11666 , n11663 , n11664 );
xor ( n11667 , n11574 , n11583 );
and ( n11668 , n830 , n6845 );
and ( n11669 , n11667 , n11668 );
xor ( n11670 , n11667 , n11668 );
xor ( n11671 , n11578 , n11581 );
and ( n11672 , n831 , n6845 );
and ( n11673 , n11671 , n11672 );
and ( n11674 , n11670 , n11673 );
or ( n11675 , n11669 , n11674 );
and ( n11676 , n11666 , n11675 );
or ( n11677 , n11665 , n11676 );
and ( n11678 , n11662 , n11677 );
or ( n11679 , n11661 , n11678 );
and ( n11680 , n11658 , n11679 );
or ( n11681 , n11657 , n11680 );
and ( n11682 , n11654 , n11681 );
or ( n11683 , n11653 , n11682 );
and ( n11684 , n11650 , n11683 );
or ( n11685 , n11649 , n11684 );
and ( n11686 , n11646 , n11685 );
or ( n11687 , n11645 , n11686 );
and ( n11688 , n11642 , n11687 );
or ( n11689 , n11641 , n11688 );
and ( n11690 , n11638 , n11689 );
or ( n11691 , n11637 , n11690 );
and ( n11692 , n11634 , n11691 );
or ( n11693 , n11633 , n11692 );
and ( n11694 , n11630 , n11693 );
or ( n11695 , n11629 , n11694 );
and ( n11696 , n11626 , n11695 );
or ( n11697 , n11625 , n11696 );
and ( n11698 , n11622 , n11697 );
or ( n11699 , n11621 , n11698 );
and ( n11700 , n11618 , n11699 );
or ( n11701 , n11617 , n11700 );
and ( n11702 , n11614 , n11701 );
or ( n11703 , n11613 , n11702 );
and ( n11704 , n816 , n6842 );
and ( n11705 , n11703 , n11704 );
xor ( n11706 , n11703 , n11704 );
xor ( n11707 , n11614 , n11701 );
and ( n11708 , n817 , n6842 );
and ( n11709 , n11707 , n11708 );
xor ( n11710 , n11707 , n11708 );
xor ( n11711 , n11618 , n11699 );
and ( n11712 , n818 , n6842 );
and ( n11713 , n11711 , n11712 );
xor ( n11714 , n11711 , n11712 );
xor ( n11715 , n11622 , n11697 );
and ( n11716 , n819 , n6842 );
and ( n11717 , n11715 , n11716 );
xor ( n11718 , n11715 , n11716 );
xor ( n11719 , n11626 , n11695 );
and ( n11720 , n820 , n6842 );
and ( n11721 , n11719 , n11720 );
xor ( n11722 , n11719 , n11720 );
xor ( n11723 , n11630 , n11693 );
and ( n11724 , n821 , n6842 );
and ( n11725 , n11723 , n11724 );
xor ( n11726 , n11723 , n11724 );
xor ( n11727 , n11634 , n11691 );
and ( n11728 , n822 , n6842 );
and ( n11729 , n11727 , n11728 );
xor ( n11730 , n11727 , n11728 );
xor ( n11731 , n11638 , n11689 );
and ( n11732 , n823 , n6842 );
and ( n11733 , n11731 , n11732 );
xor ( n11734 , n11731 , n11732 );
xor ( n11735 , n11642 , n11687 );
and ( n11736 , n824 , n6842 );
and ( n11737 , n11735 , n11736 );
xor ( n11738 , n11735 , n11736 );
xor ( n11739 , n11646 , n11685 );
and ( n11740 , n825 , n6842 );
and ( n11741 , n11739 , n11740 );
xor ( n11742 , n11739 , n11740 );
xor ( n11743 , n11650 , n11683 );
and ( n11744 , n826 , n6842 );
and ( n11745 , n11743 , n11744 );
xor ( n11746 , n11743 , n11744 );
xor ( n11747 , n11654 , n11681 );
and ( n11748 , n827 , n6842 );
and ( n11749 , n11747 , n11748 );
xor ( n11750 , n11747 , n11748 );
xor ( n11751 , n11658 , n11679 );
and ( n11752 , n828 , n6842 );
and ( n11753 , n11751 , n11752 );
xor ( n11754 , n11751 , n11752 );
xor ( n11755 , n11662 , n11677 );
and ( n11756 , n829 , n6842 );
and ( n11757 , n11755 , n11756 );
xor ( n11758 , n11755 , n11756 );
xor ( n11759 , n11666 , n11675 );
and ( n11760 , n830 , n6842 );
and ( n11761 , n11759 , n11760 );
xor ( n11762 , n11759 , n11760 );
xor ( n11763 , n11670 , n11673 );
and ( n11764 , n831 , n6842 );
and ( n11765 , n11763 , n11764 );
and ( n11766 , n11762 , n11765 );
or ( n11767 , n11761 , n11766 );
and ( n11768 , n11758 , n11767 );
or ( n11769 , n11757 , n11768 );
and ( n11770 , n11754 , n11769 );
or ( n11771 , n11753 , n11770 );
and ( n11772 , n11750 , n11771 );
or ( n11773 , n11749 , n11772 );
and ( n11774 , n11746 , n11773 );
or ( n11775 , n11745 , n11774 );
and ( n11776 , n11742 , n11775 );
or ( n11777 , n11741 , n11776 );
and ( n11778 , n11738 , n11777 );
or ( n11779 , n11737 , n11778 );
and ( n11780 , n11734 , n11779 );
or ( n11781 , n11733 , n11780 );
and ( n11782 , n11730 , n11781 );
or ( n11783 , n11729 , n11782 );
and ( n11784 , n11726 , n11783 );
or ( n11785 , n11725 , n11784 );
and ( n11786 , n11722 , n11785 );
or ( n11787 , n11721 , n11786 );
and ( n11788 , n11718 , n11787 );
or ( n11789 , n11717 , n11788 );
and ( n11790 , n11714 , n11789 );
or ( n11791 , n11713 , n11790 );
and ( n11792 , n11710 , n11791 );
or ( n11793 , n11709 , n11792 );
and ( n11794 , n11706 , n11793 );
or ( n11795 , n11705 , n11794 );
and ( n11796 , n816 , n6839 );
and ( n11797 , n11795 , n11796 );
xor ( n11798 , n11795 , n11796 );
xor ( n11799 , n11706 , n11793 );
and ( n11800 , n817 , n6839 );
and ( n11801 , n11799 , n11800 );
xor ( n11802 , n11799 , n11800 );
xor ( n11803 , n11710 , n11791 );
and ( n11804 , n818 , n6839 );
and ( n11805 , n11803 , n11804 );
xor ( n11806 , n11803 , n11804 );
xor ( n11807 , n11714 , n11789 );
and ( n11808 , n819 , n6839 );
and ( n11809 , n11807 , n11808 );
xor ( n11810 , n11807 , n11808 );
xor ( n11811 , n11718 , n11787 );
and ( n11812 , n820 , n6839 );
and ( n11813 , n11811 , n11812 );
xor ( n11814 , n11811 , n11812 );
xor ( n11815 , n11722 , n11785 );
and ( n11816 , n821 , n6839 );
and ( n11817 , n11815 , n11816 );
xor ( n11818 , n11815 , n11816 );
xor ( n11819 , n11726 , n11783 );
and ( n11820 , n822 , n6839 );
and ( n11821 , n11819 , n11820 );
xor ( n11822 , n11819 , n11820 );
xor ( n11823 , n11730 , n11781 );
and ( n11824 , n823 , n6839 );
and ( n11825 , n11823 , n11824 );
xor ( n11826 , n11823 , n11824 );
xor ( n11827 , n11734 , n11779 );
and ( n11828 , n824 , n6839 );
and ( n11829 , n11827 , n11828 );
xor ( n11830 , n11827 , n11828 );
xor ( n11831 , n11738 , n11777 );
and ( n11832 , n825 , n6839 );
and ( n11833 , n11831 , n11832 );
xor ( n11834 , n11831 , n11832 );
xor ( n11835 , n11742 , n11775 );
and ( n11836 , n826 , n6839 );
and ( n11837 , n11835 , n11836 );
xor ( n11838 , n11835 , n11836 );
xor ( n11839 , n11746 , n11773 );
and ( n11840 , n827 , n6839 );
and ( n11841 , n11839 , n11840 );
xor ( n11842 , n11839 , n11840 );
xor ( n11843 , n11750 , n11771 );
and ( n11844 , n828 , n6839 );
and ( n11845 , n11843 , n11844 );
xor ( n11846 , n11843 , n11844 );
xor ( n11847 , n11754 , n11769 );
and ( n11848 , n829 , n6839 );
and ( n11849 , n11847 , n11848 );
xor ( n11850 , n11847 , n11848 );
xor ( n11851 , n11758 , n11767 );
and ( n11852 , n830 , n6839 );
and ( n11853 , n11851 , n11852 );
xor ( n11854 , n11851 , n11852 );
xor ( n11855 , n11762 , n11765 );
and ( n11856 , n831 , n6839 );
and ( n11857 , n11855 , n11856 );
and ( n11858 , n11854 , n11857 );
or ( n11859 , n11853 , n11858 );
and ( n11860 , n11850 , n11859 );
or ( n11861 , n11849 , n11860 );
and ( n11862 , n11846 , n11861 );
or ( n11863 , n11845 , n11862 );
and ( n11864 , n11842 , n11863 );
or ( n11865 , n11841 , n11864 );
and ( n11866 , n11838 , n11865 );
or ( n11867 , n11837 , n11866 );
and ( n11868 , n11834 , n11867 );
or ( n11869 , n11833 , n11868 );
and ( n11870 , n11830 , n11869 );
or ( n11871 , n11829 , n11870 );
and ( n11872 , n11826 , n11871 );
or ( n11873 , n11825 , n11872 );
and ( n11874 , n11822 , n11873 );
or ( n11875 , n11821 , n11874 );
and ( n11876 , n11818 , n11875 );
or ( n11877 , n11817 , n11876 );
and ( n11878 , n11814 , n11877 );
or ( n11879 , n11813 , n11878 );
and ( n11880 , n11810 , n11879 );
or ( n11881 , n11809 , n11880 );
and ( n11882 , n11806 , n11881 );
or ( n11883 , n11805 , n11882 );
and ( n11884 , n11802 , n11883 );
or ( n11885 , n11801 , n11884 );
and ( n11886 , n11798 , n11885 );
or ( n11887 , n11797 , n11886 );
and ( n11888 , n816 , n6836 );
and ( n11889 , n11887 , n11888 );
xor ( n11890 , n11887 , n11888 );
xor ( n11891 , n11798 , n11885 );
and ( n11892 , n817 , n6836 );
and ( n11893 , n11891 , n11892 );
xor ( n11894 , n11891 , n11892 );
xor ( n11895 , n11802 , n11883 );
and ( n11896 , n818 , n6836 );
and ( n11897 , n11895 , n11896 );
xor ( n11898 , n11895 , n11896 );
xor ( n11899 , n11806 , n11881 );
and ( n11900 , n819 , n6836 );
and ( n11901 , n11899 , n11900 );
xor ( n11902 , n11899 , n11900 );
xor ( n11903 , n11810 , n11879 );
and ( n11904 , n820 , n6836 );
and ( n11905 , n11903 , n11904 );
xor ( n11906 , n11903 , n11904 );
xor ( n11907 , n11814 , n11877 );
and ( n11908 , n821 , n6836 );
and ( n11909 , n11907 , n11908 );
xor ( n11910 , n11907 , n11908 );
xor ( n11911 , n11818 , n11875 );
and ( n11912 , n822 , n6836 );
and ( n11913 , n11911 , n11912 );
xor ( n11914 , n11911 , n11912 );
xor ( n11915 , n11822 , n11873 );
and ( n11916 , n823 , n6836 );
and ( n11917 , n11915 , n11916 );
xor ( n11918 , n11915 , n11916 );
xor ( n11919 , n11826 , n11871 );
and ( n11920 , n824 , n6836 );
and ( n11921 , n11919 , n11920 );
xor ( n11922 , n11919 , n11920 );
xor ( n11923 , n11830 , n11869 );
and ( n11924 , n825 , n6836 );
and ( n11925 , n11923 , n11924 );
xor ( n11926 , n11923 , n11924 );
xor ( n11927 , n11834 , n11867 );
and ( n11928 , n826 , n6836 );
and ( n11929 , n11927 , n11928 );
xor ( n11930 , n11927 , n11928 );
xor ( n11931 , n11838 , n11865 );
and ( n11932 , n827 , n6836 );
and ( n11933 , n11931 , n11932 );
xor ( n11934 , n11931 , n11932 );
xor ( n11935 , n11842 , n11863 );
and ( n11936 , n828 , n6836 );
and ( n11937 , n11935 , n11936 );
xor ( n11938 , n11935 , n11936 );
xor ( n11939 , n11846 , n11861 );
and ( n11940 , n829 , n6836 );
and ( n11941 , n11939 , n11940 );
xor ( n11942 , n11939 , n11940 );
xor ( n11943 , n11850 , n11859 );
and ( n11944 , n830 , n6836 );
and ( n11945 , n11943 , n11944 );
xor ( n11946 , n11943 , n11944 );
xor ( n11947 , n11854 , n11857 );
and ( n11948 , n831 , n6836 );
and ( n11949 , n11947 , n11948 );
and ( n11950 , n11946 , n11949 );
or ( n11951 , n11945 , n11950 );
and ( n11952 , n11942 , n11951 );
or ( n11953 , n11941 , n11952 );
and ( n11954 , n11938 , n11953 );
or ( n11955 , n11937 , n11954 );
and ( n11956 , n11934 , n11955 );
or ( n11957 , n11933 , n11956 );
and ( n11958 , n11930 , n11957 );
or ( n11959 , n11929 , n11958 );
and ( n11960 , n11926 , n11959 );
or ( n11961 , n11925 , n11960 );
and ( n11962 , n11922 , n11961 );
or ( n11963 , n11921 , n11962 );
and ( n11964 , n11918 , n11963 );
or ( n11965 , n11917 , n11964 );
and ( n11966 , n11914 , n11965 );
or ( n11967 , n11913 , n11966 );
and ( n11968 , n11910 , n11967 );
or ( n11969 , n11909 , n11968 );
and ( n11970 , n11906 , n11969 );
or ( n11971 , n11905 , n11970 );
and ( n11972 , n11902 , n11971 );
or ( n11973 , n11901 , n11972 );
and ( n11974 , n11898 , n11973 );
or ( n11975 , n11897 , n11974 );
and ( n11976 , n11894 , n11975 );
or ( n11977 , n11893 , n11976 );
and ( n11978 , n11890 , n11977 );
or ( n11979 , n11889 , n11978 );
and ( n11980 , n816 , n6833 );
and ( n11981 , n11979 , n11980 );
xor ( n11982 , n11979 , n11980 );
xor ( n11983 , n11890 , n11977 );
and ( n11984 , n817 , n6833 );
and ( n11985 , n11983 , n11984 );
xor ( n11986 , n11983 , n11984 );
xor ( n11987 , n11894 , n11975 );
and ( n11988 , n818 , n6833 );
and ( n11989 , n11987 , n11988 );
xor ( n11990 , n11987 , n11988 );
xor ( n11991 , n11898 , n11973 );
and ( n11992 , n819 , n6833 );
and ( n11993 , n11991 , n11992 );
xor ( n11994 , n11991 , n11992 );
xor ( n11995 , n11902 , n11971 );
and ( n11996 , n820 , n6833 );
and ( n11997 , n11995 , n11996 );
xor ( n11998 , n11995 , n11996 );
xor ( n11999 , n11906 , n11969 );
and ( n12000 , n821 , n6833 );
and ( n12001 , n11999 , n12000 );
xor ( n12002 , n11999 , n12000 );
xor ( n12003 , n11910 , n11967 );
and ( n12004 , n822 , n6833 );
and ( n12005 , n12003 , n12004 );
xor ( n12006 , n12003 , n12004 );
xor ( n12007 , n11914 , n11965 );
and ( n12008 , n823 , n6833 );
and ( n12009 , n12007 , n12008 );
xor ( n12010 , n12007 , n12008 );
xor ( n12011 , n11918 , n11963 );
and ( n12012 , n824 , n6833 );
and ( n12013 , n12011 , n12012 );
xor ( n12014 , n12011 , n12012 );
xor ( n12015 , n11922 , n11961 );
and ( n12016 , n825 , n6833 );
and ( n12017 , n12015 , n12016 );
xor ( n12018 , n12015 , n12016 );
xor ( n12019 , n11926 , n11959 );
and ( n12020 , n826 , n6833 );
and ( n12021 , n12019 , n12020 );
xor ( n12022 , n12019 , n12020 );
xor ( n12023 , n11930 , n11957 );
and ( n12024 , n827 , n6833 );
and ( n12025 , n12023 , n12024 );
xor ( n12026 , n12023 , n12024 );
xor ( n12027 , n11934 , n11955 );
and ( n12028 , n828 , n6833 );
and ( n12029 , n12027 , n12028 );
xor ( n12030 , n12027 , n12028 );
xor ( n12031 , n11938 , n11953 );
and ( n12032 , n829 , n6833 );
and ( n12033 , n12031 , n12032 );
xor ( n12034 , n12031 , n12032 );
xor ( n12035 , n11942 , n11951 );
and ( n12036 , n830 , n6833 );
and ( n12037 , n12035 , n12036 );
xor ( n12038 , n12035 , n12036 );
xor ( n12039 , n11946 , n11949 );
and ( n12040 , n831 , n6833 );
and ( n12041 , n12039 , n12040 );
and ( n12042 , n12038 , n12041 );
or ( n12043 , n12037 , n12042 );
and ( n12044 , n12034 , n12043 );
or ( n12045 , n12033 , n12044 );
and ( n12046 , n12030 , n12045 );
or ( n12047 , n12029 , n12046 );
and ( n12048 , n12026 , n12047 );
or ( n12049 , n12025 , n12048 );
and ( n12050 , n12022 , n12049 );
or ( n12051 , n12021 , n12050 );
and ( n12052 , n12018 , n12051 );
or ( n12053 , n12017 , n12052 );
and ( n12054 , n12014 , n12053 );
or ( n12055 , n12013 , n12054 );
and ( n12056 , n12010 , n12055 );
or ( n12057 , n12009 , n12056 );
and ( n12058 , n12006 , n12057 );
or ( n12059 , n12005 , n12058 );
and ( n12060 , n12002 , n12059 );
or ( n12061 , n12001 , n12060 );
and ( n12062 , n11998 , n12061 );
or ( n12063 , n11997 , n12062 );
and ( n12064 , n11994 , n12063 );
or ( n12065 , n11993 , n12064 );
and ( n12066 , n11990 , n12065 );
or ( n12067 , n11989 , n12066 );
and ( n12068 , n11986 , n12067 );
or ( n12069 , n11985 , n12068 );
and ( n12070 , n11982 , n12069 );
or ( n12071 , n11981 , n12070 );
and ( n12072 , n816 , n6830 );
and ( n12073 , n12071 , n12072 );
xor ( n12074 , n12071 , n12072 );
xor ( n12075 , n11982 , n12069 );
and ( n12076 , n817 , n6830 );
and ( n12077 , n12075 , n12076 );
xor ( n12078 , n12075 , n12076 );
xor ( n12079 , n11986 , n12067 );
and ( n12080 , n818 , n6830 );
and ( n12081 , n12079 , n12080 );
xor ( n12082 , n12079 , n12080 );
xor ( n12083 , n11990 , n12065 );
and ( n12084 , n819 , n6830 );
and ( n12085 , n12083 , n12084 );
xor ( n12086 , n12083 , n12084 );
xor ( n12087 , n11994 , n12063 );
and ( n12088 , n820 , n6830 );
and ( n12089 , n12087 , n12088 );
xor ( n12090 , n12087 , n12088 );
xor ( n12091 , n11998 , n12061 );
and ( n12092 , n821 , n6830 );
and ( n12093 , n12091 , n12092 );
xor ( n12094 , n12091 , n12092 );
xor ( n12095 , n12002 , n12059 );
and ( n12096 , n822 , n6830 );
and ( n12097 , n12095 , n12096 );
xor ( n12098 , n12095 , n12096 );
xor ( n12099 , n12006 , n12057 );
and ( n12100 , n823 , n6830 );
and ( n12101 , n12099 , n12100 );
xor ( n12102 , n12099 , n12100 );
xor ( n12103 , n12010 , n12055 );
and ( n12104 , n824 , n6830 );
and ( n12105 , n12103 , n12104 );
xor ( n12106 , n12103 , n12104 );
xor ( n12107 , n12014 , n12053 );
and ( n12108 , n825 , n6830 );
and ( n12109 , n12107 , n12108 );
xor ( n12110 , n12107 , n12108 );
xor ( n12111 , n12018 , n12051 );
and ( n12112 , n826 , n6830 );
and ( n12113 , n12111 , n12112 );
xor ( n12114 , n12111 , n12112 );
xor ( n12115 , n12022 , n12049 );
and ( n12116 , n827 , n6830 );
and ( n12117 , n12115 , n12116 );
xor ( n12118 , n12115 , n12116 );
xor ( n12119 , n12026 , n12047 );
and ( n12120 , n828 , n6830 );
and ( n12121 , n12119 , n12120 );
xor ( n12122 , n12119 , n12120 );
xor ( n12123 , n12030 , n12045 );
and ( n12124 , n829 , n6830 );
and ( n12125 , n12123 , n12124 );
xor ( n12126 , n12123 , n12124 );
xor ( n12127 , n12034 , n12043 );
and ( n12128 , n830 , n6830 );
and ( n12129 , n12127 , n12128 );
xor ( n12130 , n12127 , n12128 );
xor ( n12131 , n12038 , n12041 );
and ( n12132 , n831 , n6830 );
and ( n12133 , n12131 , n12132 );
and ( n12134 , n12130 , n12133 );
or ( n12135 , n12129 , n12134 );
and ( n12136 , n12126 , n12135 );
or ( n12137 , n12125 , n12136 );
and ( n12138 , n12122 , n12137 );
or ( n12139 , n12121 , n12138 );
and ( n12140 , n12118 , n12139 );
or ( n12141 , n12117 , n12140 );
and ( n12142 , n12114 , n12141 );
or ( n12143 , n12113 , n12142 );
and ( n12144 , n12110 , n12143 );
or ( n12145 , n12109 , n12144 );
and ( n12146 , n12106 , n12145 );
or ( n12147 , n12105 , n12146 );
and ( n12148 , n12102 , n12147 );
or ( n12149 , n12101 , n12148 );
and ( n12150 , n12098 , n12149 );
or ( n12151 , n12097 , n12150 );
and ( n12152 , n12094 , n12151 );
or ( n12153 , n12093 , n12152 );
and ( n12154 , n12090 , n12153 );
or ( n12155 , n12089 , n12154 );
and ( n12156 , n12086 , n12155 );
or ( n12157 , n12085 , n12156 );
and ( n12158 , n12082 , n12157 );
or ( n12159 , n12081 , n12158 );
and ( n12160 , n12078 , n12159 );
or ( n12161 , n12077 , n12160 );
and ( n12162 , n12074 , n12161 );
or ( n12163 , n12073 , n12162 );
and ( n12164 , n816 , n6827 );
and ( n12165 , n12163 , n12164 );
xor ( n12166 , n12163 , n12164 );
xor ( n12167 , n12074 , n12161 );
and ( n12168 , n817 , n6827 );
and ( n12169 , n12167 , n12168 );
xor ( n12170 , n12167 , n12168 );
xor ( n12171 , n12078 , n12159 );
and ( n12172 , n818 , n6827 );
and ( n12173 , n12171 , n12172 );
xor ( n12174 , n12171 , n12172 );
xor ( n12175 , n12082 , n12157 );
and ( n12176 , n819 , n6827 );
and ( n12177 , n12175 , n12176 );
xor ( n12178 , n12175 , n12176 );
xor ( n12179 , n12086 , n12155 );
and ( n12180 , n820 , n6827 );
and ( n12181 , n12179 , n12180 );
xor ( n12182 , n12179 , n12180 );
xor ( n12183 , n12090 , n12153 );
and ( n12184 , n821 , n6827 );
and ( n12185 , n12183 , n12184 );
xor ( n12186 , n12183 , n12184 );
xor ( n12187 , n12094 , n12151 );
and ( n12188 , n822 , n6827 );
and ( n12189 , n12187 , n12188 );
xor ( n12190 , n12187 , n12188 );
xor ( n12191 , n12098 , n12149 );
and ( n12192 , n823 , n6827 );
and ( n12193 , n12191 , n12192 );
xor ( n12194 , n12191 , n12192 );
xor ( n12195 , n12102 , n12147 );
and ( n12196 , n824 , n6827 );
and ( n12197 , n12195 , n12196 );
xor ( n12198 , n12195 , n12196 );
xor ( n12199 , n12106 , n12145 );
and ( n12200 , n825 , n6827 );
and ( n12201 , n12199 , n12200 );
xor ( n12202 , n12199 , n12200 );
xor ( n12203 , n12110 , n12143 );
and ( n12204 , n826 , n6827 );
and ( n12205 , n12203 , n12204 );
xor ( n12206 , n12203 , n12204 );
xor ( n12207 , n12114 , n12141 );
and ( n12208 , n827 , n6827 );
and ( n12209 , n12207 , n12208 );
xor ( n12210 , n12207 , n12208 );
xor ( n12211 , n12118 , n12139 );
and ( n12212 , n828 , n6827 );
and ( n12213 , n12211 , n12212 );
xor ( n12214 , n12211 , n12212 );
xor ( n12215 , n12122 , n12137 );
and ( n12216 , n829 , n6827 );
and ( n12217 , n12215 , n12216 );
xor ( n12218 , n12215 , n12216 );
xor ( n12219 , n12126 , n12135 );
and ( n12220 , n830 , n6827 );
and ( n12221 , n12219 , n12220 );
xor ( n12222 , n12219 , n12220 );
xor ( n12223 , n12130 , n12133 );
and ( n12224 , n831 , n6827 );
and ( n12225 , n12223 , n12224 );
and ( n12226 , n12222 , n12225 );
or ( n12227 , n12221 , n12226 );
and ( n12228 , n12218 , n12227 );
or ( n12229 , n12217 , n12228 );
and ( n12230 , n12214 , n12229 );
or ( n12231 , n12213 , n12230 );
and ( n12232 , n12210 , n12231 );
or ( n12233 , n12209 , n12232 );
and ( n12234 , n12206 , n12233 );
or ( n12235 , n12205 , n12234 );
and ( n12236 , n12202 , n12235 );
or ( n12237 , n12201 , n12236 );
and ( n12238 , n12198 , n12237 );
or ( n12239 , n12197 , n12238 );
and ( n12240 , n12194 , n12239 );
or ( n12241 , n12193 , n12240 );
and ( n12242 , n12190 , n12241 );
or ( n12243 , n12189 , n12242 );
and ( n12244 , n12186 , n12243 );
or ( n12245 , n12185 , n12244 );
and ( n12246 , n12182 , n12245 );
or ( n12247 , n12181 , n12246 );
and ( n12248 , n12178 , n12247 );
or ( n12249 , n12177 , n12248 );
and ( n12250 , n12174 , n12249 );
or ( n12251 , n12173 , n12250 );
and ( n12252 , n12170 , n12251 );
or ( n12253 , n12169 , n12252 );
and ( n12254 , n12166 , n12253 );
or ( n12255 , n12165 , n12254 );
and ( n12256 , n816 , n6824 );
and ( n12257 , n12255 , n12256 );
xor ( n12258 , n12255 , n12256 );
xor ( n12259 , n12166 , n12253 );
and ( n12260 , n817 , n6824 );
and ( n12261 , n12259 , n12260 );
xor ( n12262 , n12259 , n12260 );
xor ( n12263 , n12170 , n12251 );
and ( n12264 , n818 , n6824 );
and ( n12265 , n12263 , n12264 );
xor ( n12266 , n12263 , n12264 );
xor ( n12267 , n12174 , n12249 );
and ( n12268 , n819 , n6824 );
and ( n12269 , n12267 , n12268 );
xor ( n12270 , n12267 , n12268 );
xor ( n12271 , n12178 , n12247 );
and ( n12272 , n820 , n6824 );
and ( n12273 , n12271 , n12272 );
xor ( n12274 , n12271 , n12272 );
xor ( n12275 , n12182 , n12245 );
and ( n12276 , n821 , n6824 );
and ( n12277 , n12275 , n12276 );
xor ( n12278 , n12275 , n12276 );
xor ( n12279 , n12186 , n12243 );
and ( n12280 , n822 , n6824 );
and ( n12281 , n12279 , n12280 );
xor ( n12282 , n12279 , n12280 );
xor ( n12283 , n12190 , n12241 );
and ( n12284 , n823 , n6824 );
and ( n12285 , n12283 , n12284 );
xor ( n12286 , n12283 , n12284 );
xor ( n12287 , n12194 , n12239 );
and ( n12288 , n824 , n6824 );
and ( n12289 , n12287 , n12288 );
xor ( n12290 , n12287 , n12288 );
xor ( n12291 , n12198 , n12237 );
and ( n12292 , n825 , n6824 );
and ( n12293 , n12291 , n12292 );
xor ( n12294 , n12291 , n12292 );
xor ( n12295 , n12202 , n12235 );
and ( n12296 , n826 , n6824 );
and ( n12297 , n12295 , n12296 );
xor ( n12298 , n12295 , n12296 );
xor ( n12299 , n12206 , n12233 );
and ( n12300 , n827 , n6824 );
and ( n12301 , n12299 , n12300 );
xor ( n12302 , n12299 , n12300 );
xor ( n12303 , n12210 , n12231 );
and ( n12304 , n828 , n6824 );
and ( n12305 , n12303 , n12304 );
xor ( n12306 , n12303 , n12304 );
xor ( n12307 , n12214 , n12229 );
and ( n12308 , n829 , n6824 );
and ( n12309 , n12307 , n12308 );
xor ( n12310 , n12307 , n12308 );
xor ( n12311 , n12218 , n12227 );
and ( n12312 , n830 , n6824 );
and ( n12313 , n12311 , n12312 );
xor ( n12314 , n12311 , n12312 );
xor ( n12315 , n12222 , n12225 );
and ( n12316 , n831 , n6824 );
and ( n12317 , n12315 , n12316 );
and ( n12318 , n12314 , n12317 );
or ( n12319 , n12313 , n12318 );
and ( n12320 , n12310 , n12319 );
or ( n12321 , n12309 , n12320 );
and ( n12322 , n12306 , n12321 );
or ( n12323 , n12305 , n12322 );
and ( n12324 , n12302 , n12323 );
or ( n12325 , n12301 , n12324 );
and ( n12326 , n12298 , n12325 );
or ( n12327 , n12297 , n12326 );
and ( n12328 , n12294 , n12327 );
or ( n12329 , n12293 , n12328 );
and ( n12330 , n12290 , n12329 );
or ( n12331 , n12289 , n12330 );
and ( n12332 , n12286 , n12331 );
or ( n12333 , n12285 , n12332 );
and ( n12334 , n12282 , n12333 );
or ( n12335 , n12281 , n12334 );
and ( n12336 , n12278 , n12335 );
or ( n12337 , n12277 , n12336 );
and ( n12338 , n12274 , n12337 );
or ( n12339 , n12273 , n12338 );
and ( n12340 , n12270 , n12339 );
or ( n12341 , n12269 , n12340 );
and ( n12342 , n12266 , n12341 );
or ( n12343 , n12265 , n12342 );
and ( n12344 , n12262 , n12343 );
or ( n12345 , n12261 , n12344 );
and ( n12346 , n12258 , n12345 );
or ( n12347 , n12257 , n12346 );
and ( n12348 , n816 , n6821 );
and ( n12349 , n12347 , n12348 );
xor ( n12350 , n12347 , n12348 );
xor ( n12351 , n12258 , n12345 );
and ( n12352 , n817 , n6821 );
and ( n12353 , n12351 , n12352 );
xor ( n12354 , n12351 , n12352 );
xor ( n12355 , n12262 , n12343 );
and ( n12356 , n818 , n6821 );
and ( n12357 , n12355 , n12356 );
xor ( n12358 , n12355 , n12356 );
xor ( n12359 , n12266 , n12341 );
and ( n12360 , n819 , n6821 );
and ( n12361 , n12359 , n12360 );
xor ( n12362 , n12359 , n12360 );
xor ( n12363 , n12270 , n12339 );
and ( n12364 , n820 , n6821 );
and ( n12365 , n12363 , n12364 );
xor ( n12366 , n12363 , n12364 );
xor ( n12367 , n12274 , n12337 );
and ( n12368 , n821 , n6821 );
and ( n12369 , n12367 , n12368 );
xor ( n12370 , n12367 , n12368 );
xor ( n12371 , n12278 , n12335 );
and ( n12372 , n822 , n6821 );
and ( n12373 , n12371 , n12372 );
xor ( n12374 , n12371 , n12372 );
xor ( n12375 , n12282 , n12333 );
and ( n12376 , n823 , n6821 );
and ( n12377 , n12375 , n12376 );
xor ( n12378 , n12375 , n12376 );
xor ( n12379 , n12286 , n12331 );
and ( n12380 , n824 , n6821 );
and ( n12381 , n12379 , n12380 );
xor ( n12382 , n12379 , n12380 );
xor ( n12383 , n12290 , n12329 );
and ( n12384 , n825 , n6821 );
and ( n12385 , n12383 , n12384 );
xor ( n12386 , n12383 , n12384 );
xor ( n12387 , n12294 , n12327 );
and ( n12388 , n826 , n6821 );
and ( n12389 , n12387 , n12388 );
xor ( n12390 , n12387 , n12388 );
xor ( n12391 , n12298 , n12325 );
and ( n12392 , n827 , n6821 );
and ( n12393 , n12391 , n12392 );
xor ( n12394 , n12391 , n12392 );
xor ( n12395 , n12302 , n12323 );
and ( n12396 , n828 , n6821 );
and ( n12397 , n12395 , n12396 );
xor ( n12398 , n12395 , n12396 );
xor ( n12399 , n12306 , n12321 );
and ( n12400 , n829 , n6821 );
and ( n12401 , n12399 , n12400 );
xor ( n12402 , n12399 , n12400 );
xor ( n12403 , n12310 , n12319 );
and ( n12404 , n830 , n6821 );
and ( n12405 , n12403 , n12404 );
xor ( n12406 , n12403 , n12404 );
xor ( n12407 , n12314 , n12317 );
and ( n12408 , n831 , n6821 );
and ( n12409 , n12407 , n12408 );
and ( n12410 , n12406 , n12409 );
or ( n12411 , n12405 , n12410 );
and ( n12412 , n12402 , n12411 );
or ( n12413 , n12401 , n12412 );
and ( n12414 , n12398 , n12413 );
or ( n12415 , n12397 , n12414 );
and ( n12416 , n12394 , n12415 );
or ( n12417 , n12393 , n12416 );
and ( n12418 , n12390 , n12417 );
or ( n12419 , n12389 , n12418 );
and ( n12420 , n12386 , n12419 );
or ( n12421 , n12385 , n12420 );
and ( n12422 , n12382 , n12421 );
or ( n12423 , n12381 , n12422 );
and ( n12424 , n12378 , n12423 );
or ( n12425 , n12377 , n12424 );
and ( n12426 , n12374 , n12425 );
or ( n12427 , n12373 , n12426 );
and ( n12428 , n12370 , n12427 );
or ( n12429 , n12369 , n12428 );
and ( n12430 , n12366 , n12429 );
or ( n12431 , n12365 , n12430 );
and ( n12432 , n12362 , n12431 );
or ( n12433 , n12361 , n12432 );
and ( n12434 , n12358 , n12433 );
or ( n12435 , n12357 , n12434 );
and ( n12436 , n12354 , n12435 );
or ( n12437 , n12353 , n12436 );
and ( n12438 , n12350 , n12437 );
or ( n12439 , n12349 , n12438 );
and ( n12440 , n816 , n6818 );
and ( n12441 , n12439 , n12440 );
xor ( n12442 , n12439 , n12440 );
xor ( n12443 , n12350 , n12437 );
and ( n12444 , n817 , n6818 );
and ( n12445 , n12443 , n12444 );
xor ( n12446 , n12443 , n12444 );
xor ( n12447 , n12354 , n12435 );
and ( n12448 , n818 , n6818 );
and ( n12449 , n12447 , n12448 );
xor ( n12450 , n12447 , n12448 );
xor ( n12451 , n12358 , n12433 );
and ( n12452 , n819 , n6818 );
and ( n12453 , n12451 , n12452 );
xor ( n12454 , n12451 , n12452 );
xor ( n12455 , n12362 , n12431 );
and ( n12456 , n820 , n6818 );
and ( n12457 , n12455 , n12456 );
xor ( n12458 , n12455 , n12456 );
xor ( n12459 , n12366 , n12429 );
and ( n12460 , n821 , n6818 );
and ( n12461 , n12459 , n12460 );
xor ( n12462 , n12459 , n12460 );
xor ( n12463 , n12370 , n12427 );
and ( n12464 , n822 , n6818 );
and ( n12465 , n12463 , n12464 );
xor ( n12466 , n12463 , n12464 );
xor ( n12467 , n12374 , n12425 );
and ( n12468 , n823 , n6818 );
and ( n12469 , n12467 , n12468 );
xor ( n12470 , n12467 , n12468 );
xor ( n12471 , n12378 , n12423 );
and ( n12472 , n824 , n6818 );
and ( n12473 , n12471 , n12472 );
xor ( n12474 , n12471 , n12472 );
xor ( n12475 , n12382 , n12421 );
and ( n12476 , n825 , n6818 );
and ( n12477 , n12475 , n12476 );
xor ( n12478 , n12475 , n12476 );
xor ( n12479 , n12386 , n12419 );
and ( n12480 , n826 , n6818 );
and ( n12481 , n12479 , n12480 );
xor ( n12482 , n12479 , n12480 );
xor ( n12483 , n12390 , n12417 );
and ( n12484 , n827 , n6818 );
and ( n12485 , n12483 , n12484 );
xor ( n12486 , n12483 , n12484 );
xor ( n12487 , n12394 , n12415 );
and ( n12488 , n828 , n6818 );
and ( n12489 , n12487 , n12488 );
xor ( n12490 , n12487 , n12488 );
xor ( n12491 , n12398 , n12413 );
and ( n12492 , n829 , n6818 );
and ( n12493 , n12491 , n12492 );
xor ( n12494 , n12491 , n12492 );
xor ( n12495 , n12402 , n12411 );
and ( n12496 , n830 , n6818 );
and ( n12497 , n12495 , n12496 );
xor ( n12498 , n12495 , n12496 );
xor ( n12499 , n12406 , n12409 );
and ( n12500 , n831 , n6818 );
and ( n12501 , n12499 , n12500 );
and ( n12502 , n12498 , n12501 );
or ( n12503 , n12497 , n12502 );
and ( n12504 , n12494 , n12503 );
or ( n12505 , n12493 , n12504 );
and ( n12506 , n12490 , n12505 );
or ( n12507 , n12489 , n12506 );
and ( n12508 , n12486 , n12507 );
or ( n12509 , n12485 , n12508 );
and ( n12510 , n12482 , n12509 );
or ( n12511 , n12481 , n12510 );
and ( n12512 , n12478 , n12511 );
or ( n12513 , n12477 , n12512 );
and ( n12514 , n12474 , n12513 );
or ( n12515 , n12473 , n12514 );
and ( n12516 , n12470 , n12515 );
or ( n12517 , n12469 , n12516 );
and ( n12518 , n12466 , n12517 );
or ( n12519 , n12465 , n12518 );
and ( n12520 , n12462 , n12519 );
or ( n12521 , n12461 , n12520 );
and ( n12522 , n12458 , n12521 );
or ( n12523 , n12457 , n12522 );
and ( n12524 , n12454 , n12523 );
or ( n12525 , n12453 , n12524 );
and ( n12526 , n12450 , n12525 );
or ( n12527 , n12449 , n12526 );
and ( n12528 , n12446 , n12527 );
or ( n12529 , n12445 , n12528 );
and ( n12530 , n12442 , n12529 );
or ( n12531 , n12441 , n12530 );
and ( n12532 , n816 , n6815 );
and ( n12533 , n12531 , n12532 );
xor ( n12534 , n12531 , n12532 );
xor ( n12535 , n12442 , n12529 );
and ( n12536 , n817 , n6815 );
and ( n12537 , n12535 , n12536 );
xor ( n12538 , n12535 , n12536 );
xor ( n12539 , n12446 , n12527 );
and ( n12540 , n818 , n6815 );
and ( n12541 , n12539 , n12540 );
xor ( n12542 , n12539 , n12540 );
xor ( n12543 , n12450 , n12525 );
and ( n12544 , n819 , n6815 );
and ( n12545 , n12543 , n12544 );
xor ( n12546 , n12543 , n12544 );
xor ( n12547 , n12454 , n12523 );
and ( n12548 , n820 , n6815 );
and ( n12549 , n12547 , n12548 );
xor ( n12550 , n12547 , n12548 );
xor ( n12551 , n12458 , n12521 );
and ( n12552 , n821 , n6815 );
and ( n12553 , n12551 , n12552 );
xor ( n12554 , n12551 , n12552 );
xor ( n12555 , n12462 , n12519 );
and ( n12556 , n822 , n6815 );
and ( n12557 , n12555 , n12556 );
xor ( n12558 , n12555 , n12556 );
xor ( n12559 , n12466 , n12517 );
and ( n12560 , n823 , n6815 );
and ( n12561 , n12559 , n12560 );
xor ( n12562 , n12559 , n12560 );
xor ( n12563 , n12470 , n12515 );
and ( n12564 , n824 , n6815 );
and ( n12565 , n12563 , n12564 );
xor ( n12566 , n12563 , n12564 );
xor ( n12567 , n12474 , n12513 );
and ( n12568 , n825 , n6815 );
and ( n12569 , n12567 , n12568 );
xor ( n12570 , n12567 , n12568 );
xor ( n12571 , n12478 , n12511 );
and ( n12572 , n826 , n6815 );
and ( n12573 , n12571 , n12572 );
xor ( n12574 , n12571 , n12572 );
xor ( n12575 , n12482 , n12509 );
and ( n12576 , n827 , n6815 );
and ( n12577 , n12575 , n12576 );
xor ( n12578 , n12575 , n12576 );
xor ( n12579 , n12486 , n12507 );
and ( n12580 , n828 , n6815 );
and ( n12581 , n12579 , n12580 );
xor ( n12582 , n12579 , n12580 );
xor ( n12583 , n12490 , n12505 );
and ( n12584 , n829 , n6815 );
and ( n12585 , n12583 , n12584 );
xor ( n12586 , n12583 , n12584 );
xor ( n12587 , n12494 , n12503 );
and ( n12588 , n830 , n6815 );
and ( n12589 , n12587 , n12588 );
xor ( n12590 , n12587 , n12588 );
xor ( n12591 , n12498 , n12501 );
and ( n12592 , n831 , n6815 );
and ( n12593 , n12591 , n12592 );
and ( n12594 , n12590 , n12593 );
or ( n12595 , n12589 , n12594 );
and ( n12596 , n12586 , n12595 );
or ( n12597 , n12585 , n12596 );
and ( n12598 , n12582 , n12597 );
or ( n12599 , n12581 , n12598 );
and ( n12600 , n12578 , n12599 );
or ( n12601 , n12577 , n12600 );
and ( n12602 , n12574 , n12601 );
or ( n12603 , n12573 , n12602 );
and ( n12604 , n12570 , n12603 );
or ( n12605 , n12569 , n12604 );
and ( n12606 , n12566 , n12605 );
or ( n12607 , n12565 , n12606 );
and ( n12608 , n12562 , n12607 );
or ( n12609 , n12561 , n12608 );
and ( n12610 , n12558 , n12609 );
or ( n12611 , n12557 , n12610 );
and ( n12612 , n12554 , n12611 );
or ( n12613 , n12553 , n12612 );
and ( n12614 , n12550 , n12613 );
or ( n12615 , n12549 , n12614 );
and ( n12616 , n12546 , n12615 );
or ( n12617 , n12545 , n12616 );
and ( n12618 , n12542 , n12617 );
or ( n12619 , n12541 , n12618 );
and ( n12620 , n12538 , n12619 );
or ( n12621 , n12537 , n12620 );
and ( n12622 , n12534 , n12621 );
or ( n12623 , n12533 , n12622 );
and ( n12624 , n816 , n6812 );
and ( n12625 , n12623 , n12624 );
xor ( n12626 , n12623 , n12624 );
xor ( n12627 , n12534 , n12621 );
and ( n12628 , n817 , n6812 );
and ( n12629 , n12627 , n12628 );
xor ( n12630 , n12627 , n12628 );
xor ( n12631 , n12538 , n12619 );
and ( n12632 , n818 , n6812 );
and ( n12633 , n12631 , n12632 );
xor ( n12634 , n12631 , n12632 );
xor ( n12635 , n12542 , n12617 );
and ( n12636 , n819 , n6812 );
and ( n12637 , n12635 , n12636 );
xor ( n12638 , n12635 , n12636 );
xor ( n12639 , n12546 , n12615 );
and ( n12640 , n820 , n6812 );
and ( n12641 , n12639 , n12640 );
xor ( n12642 , n12639 , n12640 );
xor ( n12643 , n12550 , n12613 );
and ( n12644 , n821 , n6812 );
and ( n12645 , n12643 , n12644 );
xor ( n12646 , n12643 , n12644 );
xor ( n12647 , n12554 , n12611 );
and ( n12648 , n822 , n6812 );
and ( n12649 , n12647 , n12648 );
xor ( n12650 , n12647 , n12648 );
xor ( n12651 , n12558 , n12609 );
and ( n12652 , n823 , n6812 );
and ( n12653 , n12651 , n12652 );
xor ( n12654 , n12651 , n12652 );
xor ( n12655 , n12562 , n12607 );
and ( n12656 , n824 , n6812 );
and ( n12657 , n12655 , n12656 );
xor ( n12658 , n12655 , n12656 );
xor ( n12659 , n12566 , n12605 );
and ( n12660 , n825 , n6812 );
and ( n12661 , n12659 , n12660 );
xor ( n12662 , n12659 , n12660 );
xor ( n12663 , n12570 , n12603 );
and ( n12664 , n826 , n6812 );
and ( n12665 , n12663 , n12664 );
xor ( n12666 , n12663 , n12664 );
xor ( n12667 , n12574 , n12601 );
and ( n12668 , n827 , n6812 );
and ( n12669 , n12667 , n12668 );
xor ( n12670 , n12667 , n12668 );
xor ( n12671 , n12578 , n12599 );
and ( n12672 , n828 , n6812 );
and ( n12673 , n12671 , n12672 );
xor ( n12674 , n12671 , n12672 );
xor ( n12675 , n12582 , n12597 );
and ( n12676 , n829 , n6812 );
and ( n12677 , n12675 , n12676 );
xor ( n12678 , n12675 , n12676 );
xor ( n12679 , n12586 , n12595 );
and ( n12680 , n830 , n6812 );
and ( n12681 , n12679 , n12680 );
xor ( n12682 , n12679 , n12680 );
xor ( n12683 , n12590 , n12593 );
and ( n12684 , n831 , n6812 );
and ( n12685 , n12683 , n12684 );
and ( n12686 , n12682 , n12685 );
or ( n12687 , n12681 , n12686 );
and ( n12688 , n12678 , n12687 );
or ( n12689 , n12677 , n12688 );
and ( n12690 , n12674 , n12689 );
or ( n12691 , n12673 , n12690 );
and ( n12692 , n12670 , n12691 );
or ( n12693 , n12669 , n12692 );
and ( n12694 , n12666 , n12693 );
or ( n12695 , n12665 , n12694 );
and ( n12696 , n12662 , n12695 );
or ( n12697 , n12661 , n12696 );
and ( n12698 , n12658 , n12697 );
or ( n12699 , n12657 , n12698 );
and ( n12700 , n12654 , n12699 );
or ( n12701 , n12653 , n12700 );
and ( n12702 , n12650 , n12701 );
or ( n12703 , n12649 , n12702 );
and ( n12704 , n12646 , n12703 );
or ( n12705 , n12645 , n12704 );
and ( n12706 , n12642 , n12705 );
or ( n12707 , n12641 , n12706 );
and ( n12708 , n12638 , n12707 );
or ( n12709 , n12637 , n12708 );
and ( n12710 , n12634 , n12709 );
or ( n12711 , n12633 , n12710 );
and ( n12712 , n12630 , n12711 );
or ( n12713 , n12629 , n12712 );
and ( n12714 , n12626 , n12713 );
or ( n12715 , n12625 , n12714 );
and ( n12716 , n816 , n6809 );
and ( n12717 , n12715 , n12716 );
xor ( n12718 , n12715 , n12716 );
xor ( n12719 , n12626 , n12713 );
and ( n12720 , n817 , n6809 );
and ( n12721 , n12719 , n12720 );
xor ( n12722 , n12719 , n12720 );
xor ( n12723 , n12630 , n12711 );
and ( n12724 , n818 , n6809 );
and ( n12725 , n12723 , n12724 );
xor ( n12726 , n12723 , n12724 );
xor ( n12727 , n12634 , n12709 );
and ( n12728 , n819 , n6809 );
and ( n12729 , n12727 , n12728 );
xor ( n12730 , n12727 , n12728 );
xor ( n12731 , n12638 , n12707 );
and ( n12732 , n820 , n6809 );
and ( n12733 , n12731 , n12732 );
xor ( n12734 , n12731 , n12732 );
xor ( n12735 , n12642 , n12705 );
and ( n12736 , n821 , n6809 );
and ( n12737 , n12735 , n12736 );
xor ( n12738 , n12735 , n12736 );
xor ( n12739 , n12646 , n12703 );
and ( n12740 , n822 , n6809 );
and ( n12741 , n12739 , n12740 );
xor ( n12742 , n12739 , n12740 );
xor ( n12743 , n12650 , n12701 );
and ( n12744 , n823 , n6809 );
and ( n12745 , n12743 , n12744 );
xor ( n12746 , n12743 , n12744 );
xor ( n12747 , n12654 , n12699 );
and ( n12748 , n824 , n6809 );
and ( n12749 , n12747 , n12748 );
xor ( n12750 , n12747 , n12748 );
xor ( n12751 , n12658 , n12697 );
and ( n12752 , n825 , n6809 );
and ( n12753 , n12751 , n12752 );
xor ( n12754 , n12751 , n12752 );
xor ( n12755 , n12662 , n12695 );
and ( n12756 , n826 , n6809 );
and ( n12757 , n12755 , n12756 );
xor ( n12758 , n12755 , n12756 );
xor ( n12759 , n12666 , n12693 );
and ( n12760 , n827 , n6809 );
and ( n12761 , n12759 , n12760 );
xor ( n12762 , n12759 , n12760 );
xor ( n12763 , n12670 , n12691 );
and ( n12764 , n828 , n6809 );
and ( n12765 , n12763 , n12764 );
xor ( n12766 , n12763 , n12764 );
xor ( n12767 , n12674 , n12689 );
and ( n12768 , n829 , n6809 );
and ( n12769 , n12767 , n12768 );
xor ( n12770 , n12767 , n12768 );
xor ( n12771 , n12678 , n12687 );
and ( n12772 , n830 , n6809 );
and ( n12773 , n12771 , n12772 );
xor ( n12774 , n12771 , n12772 );
xor ( n12775 , n12682 , n12685 );
and ( n12776 , n831 , n6809 );
and ( n12777 , n12775 , n12776 );
and ( n12778 , n12774 , n12777 );
or ( n12779 , n12773 , n12778 );
and ( n12780 , n12770 , n12779 );
or ( n12781 , n12769 , n12780 );
and ( n12782 , n12766 , n12781 );
or ( n12783 , n12765 , n12782 );
and ( n12784 , n12762 , n12783 );
or ( n12785 , n12761 , n12784 );
and ( n12786 , n12758 , n12785 );
or ( n12787 , n12757 , n12786 );
and ( n12788 , n12754 , n12787 );
or ( n12789 , n12753 , n12788 );
and ( n12790 , n12750 , n12789 );
or ( n12791 , n12749 , n12790 );
and ( n12792 , n12746 , n12791 );
or ( n12793 , n12745 , n12792 );
and ( n12794 , n12742 , n12793 );
or ( n12795 , n12741 , n12794 );
and ( n12796 , n12738 , n12795 );
or ( n12797 , n12737 , n12796 );
and ( n12798 , n12734 , n12797 );
or ( n12799 , n12733 , n12798 );
and ( n12800 , n12730 , n12799 );
or ( n12801 , n12729 , n12800 );
and ( n12802 , n12726 , n12801 );
or ( n12803 , n12725 , n12802 );
and ( n12804 , n12722 , n12803 );
or ( n12805 , n12721 , n12804 );
and ( n12806 , n12718 , n12805 );
or ( n12807 , n12717 , n12806 );
and ( n12808 , n816 , n6806 );
and ( n12809 , n12807 , n12808 );
xor ( n12810 , n12807 , n12808 );
xor ( n12811 , n12718 , n12805 );
and ( n12812 , n817 , n6806 );
and ( n12813 , n12811 , n12812 );
xor ( n12814 , n12811 , n12812 );
xor ( n12815 , n12722 , n12803 );
and ( n12816 , n818 , n6806 );
and ( n12817 , n12815 , n12816 );
xor ( n12818 , n12815 , n12816 );
xor ( n12819 , n12726 , n12801 );
and ( n12820 , n819 , n6806 );
and ( n12821 , n12819 , n12820 );
xor ( n12822 , n12819 , n12820 );
xor ( n12823 , n12730 , n12799 );
and ( n12824 , n820 , n6806 );
and ( n12825 , n12823 , n12824 );
xor ( n12826 , n12823 , n12824 );
xor ( n12827 , n12734 , n12797 );
and ( n12828 , n821 , n6806 );
and ( n12829 , n12827 , n12828 );
xor ( n12830 , n12827 , n12828 );
xor ( n12831 , n12738 , n12795 );
and ( n12832 , n822 , n6806 );
and ( n12833 , n12831 , n12832 );
xor ( n12834 , n12831 , n12832 );
xor ( n12835 , n12742 , n12793 );
and ( n12836 , n823 , n6806 );
and ( n12837 , n12835 , n12836 );
xor ( n12838 , n12835 , n12836 );
xor ( n12839 , n12746 , n12791 );
and ( n12840 , n824 , n6806 );
and ( n12841 , n12839 , n12840 );
xor ( n12842 , n12839 , n12840 );
xor ( n12843 , n12750 , n12789 );
and ( n12844 , n825 , n6806 );
and ( n12845 , n12843 , n12844 );
xor ( n12846 , n12843 , n12844 );
xor ( n12847 , n12754 , n12787 );
and ( n12848 , n826 , n6806 );
and ( n12849 , n12847 , n12848 );
xor ( n12850 , n12847 , n12848 );
xor ( n12851 , n12758 , n12785 );
and ( n12852 , n827 , n6806 );
and ( n12853 , n12851 , n12852 );
xor ( n12854 , n12851 , n12852 );
xor ( n12855 , n12762 , n12783 );
and ( n12856 , n828 , n6806 );
and ( n12857 , n12855 , n12856 );
xor ( n12858 , n12855 , n12856 );
xor ( n12859 , n12766 , n12781 );
and ( n12860 , n829 , n6806 );
and ( n12861 , n12859 , n12860 );
xor ( n12862 , n12859 , n12860 );
xor ( n12863 , n12770 , n12779 );
and ( n12864 , n830 , n6806 );
and ( n12865 , n12863 , n12864 );
xor ( n12866 , n12863 , n12864 );
xor ( n12867 , n12774 , n12777 );
and ( n12868 , n831 , n6806 );
and ( n12869 , n12867 , n12868 );
and ( n12870 , n12866 , n12869 );
or ( n12871 , n12865 , n12870 );
and ( n12872 , n12862 , n12871 );
or ( n12873 , n12861 , n12872 );
and ( n12874 , n12858 , n12873 );
or ( n12875 , n12857 , n12874 );
and ( n12876 , n12854 , n12875 );
or ( n12877 , n12853 , n12876 );
and ( n12878 , n12850 , n12877 );
or ( n12879 , n12849 , n12878 );
and ( n12880 , n12846 , n12879 );
or ( n12881 , n12845 , n12880 );
and ( n12882 , n12842 , n12881 );
or ( n12883 , n12841 , n12882 );
and ( n12884 , n12838 , n12883 );
or ( n12885 , n12837 , n12884 );
and ( n12886 , n12834 , n12885 );
or ( n12887 , n12833 , n12886 );
and ( n12888 , n12830 , n12887 );
or ( n12889 , n12829 , n12888 );
and ( n12890 , n12826 , n12889 );
or ( n12891 , n12825 , n12890 );
and ( n12892 , n12822 , n12891 );
or ( n12893 , n12821 , n12892 );
and ( n12894 , n12818 , n12893 );
or ( n12895 , n12817 , n12894 );
and ( n12896 , n12814 , n12895 );
or ( n12897 , n12813 , n12896 );
and ( n12898 , n12810 , n12897 );
or ( n12899 , n12809 , n12898 );
and ( n12900 , n816 , n6803 );
and ( n12901 , n12899 , n12900 );
xor ( n12902 , n12899 , n12900 );
xor ( n12903 , n12810 , n12897 );
and ( n12904 , n817 , n6803 );
and ( n12905 , n12903 , n12904 );
xor ( n12906 , n12903 , n12904 );
xor ( n12907 , n12814 , n12895 );
and ( n12908 , n818 , n6803 );
and ( n12909 , n12907 , n12908 );
xor ( n12910 , n12907 , n12908 );
xor ( n12911 , n12818 , n12893 );
and ( n12912 , n819 , n6803 );
and ( n12913 , n12911 , n12912 );
xor ( n12914 , n12911 , n12912 );
xor ( n12915 , n12822 , n12891 );
and ( n12916 , n820 , n6803 );
and ( n12917 , n12915 , n12916 );
xor ( n12918 , n12915 , n12916 );
xor ( n12919 , n12826 , n12889 );
and ( n12920 , n821 , n6803 );
and ( n12921 , n12919 , n12920 );
xor ( n12922 , n12919 , n12920 );
xor ( n12923 , n12830 , n12887 );
and ( n12924 , n822 , n6803 );
and ( n12925 , n12923 , n12924 );
xor ( n12926 , n12923 , n12924 );
xor ( n12927 , n12834 , n12885 );
and ( n12928 , n823 , n6803 );
and ( n12929 , n12927 , n12928 );
xor ( n12930 , n12927 , n12928 );
xor ( n12931 , n12838 , n12883 );
and ( n12932 , n824 , n6803 );
and ( n12933 , n12931 , n12932 );
xor ( n12934 , n12931 , n12932 );
xor ( n12935 , n12842 , n12881 );
and ( n12936 , n825 , n6803 );
and ( n12937 , n12935 , n12936 );
xor ( n12938 , n12935 , n12936 );
xor ( n12939 , n12846 , n12879 );
and ( n12940 , n826 , n6803 );
and ( n12941 , n12939 , n12940 );
xor ( n12942 , n12939 , n12940 );
xor ( n12943 , n12850 , n12877 );
and ( n12944 , n827 , n6803 );
and ( n12945 , n12943 , n12944 );
xor ( n12946 , n12943 , n12944 );
xor ( n12947 , n12854 , n12875 );
and ( n12948 , n828 , n6803 );
and ( n12949 , n12947 , n12948 );
xor ( n12950 , n12947 , n12948 );
xor ( n12951 , n12858 , n12873 );
and ( n12952 , n829 , n6803 );
and ( n12953 , n12951 , n12952 );
xor ( n12954 , n12951 , n12952 );
xor ( n12955 , n12862 , n12871 );
and ( n12956 , n830 , n6803 );
and ( n12957 , n12955 , n12956 );
xor ( n12958 , n12955 , n12956 );
xor ( n12959 , n12866 , n12869 );
and ( n12960 , n831 , n6803 );
and ( n12961 , n12959 , n12960 );
and ( n12962 , n12958 , n12961 );
or ( n12963 , n12957 , n12962 );
and ( n12964 , n12954 , n12963 );
or ( n12965 , n12953 , n12964 );
and ( n12966 , n12950 , n12965 );
or ( n12967 , n12949 , n12966 );
and ( n12968 , n12946 , n12967 );
or ( n12969 , n12945 , n12968 );
and ( n12970 , n12942 , n12969 );
or ( n12971 , n12941 , n12970 );
and ( n12972 , n12938 , n12971 );
or ( n12973 , n12937 , n12972 );
and ( n12974 , n12934 , n12973 );
or ( n12975 , n12933 , n12974 );
and ( n12976 , n12930 , n12975 );
or ( n12977 , n12929 , n12976 );
and ( n12978 , n12926 , n12977 );
or ( n12979 , n12925 , n12978 );
and ( n12980 , n12922 , n12979 );
or ( n12981 , n12921 , n12980 );
and ( n12982 , n12918 , n12981 );
or ( n12983 , n12917 , n12982 );
and ( n12984 , n12914 , n12983 );
or ( n12985 , n12913 , n12984 );
and ( n12986 , n12910 , n12985 );
or ( n12987 , n12909 , n12986 );
and ( n12988 , n12906 , n12987 );
or ( n12989 , n12905 , n12988 );
and ( n12990 , n12902 , n12989 );
or ( n12991 , n12901 , n12990 );
and ( n12992 , n816 , n6800 );
and ( n12993 , n12991 , n12992 );
xor ( n12994 , n12991 , n12992 );
xor ( n12995 , n12902 , n12989 );
and ( n12996 , n817 , n6800 );
and ( n12997 , n12995 , n12996 );
xor ( n12998 , n12995 , n12996 );
xor ( n12999 , n12906 , n12987 );
and ( n13000 , n818 , n6800 );
and ( n13001 , n12999 , n13000 );
xor ( n13002 , n12999 , n13000 );
xor ( n13003 , n12910 , n12985 );
and ( n13004 , n819 , n6800 );
and ( n13005 , n13003 , n13004 );
xor ( n13006 , n13003 , n13004 );
xor ( n13007 , n12914 , n12983 );
and ( n13008 , n820 , n6800 );
and ( n13009 , n13007 , n13008 );
xor ( n13010 , n13007 , n13008 );
xor ( n13011 , n12918 , n12981 );
and ( n13012 , n821 , n6800 );
and ( n13013 , n13011 , n13012 );
xor ( n13014 , n13011 , n13012 );
xor ( n13015 , n12922 , n12979 );
and ( n13016 , n822 , n6800 );
and ( n13017 , n13015 , n13016 );
xor ( n13018 , n13015 , n13016 );
xor ( n13019 , n12926 , n12977 );
and ( n13020 , n823 , n6800 );
and ( n13021 , n13019 , n13020 );
xor ( n13022 , n13019 , n13020 );
xor ( n13023 , n12930 , n12975 );
and ( n13024 , n824 , n6800 );
and ( n13025 , n13023 , n13024 );
xor ( n13026 , n13023 , n13024 );
xor ( n13027 , n12934 , n12973 );
and ( n13028 , n825 , n6800 );
and ( n13029 , n13027 , n13028 );
xor ( n13030 , n13027 , n13028 );
xor ( n13031 , n12938 , n12971 );
and ( n13032 , n826 , n6800 );
and ( n13033 , n13031 , n13032 );
xor ( n13034 , n13031 , n13032 );
xor ( n13035 , n12942 , n12969 );
and ( n13036 , n827 , n6800 );
and ( n13037 , n13035 , n13036 );
xor ( n13038 , n13035 , n13036 );
xor ( n13039 , n12946 , n12967 );
and ( n13040 , n828 , n6800 );
and ( n13041 , n13039 , n13040 );
xor ( n13042 , n13039 , n13040 );
xor ( n13043 , n12950 , n12965 );
and ( n13044 , n829 , n6800 );
and ( n13045 , n13043 , n13044 );
xor ( n13046 , n13043 , n13044 );
xor ( n13047 , n12954 , n12963 );
and ( n13048 , n830 , n6800 );
and ( n13049 , n13047 , n13048 );
xor ( n13050 , n13047 , n13048 );
xor ( n13051 , n12958 , n12961 );
and ( n13052 , n831 , n6800 );
and ( n13053 , n13051 , n13052 );
and ( n13054 , n13050 , n13053 );
or ( n13055 , n13049 , n13054 );
and ( n13056 , n13046 , n13055 );
or ( n13057 , n13045 , n13056 );
and ( n13058 , n13042 , n13057 );
or ( n13059 , n13041 , n13058 );
and ( n13060 , n13038 , n13059 );
or ( n13061 , n13037 , n13060 );
and ( n13062 , n13034 , n13061 );
or ( n13063 , n13033 , n13062 );
and ( n13064 , n13030 , n13063 );
or ( n13065 , n13029 , n13064 );
and ( n13066 , n13026 , n13065 );
or ( n13067 , n13025 , n13066 );
and ( n13068 , n13022 , n13067 );
or ( n13069 , n13021 , n13068 );
and ( n13070 , n13018 , n13069 );
or ( n13071 , n13017 , n13070 );
and ( n13072 , n13014 , n13071 );
or ( n13073 , n13013 , n13072 );
and ( n13074 , n13010 , n13073 );
or ( n13075 , n13009 , n13074 );
and ( n13076 , n13006 , n13075 );
or ( n13077 , n13005 , n13076 );
and ( n13078 , n13002 , n13077 );
or ( n13079 , n13001 , n13078 );
and ( n13080 , n12998 , n13079 );
or ( n13081 , n12997 , n13080 );
and ( n13082 , n12994 , n13081 );
or ( n13083 , n12993 , n13082 );
and ( n13084 , n816 , n6797 );
and ( n13085 , n13083 , n13084 );
xor ( n13086 , n13083 , n13084 );
xor ( n13087 , n12994 , n13081 );
and ( n13088 , n817 , n6797 );
and ( n13089 , n13087 , n13088 );
xor ( n13090 , n13087 , n13088 );
xor ( n13091 , n12998 , n13079 );
and ( n13092 , n818 , n6797 );
and ( n13093 , n13091 , n13092 );
xor ( n13094 , n13091 , n13092 );
xor ( n13095 , n13002 , n13077 );
and ( n13096 , n819 , n6797 );
and ( n13097 , n13095 , n13096 );
xor ( n13098 , n13095 , n13096 );
xor ( n13099 , n13006 , n13075 );
and ( n13100 , n820 , n6797 );
and ( n13101 , n13099 , n13100 );
xor ( n13102 , n13099 , n13100 );
xor ( n13103 , n13010 , n13073 );
and ( n13104 , n821 , n6797 );
and ( n13105 , n13103 , n13104 );
xor ( n13106 , n13103 , n13104 );
xor ( n13107 , n13014 , n13071 );
and ( n13108 , n822 , n6797 );
and ( n13109 , n13107 , n13108 );
xor ( n13110 , n13107 , n13108 );
xor ( n13111 , n13018 , n13069 );
and ( n13112 , n823 , n6797 );
and ( n13113 , n13111 , n13112 );
xor ( n13114 , n13111 , n13112 );
xor ( n13115 , n13022 , n13067 );
and ( n13116 , n824 , n6797 );
and ( n13117 , n13115 , n13116 );
xor ( n13118 , n13115 , n13116 );
xor ( n13119 , n13026 , n13065 );
and ( n13120 , n825 , n6797 );
and ( n13121 , n13119 , n13120 );
xor ( n13122 , n13119 , n13120 );
xor ( n13123 , n13030 , n13063 );
and ( n13124 , n826 , n6797 );
and ( n13125 , n13123 , n13124 );
xor ( n13126 , n13123 , n13124 );
xor ( n13127 , n13034 , n13061 );
and ( n13128 , n827 , n6797 );
and ( n13129 , n13127 , n13128 );
xor ( n13130 , n13127 , n13128 );
xor ( n13131 , n13038 , n13059 );
and ( n13132 , n828 , n6797 );
and ( n13133 , n13131 , n13132 );
xor ( n13134 , n13131 , n13132 );
xor ( n13135 , n13042 , n13057 );
and ( n13136 , n829 , n6797 );
and ( n13137 , n13135 , n13136 );
xor ( n13138 , n13135 , n13136 );
xor ( n13139 , n13046 , n13055 );
and ( n13140 , n830 , n6797 );
and ( n13141 , n13139 , n13140 );
xor ( n13142 , n13139 , n13140 );
xor ( n13143 , n13050 , n13053 );
and ( n13144 , n831 , n6797 );
and ( n13145 , n13143 , n13144 );
and ( n13146 , n13142 , n13145 );
or ( n13147 , n13141 , n13146 );
and ( n13148 , n13138 , n13147 );
or ( n13149 , n13137 , n13148 );
and ( n13150 , n13134 , n13149 );
or ( n13151 , n13133 , n13150 );
and ( n13152 , n13130 , n13151 );
or ( n13153 , n13129 , n13152 );
and ( n13154 , n13126 , n13153 );
or ( n13155 , n13125 , n13154 );
and ( n13156 , n13122 , n13155 );
or ( n13157 , n13121 , n13156 );
and ( n13158 , n13118 , n13157 );
or ( n13159 , n13117 , n13158 );
and ( n13160 , n13114 , n13159 );
or ( n13161 , n13113 , n13160 );
and ( n13162 , n13110 , n13161 );
or ( n13163 , n13109 , n13162 );
and ( n13164 , n13106 , n13163 );
or ( n13165 , n13105 , n13164 );
and ( n13166 , n13102 , n13165 );
or ( n13167 , n13101 , n13166 );
and ( n13168 , n13098 , n13167 );
or ( n13169 , n13097 , n13168 );
and ( n13170 , n13094 , n13169 );
or ( n13171 , n13093 , n13170 );
and ( n13172 , n13090 , n13171 );
or ( n13173 , n13089 , n13172 );
and ( n13174 , n13086 , n13173 );
or ( n13175 , n13085 , n13174 );
and ( n13176 , n816 , n6794 );
and ( n13177 , n13175 , n13176 );
xor ( n13178 , n13175 , n13176 );
xor ( n13179 , n13086 , n13173 );
and ( n13180 , n817 , n6794 );
and ( n13181 , n13179 , n13180 );
xor ( n13182 , n13179 , n13180 );
xor ( n13183 , n13090 , n13171 );
and ( n13184 , n818 , n6794 );
and ( n13185 , n13183 , n13184 );
xor ( n13186 , n13183 , n13184 );
xor ( n13187 , n13094 , n13169 );
and ( n13188 , n819 , n6794 );
and ( n13189 , n13187 , n13188 );
xor ( n13190 , n13187 , n13188 );
xor ( n13191 , n13098 , n13167 );
and ( n13192 , n820 , n6794 );
and ( n13193 , n13191 , n13192 );
xor ( n13194 , n13191 , n13192 );
xor ( n13195 , n13102 , n13165 );
and ( n13196 , n821 , n6794 );
and ( n13197 , n13195 , n13196 );
xor ( n13198 , n13195 , n13196 );
xor ( n13199 , n13106 , n13163 );
and ( n13200 , n822 , n6794 );
and ( n13201 , n13199 , n13200 );
xor ( n13202 , n13199 , n13200 );
xor ( n13203 , n13110 , n13161 );
and ( n13204 , n823 , n6794 );
and ( n13205 , n13203 , n13204 );
xor ( n13206 , n13203 , n13204 );
xor ( n13207 , n13114 , n13159 );
and ( n13208 , n824 , n6794 );
and ( n13209 , n13207 , n13208 );
xor ( n13210 , n13207 , n13208 );
xor ( n13211 , n13118 , n13157 );
and ( n13212 , n825 , n6794 );
and ( n13213 , n13211 , n13212 );
xor ( n13214 , n13211 , n13212 );
xor ( n13215 , n13122 , n13155 );
and ( n13216 , n826 , n6794 );
and ( n13217 , n13215 , n13216 );
xor ( n13218 , n13215 , n13216 );
xor ( n13219 , n13126 , n13153 );
and ( n13220 , n827 , n6794 );
and ( n13221 , n13219 , n13220 );
xor ( n13222 , n13219 , n13220 );
xor ( n13223 , n13130 , n13151 );
and ( n13224 , n828 , n6794 );
and ( n13225 , n13223 , n13224 );
xor ( n13226 , n13223 , n13224 );
xor ( n13227 , n13134 , n13149 );
and ( n13228 , n829 , n6794 );
and ( n13229 , n13227 , n13228 );
xor ( n13230 , n13227 , n13228 );
xor ( n13231 , n13138 , n13147 );
and ( n13232 , n830 , n6794 );
and ( n13233 , n13231 , n13232 );
xor ( n13234 , n13231 , n13232 );
xor ( n13235 , n13142 , n13145 );
and ( n13236 , n831 , n6794 );
and ( n13237 , n13235 , n13236 );
and ( n13238 , n13234 , n13237 );
or ( n13239 , n13233 , n13238 );
and ( n13240 , n13230 , n13239 );
or ( n13241 , n13229 , n13240 );
and ( n13242 , n13226 , n13241 );
or ( n13243 , n13225 , n13242 );
and ( n13244 , n13222 , n13243 );
or ( n13245 , n13221 , n13244 );
and ( n13246 , n13218 , n13245 );
or ( n13247 , n13217 , n13246 );
and ( n13248 , n13214 , n13247 );
or ( n13249 , n13213 , n13248 );
and ( n13250 , n13210 , n13249 );
or ( n13251 , n13209 , n13250 );
and ( n13252 , n13206 , n13251 );
or ( n13253 , n13205 , n13252 );
and ( n13254 , n13202 , n13253 );
or ( n13255 , n13201 , n13254 );
and ( n13256 , n13198 , n13255 );
or ( n13257 , n13197 , n13256 );
and ( n13258 , n13194 , n13257 );
or ( n13259 , n13193 , n13258 );
and ( n13260 , n13190 , n13259 );
or ( n13261 , n13189 , n13260 );
and ( n13262 , n13186 , n13261 );
or ( n13263 , n13185 , n13262 );
and ( n13264 , n13182 , n13263 );
or ( n13265 , n13181 , n13264 );
and ( n13266 , n13178 , n13265 );
or ( n13267 , n13177 , n13266 );
and ( n13268 , n816 , n6791 );
and ( n13269 , n13267 , n13268 );
xor ( n13270 , n13267 , n13268 );
xor ( n13271 , n13178 , n13265 );
and ( n13272 , n817 , n6791 );
and ( n13273 , n13271 , n13272 );
xor ( n13274 , n13271 , n13272 );
xor ( n13275 , n13182 , n13263 );
and ( n13276 , n818 , n6791 );
and ( n13277 , n13275 , n13276 );
xor ( n13278 , n13275 , n13276 );
xor ( n13279 , n13186 , n13261 );
and ( n13280 , n819 , n6791 );
and ( n13281 , n13279 , n13280 );
xor ( n13282 , n13279 , n13280 );
xor ( n13283 , n13190 , n13259 );
and ( n13284 , n820 , n6791 );
and ( n13285 , n13283 , n13284 );
xor ( n13286 , n13283 , n13284 );
xor ( n13287 , n13194 , n13257 );
and ( n13288 , n821 , n6791 );
and ( n13289 , n13287 , n13288 );
xor ( n13290 , n13287 , n13288 );
xor ( n13291 , n13198 , n13255 );
and ( n13292 , n822 , n6791 );
and ( n13293 , n13291 , n13292 );
xor ( n13294 , n13291 , n13292 );
xor ( n13295 , n13202 , n13253 );
and ( n13296 , n823 , n6791 );
and ( n13297 , n13295 , n13296 );
xor ( n13298 , n13295 , n13296 );
xor ( n13299 , n13206 , n13251 );
and ( n13300 , n824 , n6791 );
and ( n13301 , n13299 , n13300 );
xor ( n13302 , n13299 , n13300 );
xor ( n13303 , n13210 , n13249 );
and ( n13304 , n825 , n6791 );
and ( n13305 , n13303 , n13304 );
xor ( n13306 , n13303 , n13304 );
xor ( n13307 , n13214 , n13247 );
and ( n13308 , n826 , n6791 );
and ( n13309 , n13307 , n13308 );
xor ( n13310 , n13307 , n13308 );
xor ( n13311 , n13218 , n13245 );
and ( n13312 , n827 , n6791 );
and ( n13313 , n13311 , n13312 );
xor ( n13314 , n13311 , n13312 );
xor ( n13315 , n13222 , n13243 );
and ( n13316 , n828 , n6791 );
and ( n13317 , n13315 , n13316 );
xor ( n13318 , n13315 , n13316 );
xor ( n13319 , n13226 , n13241 );
and ( n13320 , n829 , n6791 );
and ( n13321 , n13319 , n13320 );
xor ( n13322 , n13319 , n13320 );
xor ( n13323 , n13230 , n13239 );
and ( n13324 , n830 , n6791 );
and ( n13325 , n13323 , n13324 );
xor ( n13326 , n13323 , n13324 );
xor ( n13327 , n13234 , n13237 );
and ( n13328 , n831 , n6791 );
and ( n13329 , n13327 , n13328 );
and ( n13330 , n13326 , n13329 );
or ( n13331 , n13325 , n13330 );
and ( n13332 , n13322 , n13331 );
or ( n13333 , n13321 , n13332 );
and ( n13334 , n13318 , n13333 );
or ( n13335 , n13317 , n13334 );
and ( n13336 , n13314 , n13335 );
or ( n13337 , n13313 , n13336 );
and ( n13338 , n13310 , n13337 );
or ( n13339 , n13309 , n13338 );
and ( n13340 , n13306 , n13339 );
or ( n13341 , n13305 , n13340 );
and ( n13342 , n13302 , n13341 );
or ( n13343 , n13301 , n13342 );
and ( n13344 , n13298 , n13343 );
or ( n13345 , n13297 , n13344 );
and ( n13346 , n13294 , n13345 );
or ( n13347 , n13293 , n13346 );
and ( n13348 , n13290 , n13347 );
or ( n13349 , n13289 , n13348 );
and ( n13350 , n13286 , n13349 );
or ( n13351 , n13285 , n13350 );
and ( n13352 , n13282 , n13351 );
or ( n13353 , n13281 , n13352 );
and ( n13354 , n13278 , n13353 );
or ( n13355 , n13277 , n13354 );
and ( n13356 , n13274 , n13355 );
or ( n13357 , n13273 , n13356 );
and ( n13358 , n13270 , n13357 );
or ( n13359 , n13269 , n13358 );
and ( n13360 , n816 , n6788 );
and ( n13361 , n13359 , n13360 );
xor ( n13362 , n13359 , n13360 );
xor ( n13363 , n13270 , n13357 );
and ( n13364 , n817 , n6788 );
and ( n13365 , n13363 , n13364 );
xor ( n13366 , n13363 , n13364 );
xor ( n13367 , n13274 , n13355 );
and ( n13368 , n818 , n6788 );
and ( n13369 , n13367 , n13368 );
xor ( n13370 , n13367 , n13368 );
xor ( n13371 , n13278 , n13353 );
and ( n13372 , n819 , n6788 );
and ( n13373 , n13371 , n13372 );
xor ( n13374 , n13371 , n13372 );
xor ( n13375 , n13282 , n13351 );
and ( n13376 , n820 , n6788 );
and ( n13377 , n13375 , n13376 );
xor ( n13378 , n13375 , n13376 );
xor ( n13379 , n13286 , n13349 );
and ( n13380 , n821 , n6788 );
and ( n13381 , n13379 , n13380 );
xor ( n13382 , n13379 , n13380 );
xor ( n13383 , n13290 , n13347 );
and ( n13384 , n822 , n6788 );
and ( n13385 , n13383 , n13384 );
xor ( n13386 , n13383 , n13384 );
xor ( n13387 , n13294 , n13345 );
and ( n13388 , n823 , n6788 );
and ( n13389 , n13387 , n13388 );
xor ( n13390 , n13387 , n13388 );
xor ( n13391 , n13298 , n13343 );
and ( n13392 , n824 , n6788 );
and ( n13393 , n13391 , n13392 );
xor ( n13394 , n13391 , n13392 );
xor ( n13395 , n13302 , n13341 );
and ( n13396 , n825 , n6788 );
and ( n13397 , n13395 , n13396 );
xor ( n13398 , n13395 , n13396 );
xor ( n13399 , n13306 , n13339 );
and ( n13400 , n826 , n6788 );
and ( n13401 , n13399 , n13400 );
xor ( n13402 , n13399 , n13400 );
xor ( n13403 , n13310 , n13337 );
and ( n13404 , n827 , n6788 );
and ( n13405 , n13403 , n13404 );
xor ( n13406 , n13403 , n13404 );
xor ( n13407 , n13314 , n13335 );
and ( n13408 , n828 , n6788 );
and ( n13409 , n13407 , n13408 );
xor ( n13410 , n13407 , n13408 );
xor ( n13411 , n13318 , n13333 );
and ( n13412 , n829 , n6788 );
and ( n13413 , n13411 , n13412 );
xor ( n13414 , n13411 , n13412 );
xor ( n13415 , n13322 , n13331 );
and ( n13416 , n830 , n6788 );
and ( n13417 , n13415 , n13416 );
xor ( n13418 , n13415 , n13416 );
xor ( n13419 , n13326 , n13329 );
and ( n13420 , n831 , n6788 );
and ( n13421 , n13419 , n13420 );
and ( n13422 , n13418 , n13421 );
or ( n13423 , n13417 , n13422 );
and ( n13424 , n13414 , n13423 );
or ( n13425 , n13413 , n13424 );
and ( n13426 , n13410 , n13425 );
or ( n13427 , n13409 , n13426 );
and ( n13428 , n13406 , n13427 );
or ( n13429 , n13405 , n13428 );
and ( n13430 , n13402 , n13429 );
or ( n13431 , n13401 , n13430 );
and ( n13432 , n13398 , n13431 );
or ( n13433 , n13397 , n13432 );
and ( n13434 , n13394 , n13433 );
or ( n13435 , n13393 , n13434 );
and ( n13436 , n13390 , n13435 );
or ( n13437 , n13389 , n13436 );
and ( n13438 , n13386 , n13437 );
or ( n13439 , n13385 , n13438 );
and ( n13440 , n13382 , n13439 );
or ( n13441 , n13381 , n13440 );
and ( n13442 , n13378 , n13441 );
or ( n13443 , n13377 , n13442 );
and ( n13444 , n13374 , n13443 );
or ( n13445 , n13373 , n13444 );
and ( n13446 , n13370 , n13445 );
or ( n13447 , n13369 , n13446 );
and ( n13448 , n13366 , n13447 );
or ( n13449 , n13365 , n13448 );
and ( n13450 , n13362 , n13449 );
or ( n13451 , n13361 , n13450 );
and ( n13452 , n816 , n6785 );
and ( n13453 , n13451 , n13452 );
xor ( n13454 , n13451 , n13452 );
xor ( n13455 , n13362 , n13449 );
and ( n13456 , n817 , n6785 );
and ( n13457 , n13455 , n13456 );
xor ( n13458 , n13455 , n13456 );
xor ( n13459 , n13366 , n13447 );
and ( n13460 , n818 , n6785 );
and ( n13461 , n13459 , n13460 );
xor ( n13462 , n13459 , n13460 );
xor ( n13463 , n13370 , n13445 );
and ( n13464 , n819 , n6785 );
and ( n13465 , n13463 , n13464 );
xor ( n13466 , n13463 , n13464 );
xor ( n13467 , n13374 , n13443 );
and ( n13468 , n820 , n6785 );
and ( n13469 , n13467 , n13468 );
xor ( n13470 , n13467 , n13468 );
xor ( n13471 , n13378 , n13441 );
and ( n13472 , n821 , n6785 );
and ( n13473 , n13471 , n13472 );
xor ( n13474 , n13471 , n13472 );
xor ( n13475 , n13382 , n13439 );
and ( n13476 , n822 , n6785 );
and ( n13477 , n13475 , n13476 );
xor ( n13478 , n13475 , n13476 );
xor ( n13479 , n13386 , n13437 );
and ( n13480 , n823 , n6785 );
and ( n13481 , n13479 , n13480 );
xor ( n13482 , n13479 , n13480 );
xor ( n13483 , n13390 , n13435 );
and ( n13484 , n824 , n6785 );
and ( n13485 , n13483 , n13484 );
xor ( n13486 , n13483 , n13484 );
xor ( n13487 , n13394 , n13433 );
and ( n13488 , n825 , n6785 );
and ( n13489 , n13487 , n13488 );
xor ( n13490 , n13487 , n13488 );
xor ( n13491 , n13398 , n13431 );
and ( n13492 , n826 , n6785 );
and ( n13493 , n13491 , n13492 );
xor ( n13494 , n13491 , n13492 );
xor ( n13495 , n13402 , n13429 );
and ( n13496 , n827 , n6785 );
and ( n13497 , n13495 , n13496 );
xor ( n13498 , n13495 , n13496 );
xor ( n13499 , n13406 , n13427 );
and ( n13500 , n828 , n6785 );
and ( n13501 , n13499 , n13500 );
xor ( n13502 , n13499 , n13500 );
xor ( n13503 , n13410 , n13425 );
and ( n13504 , n829 , n6785 );
and ( n13505 , n13503 , n13504 );
xor ( n13506 , n13503 , n13504 );
xor ( n13507 , n13414 , n13423 );
and ( n13508 , n830 , n6785 );
and ( n13509 , n13507 , n13508 );
xor ( n13510 , n13507 , n13508 );
xor ( n13511 , n13418 , n13421 );
and ( n13512 , n831 , n6785 );
and ( n13513 , n13511 , n13512 );
and ( n13514 , n13510 , n13513 );
or ( n13515 , n13509 , n13514 );
and ( n13516 , n13506 , n13515 );
or ( n13517 , n13505 , n13516 );
and ( n13518 , n13502 , n13517 );
or ( n13519 , n13501 , n13518 );
and ( n13520 , n13498 , n13519 );
or ( n13521 , n13497 , n13520 );
and ( n13522 , n13494 , n13521 );
or ( n13523 , n13493 , n13522 );
and ( n13524 , n13490 , n13523 );
or ( n13525 , n13489 , n13524 );
and ( n13526 , n13486 , n13525 );
or ( n13527 , n13485 , n13526 );
and ( n13528 , n13482 , n13527 );
or ( n13529 , n13481 , n13528 );
and ( n13530 , n13478 , n13529 );
or ( n13531 , n13477 , n13530 );
and ( n13532 , n13474 , n13531 );
or ( n13533 , n13473 , n13532 );
and ( n13534 , n13470 , n13533 );
or ( n13535 , n13469 , n13534 );
and ( n13536 , n13466 , n13535 );
or ( n13537 , n13465 , n13536 );
and ( n13538 , n13462 , n13537 );
or ( n13539 , n13461 , n13538 );
and ( n13540 , n13458 , n13539 );
or ( n13541 , n13457 , n13540 );
and ( n13542 , n13454 , n13541 );
or ( n13543 , n13453 , n13542 );
and ( n13544 , n816 , n6782 );
and ( n13545 , n13543 , n13544 );
xor ( n13546 , n13543 , n13544 );
xor ( n13547 , n13454 , n13541 );
and ( n13548 , n817 , n6782 );
and ( n13549 , n13547 , n13548 );
xor ( n13550 , n13547 , n13548 );
xor ( n13551 , n13458 , n13539 );
and ( n13552 , n818 , n6782 );
and ( n13553 , n13551 , n13552 );
xor ( n13554 , n13551 , n13552 );
xor ( n13555 , n13462 , n13537 );
and ( n13556 , n819 , n6782 );
and ( n13557 , n13555 , n13556 );
xor ( n13558 , n13555 , n13556 );
xor ( n13559 , n13466 , n13535 );
and ( n13560 , n820 , n6782 );
and ( n13561 , n13559 , n13560 );
xor ( n13562 , n13559 , n13560 );
xor ( n13563 , n13470 , n13533 );
and ( n13564 , n821 , n6782 );
and ( n13565 , n13563 , n13564 );
xor ( n13566 , n13563 , n13564 );
xor ( n13567 , n13474 , n13531 );
and ( n13568 , n822 , n6782 );
and ( n13569 , n13567 , n13568 );
xor ( n13570 , n13567 , n13568 );
xor ( n13571 , n13478 , n13529 );
and ( n13572 , n823 , n6782 );
and ( n13573 , n13571 , n13572 );
xor ( n13574 , n13571 , n13572 );
xor ( n13575 , n13482 , n13527 );
and ( n13576 , n824 , n6782 );
and ( n13577 , n13575 , n13576 );
xor ( n13578 , n13575 , n13576 );
xor ( n13579 , n13486 , n13525 );
and ( n13580 , n825 , n6782 );
and ( n13581 , n13579 , n13580 );
xor ( n13582 , n13579 , n13580 );
xor ( n13583 , n13490 , n13523 );
and ( n13584 , n826 , n6782 );
and ( n13585 , n13583 , n13584 );
xor ( n13586 , n13583 , n13584 );
xor ( n13587 , n13494 , n13521 );
and ( n13588 , n827 , n6782 );
and ( n13589 , n13587 , n13588 );
xor ( n13590 , n13587 , n13588 );
xor ( n13591 , n13498 , n13519 );
and ( n13592 , n828 , n6782 );
and ( n13593 , n13591 , n13592 );
xor ( n13594 , n13591 , n13592 );
xor ( n13595 , n13502 , n13517 );
and ( n13596 , n829 , n6782 );
and ( n13597 , n13595 , n13596 );
xor ( n13598 , n13595 , n13596 );
xor ( n13599 , n13506 , n13515 );
and ( n13600 , n830 , n6782 );
and ( n13601 , n13599 , n13600 );
xor ( n13602 , n13599 , n13600 );
xor ( n13603 , n13510 , n13513 );
and ( n13604 , n831 , n6782 );
and ( n13605 , n13603 , n13604 );
and ( n13606 , n13602 , n13605 );
or ( n13607 , n13601 , n13606 );
and ( n13608 , n13598 , n13607 );
or ( n13609 , n13597 , n13608 );
and ( n13610 , n13594 , n13609 );
or ( n13611 , n13593 , n13610 );
and ( n13612 , n13590 , n13611 );
or ( n13613 , n13589 , n13612 );
and ( n13614 , n13586 , n13613 );
or ( n13615 , n13585 , n13614 );
and ( n13616 , n13582 , n13615 );
or ( n13617 , n13581 , n13616 );
and ( n13618 , n13578 , n13617 );
or ( n13619 , n13577 , n13618 );
and ( n13620 , n13574 , n13619 );
or ( n13621 , n13573 , n13620 );
and ( n13622 , n13570 , n13621 );
or ( n13623 , n13569 , n13622 );
and ( n13624 , n13566 , n13623 );
or ( n13625 , n13565 , n13624 );
and ( n13626 , n13562 , n13625 );
or ( n13627 , n13561 , n13626 );
and ( n13628 , n13558 , n13627 );
or ( n13629 , n13557 , n13628 );
and ( n13630 , n13554 , n13629 );
or ( n13631 , n13553 , n13630 );
and ( n13632 , n13550 , n13631 );
or ( n13633 , n13549 , n13632 );
and ( n13634 , n13546 , n13633 );
or ( n13635 , n13545 , n13634 );
and ( n13636 , n816 , n6779 );
and ( n13637 , n13635 , n13636 );
xor ( n13638 , n13635 , n13636 );
xor ( n13639 , n13546 , n13633 );
and ( n13640 , n817 , n6779 );
and ( n13641 , n13639 , n13640 );
xor ( n13642 , n13639 , n13640 );
xor ( n13643 , n13550 , n13631 );
and ( n13644 , n818 , n6779 );
and ( n13645 , n13643 , n13644 );
xor ( n13646 , n13643 , n13644 );
xor ( n13647 , n13554 , n13629 );
and ( n13648 , n819 , n6779 );
and ( n13649 , n13647 , n13648 );
xor ( n13650 , n13647 , n13648 );
xor ( n13651 , n13558 , n13627 );
and ( n13652 , n820 , n6779 );
and ( n13653 , n13651 , n13652 );
xor ( n13654 , n13651 , n13652 );
xor ( n13655 , n13562 , n13625 );
and ( n13656 , n821 , n6779 );
and ( n13657 , n13655 , n13656 );
xor ( n13658 , n13655 , n13656 );
xor ( n13659 , n13566 , n13623 );
and ( n13660 , n822 , n6779 );
and ( n13661 , n13659 , n13660 );
xor ( n13662 , n13659 , n13660 );
xor ( n13663 , n13570 , n13621 );
and ( n13664 , n823 , n6779 );
and ( n13665 , n13663 , n13664 );
xor ( n13666 , n13663 , n13664 );
xor ( n13667 , n13574 , n13619 );
and ( n13668 , n824 , n6779 );
and ( n13669 , n13667 , n13668 );
xor ( n13670 , n13667 , n13668 );
xor ( n13671 , n13578 , n13617 );
and ( n13672 , n825 , n6779 );
and ( n13673 , n13671 , n13672 );
xor ( n13674 , n13671 , n13672 );
xor ( n13675 , n13582 , n13615 );
and ( n13676 , n826 , n6779 );
and ( n13677 , n13675 , n13676 );
xor ( n13678 , n13675 , n13676 );
xor ( n13679 , n13586 , n13613 );
and ( n13680 , n827 , n6779 );
and ( n13681 , n13679 , n13680 );
xor ( n13682 , n13679 , n13680 );
xor ( n13683 , n13590 , n13611 );
and ( n13684 , n828 , n6779 );
and ( n13685 , n13683 , n13684 );
xor ( n13686 , n13683 , n13684 );
xor ( n13687 , n13594 , n13609 );
and ( n13688 , n829 , n6779 );
and ( n13689 , n13687 , n13688 );
xor ( n13690 , n13687 , n13688 );
xor ( n13691 , n13598 , n13607 );
and ( n13692 , n830 , n6779 );
and ( n13693 , n13691 , n13692 );
xor ( n13694 , n13691 , n13692 );
xor ( n13695 , n13602 , n13605 );
and ( n13696 , n831 , n6779 );
and ( n13697 , n13695 , n13696 );
and ( n13698 , n13694 , n13697 );
or ( n13699 , n13693 , n13698 );
and ( n13700 , n13690 , n13699 );
or ( n13701 , n13689 , n13700 );
and ( n13702 , n13686 , n13701 );
or ( n13703 , n13685 , n13702 );
and ( n13704 , n13682 , n13703 );
or ( n13705 , n13681 , n13704 );
and ( n13706 , n13678 , n13705 );
or ( n13707 , n13677 , n13706 );
and ( n13708 , n13674 , n13707 );
or ( n13709 , n13673 , n13708 );
and ( n13710 , n13670 , n13709 );
or ( n13711 , n13669 , n13710 );
and ( n13712 , n13666 , n13711 );
or ( n13713 , n13665 , n13712 );
and ( n13714 , n13662 , n13713 );
or ( n13715 , n13661 , n13714 );
and ( n13716 , n13658 , n13715 );
or ( n13717 , n13657 , n13716 );
and ( n13718 , n13654 , n13717 );
or ( n13719 , n13653 , n13718 );
and ( n13720 , n13650 , n13719 );
or ( n13721 , n13649 , n13720 );
and ( n13722 , n13646 , n13721 );
or ( n13723 , n13645 , n13722 );
and ( n13724 , n13642 , n13723 );
or ( n13725 , n13641 , n13724 );
and ( n13726 , n13638 , n13725 );
or ( n13727 , n13637 , n13726 );
and ( n13728 , n816 , n6776 );
and ( n13729 , n13727 , n13728 );
xor ( n13730 , n13727 , n13728 );
xor ( n13731 , n13638 , n13725 );
and ( n13732 , n817 , n6776 );
and ( n13733 , n13731 , n13732 );
xor ( n13734 , n13731 , n13732 );
xor ( n13735 , n13642 , n13723 );
and ( n13736 , n818 , n6776 );
and ( n13737 , n13735 , n13736 );
xor ( n13738 , n13735 , n13736 );
xor ( n13739 , n13646 , n13721 );
and ( n13740 , n819 , n6776 );
and ( n13741 , n13739 , n13740 );
xor ( n13742 , n13739 , n13740 );
xor ( n13743 , n13650 , n13719 );
and ( n13744 , n820 , n6776 );
and ( n13745 , n13743 , n13744 );
xor ( n13746 , n13743 , n13744 );
xor ( n13747 , n13654 , n13717 );
and ( n13748 , n821 , n6776 );
and ( n13749 , n13747 , n13748 );
xor ( n13750 , n13747 , n13748 );
xor ( n13751 , n13658 , n13715 );
and ( n13752 , n822 , n6776 );
and ( n13753 , n13751 , n13752 );
xor ( n13754 , n13751 , n13752 );
xor ( n13755 , n13662 , n13713 );
and ( n13756 , n823 , n6776 );
and ( n13757 , n13755 , n13756 );
xor ( n13758 , n13755 , n13756 );
xor ( n13759 , n13666 , n13711 );
and ( n13760 , n824 , n6776 );
and ( n13761 , n13759 , n13760 );
xor ( n13762 , n13759 , n13760 );
xor ( n13763 , n13670 , n13709 );
and ( n13764 , n825 , n6776 );
and ( n13765 , n13763 , n13764 );
xor ( n13766 , n13763 , n13764 );
xor ( n13767 , n13674 , n13707 );
and ( n13768 , n826 , n6776 );
and ( n13769 , n13767 , n13768 );
xor ( n13770 , n13767 , n13768 );
xor ( n13771 , n13678 , n13705 );
and ( n13772 , n827 , n6776 );
and ( n13773 , n13771 , n13772 );
xor ( n13774 , n13771 , n13772 );
xor ( n13775 , n13682 , n13703 );
and ( n13776 , n828 , n6776 );
and ( n13777 , n13775 , n13776 );
xor ( n13778 , n13775 , n13776 );
xor ( n13779 , n13686 , n13701 );
and ( n13780 , n829 , n6776 );
and ( n13781 , n13779 , n13780 );
xor ( n13782 , n13779 , n13780 );
xor ( n13783 , n13690 , n13699 );
and ( n13784 , n830 , n6776 );
and ( n13785 , n13783 , n13784 );
xor ( n13786 , n13783 , n13784 );
xor ( n13787 , n13694 , n13697 );
and ( n13788 , n831 , n6776 );
and ( n13789 , n13787 , n13788 );
and ( n13790 , n13786 , n13789 );
or ( n13791 , n13785 , n13790 );
and ( n13792 , n13782 , n13791 );
or ( n13793 , n13781 , n13792 );
and ( n13794 , n13778 , n13793 );
or ( n13795 , n13777 , n13794 );
and ( n13796 , n13774 , n13795 );
or ( n13797 , n13773 , n13796 );
and ( n13798 , n13770 , n13797 );
or ( n13799 , n13769 , n13798 );
and ( n13800 , n13766 , n13799 );
or ( n13801 , n13765 , n13800 );
and ( n13802 , n13762 , n13801 );
or ( n13803 , n13761 , n13802 );
and ( n13804 , n13758 , n13803 );
or ( n13805 , n13757 , n13804 );
and ( n13806 , n13754 , n13805 );
or ( n13807 , n13753 , n13806 );
and ( n13808 , n13750 , n13807 );
or ( n13809 , n13749 , n13808 );
and ( n13810 , n13746 , n13809 );
or ( n13811 , n13745 , n13810 );
and ( n13812 , n13742 , n13811 );
or ( n13813 , n13741 , n13812 );
and ( n13814 , n13738 , n13813 );
or ( n13815 , n13737 , n13814 );
and ( n13816 , n13734 , n13815 );
or ( n13817 , n13733 , n13816 );
and ( n13818 , n13730 , n13817 );
or ( n13819 , n13729 , n13818 );
and ( n13820 , n816 , n6773 );
and ( n13821 , n13819 , n13820 );
xor ( n13822 , n13819 , n13820 );
xor ( n13823 , n13730 , n13817 );
and ( n13824 , n817 , n6773 );
and ( n13825 , n13823 , n13824 );
xor ( n13826 , n13823 , n13824 );
xor ( n13827 , n13734 , n13815 );
and ( n13828 , n818 , n6773 );
and ( n13829 , n13827 , n13828 );
xor ( n13830 , n13827 , n13828 );
xor ( n13831 , n13738 , n13813 );
and ( n13832 , n819 , n6773 );
and ( n13833 , n13831 , n13832 );
xor ( n13834 , n13831 , n13832 );
xor ( n13835 , n13742 , n13811 );
and ( n13836 , n820 , n6773 );
and ( n13837 , n13835 , n13836 );
xor ( n13838 , n13835 , n13836 );
xor ( n13839 , n13746 , n13809 );
and ( n13840 , n821 , n6773 );
and ( n13841 , n13839 , n13840 );
xor ( n13842 , n13839 , n13840 );
xor ( n13843 , n13750 , n13807 );
and ( n13844 , n822 , n6773 );
and ( n13845 , n13843 , n13844 );
xor ( n13846 , n13843 , n13844 );
xor ( n13847 , n13754 , n13805 );
and ( n13848 , n823 , n6773 );
and ( n13849 , n13847 , n13848 );
xor ( n13850 , n13847 , n13848 );
xor ( n13851 , n13758 , n13803 );
and ( n13852 , n824 , n6773 );
and ( n13853 , n13851 , n13852 );
xor ( n13854 , n13851 , n13852 );
xor ( n13855 , n13762 , n13801 );
and ( n13856 , n825 , n6773 );
and ( n13857 , n13855 , n13856 );
xor ( n13858 , n13855 , n13856 );
xor ( n13859 , n13766 , n13799 );
and ( n13860 , n826 , n6773 );
and ( n13861 , n13859 , n13860 );
xor ( n13862 , n13859 , n13860 );
xor ( n13863 , n13770 , n13797 );
and ( n13864 , n827 , n6773 );
and ( n13865 , n13863 , n13864 );
xor ( n13866 , n13863 , n13864 );
xor ( n13867 , n13774 , n13795 );
and ( n13868 , n828 , n6773 );
and ( n13869 , n13867 , n13868 );
xor ( n13870 , n13867 , n13868 );
xor ( n13871 , n13778 , n13793 );
and ( n13872 , n829 , n6773 );
and ( n13873 , n13871 , n13872 );
xor ( n13874 , n13871 , n13872 );
xor ( n13875 , n13782 , n13791 );
and ( n13876 , n830 , n6773 );
and ( n13877 , n13875 , n13876 );
xor ( n13878 , n13875 , n13876 );
xor ( n13879 , n13786 , n13789 );
and ( n13880 , n831 , n6773 );
and ( n13881 , n13879 , n13880 );
and ( n13882 , n13878 , n13881 );
or ( n13883 , n13877 , n13882 );
and ( n13884 , n13874 , n13883 );
or ( n13885 , n13873 , n13884 );
and ( n13886 , n13870 , n13885 );
or ( n13887 , n13869 , n13886 );
and ( n13888 , n13866 , n13887 );
or ( n13889 , n13865 , n13888 );
and ( n13890 , n13862 , n13889 );
or ( n13891 , n13861 , n13890 );
and ( n13892 , n13858 , n13891 );
or ( n13893 , n13857 , n13892 );
and ( n13894 , n13854 , n13893 );
or ( n13895 , n13853 , n13894 );
and ( n13896 , n13850 , n13895 );
or ( n13897 , n13849 , n13896 );
and ( n13898 , n13846 , n13897 );
or ( n13899 , n13845 , n13898 );
and ( n13900 , n13842 , n13899 );
or ( n13901 , n13841 , n13900 );
and ( n13902 , n13838 , n13901 );
or ( n13903 , n13837 , n13902 );
and ( n13904 , n13834 , n13903 );
or ( n13905 , n13833 , n13904 );
and ( n13906 , n13830 , n13905 );
or ( n13907 , n13829 , n13906 );
and ( n13908 , n13826 , n13907 );
or ( n13909 , n13825 , n13908 );
and ( n13910 , n13822 , n13909 );
or ( n13911 , n13821 , n13910 );
and ( n13912 , n816 , n6770 );
and ( n13913 , n13911 , n13912 );
xor ( n13914 , n13911 , n13912 );
xor ( n13915 , n13822 , n13909 );
and ( n13916 , n817 , n6770 );
and ( n13917 , n13915 , n13916 );
xor ( n13918 , n13915 , n13916 );
xor ( n13919 , n13826 , n13907 );
and ( n13920 , n818 , n6770 );
and ( n13921 , n13919 , n13920 );
xor ( n13922 , n13919 , n13920 );
xor ( n13923 , n13830 , n13905 );
and ( n13924 , n819 , n6770 );
and ( n13925 , n13923 , n13924 );
xor ( n13926 , n13923 , n13924 );
xor ( n13927 , n13834 , n13903 );
and ( n13928 , n820 , n6770 );
and ( n13929 , n13927 , n13928 );
xor ( n13930 , n13927 , n13928 );
xor ( n13931 , n13838 , n13901 );
and ( n13932 , n821 , n6770 );
and ( n13933 , n13931 , n13932 );
xor ( n13934 , n13931 , n13932 );
xor ( n13935 , n13842 , n13899 );
and ( n13936 , n822 , n6770 );
and ( n13937 , n13935 , n13936 );
xor ( n13938 , n13935 , n13936 );
xor ( n13939 , n13846 , n13897 );
and ( n13940 , n823 , n6770 );
and ( n13941 , n13939 , n13940 );
xor ( n13942 , n13939 , n13940 );
xor ( n13943 , n13850 , n13895 );
and ( n13944 , n824 , n6770 );
and ( n13945 , n13943 , n13944 );
xor ( n13946 , n13943 , n13944 );
xor ( n13947 , n13854 , n13893 );
and ( n13948 , n825 , n6770 );
and ( n13949 , n13947 , n13948 );
xor ( n13950 , n13947 , n13948 );
xor ( n13951 , n13858 , n13891 );
and ( n13952 , n826 , n6770 );
and ( n13953 , n13951 , n13952 );
xor ( n13954 , n13951 , n13952 );
xor ( n13955 , n13862 , n13889 );
and ( n13956 , n827 , n6770 );
and ( n13957 , n13955 , n13956 );
xor ( n13958 , n13955 , n13956 );
xor ( n13959 , n13866 , n13887 );
and ( n13960 , n828 , n6770 );
and ( n13961 , n13959 , n13960 );
xor ( n13962 , n13959 , n13960 );
xor ( n13963 , n13870 , n13885 );
and ( n13964 , n829 , n6770 );
and ( n13965 , n13963 , n13964 );
xor ( n13966 , n13963 , n13964 );
xor ( n13967 , n13874 , n13883 );
and ( n13968 , n830 , n6770 );
and ( n13969 , n13967 , n13968 );
xor ( n13970 , n13967 , n13968 );
xor ( n13971 , n13878 , n13881 );
and ( n13972 , n831 , n6770 );
and ( n13973 , n13971 , n13972 );
and ( n13974 , n13970 , n13973 );
or ( n13975 , n13969 , n13974 );
and ( n13976 , n13966 , n13975 );
or ( n13977 , n13965 , n13976 );
and ( n13978 , n13962 , n13977 );
or ( n13979 , n13961 , n13978 );
and ( n13980 , n13958 , n13979 );
or ( n13981 , n13957 , n13980 );
and ( n13982 , n13954 , n13981 );
or ( n13983 , n13953 , n13982 );
and ( n13984 , n13950 , n13983 );
or ( n13985 , n13949 , n13984 );
and ( n13986 , n13946 , n13985 );
or ( n13987 , n13945 , n13986 );
and ( n13988 , n13942 , n13987 );
or ( n13989 , n13941 , n13988 );
and ( n13990 , n13938 , n13989 );
or ( n13991 , n13937 , n13990 );
and ( n13992 , n13934 , n13991 );
or ( n13993 , n13933 , n13992 );
and ( n13994 , n13930 , n13993 );
or ( n13995 , n13929 , n13994 );
and ( n13996 , n13926 , n13995 );
or ( n13997 , n13925 , n13996 );
and ( n13998 , n13922 , n13997 );
or ( n13999 , n13921 , n13998 );
and ( n14000 , n13918 , n13999 );
or ( n14001 , n13917 , n14000 );
and ( n14002 , n13914 , n14001 );
or ( n14003 , n13913 , n14002 );
and ( n14004 , n816 , n6767 );
and ( n14005 , n14003 , n14004 );
xor ( n14006 , n14003 , n14004 );
xor ( n14007 , n13914 , n14001 );
and ( n14008 , n817 , n6767 );
and ( n14009 , n14007 , n14008 );
xor ( n14010 , n14007 , n14008 );
xor ( n14011 , n13918 , n13999 );
and ( n14012 , n818 , n6767 );
and ( n14013 , n14011 , n14012 );
xor ( n14014 , n14011 , n14012 );
xor ( n14015 , n13922 , n13997 );
and ( n14016 , n819 , n6767 );
and ( n14017 , n14015 , n14016 );
xor ( n14018 , n14015 , n14016 );
xor ( n14019 , n13926 , n13995 );
and ( n14020 , n820 , n6767 );
and ( n14021 , n14019 , n14020 );
xor ( n14022 , n14019 , n14020 );
xor ( n14023 , n13930 , n13993 );
and ( n14024 , n821 , n6767 );
and ( n14025 , n14023 , n14024 );
xor ( n14026 , n14023 , n14024 );
xor ( n14027 , n13934 , n13991 );
and ( n14028 , n822 , n6767 );
and ( n14029 , n14027 , n14028 );
xor ( n14030 , n14027 , n14028 );
xor ( n14031 , n13938 , n13989 );
and ( n14032 , n823 , n6767 );
and ( n14033 , n14031 , n14032 );
xor ( n14034 , n14031 , n14032 );
xor ( n14035 , n13942 , n13987 );
and ( n14036 , n824 , n6767 );
and ( n14037 , n14035 , n14036 );
xor ( n14038 , n14035 , n14036 );
xor ( n14039 , n13946 , n13985 );
and ( n14040 , n825 , n6767 );
and ( n14041 , n14039 , n14040 );
xor ( n14042 , n14039 , n14040 );
xor ( n14043 , n13950 , n13983 );
and ( n14044 , n826 , n6767 );
and ( n14045 , n14043 , n14044 );
xor ( n14046 , n14043 , n14044 );
xor ( n14047 , n13954 , n13981 );
and ( n14048 , n827 , n6767 );
and ( n14049 , n14047 , n14048 );
xor ( n14050 , n14047 , n14048 );
xor ( n14051 , n13958 , n13979 );
and ( n14052 , n828 , n6767 );
and ( n14053 , n14051 , n14052 );
xor ( n14054 , n14051 , n14052 );
xor ( n14055 , n13962 , n13977 );
and ( n14056 , n829 , n6767 );
and ( n14057 , n14055 , n14056 );
xor ( n14058 , n14055 , n14056 );
xor ( n14059 , n13966 , n13975 );
and ( n14060 , n830 , n6767 );
and ( n14061 , n14059 , n14060 );
xor ( n14062 , n14059 , n14060 );
xor ( n14063 , n13970 , n13973 );
and ( n14064 , n831 , n6767 );
and ( n14065 , n14063 , n14064 );
and ( n14066 , n14062 , n14065 );
or ( n14067 , n14061 , n14066 );
and ( n14068 , n14058 , n14067 );
or ( n14069 , n14057 , n14068 );
and ( n14070 , n14054 , n14069 );
or ( n14071 , n14053 , n14070 );
and ( n14072 , n14050 , n14071 );
or ( n14073 , n14049 , n14072 );
and ( n14074 , n14046 , n14073 );
or ( n14075 , n14045 , n14074 );
and ( n14076 , n14042 , n14075 );
or ( n14077 , n14041 , n14076 );
and ( n14078 , n14038 , n14077 );
or ( n14079 , n14037 , n14078 );
and ( n14080 , n14034 , n14079 );
or ( n14081 , n14033 , n14080 );
and ( n14082 , n14030 , n14081 );
or ( n14083 , n14029 , n14082 );
and ( n14084 , n14026 , n14083 );
or ( n14085 , n14025 , n14084 );
and ( n14086 , n14022 , n14085 );
or ( n14087 , n14021 , n14086 );
and ( n14088 , n14018 , n14087 );
or ( n14089 , n14017 , n14088 );
and ( n14090 , n14014 , n14089 );
or ( n14091 , n14013 , n14090 );
and ( n14092 , n14010 , n14091 );
or ( n14093 , n14009 , n14092 );
and ( n14094 , n14006 , n14093 );
or ( n14095 , n14005 , n14094 );
and ( n14096 , n816 , n6764 );
and ( n14097 , n14095 , n14096 );
xor ( n14098 , n14095 , n14096 );
xor ( n14099 , n14006 , n14093 );
and ( n14100 , n817 , n6764 );
and ( n14101 , n14099 , n14100 );
xor ( n14102 , n14099 , n14100 );
xor ( n14103 , n14010 , n14091 );
and ( n14104 , n818 , n6764 );
and ( n14105 , n14103 , n14104 );
xor ( n14106 , n14103 , n14104 );
xor ( n14107 , n14014 , n14089 );
and ( n14108 , n819 , n6764 );
and ( n14109 , n14107 , n14108 );
xor ( n14110 , n14107 , n14108 );
xor ( n14111 , n14018 , n14087 );
and ( n14112 , n820 , n6764 );
and ( n14113 , n14111 , n14112 );
xor ( n14114 , n14111 , n14112 );
xor ( n14115 , n14022 , n14085 );
and ( n14116 , n821 , n6764 );
and ( n14117 , n14115 , n14116 );
xor ( n14118 , n14115 , n14116 );
xor ( n14119 , n14026 , n14083 );
and ( n14120 , n822 , n6764 );
and ( n14121 , n14119 , n14120 );
xor ( n14122 , n14119 , n14120 );
xor ( n14123 , n14030 , n14081 );
and ( n14124 , n823 , n6764 );
and ( n14125 , n14123 , n14124 );
xor ( n14126 , n14123 , n14124 );
xor ( n14127 , n14034 , n14079 );
and ( n14128 , n824 , n6764 );
and ( n14129 , n14127 , n14128 );
xor ( n14130 , n14127 , n14128 );
xor ( n14131 , n14038 , n14077 );
and ( n14132 , n825 , n6764 );
and ( n14133 , n14131 , n14132 );
xor ( n14134 , n14131 , n14132 );
xor ( n14135 , n14042 , n14075 );
and ( n14136 , n826 , n6764 );
and ( n14137 , n14135 , n14136 );
xor ( n14138 , n14135 , n14136 );
xor ( n14139 , n14046 , n14073 );
and ( n14140 , n827 , n6764 );
and ( n14141 , n14139 , n14140 );
xor ( n14142 , n14139 , n14140 );
xor ( n14143 , n14050 , n14071 );
and ( n14144 , n828 , n6764 );
and ( n14145 , n14143 , n14144 );
xor ( n14146 , n14143 , n14144 );
xor ( n14147 , n14054 , n14069 );
and ( n14148 , n829 , n6764 );
and ( n14149 , n14147 , n14148 );
xor ( n14150 , n14147 , n14148 );
xor ( n14151 , n14058 , n14067 );
and ( n14152 , n830 , n6764 );
and ( n14153 , n14151 , n14152 );
xor ( n14154 , n14151 , n14152 );
xor ( n14155 , n14062 , n14065 );
and ( n14156 , n831 , n6764 );
and ( n14157 , n14155 , n14156 );
and ( n14158 , n14154 , n14157 );
or ( n14159 , n14153 , n14158 );
and ( n14160 , n14150 , n14159 );
or ( n14161 , n14149 , n14160 );
and ( n14162 , n14146 , n14161 );
or ( n14163 , n14145 , n14162 );
and ( n14164 , n14142 , n14163 );
or ( n14165 , n14141 , n14164 );
and ( n14166 , n14138 , n14165 );
or ( n14167 , n14137 , n14166 );
and ( n14168 , n14134 , n14167 );
or ( n14169 , n14133 , n14168 );
and ( n14170 , n14130 , n14169 );
or ( n14171 , n14129 , n14170 );
and ( n14172 , n14126 , n14171 );
or ( n14173 , n14125 , n14172 );
and ( n14174 , n14122 , n14173 );
or ( n14175 , n14121 , n14174 );
and ( n14176 , n14118 , n14175 );
or ( n14177 , n14117 , n14176 );
and ( n14178 , n14114 , n14177 );
or ( n14179 , n14113 , n14178 );
and ( n14180 , n14110 , n14179 );
or ( n14181 , n14109 , n14180 );
and ( n14182 , n14106 , n14181 );
or ( n14183 , n14105 , n14182 );
and ( n14184 , n14102 , n14183 );
or ( n14185 , n14101 , n14184 );
and ( n14186 , n14098 , n14185 );
or ( n14187 , n14097 , n14186 );
and ( n14188 , n816 , n6761 );
and ( n14189 , n14187 , n14188 );
xor ( n14190 , n14187 , n14188 );
xor ( n14191 , n14098 , n14185 );
and ( n14192 , n817 , n6761 );
and ( n14193 , n14191 , n14192 );
xor ( n14194 , n14191 , n14192 );
xor ( n14195 , n14102 , n14183 );
and ( n14196 , n818 , n6761 );
and ( n14197 , n14195 , n14196 );
xor ( n14198 , n14195 , n14196 );
xor ( n14199 , n14106 , n14181 );
and ( n14200 , n819 , n6761 );
and ( n14201 , n14199 , n14200 );
xor ( n14202 , n14199 , n14200 );
xor ( n14203 , n14110 , n14179 );
and ( n14204 , n820 , n6761 );
and ( n14205 , n14203 , n14204 );
xor ( n14206 , n14203 , n14204 );
xor ( n14207 , n14114 , n14177 );
and ( n14208 , n821 , n6761 );
and ( n14209 , n14207 , n14208 );
xor ( n14210 , n14207 , n14208 );
xor ( n14211 , n14118 , n14175 );
and ( n14212 , n822 , n6761 );
and ( n14213 , n14211 , n14212 );
xor ( n14214 , n14211 , n14212 );
xor ( n14215 , n14122 , n14173 );
and ( n14216 , n823 , n6761 );
and ( n14217 , n14215 , n14216 );
xor ( n14218 , n14215 , n14216 );
xor ( n14219 , n14126 , n14171 );
and ( n14220 , n824 , n6761 );
and ( n14221 , n14219 , n14220 );
xor ( n14222 , n14219 , n14220 );
xor ( n14223 , n14130 , n14169 );
and ( n14224 , n825 , n6761 );
and ( n14225 , n14223 , n14224 );
xor ( n14226 , n14223 , n14224 );
xor ( n14227 , n14134 , n14167 );
and ( n14228 , n826 , n6761 );
and ( n14229 , n14227 , n14228 );
xor ( n14230 , n14227 , n14228 );
xor ( n14231 , n14138 , n14165 );
and ( n14232 , n827 , n6761 );
and ( n14233 , n14231 , n14232 );
xor ( n14234 , n14231 , n14232 );
xor ( n14235 , n14142 , n14163 );
and ( n14236 , n828 , n6761 );
and ( n14237 , n14235 , n14236 );
xor ( n14238 , n14235 , n14236 );
xor ( n14239 , n14146 , n14161 );
and ( n14240 , n829 , n6761 );
and ( n14241 , n14239 , n14240 );
xor ( n14242 , n14239 , n14240 );
xor ( n14243 , n14150 , n14159 );
and ( n14244 , n830 , n6761 );
and ( n14245 , n14243 , n14244 );
xor ( n14246 , n14243 , n14244 );
xor ( n14247 , n14154 , n14157 );
and ( n14248 , n831 , n6761 );
and ( n14249 , n14247 , n14248 );
and ( n14250 , n14246 , n14249 );
or ( n14251 , n14245 , n14250 );
and ( n14252 , n14242 , n14251 );
or ( n14253 , n14241 , n14252 );
and ( n14254 , n14238 , n14253 );
or ( n14255 , n14237 , n14254 );
and ( n14256 , n14234 , n14255 );
or ( n14257 , n14233 , n14256 );
and ( n14258 , n14230 , n14257 );
or ( n14259 , n14229 , n14258 );
and ( n14260 , n14226 , n14259 );
or ( n14261 , n14225 , n14260 );
and ( n14262 , n14222 , n14261 );
or ( n14263 , n14221 , n14262 );
and ( n14264 , n14218 , n14263 );
or ( n14265 , n14217 , n14264 );
and ( n14266 , n14214 , n14265 );
or ( n14267 , n14213 , n14266 );
and ( n14268 , n14210 , n14267 );
or ( n14269 , n14209 , n14268 );
and ( n14270 , n14206 , n14269 );
or ( n14271 , n14205 , n14270 );
and ( n14272 , n14202 , n14271 );
or ( n14273 , n14201 , n14272 );
and ( n14274 , n14198 , n14273 );
or ( n14275 , n14197 , n14274 );
and ( n14276 , n14194 , n14275 );
or ( n14277 , n14193 , n14276 );
and ( n14278 , n14190 , n14277 );
or ( n14279 , n14189 , n14278 );
and ( n14280 , n816 , n6758 );
and ( n14281 , n14279 , n14280 );
xor ( n14282 , n14279 , n14280 );
xor ( n14283 , n14190 , n14277 );
and ( n14284 , n817 , n6758 );
and ( n14285 , n14283 , n14284 );
xor ( n14286 , n14283 , n14284 );
xor ( n14287 , n14194 , n14275 );
and ( n14288 , n818 , n6758 );
and ( n14289 , n14287 , n14288 );
xor ( n14290 , n14287 , n14288 );
xor ( n14291 , n14198 , n14273 );
and ( n14292 , n819 , n6758 );
and ( n14293 , n14291 , n14292 );
xor ( n14294 , n14291 , n14292 );
xor ( n14295 , n14202 , n14271 );
and ( n14296 , n820 , n6758 );
and ( n14297 , n14295 , n14296 );
xor ( n14298 , n14295 , n14296 );
xor ( n14299 , n14206 , n14269 );
and ( n14300 , n821 , n6758 );
and ( n14301 , n14299 , n14300 );
xor ( n14302 , n14299 , n14300 );
xor ( n14303 , n14210 , n14267 );
and ( n14304 , n822 , n6758 );
and ( n14305 , n14303 , n14304 );
xor ( n14306 , n14303 , n14304 );
xor ( n14307 , n14214 , n14265 );
and ( n14308 , n823 , n6758 );
and ( n14309 , n14307 , n14308 );
xor ( n14310 , n14307 , n14308 );
xor ( n14311 , n14218 , n14263 );
and ( n14312 , n824 , n6758 );
and ( n14313 , n14311 , n14312 );
xor ( n14314 , n14311 , n14312 );
xor ( n14315 , n14222 , n14261 );
and ( n14316 , n825 , n6758 );
and ( n14317 , n14315 , n14316 );
xor ( n14318 , n14315 , n14316 );
xor ( n14319 , n14226 , n14259 );
and ( n14320 , n826 , n6758 );
and ( n14321 , n14319 , n14320 );
xor ( n14322 , n14319 , n14320 );
xor ( n14323 , n14230 , n14257 );
and ( n14324 , n827 , n6758 );
and ( n14325 , n14323 , n14324 );
xor ( n14326 , n14323 , n14324 );
xor ( n14327 , n14234 , n14255 );
and ( n14328 , n828 , n6758 );
and ( n14329 , n14327 , n14328 );
xor ( n14330 , n14327 , n14328 );
xor ( n14331 , n14238 , n14253 );
and ( n14332 , n829 , n6758 );
and ( n14333 , n14331 , n14332 );
xor ( n14334 , n14331 , n14332 );
xor ( n14335 , n14242 , n14251 );
and ( n14336 , n830 , n6758 );
and ( n14337 , n14335 , n14336 );
xor ( n14338 , n14335 , n14336 );
xor ( n14339 , n14246 , n14249 );
and ( n14340 , n831 , n6758 );
and ( n14341 , n14339 , n14340 );
and ( n14342 , n14338 , n14341 );
or ( n14343 , n14337 , n14342 );
and ( n14344 , n14334 , n14343 );
or ( n14345 , n14333 , n14344 );
and ( n14346 , n14330 , n14345 );
or ( n14347 , n14329 , n14346 );
and ( n14348 , n14326 , n14347 );
or ( n14349 , n14325 , n14348 );
and ( n14350 , n14322 , n14349 );
or ( n14351 , n14321 , n14350 );
and ( n14352 , n14318 , n14351 );
or ( n14353 , n14317 , n14352 );
and ( n14354 , n14314 , n14353 );
or ( n14355 , n14313 , n14354 );
and ( n14356 , n14310 , n14355 );
or ( n14357 , n14309 , n14356 );
and ( n14358 , n14306 , n14357 );
or ( n14359 , n14305 , n14358 );
and ( n14360 , n14302 , n14359 );
or ( n14361 , n14301 , n14360 );
and ( n14362 , n14298 , n14361 );
or ( n14363 , n14297 , n14362 );
and ( n14364 , n14294 , n14363 );
or ( n14365 , n14293 , n14364 );
and ( n14366 , n14290 , n14365 );
or ( n14367 , n14289 , n14366 );
and ( n14368 , n14286 , n14367 );
or ( n14369 , n14285 , n14368 );
and ( n14370 , n14282 , n14369 );
or ( n14371 , n14281 , n14370 );
and ( n14372 , n816 , n6755 );
and ( n14373 , n14371 , n14372 );
xor ( n14374 , n14371 , n14372 );
xor ( n14375 , n14282 , n14369 );
and ( n14376 , n817 , n6755 );
and ( n14377 , n14375 , n14376 );
xor ( n14378 , n14375 , n14376 );
xor ( n14379 , n14286 , n14367 );
and ( n14380 , n818 , n6755 );
and ( n14381 , n14379 , n14380 );
xor ( n14382 , n14379 , n14380 );
xor ( n14383 , n14290 , n14365 );
and ( n14384 , n819 , n6755 );
and ( n14385 , n14383 , n14384 );
xor ( n14386 , n14383 , n14384 );
xor ( n14387 , n14294 , n14363 );
and ( n14388 , n820 , n6755 );
and ( n14389 , n14387 , n14388 );
xor ( n14390 , n14387 , n14388 );
xor ( n14391 , n14298 , n14361 );
and ( n14392 , n821 , n6755 );
and ( n14393 , n14391 , n14392 );
xor ( n14394 , n14391 , n14392 );
xor ( n14395 , n14302 , n14359 );
and ( n14396 , n822 , n6755 );
and ( n14397 , n14395 , n14396 );
xor ( n14398 , n14395 , n14396 );
xor ( n14399 , n14306 , n14357 );
and ( n14400 , n823 , n6755 );
and ( n14401 , n14399 , n14400 );
xor ( n14402 , n14399 , n14400 );
xor ( n14403 , n14310 , n14355 );
and ( n14404 , n824 , n6755 );
and ( n14405 , n14403 , n14404 );
xor ( n14406 , n14403 , n14404 );
xor ( n14407 , n14314 , n14353 );
and ( n14408 , n825 , n6755 );
and ( n14409 , n14407 , n14408 );
xor ( n14410 , n14407 , n14408 );
xor ( n14411 , n14318 , n14351 );
and ( n14412 , n826 , n6755 );
and ( n14413 , n14411 , n14412 );
xor ( n14414 , n14411 , n14412 );
xor ( n14415 , n14322 , n14349 );
and ( n14416 , n827 , n6755 );
and ( n14417 , n14415 , n14416 );
xor ( n14418 , n14415 , n14416 );
xor ( n14419 , n14326 , n14347 );
and ( n14420 , n828 , n6755 );
and ( n14421 , n14419 , n14420 );
xor ( n14422 , n14419 , n14420 );
xor ( n14423 , n14330 , n14345 );
and ( n14424 , n829 , n6755 );
and ( n14425 , n14423 , n14424 );
xor ( n14426 , n14423 , n14424 );
xor ( n14427 , n14334 , n14343 );
and ( n14428 , n830 , n6755 );
and ( n14429 , n14427 , n14428 );
xor ( n14430 , n14427 , n14428 );
xor ( n14431 , n14338 , n14341 );
and ( n14432 , n831 , n6755 );
and ( n14433 , n14431 , n14432 );
and ( n14434 , n14430 , n14433 );
or ( n14435 , n14429 , n14434 );
and ( n14436 , n14426 , n14435 );
or ( n14437 , n14425 , n14436 );
and ( n14438 , n14422 , n14437 );
or ( n14439 , n14421 , n14438 );
and ( n14440 , n14418 , n14439 );
or ( n14441 , n14417 , n14440 );
and ( n14442 , n14414 , n14441 );
or ( n14443 , n14413 , n14442 );
and ( n14444 , n14410 , n14443 );
or ( n14445 , n14409 , n14444 );
and ( n14446 , n14406 , n14445 );
or ( n14447 , n14405 , n14446 );
and ( n14448 , n14402 , n14447 );
or ( n14449 , n14401 , n14448 );
and ( n14450 , n14398 , n14449 );
or ( n14451 , n14397 , n14450 );
and ( n14452 , n14394 , n14451 );
or ( n14453 , n14393 , n14452 );
and ( n14454 , n14390 , n14453 );
or ( n14455 , n14389 , n14454 );
and ( n14456 , n14386 , n14455 );
or ( n14457 , n14385 , n14456 );
and ( n14458 , n14382 , n14457 );
or ( n14459 , n14381 , n14458 );
and ( n14460 , n14378 , n14459 );
or ( n14461 , n14377 , n14460 );
and ( n14462 , n14374 , n14461 );
or ( n14463 , n14373 , n14462 );
and ( n14464 , n816 , n6752 );
and ( n14465 , n14463 , n14464 );
xor ( n14466 , n14463 , n14464 );
xor ( n14467 , n14374 , n14461 );
and ( n14468 , n817 , n6752 );
and ( n14469 , n14467 , n14468 );
xor ( n14470 , n14467 , n14468 );
xor ( n14471 , n14378 , n14459 );
and ( n14472 , n818 , n6752 );
and ( n14473 , n14471 , n14472 );
xor ( n14474 , n14471 , n14472 );
xor ( n14475 , n14382 , n14457 );
and ( n14476 , n819 , n6752 );
and ( n14477 , n14475 , n14476 );
xor ( n14478 , n14475 , n14476 );
xor ( n14479 , n14386 , n14455 );
and ( n14480 , n820 , n6752 );
and ( n14481 , n14479 , n14480 );
xor ( n14482 , n14479 , n14480 );
xor ( n14483 , n14390 , n14453 );
and ( n14484 , n821 , n6752 );
and ( n14485 , n14483 , n14484 );
xor ( n14486 , n14483 , n14484 );
xor ( n14487 , n14394 , n14451 );
and ( n14488 , n822 , n6752 );
and ( n14489 , n14487 , n14488 );
xor ( n14490 , n14487 , n14488 );
xor ( n14491 , n14398 , n14449 );
and ( n14492 , n823 , n6752 );
and ( n14493 , n14491 , n14492 );
xor ( n14494 , n14491 , n14492 );
xor ( n14495 , n14402 , n14447 );
and ( n14496 , n824 , n6752 );
and ( n14497 , n14495 , n14496 );
xor ( n14498 , n14495 , n14496 );
xor ( n14499 , n14406 , n14445 );
and ( n14500 , n825 , n6752 );
and ( n14501 , n14499 , n14500 );
xor ( n14502 , n14499 , n14500 );
xor ( n14503 , n14410 , n14443 );
and ( n14504 , n826 , n6752 );
and ( n14505 , n14503 , n14504 );
xor ( n14506 , n14503 , n14504 );
xor ( n14507 , n14414 , n14441 );
and ( n14508 , n827 , n6752 );
and ( n14509 , n14507 , n14508 );
xor ( n14510 , n14507 , n14508 );
xor ( n14511 , n14418 , n14439 );
and ( n14512 , n828 , n6752 );
and ( n14513 , n14511 , n14512 );
xor ( n14514 , n14511 , n14512 );
xor ( n14515 , n14422 , n14437 );
and ( n14516 , n829 , n6752 );
and ( n14517 , n14515 , n14516 );
xor ( n14518 , n14515 , n14516 );
xor ( n14519 , n14426 , n14435 );
and ( n14520 , n830 , n6752 );
and ( n14521 , n14519 , n14520 );
xor ( n14522 , n14519 , n14520 );
xor ( n14523 , n14430 , n14433 );
and ( n14524 , n831 , n6752 );
and ( n14525 , n14523 , n14524 );
and ( n14526 , n14522 , n14525 );
or ( n14527 , n14521 , n14526 );
and ( n14528 , n14518 , n14527 );
or ( n14529 , n14517 , n14528 );
and ( n14530 , n14514 , n14529 );
or ( n14531 , n14513 , n14530 );
and ( n14532 , n14510 , n14531 );
or ( n14533 , n14509 , n14532 );
and ( n14534 , n14506 , n14533 );
or ( n14535 , n14505 , n14534 );
and ( n14536 , n14502 , n14535 );
or ( n14537 , n14501 , n14536 );
and ( n14538 , n14498 , n14537 );
or ( n14539 , n14497 , n14538 );
and ( n14540 , n14494 , n14539 );
or ( n14541 , n14493 , n14540 );
and ( n14542 , n14490 , n14541 );
or ( n14543 , n14489 , n14542 );
and ( n14544 , n14486 , n14543 );
or ( n14545 , n14485 , n14544 );
and ( n14546 , n14482 , n14545 );
or ( n14547 , n14481 , n14546 );
and ( n14548 , n14478 , n14547 );
or ( n14549 , n14477 , n14548 );
and ( n14550 , n14474 , n14549 );
or ( n14551 , n14473 , n14550 );
and ( n14552 , n14470 , n14551 );
or ( n14553 , n14469 , n14552 );
and ( n14554 , n14466 , n14553 );
or ( n14555 , n14465 , n14554 );
and ( n14556 , n816 , n6749 );
and ( n14557 , n14555 , n14556 );
xor ( n14558 , n14555 , n14556 );
xor ( n14559 , n14466 , n14553 );
and ( n14560 , n817 , n6749 );
and ( n14561 , n14559 , n14560 );
xor ( n14562 , n14559 , n14560 );
xor ( n14563 , n14470 , n14551 );
and ( n14564 , n818 , n6749 );
and ( n14565 , n14563 , n14564 );
xor ( n14566 , n14563 , n14564 );
xor ( n14567 , n14474 , n14549 );
and ( n14568 , n819 , n6749 );
and ( n14569 , n14567 , n14568 );
xor ( n14570 , n14567 , n14568 );
xor ( n14571 , n14478 , n14547 );
and ( n14572 , n820 , n6749 );
and ( n14573 , n14571 , n14572 );
xor ( n14574 , n14571 , n14572 );
xor ( n14575 , n14482 , n14545 );
and ( n14576 , n821 , n6749 );
and ( n14577 , n14575 , n14576 );
xor ( n14578 , n14575 , n14576 );
xor ( n14579 , n14486 , n14543 );
and ( n14580 , n822 , n6749 );
and ( n14581 , n14579 , n14580 );
xor ( n14582 , n14579 , n14580 );
xor ( n14583 , n14490 , n14541 );
and ( n14584 , n823 , n6749 );
and ( n14585 , n14583 , n14584 );
xor ( n14586 , n14583 , n14584 );
xor ( n14587 , n14494 , n14539 );
and ( n14588 , n824 , n6749 );
and ( n14589 , n14587 , n14588 );
xor ( n14590 , n14587 , n14588 );
xor ( n14591 , n14498 , n14537 );
and ( n14592 , n825 , n6749 );
and ( n14593 , n14591 , n14592 );
xor ( n14594 , n14591 , n14592 );
xor ( n14595 , n14502 , n14535 );
and ( n14596 , n826 , n6749 );
and ( n14597 , n14595 , n14596 );
xor ( n14598 , n14595 , n14596 );
xor ( n14599 , n14506 , n14533 );
and ( n14600 , n827 , n6749 );
and ( n14601 , n14599 , n14600 );
xor ( n14602 , n14599 , n14600 );
xor ( n14603 , n14510 , n14531 );
and ( n14604 , n828 , n6749 );
and ( n14605 , n14603 , n14604 );
xor ( n14606 , n14603 , n14604 );
xor ( n14607 , n14514 , n14529 );
and ( n14608 , n829 , n6749 );
and ( n14609 , n14607 , n14608 );
xor ( n14610 , n14607 , n14608 );
xor ( n14611 , n14518 , n14527 );
and ( n14612 , n830 , n6749 );
and ( n14613 , n14611 , n14612 );
xor ( n14614 , n14611 , n14612 );
xor ( n14615 , n14522 , n14525 );
and ( n14616 , n831 , n6749 );
and ( n14617 , n14615 , n14616 );
and ( n14618 , n14614 , n14617 );
or ( n14619 , n14613 , n14618 );
and ( n14620 , n14610 , n14619 );
or ( n14621 , n14609 , n14620 );
and ( n14622 , n14606 , n14621 );
or ( n14623 , n14605 , n14622 );
and ( n14624 , n14602 , n14623 );
or ( n14625 , n14601 , n14624 );
and ( n14626 , n14598 , n14625 );
or ( n14627 , n14597 , n14626 );
and ( n14628 , n14594 , n14627 );
or ( n14629 , n14593 , n14628 );
and ( n14630 , n14590 , n14629 );
or ( n14631 , n14589 , n14630 );
and ( n14632 , n14586 , n14631 );
or ( n14633 , n14585 , n14632 );
and ( n14634 , n14582 , n14633 );
or ( n14635 , n14581 , n14634 );
and ( n14636 , n14578 , n14635 );
or ( n14637 , n14577 , n14636 );
and ( n14638 , n14574 , n14637 );
or ( n14639 , n14573 , n14638 );
and ( n14640 , n14570 , n14639 );
or ( n14641 , n14569 , n14640 );
and ( n14642 , n14566 , n14641 );
or ( n14643 , n14565 , n14642 );
and ( n14644 , n14562 , n14643 );
or ( n14645 , n14561 , n14644 );
and ( n14646 , n14558 , n14645 );
or ( n14647 , n14557 , n14646 );
and ( n14648 , n816 , n6746 );
and ( n14649 , n14647 , n14648 );
xor ( n14650 , n14647 , n14648 );
xor ( n14651 , n14558 , n14645 );
and ( n14652 , n817 , n6746 );
and ( n14653 , n14651 , n14652 );
xor ( n14654 , n14651 , n14652 );
xor ( n14655 , n14562 , n14643 );
and ( n14656 , n818 , n6746 );
and ( n14657 , n14655 , n14656 );
xor ( n14658 , n14655 , n14656 );
xor ( n14659 , n14566 , n14641 );
and ( n14660 , n819 , n6746 );
and ( n14661 , n14659 , n14660 );
xor ( n14662 , n14659 , n14660 );
xor ( n14663 , n14570 , n14639 );
and ( n14664 , n820 , n6746 );
and ( n14665 , n14663 , n14664 );
xor ( n14666 , n14663 , n14664 );
xor ( n14667 , n14574 , n14637 );
and ( n14668 , n821 , n6746 );
and ( n14669 , n14667 , n14668 );
xor ( n14670 , n14667 , n14668 );
xor ( n14671 , n14578 , n14635 );
and ( n14672 , n822 , n6746 );
and ( n14673 , n14671 , n14672 );
xor ( n14674 , n14671 , n14672 );
xor ( n14675 , n14582 , n14633 );
and ( n14676 , n823 , n6746 );
and ( n14677 , n14675 , n14676 );
xor ( n14678 , n14675 , n14676 );
xor ( n14679 , n14586 , n14631 );
and ( n14680 , n824 , n6746 );
and ( n14681 , n14679 , n14680 );
xor ( n14682 , n14679 , n14680 );
xor ( n14683 , n14590 , n14629 );
and ( n14684 , n825 , n6746 );
and ( n14685 , n14683 , n14684 );
xor ( n14686 , n14683 , n14684 );
xor ( n14687 , n14594 , n14627 );
and ( n14688 , n826 , n6746 );
and ( n14689 , n14687 , n14688 );
xor ( n14690 , n14687 , n14688 );
xor ( n14691 , n14598 , n14625 );
and ( n14692 , n827 , n6746 );
and ( n14693 , n14691 , n14692 );
xor ( n14694 , n14691 , n14692 );
xor ( n14695 , n14602 , n14623 );
and ( n14696 , n828 , n6746 );
and ( n14697 , n14695 , n14696 );
xor ( n14698 , n14695 , n14696 );
xor ( n14699 , n14606 , n14621 );
and ( n14700 , n829 , n6746 );
and ( n14701 , n14699 , n14700 );
xor ( n14702 , n14699 , n14700 );
xor ( n14703 , n14610 , n14619 );
and ( n14704 , n830 , n6746 );
and ( n14705 , n14703 , n14704 );
xor ( n14706 , n14703 , n14704 );
xor ( n14707 , n14614 , n14617 );
and ( n14708 , n831 , n6746 );
and ( n14709 , n14707 , n14708 );
and ( n14710 , n14706 , n14709 );
or ( n14711 , n14705 , n14710 );
and ( n14712 , n14702 , n14711 );
or ( n14713 , n14701 , n14712 );
and ( n14714 , n14698 , n14713 );
or ( n14715 , n14697 , n14714 );
and ( n14716 , n14694 , n14715 );
or ( n14717 , n14693 , n14716 );
and ( n14718 , n14690 , n14717 );
or ( n14719 , n14689 , n14718 );
and ( n14720 , n14686 , n14719 );
or ( n14721 , n14685 , n14720 );
and ( n14722 , n14682 , n14721 );
or ( n14723 , n14681 , n14722 );
and ( n14724 , n14678 , n14723 );
or ( n14725 , n14677 , n14724 );
and ( n14726 , n14674 , n14725 );
or ( n14727 , n14673 , n14726 );
and ( n14728 , n14670 , n14727 );
or ( n14729 , n14669 , n14728 );
and ( n14730 , n14666 , n14729 );
or ( n14731 , n14665 , n14730 );
and ( n14732 , n14662 , n14731 );
or ( n14733 , n14661 , n14732 );
and ( n14734 , n14658 , n14733 );
or ( n14735 , n14657 , n14734 );
and ( n14736 , n14654 , n14735 );
or ( n14737 , n14653 , n14736 );
and ( n14738 , n14650 , n14737 );
or ( n14739 , n14649 , n14738 );
and ( n14740 , n816 , n6743 );
and ( n14741 , n14739 , n14740 );
xor ( n14742 , n14739 , n14740 );
xor ( n14743 , n14650 , n14737 );
and ( n14744 , n817 , n6743 );
and ( n14745 , n14743 , n14744 );
xor ( n14746 , n14743 , n14744 );
xor ( n14747 , n14654 , n14735 );
and ( n14748 , n818 , n6743 );
and ( n14749 , n14747 , n14748 );
xor ( n14750 , n14747 , n14748 );
xor ( n14751 , n14658 , n14733 );
and ( n14752 , n819 , n6743 );
and ( n14753 , n14751 , n14752 );
xor ( n14754 , n14751 , n14752 );
xor ( n14755 , n14662 , n14731 );
and ( n14756 , n820 , n6743 );
and ( n14757 , n14755 , n14756 );
xor ( n14758 , n14755 , n14756 );
xor ( n14759 , n14666 , n14729 );
and ( n14760 , n821 , n6743 );
and ( n14761 , n14759 , n14760 );
xor ( n14762 , n14759 , n14760 );
xor ( n14763 , n14670 , n14727 );
and ( n14764 , n822 , n6743 );
and ( n14765 , n14763 , n14764 );
xor ( n14766 , n14763 , n14764 );
xor ( n14767 , n14674 , n14725 );
and ( n14768 , n823 , n6743 );
and ( n14769 , n14767 , n14768 );
xor ( n14770 , n14767 , n14768 );
xor ( n14771 , n14678 , n14723 );
and ( n14772 , n824 , n6743 );
and ( n14773 , n14771 , n14772 );
xor ( n14774 , n14771 , n14772 );
xor ( n14775 , n14682 , n14721 );
and ( n14776 , n825 , n6743 );
and ( n14777 , n14775 , n14776 );
xor ( n14778 , n14775 , n14776 );
xor ( n14779 , n14686 , n14719 );
and ( n14780 , n826 , n6743 );
and ( n14781 , n14779 , n14780 );
xor ( n14782 , n14779 , n14780 );
xor ( n14783 , n14690 , n14717 );
and ( n14784 , n827 , n6743 );
and ( n14785 , n14783 , n14784 );
xor ( n14786 , n14783 , n14784 );
xor ( n14787 , n14694 , n14715 );
and ( n14788 , n828 , n6743 );
and ( n14789 , n14787 , n14788 );
xor ( n14790 , n14787 , n14788 );
xor ( n14791 , n14698 , n14713 );
and ( n14792 , n829 , n6743 );
and ( n14793 , n14791 , n14792 );
xor ( n14794 , n14791 , n14792 );
xor ( n14795 , n14702 , n14711 );
and ( n14796 , n830 , n6743 );
and ( n14797 , n14795 , n14796 );
xor ( n14798 , n14795 , n14796 );
xor ( n14799 , n14706 , n14709 );
and ( n14800 , n831 , n6743 );
and ( n14801 , n14799 , n14800 );
and ( n14802 , n14798 , n14801 );
or ( n14803 , n14797 , n14802 );
and ( n14804 , n14794 , n14803 );
or ( n14805 , n14793 , n14804 );
and ( n14806 , n14790 , n14805 );
or ( n14807 , n14789 , n14806 );
and ( n14808 , n14786 , n14807 );
or ( n14809 , n14785 , n14808 );
and ( n14810 , n14782 , n14809 );
or ( n14811 , n14781 , n14810 );
and ( n14812 , n14778 , n14811 );
or ( n14813 , n14777 , n14812 );
and ( n14814 , n14774 , n14813 );
or ( n14815 , n14773 , n14814 );
and ( n14816 , n14770 , n14815 );
or ( n14817 , n14769 , n14816 );
and ( n14818 , n14766 , n14817 );
or ( n14819 , n14765 , n14818 );
and ( n14820 , n14762 , n14819 );
or ( n14821 , n14761 , n14820 );
and ( n14822 , n14758 , n14821 );
or ( n14823 , n14757 , n14822 );
and ( n14824 , n14754 , n14823 );
or ( n14825 , n14753 , n14824 );
and ( n14826 , n14750 , n14825 );
or ( n14827 , n14749 , n14826 );
and ( n14828 , n14746 , n14827 );
or ( n14829 , n14745 , n14828 );
and ( n14830 , n14742 , n14829 );
or ( n14831 , n14741 , n14830 );
and ( n14832 , n816 , n6740 );
and ( n14833 , n14831 , n14832 );
xor ( n14834 , n14831 , n14832 );
xor ( n14835 , n14742 , n14829 );
and ( n14836 , n817 , n6740 );
and ( n14837 , n14835 , n14836 );
xor ( n14838 , n14835 , n14836 );
xor ( n14839 , n14746 , n14827 );
and ( n14840 , n818 , n6740 );
and ( n14841 , n14839 , n14840 );
xor ( n14842 , n14839 , n14840 );
xor ( n14843 , n14750 , n14825 );
and ( n14844 , n819 , n6740 );
and ( n14845 , n14843 , n14844 );
xor ( n14846 , n14843 , n14844 );
xor ( n14847 , n14754 , n14823 );
and ( n14848 , n820 , n6740 );
and ( n14849 , n14847 , n14848 );
xor ( n14850 , n14847 , n14848 );
xor ( n14851 , n14758 , n14821 );
and ( n14852 , n821 , n6740 );
and ( n14853 , n14851 , n14852 );
xor ( n14854 , n14851 , n14852 );
xor ( n14855 , n14762 , n14819 );
and ( n14856 , n822 , n6740 );
and ( n14857 , n14855 , n14856 );
xor ( n14858 , n14855 , n14856 );
xor ( n14859 , n14766 , n14817 );
and ( n14860 , n823 , n6740 );
and ( n14861 , n14859 , n14860 );
xor ( n14862 , n14859 , n14860 );
xor ( n14863 , n14770 , n14815 );
and ( n14864 , n824 , n6740 );
and ( n14865 , n14863 , n14864 );
xor ( n14866 , n14863 , n14864 );
xor ( n14867 , n14774 , n14813 );
and ( n14868 , n825 , n6740 );
and ( n14869 , n14867 , n14868 );
xor ( n14870 , n14867 , n14868 );
xor ( n14871 , n14778 , n14811 );
and ( n14872 , n826 , n6740 );
and ( n14873 , n14871 , n14872 );
xor ( n14874 , n14871 , n14872 );
xor ( n14875 , n14782 , n14809 );
and ( n14876 , n827 , n6740 );
and ( n14877 , n14875 , n14876 );
xor ( n14878 , n14875 , n14876 );
xor ( n14879 , n14786 , n14807 );
and ( n14880 , n828 , n6740 );
and ( n14881 , n14879 , n14880 );
xor ( n14882 , n14879 , n14880 );
xor ( n14883 , n14790 , n14805 );
and ( n14884 , n829 , n6740 );
and ( n14885 , n14883 , n14884 );
xor ( n14886 , n14883 , n14884 );
xor ( n14887 , n14794 , n14803 );
and ( n14888 , n830 , n6740 );
and ( n14889 , n14887 , n14888 );
xor ( n14890 , n14887 , n14888 );
xor ( n14891 , n14798 , n14801 );
and ( n14892 , n831 , n6740 );
and ( n14893 , n14891 , n14892 );
and ( n14894 , n14890 , n14893 );
or ( n14895 , n14889 , n14894 );
and ( n14896 , n14886 , n14895 );
or ( n14897 , n14885 , n14896 );
and ( n14898 , n14882 , n14897 );
or ( n14899 , n14881 , n14898 );
and ( n14900 , n14878 , n14899 );
or ( n14901 , n14877 , n14900 );
and ( n14902 , n14874 , n14901 );
or ( n14903 , n14873 , n14902 );
and ( n14904 , n14870 , n14903 );
or ( n14905 , n14869 , n14904 );
and ( n14906 , n14866 , n14905 );
or ( n14907 , n14865 , n14906 );
and ( n14908 , n14862 , n14907 );
or ( n14909 , n14861 , n14908 );
and ( n14910 , n14858 , n14909 );
or ( n14911 , n14857 , n14910 );
and ( n14912 , n14854 , n14911 );
or ( n14913 , n14853 , n14912 );
and ( n14914 , n14850 , n14913 );
or ( n14915 , n14849 , n14914 );
and ( n14916 , n14846 , n14915 );
or ( n14917 , n14845 , n14916 );
and ( n14918 , n14842 , n14917 );
or ( n14919 , n14841 , n14918 );
and ( n14920 , n14838 , n14919 );
or ( n14921 , n14837 , n14920 );
and ( n14922 , n14834 , n14921 );
or ( n14923 , n14833 , n14922 );
and ( n14924 , n816 , n6737 );
and ( n14925 , n14923 , n14924 );
xor ( n14926 , n14923 , n14924 );
xor ( n14927 , n14834 , n14921 );
and ( n14928 , n817 , n6737 );
and ( n14929 , n14927 , n14928 );
xor ( n14930 , n14927 , n14928 );
xor ( n14931 , n14838 , n14919 );
and ( n14932 , n818 , n6737 );
and ( n14933 , n14931 , n14932 );
xor ( n14934 , n14931 , n14932 );
xor ( n14935 , n14842 , n14917 );
and ( n14936 , n819 , n6737 );
and ( n14937 , n14935 , n14936 );
xor ( n14938 , n14935 , n14936 );
xor ( n14939 , n14846 , n14915 );
and ( n14940 , n820 , n6737 );
and ( n14941 , n14939 , n14940 );
xor ( n14942 , n14939 , n14940 );
xor ( n14943 , n14850 , n14913 );
and ( n14944 , n821 , n6737 );
and ( n14945 , n14943 , n14944 );
xor ( n14946 , n14943 , n14944 );
xor ( n14947 , n14854 , n14911 );
and ( n14948 , n822 , n6737 );
and ( n14949 , n14947 , n14948 );
xor ( n14950 , n14947 , n14948 );
xor ( n14951 , n14858 , n14909 );
and ( n14952 , n823 , n6737 );
and ( n14953 , n14951 , n14952 );
xor ( n14954 , n14951 , n14952 );
xor ( n14955 , n14862 , n14907 );
and ( n14956 , n824 , n6737 );
and ( n14957 , n14955 , n14956 );
xor ( n14958 , n14955 , n14956 );
xor ( n14959 , n14866 , n14905 );
and ( n14960 , n825 , n6737 );
and ( n14961 , n14959 , n14960 );
xor ( n14962 , n14959 , n14960 );
xor ( n14963 , n14870 , n14903 );
and ( n14964 , n826 , n6737 );
and ( n14965 , n14963 , n14964 );
xor ( n14966 , n14963 , n14964 );
xor ( n14967 , n14874 , n14901 );
and ( n14968 , n827 , n6737 );
and ( n14969 , n14967 , n14968 );
xor ( n14970 , n14967 , n14968 );
xor ( n14971 , n14878 , n14899 );
and ( n14972 , n828 , n6737 );
and ( n14973 , n14971 , n14972 );
xor ( n14974 , n14971 , n14972 );
xor ( n14975 , n14882 , n14897 );
and ( n14976 , n829 , n6737 );
and ( n14977 , n14975 , n14976 );
xor ( n14978 , n14975 , n14976 );
xor ( n14979 , n14886 , n14895 );
and ( n14980 , n830 , n6737 );
and ( n14981 , n14979 , n14980 );
xor ( n14982 , n14979 , n14980 );
xor ( n14983 , n14890 , n14893 );
and ( n14984 , n831 , n6737 );
and ( n14985 , n14983 , n14984 );
and ( n14986 , n14982 , n14985 );
or ( n14987 , n14981 , n14986 );
and ( n14988 , n14978 , n14987 );
or ( n14989 , n14977 , n14988 );
and ( n14990 , n14974 , n14989 );
or ( n14991 , n14973 , n14990 );
and ( n14992 , n14970 , n14991 );
or ( n14993 , n14969 , n14992 );
and ( n14994 , n14966 , n14993 );
or ( n14995 , n14965 , n14994 );
and ( n14996 , n14962 , n14995 );
or ( n14997 , n14961 , n14996 );
and ( n14998 , n14958 , n14997 );
or ( n14999 , n14957 , n14998 );
and ( n15000 , n14954 , n14999 );
or ( n15001 , n14953 , n15000 );
and ( n15002 , n14950 , n15001 );
or ( n15003 , n14949 , n15002 );
and ( n15004 , n14946 , n15003 );
or ( n15005 , n14945 , n15004 );
and ( n15006 , n14942 , n15005 );
or ( n15007 , n14941 , n15006 );
and ( n15008 , n14938 , n15007 );
or ( n15009 , n14937 , n15008 );
and ( n15010 , n14934 , n15009 );
or ( n15011 , n14933 , n15010 );
and ( n15012 , n14930 , n15011 );
or ( n15013 , n14929 , n15012 );
and ( n15014 , n14926 , n15013 );
or ( n15015 , n14925 , n15014 );
and ( n15016 , n816 , n6734 );
and ( n15017 , n15015 , n15016 );
xor ( n15018 , n15015 , n15016 );
xor ( n15019 , n14926 , n15013 );
and ( n15020 , n817 , n6734 );
and ( n15021 , n15019 , n15020 );
xor ( n15022 , n15019 , n15020 );
xor ( n15023 , n14930 , n15011 );
and ( n15024 , n818 , n6734 );
and ( n15025 , n15023 , n15024 );
xor ( n15026 , n15023 , n15024 );
xor ( n15027 , n14934 , n15009 );
and ( n15028 , n819 , n6734 );
and ( n15029 , n15027 , n15028 );
xor ( n15030 , n15027 , n15028 );
xor ( n15031 , n14938 , n15007 );
and ( n15032 , n820 , n6734 );
and ( n15033 , n15031 , n15032 );
xor ( n15034 , n15031 , n15032 );
xor ( n15035 , n14942 , n15005 );
and ( n15036 , n821 , n6734 );
and ( n15037 , n15035 , n15036 );
xor ( n15038 , n15035 , n15036 );
xor ( n15039 , n14946 , n15003 );
and ( n15040 , n822 , n6734 );
and ( n15041 , n15039 , n15040 );
xor ( n15042 , n15039 , n15040 );
xor ( n15043 , n14950 , n15001 );
and ( n15044 , n823 , n6734 );
and ( n15045 , n15043 , n15044 );
xor ( n15046 , n15043 , n15044 );
xor ( n15047 , n14954 , n14999 );
and ( n15048 , n824 , n6734 );
and ( n15049 , n15047 , n15048 );
xor ( n15050 , n15047 , n15048 );
xor ( n15051 , n14958 , n14997 );
and ( n15052 , n825 , n6734 );
and ( n15053 , n15051 , n15052 );
xor ( n15054 , n15051 , n15052 );
xor ( n15055 , n14962 , n14995 );
and ( n15056 , n826 , n6734 );
and ( n15057 , n15055 , n15056 );
xor ( n15058 , n15055 , n15056 );
xor ( n15059 , n14966 , n14993 );
and ( n15060 , n827 , n6734 );
and ( n15061 , n15059 , n15060 );
xor ( n15062 , n15059 , n15060 );
xor ( n15063 , n14970 , n14991 );
and ( n15064 , n828 , n6734 );
and ( n15065 , n15063 , n15064 );
xor ( n15066 , n15063 , n15064 );
xor ( n15067 , n14974 , n14989 );
and ( n15068 , n829 , n6734 );
and ( n15069 , n15067 , n15068 );
xor ( n15070 , n15067 , n15068 );
xor ( n15071 , n14978 , n14987 );
and ( n15072 , n830 , n6734 );
and ( n15073 , n15071 , n15072 );
xor ( n15074 , n15071 , n15072 );
xor ( n15075 , n14982 , n14985 );
and ( n15076 , n831 , n6734 );
and ( n15077 , n15075 , n15076 );
and ( n15078 , n15074 , n15077 );
or ( n15079 , n15073 , n15078 );
and ( n15080 , n15070 , n15079 );
or ( n15081 , n15069 , n15080 );
and ( n15082 , n15066 , n15081 );
or ( n15083 , n15065 , n15082 );
and ( n15084 , n15062 , n15083 );
or ( n15085 , n15061 , n15084 );
and ( n15086 , n15058 , n15085 );
or ( n15087 , n15057 , n15086 );
and ( n15088 , n15054 , n15087 );
or ( n15089 , n15053 , n15088 );
and ( n15090 , n15050 , n15089 );
or ( n15091 , n15049 , n15090 );
and ( n15092 , n15046 , n15091 );
or ( n15093 , n15045 , n15092 );
and ( n15094 , n15042 , n15093 );
or ( n15095 , n15041 , n15094 );
and ( n15096 , n15038 , n15095 );
or ( n15097 , n15037 , n15096 );
and ( n15098 , n15034 , n15097 );
or ( n15099 , n15033 , n15098 );
and ( n15100 , n15030 , n15099 );
or ( n15101 , n15029 , n15100 );
and ( n15102 , n15026 , n15101 );
or ( n15103 , n15025 , n15102 );
and ( n15104 , n15022 , n15103 );
or ( n15105 , n15021 , n15104 );
and ( n15106 , n15018 , n15105 );
or ( n15107 , n15017 , n15106 );
and ( n15108 , n816 , n6731 );
and ( n15109 , n15107 , n15108 );
xor ( n15110 , n15107 , n15108 );
xor ( n15111 , n15018 , n15105 );
and ( n15112 , n817 , n6731 );
and ( n15113 , n15111 , n15112 );
xor ( n15114 , n15111 , n15112 );
xor ( n15115 , n15022 , n15103 );
and ( n15116 , n818 , n6731 );
and ( n15117 , n15115 , n15116 );
xor ( n15118 , n15115 , n15116 );
xor ( n15119 , n15026 , n15101 );
and ( n15120 , n819 , n6731 );
and ( n15121 , n15119 , n15120 );
xor ( n15122 , n15119 , n15120 );
xor ( n15123 , n15030 , n15099 );
and ( n15124 , n820 , n6731 );
and ( n15125 , n15123 , n15124 );
xor ( n15126 , n15123 , n15124 );
xor ( n15127 , n15034 , n15097 );
and ( n15128 , n821 , n6731 );
and ( n15129 , n15127 , n15128 );
xor ( n15130 , n15127 , n15128 );
xor ( n15131 , n15038 , n15095 );
and ( n15132 , n822 , n6731 );
and ( n15133 , n15131 , n15132 );
xor ( n15134 , n15131 , n15132 );
xor ( n15135 , n15042 , n15093 );
and ( n15136 , n823 , n6731 );
and ( n15137 , n15135 , n15136 );
xor ( n15138 , n15135 , n15136 );
xor ( n15139 , n15046 , n15091 );
and ( n15140 , n824 , n6731 );
and ( n15141 , n15139 , n15140 );
xor ( n15142 , n15139 , n15140 );
xor ( n15143 , n15050 , n15089 );
and ( n15144 , n825 , n6731 );
and ( n15145 , n15143 , n15144 );
xor ( n15146 , n15143 , n15144 );
xor ( n15147 , n15054 , n15087 );
and ( n15148 , n826 , n6731 );
and ( n15149 , n15147 , n15148 );
xor ( n15150 , n15147 , n15148 );
xor ( n15151 , n15058 , n15085 );
and ( n15152 , n827 , n6731 );
and ( n15153 , n15151 , n15152 );
xor ( n15154 , n15151 , n15152 );
xor ( n15155 , n15062 , n15083 );
and ( n15156 , n828 , n6731 );
and ( n15157 , n15155 , n15156 );
xor ( n15158 , n15155 , n15156 );
xor ( n15159 , n15066 , n15081 );
and ( n15160 , n829 , n6731 );
and ( n15161 , n15159 , n15160 );
xor ( n15162 , n15159 , n15160 );
xor ( n15163 , n15070 , n15079 );
and ( n15164 , n830 , n6731 );
and ( n15165 , n15163 , n15164 );
xor ( n15166 , n15163 , n15164 );
xor ( n15167 , n15074 , n15077 );
and ( n15168 , n831 , n6731 );
and ( n15169 , n15167 , n15168 );
and ( n15170 , n15166 , n15169 );
or ( n15171 , n15165 , n15170 );
and ( n15172 , n15162 , n15171 );
or ( n15173 , n15161 , n15172 );
and ( n15174 , n15158 , n15173 );
or ( n15175 , n15157 , n15174 );
and ( n15176 , n15154 , n15175 );
or ( n15177 , n15153 , n15176 );
and ( n15178 , n15150 , n15177 );
or ( n15179 , n15149 , n15178 );
and ( n15180 , n15146 , n15179 );
or ( n15181 , n15145 , n15180 );
and ( n15182 , n15142 , n15181 );
or ( n15183 , n15141 , n15182 );
and ( n15184 , n15138 , n15183 );
or ( n15185 , n15137 , n15184 );
and ( n15186 , n15134 , n15185 );
or ( n15187 , n15133 , n15186 );
and ( n15188 , n15130 , n15187 );
or ( n15189 , n15129 , n15188 );
and ( n15190 , n15126 , n15189 );
or ( n15191 , n15125 , n15190 );
and ( n15192 , n15122 , n15191 );
or ( n15193 , n15121 , n15192 );
and ( n15194 , n15118 , n15193 );
or ( n15195 , n15117 , n15194 );
and ( n15196 , n15114 , n15195 );
or ( n15197 , n15113 , n15196 );
and ( n15198 , n15110 , n15197 );
or ( n15199 , n15109 , n15198 );
and ( n15200 , n816 , n6728 );
and ( n15201 , n15199 , n15200 );
xor ( n15202 , n15199 , n15200 );
xor ( n15203 , n15110 , n15197 );
and ( n15204 , n817 , n6728 );
and ( n15205 , n15203 , n15204 );
xor ( n15206 , n15203 , n15204 );
xor ( n15207 , n15114 , n15195 );
and ( n15208 , n818 , n6728 );
and ( n15209 , n15207 , n15208 );
xor ( n15210 , n15207 , n15208 );
xor ( n15211 , n15118 , n15193 );
and ( n15212 , n819 , n6728 );
and ( n15213 , n15211 , n15212 );
xor ( n15214 , n15211 , n15212 );
xor ( n15215 , n15122 , n15191 );
and ( n15216 , n820 , n6728 );
and ( n15217 , n15215 , n15216 );
xor ( n15218 , n15215 , n15216 );
xor ( n15219 , n15126 , n15189 );
and ( n15220 , n821 , n6728 );
and ( n15221 , n15219 , n15220 );
xor ( n15222 , n15219 , n15220 );
xor ( n15223 , n15130 , n15187 );
and ( n15224 , n822 , n6728 );
and ( n15225 , n15223 , n15224 );
xor ( n15226 , n15223 , n15224 );
xor ( n15227 , n15134 , n15185 );
and ( n15228 , n823 , n6728 );
and ( n15229 , n15227 , n15228 );
xor ( n15230 , n15227 , n15228 );
xor ( n15231 , n15138 , n15183 );
and ( n15232 , n824 , n6728 );
and ( n15233 , n15231 , n15232 );
xor ( n15234 , n15231 , n15232 );
xor ( n15235 , n15142 , n15181 );
and ( n15236 , n825 , n6728 );
and ( n15237 , n15235 , n15236 );
xor ( n15238 , n15235 , n15236 );
xor ( n15239 , n15146 , n15179 );
and ( n15240 , n826 , n6728 );
and ( n15241 , n15239 , n15240 );
xor ( n15242 , n15239 , n15240 );
xor ( n15243 , n15150 , n15177 );
and ( n15244 , n827 , n6728 );
and ( n15245 , n15243 , n15244 );
xor ( n15246 , n15243 , n15244 );
xor ( n15247 , n15154 , n15175 );
and ( n15248 , n828 , n6728 );
and ( n15249 , n15247 , n15248 );
xor ( n15250 , n15247 , n15248 );
xor ( n15251 , n15158 , n15173 );
and ( n15252 , n829 , n6728 );
and ( n15253 , n15251 , n15252 );
xor ( n15254 , n15251 , n15252 );
xor ( n15255 , n15162 , n15171 );
and ( n15256 , n830 , n6728 );
and ( n15257 , n15255 , n15256 );
xor ( n15258 , n15255 , n15256 );
xor ( n15259 , n15166 , n15169 );
and ( n15260 , n831 , n6728 );
and ( n15261 , n15259 , n15260 );
and ( n15262 , n15258 , n15261 );
or ( n15263 , n15257 , n15262 );
and ( n15264 , n15254 , n15263 );
or ( n15265 , n15253 , n15264 );
and ( n15266 , n15250 , n15265 );
or ( n15267 , n15249 , n15266 );
and ( n15268 , n15246 , n15267 );
or ( n15269 , n15245 , n15268 );
and ( n15270 , n15242 , n15269 );
or ( n15271 , n15241 , n15270 );
and ( n15272 , n15238 , n15271 );
or ( n15273 , n15237 , n15272 );
and ( n15274 , n15234 , n15273 );
or ( n15275 , n15233 , n15274 );
and ( n15276 , n15230 , n15275 );
or ( n15277 , n15229 , n15276 );
and ( n15278 , n15226 , n15277 );
or ( n15279 , n15225 , n15278 );
and ( n15280 , n15222 , n15279 );
or ( n15281 , n15221 , n15280 );
and ( n15282 , n15218 , n15281 );
or ( n15283 , n15217 , n15282 );
and ( n15284 , n15214 , n15283 );
or ( n15285 , n15213 , n15284 );
and ( n15286 , n15210 , n15285 );
or ( n15287 , n15209 , n15286 );
and ( n15288 , n15206 , n15287 );
or ( n15289 , n15205 , n15288 );
and ( n15290 , n15202 , n15289 );
or ( n15291 , n15201 , n15290 );
and ( n15292 , n816 , n6725 );
and ( n15293 , n15291 , n15292 );
xor ( n15294 , n15291 , n15292 );
xor ( n15295 , n15202 , n15289 );
and ( n15296 , n817 , n6725 );
and ( n15297 , n15295 , n15296 );
xor ( n15298 , n15295 , n15296 );
xor ( n15299 , n15206 , n15287 );
and ( n15300 , n818 , n6725 );
and ( n15301 , n15299 , n15300 );
xor ( n15302 , n15299 , n15300 );
xor ( n15303 , n15210 , n15285 );
and ( n15304 , n819 , n6725 );
and ( n15305 , n15303 , n15304 );
xor ( n15306 , n15303 , n15304 );
xor ( n15307 , n15214 , n15283 );
and ( n15308 , n820 , n6725 );
and ( n15309 , n15307 , n15308 );
xor ( n15310 , n15307 , n15308 );
xor ( n15311 , n15218 , n15281 );
and ( n15312 , n821 , n6725 );
and ( n15313 , n15311 , n15312 );
xor ( n15314 , n15311 , n15312 );
xor ( n15315 , n15222 , n15279 );
and ( n15316 , n822 , n6725 );
and ( n15317 , n15315 , n15316 );
xor ( n15318 , n15315 , n15316 );
xor ( n15319 , n15226 , n15277 );
and ( n15320 , n823 , n6725 );
and ( n15321 , n15319 , n15320 );
xor ( n15322 , n15319 , n15320 );
xor ( n15323 , n15230 , n15275 );
and ( n15324 , n824 , n6725 );
and ( n15325 , n15323 , n15324 );
xor ( n15326 , n15323 , n15324 );
xor ( n15327 , n15234 , n15273 );
and ( n15328 , n825 , n6725 );
and ( n15329 , n15327 , n15328 );
xor ( n15330 , n15327 , n15328 );
xor ( n15331 , n15238 , n15271 );
and ( n15332 , n826 , n6725 );
and ( n15333 , n15331 , n15332 );
xor ( n15334 , n15331 , n15332 );
xor ( n15335 , n15242 , n15269 );
and ( n15336 , n827 , n6725 );
and ( n15337 , n15335 , n15336 );
xor ( n15338 , n15335 , n15336 );
xor ( n15339 , n15246 , n15267 );
and ( n15340 , n828 , n6725 );
and ( n15341 , n15339 , n15340 );
xor ( n15342 , n15339 , n15340 );
xor ( n15343 , n15250 , n15265 );
and ( n15344 , n829 , n6725 );
and ( n15345 , n15343 , n15344 );
xor ( n15346 , n15343 , n15344 );
xor ( n15347 , n15254 , n15263 );
and ( n15348 , n830 , n6725 );
and ( n15349 , n15347 , n15348 );
xor ( n15350 , n15347 , n15348 );
xor ( n15351 , n15258 , n15261 );
and ( n15352 , n831 , n6725 );
and ( n15353 , n15351 , n15352 );
and ( n15354 , n15350 , n15353 );
or ( n15355 , n15349 , n15354 );
and ( n15356 , n15346 , n15355 );
or ( n15357 , n15345 , n15356 );
and ( n15358 , n15342 , n15357 );
or ( n15359 , n15341 , n15358 );
and ( n15360 , n15338 , n15359 );
or ( n15361 , n15337 , n15360 );
and ( n15362 , n15334 , n15361 );
or ( n15363 , n15333 , n15362 );
and ( n15364 , n15330 , n15363 );
or ( n15365 , n15329 , n15364 );
and ( n15366 , n15326 , n15365 );
or ( n15367 , n15325 , n15366 );
and ( n15368 , n15322 , n15367 );
or ( n15369 , n15321 , n15368 );
and ( n15370 , n15318 , n15369 );
or ( n15371 , n15317 , n15370 );
and ( n15372 , n15314 , n15371 );
or ( n15373 , n15313 , n15372 );
and ( n15374 , n15310 , n15373 );
or ( n15375 , n15309 , n15374 );
and ( n15376 , n15306 , n15375 );
or ( n15377 , n15305 , n15376 );
and ( n15378 , n15302 , n15377 );
or ( n15379 , n15301 , n15378 );
and ( n15380 , n15298 , n15379 );
or ( n15381 , n15297 , n15380 );
and ( n15382 , n15294 , n15381 );
or ( n15383 , n15293 , n15382 );
and ( n15384 , n816 , n6722 );
and ( n15385 , n15383 , n15384 );
xor ( n15386 , n15383 , n15384 );
xor ( n15387 , n15294 , n15381 );
and ( n15388 , n817 , n6722 );
and ( n15389 , n15387 , n15388 );
xor ( n15390 , n15387 , n15388 );
xor ( n15391 , n15298 , n15379 );
and ( n15392 , n818 , n6722 );
and ( n15393 , n15391 , n15392 );
xor ( n15394 , n15391 , n15392 );
xor ( n15395 , n15302 , n15377 );
and ( n15396 , n819 , n6722 );
and ( n15397 , n15395 , n15396 );
xor ( n15398 , n15395 , n15396 );
xor ( n15399 , n15306 , n15375 );
and ( n15400 , n820 , n6722 );
and ( n15401 , n15399 , n15400 );
xor ( n15402 , n15399 , n15400 );
xor ( n15403 , n15310 , n15373 );
and ( n15404 , n821 , n6722 );
and ( n15405 , n15403 , n15404 );
xor ( n15406 , n15403 , n15404 );
xor ( n15407 , n15314 , n15371 );
and ( n15408 , n822 , n6722 );
and ( n15409 , n15407 , n15408 );
xor ( n15410 , n15407 , n15408 );
xor ( n15411 , n15318 , n15369 );
and ( n15412 , n823 , n6722 );
and ( n15413 , n15411 , n15412 );
xor ( n15414 , n15411 , n15412 );
xor ( n15415 , n15322 , n15367 );
and ( n15416 , n824 , n6722 );
and ( n15417 , n15415 , n15416 );
xor ( n15418 , n15415 , n15416 );
xor ( n15419 , n15326 , n15365 );
and ( n15420 , n825 , n6722 );
and ( n15421 , n15419 , n15420 );
xor ( n15422 , n15419 , n15420 );
xor ( n15423 , n15330 , n15363 );
and ( n15424 , n826 , n6722 );
and ( n15425 , n15423 , n15424 );
xor ( n15426 , n15423 , n15424 );
xor ( n15427 , n15334 , n15361 );
and ( n15428 , n827 , n6722 );
and ( n15429 , n15427 , n15428 );
xor ( n15430 , n15427 , n15428 );
xor ( n15431 , n15338 , n15359 );
and ( n15432 , n828 , n6722 );
and ( n15433 , n15431 , n15432 );
xor ( n15434 , n15431 , n15432 );
xor ( n15435 , n15342 , n15357 );
and ( n15436 , n829 , n6722 );
and ( n15437 , n15435 , n15436 );
xor ( n15438 , n15435 , n15436 );
xor ( n15439 , n15346 , n15355 );
and ( n15440 , n830 , n6722 );
and ( n15441 , n15439 , n15440 );
xor ( n15442 , n15439 , n15440 );
xor ( n15443 , n15350 , n15353 );
and ( n15444 , n831 , n6722 );
and ( n15445 , n15443 , n15444 );
and ( n15446 , n15442 , n15445 );
or ( n15447 , n15441 , n15446 );
and ( n15448 , n15438 , n15447 );
or ( n15449 , n15437 , n15448 );
and ( n15450 , n15434 , n15449 );
or ( n15451 , n15433 , n15450 );
and ( n15452 , n15430 , n15451 );
or ( n15453 , n15429 , n15452 );
and ( n15454 , n15426 , n15453 );
or ( n15455 , n15425 , n15454 );
and ( n15456 , n15422 , n15455 );
or ( n15457 , n15421 , n15456 );
and ( n15458 , n15418 , n15457 );
or ( n15459 , n15417 , n15458 );
and ( n15460 , n15414 , n15459 );
or ( n15461 , n15413 , n15460 );
and ( n15462 , n15410 , n15461 );
or ( n15463 , n15409 , n15462 );
and ( n15464 , n15406 , n15463 );
or ( n15465 , n15405 , n15464 );
and ( n15466 , n15402 , n15465 );
or ( n15467 , n15401 , n15466 );
and ( n15468 , n15398 , n15467 );
or ( n15469 , n15397 , n15468 );
and ( n15470 , n15394 , n15469 );
or ( n15471 , n15393 , n15470 );
and ( n15472 , n15390 , n15471 );
or ( n15473 , n15389 , n15472 );
and ( n15474 , n15386 , n15473 );
or ( n15475 , n15385 , n15474 );
and ( n15476 , n816 , n6719 );
and ( n15477 , n15475 , n15476 );
xor ( n15478 , n15475 , n15476 );
xor ( n15479 , n15386 , n15473 );
and ( n15480 , n817 , n6719 );
and ( n15481 , n15479 , n15480 );
xor ( n15482 , n15479 , n15480 );
xor ( n15483 , n15390 , n15471 );
and ( n15484 , n818 , n6719 );
and ( n15485 , n15483 , n15484 );
xor ( n15486 , n15483 , n15484 );
xor ( n15487 , n15394 , n15469 );
and ( n15488 , n819 , n6719 );
and ( n15489 , n15487 , n15488 );
xor ( n15490 , n15487 , n15488 );
xor ( n15491 , n15398 , n15467 );
and ( n15492 , n820 , n6719 );
and ( n15493 , n15491 , n15492 );
xor ( n15494 , n15491 , n15492 );
xor ( n15495 , n15402 , n15465 );
and ( n15496 , n821 , n6719 );
and ( n15497 , n15495 , n15496 );
xor ( n15498 , n15495 , n15496 );
xor ( n15499 , n15406 , n15463 );
and ( n15500 , n822 , n6719 );
and ( n15501 , n15499 , n15500 );
xor ( n15502 , n15499 , n15500 );
xor ( n15503 , n15410 , n15461 );
and ( n15504 , n823 , n6719 );
and ( n15505 , n15503 , n15504 );
xor ( n15506 , n15503 , n15504 );
xor ( n15507 , n15414 , n15459 );
and ( n15508 , n824 , n6719 );
and ( n15509 , n15507 , n15508 );
xor ( n15510 , n15507 , n15508 );
xor ( n15511 , n15418 , n15457 );
and ( n15512 , n825 , n6719 );
and ( n15513 , n15511 , n15512 );
xor ( n15514 , n15511 , n15512 );
xor ( n15515 , n15422 , n15455 );
and ( n15516 , n826 , n6719 );
and ( n15517 , n15515 , n15516 );
xor ( n15518 , n15515 , n15516 );
xor ( n15519 , n15426 , n15453 );
and ( n15520 , n827 , n6719 );
and ( n15521 , n15519 , n15520 );
xor ( n15522 , n15519 , n15520 );
xor ( n15523 , n15430 , n15451 );
and ( n15524 , n828 , n6719 );
and ( n15525 , n15523 , n15524 );
xor ( n15526 , n15523 , n15524 );
xor ( n15527 , n15434 , n15449 );
and ( n15528 , n829 , n6719 );
and ( n15529 , n15527 , n15528 );
xor ( n15530 , n15527 , n15528 );
xor ( n15531 , n15438 , n15447 );
and ( n15532 , n830 , n6719 );
and ( n15533 , n15531 , n15532 );
xor ( n15534 , n15531 , n15532 );
xor ( n15535 , n15442 , n15445 );
and ( n15536 , n831 , n6719 );
and ( n15537 , n15535 , n15536 );
and ( n15538 , n15534 , n15537 );
or ( n15539 , n15533 , n15538 );
and ( n15540 , n15530 , n15539 );
or ( n15541 , n15529 , n15540 );
and ( n15542 , n15526 , n15541 );
or ( n15543 , n15525 , n15542 );
and ( n15544 , n15522 , n15543 );
or ( n15545 , n15521 , n15544 );
and ( n15546 , n15518 , n15545 );
or ( n15547 , n15517 , n15546 );
and ( n15548 , n15514 , n15547 );
or ( n15549 , n15513 , n15548 );
and ( n15550 , n15510 , n15549 );
or ( n15551 , n15509 , n15550 );
and ( n15552 , n15506 , n15551 );
or ( n15553 , n15505 , n15552 );
and ( n15554 , n15502 , n15553 );
or ( n15555 , n15501 , n15554 );
and ( n15556 , n15498 , n15555 );
or ( n15557 , n15497 , n15556 );
and ( n15558 , n15494 , n15557 );
or ( n15559 , n15493 , n15558 );
and ( n15560 , n15490 , n15559 );
or ( n15561 , n15489 , n15560 );
and ( n15562 , n15486 , n15561 );
or ( n15563 , n15485 , n15562 );
and ( n15564 , n15482 , n15563 );
or ( n15565 , n15481 , n15564 );
and ( n15566 , n15478 , n15565 );
or ( n15567 , n15477 , n15566 );
and ( n15568 , n816 , n6716 );
and ( n15569 , n15567 , n15568 );
xor ( n15570 , n15567 , n15568 );
xor ( n15571 , n15478 , n15565 );
and ( n15572 , n817 , n6716 );
and ( n15573 , n15571 , n15572 );
xor ( n15574 , n15571 , n15572 );
xor ( n15575 , n15482 , n15563 );
and ( n15576 , n818 , n6716 );
and ( n15577 , n15575 , n15576 );
xor ( n15578 , n15575 , n15576 );
xor ( n15579 , n15486 , n15561 );
and ( n15580 , n819 , n6716 );
and ( n15581 , n15579 , n15580 );
xor ( n15582 , n15579 , n15580 );
xor ( n15583 , n15490 , n15559 );
and ( n15584 , n820 , n6716 );
and ( n15585 , n15583 , n15584 );
xor ( n15586 , n15583 , n15584 );
xor ( n15587 , n15494 , n15557 );
and ( n15588 , n821 , n6716 );
and ( n15589 , n15587 , n15588 );
xor ( n15590 , n15587 , n15588 );
xor ( n15591 , n15498 , n15555 );
and ( n15592 , n822 , n6716 );
and ( n15593 , n15591 , n15592 );
xor ( n15594 , n15591 , n15592 );
xor ( n15595 , n15502 , n15553 );
and ( n15596 , n823 , n6716 );
and ( n15597 , n15595 , n15596 );
xor ( n15598 , n15595 , n15596 );
xor ( n15599 , n15506 , n15551 );
and ( n15600 , n824 , n6716 );
and ( n15601 , n15599 , n15600 );
xor ( n15602 , n15599 , n15600 );
xor ( n15603 , n15510 , n15549 );
and ( n15604 , n825 , n6716 );
and ( n15605 , n15603 , n15604 );
xor ( n15606 , n15603 , n15604 );
xor ( n15607 , n15514 , n15547 );
and ( n15608 , n826 , n6716 );
and ( n15609 , n15607 , n15608 );
xor ( n15610 , n15607 , n15608 );
xor ( n15611 , n15518 , n15545 );
and ( n15612 , n827 , n6716 );
and ( n15613 , n15611 , n15612 );
xor ( n15614 , n15611 , n15612 );
xor ( n15615 , n15522 , n15543 );
and ( n15616 , n828 , n6716 );
and ( n15617 , n15615 , n15616 );
xor ( n15618 , n15615 , n15616 );
xor ( n15619 , n15526 , n15541 );
and ( n15620 , n829 , n6716 );
and ( n15621 , n15619 , n15620 );
xor ( n15622 , n15619 , n15620 );
xor ( n15623 , n15530 , n15539 );
and ( n15624 , n830 , n6716 );
and ( n15625 , n15623 , n15624 );
xor ( n15626 , n15623 , n15624 );
xor ( n15627 , n15534 , n15537 );
and ( n15628 , n831 , n6716 );
and ( n15629 , n15627 , n15628 );
and ( n15630 , n15626 , n15629 );
or ( n15631 , n15625 , n15630 );
and ( n15632 , n15622 , n15631 );
or ( n15633 , n15621 , n15632 );
and ( n15634 , n15618 , n15633 );
or ( n15635 , n15617 , n15634 );
and ( n15636 , n15614 , n15635 );
or ( n15637 , n15613 , n15636 );
and ( n15638 , n15610 , n15637 );
or ( n15639 , n15609 , n15638 );
and ( n15640 , n15606 , n15639 );
or ( n15641 , n15605 , n15640 );
and ( n15642 , n15602 , n15641 );
or ( n15643 , n15601 , n15642 );
and ( n15644 , n15598 , n15643 );
or ( n15645 , n15597 , n15644 );
and ( n15646 , n15594 , n15645 );
or ( n15647 , n15593 , n15646 );
and ( n15648 , n15590 , n15647 );
or ( n15649 , n15589 , n15648 );
and ( n15650 , n15586 , n15649 );
or ( n15651 , n15585 , n15650 );
and ( n15652 , n15582 , n15651 );
or ( n15653 , n15581 , n15652 );
and ( n15654 , n15578 , n15653 );
or ( n15655 , n15577 , n15654 );
and ( n15656 , n15574 , n15655 );
or ( n15657 , n15573 , n15656 );
and ( n15658 , n15570 , n15657 );
or ( n15659 , n15569 , n15658 );
and ( n15660 , n816 , n6713 );
and ( n15661 , n15659 , n15660 );
xor ( n15662 , n15659 , n15660 );
xor ( n15663 , n15570 , n15657 );
and ( n15664 , n817 , n6713 );
and ( n15665 , n15663 , n15664 );
xor ( n15666 , n15663 , n15664 );
xor ( n15667 , n15574 , n15655 );
and ( n15668 , n818 , n6713 );
and ( n15669 , n15667 , n15668 );
xor ( n15670 , n15667 , n15668 );
xor ( n15671 , n15578 , n15653 );
and ( n15672 , n819 , n6713 );
and ( n15673 , n15671 , n15672 );
xor ( n15674 , n15671 , n15672 );
xor ( n15675 , n15582 , n15651 );
and ( n15676 , n820 , n6713 );
and ( n15677 , n15675 , n15676 );
xor ( n15678 , n15675 , n15676 );
xor ( n15679 , n15586 , n15649 );
and ( n15680 , n821 , n6713 );
and ( n15681 , n15679 , n15680 );
xor ( n15682 , n15679 , n15680 );
xor ( n15683 , n15590 , n15647 );
and ( n15684 , n822 , n6713 );
and ( n15685 , n15683 , n15684 );
xor ( n15686 , n15683 , n15684 );
xor ( n15687 , n15594 , n15645 );
and ( n15688 , n823 , n6713 );
and ( n15689 , n15687 , n15688 );
xor ( n15690 , n15687 , n15688 );
xor ( n15691 , n15598 , n15643 );
and ( n15692 , n824 , n6713 );
and ( n15693 , n15691 , n15692 );
xor ( n15694 , n15691 , n15692 );
xor ( n15695 , n15602 , n15641 );
and ( n15696 , n825 , n6713 );
and ( n15697 , n15695 , n15696 );
xor ( n15698 , n15695 , n15696 );
xor ( n15699 , n15606 , n15639 );
and ( n15700 , n826 , n6713 );
and ( n15701 , n15699 , n15700 );
xor ( n15702 , n15699 , n15700 );
xor ( n15703 , n15610 , n15637 );
and ( n15704 , n827 , n6713 );
and ( n15705 , n15703 , n15704 );
xor ( n15706 , n15703 , n15704 );
xor ( n15707 , n15614 , n15635 );
and ( n15708 , n828 , n6713 );
and ( n15709 , n15707 , n15708 );
xor ( n15710 , n15707 , n15708 );
xor ( n15711 , n15618 , n15633 );
and ( n15712 , n829 , n6713 );
and ( n15713 , n15711 , n15712 );
xor ( n15714 , n15711 , n15712 );
xor ( n15715 , n15622 , n15631 );
and ( n15716 , n830 , n6713 );
and ( n15717 , n15715 , n15716 );
xor ( n15718 , n15715 , n15716 );
xor ( n15719 , n15626 , n15629 );
and ( n15720 , n831 , n6713 );
and ( n15721 , n15719 , n15720 );
and ( n15722 , n15718 , n15721 );
or ( n15723 , n15717 , n15722 );
and ( n15724 , n15714 , n15723 );
or ( n15725 , n15713 , n15724 );
and ( n15726 , n15710 , n15725 );
or ( n15727 , n15709 , n15726 );
and ( n15728 , n15706 , n15727 );
or ( n15729 , n15705 , n15728 );
and ( n15730 , n15702 , n15729 );
or ( n15731 , n15701 , n15730 );
and ( n15732 , n15698 , n15731 );
or ( n15733 , n15697 , n15732 );
and ( n15734 , n15694 , n15733 );
or ( n15735 , n15693 , n15734 );
and ( n15736 , n15690 , n15735 );
or ( n15737 , n15689 , n15736 );
and ( n15738 , n15686 , n15737 );
or ( n15739 , n15685 , n15738 );
and ( n15740 , n15682 , n15739 );
or ( n15741 , n15681 , n15740 );
and ( n15742 , n15678 , n15741 );
or ( n15743 , n15677 , n15742 );
and ( n15744 , n15674 , n15743 );
or ( n15745 , n15673 , n15744 );
and ( n15746 , n15670 , n15745 );
or ( n15747 , n15669 , n15746 );
and ( n15748 , n15666 , n15747 );
or ( n15749 , n15665 , n15748 );
and ( n15750 , n15662 , n15749 );
or ( n15751 , n15661 , n15750 );
and ( n15752 , n816 , n6710 );
and ( n15753 , n15751 , n15752 );
xor ( n15754 , n15751 , n15752 );
xor ( n15755 , n15662 , n15749 );
and ( n15756 , n817 , n6710 );
and ( n15757 , n15755 , n15756 );
xor ( n15758 , n15755 , n15756 );
xor ( n15759 , n15666 , n15747 );
and ( n15760 , n818 , n6710 );
and ( n15761 , n15759 , n15760 );
xor ( n15762 , n15759 , n15760 );
xor ( n15763 , n15670 , n15745 );
and ( n15764 , n819 , n6710 );
and ( n15765 , n15763 , n15764 );
xor ( n15766 , n15763 , n15764 );
xor ( n15767 , n15674 , n15743 );
and ( n15768 , n820 , n6710 );
and ( n15769 , n15767 , n15768 );
xor ( n15770 , n15767 , n15768 );
xor ( n15771 , n15678 , n15741 );
and ( n15772 , n821 , n6710 );
and ( n15773 , n15771 , n15772 );
xor ( n15774 , n15771 , n15772 );
xor ( n15775 , n15682 , n15739 );
and ( n15776 , n822 , n6710 );
and ( n15777 , n15775 , n15776 );
xor ( n15778 , n15775 , n15776 );
xor ( n15779 , n15686 , n15737 );
and ( n15780 , n823 , n6710 );
and ( n15781 , n15779 , n15780 );
xor ( n15782 , n15779 , n15780 );
xor ( n15783 , n15690 , n15735 );
and ( n15784 , n824 , n6710 );
and ( n15785 , n15783 , n15784 );
xor ( n15786 , n15783 , n15784 );
xor ( n15787 , n15694 , n15733 );
and ( n15788 , n825 , n6710 );
and ( n15789 , n15787 , n15788 );
xor ( n15790 , n15787 , n15788 );
xor ( n15791 , n15698 , n15731 );
and ( n15792 , n826 , n6710 );
and ( n15793 , n15791 , n15792 );
xor ( n15794 , n15791 , n15792 );
xor ( n15795 , n15702 , n15729 );
and ( n15796 , n827 , n6710 );
and ( n15797 , n15795 , n15796 );
xor ( n15798 , n15795 , n15796 );
xor ( n15799 , n15706 , n15727 );
and ( n15800 , n828 , n6710 );
and ( n15801 , n15799 , n15800 );
xor ( n15802 , n15799 , n15800 );
xor ( n15803 , n15710 , n15725 );
and ( n15804 , n829 , n6710 );
and ( n15805 , n15803 , n15804 );
xor ( n15806 , n15803 , n15804 );
xor ( n15807 , n15714 , n15723 );
and ( n15808 , n830 , n6710 );
and ( n15809 , n15807 , n15808 );
xor ( n15810 , n15807 , n15808 );
xor ( n15811 , n15718 , n15721 );
and ( n15812 , n831 , n6710 );
and ( n15813 , n15811 , n15812 );
and ( n15814 , n15810 , n15813 );
or ( n15815 , n15809 , n15814 );
and ( n15816 , n15806 , n15815 );
or ( n15817 , n15805 , n15816 );
and ( n15818 , n15802 , n15817 );
or ( n15819 , n15801 , n15818 );
and ( n15820 , n15798 , n15819 );
or ( n15821 , n15797 , n15820 );
and ( n15822 , n15794 , n15821 );
or ( n15823 , n15793 , n15822 );
and ( n15824 , n15790 , n15823 );
or ( n15825 , n15789 , n15824 );
and ( n15826 , n15786 , n15825 );
or ( n15827 , n15785 , n15826 );
and ( n15828 , n15782 , n15827 );
or ( n15829 , n15781 , n15828 );
and ( n15830 , n15778 , n15829 );
or ( n15831 , n15777 , n15830 );
and ( n15832 , n15774 , n15831 );
or ( n15833 , n15773 , n15832 );
and ( n15834 , n15770 , n15833 );
or ( n15835 , n15769 , n15834 );
and ( n15836 , n15766 , n15835 );
or ( n15837 , n15765 , n15836 );
and ( n15838 , n15762 , n15837 );
or ( n15839 , n15761 , n15838 );
and ( n15840 , n15758 , n15839 );
or ( n15841 , n15757 , n15840 );
and ( n15842 , n15754 , n15841 );
or ( n15843 , n15753 , n15842 );
and ( n15844 , n816 , n6707 );
and ( n15845 , n15843 , n15844 );
xor ( n15846 , n15843 , n15844 );
xor ( n15847 , n15754 , n15841 );
and ( n15848 , n817 , n6707 );
and ( n15849 , n15847 , n15848 );
xor ( n15850 , n15847 , n15848 );
xor ( n15851 , n15758 , n15839 );
and ( n15852 , n818 , n6707 );
and ( n15853 , n15851 , n15852 );
xor ( n15854 , n15851 , n15852 );
xor ( n15855 , n15762 , n15837 );
and ( n15856 , n819 , n6707 );
and ( n15857 , n15855 , n15856 );
xor ( n15858 , n15855 , n15856 );
xor ( n15859 , n15766 , n15835 );
and ( n15860 , n820 , n6707 );
and ( n15861 , n15859 , n15860 );
xor ( n15862 , n15859 , n15860 );
xor ( n15863 , n15770 , n15833 );
and ( n15864 , n821 , n6707 );
and ( n15865 , n15863 , n15864 );
xor ( n15866 , n15863 , n15864 );
xor ( n15867 , n15774 , n15831 );
and ( n15868 , n822 , n6707 );
and ( n15869 , n15867 , n15868 );
xor ( n15870 , n15867 , n15868 );
xor ( n15871 , n15778 , n15829 );
and ( n15872 , n823 , n6707 );
and ( n15873 , n15871 , n15872 );
xor ( n15874 , n15871 , n15872 );
xor ( n15875 , n15782 , n15827 );
and ( n15876 , n824 , n6707 );
and ( n15877 , n15875 , n15876 );
xor ( n15878 , n15875 , n15876 );
xor ( n15879 , n15786 , n15825 );
and ( n15880 , n825 , n6707 );
and ( n15881 , n15879 , n15880 );
xor ( n15882 , n15879 , n15880 );
xor ( n15883 , n15790 , n15823 );
and ( n15884 , n826 , n6707 );
and ( n15885 , n15883 , n15884 );
xor ( n15886 , n15883 , n15884 );
xor ( n15887 , n15794 , n15821 );
and ( n15888 , n827 , n6707 );
and ( n15889 , n15887 , n15888 );
xor ( n15890 , n15887 , n15888 );
xor ( n15891 , n15798 , n15819 );
and ( n15892 , n828 , n6707 );
and ( n15893 , n15891 , n15892 );
xor ( n15894 , n15891 , n15892 );
xor ( n15895 , n15802 , n15817 );
and ( n15896 , n829 , n6707 );
and ( n15897 , n15895 , n15896 );
xor ( n15898 , n15895 , n15896 );
xor ( n15899 , n15806 , n15815 );
and ( n15900 , n830 , n6707 );
and ( n15901 , n15899 , n15900 );
xor ( n15902 , n15899 , n15900 );
xor ( n15903 , n15810 , n15813 );
and ( n15904 , n831 , n6707 );
and ( n15905 , n15903 , n15904 );
and ( n15906 , n15902 , n15905 );
or ( n15907 , n15901 , n15906 );
and ( n15908 , n15898 , n15907 );
or ( n15909 , n15897 , n15908 );
and ( n15910 , n15894 , n15909 );
or ( n15911 , n15893 , n15910 );
and ( n15912 , n15890 , n15911 );
or ( n15913 , n15889 , n15912 );
and ( n15914 , n15886 , n15913 );
or ( n15915 , n15885 , n15914 );
and ( n15916 , n15882 , n15915 );
or ( n15917 , n15881 , n15916 );
and ( n15918 , n15878 , n15917 );
or ( n15919 , n15877 , n15918 );
and ( n15920 , n15874 , n15919 );
or ( n15921 , n15873 , n15920 );
and ( n15922 , n15870 , n15921 );
or ( n15923 , n15869 , n15922 );
and ( n15924 , n15866 , n15923 );
or ( n15925 , n15865 , n15924 );
and ( n15926 , n15862 , n15925 );
or ( n15927 , n15861 , n15926 );
and ( n15928 , n15858 , n15927 );
or ( n15929 , n15857 , n15928 );
and ( n15930 , n15854 , n15929 );
or ( n15931 , n15853 , n15930 );
and ( n15932 , n15850 , n15931 );
or ( n15933 , n15849 , n15932 );
and ( n15934 , n15846 , n15933 );
or ( n15935 , n15845 , n15934 );
and ( n15936 , n816 , n6704 );
and ( n15937 , n15935 , n15936 );
xor ( n15938 , n15935 , n15936 );
xor ( n15939 , n15846 , n15933 );
and ( n15940 , n817 , n6704 );
and ( n15941 , n15939 , n15940 );
xor ( n15942 , n15939 , n15940 );
xor ( n15943 , n15850 , n15931 );
and ( n15944 , n818 , n6704 );
and ( n15945 , n15943 , n15944 );
xor ( n15946 , n15943 , n15944 );
xor ( n15947 , n15854 , n15929 );
and ( n15948 , n819 , n6704 );
and ( n15949 , n15947 , n15948 );
xor ( n15950 , n15947 , n15948 );
xor ( n15951 , n15858 , n15927 );
and ( n15952 , n820 , n6704 );
and ( n15953 , n15951 , n15952 );
xor ( n15954 , n15951 , n15952 );
xor ( n15955 , n15862 , n15925 );
and ( n15956 , n821 , n6704 );
and ( n15957 , n15955 , n15956 );
xor ( n15958 , n15955 , n15956 );
xor ( n15959 , n15866 , n15923 );
and ( n15960 , n822 , n6704 );
and ( n15961 , n15959 , n15960 );
xor ( n15962 , n15959 , n15960 );
xor ( n15963 , n15870 , n15921 );
and ( n15964 , n823 , n6704 );
and ( n15965 , n15963 , n15964 );
xor ( n15966 , n15963 , n15964 );
xor ( n15967 , n15874 , n15919 );
and ( n15968 , n824 , n6704 );
and ( n15969 , n15967 , n15968 );
xor ( n15970 , n15967 , n15968 );
xor ( n15971 , n15878 , n15917 );
and ( n15972 , n825 , n6704 );
and ( n15973 , n15971 , n15972 );
xor ( n15974 , n15971 , n15972 );
xor ( n15975 , n15882 , n15915 );
and ( n15976 , n826 , n6704 );
and ( n15977 , n15975 , n15976 );
xor ( n15978 , n15975 , n15976 );
xor ( n15979 , n15886 , n15913 );
and ( n15980 , n827 , n6704 );
and ( n15981 , n15979 , n15980 );
xor ( n15982 , n15979 , n15980 );
xor ( n15983 , n15890 , n15911 );
and ( n15984 , n828 , n6704 );
and ( n15985 , n15983 , n15984 );
xor ( n15986 , n15983 , n15984 );
xor ( n15987 , n15894 , n15909 );
and ( n15988 , n829 , n6704 );
and ( n15989 , n15987 , n15988 );
xor ( n15990 , n15987 , n15988 );
xor ( n15991 , n15898 , n15907 );
and ( n15992 , n830 , n6704 );
and ( n15993 , n15991 , n15992 );
xor ( n15994 , n15991 , n15992 );
xor ( n15995 , n15902 , n15905 );
and ( n15996 , n831 , n6704 );
and ( n15997 , n15995 , n15996 );
and ( n15998 , n15994 , n15997 );
or ( n15999 , n15993 , n15998 );
and ( n16000 , n15990 , n15999 );
or ( n16001 , n15989 , n16000 );
and ( n16002 , n15986 , n16001 );
or ( n16003 , n15985 , n16002 );
and ( n16004 , n15982 , n16003 );
or ( n16005 , n15981 , n16004 );
and ( n16006 , n15978 , n16005 );
or ( n16007 , n15977 , n16006 );
and ( n16008 , n15974 , n16007 );
or ( n16009 , n15973 , n16008 );
and ( n16010 , n15970 , n16009 );
or ( n16011 , n15969 , n16010 );
and ( n16012 , n15966 , n16011 );
or ( n16013 , n15965 , n16012 );
and ( n16014 , n15962 , n16013 );
or ( n16015 , n15961 , n16014 );
and ( n16016 , n15958 , n16015 );
or ( n16017 , n15957 , n16016 );
and ( n16018 , n15954 , n16017 );
or ( n16019 , n15953 , n16018 );
and ( n16020 , n15950 , n16019 );
or ( n16021 , n15949 , n16020 );
and ( n16022 , n15946 , n16021 );
or ( n16023 , n15945 , n16022 );
and ( n16024 , n15942 , n16023 );
or ( n16025 , n15941 , n16024 );
and ( n16026 , n15938 , n16025 );
or ( n16027 , n15937 , n16026 );
and ( n16028 , n816 , n6701 );
and ( n16029 , n16027 , n16028 );
xor ( n16030 , n16027 , n16028 );
xor ( n16031 , n15938 , n16025 );
and ( n16032 , n817 , n6701 );
and ( n16033 , n16031 , n16032 );
xor ( n16034 , n16031 , n16032 );
xor ( n16035 , n15942 , n16023 );
and ( n16036 , n818 , n6701 );
and ( n16037 , n16035 , n16036 );
xor ( n16038 , n16035 , n16036 );
xor ( n16039 , n15946 , n16021 );
and ( n16040 , n819 , n6701 );
and ( n16041 , n16039 , n16040 );
xor ( n16042 , n16039 , n16040 );
xor ( n16043 , n15950 , n16019 );
and ( n16044 , n820 , n6701 );
and ( n16045 , n16043 , n16044 );
xor ( n16046 , n16043 , n16044 );
xor ( n16047 , n15954 , n16017 );
and ( n16048 , n821 , n6701 );
and ( n16049 , n16047 , n16048 );
xor ( n16050 , n16047 , n16048 );
xor ( n16051 , n15958 , n16015 );
and ( n16052 , n822 , n6701 );
and ( n16053 , n16051 , n16052 );
xor ( n16054 , n16051 , n16052 );
xor ( n16055 , n15962 , n16013 );
and ( n16056 , n823 , n6701 );
and ( n16057 , n16055 , n16056 );
xor ( n16058 , n16055 , n16056 );
xor ( n16059 , n15966 , n16011 );
and ( n16060 , n824 , n6701 );
and ( n16061 , n16059 , n16060 );
xor ( n16062 , n16059 , n16060 );
xor ( n16063 , n15970 , n16009 );
and ( n16064 , n825 , n6701 );
and ( n16065 , n16063 , n16064 );
xor ( n16066 , n16063 , n16064 );
xor ( n16067 , n15974 , n16007 );
and ( n16068 , n826 , n6701 );
and ( n16069 , n16067 , n16068 );
xor ( n16070 , n16067 , n16068 );
xor ( n16071 , n15978 , n16005 );
and ( n16072 , n827 , n6701 );
and ( n16073 , n16071 , n16072 );
xor ( n16074 , n16071 , n16072 );
xor ( n16075 , n15982 , n16003 );
and ( n16076 , n828 , n6701 );
and ( n16077 , n16075 , n16076 );
xor ( n16078 , n16075 , n16076 );
xor ( n16079 , n15986 , n16001 );
and ( n16080 , n829 , n6701 );
and ( n16081 , n16079 , n16080 );
xor ( n16082 , n16079 , n16080 );
xor ( n16083 , n15990 , n15999 );
and ( n16084 , n830 , n6701 );
and ( n16085 , n16083 , n16084 );
xor ( n16086 , n16083 , n16084 );
xor ( n16087 , n15994 , n15997 );
and ( n16088 , n831 , n6701 );
and ( n16089 , n16087 , n16088 );
and ( n16090 , n16086 , n16089 );
or ( n16091 , n16085 , n16090 );
and ( n16092 , n16082 , n16091 );
or ( n16093 , n16081 , n16092 );
and ( n16094 , n16078 , n16093 );
or ( n16095 , n16077 , n16094 );
and ( n16096 , n16074 , n16095 );
or ( n16097 , n16073 , n16096 );
and ( n16098 , n16070 , n16097 );
or ( n16099 , n16069 , n16098 );
and ( n16100 , n16066 , n16099 );
or ( n16101 , n16065 , n16100 );
and ( n16102 , n16062 , n16101 );
or ( n16103 , n16061 , n16102 );
and ( n16104 , n16058 , n16103 );
or ( n16105 , n16057 , n16104 );
and ( n16106 , n16054 , n16105 );
or ( n16107 , n16053 , n16106 );
and ( n16108 , n16050 , n16107 );
or ( n16109 , n16049 , n16108 );
and ( n16110 , n16046 , n16109 );
or ( n16111 , n16045 , n16110 );
and ( n16112 , n16042 , n16111 );
or ( n16113 , n16041 , n16112 );
and ( n16114 , n16038 , n16113 );
or ( n16115 , n16037 , n16114 );
and ( n16116 , n16034 , n16115 );
or ( n16117 , n16033 , n16116 );
and ( n16118 , n16030 , n16117 );
or ( n16119 , n16029 , n16118 );
and ( n16120 , n816 , n6698 );
and ( n16121 , n16119 , n16120 );
xor ( n16122 , n16119 , n16120 );
xor ( n16123 , n16030 , n16117 );
and ( n16124 , n817 , n6698 );
and ( n16125 , n16123 , n16124 );
xor ( n16126 , n16123 , n16124 );
xor ( n16127 , n16034 , n16115 );
and ( n16128 , n818 , n6698 );
and ( n16129 , n16127 , n16128 );
xor ( n16130 , n16127 , n16128 );
xor ( n16131 , n16038 , n16113 );
and ( n16132 , n819 , n6698 );
and ( n16133 , n16131 , n16132 );
xor ( n16134 , n16131 , n16132 );
xor ( n16135 , n16042 , n16111 );
and ( n16136 , n820 , n6698 );
and ( n16137 , n16135 , n16136 );
xor ( n16138 , n16135 , n16136 );
xor ( n16139 , n16046 , n16109 );
and ( n16140 , n821 , n6698 );
and ( n16141 , n16139 , n16140 );
xor ( n16142 , n16139 , n16140 );
xor ( n16143 , n16050 , n16107 );
and ( n16144 , n822 , n6698 );
and ( n16145 , n16143 , n16144 );
xor ( n16146 , n16143 , n16144 );
xor ( n16147 , n16054 , n16105 );
and ( n16148 , n823 , n6698 );
and ( n16149 , n16147 , n16148 );
xor ( n16150 , n16147 , n16148 );
xor ( n16151 , n16058 , n16103 );
and ( n16152 , n824 , n6698 );
and ( n16153 , n16151 , n16152 );
xor ( n16154 , n16151 , n16152 );
xor ( n16155 , n16062 , n16101 );
and ( n16156 , n825 , n6698 );
and ( n16157 , n16155 , n16156 );
xor ( n16158 , n16155 , n16156 );
xor ( n16159 , n16066 , n16099 );
and ( n16160 , n826 , n6698 );
and ( n16161 , n16159 , n16160 );
xor ( n16162 , n16159 , n16160 );
xor ( n16163 , n16070 , n16097 );
and ( n16164 , n827 , n6698 );
and ( n16165 , n16163 , n16164 );
xor ( n16166 , n16163 , n16164 );
xor ( n16167 , n16074 , n16095 );
and ( n16168 , n828 , n6698 );
and ( n16169 , n16167 , n16168 );
xor ( n16170 , n16167 , n16168 );
xor ( n16171 , n16078 , n16093 );
and ( n16172 , n829 , n6698 );
and ( n16173 , n16171 , n16172 );
xor ( n16174 , n16171 , n16172 );
xor ( n16175 , n16082 , n16091 );
and ( n16176 , n830 , n6698 );
and ( n16177 , n16175 , n16176 );
xor ( n16178 , n16175 , n16176 );
xor ( n16179 , n16086 , n16089 );
and ( n16180 , n831 , n6698 );
and ( n16181 , n16179 , n16180 );
and ( n16182 , n16178 , n16181 );
or ( n16183 , n16177 , n16182 );
and ( n16184 , n16174 , n16183 );
or ( n16185 , n16173 , n16184 );
and ( n16186 , n16170 , n16185 );
or ( n16187 , n16169 , n16186 );
and ( n16188 , n16166 , n16187 );
or ( n16189 , n16165 , n16188 );
and ( n16190 , n16162 , n16189 );
or ( n16191 , n16161 , n16190 );
and ( n16192 , n16158 , n16191 );
or ( n16193 , n16157 , n16192 );
and ( n16194 , n16154 , n16193 );
or ( n16195 , n16153 , n16194 );
and ( n16196 , n16150 , n16195 );
or ( n16197 , n16149 , n16196 );
and ( n16198 , n16146 , n16197 );
or ( n16199 , n16145 , n16198 );
and ( n16200 , n16142 , n16199 );
or ( n16201 , n16141 , n16200 );
and ( n16202 , n16138 , n16201 );
or ( n16203 , n16137 , n16202 );
and ( n16204 , n16134 , n16203 );
or ( n16205 , n16133 , n16204 );
and ( n16206 , n16130 , n16205 );
or ( n16207 , n16129 , n16206 );
and ( n16208 , n16126 , n16207 );
or ( n16209 , n16125 , n16208 );
and ( n16210 , n16122 , n16209 );
or ( n16211 , n16121 , n16210 );
and ( n16212 , n816 , n6695 );
and ( n16213 , n16211 , n16212 );
xor ( n16214 , n16211 , n16212 );
xor ( n16215 , n16122 , n16209 );
and ( n16216 , n817 , n6695 );
and ( n16217 , n16215 , n16216 );
xor ( n16218 , n16215 , n16216 );
xor ( n16219 , n16126 , n16207 );
and ( n16220 , n818 , n6695 );
and ( n16221 , n16219 , n16220 );
xor ( n16222 , n16219 , n16220 );
xor ( n16223 , n16130 , n16205 );
and ( n16224 , n819 , n6695 );
and ( n16225 , n16223 , n16224 );
xor ( n16226 , n16223 , n16224 );
xor ( n16227 , n16134 , n16203 );
and ( n16228 , n820 , n6695 );
and ( n16229 , n16227 , n16228 );
xor ( n16230 , n16227 , n16228 );
xor ( n16231 , n16138 , n16201 );
and ( n16232 , n821 , n6695 );
and ( n16233 , n16231 , n16232 );
xor ( n16234 , n16231 , n16232 );
xor ( n16235 , n16142 , n16199 );
and ( n16236 , n822 , n6695 );
and ( n16237 , n16235 , n16236 );
xor ( n16238 , n16235 , n16236 );
xor ( n16239 , n16146 , n16197 );
and ( n16240 , n823 , n6695 );
and ( n16241 , n16239 , n16240 );
xor ( n16242 , n16239 , n16240 );
xor ( n16243 , n16150 , n16195 );
and ( n16244 , n824 , n6695 );
and ( n16245 , n16243 , n16244 );
xor ( n16246 , n16243 , n16244 );
xor ( n16247 , n16154 , n16193 );
and ( n16248 , n825 , n6695 );
and ( n16249 , n16247 , n16248 );
xor ( n16250 , n16247 , n16248 );
xor ( n16251 , n16158 , n16191 );
and ( n16252 , n826 , n6695 );
and ( n16253 , n16251 , n16252 );
xor ( n16254 , n16251 , n16252 );
xor ( n16255 , n16162 , n16189 );
and ( n16256 , n827 , n6695 );
and ( n16257 , n16255 , n16256 );
xor ( n16258 , n16255 , n16256 );
xor ( n16259 , n16166 , n16187 );
and ( n16260 , n828 , n6695 );
and ( n16261 , n16259 , n16260 );
xor ( n16262 , n16259 , n16260 );
xor ( n16263 , n16170 , n16185 );
and ( n16264 , n829 , n6695 );
and ( n16265 , n16263 , n16264 );
xor ( n16266 , n16263 , n16264 );
xor ( n16267 , n16174 , n16183 );
and ( n16268 , n830 , n6695 );
and ( n16269 , n16267 , n16268 );
xor ( n16270 , n16267 , n16268 );
xor ( n16271 , n16178 , n16181 );
and ( n16272 , n831 , n6695 );
and ( n16273 , n16271 , n16272 );
and ( n16274 , n16270 , n16273 );
or ( n16275 , n16269 , n16274 );
and ( n16276 , n16266 , n16275 );
or ( n16277 , n16265 , n16276 );
and ( n16278 , n16262 , n16277 );
or ( n16279 , n16261 , n16278 );
and ( n16280 , n16258 , n16279 );
or ( n16281 , n16257 , n16280 );
and ( n16282 , n16254 , n16281 );
or ( n16283 , n16253 , n16282 );
and ( n16284 , n16250 , n16283 );
or ( n16285 , n16249 , n16284 );
and ( n16286 , n16246 , n16285 );
or ( n16287 , n16245 , n16286 );
and ( n16288 , n16242 , n16287 );
or ( n16289 , n16241 , n16288 );
and ( n16290 , n16238 , n16289 );
or ( n16291 , n16237 , n16290 );
and ( n16292 , n16234 , n16291 );
or ( n16293 , n16233 , n16292 );
and ( n16294 , n16230 , n16293 );
or ( n16295 , n16229 , n16294 );
and ( n16296 , n16226 , n16295 );
or ( n16297 , n16225 , n16296 );
and ( n16298 , n16222 , n16297 );
or ( n16299 , n16221 , n16298 );
and ( n16300 , n16218 , n16299 );
or ( n16301 , n16217 , n16300 );
and ( n16302 , n16214 , n16301 );
or ( n16303 , n16213 , n16302 );
and ( n16304 , n816 , n6692 );
and ( n16305 , n16303 , n16304 );
xor ( n16306 , n16303 , n16304 );
xor ( n16307 , n16214 , n16301 );
and ( n16308 , n817 , n6692 );
and ( n16309 , n16307 , n16308 );
xor ( n16310 , n16307 , n16308 );
xor ( n16311 , n16218 , n16299 );
and ( n16312 , n818 , n6692 );
and ( n16313 , n16311 , n16312 );
xor ( n16314 , n16311 , n16312 );
xor ( n16315 , n16222 , n16297 );
and ( n16316 , n819 , n6692 );
and ( n16317 , n16315 , n16316 );
xor ( n16318 , n16315 , n16316 );
xor ( n16319 , n16226 , n16295 );
and ( n16320 , n820 , n6692 );
and ( n16321 , n16319 , n16320 );
xor ( n16322 , n16319 , n16320 );
xor ( n16323 , n16230 , n16293 );
and ( n16324 , n821 , n6692 );
and ( n16325 , n16323 , n16324 );
xor ( n16326 , n16323 , n16324 );
xor ( n16327 , n16234 , n16291 );
and ( n16328 , n822 , n6692 );
and ( n16329 , n16327 , n16328 );
xor ( n16330 , n16327 , n16328 );
xor ( n16331 , n16238 , n16289 );
and ( n16332 , n823 , n6692 );
and ( n16333 , n16331 , n16332 );
xor ( n16334 , n16331 , n16332 );
xor ( n16335 , n16242 , n16287 );
and ( n16336 , n824 , n6692 );
and ( n16337 , n16335 , n16336 );
xor ( n16338 , n16335 , n16336 );
xor ( n16339 , n16246 , n16285 );
and ( n16340 , n825 , n6692 );
and ( n16341 , n16339 , n16340 );
xor ( n16342 , n16339 , n16340 );
xor ( n16343 , n16250 , n16283 );
and ( n16344 , n826 , n6692 );
and ( n16345 , n16343 , n16344 );
xor ( n16346 , n16343 , n16344 );
xor ( n16347 , n16254 , n16281 );
and ( n16348 , n827 , n6692 );
and ( n16349 , n16347 , n16348 );
xor ( n16350 , n16347 , n16348 );
xor ( n16351 , n16258 , n16279 );
and ( n16352 , n828 , n6692 );
and ( n16353 , n16351 , n16352 );
xor ( n16354 , n16351 , n16352 );
xor ( n16355 , n16262 , n16277 );
and ( n16356 , n829 , n6692 );
and ( n16357 , n16355 , n16356 );
xor ( n16358 , n16355 , n16356 );
xor ( n16359 , n16266 , n16275 );
and ( n16360 , n830 , n6692 );
and ( n16361 , n16359 , n16360 );
xor ( n16362 , n16359 , n16360 );
xor ( n16363 , n16270 , n16273 );
and ( n16364 , n831 , n6692 );
and ( n16365 , n16363 , n16364 );
and ( n16366 , n16362 , n16365 );
or ( n16367 , n16361 , n16366 );
and ( n16368 , n16358 , n16367 );
or ( n16369 , n16357 , n16368 );
and ( n16370 , n16354 , n16369 );
or ( n16371 , n16353 , n16370 );
and ( n16372 , n16350 , n16371 );
or ( n16373 , n16349 , n16372 );
and ( n16374 , n16346 , n16373 );
or ( n16375 , n16345 , n16374 );
and ( n16376 , n16342 , n16375 );
or ( n16377 , n16341 , n16376 );
and ( n16378 , n16338 , n16377 );
or ( n16379 , n16337 , n16378 );
and ( n16380 , n16334 , n16379 );
or ( n16381 , n16333 , n16380 );
and ( n16382 , n16330 , n16381 );
or ( n16383 , n16329 , n16382 );
and ( n16384 , n16326 , n16383 );
or ( n16385 , n16325 , n16384 );
and ( n16386 , n16322 , n16385 );
or ( n16387 , n16321 , n16386 );
and ( n16388 , n16318 , n16387 );
or ( n16389 , n16317 , n16388 );
and ( n16390 , n16314 , n16389 );
or ( n16391 , n16313 , n16390 );
and ( n16392 , n16310 , n16391 );
or ( n16393 , n16309 , n16392 );
and ( n16394 , n16306 , n16393 );
or ( n16395 , n16305 , n16394 );
and ( n16396 , n816 , n6689 );
and ( n16397 , n16395 , n16396 );
xor ( n16398 , n16395 , n16396 );
xor ( n16399 , n16306 , n16393 );
and ( n16400 , n817 , n6689 );
and ( n16401 , n16399 , n16400 );
xor ( n16402 , n16399 , n16400 );
xor ( n16403 , n16310 , n16391 );
and ( n16404 , n818 , n6689 );
and ( n16405 , n16403 , n16404 );
xor ( n16406 , n16403 , n16404 );
xor ( n16407 , n16314 , n16389 );
and ( n16408 , n819 , n6689 );
and ( n16409 , n16407 , n16408 );
xor ( n16410 , n16407 , n16408 );
xor ( n16411 , n16318 , n16387 );
and ( n16412 , n820 , n6689 );
and ( n16413 , n16411 , n16412 );
xor ( n16414 , n16411 , n16412 );
xor ( n16415 , n16322 , n16385 );
and ( n16416 , n821 , n6689 );
and ( n16417 , n16415 , n16416 );
xor ( n16418 , n16415 , n16416 );
xor ( n16419 , n16326 , n16383 );
and ( n16420 , n822 , n6689 );
and ( n16421 , n16419 , n16420 );
xor ( n16422 , n16419 , n16420 );
xor ( n16423 , n16330 , n16381 );
and ( n16424 , n823 , n6689 );
and ( n16425 , n16423 , n16424 );
xor ( n16426 , n16423 , n16424 );
xor ( n16427 , n16334 , n16379 );
and ( n16428 , n824 , n6689 );
and ( n16429 , n16427 , n16428 );
xor ( n16430 , n16427 , n16428 );
xor ( n16431 , n16338 , n16377 );
and ( n16432 , n825 , n6689 );
and ( n16433 , n16431 , n16432 );
xor ( n16434 , n16431 , n16432 );
xor ( n16435 , n16342 , n16375 );
and ( n16436 , n826 , n6689 );
and ( n16437 , n16435 , n16436 );
xor ( n16438 , n16435 , n16436 );
xor ( n16439 , n16346 , n16373 );
and ( n16440 , n827 , n6689 );
and ( n16441 , n16439 , n16440 );
xor ( n16442 , n16439 , n16440 );
xor ( n16443 , n16350 , n16371 );
and ( n16444 , n828 , n6689 );
and ( n16445 , n16443 , n16444 );
xor ( n16446 , n16443 , n16444 );
xor ( n16447 , n16354 , n16369 );
and ( n16448 , n829 , n6689 );
and ( n16449 , n16447 , n16448 );
xor ( n16450 , n16447 , n16448 );
xor ( n16451 , n16358 , n16367 );
and ( n16452 , n830 , n6689 );
and ( n16453 , n16451 , n16452 );
xor ( n16454 , n16451 , n16452 );
xor ( n16455 , n16362 , n16365 );
and ( n16456 , n831 , n6689 );
and ( n16457 , n16455 , n16456 );
and ( n16458 , n16454 , n16457 );
or ( n16459 , n16453 , n16458 );
and ( n16460 , n16450 , n16459 );
or ( n16461 , n16449 , n16460 );
and ( n16462 , n16446 , n16461 );
or ( n16463 , n16445 , n16462 );
and ( n16464 , n16442 , n16463 );
or ( n16465 , n16441 , n16464 );
and ( n16466 , n16438 , n16465 );
or ( n16467 , n16437 , n16466 );
and ( n16468 , n16434 , n16467 );
or ( n16469 , n16433 , n16468 );
and ( n16470 , n16430 , n16469 );
or ( n16471 , n16429 , n16470 );
and ( n16472 , n16426 , n16471 );
or ( n16473 , n16425 , n16472 );
and ( n16474 , n16422 , n16473 );
or ( n16475 , n16421 , n16474 );
and ( n16476 , n16418 , n16475 );
or ( n16477 , n16417 , n16476 );
and ( n16478 , n16414 , n16477 );
or ( n16479 , n16413 , n16478 );
and ( n16480 , n16410 , n16479 );
or ( n16481 , n16409 , n16480 );
and ( n16482 , n16406 , n16481 );
or ( n16483 , n16405 , n16482 );
and ( n16484 , n16402 , n16483 );
or ( n16485 , n16401 , n16484 );
and ( n16486 , n16398 , n16485 );
or ( n16487 , n16397 , n16486 );
and ( n16488 , n816 , n6686 );
and ( n16489 , n16487 , n16488 );
xor ( n16490 , n16487 , n16488 );
xor ( n16491 , n16398 , n16485 );
and ( n16492 , n817 , n6686 );
and ( n16493 , n16491 , n16492 );
xor ( n16494 , n16491 , n16492 );
xor ( n16495 , n16402 , n16483 );
and ( n16496 , n818 , n6686 );
and ( n16497 , n16495 , n16496 );
xor ( n16498 , n16495 , n16496 );
xor ( n16499 , n16406 , n16481 );
and ( n16500 , n819 , n6686 );
and ( n16501 , n16499 , n16500 );
xor ( n16502 , n16499 , n16500 );
xor ( n16503 , n16410 , n16479 );
and ( n16504 , n820 , n6686 );
and ( n16505 , n16503 , n16504 );
xor ( n16506 , n16503 , n16504 );
xor ( n16507 , n16414 , n16477 );
and ( n16508 , n821 , n6686 );
and ( n16509 , n16507 , n16508 );
xor ( n16510 , n16507 , n16508 );
xor ( n16511 , n16418 , n16475 );
and ( n16512 , n822 , n6686 );
and ( n16513 , n16511 , n16512 );
xor ( n16514 , n16511 , n16512 );
xor ( n16515 , n16422 , n16473 );
and ( n16516 , n823 , n6686 );
and ( n16517 , n16515 , n16516 );
xor ( n16518 , n16515 , n16516 );
xor ( n16519 , n16426 , n16471 );
and ( n16520 , n824 , n6686 );
and ( n16521 , n16519 , n16520 );
xor ( n16522 , n16519 , n16520 );
xor ( n16523 , n16430 , n16469 );
and ( n16524 , n825 , n6686 );
and ( n16525 , n16523 , n16524 );
xor ( n16526 , n16523 , n16524 );
xor ( n16527 , n16434 , n16467 );
and ( n16528 , n826 , n6686 );
and ( n16529 , n16527 , n16528 );
xor ( n16530 , n16527 , n16528 );
xor ( n16531 , n16438 , n16465 );
and ( n16532 , n827 , n6686 );
and ( n16533 , n16531 , n16532 );
xor ( n16534 , n16531 , n16532 );
xor ( n16535 , n16442 , n16463 );
and ( n16536 , n828 , n6686 );
and ( n16537 , n16535 , n16536 );
xor ( n16538 , n16535 , n16536 );
xor ( n16539 , n16446 , n16461 );
and ( n16540 , n829 , n6686 );
and ( n16541 , n16539 , n16540 );
xor ( n16542 , n16539 , n16540 );
xor ( n16543 , n16450 , n16459 );
and ( n16544 , n830 , n6686 );
and ( n16545 , n16543 , n16544 );
xor ( n16546 , n16543 , n16544 );
xor ( n16547 , n16454 , n16457 );
and ( n16548 , n831 , n6686 );
and ( n16549 , n16547 , n16548 );
and ( n16550 , n16546 , n16549 );
or ( n16551 , n16545 , n16550 );
and ( n16552 , n16542 , n16551 );
or ( n16553 , n16541 , n16552 );
and ( n16554 , n16538 , n16553 );
or ( n16555 , n16537 , n16554 );
and ( n16556 , n16534 , n16555 );
or ( n16557 , n16533 , n16556 );
and ( n16558 , n16530 , n16557 );
or ( n16559 , n16529 , n16558 );
and ( n16560 , n16526 , n16559 );
or ( n16561 , n16525 , n16560 );
and ( n16562 , n16522 , n16561 );
or ( n16563 , n16521 , n16562 );
and ( n16564 , n16518 , n16563 );
or ( n16565 , n16517 , n16564 );
and ( n16566 , n16514 , n16565 );
or ( n16567 , n16513 , n16566 );
and ( n16568 , n16510 , n16567 );
or ( n16569 , n16509 , n16568 );
and ( n16570 , n16506 , n16569 );
or ( n16571 , n16505 , n16570 );
and ( n16572 , n16502 , n16571 );
or ( n16573 , n16501 , n16572 );
and ( n16574 , n16498 , n16573 );
or ( n16575 , n16497 , n16574 );
and ( n16576 , n16494 , n16575 );
or ( n16577 , n16493 , n16576 );
and ( n16578 , n16490 , n16577 );
or ( n16579 , n16489 , n16578 );
and ( n16580 , n816 , n6683 );
and ( n16581 , n16579 , n16580 );
xor ( n16582 , n16579 , n16580 );
xor ( n16583 , n16490 , n16577 );
and ( n16584 , n817 , n6683 );
and ( n16585 , n16583 , n16584 );
xor ( n16586 , n16583 , n16584 );
xor ( n16587 , n16494 , n16575 );
and ( n16588 , n818 , n6683 );
and ( n16589 , n16587 , n16588 );
xor ( n16590 , n16587 , n16588 );
xor ( n16591 , n16498 , n16573 );
and ( n16592 , n819 , n6683 );
and ( n16593 , n16591 , n16592 );
xor ( n16594 , n16591 , n16592 );
xor ( n16595 , n16502 , n16571 );
and ( n16596 , n820 , n6683 );
and ( n16597 , n16595 , n16596 );
xor ( n16598 , n16595 , n16596 );
xor ( n16599 , n16506 , n16569 );
and ( n16600 , n821 , n6683 );
and ( n16601 , n16599 , n16600 );
xor ( n16602 , n16599 , n16600 );
xor ( n16603 , n16510 , n16567 );
and ( n16604 , n822 , n6683 );
and ( n16605 , n16603 , n16604 );
xor ( n16606 , n16603 , n16604 );
xor ( n16607 , n16514 , n16565 );
and ( n16608 , n823 , n6683 );
and ( n16609 , n16607 , n16608 );
xor ( n16610 , n16607 , n16608 );
xor ( n16611 , n16518 , n16563 );
and ( n16612 , n824 , n6683 );
and ( n16613 , n16611 , n16612 );
xor ( n16614 , n16611 , n16612 );
xor ( n16615 , n16522 , n16561 );
and ( n16616 , n825 , n6683 );
and ( n16617 , n16615 , n16616 );
xor ( n16618 , n16615 , n16616 );
xor ( n16619 , n16526 , n16559 );
and ( n16620 , n826 , n6683 );
and ( n16621 , n16619 , n16620 );
xor ( n16622 , n16619 , n16620 );
xor ( n16623 , n16530 , n16557 );
and ( n16624 , n827 , n6683 );
and ( n16625 , n16623 , n16624 );
xor ( n16626 , n16623 , n16624 );
xor ( n16627 , n16534 , n16555 );
and ( n16628 , n828 , n6683 );
and ( n16629 , n16627 , n16628 );
xor ( n16630 , n16627 , n16628 );
xor ( n16631 , n16538 , n16553 );
and ( n16632 , n829 , n6683 );
and ( n16633 , n16631 , n16632 );
xor ( n16634 , n16631 , n16632 );
xor ( n16635 , n16542 , n16551 );
and ( n16636 , n830 , n6683 );
and ( n16637 , n16635 , n16636 );
xor ( n16638 , n16635 , n16636 );
xor ( n16639 , n16546 , n16549 );
and ( n16640 , n831 , n6683 );
and ( n16641 , n16639 , n16640 );
and ( n16642 , n16638 , n16641 );
or ( n16643 , n16637 , n16642 );
and ( n16644 , n16634 , n16643 );
or ( n16645 , n16633 , n16644 );
and ( n16646 , n16630 , n16645 );
or ( n16647 , n16629 , n16646 );
and ( n16648 , n16626 , n16647 );
or ( n16649 , n16625 , n16648 );
and ( n16650 , n16622 , n16649 );
or ( n16651 , n16621 , n16650 );
and ( n16652 , n16618 , n16651 );
or ( n16653 , n16617 , n16652 );
and ( n16654 , n16614 , n16653 );
or ( n16655 , n16613 , n16654 );
and ( n16656 , n16610 , n16655 );
or ( n16657 , n16609 , n16656 );
and ( n16658 , n16606 , n16657 );
or ( n16659 , n16605 , n16658 );
and ( n16660 , n16602 , n16659 );
or ( n16661 , n16601 , n16660 );
and ( n16662 , n16598 , n16661 );
or ( n16663 , n16597 , n16662 );
and ( n16664 , n16594 , n16663 );
or ( n16665 , n16593 , n16664 );
and ( n16666 , n16590 , n16665 );
or ( n16667 , n16589 , n16666 );
and ( n16668 , n16586 , n16667 );
or ( n16669 , n16585 , n16668 );
and ( n16670 , n16582 , n16669 );
or ( n16671 , n16581 , n16670 );
and ( n16672 , n816 , n6680 );
and ( n16673 , n16671 , n16672 );
xor ( n16674 , n16671 , n16672 );
xor ( n16675 , n16582 , n16669 );
and ( n16676 , n817 , n6680 );
and ( n16677 , n16675 , n16676 );
xor ( n16678 , n16675 , n16676 );
xor ( n16679 , n16586 , n16667 );
and ( n16680 , n818 , n6680 );
and ( n16681 , n16679 , n16680 );
xor ( n16682 , n16679 , n16680 );
xor ( n16683 , n16590 , n16665 );
and ( n16684 , n819 , n6680 );
and ( n16685 , n16683 , n16684 );
xor ( n16686 , n16683 , n16684 );
xor ( n16687 , n16594 , n16663 );
and ( n16688 , n820 , n6680 );
and ( n16689 , n16687 , n16688 );
xor ( n16690 , n16687 , n16688 );
xor ( n16691 , n16598 , n16661 );
and ( n16692 , n821 , n6680 );
and ( n16693 , n16691 , n16692 );
xor ( n16694 , n16691 , n16692 );
xor ( n16695 , n16602 , n16659 );
and ( n16696 , n822 , n6680 );
and ( n16697 , n16695 , n16696 );
xor ( n16698 , n16695 , n16696 );
xor ( n16699 , n16606 , n16657 );
and ( n16700 , n823 , n6680 );
and ( n16701 , n16699 , n16700 );
xor ( n16702 , n16699 , n16700 );
xor ( n16703 , n16610 , n16655 );
and ( n16704 , n824 , n6680 );
and ( n16705 , n16703 , n16704 );
xor ( n16706 , n16703 , n16704 );
xor ( n16707 , n16614 , n16653 );
and ( n16708 , n825 , n6680 );
and ( n16709 , n16707 , n16708 );
xor ( n16710 , n16707 , n16708 );
xor ( n16711 , n16618 , n16651 );
and ( n16712 , n826 , n6680 );
and ( n16713 , n16711 , n16712 );
xor ( n16714 , n16711 , n16712 );
xor ( n16715 , n16622 , n16649 );
and ( n16716 , n827 , n6680 );
and ( n16717 , n16715 , n16716 );
xor ( n16718 , n16715 , n16716 );
xor ( n16719 , n16626 , n16647 );
and ( n16720 , n828 , n6680 );
and ( n16721 , n16719 , n16720 );
xor ( n16722 , n16719 , n16720 );
xor ( n16723 , n16630 , n16645 );
and ( n16724 , n829 , n6680 );
and ( n16725 , n16723 , n16724 );
xor ( n16726 , n16723 , n16724 );
xor ( n16727 , n16634 , n16643 );
and ( n16728 , n830 , n6680 );
and ( n16729 , n16727 , n16728 );
xor ( n16730 , n16727 , n16728 );
xor ( n16731 , n16638 , n16641 );
and ( n16732 , n831 , n6680 );
and ( n16733 , n16731 , n16732 );
and ( n16734 , n16730 , n16733 );
or ( n16735 , n16729 , n16734 );
and ( n16736 , n16726 , n16735 );
or ( n16737 , n16725 , n16736 );
and ( n16738 , n16722 , n16737 );
or ( n16739 , n16721 , n16738 );
and ( n16740 , n16718 , n16739 );
or ( n16741 , n16717 , n16740 );
and ( n16742 , n16714 , n16741 );
or ( n16743 , n16713 , n16742 );
and ( n16744 , n16710 , n16743 );
or ( n16745 , n16709 , n16744 );
and ( n16746 , n16706 , n16745 );
or ( n16747 , n16705 , n16746 );
and ( n16748 , n16702 , n16747 );
or ( n16749 , n16701 , n16748 );
and ( n16750 , n16698 , n16749 );
or ( n16751 , n16697 , n16750 );
and ( n16752 , n16694 , n16751 );
or ( n16753 , n16693 , n16752 );
and ( n16754 , n16690 , n16753 );
or ( n16755 , n16689 , n16754 );
and ( n16756 , n16686 , n16755 );
or ( n16757 , n16685 , n16756 );
and ( n16758 , n16682 , n16757 );
or ( n16759 , n16681 , n16758 );
and ( n16760 , n16678 , n16759 );
or ( n16761 , n16677 , n16760 );
and ( n16762 , n16674 , n16761 );
or ( n16763 , n16673 , n16762 );
and ( n16764 , n816 , n6677 );
and ( n16765 , n16763 , n16764 );
xor ( n16766 , n16763 , n16764 );
xor ( n16767 , n16674 , n16761 );
and ( n16768 , n817 , n6677 );
and ( n16769 , n16767 , n16768 );
xor ( n16770 , n16767 , n16768 );
xor ( n16771 , n16678 , n16759 );
and ( n16772 , n818 , n6677 );
and ( n16773 , n16771 , n16772 );
xor ( n16774 , n16771 , n16772 );
xor ( n16775 , n16682 , n16757 );
and ( n16776 , n819 , n6677 );
and ( n16777 , n16775 , n16776 );
xor ( n16778 , n16775 , n16776 );
xor ( n16779 , n16686 , n16755 );
and ( n16780 , n820 , n6677 );
and ( n16781 , n16779 , n16780 );
xor ( n16782 , n16779 , n16780 );
xor ( n16783 , n16690 , n16753 );
and ( n16784 , n821 , n6677 );
and ( n16785 , n16783 , n16784 );
xor ( n16786 , n16783 , n16784 );
xor ( n16787 , n16694 , n16751 );
and ( n16788 , n822 , n6677 );
and ( n16789 , n16787 , n16788 );
xor ( n16790 , n16787 , n16788 );
xor ( n16791 , n16698 , n16749 );
and ( n16792 , n823 , n6677 );
and ( n16793 , n16791 , n16792 );
xor ( n16794 , n16791 , n16792 );
xor ( n16795 , n16702 , n16747 );
and ( n16796 , n824 , n6677 );
and ( n16797 , n16795 , n16796 );
xor ( n16798 , n16795 , n16796 );
xor ( n16799 , n16706 , n16745 );
and ( n16800 , n825 , n6677 );
and ( n16801 , n16799 , n16800 );
xor ( n16802 , n16799 , n16800 );
xor ( n16803 , n16710 , n16743 );
and ( n16804 , n826 , n6677 );
and ( n16805 , n16803 , n16804 );
xor ( n16806 , n16803 , n16804 );
xor ( n16807 , n16714 , n16741 );
and ( n16808 , n827 , n6677 );
and ( n16809 , n16807 , n16808 );
xor ( n16810 , n16807 , n16808 );
xor ( n16811 , n16718 , n16739 );
and ( n16812 , n828 , n6677 );
and ( n16813 , n16811 , n16812 );
xor ( n16814 , n16811 , n16812 );
xor ( n16815 , n16722 , n16737 );
and ( n16816 , n829 , n6677 );
and ( n16817 , n16815 , n16816 );
xor ( n16818 , n16815 , n16816 );
xor ( n16819 , n16726 , n16735 );
and ( n16820 , n830 , n6677 );
and ( n16821 , n16819 , n16820 );
xor ( n16822 , n16819 , n16820 );
xor ( n16823 , n16730 , n16733 );
and ( n16824 , n831 , n6677 );
and ( n16825 , n16823 , n16824 );
and ( n16826 , n16822 , n16825 );
or ( n16827 , n16821 , n16826 );
and ( n16828 , n16818 , n16827 );
or ( n16829 , n16817 , n16828 );
and ( n16830 , n16814 , n16829 );
or ( n16831 , n16813 , n16830 );
and ( n16832 , n16810 , n16831 );
or ( n16833 , n16809 , n16832 );
and ( n16834 , n16806 , n16833 );
or ( n16835 , n16805 , n16834 );
and ( n16836 , n16802 , n16835 );
or ( n16837 , n16801 , n16836 );
and ( n16838 , n16798 , n16837 );
or ( n16839 , n16797 , n16838 );
and ( n16840 , n16794 , n16839 );
or ( n16841 , n16793 , n16840 );
and ( n16842 , n16790 , n16841 );
or ( n16843 , n16789 , n16842 );
and ( n16844 , n16786 , n16843 );
or ( n16845 , n16785 , n16844 );
and ( n16846 , n16782 , n16845 );
or ( n16847 , n16781 , n16846 );
and ( n16848 , n16778 , n16847 );
or ( n16849 , n16777 , n16848 );
and ( n16850 , n16774 , n16849 );
or ( n16851 , n16773 , n16850 );
and ( n16852 , n16770 , n16851 );
or ( n16853 , n16769 , n16852 );
and ( n16854 , n16766 , n16853 );
or ( n16855 , n16765 , n16854 );
and ( n16856 , n816 , n6674 );
and ( n16857 , n16855 , n16856 );
xor ( n16858 , n16855 , n16856 );
xor ( n16859 , n16766 , n16853 );
and ( n16860 , n817 , n6674 );
and ( n16861 , n16859 , n16860 );
xor ( n16862 , n16859 , n16860 );
xor ( n16863 , n16770 , n16851 );
and ( n16864 , n818 , n6674 );
and ( n16865 , n16863 , n16864 );
xor ( n16866 , n16863 , n16864 );
xor ( n16867 , n16774 , n16849 );
and ( n16868 , n819 , n6674 );
and ( n16869 , n16867 , n16868 );
xor ( n16870 , n16867 , n16868 );
xor ( n16871 , n16778 , n16847 );
and ( n16872 , n820 , n6674 );
and ( n16873 , n16871 , n16872 );
xor ( n16874 , n16871 , n16872 );
xor ( n16875 , n16782 , n16845 );
and ( n16876 , n821 , n6674 );
and ( n16877 , n16875 , n16876 );
xor ( n16878 , n16875 , n16876 );
xor ( n16879 , n16786 , n16843 );
and ( n16880 , n822 , n6674 );
and ( n16881 , n16879 , n16880 );
xor ( n16882 , n16879 , n16880 );
xor ( n16883 , n16790 , n16841 );
and ( n16884 , n823 , n6674 );
and ( n16885 , n16883 , n16884 );
xor ( n16886 , n16883 , n16884 );
xor ( n16887 , n16794 , n16839 );
and ( n16888 , n824 , n6674 );
and ( n16889 , n16887 , n16888 );
xor ( n16890 , n16887 , n16888 );
xor ( n16891 , n16798 , n16837 );
and ( n16892 , n825 , n6674 );
and ( n16893 , n16891 , n16892 );
xor ( n16894 , n16891 , n16892 );
xor ( n16895 , n16802 , n16835 );
and ( n16896 , n826 , n6674 );
and ( n16897 , n16895 , n16896 );
xor ( n16898 , n16895 , n16896 );
xor ( n16899 , n16806 , n16833 );
and ( n16900 , n827 , n6674 );
and ( n16901 , n16899 , n16900 );
xor ( n16902 , n16899 , n16900 );
xor ( n16903 , n16810 , n16831 );
and ( n16904 , n828 , n6674 );
and ( n16905 , n16903 , n16904 );
xor ( n16906 , n16903 , n16904 );
xor ( n16907 , n16814 , n16829 );
and ( n16908 , n829 , n6674 );
and ( n16909 , n16907 , n16908 );
xor ( n16910 , n16907 , n16908 );
xor ( n16911 , n16818 , n16827 );
and ( n16912 , n830 , n6674 );
and ( n16913 , n16911 , n16912 );
xor ( n16914 , n16911 , n16912 );
xor ( n16915 , n16822 , n16825 );
and ( n16916 , n831 , n6674 );
and ( n16917 , n16915 , n16916 );
and ( n16918 , n16914 , n16917 );
or ( n16919 , n16913 , n16918 );
and ( n16920 , n16910 , n16919 );
or ( n16921 , n16909 , n16920 );
and ( n16922 , n16906 , n16921 );
or ( n16923 , n16905 , n16922 );
and ( n16924 , n16902 , n16923 );
or ( n16925 , n16901 , n16924 );
and ( n16926 , n16898 , n16925 );
or ( n16927 , n16897 , n16926 );
and ( n16928 , n16894 , n16927 );
or ( n16929 , n16893 , n16928 );
and ( n16930 , n16890 , n16929 );
or ( n16931 , n16889 , n16930 );
and ( n16932 , n16886 , n16931 );
or ( n16933 , n16885 , n16932 );
and ( n16934 , n16882 , n16933 );
or ( n16935 , n16881 , n16934 );
and ( n16936 , n16878 , n16935 );
or ( n16937 , n16877 , n16936 );
and ( n16938 , n16874 , n16937 );
or ( n16939 , n16873 , n16938 );
and ( n16940 , n16870 , n16939 );
or ( n16941 , n16869 , n16940 );
and ( n16942 , n16866 , n16941 );
or ( n16943 , n16865 , n16942 );
and ( n16944 , n16862 , n16943 );
or ( n16945 , n16861 , n16944 );
and ( n16946 , n16858 , n16945 );
or ( n16947 , n16857 , n16946 );
and ( n16948 , n816 , n6671 );
and ( n16949 , n16947 , n16948 );
xor ( n16950 , n16947 , n16948 );
xor ( n16951 , n16858 , n16945 );
and ( n16952 , n817 , n6671 );
and ( n16953 , n16951 , n16952 );
xor ( n16954 , n16951 , n16952 );
xor ( n16955 , n16862 , n16943 );
and ( n16956 , n818 , n6671 );
and ( n16957 , n16955 , n16956 );
xor ( n16958 , n16955 , n16956 );
xor ( n16959 , n16866 , n16941 );
and ( n16960 , n819 , n6671 );
and ( n16961 , n16959 , n16960 );
xor ( n16962 , n16959 , n16960 );
xor ( n16963 , n16870 , n16939 );
and ( n16964 , n820 , n6671 );
and ( n16965 , n16963 , n16964 );
xor ( n16966 , n16963 , n16964 );
xor ( n16967 , n16874 , n16937 );
and ( n16968 , n821 , n6671 );
and ( n16969 , n16967 , n16968 );
xor ( n16970 , n16967 , n16968 );
xor ( n16971 , n16878 , n16935 );
and ( n16972 , n822 , n6671 );
and ( n16973 , n16971 , n16972 );
xor ( n16974 , n16971 , n16972 );
xor ( n16975 , n16882 , n16933 );
and ( n16976 , n823 , n6671 );
and ( n16977 , n16975 , n16976 );
xor ( n16978 , n16975 , n16976 );
xor ( n16979 , n16886 , n16931 );
and ( n16980 , n824 , n6671 );
and ( n16981 , n16979 , n16980 );
xor ( n16982 , n16979 , n16980 );
xor ( n16983 , n16890 , n16929 );
and ( n16984 , n825 , n6671 );
and ( n16985 , n16983 , n16984 );
xor ( n16986 , n16983 , n16984 );
xor ( n16987 , n16894 , n16927 );
and ( n16988 , n826 , n6671 );
and ( n16989 , n16987 , n16988 );
xor ( n16990 , n16987 , n16988 );
xor ( n16991 , n16898 , n16925 );
and ( n16992 , n827 , n6671 );
and ( n16993 , n16991 , n16992 );
xor ( n16994 , n16991 , n16992 );
xor ( n16995 , n16902 , n16923 );
and ( n16996 , n828 , n6671 );
and ( n16997 , n16995 , n16996 );
xor ( n16998 , n16995 , n16996 );
xor ( n16999 , n16906 , n16921 );
and ( n17000 , n829 , n6671 );
and ( n17001 , n16999 , n17000 );
xor ( n17002 , n16999 , n17000 );
xor ( n17003 , n16910 , n16919 );
and ( n17004 , n830 , n6671 );
and ( n17005 , n17003 , n17004 );
xor ( n17006 , n17003 , n17004 );
xor ( n17007 , n16914 , n16917 );
and ( n17008 , n831 , n6671 );
and ( n17009 , n17007 , n17008 );
and ( n17010 , n17006 , n17009 );
or ( n17011 , n17005 , n17010 );
and ( n17012 , n17002 , n17011 );
or ( n17013 , n17001 , n17012 );
and ( n17014 , n16998 , n17013 );
or ( n17015 , n16997 , n17014 );
and ( n17016 , n16994 , n17015 );
or ( n17017 , n16993 , n17016 );
and ( n17018 , n16990 , n17017 );
or ( n17019 , n16989 , n17018 );
and ( n17020 , n16986 , n17019 );
or ( n17021 , n16985 , n17020 );
and ( n17022 , n16982 , n17021 );
or ( n17023 , n16981 , n17022 );
and ( n17024 , n16978 , n17023 );
or ( n17025 , n16977 , n17024 );
and ( n17026 , n16974 , n17025 );
or ( n17027 , n16973 , n17026 );
and ( n17028 , n16970 , n17027 );
or ( n17029 , n16969 , n17028 );
and ( n17030 , n16966 , n17029 );
or ( n17031 , n16965 , n17030 );
and ( n17032 , n16962 , n17031 );
or ( n17033 , n16961 , n17032 );
and ( n17034 , n16958 , n17033 );
or ( n17035 , n16957 , n17034 );
and ( n17036 , n16954 , n17035 );
or ( n17037 , n16953 , n17036 );
and ( n17038 , n16950 , n17037 );
or ( n17039 , n16949 , n17038 );
and ( n17040 , n816 , n6668 );
and ( n17041 , n17039 , n17040 );
xor ( n17042 , n17039 , n17040 );
xor ( n17043 , n16950 , n17037 );
and ( n17044 , n817 , n6668 );
and ( n17045 , n17043 , n17044 );
xor ( n17046 , n17043 , n17044 );
xor ( n17047 , n16954 , n17035 );
and ( n17048 , n818 , n6668 );
and ( n17049 , n17047 , n17048 );
xor ( n17050 , n17047 , n17048 );
xor ( n17051 , n16958 , n17033 );
and ( n17052 , n819 , n6668 );
and ( n17053 , n17051 , n17052 );
xor ( n17054 , n17051 , n17052 );
xor ( n17055 , n16962 , n17031 );
and ( n17056 , n820 , n6668 );
and ( n17057 , n17055 , n17056 );
xor ( n17058 , n17055 , n17056 );
xor ( n17059 , n16966 , n17029 );
and ( n17060 , n821 , n6668 );
and ( n17061 , n17059 , n17060 );
xor ( n17062 , n17059 , n17060 );
xor ( n17063 , n16970 , n17027 );
and ( n17064 , n822 , n6668 );
and ( n17065 , n17063 , n17064 );
xor ( n17066 , n17063 , n17064 );
xor ( n17067 , n16974 , n17025 );
and ( n17068 , n823 , n6668 );
and ( n17069 , n17067 , n17068 );
xor ( n17070 , n17067 , n17068 );
xor ( n17071 , n16978 , n17023 );
and ( n17072 , n824 , n6668 );
and ( n17073 , n17071 , n17072 );
xor ( n17074 , n17071 , n17072 );
xor ( n17075 , n16982 , n17021 );
and ( n17076 , n825 , n6668 );
and ( n17077 , n17075 , n17076 );
xor ( n17078 , n17075 , n17076 );
xor ( n17079 , n16986 , n17019 );
and ( n17080 , n826 , n6668 );
and ( n17081 , n17079 , n17080 );
xor ( n17082 , n17079 , n17080 );
xor ( n17083 , n16990 , n17017 );
and ( n17084 , n827 , n6668 );
and ( n17085 , n17083 , n17084 );
xor ( n17086 , n17083 , n17084 );
xor ( n17087 , n16994 , n17015 );
and ( n17088 , n828 , n6668 );
and ( n17089 , n17087 , n17088 );
xor ( n17090 , n17087 , n17088 );
xor ( n17091 , n16998 , n17013 );
and ( n17092 , n829 , n6668 );
and ( n17093 , n17091 , n17092 );
xor ( n17094 , n17091 , n17092 );
xor ( n17095 , n17002 , n17011 );
and ( n17096 , n830 , n6668 );
and ( n17097 , n17095 , n17096 );
xor ( n17098 , n17095 , n17096 );
xor ( n17099 , n17006 , n17009 );
and ( n17100 , n831 , n6668 );
and ( n17101 , n17099 , n17100 );
and ( n17102 , n17098 , n17101 );
or ( n17103 , n17097 , n17102 );
and ( n17104 , n17094 , n17103 );
or ( n17105 , n17093 , n17104 );
and ( n17106 , n17090 , n17105 );
or ( n17107 , n17089 , n17106 );
and ( n17108 , n17086 , n17107 );
or ( n17109 , n17085 , n17108 );
and ( n17110 , n17082 , n17109 );
or ( n17111 , n17081 , n17110 );
and ( n17112 , n17078 , n17111 );
or ( n17113 , n17077 , n17112 );
and ( n17114 , n17074 , n17113 );
or ( n17115 , n17073 , n17114 );
and ( n17116 , n17070 , n17115 );
or ( n17117 , n17069 , n17116 );
and ( n17118 , n17066 , n17117 );
or ( n17119 , n17065 , n17118 );
and ( n17120 , n17062 , n17119 );
or ( n17121 , n17061 , n17120 );
and ( n17122 , n17058 , n17121 );
or ( n17123 , n17057 , n17122 );
and ( n17124 , n17054 , n17123 );
or ( n17125 , n17053 , n17124 );
and ( n17126 , n17050 , n17125 );
or ( n17127 , n17049 , n17126 );
and ( n17128 , n17046 , n17127 );
or ( n17129 , n17045 , n17128 );
and ( n17130 , n17042 , n17129 );
or ( n17131 , n17041 , n17130 );
and ( n17132 , n816 , n6665 );
xor ( n17133 , n17131 , n17132 );
xor ( n17134 , n17042 , n17129 );
and ( n17135 , n817 , n6665 );
and ( n17136 , n17134 , n17135 );
xor ( n17137 , n17134 , n17135 );
xor ( n17138 , n17046 , n17127 );
and ( n17139 , n818 , n6665 );
and ( n17140 , n17138 , n17139 );
xor ( n17141 , n17138 , n17139 );
xor ( n17142 , n17050 , n17125 );
and ( n17143 , n819 , n6665 );
and ( n17144 , n17142 , n17143 );
xor ( n17145 , n17142 , n17143 );
xor ( n17146 , n17054 , n17123 );
and ( n17147 , n820 , n6665 );
and ( n17148 , n17146 , n17147 );
xor ( n17149 , n17146 , n17147 );
xor ( n17150 , n17058 , n17121 );
and ( n17151 , n821 , n6665 );
and ( n17152 , n17150 , n17151 );
xor ( n17153 , n17150 , n17151 );
xor ( n17154 , n17062 , n17119 );
and ( n17155 , n822 , n6665 );
and ( n17156 , n17154 , n17155 );
xor ( n17157 , n17154 , n17155 );
xor ( n17158 , n17066 , n17117 );
and ( n17159 , n823 , n6665 );
and ( n17160 , n17158 , n17159 );
xor ( n17161 , n17158 , n17159 );
xor ( n17162 , n17070 , n17115 );
and ( n17163 , n824 , n6665 );
and ( n17164 , n17162 , n17163 );
xor ( n17165 , n17162 , n17163 );
xor ( n17166 , n17074 , n17113 );
and ( n17167 , n825 , n6665 );
and ( n17168 , n17166 , n17167 );
xor ( n17169 , n17166 , n17167 );
xor ( n17170 , n17078 , n17111 );
and ( n17171 , n826 , n6665 );
and ( n17172 , n17170 , n17171 );
xor ( n17173 , n17170 , n17171 );
xor ( n17174 , n17082 , n17109 );
and ( n17175 , n827 , n6665 );
and ( n17176 , n17174 , n17175 );
xor ( n17177 , n17174 , n17175 );
xor ( n17178 , n17086 , n17107 );
and ( n17179 , n828 , n6665 );
and ( n17180 , n17178 , n17179 );
xor ( n17181 , n17178 , n17179 );
xor ( n17182 , n17090 , n17105 );
and ( n17183 , n829 , n6665 );
and ( n17184 , n17182 , n17183 );
xor ( n17185 , n17182 , n17183 );
xor ( n17186 , n17094 , n17103 );
and ( n17187 , n830 , n6665 );
and ( n17188 , n17186 , n17187 );
xor ( n17189 , n17186 , n17187 );
xor ( n17190 , n17098 , n17101 );
and ( n17191 , n831 , n6665 );
and ( n17192 , n17190 , n17191 );
and ( n17193 , n17189 , n17192 );
or ( n17194 , n17188 , n17193 );
and ( n17195 , n17185 , n17194 );
or ( n17196 , n17184 , n17195 );
and ( n17197 , n17181 , n17196 );
or ( n17198 , n17180 , n17197 );
and ( n17199 , n17177 , n17198 );
or ( n17200 , n17176 , n17199 );
and ( n17201 , n17173 , n17200 );
or ( n17202 , n17172 , n17201 );
and ( n17203 , n17169 , n17202 );
or ( n17204 , n17168 , n17203 );
and ( n17205 , n17165 , n17204 );
or ( n17206 , n17164 , n17205 );
and ( n17207 , n17161 , n17206 );
or ( n17208 , n17160 , n17207 );
and ( n17209 , n17157 , n17208 );
or ( n17210 , n17156 , n17209 );
and ( n17211 , n17153 , n17210 );
or ( n17212 , n17152 , n17211 );
and ( n17213 , n17149 , n17212 );
or ( n17214 , n17148 , n17213 );
and ( n17215 , n17145 , n17214 );
or ( n17216 , n17144 , n17215 );
and ( n17217 , n17141 , n17216 );
or ( n17218 , n17140 , n17217 );
and ( n17219 , n17137 , n17218 );
or ( n17220 , n17136 , n17219 );
xor ( n17221 , n17133 , n17220 );
and ( n17222 , n817 , n6662 );
xor ( n17223 , n17221 , n17222 );
xor ( n17224 , n17137 , n17218 );
and ( n17225 , n818 , n6662 );
and ( n17226 , n17224 , n17225 );
xor ( n17227 , n17224 , n17225 );
xor ( n17228 , n17141 , n17216 );
and ( n17229 , n819 , n6662 );
and ( n17230 , n17228 , n17229 );
xor ( n17231 , n17228 , n17229 );
xor ( n17232 , n17145 , n17214 );
and ( n17233 , n820 , n6662 );
and ( n17234 , n17232 , n17233 );
xor ( n17235 , n17232 , n17233 );
xor ( n17236 , n17149 , n17212 );
and ( n17237 , n821 , n6662 );
and ( n17238 , n17236 , n17237 );
xor ( n17239 , n17236 , n17237 );
xor ( n17240 , n17153 , n17210 );
and ( n17241 , n822 , n6662 );
and ( n17242 , n17240 , n17241 );
xor ( n17243 , n17240 , n17241 );
xor ( n17244 , n17157 , n17208 );
and ( n17245 , n823 , n6662 );
and ( n17246 , n17244 , n17245 );
xor ( n17247 , n17244 , n17245 );
xor ( n17248 , n17161 , n17206 );
and ( n17249 , n824 , n6662 );
and ( n17250 , n17248 , n17249 );
xor ( n17251 , n17248 , n17249 );
xor ( n17252 , n17165 , n17204 );
and ( n17253 , n825 , n6662 );
and ( n17254 , n17252 , n17253 );
xor ( n17255 , n17252 , n17253 );
xor ( n17256 , n17169 , n17202 );
and ( n17257 , n826 , n6662 );
and ( n17258 , n17256 , n17257 );
xor ( n17259 , n17256 , n17257 );
xor ( n17260 , n17173 , n17200 );
and ( n17261 , n827 , n6662 );
and ( n17262 , n17260 , n17261 );
xor ( n17263 , n17260 , n17261 );
xor ( n17264 , n17177 , n17198 );
and ( n17265 , n828 , n6662 );
and ( n17266 , n17264 , n17265 );
xor ( n17267 , n17264 , n17265 );
xor ( n17268 , n17181 , n17196 );
and ( n17269 , n829 , n6662 );
and ( n17270 , n17268 , n17269 );
xor ( n17271 , n17268 , n17269 );
xor ( n17272 , n17185 , n17194 );
and ( n17273 , n830 , n6662 );
and ( n17274 , n17272 , n17273 );
xor ( n17275 , n17272 , n17273 );
xor ( n17276 , n17189 , n17192 );
and ( n17277 , n831 , n6662 );
and ( n17278 , n17276 , n17277 );
and ( n17279 , n17275 , n17278 );
or ( n17280 , n17274 , n17279 );
and ( n17281 , n17271 , n17280 );
or ( n17282 , n17270 , n17281 );
and ( n17283 , n17267 , n17282 );
or ( n17284 , n17266 , n17283 );
and ( n17285 , n17263 , n17284 );
or ( n17286 , n17262 , n17285 );
and ( n17287 , n17259 , n17286 );
or ( n17288 , n17258 , n17287 );
and ( n17289 , n17255 , n17288 );
or ( n17290 , n17254 , n17289 );
and ( n17291 , n17251 , n17290 );
or ( n17292 , n17250 , n17291 );
and ( n17293 , n17247 , n17292 );
or ( n17294 , n17246 , n17293 );
and ( n17295 , n17243 , n17294 );
or ( n17296 , n17242 , n17295 );
and ( n17297 , n17239 , n17296 );
or ( n17298 , n17238 , n17297 );
and ( n17299 , n17235 , n17298 );
or ( n17300 , n17234 , n17299 );
and ( n17301 , n17231 , n17300 );
or ( n17302 , n17230 , n17301 );
and ( n17303 , n17227 , n17302 );
or ( n17304 , n17226 , n17303 );
xor ( n17305 , n17223 , n17304 );
and ( n17306 , n818 , n6659 );
xor ( n17307 , n17305 , n17306 );
xor ( n17308 , n17227 , n17302 );
and ( n17309 , n819 , n6659 );
and ( n17310 , n17308 , n17309 );
xor ( n17311 , n17308 , n17309 );
xor ( n17312 , n17231 , n17300 );
and ( n17313 , n820 , n6659 );
and ( n17314 , n17312 , n17313 );
xor ( n17315 , n17312 , n17313 );
xor ( n17316 , n17235 , n17298 );
and ( n17317 , n821 , n6659 );
and ( n17318 , n17316 , n17317 );
xor ( n17319 , n17316 , n17317 );
xor ( n17320 , n17239 , n17296 );
and ( n17321 , n822 , n6659 );
and ( n17322 , n17320 , n17321 );
xor ( n17323 , n17320 , n17321 );
xor ( n17324 , n17243 , n17294 );
and ( n17325 , n823 , n6659 );
and ( n17326 , n17324 , n17325 );
xor ( n17327 , n17324 , n17325 );
xor ( n17328 , n17247 , n17292 );
and ( n17329 , n824 , n6659 );
and ( n17330 , n17328 , n17329 );
xor ( n17331 , n17328 , n17329 );
xor ( n17332 , n17251 , n17290 );
and ( n17333 , n825 , n6659 );
and ( n17334 , n17332 , n17333 );
xor ( n17335 , n17332 , n17333 );
xor ( n17336 , n17255 , n17288 );
and ( n17337 , n826 , n6659 );
and ( n17338 , n17336 , n17337 );
xor ( n17339 , n17336 , n17337 );
xor ( n17340 , n17259 , n17286 );
and ( n17341 , n827 , n6659 );
and ( n17342 , n17340 , n17341 );
xor ( n17343 , n17340 , n17341 );
xor ( n17344 , n17263 , n17284 );
and ( n17345 , n828 , n6659 );
and ( n17346 , n17344 , n17345 );
xor ( n17347 , n17344 , n17345 );
xor ( n17348 , n17267 , n17282 );
and ( n17349 , n829 , n6659 );
and ( n17350 , n17348 , n17349 );
xor ( n17351 , n17348 , n17349 );
xor ( n17352 , n17271 , n17280 );
and ( n17353 , n830 , n6659 );
and ( n17354 , n17352 , n17353 );
xor ( n17355 , n17352 , n17353 );
xor ( n17356 , n17275 , n17278 );
and ( n17357 , n831 , n6659 );
and ( n17358 , n17356 , n17357 );
and ( n17359 , n17355 , n17358 );
or ( n17360 , n17354 , n17359 );
and ( n17361 , n17351 , n17360 );
or ( n17362 , n17350 , n17361 );
and ( n17363 , n17347 , n17362 );
or ( n17364 , n17346 , n17363 );
and ( n17365 , n17343 , n17364 );
or ( n17366 , n17342 , n17365 );
and ( n17367 , n17339 , n17366 );
or ( n17368 , n17338 , n17367 );
and ( n17369 , n17335 , n17368 );
or ( n17370 , n17334 , n17369 );
and ( n17371 , n17331 , n17370 );
or ( n17372 , n17330 , n17371 );
and ( n17373 , n17327 , n17372 );
or ( n17374 , n17326 , n17373 );
and ( n17375 , n17323 , n17374 );
or ( n17376 , n17322 , n17375 );
and ( n17377 , n17319 , n17376 );
or ( n17378 , n17318 , n17377 );
and ( n17379 , n17315 , n17378 );
or ( n17380 , n17314 , n17379 );
and ( n17381 , n17311 , n17380 );
or ( n17382 , n17310 , n17381 );
xor ( n17383 , n17307 , n17382 );
and ( n17384 , n819 , n6656 );
xor ( n17385 , n17383 , n17384 );
xor ( n17386 , n17311 , n17380 );
and ( n17387 , n820 , n6656 );
and ( n17388 , n17386 , n17387 );
xor ( n17389 , n17386 , n17387 );
xor ( n17390 , n17315 , n17378 );
and ( n17391 , n821 , n6656 );
and ( n17392 , n17390 , n17391 );
xor ( n17393 , n17390 , n17391 );
xor ( n17394 , n17319 , n17376 );
and ( n17395 , n822 , n6656 );
and ( n17396 , n17394 , n17395 );
xor ( n17397 , n17394 , n17395 );
xor ( n17398 , n17323 , n17374 );
and ( n17399 , n823 , n6656 );
and ( n17400 , n17398 , n17399 );
xor ( n17401 , n17398 , n17399 );
xor ( n17402 , n17327 , n17372 );
and ( n17403 , n824 , n6656 );
and ( n17404 , n17402 , n17403 );
xor ( n17405 , n17402 , n17403 );
xor ( n17406 , n17331 , n17370 );
and ( n17407 , n825 , n6656 );
and ( n17408 , n17406 , n17407 );
xor ( n17409 , n17406 , n17407 );
xor ( n17410 , n17335 , n17368 );
and ( n17411 , n826 , n6656 );
and ( n17412 , n17410 , n17411 );
xor ( n17413 , n17410 , n17411 );
xor ( n17414 , n17339 , n17366 );
and ( n17415 , n827 , n6656 );
and ( n17416 , n17414 , n17415 );
xor ( n17417 , n17414 , n17415 );
xor ( n17418 , n17343 , n17364 );
and ( n17419 , n828 , n6656 );
and ( n17420 , n17418 , n17419 );
xor ( n17421 , n17418 , n17419 );
xor ( n17422 , n17347 , n17362 );
and ( n17423 , n829 , n6656 );
and ( n17424 , n17422 , n17423 );
xor ( n17425 , n17422 , n17423 );
xor ( n17426 , n17351 , n17360 );
and ( n17427 , n830 , n6656 );
and ( n17428 , n17426 , n17427 );
xor ( n17429 , n17426 , n17427 );
xor ( n17430 , n17355 , n17358 );
and ( n17431 , n831 , n6656 );
and ( n17432 , n17430 , n17431 );
and ( n17433 , n17429 , n17432 );
or ( n17434 , n17428 , n17433 );
and ( n17435 , n17425 , n17434 );
or ( n17436 , n17424 , n17435 );
and ( n17437 , n17421 , n17436 );
or ( n17438 , n17420 , n17437 );
and ( n17439 , n17417 , n17438 );
or ( n17440 , n17416 , n17439 );
and ( n17441 , n17413 , n17440 );
or ( n17442 , n17412 , n17441 );
and ( n17443 , n17409 , n17442 );
or ( n17444 , n17408 , n17443 );
and ( n17445 , n17405 , n17444 );
or ( n17446 , n17404 , n17445 );
and ( n17447 , n17401 , n17446 );
or ( n17448 , n17400 , n17447 );
and ( n17449 , n17397 , n17448 );
or ( n17450 , n17396 , n17449 );
and ( n17451 , n17393 , n17450 );
or ( n17452 , n17392 , n17451 );
and ( n17453 , n17389 , n17452 );
or ( n17454 , n17388 , n17453 );
xor ( n17455 , n17385 , n17454 );
and ( n17456 , n820 , n6653 );
xor ( n17457 , n17455 , n17456 );
xor ( n17458 , n17389 , n17452 );
and ( n17459 , n821 , n6653 );
and ( n17460 , n17458 , n17459 );
xor ( n17461 , n17458 , n17459 );
xor ( n17462 , n17393 , n17450 );
and ( n17463 , n822 , n6653 );
and ( n17464 , n17462 , n17463 );
xor ( n17465 , n17462 , n17463 );
xor ( n17466 , n17397 , n17448 );
and ( n17467 , n823 , n6653 );
and ( n17468 , n17466 , n17467 );
xor ( n17469 , n17466 , n17467 );
xor ( n17470 , n17401 , n17446 );
and ( n17471 , n824 , n6653 );
and ( n17472 , n17470 , n17471 );
xor ( n17473 , n17470 , n17471 );
xor ( n17474 , n17405 , n17444 );
and ( n17475 , n825 , n6653 );
and ( n17476 , n17474 , n17475 );
xor ( n17477 , n17474 , n17475 );
xor ( n17478 , n17409 , n17442 );
and ( n17479 , n826 , n6653 );
and ( n17480 , n17478 , n17479 );
xor ( n17481 , n17478 , n17479 );
xor ( n17482 , n17413 , n17440 );
and ( n17483 , n827 , n6653 );
and ( n17484 , n17482 , n17483 );
xor ( n17485 , n17482 , n17483 );
xor ( n17486 , n17417 , n17438 );
and ( n17487 , n828 , n6653 );
and ( n17488 , n17486 , n17487 );
xor ( n17489 , n17486 , n17487 );
xor ( n17490 , n17421 , n17436 );
and ( n17491 , n829 , n6653 );
and ( n17492 , n17490 , n17491 );
xor ( n17493 , n17490 , n17491 );
xor ( n17494 , n17425 , n17434 );
and ( n17495 , n830 , n6653 );
and ( n17496 , n17494 , n17495 );
xor ( n17497 , n17494 , n17495 );
xor ( n17498 , n17429 , n17432 );
and ( n17499 , n831 , n6653 );
and ( n17500 , n17498 , n17499 );
and ( n17501 , n17497 , n17500 );
or ( n17502 , n17496 , n17501 );
and ( n17503 , n17493 , n17502 );
or ( n17504 , n17492 , n17503 );
and ( n17505 , n17489 , n17504 );
or ( n17506 , n17488 , n17505 );
and ( n17507 , n17485 , n17506 );
or ( n17508 , n17484 , n17507 );
and ( n17509 , n17481 , n17508 );
or ( n17510 , n17480 , n17509 );
and ( n17511 , n17477 , n17510 );
or ( n17512 , n17476 , n17511 );
and ( n17513 , n17473 , n17512 );
or ( n17514 , n17472 , n17513 );
and ( n17515 , n17469 , n17514 );
or ( n17516 , n17468 , n17515 );
and ( n17517 , n17465 , n17516 );
or ( n17518 , n17464 , n17517 );
and ( n17519 , n17461 , n17518 );
or ( n17520 , n17460 , n17519 );
xor ( n17521 , n17457 , n17520 );
and ( n17522 , n821 , n6650 );
xor ( n17523 , n17521 , n17522 );
xor ( n17524 , n17461 , n17518 );
and ( n17525 , n822 , n6650 );
and ( n17526 , n17524 , n17525 );
xor ( n17527 , n17524 , n17525 );
xor ( n17528 , n17465 , n17516 );
and ( n17529 , n823 , n6650 );
and ( n17530 , n17528 , n17529 );
xor ( n17531 , n17528 , n17529 );
xor ( n17532 , n17469 , n17514 );
and ( n17533 , n824 , n6650 );
and ( n17534 , n17532 , n17533 );
xor ( n17535 , n17532 , n17533 );
xor ( n17536 , n17473 , n17512 );
and ( n17537 , n825 , n6650 );
and ( n17538 , n17536 , n17537 );
xor ( n17539 , n17536 , n17537 );
xor ( n17540 , n17477 , n17510 );
and ( n17541 , n826 , n6650 );
and ( n17542 , n17540 , n17541 );
xor ( n17543 , n17540 , n17541 );
xor ( n17544 , n17481 , n17508 );
and ( n17545 , n827 , n6650 );
and ( n17546 , n17544 , n17545 );
xor ( n17547 , n17544 , n17545 );
xor ( n17548 , n17485 , n17506 );
and ( n17549 , n828 , n6650 );
and ( n17550 , n17548 , n17549 );
xor ( n17551 , n17548 , n17549 );
xor ( n17552 , n17489 , n17504 );
and ( n17553 , n829 , n6650 );
and ( n17554 , n17552 , n17553 );
xor ( n17555 , n17552 , n17553 );
xor ( n17556 , n17493 , n17502 );
and ( n17557 , n830 , n6650 );
and ( n17558 , n17556 , n17557 );
xor ( n17559 , n17556 , n17557 );
xor ( n17560 , n17497 , n17500 );
and ( n17561 , n831 , n6650 );
and ( n17562 , n17560 , n17561 );
and ( n17563 , n17559 , n17562 );
or ( n17564 , n17558 , n17563 );
and ( n17565 , n17555 , n17564 );
or ( n17566 , n17554 , n17565 );
and ( n17567 , n17551 , n17566 );
or ( n17568 , n17550 , n17567 );
and ( n17569 , n17547 , n17568 );
or ( n17570 , n17546 , n17569 );
and ( n17571 , n17543 , n17570 );
or ( n17572 , n17542 , n17571 );
and ( n17573 , n17539 , n17572 );
or ( n17574 , n17538 , n17573 );
and ( n17575 , n17535 , n17574 );
or ( n17576 , n17534 , n17575 );
and ( n17577 , n17531 , n17576 );
or ( n17578 , n17530 , n17577 );
and ( n17579 , n17527 , n17578 );
or ( n17580 , n17526 , n17579 );
xor ( n17581 , n17523 , n17580 );
and ( n17582 , n822 , n6647 );
xor ( n17583 , n17581 , n17582 );
xor ( n17584 , n17527 , n17578 );
and ( n17585 , n823 , n6647 );
and ( n17586 , n17584 , n17585 );
xor ( n17587 , n17584 , n17585 );
xor ( n17588 , n17531 , n17576 );
and ( n17589 , n824 , n6647 );
and ( n17590 , n17588 , n17589 );
xor ( n17591 , n17588 , n17589 );
xor ( n17592 , n17535 , n17574 );
and ( n17593 , n825 , n6647 );
and ( n17594 , n17592 , n17593 );
xor ( n17595 , n17592 , n17593 );
xor ( n17596 , n17539 , n17572 );
and ( n17597 , n826 , n6647 );
and ( n17598 , n17596 , n17597 );
xor ( n17599 , n17596 , n17597 );
xor ( n17600 , n17543 , n17570 );
and ( n17601 , n827 , n6647 );
and ( n17602 , n17600 , n17601 );
xor ( n17603 , n17600 , n17601 );
xor ( n17604 , n17547 , n17568 );
and ( n17605 , n828 , n6647 );
and ( n17606 , n17604 , n17605 );
xor ( n17607 , n17604 , n17605 );
xor ( n17608 , n17551 , n17566 );
and ( n17609 , n829 , n6647 );
and ( n17610 , n17608 , n17609 );
xor ( n17611 , n17608 , n17609 );
xor ( n17612 , n17555 , n17564 );
and ( n17613 , n830 , n6647 );
and ( n17614 , n17612 , n17613 );
xor ( n17615 , n17612 , n17613 );
xor ( n17616 , n17559 , n17562 );
and ( n17617 , n831 , n6647 );
and ( n17618 , n17616 , n17617 );
and ( n17619 , n17615 , n17618 );
or ( n17620 , n17614 , n17619 );
and ( n17621 , n17611 , n17620 );
or ( n17622 , n17610 , n17621 );
and ( n17623 , n17607 , n17622 );
or ( n17624 , n17606 , n17623 );
and ( n17625 , n17603 , n17624 );
or ( n17626 , n17602 , n17625 );
and ( n17627 , n17599 , n17626 );
or ( n17628 , n17598 , n17627 );
and ( n17629 , n17595 , n17628 );
or ( n17630 , n17594 , n17629 );
and ( n17631 , n17591 , n17630 );
or ( n17632 , n17590 , n17631 );
and ( n17633 , n17587 , n17632 );
or ( n17634 , n17586 , n17633 );
xor ( n17635 , n17583 , n17634 );
and ( n17636 , n823 , n6644 );
xor ( n17637 , n17635 , n17636 );
xor ( n17638 , n17587 , n17632 );
and ( n17639 , n824 , n6644 );
and ( n17640 , n17638 , n17639 );
xor ( n17641 , n17638 , n17639 );
xor ( n17642 , n17591 , n17630 );
and ( n17643 , n825 , n6644 );
and ( n17644 , n17642 , n17643 );
xor ( n17645 , n17642 , n17643 );
xor ( n17646 , n17595 , n17628 );
and ( n17647 , n826 , n6644 );
and ( n17648 , n17646 , n17647 );
xor ( n17649 , n17646 , n17647 );
xor ( n17650 , n17599 , n17626 );
and ( n17651 , n827 , n6644 );
and ( n17652 , n17650 , n17651 );
xor ( n17653 , n17650 , n17651 );
xor ( n17654 , n17603 , n17624 );
and ( n17655 , n828 , n6644 );
and ( n17656 , n17654 , n17655 );
xor ( n17657 , n17654 , n17655 );
xor ( n17658 , n17607 , n17622 );
and ( n17659 , n829 , n6644 );
and ( n17660 , n17658 , n17659 );
xor ( n17661 , n17658 , n17659 );
xor ( n17662 , n17611 , n17620 );
and ( n17663 , n830 , n6644 );
and ( n17664 , n17662 , n17663 );
xor ( n17665 , n17662 , n17663 );
xor ( n17666 , n17615 , n17618 );
and ( n17667 , n831 , n6644 );
and ( n17668 , n17666 , n17667 );
and ( n17669 , n17665 , n17668 );
or ( n17670 , n17664 , n17669 );
and ( n17671 , n17661 , n17670 );
or ( n17672 , n17660 , n17671 );
and ( n17673 , n17657 , n17672 );
or ( n17674 , n17656 , n17673 );
and ( n17675 , n17653 , n17674 );
or ( n17676 , n17652 , n17675 );
and ( n17677 , n17649 , n17676 );
or ( n17678 , n17648 , n17677 );
and ( n17679 , n17645 , n17678 );
or ( n17680 , n17644 , n17679 );
and ( n17681 , n17641 , n17680 );
or ( n17682 , n17640 , n17681 );
xor ( n17683 , n17637 , n17682 );
and ( n17684 , n824 , n6641 );
xor ( n17685 , n17683 , n17684 );
xor ( n17686 , n17641 , n17680 );
and ( n17687 , n825 , n6641 );
and ( n17688 , n17686 , n17687 );
xor ( n17689 , n17686 , n17687 );
xor ( n17690 , n17645 , n17678 );
and ( n17691 , n826 , n6641 );
and ( n17692 , n17690 , n17691 );
xor ( n17693 , n17690 , n17691 );
xor ( n17694 , n17649 , n17676 );
and ( n17695 , n827 , n6641 );
and ( n17696 , n17694 , n17695 );
xor ( n17697 , n17694 , n17695 );
xor ( n17698 , n17653 , n17674 );
and ( n17699 , n828 , n6641 );
and ( n17700 , n17698 , n17699 );
xor ( n17701 , n17698 , n17699 );
xor ( n17702 , n17657 , n17672 );
and ( n17703 , n829 , n6641 );
and ( n17704 , n17702 , n17703 );
xor ( n17705 , n17702 , n17703 );
xor ( n17706 , n17661 , n17670 );
and ( n17707 , n830 , n6641 );
and ( n17708 , n17706 , n17707 );
xor ( n17709 , n17706 , n17707 );
xor ( n17710 , n17665 , n17668 );
and ( n17711 , n831 , n6641 );
and ( n17712 , n17710 , n17711 );
and ( n17713 , n17709 , n17712 );
or ( n17714 , n17708 , n17713 );
and ( n17715 , n17705 , n17714 );
or ( n17716 , n17704 , n17715 );
and ( n17717 , n17701 , n17716 );
or ( n17718 , n17700 , n17717 );
and ( n17719 , n17697 , n17718 );
or ( n17720 , n17696 , n17719 );
and ( n17721 , n17693 , n17720 );
or ( n17722 , n17692 , n17721 );
and ( n17723 , n17689 , n17722 );
or ( n17724 , n17688 , n17723 );
xor ( n17725 , n17685 , n17724 );
and ( n17726 , n825 , n6638 );
xor ( n17727 , n17725 , n17726 );
xor ( n17728 , n17689 , n17722 );
and ( n17729 , n826 , n6638 );
and ( n17730 , n17728 , n17729 );
xor ( n17731 , n17728 , n17729 );
xor ( n17732 , n17693 , n17720 );
and ( n17733 , n827 , n6638 );
and ( n17734 , n17732 , n17733 );
xor ( n17735 , n17732 , n17733 );
xor ( n17736 , n17697 , n17718 );
and ( n17737 , n828 , n6638 );
and ( n17738 , n17736 , n17737 );
xor ( n17739 , n17736 , n17737 );
xor ( n17740 , n17701 , n17716 );
and ( n17741 , n829 , n6638 );
and ( n17742 , n17740 , n17741 );
xor ( n17743 , n17740 , n17741 );
xor ( n17744 , n17705 , n17714 );
and ( n17745 , n830 , n6638 );
and ( n17746 , n17744 , n17745 );
xor ( n17747 , n17744 , n17745 );
xor ( n17748 , n17709 , n17712 );
and ( n17749 , n831 , n6638 );
and ( n17750 , n17748 , n17749 );
and ( n17751 , n17747 , n17750 );
or ( n17752 , n17746 , n17751 );
and ( n17753 , n17743 , n17752 );
or ( n17754 , n17742 , n17753 );
and ( n17755 , n17739 , n17754 );
or ( n17756 , n17738 , n17755 );
and ( n17757 , n17735 , n17756 );
or ( n17758 , n17734 , n17757 );
and ( n17759 , n17731 , n17758 );
or ( n17760 , n17730 , n17759 );
xor ( n17761 , n17727 , n17760 );
and ( n17762 , n826 , n6635 );
xor ( n17763 , n17761 , n17762 );
xor ( n17764 , n17731 , n17758 );
and ( n17765 , n827 , n6635 );
and ( n17766 , n17764 , n17765 );
xor ( n17767 , n17764 , n17765 );
xor ( n17768 , n17735 , n17756 );
and ( n17769 , n828 , n6635 );
and ( n17770 , n17768 , n17769 );
xor ( n17771 , n17768 , n17769 );
xor ( n17772 , n17739 , n17754 );
and ( n17773 , n829 , n6635 );
and ( n17774 , n17772 , n17773 );
xor ( n17775 , n17772 , n17773 );
xor ( n17776 , n17743 , n17752 );
and ( n17777 , n830 , n6635 );
and ( n17778 , n17776 , n17777 );
xor ( n17779 , n17776 , n17777 );
xor ( n17780 , n17747 , n17750 );
and ( n17781 , n831 , n6635 );
and ( n17782 , n17780 , n17781 );
and ( n17783 , n17779 , n17782 );
or ( n17784 , n17778 , n17783 );
and ( n17785 , n17775 , n17784 );
or ( n17786 , n17774 , n17785 );
and ( n17787 , n17771 , n17786 );
or ( n17788 , n17770 , n17787 );
and ( n17789 , n17767 , n17788 );
or ( n17790 , n17766 , n17789 );
xor ( n17791 , n17763 , n17790 );
and ( n17792 , n827 , n6632 );
xor ( n17793 , n17791 , n17792 );
xor ( n17794 , n17767 , n17788 );
and ( n17795 , n828 , n6632 );
and ( n17796 , n17794 , n17795 );
xor ( n17797 , n17794 , n17795 );
xor ( n17798 , n17771 , n17786 );
and ( n17799 , n829 , n6632 );
and ( n17800 , n17798 , n17799 );
xor ( n17801 , n17798 , n17799 );
xor ( n17802 , n17775 , n17784 );
and ( n17803 , n830 , n6632 );
and ( n17804 , n17802 , n17803 );
xor ( n17805 , n17802 , n17803 );
xor ( n17806 , n17779 , n17782 );
and ( n17807 , n831 , n6632 );
and ( n17808 , n17806 , n17807 );
and ( n17809 , n17805 , n17808 );
or ( n17810 , n17804 , n17809 );
and ( n17811 , n17801 , n17810 );
or ( n17812 , n17800 , n17811 );
and ( n17813 , n17797 , n17812 );
or ( n17814 , n17796 , n17813 );
xor ( n17815 , n17793 , n17814 );
and ( n17816 , n828 , n6629 );
xor ( n17817 , n17815 , n17816 );
xor ( n17818 , n17797 , n17812 );
and ( n17819 , n829 , n6629 );
and ( n17820 , n17818 , n17819 );
xor ( n17821 , n17818 , n17819 );
xor ( n17822 , n17801 , n17810 );
and ( n17823 , n830 , n6629 );
and ( n17824 , n17822 , n17823 );
xor ( n17825 , n17822 , n17823 );
xor ( n17826 , n17805 , n17808 );
and ( n17827 , n831 , n6629 );
and ( n17828 , n17826 , n17827 );
and ( n17829 , n17825 , n17828 );
or ( n17830 , n17824 , n17829 );
and ( n17831 , n17821 , n17830 );
or ( n17832 , n17820 , n17831 );
xor ( n17833 , n17817 , n17832 );
and ( n17834 , n829 , n6626 );
xor ( n17835 , n17833 , n17834 );
xor ( n17836 , n17821 , n17830 );
and ( n17837 , n830 , n6626 );
and ( n17838 , n17836 , n17837 );
xor ( n17839 , n17836 , n17837 );
xor ( n17840 , n17825 , n17828 );
and ( n17841 , n831 , n6626 );
and ( n17842 , n17840 , n17841 );
and ( n17843 , n17839 , n17842 );
or ( n17844 , n17838 , n17843 );
xor ( n17845 , n17835 , n17844 );
and ( n17846 , n830 , n6623 );
xor ( n17847 , n17845 , n17846 );
xor ( n17848 , n17839 , n17842 );
and ( n17849 , n831 , n6623 );
and ( n17850 , n17848 , n17849 );
xor ( n17851 , n17847 , n17850 );
and ( n17852 , n831 , n6620 );
xor ( n17853 , n17851 , n17852 );
buf ( n17854 , n17853 );
xor ( n17855 , n17848 , n17849 );
buf ( n17856 , n17855 );
xor ( n17857 , n17840 , n17841 );
buf ( n17858 , n17857 );
xor ( n17859 , n17826 , n17827 );
buf ( n17860 , n17859 );
xor ( n17861 , n17806 , n17807 );
buf ( n17862 , n17861 );
xor ( n17863 , n17780 , n17781 );
buf ( n17864 , n17863 );
xor ( n17865 , n17748 , n17749 );
buf ( n17866 , n17865 );
xor ( n17867 , n17710 , n17711 );
buf ( n17868 , n17867 );
xor ( n17869 , n17666 , n17667 );
buf ( n17870 , n17869 );
xor ( n17871 , n17616 , n17617 );
buf ( n17872 , n17871 );
xor ( n17873 , n17560 , n17561 );
buf ( n17874 , n17873 );
xor ( n17875 , n17498 , n17499 );
buf ( n17876 , n17875 );
xor ( n17877 , n17430 , n17431 );
buf ( n17878 , n17877 );
xor ( n17879 , n17356 , n17357 );
buf ( n17880 , n17879 );
xor ( n17881 , n17276 , n17277 );
buf ( n17882 , n17881 );
xor ( n17883 , n17190 , n17191 );
buf ( n17884 , n17883 );
xor ( n17885 , n17099 , n17100 );
buf ( n17886 , n17885 );
xor ( n17887 , n17007 , n17008 );
buf ( n17888 , n17887 );
xor ( n17889 , n16915 , n16916 );
buf ( n17890 , n17889 );
xor ( n17891 , n16823 , n16824 );
buf ( n17892 , n17891 );
xor ( n17893 , n16731 , n16732 );
buf ( n17894 , n17893 );
xor ( n17895 , n16639 , n16640 );
buf ( n17896 , n17895 );
xor ( n17897 , n16547 , n16548 );
buf ( n17898 , n17897 );
xor ( n17899 , n16455 , n16456 );
buf ( n17900 , n17899 );
xor ( n17901 , n16363 , n16364 );
buf ( n17902 , n17901 );
xor ( n17903 , n16271 , n16272 );
buf ( n17904 , n17903 );
xor ( n17905 , n16179 , n16180 );
buf ( n17906 , n17905 );
xor ( n17907 , n16087 , n16088 );
buf ( n17908 , n17907 );
xor ( n17909 , n15995 , n15996 );
buf ( n17910 , n17909 );
xor ( n17911 , n15903 , n15904 );
buf ( n17912 , n17911 );
xor ( n17913 , n15811 , n15812 );
buf ( n17914 , n17913 );
xor ( n17915 , n15719 , n15720 );
buf ( n17916 , n17915 );
xor ( n17917 , n15627 , n15628 );
buf ( n17918 , n17917 );
xor ( n17919 , n15535 , n15536 );
buf ( n17920 , n17919 );
xor ( n17921 , n15443 , n15444 );
buf ( n17922 , n17921 );
xor ( n17923 , n15351 , n15352 );
buf ( n17924 , n17923 );
xor ( n17925 , n15259 , n15260 );
buf ( n17926 , n17925 );
xor ( n17927 , n15167 , n15168 );
buf ( n17928 , n17927 );
xor ( n17929 , n15075 , n15076 );
buf ( n17930 , n17929 );
xor ( n17931 , n14983 , n14984 );
buf ( n17932 , n17931 );
xor ( n17933 , n14891 , n14892 );
buf ( n17934 , n17933 );
xor ( n17935 , n14799 , n14800 );
buf ( n17936 , n17935 );
xor ( n17937 , n14707 , n14708 );
buf ( n17938 , n17937 );
xor ( n17939 , n14615 , n14616 );
buf ( n17940 , n17939 );
xor ( n17941 , n14523 , n14524 );
buf ( n17942 , n17941 );
xor ( n17943 , n14431 , n14432 );
buf ( n17944 , n17943 );
xor ( n17945 , n14339 , n14340 );
buf ( n17946 , n17945 );
xor ( n17947 , n14247 , n14248 );
buf ( n17948 , n17947 );
xor ( n17949 , n14155 , n14156 );
buf ( n17950 , n17949 );
xor ( n17951 , n14063 , n14064 );
buf ( n17952 , n17951 );
xor ( n17953 , n13971 , n13972 );
buf ( n17954 , n17953 );
xor ( n17955 , n13879 , n13880 );
buf ( n17956 , n17955 );
xor ( n17957 , n13787 , n13788 );
buf ( n17958 , n17957 );
xor ( n17959 , n13695 , n13696 );
buf ( n17960 , n17959 );
xor ( n17961 , n13603 , n13604 );
buf ( n17962 , n17961 );
xor ( n17963 , n13511 , n13512 );
buf ( n17964 , n17963 );
xor ( n17965 , n13419 , n13420 );
buf ( n17966 , n17965 );
xor ( n17967 , n13327 , n13328 );
buf ( n17968 , n17967 );
xor ( n17969 , n13235 , n13236 );
buf ( n17970 , n17969 );
xor ( n17971 , n13143 , n13144 );
buf ( n17972 , n17971 );
xor ( n17973 , n13051 , n13052 );
buf ( n17974 , n17973 );
xor ( n17975 , n12959 , n12960 );
buf ( n17976 , n17975 );
xor ( n17977 , n12867 , n12868 );
buf ( n17978 , n17977 );
xor ( n17979 , n12775 , n12776 );
buf ( n17980 , n17979 );
xor ( n17981 , n12683 , n12684 );
buf ( n17982 , n17981 );
xor ( n17983 , n12591 , n12592 );
buf ( n17984 , n17983 );
xor ( n17985 , n12499 , n12500 );
buf ( n17986 , n17985 );
xor ( n17987 , n12407 , n12408 );
buf ( n17988 , n17987 );
xor ( n17989 , n12315 , n12316 );
buf ( n17990 , n17989 );
xor ( n17991 , n12223 , n12224 );
buf ( n17992 , n17991 );
xor ( n17993 , n12131 , n12132 );
buf ( n17994 , n17993 );
xor ( n17995 , n12039 , n12040 );
buf ( n17996 , n17995 );
xor ( n17997 , n11947 , n11948 );
buf ( n17998 , n17997 );
xor ( n17999 , n11855 , n11856 );
buf ( n18000 , n17999 );
xor ( n18001 , n11763 , n11764 );
buf ( n18002 , n18001 );
xor ( n18003 , n11671 , n11672 );
buf ( n18004 , n18003 );
xor ( n18005 , n11579 , n11580 );
buf ( n18006 , n18005 );
xor ( n18007 , n11487 , n11488 );
buf ( n18008 , n18007 );
xor ( n18009 , n11395 , n11396 );
buf ( n18010 , n18009 );
xor ( n18011 , n11303 , n11304 );
buf ( n18012 , n18011 );
xor ( n18013 , n11211 , n11212 );
buf ( n18014 , n18013 );
xor ( n18015 , n11119 , n11120 );
buf ( n18016 , n18015 );
xor ( n18017 , n11027 , n11028 );
buf ( n18018 , n18017 );
xor ( n18019 , n10935 , n10936 );
buf ( n18020 , n18019 );
xor ( n18021 , n10843 , n10844 );
buf ( n18022 , n18021 );
xor ( n18023 , n10751 , n10752 );
buf ( n18024 , n18023 );
xor ( n18025 , n10659 , n10660 );
buf ( n18026 , n18025 );
xor ( n18027 , n10567 , n10568 );
buf ( n18028 , n18027 );
xor ( n18029 , n10475 , n10476 );
buf ( n18030 , n18029 );
xor ( n18031 , n10383 , n10384 );
buf ( n18032 , n18031 );
xor ( n18033 , n10291 , n10292 );
buf ( n18034 , n18033 );
xor ( n18035 , n10199 , n10200 );
buf ( n18036 , n18035 );
xor ( n18037 , n10107 , n10108 );
buf ( n18038 , n18037 );
xor ( n18039 , n10015 , n10016 );
buf ( n18040 , n18039 );
xor ( n18041 , n9923 , n9924 );
buf ( n18042 , n18041 );
xor ( n18043 , n9831 , n9832 );
buf ( n18044 , n18043 );
xor ( n18045 , n9739 , n9740 );
buf ( n18046 , n18045 );
xor ( n18047 , n9647 , n9648 );
buf ( n18048 , n18047 );
xor ( n18049 , n9555 , n9556 );
buf ( n18050 , n18049 );
xor ( n18051 , n9463 , n9464 );
buf ( n18052 , n18051 );
xor ( n18053 , n9371 , n9372 );
buf ( n18054 , n18053 );
xor ( n18055 , n9279 , n9280 );
buf ( n18056 , n18055 );
xor ( n18057 , n9187 , n9188 );
buf ( n18058 , n18057 );
xor ( n18059 , n9095 , n9096 );
buf ( n18060 , n18059 );
xor ( n18061 , n9003 , n9004 );
buf ( n18062 , n18061 );
xor ( n18063 , n8911 , n8912 );
buf ( n18064 , n18063 );
xor ( n18065 , n8819 , n8820 );
buf ( n18066 , n18065 );
xor ( n18067 , n8727 , n8728 );
buf ( n18068 , n18067 );
xor ( n18069 , n8635 , n8636 );
buf ( n18070 , n18069 );
xor ( n18071 , n8543 , n8544 );
buf ( n18072 , n18071 );
xor ( n18073 , n8451 , n8452 );
buf ( n18074 , n18073 );
xor ( n18075 , n8359 , n8360 );
buf ( n18076 , n18075 );
xor ( n18077 , n8267 , n8268 );
buf ( n18078 , n18077 );
xor ( n18079 , n8175 , n8176 );
buf ( n18080 , n18079 );
xor ( n18081 , n8083 , n8084 );
buf ( n18082 , n18081 );
xor ( n18083 , n7991 , n7992 );
buf ( n18084 , n18083 );
xor ( n18085 , n7899 , n7900 );
buf ( n18086 , n18085 );
xor ( n18087 , n7807 , n7808 );
buf ( n18088 , n18087 );
xor ( n18089 , n7715 , n7716 );
buf ( n18090 , n18089 );
xor ( n18091 , n7623 , n7624 );
buf ( n18092 , n18091 );
xor ( n18093 , n7531 , n7532 );
buf ( n18094 , n18093 );
xor ( n18095 , n7439 , n7440 );
buf ( n18096 , n18095 );
xor ( n18097 , n7347 , n7348 );
buf ( n18098 , n18097 );
xor ( n18099 , n7255 , n7256 );
buf ( n18100 , n18099 );
xor ( n18101 , n7163 , n7164 );
buf ( n18102 , n18101 );
xor ( n18103 , n7072 , n7073 );
buf ( n18104 , n18103 );
and ( n18105 , n831 , n7014 );
buf ( n18106 , n18105 );
buf ( n18107 , n576 );
buf ( n18108 , n577 );
buf ( n18109 , n578 );
buf ( n18110 , n579 );
buf ( n18111 , n580 );
buf ( n18112 , n581 );
buf ( n18113 , n582 );
buf ( n18114 , n583 );
buf ( n18115 , n584 );
buf ( n18116 , n585 );
buf ( n18117 , n586 );
buf ( n18118 , n587 );
buf ( n18119 , n588 );
buf ( n18120 , n589 );
buf ( n18121 , n590 );
buf ( n18122 , n591 );
buf ( n18123 , n4041 );
buf ( n18124 , n5783 );
not ( n18125 , n18124 );
and ( n18126 , n18123 , n18125 );
buf ( n18127 , n5788 );
buf ( n18128 , n5791 );
not ( n18129 , n18128 );
and ( n18130 , n18127 , n18129 );
buf ( n18131 , n5796 );
buf ( n18132 , n5799 );
not ( n18133 , n18132 );
and ( n18134 , n18131 , n18133 );
buf ( n18135 , n5804 );
buf ( n18136 , n5807 );
not ( n18137 , n18136 );
and ( n18138 , n18135 , n18137 );
buf ( n18139 , n5812 );
buf ( n18140 , n5815 );
not ( n18141 , n18140 );
and ( n18142 , n18139 , n18141 );
buf ( n18143 , n5820 );
buf ( n18144 , n5823 );
not ( n18145 , n18144 );
and ( n18146 , n18143 , n18145 );
buf ( n18147 , n5828 );
buf ( n18148 , n5831 );
not ( n18149 , n18148 );
and ( n18150 , n18147 , n18149 );
buf ( n18151 , n5836 );
buf ( n18152 , n5839 );
not ( n18153 , n18152 );
and ( n18154 , n18151 , n18153 );
buf ( n18155 , n5844 );
buf ( n18156 , n5847 );
not ( n18157 , n18156 );
and ( n18158 , n18155 , n18157 );
buf ( n18159 , n5852 );
buf ( n18160 , n5855 );
not ( n18161 , n18160 );
and ( n18162 , n18159 , n18161 );
buf ( n18163 , n5860 );
buf ( n18164 , n5863 );
not ( n18165 , n18164 );
and ( n18166 , n18163 , n18165 );
buf ( n18167 , n5868 );
buf ( n18168 , n5871 );
not ( n18169 , n18168 );
and ( n18170 , n18167 , n18169 );
buf ( n18171 , n5876 );
buf ( n18172 , n5879 );
not ( n18173 , n18172 );
and ( n18174 , n18171 , n18173 );
buf ( n18175 , n5884 );
buf ( n18176 , n5887 );
not ( n18177 , n18176 );
and ( n18178 , n18175 , n18177 );
buf ( n18179 , n5892 );
buf ( n18180 , n5895 );
not ( n18181 , n18180 );
and ( n18182 , n18179 , n18181 );
buf ( n18183 , n5900 );
buf ( n18184 , n5903 );
not ( n18185 , n18184 );
and ( n18186 , n18183 , n18185 );
buf ( n18187 , n5908 );
buf ( n18188 , n5911 );
not ( n18189 , n18188 );
and ( n18190 , n18187 , n18189 );
buf ( n18191 , n5916 );
buf ( n18192 , n5919 );
not ( n18193 , n18192 );
and ( n18194 , n18191 , n18193 );
buf ( n18195 , n5924 );
buf ( n18196 , n5927 );
not ( n18197 , n18196 );
and ( n18198 , n18195 , n18197 );
buf ( n18199 , n5932 );
buf ( n18200 , n5935 );
not ( n18201 , n18200 );
and ( n18202 , n18199 , n18201 );
buf ( n18203 , n5940 );
buf ( n18204 , n5943 );
not ( n18205 , n18204 );
and ( n18206 , n18203 , n18205 );
buf ( n18207 , n5948 );
buf ( n18208 , n5951 );
not ( n18209 , n18208 );
and ( n18210 , n18207 , n18209 );
buf ( n18211 , n5956 );
buf ( n18212 , n5959 );
not ( n18213 , n18212 );
and ( n18214 , n18211 , n18213 );
buf ( n18215 , n5964 );
buf ( n18216 , n5967 );
not ( n18217 , n18216 );
and ( n18218 , n18215 , n18217 );
buf ( n18219 , n5972 );
buf ( n18220 , n5975 );
not ( n18221 , n18220 );
and ( n18222 , n18219 , n18221 );
buf ( n18223 , n5980 );
buf ( n18224 , n5983 );
not ( n18225 , n18224 );
and ( n18226 , n18223 , n18225 );
buf ( n18227 , n5988 );
buf ( n18228 , n5991 );
not ( n18229 , n18228 );
and ( n18230 , n18227 , n18229 );
buf ( n18231 , n5996 );
buf ( n18232 , n5999 );
not ( n18233 , n18232 );
and ( n18234 , n18231 , n18233 );
buf ( n18235 , n6004 );
buf ( n18236 , n6007 );
not ( n18237 , n18236 );
and ( n18238 , n18235 , n18237 );
buf ( n18239 , n6012 );
buf ( n18240 , n6015 );
not ( n18241 , n18240 );
and ( n18242 , n18239 , n18241 );
buf ( n18243 , n6020 );
buf ( n18244 , n6023 );
not ( n18245 , n18244 );
and ( n18246 , n18243 , n18245 );
buf ( n18247 , n18245 );
buf ( n18248 , n18243 );
or ( n18249 , n18246 , n18247 , n18248 );
and ( n18250 , n18241 , n18249 );
and ( n18251 , n18239 , n18249 );
or ( n18252 , n18242 , n18250 , n18251 );
and ( n18253 , n18237 , n18252 );
and ( n18254 , n18235 , n18252 );
or ( n18255 , n18238 , n18253 , n18254 );
and ( n18256 , n18233 , n18255 );
and ( n18257 , n18231 , n18255 );
or ( n18258 , n18234 , n18256 , n18257 );
and ( n18259 , n18229 , n18258 );
and ( n18260 , n18227 , n18258 );
or ( n18261 , n18230 , n18259 , n18260 );
and ( n18262 , n18225 , n18261 );
and ( n18263 , n18223 , n18261 );
or ( n18264 , n18226 , n18262 , n18263 );
and ( n18265 , n18221 , n18264 );
and ( n18266 , n18219 , n18264 );
or ( n18267 , n18222 , n18265 , n18266 );
and ( n18268 , n18217 , n18267 );
and ( n18269 , n18215 , n18267 );
or ( n18270 , n18218 , n18268 , n18269 );
and ( n18271 , n18213 , n18270 );
and ( n18272 , n18211 , n18270 );
or ( n18273 , n18214 , n18271 , n18272 );
and ( n18274 , n18209 , n18273 );
and ( n18275 , n18207 , n18273 );
or ( n18276 , n18210 , n18274 , n18275 );
and ( n18277 , n18205 , n18276 );
and ( n18278 , n18203 , n18276 );
or ( n18279 , n18206 , n18277 , n18278 );
and ( n18280 , n18201 , n18279 );
and ( n18281 , n18199 , n18279 );
or ( n18282 , n18202 , n18280 , n18281 );
and ( n18283 , n18197 , n18282 );
and ( n18284 , n18195 , n18282 );
or ( n18285 , n18198 , n18283 , n18284 );
and ( n18286 , n18193 , n18285 );
and ( n18287 , n18191 , n18285 );
or ( n18288 , n18194 , n18286 , n18287 );
and ( n18289 , n18189 , n18288 );
and ( n18290 , n18187 , n18288 );
or ( n18291 , n18190 , n18289 , n18290 );
and ( n18292 , n18185 , n18291 );
and ( n18293 , n18183 , n18291 );
or ( n18294 , n18186 , n18292 , n18293 );
and ( n18295 , n18181 , n18294 );
and ( n18296 , n18179 , n18294 );
or ( n18297 , n18182 , n18295 , n18296 );
and ( n18298 , n18177 , n18297 );
and ( n18299 , n18175 , n18297 );
or ( n18300 , n18178 , n18298 , n18299 );
and ( n18301 , n18173 , n18300 );
and ( n18302 , n18171 , n18300 );
or ( n18303 , n18174 , n18301 , n18302 );
and ( n18304 , n18169 , n18303 );
and ( n18305 , n18167 , n18303 );
or ( n18306 , n18170 , n18304 , n18305 );
and ( n18307 , n18165 , n18306 );
and ( n18308 , n18163 , n18306 );
or ( n18309 , n18166 , n18307 , n18308 );
and ( n18310 , n18161 , n18309 );
and ( n18311 , n18159 , n18309 );
or ( n18312 , n18162 , n18310 , n18311 );
and ( n18313 , n18157 , n18312 );
and ( n18314 , n18155 , n18312 );
or ( n18315 , n18158 , n18313 , n18314 );
and ( n18316 , n18153 , n18315 );
and ( n18317 , n18151 , n18315 );
or ( n18318 , n18154 , n18316 , n18317 );
and ( n18319 , n18149 , n18318 );
and ( n18320 , n18147 , n18318 );
or ( n18321 , n18150 , n18319 , n18320 );
and ( n18322 , n18145 , n18321 );
and ( n18323 , n18143 , n18321 );
or ( n18324 , n18146 , n18322 , n18323 );
and ( n18325 , n18141 , n18324 );
and ( n18326 , n18139 , n18324 );
or ( n18327 , n18142 , n18325 , n18326 );
and ( n18328 , n18137 , n18327 );
and ( n18329 , n18135 , n18327 );
or ( n18330 , n18138 , n18328 , n18329 );
and ( n18331 , n18133 , n18330 );
and ( n18332 , n18131 , n18330 );
or ( n18333 , n18134 , n18331 , n18332 );
and ( n18334 , n18129 , n18333 );
and ( n18335 , n18127 , n18333 );
or ( n18336 , n18130 , n18334 , n18335 );
and ( n18337 , n18125 , n18336 );
and ( n18338 , n18123 , n18336 );
or ( n18339 , n18126 , n18337 , n18338 );
not ( n18340 , n18339 );
buf ( n18341 , n18340 );
buf ( n18342 , n18341 );
buf ( n18343 , n18340 );
buf ( n18344 , n18343 );
buf ( n18345 , n18340 );
buf ( n18346 , n18345 );
buf ( n18347 , n18340 );
buf ( n18348 , n18347 );
buf ( n18349 , n18340 );
buf ( n18350 , n18349 );
buf ( n18351 , n18340 );
buf ( n18352 , n18351 );
buf ( n18353 , n18340 );
buf ( n18354 , n18353 );
buf ( n18355 , n18340 );
buf ( n18356 , n18355 );
buf ( n18357 , n18340 );
buf ( n18358 , n18357 );
buf ( n18359 , n18340 );
buf ( n18360 , n18359 );
buf ( n18361 , n18340 );
buf ( n18362 , n18361 );
buf ( n18363 , n18340 );
buf ( n18364 , n18363 );
buf ( n18365 , n18340 );
buf ( n18366 , n18365 );
buf ( n18367 , n18340 );
buf ( n18368 , n18367 );
buf ( n18369 , n18340 );
buf ( n18370 , n18369 );
buf ( n18371 , n18340 );
buf ( n18372 , n18371 );
buf ( n18373 , n18340 );
buf ( n18374 , n18373 );
buf ( n18375 , n18340 );
buf ( n18376 , n18375 );
buf ( n18377 , n18340 );
buf ( n18378 , n18377 );
buf ( n18379 , n18340 );
buf ( n18380 , n18379 );
buf ( n18381 , n18340 );
buf ( n18382 , n18381 );
buf ( n18383 , n18340 );
buf ( n18384 , n18383 );
buf ( n18385 , n18340 );
buf ( n18386 , n18385 );
buf ( n18387 , n18340 );
buf ( n18388 , n18387 );
buf ( n18389 , n18340 );
buf ( n18390 , n18389 );
buf ( n18391 , n18340 );
buf ( n18392 , n18391 );
buf ( n18393 , n18340 );
buf ( n18394 , n18393 );
buf ( n18395 , n18340 );
buf ( n18396 , n18395 );
buf ( n18397 , n18340 );
buf ( n18398 , n18397 );
buf ( n18399 , n18340 );
buf ( n18400 , n18399 );
buf ( n18401 , n18340 );
buf ( n18402 , n18401 );
buf ( n18403 , n18340 );
buf ( n18404 , n18403 );
buf ( n18405 , n18340 );
buf ( n18406 , n18405 );
buf ( n18407 , n18340 );
buf ( n18408 , n18407 );
buf ( n18409 , n18340 );
buf ( n18410 , n18409 );
buf ( n18411 , n18340 );
buf ( n18412 , n18411 );
buf ( n18413 , n18340 );
buf ( n18414 , n18413 );
buf ( n18415 , n18340 );
buf ( n18416 , n18415 );
buf ( n18417 , n18340 );
buf ( n18418 , n18417 );
buf ( n18419 , n18340 );
buf ( n18420 , n18419 );
buf ( n18421 , n18340 );
buf ( n18422 , n18421 );
buf ( n18423 , n18340 );
buf ( n18424 , n18423 );
buf ( n18425 , n18340 );
buf ( n18426 , n18425 );
buf ( n18427 , n18340 );
buf ( n18428 , n18427 );
buf ( n18429 , n18340 );
buf ( n18430 , n18429 );
buf ( n18431 , n18340 );
buf ( n18432 , n18431 );
buf ( n18433 , n18340 );
buf ( n18434 , n18433 );
buf ( n18435 , n18340 );
buf ( n18436 , n18435 );
buf ( n18437 , n18340 );
buf ( n18438 , n18437 );
buf ( n18439 , n18340 );
buf ( n18440 , n18439 );
buf ( n18441 , n18340 );
buf ( n18442 , n18441 );
buf ( n18443 , n18340 );
buf ( n18444 , n18443 );
buf ( n18445 , n18340 );
buf ( n18446 , n18445 );
buf ( n18447 , n18340 );
buf ( n18448 , n18447 );
buf ( n18449 , n18340 );
buf ( n18450 , n18449 );
buf ( n18451 , n18340 );
buf ( n18452 , n18451 );
buf ( n18453 , n18340 );
buf ( n18454 , n18453 );
buf ( n18455 , n18340 );
buf ( n18456 , n18455 );
buf ( n18457 , n18340 );
buf ( n18458 , n18457 );
buf ( n18459 , n18340 );
buf ( n18460 , n18459 );
buf ( n18461 , n18340 );
buf ( n18462 , n18461 );
buf ( n18463 , n18340 );
buf ( n18464 , n18463 );
buf ( n18465 , n18340 );
buf ( n18466 , n18465 );
buf ( n18467 , n18340 );
buf ( n18468 , n18467 );
buf ( n18469 , n18340 );
buf ( n18470 , n18469 );
buf ( n18471 , n18340 );
buf ( n18472 , n18471 );
buf ( n18473 , n18340 );
buf ( n18474 , n18473 );
buf ( n18475 , n18340 );
buf ( n18476 , n18475 );
buf ( n18477 , n18340 );
buf ( n18478 , n18477 );
buf ( n18479 , n18340 );
buf ( n18480 , n18479 );
buf ( n18481 , n18340 );
buf ( n18482 , n18481 );
buf ( n18483 , n18340 );
buf ( n18484 , n18483 );
buf ( n18485 , n18340 );
buf ( n18486 , n18485 );
buf ( n18487 , n18340 );
buf ( n18488 , n18487 );
buf ( n18489 , n18340 );
buf ( n18490 , n18489 );
buf ( n18491 , n18340 );
buf ( n18492 , n18491 );
buf ( n18493 , n18340 );
buf ( n18494 , n18493 );
buf ( n18495 , n18340 );
buf ( n18496 , n18495 );
buf ( n18497 , n18340 );
buf ( n18498 , n18497 );
buf ( n18499 , n18340 );
buf ( n18500 , n18499 );
buf ( n18501 , n18340 );
buf ( n18502 , n18501 );
buf ( n18503 , n18340 );
buf ( n18504 , n18503 );
buf ( n18505 , n18340 );
buf ( n18506 , n18505 );
buf ( n18507 , n18340 );
buf ( n18508 , n18507 );
buf ( n18509 , n18340 );
buf ( n18510 , n18509 );
buf ( n18511 , n18340 );
buf ( n18512 , n18511 );
buf ( n18513 , n18340 );
buf ( n18514 , n18513 );
buf ( n18515 , n18340 );
buf ( n18516 , n18515 );
buf ( n18517 , n18340 );
buf ( n18518 , n18517 );
buf ( n18519 , n18340 );
buf ( n18520 , n18519 );
buf ( n18521 , n18340 );
buf ( n18522 , n18521 );
buf ( n18523 , n18340 );
buf ( n18524 , n18523 );
buf ( n18525 , n18340 );
buf ( n18526 , n18525 );
buf ( n18527 , n18340 );
buf ( n18528 , n18527 );
buf ( n18529 , n18340 );
buf ( n18530 , n18529 );
buf ( n18531 , n18340 );
buf ( n18532 , n18531 );
xor ( n18533 , n18123 , n18125 );
xor ( n18534 , n18533 , n18336 );
buf ( n18535 , n18534 );
buf ( n18536 , n18535 );
xor ( n18537 , n18127 , n18129 );
xor ( n18538 , n18537 , n18333 );
buf ( n18539 , n18538 );
buf ( n18540 , n18539 );
xor ( n18541 , n18131 , n18133 );
xor ( n18542 , n18541 , n18330 );
buf ( n18543 , n18542 );
buf ( n18544 , n18543 );
xor ( n18545 , n18135 , n18137 );
xor ( n18546 , n18545 , n18327 );
buf ( n18547 , n18546 );
buf ( n18548 , n18547 );
xor ( n18549 , n18139 , n18141 );
xor ( n18550 , n18549 , n18324 );
buf ( n18551 , n18550 );
buf ( n18552 , n18551 );
xor ( n18553 , n18143 , n18145 );
xor ( n18554 , n18553 , n18321 );
buf ( n18555 , n18554 );
buf ( n18556 , n18555 );
xor ( n18557 , n18147 , n18149 );
xor ( n18558 , n18557 , n18318 );
buf ( n18559 , n18558 );
buf ( n18560 , n18559 );
xor ( n18561 , n18151 , n18153 );
xor ( n18562 , n18561 , n18315 );
buf ( n18563 , n18562 );
buf ( n18564 , n18563 );
xor ( n18565 , n18155 , n18157 );
xor ( n18566 , n18565 , n18312 );
buf ( n18567 , n18566 );
buf ( n18568 , n18567 );
xor ( n18569 , n18159 , n18161 );
xor ( n18570 , n18569 , n18309 );
buf ( n18571 , n18570 );
buf ( n18572 , n18571 );
xor ( n18573 , n18163 , n18165 );
xor ( n18574 , n18573 , n18306 );
buf ( n18575 , n18574 );
buf ( n18576 , n18575 );
xor ( n18577 , n18167 , n18169 );
xor ( n18578 , n18577 , n18303 );
buf ( n18579 , n18578 );
buf ( n18580 , n18579 );
xor ( n18581 , n18171 , n18173 );
xor ( n18582 , n18581 , n18300 );
buf ( n18583 , n18582 );
buf ( n18584 , n18583 );
xor ( n18585 , n18175 , n18177 );
xor ( n18586 , n18585 , n18297 );
buf ( n18587 , n18586 );
buf ( n18588 , n18587 );
xor ( n18589 , n18179 , n18181 );
xor ( n18590 , n18589 , n18294 );
buf ( n18591 , n18590 );
buf ( n18592 , n18591 );
xor ( n18593 , n18183 , n18185 );
xor ( n18594 , n18593 , n18291 );
buf ( n18595 , n18594 );
buf ( n18596 , n18595 );
xor ( n18597 , n18187 , n18189 );
xor ( n18598 , n18597 , n18288 );
buf ( n18599 , n18598 );
buf ( n18600 , n18599 );
xor ( n18601 , n18191 , n18193 );
xor ( n18602 , n18601 , n18285 );
buf ( n18603 , n18602 );
buf ( n18604 , n18603 );
xor ( n18605 , n18195 , n18197 );
xor ( n18606 , n18605 , n18282 );
buf ( n18607 , n18606 );
buf ( n18608 , n18607 );
xor ( n18609 , n18199 , n18201 );
xor ( n18610 , n18609 , n18279 );
buf ( n18611 , n18610 );
buf ( n18612 , n18611 );
xor ( n18613 , n18203 , n18205 );
xor ( n18614 , n18613 , n18276 );
buf ( n18615 , n18614 );
buf ( n18616 , n18615 );
xor ( n18617 , n18207 , n18209 );
xor ( n18618 , n18617 , n18273 );
buf ( n18619 , n18618 );
buf ( n18620 , n18619 );
xor ( n18621 , n18211 , n18213 );
xor ( n18622 , n18621 , n18270 );
buf ( n18623 , n18622 );
buf ( n18624 , n18623 );
xor ( n18625 , n18215 , n18217 );
xor ( n18626 , n18625 , n18267 );
buf ( n18627 , n18626 );
buf ( n18628 , n18627 );
xor ( n18629 , n18219 , n18221 );
xor ( n18630 , n18629 , n18264 );
buf ( n18631 , n18630 );
buf ( n18632 , n18631 );
xor ( n18633 , n18223 , n18225 );
xor ( n18634 , n18633 , n18261 );
buf ( n18635 , n18634 );
buf ( n18636 , n18635 );
xor ( n18637 , n18227 , n18229 );
xor ( n18638 , n18637 , n18258 );
buf ( n18639 , n18638 );
buf ( n18640 , n18639 );
xor ( n18641 , n18231 , n18233 );
xor ( n18642 , n18641 , n18255 );
buf ( n18643 , n18642 );
buf ( n18644 , n18643 );
xor ( n18645 , n18235 , n18237 );
xor ( n18646 , n18645 , n18252 );
buf ( n18647 , n18646 );
buf ( n18648 , n18647 );
xor ( n18649 , n18239 , n18241 );
xor ( n18650 , n18649 , n18249 );
buf ( n18651 , n18650 );
buf ( n18652 , n18651 );
xor ( n18653 , n18243 , n18245 );
not ( n18654 , n18653 );
buf ( n18655 , n18654 );
buf ( n18656 , n18655 );
and ( n18657 , n18107 , n18652 );
buf ( n18658 , n18657 );
and ( n18659 , n18107 , n18656 );
buf ( n18660 , n18659 );
and ( n18661 , n18108 , n18652 );
and ( n18662 , n18660 , n18661 );
xor ( n18663 , n18660 , n18661 );
and ( n18664 , n18108 , n18656 );
buf ( n18665 , n18664 );
buf ( n18666 , n18665 );
and ( n18667 , n18109 , n18652 );
and ( n18668 , n18666 , n18667 );
xor ( n18669 , n18666 , n18667 );
and ( n18670 , n18109 , n18656 );
buf ( n18671 , n18670 );
buf ( n18672 , n18671 );
and ( n18673 , n18110 , n18652 );
and ( n18674 , n18672 , n18673 );
xor ( n18675 , n18672 , n18673 );
and ( n18676 , n18110 , n18656 );
buf ( n18677 , n18676 );
buf ( n18678 , n18677 );
and ( n18679 , n18111 , n18652 );
and ( n18680 , n18678 , n18679 );
xor ( n18681 , n18678 , n18679 );
and ( n18682 , n18111 , n18656 );
buf ( n18683 , n18682 );
buf ( n18684 , n18683 );
and ( n18685 , n18112 , n18652 );
and ( n18686 , n18684 , n18685 );
xor ( n18687 , n18684 , n18685 );
and ( n18688 , n18112 , n18656 );
buf ( n18689 , n18688 );
buf ( n18690 , n18689 );
and ( n18691 , n18113 , n18652 );
and ( n18692 , n18690 , n18691 );
xor ( n18693 , n18690 , n18691 );
and ( n18694 , n18113 , n18656 );
buf ( n18695 , n18694 );
buf ( n18696 , n18695 );
and ( n18697 , n18114 , n18652 );
and ( n18698 , n18696 , n18697 );
xor ( n18699 , n18696 , n18697 );
and ( n18700 , n18114 , n18656 );
buf ( n18701 , n18700 );
buf ( n18702 , n18701 );
and ( n18703 , n18115 , n18652 );
and ( n18704 , n18702 , n18703 );
xor ( n18705 , n18702 , n18703 );
and ( n18706 , n18115 , n18656 );
buf ( n18707 , n18706 );
buf ( n18708 , n18707 );
and ( n18709 , n18116 , n18652 );
and ( n18710 , n18708 , n18709 );
xor ( n18711 , n18708 , n18709 );
and ( n18712 , n18116 , n18656 );
buf ( n18713 , n18712 );
buf ( n18714 , n18713 );
and ( n18715 , n18117 , n18652 );
and ( n18716 , n18714 , n18715 );
xor ( n18717 , n18714 , n18715 );
and ( n18718 , n18117 , n18656 );
buf ( n18719 , n18718 );
buf ( n18720 , n18719 );
and ( n18721 , n18118 , n18652 );
and ( n18722 , n18720 , n18721 );
xor ( n18723 , n18720 , n18721 );
and ( n18724 , n18118 , n18656 );
buf ( n18725 , n18724 );
buf ( n18726 , n18725 );
and ( n18727 , n18119 , n18652 );
and ( n18728 , n18726 , n18727 );
xor ( n18729 , n18726 , n18727 );
and ( n18730 , n18119 , n18656 );
buf ( n18731 , n18730 );
buf ( n18732 , n18731 );
and ( n18733 , n18120 , n18652 );
and ( n18734 , n18732 , n18733 );
xor ( n18735 , n18732 , n18733 );
and ( n18736 , n18120 , n18656 );
buf ( n18737 , n18736 );
buf ( n18738 , n18737 );
and ( n18739 , n18121 , n18652 );
and ( n18740 , n18738 , n18739 );
xor ( n18741 , n18738 , n18739 );
and ( n18742 , n18121 , n18656 );
buf ( n18743 , n18742 );
buf ( n18744 , n18743 );
and ( n18745 , n18122 , n18652 );
and ( n18746 , n18744 , n18745 );
and ( n18747 , n18741 , n18746 );
or ( n18748 , n18740 , n18747 );
and ( n18749 , n18735 , n18748 );
or ( n18750 , n18734 , n18749 );
and ( n18751 , n18729 , n18750 );
or ( n18752 , n18728 , n18751 );
and ( n18753 , n18723 , n18752 );
or ( n18754 , n18722 , n18753 );
and ( n18755 , n18717 , n18754 );
or ( n18756 , n18716 , n18755 );
and ( n18757 , n18711 , n18756 );
or ( n18758 , n18710 , n18757 );
and ( n18759 , n18705 , n18758 );
or ( n18760 , n18704 , n18759 );
and ( n18761 , n18699 , n18760 );
or ( n18762 , n18698 , n18761 );
and ( n18763 , n18693 , n18762 );
or ( n18764 , n18692 , n18763 );
and ( n18765 , n18687 , n18764 );
or ( n18766 , n18686 , n18765 );
and ( n18767 , n18681 , n18766 );
or ( n18768 , n18680 , n18767 );
and ( n18769 , n18675 , n18768 );
or ( n18770 , n18674 , n18769 );
and ( n18771 , n18669 , n18770 );
or ( n18772 , n18668 , n18771 );
and ( n18773 , n18663 , n18772 );
or ( n18774 , n18662 , n18773 );
and ( n18775 , n18658 , n18774 );
buf ( n18776 , n18775 );
and ( n18777 , n18107 , n18648 );
and ( n18778 , n18776 , n18777 );
xor ( n18779 , n18776 , n18777 );
xor ( n18780 , n18658 , n18774 );
and ( n18781 , n18108 , n18648 );
and ( n18782 , n18780 , n18781 );
xor ( n18783 , n18780 , n18781 );
xor ( n18784 , n18663 , n18772 );
and ( n18785 , n18109 , n18648 );
and ( n18786 , n18784 , n18785 );
xor ( n18787 , n18784 , n18785 );
xor ( n18788 , n18669 , n18770 );
and ( n18789 , n18110 , n18648 );
and ( n18790 , n18788 , n18789 );
xor ( n18791 , n18788 , n18789 );
xor ( n18792 , n18675 , n18768 );
and ( n18793 , n18111 , n18648 );
and ( n18794 , n18792 , n18793 );
xor ( n18795 , n18792 , n18793 );
xor ( n18796 , n18681 , n18766 );
and ( n18797 , n18112 , n18648 );
and ( n18798 , n18796 , n18797 );
xor ( n18799 , n18796 , n18797 );
xor ( n18800 , n18687 , n18764 );
and ( n18801 , n18113 , n18648 );
and ( n18802 , n18800 , n18801 );
xor ( n18803 , n18800 , n18801 );
xor ( n18804 , n18693 , n18762 );
and ( n18805 , n18114 , n18648 );
and ( n18806 , n18804 , n18805 );
xor ( n18807 , n18804 , n18805 );
xor ( n18808 , n18699 , n18760 );
and ( n18809 , n18115 , n18648 );
and ( n18810 , n18808 , n18809 );
xor ( n18811 , n18808 , n18809 );
xor ( n18812 , n18705 , n18758 );
and ( n18813 , n18116 , n18648 );
and ( n18814 , n18812 , n18813 );
xor ( n18815 , n18812 , n18813 );
xor ( n18816 , n18711 , n18756 );
and ( n18817 , n18117 , n18648 );
and ( n18818 , n18816 , n18817 );
xor ( n18819 , n18816 , n18817 );
xor ( n18820 , n18717 , n18754 );
and ( n18821 , n18118 , n18648 );
and ( n18822 , n18820 , n18821 );
xor ( n18823 , n18820 , n18821 );
xor ( n18824 , n18723 , n18752 );
and ( n18825 , n18119 , n18648 );
and ( n18826 , n18824 , n18825 );
xor ( n18827 , n18824 , n18825 );
xor ( n18828 , n18729 , n18750 );
and ( n18829 , n18120 , n18648 );
and ( n18830 , n18828 , n18829 );
xor ( n18831 , n18828 , n18829 );
xor ( n18832 , n18735 , n18748 );
and ( n18833 , n18121 , n18648 );
and ( n18834 , n18832 , n18833 );
xor ( n18835 , n18832 , n18833 );
xor ( n18836 , n18741 , n18746 );
and ( n18837 , n18122 , n18648 );
and ( n18838 , n18836 , n18837 );
and ( n18839 , n18835 , n18838 );
or ( n18840 , n18834 , n18839 );
and ( n18841 , n18831 , n18840 );
or ( n18842 , n18830 , n18841 );
and ( n18843 , n18827 , n18842 );
or ( n18844 , n18826 , n18843 );
and ( n18845 , n18823 , n18844 );
or ( n18846 , n18822 , n18845 );
and ( n18847 , n18819 , n18846 );
or ( n18848 , n18818 , n18847 );
and ( n18849 , n18815 , n18848 );
or ( n18850 , n18814 , n18849 );
and ( n18851 , n18811 , n18850 );
or ( n18852 , n18810 , n18851 );
and ( n18853 , n18807 , n18852 );
or ( n18854 , n18806 , n18853 );
and ( n18855 , n18803 , n18854 );
or ( n18856 , n18802 , n18855 );
and ( n18857 , n18799 , n18856 );
or ( n18858 , n18798 , n18857 );
and ( n18859 , n18795 , n18858 );
or ( n18860 , n18794 , n18859 );
and ( n18861 , n18791 , n18860 );
or ( n18862 , n18790 , n18861 );
and ( n18863 , n18787 , n18862 );
or ( n18864 , n18786 , n18863 );
and ( n18865 , n18783 , n18864 );
or ( n18866 , n18782 , n18865 );
and ( n18867 , n18779 , n18866 );
or ( n18868 , n18778 , n18867 );
and ( n18869 , n18107 , n18644 );
and ( n18870 , n18868 , n18869 );
xor ( n18871 , n18868 , n18869 );
xor ( n18872 , n18779 , n18866 );
and ( n18873 , n18108 , n18644 );
and ( n18874 , n18872 , n18873 );
xor ( n18875 , n18872 , n18873 );
xor ( n18876 , n18783 , n18864 );
and ( n18877 , n18109 , n18644 );
and ( n18878 , n18876 , n18877 );
xor ( n18879 , n18876 , n18877 );
xor ( n18880 , n18787 , n18862 );
and ( n18881 , n18110 , n18644 );
and ( n18882 , n18880 , n18881 );
xor ( n18883 , n18880 , n18881 );
xor ( n18884 , n18791 , n18860 );
and ( n18885 , n18111 , n18644 );
and ( n18886 , n18884 , n18885 );
xor ( n18887 , n18884 , n18885 );
xor ( n18888 , n18795 , n18858 );
and ( n18889 , n18112 , n18644 );
and ( n18890 , n18888 , n18889 );
xor ( n18891 , n18888 , n18889 );
xor ( n18892 , n18799 , n18856 );
and ( n18893 , n18113 , n18644 );
and ( n18894 , n18892 , n18893 );
xor ( n18895 , n18892 , n18893 );
xor ( n18896 , n18803 , n18854 );
and ( n18897 , n18114 , n18644 );
and ( n18898 , n18896 , n18897 );
xor ( n18899 , n18896 , n18897 );
xor ( n18900 , n18807 , n18852 );
and ( n18901 , n18115 , n18644 );
and ( n18902 , n18900 , n18901 );
xor ( n18903 , n18900 , n18901 );
xor ( n18904 , n18811 , n18850 );
and ( n18905 , n18116 , n18644 );
and ( n18906 , n18904 , n18905 );
xor ( n18907 , n18904 , n18905 );
xor ( n18908 , n18815 , n18848 );
and ( n18909 , n18117 , n18644 );
and ( n18910 , n18908 , n18909 );
xor ( n18911 , n18908 , n18909 );
xor ( n18912 , n18819 , n18846 );
and ( n18913 , n18118 , n18644 );
and ( n18914 , n18912 , n18913 );
xor ( n18915 , n18912 , n18913 );
xor ( n18916 , n18823 , n18844 );
and ( n18917 , n18119 , n18644 );
and ( n18918 , n18916 , n18917 );
xor ( n18919 , n18916 , n18917 );
xor ( n18920 , n18827 , n18842 );
and ( n18921 , n18120 , n18644 );
and ( n18922 , n18920 , n18921 );
xor ( n18923 , n18920 , n18921 );
xor ( n18924 , n18831 , n18840 );
and ( n18925 , n18121 , n18644 );
and ( n18926 , n18924 , n18925 );
xor ( n18927 , n18924 , n18925 );
xor ( n18928 , n18835 , n18838 );
and ( n18929 , n18122 , n18644 );
and ( n18930 , n18928 , n18929 );
and ( n18931 , n18927 , n18930 );
or ( n18932 , n18926 , n18931 );
and ( n18933 , n18923 , n18932 );
or ( n18934 , n18922 , n18933 );
and ( n18935 , n18919 , n18934 );
or ( n18936 , n18918 , n18935 );
and ( n18937 , n18915 , n18936 );
or ( n18938 , n18914 , n18937 );
and ( n18939 , n18911 , n18938 );
or ( n18940 , n18910 , n18939 );
and ( n18941 , n18907 , n18940 );
or ( n18942 , n18906 , n18941 );
and ( n18943 , n18903 , n18942 );
or ( n18944 , n18902 , n18943 );
and ( n18945 , n18899 , n18944 );
or ( n18946 , n18898 , n18945 );
and ( n18947 , n18895 , n18946 );
or ( n18948 , n18894 , n18947 );
and ( n18949 , n18891 , n18948 );
or ( n18950 , n18890 , n18949 );
and ( n18951 , n18887 , n18950 );
or ( n18952 , n18886 , n18951 );
and ( n18953 , n18883 , n18952 );
or ( n18954 , n18882 , n18953 );
and ( n18955 , n18879 , n18954 );
or ( n18956 , n18878 , n18955 );
and ( n18957 , n18875 , n18956 );
or ( n18958 , n18874 , n18957 );
and ( n18959 , n18871 , n18958 );
or ( n18960 , n18870 , n18959 );
and ( n18961 , n18107 , n18640 );
and ( n18962 , n18960 , n18961 );
xor ( n18963 , n18960 , n18961 );
xor ( n18964 , n18871 , n18958 );
and ( n18965 , n18108 , n18640 );
and ( n18966 , n18964 , n18965 );
xor ( n18967 , n18964 , n18965 );
xor ( n18968 , n18875 , n18956 );
and ( n18969 , n18109 , n18640 );
and ( n18970 , n18968 , n18969 );
xor ( n18971 , n18968 , n18969 );
xor ( n18972 , n18879 , n18954 );
and ( n18973 , n18110 , n18640 );
and ( n18974 , n18972 , n18973 );
xor ( n18975 , n18972 , n18973 );
xor ( n18976 , n18883 , n18952 );
and ( n18977 , n18111 , n18640 );
and ( n18978 , n18976 , n18977 );
xor ( n18979 , n18976 , n18977 );
xor ( n18980 , n18887 , n18950 );
and ( n18981 , n18112 , n18640 );
and ( n18982 , n18980 , n18981 );
xor ( n18983 , n18980 , n18981 );
xor ( n18984 , n18891 , n18948 );
and ( n18985 , n18113 , n18640 );
and ( n18986 , n18984 , n18985 );
xor ( n18987 , n18984 , n18985 );
xor ( n18988 , n18895 , n18946 );
and ( n18989 , n18114 , n18640 );
and ( n18990 , n18988 , n18989 );
xor ( n18991 , n18988 , n18989 );
xor ( n18992 , n18899 , n18944 );
and ( n18993 , n18115 , n18640 );
and ( n18994 , n18992 , n18993 );
xor ( n18995 , n18992 , n18993 );
xor ( n18996 , n18903 , n18942 );
and ( n18997 , n18116 , n18640 );
and ( n18998 , n18996 , n18997 );
xor ( n18999 , n18996 , n18997 );
xor ( n19000 , n18907 , n18940 );
and ( n19001 , n18117 , n18640 );
and ( n19002 , n19000 , n19001 );
xor ( n19003 , n19000 , n19001 );
xor ( n19004 , n18911 , n18938 );
and ( n19005 , n18118 , n18640 );
and ( n19006 , n19004 , n19005 );
xor ( n19007 , n19004 , n19005 );
xor ( n19008 , n18915 , n18936 );
and ( n19009 , n18119 , n18640 );
and ( n19010 , n19008 , n19009 );
xor ( n19011 , n19008 , n19009 );
xor ( n19012 , n18919 , n18934 );
and ( n19013 , n18120 , n18640 );
and ( n19014 , n19012 , n19013 );
xor ( n19015 , n19012 , n19013 );
xor ( n19016 , n18923 , n18932 );
and ( n19017 , n18121 , n18640 );
and ( n19018 , n19016 , n19017 );
xor ( n19019 , n19016 , n19017 );
xor ( n19020 , n18927 , n18930 );
and ( n19021 , n18122 , n18640 );
and ( n19022 , n19020 , n19021 );
and ( n19023 , n19019 , n19022 );
or ( n19024 , n19018 , n19023 );
and ( n19025 , n19015 , n19024 );
or ( n19026 , n19014 , n19025 );
and ( n19027 , n19011 , n19026 );
or ( n19028 , n19010 , n19027 );
and ( n19029 , n19007 , n19028 );
or ( n19030 , n19006 , n19029 );
and ( n19031 , n19003 , n19030 );
or ( n19032 , n19002 , n19031 );
and ( n19033 , n18999 , n19032 );
or ( n19034 , n18998 , n19033 );
and ( n19035 , n18995 , n19034 );
or ( n19036 , n18994 , n19035 );
and ( n19037 , n18991 , n19036 );
or ( n19038 , n18990 , n19037 );
and ( n19039 , n18987 , n19038 );
or ( n19040 , n18986 , n19039 );
and ( n19041 , n18983 , n19040 );
or ( n19042 , n18982 , n19041 );
and ( n19043 , n18979 , n19042 );
or ( n19044 , n18978 , n19043 );
and ( n19045 , n18975 , n19044 );
or ( n19046 , n18974 , n19045 );
and ( n19047 , n18971 , n19046 );
or ( n19048 , n18970 , n19047 );
and ( n19049 , n18967 , n19048 );
or ( n19050 , n18966 , n19049 );
and ( n19051 , n18963 , n19050 );
or ( n19052 , n18962 , n19051 );
and ( n19053 , n18107 , n18636 );
and ( n19054 , n19052 , n19053 );
xor ( n19055 , n19052 , n19053 );
xor ( n19056 , n18963 , n19050 );
and ( n19057 , n18108 , n18636 );
and ( n19058 , n19056 , n19057 );
xor ( n19059 , n19056 , n19057 );
xor ( n19060 , n18967 , n19048 );
and ( n19061 , n18109 , n18636 );
and ( n19062 , n19060 , n19061 );
xor ( n19063 , n19060 , n19061 );
xor ( n19064 , n18971 , n19046 );
and ( n19065 , n18110 , n18636 );
and ( n19066 , n19064 , n19065 );
xor ( n19067 , n19064 , n19065 );
xor ( n19068 , n18975 , n19044 );
and ( n19069 , n18111 , n18636 );
and ( n19070 , n19068 , n19069 );
xor ( n19071 , n19068 , n19069 );
xor ( n19072 , n18979 , n19042 );
and ( n19073 , n18112 , n18636 );
and ( n19074 , n19072 , n19073 );
xor ( n19075 , n19072 , n19073 );
xor ( n19076 , n18983 , n19040 );
and ( n19077 , n18113 , n18636 );
and ( n19078 , n19076 , n19077 );
xor ( n19079 , n19076 , n19077 );
xor ( n19080 , n18987 , n19038 );
and ( n19081 , n18114 , n18636 );
and ( n19082 , n19080 , n19081 );
xor ( n19083 , n19080 , n19081 );
xor ( n19084 , n18991 , n19036 );
and ( n19085 , n18115 , n18636 );
and ( n19086 , n19084 , n19085 );
xor ( n19087 , n19084 , n19085 );
xor ( n19088 , n18995 , n19034 );
and ( n19089 , n18116 , n18636 );
and ( n19090 , n19088 , n19089 );
xor ( n19091 , n19088 , n19089 );
xor ( n19092 , n18999 , n19032 );
and ( n19093 , n18117 , n18636 );
and ( n19094 , n19092 , n19093 );
xor ( n19095 , n19092 , n19093 );
xor ( n19096 , n19003 , n19030 );
and ( n19097 , n18118 , n18636 );
and ( n19098 , n19096 , n19097 );
xor ( n19099 , n19096 , n19097 );
xor ( n19100 , n19007 , n19028 );
and ( n19101 , n18119 , n18636 );
and ( n19102 , n19100 , n19101 );
xor ( n19103 , n19100 , n19101 );
xor ( n19104 , n19011 , n19026 );
and ( n19105 , n18120 , n18636 );
and ( n19106 , n19104 , n19105 );
xor ( n19107 , n19104 , n19105 );
xor ( n19108 , n19015 , n19024 );
and ( n19109 , n18121 , n18636 );
and ( n19110 , n19108 , n19109 );
xor ( n19111 , n19108 , n19109 );
xor ( n19112 , n19019 , n19022 );
and ( n19113 , n18122 , n18636 );
and ( n19114 , n19112 , n19113 );
and ( n19115 , n19111 , n19114 );
or ( n19116 , n19110 , n19115 );
and ( n19117 , n19107 , n19116 );
or ( n19118 , n19106 , n19117 );
and ( n19119 , n19103 , n19118 );
or ( n19120 , n19102 , n19119 );
and ( n19121 , n19099 , n19120 );
or ( n19122 , n19098 , n19121 );
and ( n19123 , n19095 , n19122 );
or ( n19124 , n19094 , n19123 );
and ( n19125 , n19091 , n19124 );
or ( n19126 , n19090 , n19125 );
and ( n19127 , n19087 , n19126 );
or ( n19128 , n19086 , n19127 );
and ( n19129 , n19083 , n19128 );
or ( n19130 , n19082 , n19129 );
and ( n19131 , n19079 , n19130 );
or ( n19132 , n19078 , n19131 );
and ( n19133 , n19075 , n19132 );
or ( n19134 , n19074 , n19133 );
and ( n19135 , n19071 , n19134 );
or ( n19136 , n19070 , n19135 );
and ( n19137 , n19067 , n19136 );
or ( n19138 , n19066 , n19137 );
and ( n19139 , n19063 , n19138 );
or ( n19140 , n19062 , n19139 );
and ( n19141 , n19059 , n19140 );
or ( n19142 , n19058 , n19141 );
and ( n19143 , n19055 , n19142 );
or ( n19144 , n19054 , n19143 );
and ( n19145 , n18107 , n18632 );
and ( n19146 , n19144 , n19145 );
xor ( n19147 , n19144 , n19145 );
xor ( n19148 , n19055 , n19142 );
and ( n19149 , n18108 , n18632 );
and ( n19150 , n19148 , n19149 );
xor ( n19151 , n19148 , n19149 );
xor ( n19152 , n19059 , n19140 );
and ( n19153 , n18109 , n18632 );
and ( n19154 , n19152 , n19153 );
xor ( n19155 , n19152 , n19153 );
xor ( n19156 , n19063 , n19138 );
and ( n19157 , n18110 , n18632 );
and ( n19158 , n19156 , n19157 );
xor ( n19159 , n19156 , n19157 );
xor ( n19160 , n19067 , n19136 );
and ( n19161 , n18111 , n18632 );
and ( n19162 , n19160 , n19161 );
xor ( n19163 , n19160 , n19161 );
xor ( n19164 , n19071 , n19134 );
and ( n19165 , n18112 , n18632 );
and ( n19166 , n19164 , n19165 );
xor ( n19167 , n19164 , n19165 );
xor ( n19168 , n19075 , n19132 );
and ( n19169 , n18113 , n18632 );
and ( n19170 , n19168 , n19169 );
xor ( n19171 , n19168 , n19169 );
xor ( n19172 , n19079 , n19130 );
and ( n19173 , n18114 , n18632 );
and ( n19174 , n19172 , n19173 );
xor ( n19175 , n19172 , n19173 );
xor ( n19176 , n19083 , n19128 );
and ( n19177 , n18115 , n18632 );
and ( n19178 , n19176 , n19177 );
xor ( n19179 , n19176 , n19177 );
xor ( n19180 , n19087 , n19126 );
and ( n19181 , n18116 , n18632 );
and ( n19182 , n19180 , n19181 );
xor ( n19183 , n19180 , n19181 );
xor ( n19184 , n19091 , n19124 );
and ( n19185 , n18117 , n18632 );
and ( n19186 , n19184 , n19185 );
xor ( n19187 , n19184 , n19185 );
xor ( n19188 , n19095 , n19122 );
and ( n19189 , n18118 , n18632 );
and ( n19190 , n19188 , n19189 );
xor ( n19191 , n19188 , n19189 );
xor ( n19192 , n19099 , n19120 );
and ( n19193 , n18119 , n18632 );
and ( n19194 , n19192 , n19193 );
xor ( n19195 , n19192 , n19193 );
xor ( n19196 , n19103 , n19118 );
and ( n19197 , n18120 , n18632 );
and ( n19198 , n19196 , n19197 );
xor ( n19199 , n19196 , n19197 );
xor ( n19200 , n19107 , n19116 );
and ( n19201 , n18121 , n18632 );
and ( n19202 , n19200 , n19201 );
xor ( n19203 , n19200 , n19201 );
xor ( n19204 , n19111 , n19114 );
and ( n19205 , n18122 , n18632 );
and ( n19206 , n19204 , n19205 );
and ( n19207 , n19203 , n19206 );
or ( n19208 , n19202 , n19207 );
and ( n19209 , n19199 , n19208 );
or ( n19210 , n19198 , n19209 );
and ( n19211 , n19195 , n19210 );
or ( n19212 , n19194 , n19211 );
and ( n19213 , n19191 , n19212 );
or ( n19214 , n19190 , n19213 );
and ( n19215 , n19187 , n19214 );
or ( n19216 , n19186 , n19215 );
and ( n19217 , n19183 , n19216 );
or ( n19218 , n19182 , n19217 );
and ( n19219 , n19179 , n19218 );
or ( n19220 , n19178 , n19219 );
and ( n19221 , n19175 , n19220 );
or ( n19222 , n19174 , n19221 );
and ( n19223 , n19171 , n19222 );
or ( n19224 , n19170 , n19223 );
and ( n19225 , n19167 , n19224 );
or ( n19226 , n19166 , n19225 );
and ( n19227 , n19163 , n19226 );
or ( n19228 , n19162 , n19227 );
and ( n19229 , n19159 , n19228 );
or ( n19230 , n19158 , n19229 );
and ( n19231 , n19155 , n19230 );
or ( n19232 , n19154 , n19231 );
and ( n19233 , n19151 , n19232 );
or ( n19234 , n19150 , n19233 );
and ( n19235 , n19147 , n19234 );
or ( n19236 , n19146 , n19235 );
and ( n19237 , n18107 , n18628 );
and ( n19238 , n19236 , n19237 );
xor ( n19239 , n19236 , n19237 );
xor ( n19240 , n19147 , n19234 );
and ( n19241 , n18108 , n18628 );
and ( n19242 , n19240 , n19241 );
xor ( n19243 , n19240 , n19241 );
xor ( n19244 , n19151 , n19232 );
and ( n19245 , n18109 , n18628 );
and ( n19246 , n19244 , n19245 );
xor ( n19247 , n19244 , n19245 );
xor ( n19248 , n19155 , n19230 );
and ( n19249 , n18110 , n18628 );
and ( n19250 , n19248 , n19249 );
xor ( n19251 , n19248 , n19249 );
xor ( n19252 , n19159 , n19228 );
and ( n19253 , n18111 , n18628 );
and ( n19254 , n19252 , n19253 );
xor ( n19255 , n19252 , n19253 );
xor ( n19256 , n19163 , n19226 );
and ( n19257 , n18112 , n18628 );
and ( n19258 , n19256 , n19257 );
xor ( n19259 , n19256 , n19257 );
xor ( n19260 , n19167 , n19224 );
and ( n19261 , n18113 , n18628 );
and ( n19262 , n19260 , n19261 );
xor ( n19263 , n19260 , n19261 );
xor ( n19264 , n19171 , n19222 );
and ( n19265 , n18114 , n18628 );
and ( n19266 , n19264 , n19265 );
xor ( n19267 , n19264 , n19265 );
xor ( n19268 , n19175 , n19220 );
and ( n19269 , n18115 , n18628 );
and ( n19270 , n19268 , n19269 );
xor ( n19271 , n19268 , n19269 );
xor ( n19272 , n19179 , n19218 );
and ( n19273 , n18116 , n18628 );
and ( n19274 , n19272 , n19273 );
xor ( n19275 , n19272 , n19273 );
xor ( n19276 , n19183 , n19216 );
and ( n19277 , n18117 , n18628 );
and ( n19278 , n19276 , n19277 );
xor ( n19279 , n19276 , n19277 );
xor ( n19280 , n19187 , n19214 );
and ( n19281 , n18118 , n18628 );
and ( n19282 , n19280 , n19281 );
xor ( n19283 , n19280 , n19281 );
xor ( n19284 , n19191 , n19212 );
and ( n19285 , n18119 , n18628 );
and ( n19286 , n19284 , n19285 );
xor ( n19287 , n19284 , n19285 );
xor ( n19288 , n19195 , n19210 );
and ( n19289 , n18120 , n18628 );
and ( n19290 , n19288 , n19289 );
xor ( n19291 , n19288 , n19289 );
xor ( n19292 , n19199 , n19208 );
and ( n19293 , n18121 , n18628 );
and ( n19294 , n19292 , n19293 );
xor ( n19295 , n19292 , n19293 );
xor ( n19296 , n19203 , n19206 );
and ( n19297 , n18122 , n18628 );
and ( n19298 , n19296 , n19297 );
and ( n19299 , n19295 , n19298 );
or ( n19300 , n19294 , n19299 );
and ( n19301 , n19291 , n19300 );
or ( n19302 , n19290 , n19301 );
and ( n19303 , n19287 , n19302 );
or ( n19304 , n19286 , n19303 );
and ( n19305 , n19283 , n19304 );
or ( n19306 , n19282 , n19305 );
and ( n19307 , n19279 , n19306 );
or ( n19308 , n19278 , n19307 );
and ( n19309 , n19275 , n19308 );
or ( n19310 , n19274 , n19309 );
and ( n19311 , n19271 , n19310 );
or ( n19312 , n19270 , n19311 );
and ( n19313 , n19267 , n19312 );
or ( n19314 , n19266 , n19313 );
and ( n19315 , n19263 , n19314 );
or ( n19316 , n19262 , n19315 );
and ( n19317 , n19259 , n19316 );
or ( n19318 , n19258 , n19317 );
and ( n19319 , n19255 , n19318 );
or ( n19320 , n19254 , n19319 );
and ( n19321 , n19251 , n19320 );
or ( n19322 , n19250 , n19321 );
and ( n19323 , n19247 , n19322 );
or ( n19324 , n19246 , n19323 );
and ( n19325 , n19243 , n19324 );
or ( n19326 , n19242 , n19325 );
and ( n19327 , n19239 , n19326 );
or ( n19328 , n19238 , n19327 );
and ( n19329 , n18107 , n18624 );
and ( n19330 , n19328 , n19329 );
xor ( n19331 , n19328 , n19329 );
xor ( n19332 , n19239 , n19326 );
and ( n19333 , n18108 , n18624 );
and ( n19334 , n19332 , n19333 );
xor ( n19335 , n19332 , n19333 );
xor ( n19336 , n19243 , n19324 );
and ( n19337 , n18109 , n18624 );
and ( n19338 , n19336 , n19337 );
xor ( n19339 , n19336 , n19337 );
xor ( n19340 , n19247 , n19322 );
and ( n19341 , n18110 , n18624 );
and ( n19342 , n19340 , n19341 );
xor ( n19343 , n19340 , n19341 );
xor ( n19344 , n19251 , n19320 );
and ( n19345 , n18111 , n18624 );
and ( n19346 , n19344 , n19345 );
xor ( n19347 , n19344 , n19345 );
xor ( n19348 , n19255 , n19318 );
and ( n19349 , n18112 , n18624 );
and ( n19350 , n19348 , n19349 );
xor ( n19351 , n19348 , n19349 );
xor ( n19352 , n19259 , n19316 );
and ( n19353 , n18113 , n18624 );
and ( n19354 , n19352 , n19353 );
xor ( n19355 , n19352 , n19353 );
xor ( n19356 , n19263 , n19314 );
and ( n19357 , n18114 , n18624 );
and ( n19358 , n19356 , n19357 );
xor ( n19359 , n19356 , n19357 );
xor ( n19360 , n19267 , n19312 );
and ( n19361 , n18115 , n18624 );
and ( n19362 , n19360 , n19361 );
xor ( n19363 , n19360 , n19361 );
xor ( n19364 , n19271 , n19310 );
and ( n19365 , n18116 , n18624 );
and ( n19366 , n19364 , n19365 );
xor ( n19367 , n19364 , n19365 );
xor ( n19368 , n19275 , n19308 );
and ( n19369 , n18117 , n18624 );
and ( n19370 , n19368 , n19369 );
xor ( n19371 , n19368 , n19369 );
xor ( n19372 , n19279 , n19306 );
and ( n19373 , n18118 , n18624 );
and ( n19374 , n19372 , n19373 );
xor ( n19375 , n19372 , n19373 );
xor ( n19376 , n19283 , n19304 );
and ( n19377 , n18119 , n18624 );
and ( n19378 , n19376 , n19377 );
xor ( n19379 , n19376 , n19377 );
xor ( n19380 , n19287 , n19302 );
and ( n19381 , n18120 , n18624 );
and ( n19382 , n19380 , n19381 );
xor ( n19383 , n19380 , n19381 );
xor ( n19384 , n19291 , n19300 );
and ( n19385 , n18121 , n18624 );
and ( n19386 , n19384 , n19385 );
xor ( n19387 , n19384 , n19385 );
xor ( n19388 , n19295 , n19298 );
and ( n19389 , n18122 , n18624 );
and ( n19390 , n19388 , n19389 );
and ( n19391 , n19387 , n19390 );
or ( n19392 , n19386 , n19391 );
and ( n19393 , n19383 , n19392 );
or ( n19394 , n19382 , n19393 );
and ( n19395 , n19379 , n19394 );
or ( n19396 , n19378 , n19395 );
and ( n19397 , n19375 , n19396 );
or ( n19398 , n19374 , n19397 );
and ( n19399 , n19371 , n19398 );
or ( n19400 , n19370 , n19399 );
and ( n19401 , n19367 , n19400 );
or ( n19402 , n19366 , n19401 );
and ( n19403 , n19363 , n19402 );
or ( n19404 , n19362 , n19403 );
and ( n19405 , n19359 , n19404 );
or ( n19406 , n19358 , n19405 );
and ( n19407 , n19355 , n19406 );
or ( n19408 , n19354 , n19407 );
and ( n19409 , n19351 , n19408 );
or ( n19410 , n19350 , n19409 );
and ( n19411 , n19347 , n19410 );
or ( n19412 , n19346 , n19411 );
and ( n19413 , n19343 , n19412 );
or ( n19414 , n19342 , n19413 );
and ( n19415 , n19339 , n19414 );
or ( n19416 , n19338 , n19415 );
and ( n19417 , n19335 , n19416 );
or ( n19418 , n19334 , n19417 );
and ( n19419 , n19331 , n19418 );
or ( n19420 , n19330 , n19419 );
and ( n19421 , n18107 , n18620 );
and ( n19422 , n19420 , n19421 );
xor ( n19423 , n19420 , n19421 );
xor ( n19424 , n19331 , n19418 );
and ( n19425 , n18108 , n18620 );
and ( n19426 , n19424 , n19425 );
xor ( n19427 , n19424 , n19425 );
xor ( n19428 , n19335 , n19416 );
and ( n19429 , n18109 , n18620 );
and ( n19430 , n19428 , n19429 );
xor ( n19431 , n19428 , n19429 );
xor ( n19432 , n19339 , n19414 );
and ( n19433 , n18110 , n18620 );
and ( n19434 , n19432 , n19433 );
xor ( n19435 , n19432 , n19433 );
xor ( n19436 , n19343 , n19412 );
and ( n19437 , n18111 , n18620 );
and ( n19438 , n19436 , n19437 );
xor ( n19439 , n19436 , n19437 );
xor ( n19440 , n19347 , n19410 );
and ( n19441 , n18112 , n18620 );
and ( n19442 , n19440 , n19441 );
xor ( n19443 , n19440 , n19441 );
xor ( n19444 , n19351 , n19408 );
and ( n19445 , n18113 , n18620 );
and ( n19446 , n19444 , n19445 );
xor ( n19447 , n19444 , n19445 );
xor ( n19448 , n19355 , n19406 );
and ( n19449 , n18114 , n18620 );
and ( n19450 , n19448 , n19449 );
xor ( n19451 , n19448 , n19449 );
xor ( n19452 , n19359 , n19404 );
and ( n19453 , n18115 , n18620 );
and ( n19454 , n19452 , n19453 );
xor ( n19455 , n19452 , n19453 );
xor ( n19456 , n19363 , n19402 );
and ( n19457 , n18116 , n18620 );
and ( n19458 , n19456 , n19457 );
xor ( n19459 , n19456 , n19457 );
xor ( n19460 , n19367 , n19400 );
and ( n19461 , n18117 , n18620 );
and ( n19462 , n19460 , n19461 );
xor ( n19463 , n19460 , n19461 );
xor ( n19464 , n19371 , n19398 );
and ( n19465 , n18118 , n18620 );
and ( n19466 , n19464 , n19465 );
xor ( n19467 , n19464 , n19465 );
xor ( n19468 , n19375 , n19396 );
and ( n19469 , n18119 , n18620 );
and ( n19470 , n19468 , n19469 );
xor ( n19471 , n19468 , n19469 );
xor ( n19472 , n19379 , n19394 );
and ( n19473 , n18120 , n18620 );
and ( n19474 , n19472 , n19473 );
xor ( n19475 , n19472 , n19473 );
xor ( n19476 , n19383 , n19392 );
and ( n19477 , n18121 , n18620 );
and ( n19478 , n19476 , n19477 );
xor ( n19479 , n19476 , n19477 );
xor ( n19480 , n19387 , n19390 );
and ( n19481 , n18122 , n18620 );
and ( n19482 , n19480 , n19481 );
and ( n19483 , n19479 , n19482 );
or ( n19484 , n19478 , n19483 );
and ( n19485 , n19475 , n19484 );
or ( n19486 , n19474 , n19485 );
and ( n19487 , n19471 , n19486 );
or ( n19488 , n19470 , n19487 );
and ( n19489 , n19467 , n19488 );
or ( n19490 , n19466 , n19489 );
and ( n19491 , n19463 , n19490 );
or ( n19492 , n19462 , n19491 );
and ( n19493 , n19459 , n19492 );
or ( n19494 , n19458 , n19493 );
and ( n19495 , n19455 , n19494 );
or ( n19496 , n19454 , n19495 );
and ( n19497 , n19451 , n19496 );
or ( n19498 , n19450 , n19497 );
and ( n19499 , n19447 , n19498 );
or ( n19500 , n19446 , n19499 );
and ( n19501 , n19443 , n19500 );
or ( n19502 , n19442 , n19501 );
and ( n19503 , n19439 , n19502 );
or ( n19504 , n19438 , n19503 );
and ( n19505 , n19435 , n19504 );
or ( n19506 , n19434 , n19505 );
and ( n19507 , n19431 , n19506 );
or ( n19508 , n19430 , n19507 );
and ( n19509 , n19427 , n19508 );
or ( n19510 , n19426 , n19509 );
and ( n19511 , n19423 , n19510 );
or ( n19512 , n19422 , n19511 );
and ( n19513 , n18107 , n18616 );
and ( n19514 , n19512 , n19513 );
xor ( n19515 , n19512 , n19513 );
xor ( n19516 , n19423 , n19510 );
and ( n19517 , n18108 , n18616 );
and ( n19518 , n19516 , n19517 );
xor ( n19519 , n19516 , n19517 );
xor ( n19520 , n19427 , n19508 );
and ( n19521 , n18109 , n18616 );
and ( n19522 , n19520 , n19521 );
xor ( n19523 , n19520 , n19521 );
xor ( n19524 , n19431 , n19506 );
and ( n19525 , n18110 , n18616 );
and ( n19526 , n19524 , n19525 );
xor ( n19527 , n19524 , n19525 );
xor ( n19528 , n19435 , n19504 );
and ( n19529 , n18111 , n18616 );
and ( n19530 , n19528 , n19529 );
xor ( n19531 , n19528 , n19529 );
xor ( n19532 , n19439 , n19502 );
and ( n19533 , n18112 , n18616 );
and ( n19534 , n19532 , n19533 );
xor ( n19535 , n19532 , n19533 );
xor ( n19536 , n19443 , n19500 );
and ( n19537 , n18113 , n18616 );
and ( n19538 , n19536 , n19537 );
xor ( n19539 , n19536 , n19537 );
xor ( n19540 , n19447 , n19498 );
and ( n19541 , n18114 , n18616 );
and ( n19542 , n19540 , n19541 );
xor ( n19543 , n19540 , n19541 );
xor ( n19544 , n19451 , n19496 );
and ( n19545 , n18115 , n18616 );
and ( n19546 , n19544 , n19545 );
xor ( n19547 , n19544 , n19545 );
xor ( n19548 , n19455 , n19494 );
and ( n19549 , n18116 , n18616 );
and ( n19550 , n19548 , n19549 );
xor ( n19551 , n19548 , n19549 );
xor ( n19552 , n19459 , n19492 );
and ( n19553 , n18117 , n18616 );
and ( n19554 , n19552 , n19553 );
xor ( n19555 , n19552 , n19553 );
xor ( n19556 , n19463 , n19490 );
and ( n19557 , n18118 , n18616 );
and ( n19558 , n19556 , n19557 );
xor ( n19559 , n19556 , n19557 );
xor ( n19560 , n19467 , n19488 );
and ( n19561 , n18119 , n18616 );
and ( n19562 , n19560 , n19561 );
xor ( n19563 , n19560 , n19561 );
xor ( n19564 , n19471 , n19486 );
and ( n19565 , n18120 , n18616 );
and ( n19566 , n19564 , n19565 );
xor ( n19567 , n19564 , n19565 );
xor ( n19568 , n19475 , n19484 );
and ( n19569 , n18121 , n18616 );
and ( n19570 , n19568 , n19569 );
xor ( n19571 , n19568 , n19569 );
xor ( n19572 , n19479 , n19482 );
and ( n19573 , n18122 , n18616 );
and ( n19574 , n19572 , n19573 );
and ( n19575 , n19571 , n19574 );
or ( n19576 , n19570 , n19575 );
and ( n19577 , n19567 , n19576 );
or ( n19578 , n19566 , n19577 );
and ( n19579 , n19563 , n19578 );
or ( n19580 , n19562 , n19579 );
and ( n19581 , n19559 , n19580 );
or ( n19582 , n19558 , n19581 );
and ( n19583 , n19555 , n19582 );
or ( n19584 , n19554 , n19583 );
and ( n19585 , n19551 , n19584 );
or ( n19586 , n19550 , n19585 );
and ( n19587 , n19547 , n19586 );
or ( n19588 , n19546 , n19587 );
and ( n19589 , n19543 , n19588 );
or ( n19590 , n19542 , n19589 );
and ( n19591 , n19539 , n19590 );
or ( n19592 , n19538 , n19591 );
and ( n19593 , n19535 , n19592 );
or ( n19594 , n19534 , n19593 );
and ( n19595 , n19531 , n19594 );
or ( n19596 , n19530 , n19595 );
and ( n19597 , n19527 , n19596 );
or ( n19598 , n19526 , n19597 );
and ( n19599 , n19523 , n19598 );
or ( n19600 , n19522 , n19599 );
and ( n19601 , n19519 , n19600 );
or ( n19602 , n19518 , n19601 );
and ( n19603 , n19515 , n19602 );
or ( n19604 , n19514 , n19603 );
and ( n19605 , n18107 , n18612 );
and ( n19606 , n19604 , n19605 );
xor ( n19607 , n19604 , n19605 );
xor ( n19608 , n19515 , n19602 );
and ( n19609 , n18108 , n18612 );
and ( n19610 , n19608 , n19609 );
xor ( n19611 , n19608 , n19609 );
xor ( n19612 , n19519 , n19600 );
and ( n19613 , n18109 , n18612 );
and ( n19614 , n19612 , n19613 );
xor ( n19615 , n19612 , n19613 );
xor ( n19616 , n19523 , n19598 );
and ( n19617 , n18110 , n18612 );
and ( n19618 , n19616 , n19617 );
xor ( n19619 , n19616 , n19617 );
xor ( n19620 , n19527 , n19596 );
and ( n19621 , n18111 , n18612 );
and ( n19622 , n19620 , n19621 );
xor ( n19623 , n19620 , n19621 );
xor ( n19624 , n19531 , n19594 );
and ( n19625 , n18112 , n18612 );
and ( n19626 , n19624 , n19625 );
xor ( n19627 , n19624 , n19625 );
xor ( n19628 , n19535 , n19592 );
and ( n19629 , n18113 , n18612 );
and ( n19630 , n19628 , n19629 );
xor ( n19631 , n19628 , n19629 );
xor ( n19632 , n19539 , n19590 );
and ( n19633 , n18114 , n18612 );
and ( n19634 , n19632 , n19633 );
xor ( n19635 , n19632 , n19633 );
xor ( n19636 , n19543 , n19588 );
and ( n19637 , n18115 , n18612 );
and ( n19638 , n19636 , n19637 );
xor ( n19639 , n19636 , n19637 );
xor ( n19640 , n19547 , n19586 );
and ( n19641 , n18116 , n18612 );
and ( n19642 , n19640 , n19641 );
xor ( n19643 , n19640 , n19641 );
xor ( n19644 , n19551 , n19584 );
and ( n19645 , n18117 , n18612 );
and ( n19646 , n19644 , n19645 );
xor ( n19647 , n19644 , n19645 );
xor ( n19648 , n19555 , n19582 );
and ( n19649 , n18118 , n18612 );
and ( n19650 , n19648 , n19649 );
xor ( n19651 , n19648 , n19649 );
xor ( n19652 , n19559 , n19580 );
and ( n19653 , n18119 , n18612 );
and ( n19654 , n19652 , n19653 );
xor ( n19655 , n19652 , n19653 );
xor ( n19656 , n19563 , n19578 );
and ( n19657 , n18120 , n18612 );
and ( n19658 , n19656 , n19657 );
xor ( n19659 , n19656 , n19657 );
xor ( n19660 , n19567 , n19576 );
and ( n19661 , n18121 , n18612 );
and ( n19662 , n19660 , n19661 );
xor ( n19663 , n19660 , n19661 );
xor ( n19664 , n19571 , n19574 );
and ( n19665 , n18122 , n18612 );
and ( n19666 , n19664 , n19665 );
and ( n19667 , n19663 , n19666 );
or ( n19668 , n19662 , n19667 );
and ( n19669 , n19659 , n19668 );
or ( n19670 , n19658 , n19669 );
and ( n19671 , n19655 , n19670 );
or ( n19672 , n19654 , n19671 );
and ( n19673 , n19651 , n19672 );
or ( n19674 , n19650 , n19673 );
and ( n19675 , n19647 , n19674 );
or ( n19676 , n19646 , n19675 );
and ( n19677 , n19643 , n19676 );
or ( n19678 , n19642 , n19677 );
and ( n19679 , n19639 , n19678 );
or ( n19680 , n19638 , n19679 );
and ( n19681 , n19635 , n19680 );
or ( n19682 , n19634 , n19681 );
and ( n19683 , n19631 , n19682 );
or ( n19684 , n19630 , n19683 );
and ( n19685 , n19627 , n19684 );
or ( n19686 , n19626 , n19685 );
and ( n19687 , n19623 , n19686 );
or ( n19688 , n19622 , n19687 );
and ( n19689 , n19619 , n19688 );
or ( n19690 , n19618 , n19689 );
and ( n19691 , n19615 , n19690 );
or ( n19692 , n19614 , n19691 );
and ( n19693 , n19611 , n19692 );
or ( n19694 , n19610 , n19693 );
and ( n19695 , n19607 , n19694 );
or ( n19696 , n19606 , n19695 );
and ( n19697 , n18107 , n18608 );
and ( n19698 , n19696 , n19697 );
xor ( n19699 , n19696 , n19697 );
xor ( n19700 , n19607 , n19694 );
and ( n19701 , n18108 , n18608 );
and ( n19702 , n19700 , n19701 );
xor ( n19703 , n19700 , n19701 );
xor ( n19704 , n19611 , n19692 );
and ( n19705 , n18109 , n18608 );
and ( n19706 , n19704 , n19705 );
xor ( n19707 , n19704 , n19705 );
xor ( n19708 , n19615 , n19690 );
and ( n19709 , n18110 , n18608 );
and ( n19710 , n19708 , n19709 );
xor ( n19711 , n19708 , n19709 );
xor ( n19712 , n19619 , n19688 );
and ( n19713 , n18111 , n18608 );
and ( n19714 , n19712 , n19713 );
xor ( n19715 , n19712 , n19713 );
xor ( n19716 , n19623 , n19686 );
and ( n19717 , n18112 , n18608 );
and ( n19718 , n19716 , n19717 );
xor ( n19719 , n19716 , n19717 );
xor ( n19720 , n19627 , n19684 );
and ( n19721 , n18113 , n18608 );
and ( n19722 , n19720 , n19721 );
xor ( n19723 , n19720 , n19721 );
xor ( n19724 , n19631 , n19682 );
and ( n19725 , n18114 , n18608 );
and ( n19726 , n19724 , n19725 );
xor ( n19727 , n19724 , n19725 );
xor ( n19728 , n19635 , n19680 );
and ( n19729 , n18115 , n18608 );
and ( n19730 , n19728 , n19729 );
xor ( n19731 , n19728 , n19729 );
xor ( n19732 , n19639 , n19678 );
and ( n19733 , n18116 , n18608 );
and ( n19734 , n19732 , n19733 );
xor ( n19735 , n19732 , n19733 );
xor ( n19736 , n19643 , n19676 );
and ( n19737 , n18117 , n18608 );
and ( n19738 , n19736 , n19737 );
xor ( n19739 , n19736 , n19737 );
xor ( n19740 , n19647 , n19674 );
and ( n19741 , n18118 , n18608 );
and ( n19742 , n19740 , n19741 );
xor ( n19743 , n19740 , n19741 );
xor ( n19744 , n19651 , n19672 );
and ( n19745 , n18119 , n18608 );
and ( n19746 , n19744 , n19745 );
xor ( n19747 , n19744 , n19745 );
xor ( n19748 , n19655 , n19670 );
and ( n19749 , n18120 , n18608 );
and ( n19750 , n19748 , n19749 );
xor ( n19751 , n19748 , n19749 );
xor ( n19752 , n19659 , n19668 );
and ( n19753 , n18121 , n18608 );
and ( n19754 , n19752 , n19753 );
xor ( n19755 , n19752 , n19753 );
xor ( n19756 , n19663 , n19666 );
and ( n19757 , n18122 , n18608 );
and ( n19758 , n19756 , n19757 );
and ( n19759 , n19755 , n19758 );
or ( n19760 , n19754 , n19759 );
and ( n19761 , n19751 , n19760 );
or ( n19762 , n19750 , n19761 );
and ( n19763 , n19747 , n19762 );
or ( n19764 , n19746 , n19763 );
and ( n19765 , n19743 , n19764 );
or ( n19766 , n19742 , n19765 );
and ( n19767 , n19739 , n19766 );
or ( n19768 , n19738 , n19767 );
and ( n19769 , n19735 , n19768 );
or ( n19770 , n19734 , n19769 );
and ( n19771 , n19731 , n19770 );
or ( n19772 , n19730 , n19771 );
and ( n19773 , n19727 , n19772 );
or ( n19774 , n19726 , n19773 );
and ( n19775 , n19723 , n19774 );
or ( n19776 , n19722 , n19775 );
and ( n19777 , n19719 , n19776 );
or ( n19778 , n19718 , n19777 );
and ( n19779 , n19715 , n19778 );
or ( n19780 , n19714 , n19779 );
and ( n19781 , n19711 , n19780 );
or ( n19782 , n19710 , n19781 );
and ( n19783 , n19707 , n19782 );
or ( n19784 , n19706 , n19783 );
and ( n19785 , n19703 , n19784 );
or ( n19786 , n19702 , n19785 );
and ( n19787 , n19699 , n19786 );
or ( n19788 , n19698 , n19787 );
and ( n19789 , n18107 , n18604 );
and ( n19790 , n19788 , n19789 );
xor ( n19791 , n19788 , n19789 );
xor ( n19792 , n19699 , n19786 );
and ( n19793 , n18108 , n18604 );
and ( n19794 , n19792 , n19793 );
xor ( n19795 , n19792 , n19793 );
xor ( n19796 , n19703 , n19784 );
and ( n19797 , n18109 , n18604 );
and ( n19798 , n19796 , n19797 );
xor ( n19799 , n19796 , n19797 );
xor ( n19800 , n19707 , n19782 );
and ( n19801 , n18110 , n18604 );
and ( n19802 , n19800 , n19801 );
xor ( n19803 , n19800 , n19801 );
xor ( n19804 , n19711 , n19780 );
and ( n19805 , n18111 , n18604 );
and ( n19806 , n19804 , n19805 );
xor ( n19807 , n19804 , n19805 );
xor ( n19808 , n19715 , n19778 );
and ( n19809 , n18112 , n18604 );
and ( n19810 , n19808 , n19809 );
xor ( n19811 , n19808 , n19809 );
xor ( n19812 , n19719 , n19776 );
and ( n19813 , n18113 , n18604 );
and ( n19814 , n19812 , n19813 );
xor ( n19815 , n19812 , n19813 );
xor ( n19816 , n19723 , n19774 );
and ( n19817 , n18114 , n18604 );
and ( n19818 , n19816 , n19817 );
xor ( n19819 , n19816 , n19817 );
xor ( n19820 , n19727 , n19772 );
and ( n19821 , n18115 , n18604 );
and ( n19822 , n19820 , n19821 );
xor ( n19823 , n19820 , n19821 );
xor ( n19824 , n19731 , n19770 );
and ( n19825 , n18116 , n18604 );
and ( n19826 , n19824 , n19825 );
xor ( n19827 , n19824 , n19825 );
xor ( n19828 , n19735 , n19768 );
and ( n19829 , n18117 , n18604 );
and ( n19830 , n19828 , n19829 );
xor ( n19831 , n19828 , n19829 );
xor ( n19832 , n19739 , n19766 );
and ( n19833 , n18118 , n18604 );
and ( n19834 , n19832 , n19833 );
xor ( n19835 , n19832 , n19833 );
xor ( n19836 , n19743 , n19764 );
and ( n19837 , n18119 , n18604 );
and ( n19838 , n19836 , n19837 );
xor ( n19839 , n19836 , n19837 );
xor ( n19840 , n19747 , n19762 );
and ( n19841 , n18120 , n18604 );
and ( n19842 , n19840 , n19841 );
xor ( n19843 , n19840 , n19841 );
xor ( n19844 , n19751 , n19760 );
and ( n19845 , n18121 , n18604 );
and ( n19846 , n19844 , n19845 );
xor ( n19847 , n19844 , n19845 );
xor ( n19848 , n19755 , n19758 );
and ( n19849 , n18122 , n18604 );
and ( n19850 , n19848 , n19849 );
and ( n19851 , n19847 , n19850 );
or ( n19852 , n19846 , n19851 );
and ( n19853 , n19843 , n19852 );
or ( n19854 , n19842 , n19853 );
and ( n19855 , n19839 , n19854 );
or ( n19856 , n19838 , n19855 );
and ( n19857 , n19835 , n19856 );
or ( n19858 , n19834 , n19857 );
and ( n19859 , n19831 , n19858 );
or ( n19860 , n19830 , n19859 );
and ( n19861 , n19827 , n19860 );
or ( n19862 , n19826 , n19861 );
and ( n19863 , n19823 , n19862 );
or ( n19864 , n19822 , n19863 );
and ( n19865 , n19819 , n19864 );
or ( n19866 , n19818 , n19865 );
and ( n19867 , n19815 , n19866 );
or ( n19868 , n19814 , n19867 );
and ( n19869 , n19811 , n19868 );
or ( n19870 , n19810 , n19869 );
and ( n19871 , n19807 , n19870 );
or ( n19872 , n19806 , n19871 );
and ( n19873 , n19803 , n19872 );
or ( n19874 , n19802 , n19873 );
and ( n19875 , n19799 , n19874 );
or ( n19876 , n19798 , n19875 );
and ( n19877 , n19795 , n19876 );
or ( n19878 , n19794 , n19877 );
and ( n19879 , n19791 , n19878 );
or ( n19880 , n19790 , n19879 );
and ( n19881 , n18107 , n18600 );
and ( n19882 , n19880 , n19881 );
xor ( n19883 , n19880 , n19881 );
xor ( n19884 , n19791 , n19878 );
and ( n19885 , n18108 , n18600 );
and ( n19886 , n19884 , n19885 );
xor ( n19887 , n19884 , n19885 );
xor ( n19888 , n19795 , n19876 );
and ( n19889 , n18109 , n18600 );
and ( n19890 , n19888 , n19889 );
xor ( n19891 , n19888 , n19889 );
xor ( n19892 , n19799 , n19874 );
and ( n19893 , n18110 , n18600 );
and ( n19894 , n19892 , n19893 );
xor ( n19895 , n19892 , n19893 );
xor ( n19896 , n19803 , n19872 );
and ( n19897 , n18111 , n18600 );
and ( n19898 , n19896 , n19897 );
xor ( n19899 , n19896 , n19897 );
xor ( n19900 , n19807 , n19870 );
and ( n19901 , n18112 , n18600 );
and ( n19902 , n19900 , n19901 );
xor ( n19903 , n19900 , n19901 );
xor ( n19904 , n19811 , n19868 );
and ( n19905 , n18113 , n18600 );
and ( n19906 , n19904 , n19905 );
xor ( n19907 , n19904 , n19905 );
xor ( n19908 , n19815 , n19866 );
and ( n19909 , n18114 , n18600 );
and ( n19910 , n19908 , n19909 );
xor ( n19911 , n19908 , n19909 );
xor ( n19912 , n19819 , n19864 );
and ( n19913 , n18115 , n18600 );
and ( n19914 , n19912 , n19913 );
xor ( n19915 , n19912 , n19913 );
xor ( n19916 , n19823 , n19862 );
and ( n19917 , n18116 , n18600 );
and ( n19918 , n19916 , n19917 );
xor ( n19919 , n19916 , n19917 );
xor ( n19920 , n19827 , n19860 );
and ( n19921 , n18117 , n18600 );
and ( n19922 , n19920 , n19921 );
xor ( n19923 , n19920 , n19921 );
xor ( n19924 , n19831 , n19858 );
and ( n19925 , n18118 , n18600 );
and ( n19926 , n19924 , n19925 );
xor ( n19927 , n19924 , n19925 );
xor ( n19928 , n19835 , n19856 );
and ( n19929 , n18119 , n18600 );
and ( n19930 , n19928 , n19929 );
xor ( n19931 , n19928 , n19929 );
xor ( n19932 , n19839 , n19854 );
and ( n19933 , n18120 , n18600 );
and ( n19934 , n19932 , n19933 );
xor ( n19935 , n19932 , n19933 );
xor ( n19936 , n19843 , n19852 );
and ( n19937 , n18121 , n18600 );
and ( n19938 , n19936 , n19937 );
xor ( n19939 , n19936 , n19937 );
xor ( n19940 , n19847 , n19850 );
and ( n19941 , n18122 , n18600 );
and ( n19942 , n19940 , n19941 );
and ( n19943 , n19939 , n19942 );
or ( n19944 , n19938 , n19943 );
and ( n19945 , n19935 , n19944 );
or ( n19946 , n19934 , n19945 );
and ( n19947 , n19931 , n19946 );
or ( n19948 , n19930 , n19947 );
and ( n19949 , n19927 , n19948 );
or ( n19950 , n19926 , n19949 );
and ( n19951 , n19923 , n19950 );
or ( n19952 , n19922 , n19951 );
and ( n19953 , n19919 , n19952 );
or ( n19954 , n19918 , n19953 );
and ( n19955 , n19915 , n19954 );
or ( n19956 , n19914 , n19955 );
and ( n19957 , n19911 , n19956 );
or ( n19958 , n19910 , n19957 );
and ( n19959 , n19907 , n19958 );
or ( n19960 , n19906 , n19959 );
and ( n19961 , n19903 , n19960 );
or ( n19962 , n19902 , n19961 );
and ( n19963 , n19899 , n19962 );
or ( n19964 , n19898 , n19963 );
and ( n19965 , n19895 , n19964 );
or ( n19966 , n19894 , n19965 );
and ( n19967 , n19891 , n19966 );
or ( n19968 , n19890 , n19967 );
and ( n19969 , n19887 , n19968 );
or ( n19970 , n19886 , n19969 );
and ( n19971 , n19883 , n19970 );
or ( n19972 , n19882 , n19971 );
and ( n19973 , n18107 , n18596 );
and ( n19974 , n19972 , n19973 );
xor ( n19975 , n19972 , n19973 );
xor ( n19976 , n19883 , n19970 );
and ( n19977 , n18108 , n18596 );
and ( n19978 , n19976 , n19977 );
xor ( n19979 , n19976 , n19977 );
xor ( n19980 , n19887 , n19968 );
and ( n19981 , n18109 , n18596 );
and ( n19982 , n19980 , n19981 );
xor ( n19983 , n19980 , n19981 );
xor ( n19984 , n19891 , n19966 );
and ( n19985 , n18110 , n18596 );
and ( n19986 , n19984 , n19985 );
xor ( n19987 , n19984 , n19985 );
xor ( n19988 , n19895 , n19964 );
and ( n19989 , n18111 , n18596 );
and ( n19990 , n19988 , n19989 );
xor ( n19991 , n19988 , n19989 );
xor ( n19992 , n19899 , n19962 );
and ( n19993 , n18112 , n18596 );
and ( n19994 , n19992 , n19993 );
xor ( n19995 , n19992 , n19993 );
xor ( n19996 , n19903 , n19960 );
and ( n19997 , n18113 , n18596 );
and ( n19998 , n19996 , n19997 );
xor ( n19999 , n19996 , n19997 );
xor ( n20000 , n19907 , n19958 );
and ( n20001 , n18114 , n18596 );
and ( n20002 , n20000 , n20001 );
xor ( n20003 , n20000 , n20001 );
xor ( n20004 , n19911 , n19956 );
and ( n20005 , n18115 , n18596 );
and ( n20006 , n20004 , n20005 );
xor ( n20007 , n20004 , n20005 );
xor ( n20008 , n19915 , n19954 );
and ( n20009 , n18116 , n18596 );
and ( n20010 , n20008 , n20009 );
xor ( n20011 , n20008 , n20009 );
xor ( n20012 , n19919 , n19952 );
and ( n20013 , n18117 , n18596 );
and ( n20014 , n20012 , n20013 );
xor ( n20015 , n20012 , n20013 );
xor ( n20016 , n19923 , n19950 );
and ( n20017 , n18118 , n18596 );
and ( n20018 , n20016 , n20017 );
xor ( n20019 , n20016 , n20017 );
xor ( n20020 , n19927 , n19948 );
and ( n20021 , n18119 , n18596 );
and ( n20022 , n20020 , n20021 );
xor ( n20023 , n20020 , n20021 );
xor ( n20024 , n19931 , n19946 );
and ( n20025 , n18120 , n18596 );
and ( n20026 , n20024 , n20025 );
xor ( n20027 , n20024 , n20025 );
xor ( n20028 , n19935 , n19944 );
and ( n20029 , n18121 , n18596 );
and ( n20030 , n20028 , n20029 );
xor ( n20031 , n20028 , n20029 );
xor ( n20032 , n19939 , n19942 );
and ( n20033 , n18122 , n18596 );
and ( n20034 , n20032 , n20033 );
and ( n20035 , n20031 , n20034 );
or ( n20036 , n20030 , n20035 );
and ( n20037 , n20027 , n20036 );
or ( n20038 , n20026 , n20037 );
and ( n20039 , n20023 , n20038 );
or ( n20040 , n20022 , n20039 );
and ( n20041 , n20019 , n20040 );
or ( n20042 , n20018 , n20041 );
and ( n20043 , n20015 , n20042 );
or ( n20044 , n20014 , n20043 );
and ( n20045 , n20011 , n20044 );
or ( n20046 , n20010 , n20045 );
and ( n20047 , n20007 , n20046 );
or ( n20048 , n20006 , n20047 );
and ( n20049 , n20003 , n20048 );
or ( n20050 , n20002 , n20049 );
and ( n20051 , n19999 , n20050 );
or ( n20052 , n19998 , n20051 );
and ( n20053 , n19995 , n20052 );
or ( n20054 , n19994 , n20053 );
and ( n20055 , n19991 , n20054 );
or ( n20056 , n19990 , n20055 );
and ( n20057 , n19987 , n20056 );
or ( n20058 , n19986 , n20057 );
and ( n20059 , n19983 , n20058 );
or ( n20060 , n19982 , n20059 );
and ( n20061 , n19979 , n20060 );
or ( n20062 , n19978 , n20061 );
and ( n20063 , n19975 , n20062 );
or ( n20064 , n19974 , n20063 );
and ( n20065 , n18107 , n18592 );
and ( n20066 , n20064 , n20065 );
xor ( n20067 , n20064 , n20065 );
xor ( n20068 , n19975 , n20062 );
and ( n20069 , n18108 , n18592 );
and ( n20070 , n20068 , n20069 );
xor ( n20071 , n20068 , n20069 );
xor ( n20072 , n19979 , n20060 );
and ( n20073 , n18109 , n18592 );
and ( n20074 , n20072 , n20073 );
xor ( n20075 , n20072 , n20073 );
xor ( n20076 , n19983 , n20058 );
and ( n20077 , n18110 , n18592 );
and ( n20078 , n20076 , n20077 );
xor ( n20079 , n20076 , n20077 );
xor ( n20080 , n19987 , n20056 );
and ( n20081 , n18111 , n18592 );
and ( n20082 , n20080 , n20081 );
xor ( n20083 , n20080 , n20081 );
xor ( n20084 , n19991 , n20054 );
and ( n20085 , n18112 , n18592 );
and ( n20086 , n20084 , n20085 );
xor ( n20087 , n20084 , n20085 );
xor ( n20088 , n19995 , n20052 );
and ( n20089 , n18113 , n18592 );
and ( n20090 , n20088 , n20089 );
xor ( n20091 , n20088 , n20089 );
xor ( n20092 , n19999 , n20050 );
and ( n20093 , n18114 , n18592 );
and ( n20094 , n20092 , n20093 );
xor ( n20095 , n20092 , n20093 );
xor ( n20096 , n20003 , n20048 );
and ( n20097 , n18115 , n18592 );
and ( n20098 , n20096 , n20097 );
xor ( n20099 , n20096 , n20097 );
xor ( n20100 , n20007 , n20046 );
and ( n20101 , n18116 , n18592 );
and ( n20102 , n20100 , n20101 );
xor ( n20103 , n20100 , n20101 );
xor ( n20104 , n20011 , n20044 );
and ( n20105 , n18117 , n18592 );
and ( n20106 , n20104 , n20105 );
xor ( n20107 , n20104 , n20105 );
xor ( n20108 , n20015 , n20042 );
and ( n20109 , n18118 , n18592 );
and ( n20110 , n20108 , n20109 );
xor ( n20111 , n20108 , n20109 );
xor ( n20112 , n20019 , n20040 );
and ( n20113 , n18119 , n18592 );
and ( n20114 , n20112 , n20113 );
xor ( n20115 , n20112 , n20113 );
xor ( n20116 , n20023 , n20038 );
and ( n20117 , n18120 , n18592 );
and ( n20118 , n20116 , n20117 );
xor ( n20119 , n20116 , n20117 );
xor ( n20120 , n20027 , n20036 );
and ( n20121 , n18121 , n18592 );
and ( n20122 , n20120 , n20121 );
xor ( n20123 , n20120 , n20121 );
xor ( n20124 , n20031 , n20034 );
and ( n20125 , n18122 , n18592 );
and ( n20126 , n20124 , n20125 );
and ( n20127 , n20123 , n20126 );
or ( n20128 , n20122 , n20127 );
and ( n20129 , n20119 , n20128 );
or ( n20130 , n20118 , n20129 );
and ( n20131 , n20115 , n20130 );
or ( n20132 , n20114 , n20131 );
and ( n20133 , n20111 , n20132 );
or ( n20134 , n20110 , n20133 );
and ( n20135 , n20107 , n20134 );
or ( n20136 , n20106 , n20135 );
and ( n20137 , n20103 , n20136 );
or ( n20138 , n20102 , n20137 );
and ( n20139 , n20099 , n20138 );
or ( n20140 , n20098 , n20139 );
and ( n20141 , n20095 , n20140 );
or ( n20142 , n20094 , n20141 );
and ( n20143 , n20091 , n20142 );
or ( n20144 , n20090 , n20143 );
and ( n20145 , n20087 , n20144 );
or ( n20146 , n20086 , n20145 );
and ( n20147 , n20083 , n20146 );
or ( n20148 , n20082 , n20147 );
and ( n20149 , n20079 , n20148 );
or ( n20150 , n20078 , n20149 );
and ( n20151 , n20075 , n20150 );
or ( n20152 , n20074 , n20151 );
and ( n20153 , n20071 , n20152 );
or ( n20154 , n20070 , n20153 );
and ( n20155 , n20067 , n20154 );
or ( n20156 , n20066 , n20155 );
and ( n20157 , n18107 , n18588 );
and ( n20158 , n20156 , n20157 );
xor ( n20159 , n20156 , n20157 );
xor ( n20160 , n20067 , n20154 );
and ( n20161 , n18108 , n18588 );
and ( n20162 , n20160 , n20161 );
xor ( n20163 , n20160 , n20161 );
xor ( n20164 , n20071 , n20152 );
and ( n20165 , n18109 , n18588 );
and ( n20166 , n20164 , n20165 );
xor ( n20167 , n20164 , n20165 );
xor ( n20168 , n20075 , n20150 );
and ( n20169 , n18110 , n18588 );
and ( n20170 , n20168 , n20169 );
xor ( n20171 , n20168 , n20169 );
xor ( n20172 , n20079 , n20148 );
and ( n20173 , n18111 , n18588 );
and ( n20174 , n20172 , n20173 );
xor ( n20175 , n20172 , n20173 );
xor ( n20176 , n20083 , n20146 );
and ( n20177 , n18112 , n18588 );
and ( n20178 , n20176 , n20177 );
xor ( n20179 , n20176 , n20177 );
xor ( n20180 , n20087 , n20144 );
and ( n20181 , n18113 , n18588 );
and ( n20182 , n20180 , n20181 );
xor ( n20183 , n20180 , n20181 );
xor ( n20184 , n20091 , n20142 );
and ( n20185 , n18114 , n18588 );
and ( n20186 , n20184 , n20185 );
xor ( n20187 , n20184 , n20185 );
xor ( n20188 , n20095 , n20140 );
and ( n20189 , n18115 , n18588 );
and ( n20190 , n20188 , n20189 );
xor ( n20191 , n20188 , n20189 );
xor ( n20192 , n20099 , n20138 );
and ( n20193 , n18116 , n18588 );
and ( n20194 , n20192 , n20193 );
xor ( n20195 , n20192 , n20193 );
xor ( n20196 , n20103 , n20136 );
and ( n20197 , n18117 , n18588 );
and ( n20198 , n20196 , n20197 );
xor ( n20199 , n20196 , n20197 );
xor ( n20200 , n20107 , n20134 );
and ( n20201 , n18118 , n18588 );
and ( n20202 , n20200 , n20201 );
xor ( n20203 , n20200 , n20201 );
xor ( n20204 , n20111 , n20132 );
and ( n20205 , n18119 , n18588 );
and ( n20206 , n20204 , n20205 );
xor ( n20207 , n20204 , n20205 );
xor ( n20208 , n20115 , n20130 );
and ( n20209 , n18120 , n18588 );
and ( n20210 , n20208 , n20209 );
xor ( n20211 , n20208 , n20209 );
xor ( n20212 , n20119 , n20128 );
and ( n20213 , n18121 , n18588 );
and ( n20214 , n20212 , n20213 );
xor ( n20215 , n20212 , n20213 );
xor ( n20216 , n20123 , n20126 );
and ( n20217 , n18122 , n18588 );
and ( n20218 , n20216 , n20217 );
and ( n20219 , n20215 , n20218 );
or ( n20220 , n20214 , n20219 );
and ( n20221 , n20211 , n20220 );
or ( n20222 , n20210 , n20221 );
and ( n20223 , n20207 , n20222 );
or ( n20224 , n20206 , n20223 );
and ( n20225 , n20203 , n20224 );
or ( n20226 , n20202 , n20225 );
and ( n20227 , n20199 , n20226 );
or ( n20228 , n20198 , n20227 );
and ( n20229 , n20195 , n20228 );
or ( n20230 , n20194 , n20229 );
and ( n20231 , n20191 , n20230 );
or ( n20232 , n20190 , n20231 );
and ( n20233 , n20187 , n20232 );
or ( n20234 , n20186 , n20233 );
and ( n20235 , n20183 , n20234 );
or ( n20236 , n20182 , n20235 );
and ( n20237 , n20179 , n20236 );
or ( n20238 , n20178 , n20237 );
and ( n20239 , n20175 , n20238 );
or ( n20240 , n20174 , n20239 );
and ( n20241 , n20171 , n20240 );
or ( n20242 , n20170 , n20241 );
and ( n20243 , n20167 , n20242 );
or ( n20244 , n20166 , n20243 );
and ( n20245 , n20163 , n20244 );
or ( n20246 , n20162 , n20245 );
and ( n20247 , n20159 , n20246 );
or ( n20248 , n20158 , n20247 );
and ( n20249 , n18107 , n18584 );
and ( n20250 , n20248 , n20249 );
xor ( n20251 , n20248 , n20249 );
xor ( n20252 , n20159 , n20246 );
and ( n20253 , n18108 , n18584 );
and ( n20254 , n20252 , n20253 );
xor ( n20255 , n20252 , n20253 );
xor ( n20256 , n20163 , n20244 );
and ( n20257 , n18109 , n18584 );
and ( n20258 , n20256 , n20257 );
xor ( n20259 , n20256 , n20257 );
xor ( n20260 , n20167 , n20242 );
and ( n20261 , n18110 , n18584 );
and ( n20262 , n20260 , n20261 );
xor ( n20263 , n20260 , n20261 );
xor ( n20264 , n20171 , n20240 );
and ( n20265 , n18111 , n18584 );
and ( n20266 , n20264 , n20265 );
xor ( n20267 , n20264 , n20265 );
xor ( n20268 , n20175 , n20238 );
and ( n20269 , n18112 , n18584 );
and ( n20270 , n20268 , n20269 );
xor ( n20271 , n20268 , n20269 );
xor ( n20272 , n20179 , n20236 );
and ( n20273 , n18113 , n18584 );
and ( n20274 , n20272 , n20273 );
xor ( n20275 , n20272 , n20273 );
xor ( n20276 , n20183 , n20234 );
and ( n20277 , n18114 , n18584 );
and ( n20278 , n20276 , n20277 );
xor ( n20279 , n20276 , n20277 );
xor ( n20280 , n20187 , n20232 );
and ( n20281 , n18115 , n18584 );
and ( n20282 , n20280 , n20281 );
xor ( n20283 , n20280 , n20281 );
xor ( n20284 , n20191 , n20230 );
and ( n20285 , n18116 , n18584 );
and ( n20286 , n20284 , n20285 );
xor ( n20287 , n20284 , n20285 );
xor ( n20288 , n20195 , n20228 );
and ( n20289 , n18117 , n18584 );
and ( n20290 , n20288 , n20289 );
xor ( n20291 , n20288 , n20289 );
xor ( n20292 , n20199 , n20226 );
and ( n20293 , n18118 , n18584 );
and ( n20294 , n20292 , n20293 );
xor ( n20295 , n20292 , n20293 );
xor ( n20296 , n20203 , n20224 );
and ( n20297 , n18119 , n18584 );
and ( n20298 , n20296 , n20297 );
xor ( n20299 , n20296 , n20297 );
xor ( n20300 , n20207 , n20222 );
and ( n20301 , n18120 , n18584 );
and ( n20302 , n20300 , n20301 );
xor ( n20303 , n20300 , n20301 );
xor ( n20304 , n20211 , n20220 );
and ( n20305 , n18121 , n18584 );
and ( n20306 , n20304 , n20305 );
xor ( n20307 , n20304 , n20305 );
xor ( n20308 , n20215 , n20218 );
and ( n20309 , n18122 , n18584 );
and ( n20310 , n20308 , n20309 );
and ( n20311 , n20307 , n20310 );
or ( n20312 , n20306 , n20311 );
and ( n20313 , n20303 , n20312 );
or ( n20314 , n20302 , n20313 );
and ( n20315 , n20299 , n20314 );
or ( n20316 , n20298 , n20315 );
and ( n20317 , n20295 , n20316 );
or ( n20318 , n20294 , n20317 );
and ( n20319 , n20291 , n20318 );
or ( n20320 , n20290 , n20319 );
and ( n20321 , n20287 , n20320 );
or ( n20322 , n20286 , n20321 );
and ( n20323 , n20283 , n20322 );
or ( n20324 , n20282 , n20323 );
and ( n20325 , n20279 , n20324 );
or ( n20326 , n20278 , n20325 );
and ( n20327 , n20275 , n20326 );
or ( n20328 , n20274 , n20327 );
and ( n20329 , n20271 , n20328 );
or ( n20330 , n20270 , n20329 );
and ( n20331 , n20267 , n20330 );
or ( n20332 , n20266 , n20331 );
and ( n20333 , n20263 , n20332 );
or ( n20334 , n20262 , n20333 );
and ( n20335 , n20259 , n20334 );
or ( n20336 , n20258 , n20335 );
and ( n20337 , n20255 , n20336 );
or ( n20338 , n20254 , n20337 );
and ( n20339 , n20251 , n20338 );
or ( n20340 , n20250 , n20339 );
and ( n20341 , n18107 , n18580 );
and ( n20342 , n20340 , n20341 );
xor ( n20343 , n20340 , n20341 );
xor ( n20344 , n20251 , n20338 );
and ( n20345 , n18108 , n18580 );
and ( n20346 , n20344 , n20345 );
xor ( n20347 , n20344 , n20345 );
xor ( n20348 , n20255 , n20336 );
and ( n20349 , n18109 , n18580 );
and ( n20350 , n20348 , n20349 );
xor ( n20351 , n20348 , n20349 );
xor ( n20352 , n20259 , n20334 );
and ( n20353 , n18110 , n18580 );
and ( n20354 , n20352 , n20353 );
xor ( n20355 , n20352 , n20353 );
xor ( n20356 , n20263 , n20332 );
and ( n20357 , n18111 , n18580 );
and ( n20358 , n20356 , n20357 );
xor ( n20359 , n20356 , n20357 );
xor ( n20360 , n20267 , n20330 );
and ( n20361 , n18112 , n18580 );
and ( n20362 , n20360 , n20361 );
xor ( n20363 , n20360 , n20361 );
xor ( n20364 , n20271 , n20328 );
and ( n20365 , n18113 , n18580 );
and ( n20366 , n20364 , n20365 );
xor ( n20367 , n20364 , n20365 );
xor ( n20368 , n20275 , n20326 );
and ( n20369 , n18114 , n18580 );
and ( n20370 , n20368 , n20369 );
xor ( n20371 , n20368 , n20369 );
xor ( n20372 , n20279 , n20324 );
and ( n20373 , n18115 , n18580 );
and ( n20374 , n20372 , n20373 );
xor ( n20375 , n20372 , n20373 );
xor ( n20376 , n20283 , n20322 );
and ( n20377 , n18116 , n18580 );
and ( n20378 , n20376 , n20377 );
xor ( n20379 , n20376 , n20377 );
xor ( n20380 , n20287 , n20320 );
and ( n20381 , n18117 , n18580 );
and ( n20382 , n20380 , n20381 );
xor ( n20383 , n20380 , n20381 );
xor ( n20384 , n20291 , n20318 );
and ( n20385 , n18118 , n18580 );
and ( n20386 , n20384 , n20385 );
xor ( n20387 , n20384 , n20385 );
xor ( n20388 , n20295 , n20316 );
and ( n20389 , n18119 , n18580 );
and ( n20390 , n20388 , n20389 );
xor ( n20391 , n20388 , n20389 );
xor ( n20392 , n20299 , n20314 );
and ( n20393 , n18120 , n18580 );
and ( n20394 , n20392 , n20393 );
xor ( n20395 , n20392 , n20393 );
xor ( n20396 , n20303 , n20312 );
and ( n20397 , n18121 , n18580 );
and ( n20398 , n20396 , n20397 );
xor ( n20399 , n20396 , n20397 );
xor ( n20400 , n20307 , n20310 );
and ( n20401 , n18122 , n18580 );
and ( n20402 , n20400 , n20401 );
and ( n20403 , n20399 , n20402 );
or ( n20404 , n20398 , n20403 );
and ( n20405 , n20395 , n20404 );
or ( n20406 , n20394 , n20405 );
and ( n20407 , n20391 , n20406 );
or ( n20408 , n20390 , n20407 );
and ( n20409 , n20387 , n20408 );
or ( n20410 , n20386 , n20409 );
and ( n20411 , n20383 , n20410 );
or ( n20412 , n20382 , n20411 );
and ( n20413 , n20379 , n20412 );
or ( n20414 , n20378 , n20413 );
and ( n20415 , n20375 , n20414 );
or ( n20416 , n20374 , n20415 );
and ( n20417 , n20371 , n20416 );
or ( n20418 , n20370 , n20417 );
and ( n20419 , n20367 , n20418 );
or ( n20420 , n20366 , n20419 );
and ( n20421 , n20363 , n20420 );
or ( n20422 , n20362 , n20421 );
and ( n20423 , n20359 , n20422 );
or ( n20424 , n20358 , n20423 );
and ( n20425 , n20355 , n20424 );
or ( n20426 , n20354 , n20425 );
and ( n20427 , n20351 , n20426 );
or ( n20428 , n20350 , n20427 );
and ( n20429 , n20347 , n20428 );
or ( n20430 , n20346 , n20429 );
and ( n20431 , n20343 , n20430 );
or ( n20432 , n20342 , n20431 );
and ( n20433 , n18107 , n18576 );
and ( n20434 , n20432 , n20433 );
xor ( n20435 , n20432 , n20433 );
xor ( n20436 , n20343 , n20430 );
and ( n20437 , n18108 , n18576 );
and ( n20438 , n20436 , n20437 );
xor ( n20439 , n20436 , n20437 );
xor ( n20440 , n20347 , n20428 );
and ( n20441 , n18109 , n18576 );
and ( n20442 , n20440 , n20441 );
xor ( n20443 , n20440 , n20441 );
xor ( n20444 , n20351 , n20426 );
and ( n20445 , n18110 , n18576 );
and ( n20446 , n20444 , n20445 );
xor ( n20447 , n20444 , n20445 );
xor ( n20448 , n20355 , n20424 );
and ( n20449 , n18111 , n18576 );
and ( n20450 , n20448 , n20449 );
xor ( n20451 , n20448 , n20449 );
xor ( n20452 , n20359 , n20422 );
and ( n20453 , n18112 , n18576 );
and ( n20454 , n20452 , n20453 );
xor ( n20455 , n20452 , n20453 );
xor ( n20456 , n20363 , n20420 );
and ( n20457 , n18113 , n18576 );
and ( n20458 , n20456 , n20457 );
xor ( n20459 , n20456 , n20457 );
xor ( n20460 , n20367 , n20418 );
and ( n20461 , n18114 , n18576 );
and ( n20462 , n20460 , n20461 );
xor ( n20463 , n20460 , n20461 );
xor ( n20464 , n20371 , n20416 );
and ( n20465 , n18115 , n18576 );
and ( n20466 , n20464 , n20465 );
xor ( n20467 , n20464 , n20465 );
xor ( n20468 , n20375 , n20414 );
and ( n20469 , n18116 , n18576 );
and ( n20470 , n20468 , n20469 );
xor ( n20471 , n20468 , n20469 );
xor ( n20472 , n20379 , n20412 );
and ( n20473 , n18117 , n18576 );
and ( n20474 , n20472 , n20473 );
xor ( n20475 , n20472 , n20473 );
xor ( n20476 , n20383 , n20410 );
and ( n20477 , n18118 , n18576 );
and ( n20478 , n20476 , n20477 );
xor ( n20479 , n20476 , n20477 );
xor ( n20480 , n20387 , n20408 );
and ( n20481 , n18119 , n18576 );
and ( n20482 , n20480 , n20481 );
xor ( n20483 , n20480 , n20481 );
xor ( n20484 , n20391 , n20406 );
and ( n20485 , n18120 , n18576 );
and ( n20486 , n20484 , n20485 );
xor ( n20487 , n20484 , n20485 );
xor ( n20488 , n20395 , n20404 );
and ( n20489 , n18121 , n18576 );
and ( n20490 , n20488 , n20489 );
xor ( n20491 , n20488 , n20489 );
xor ( n20492 , n20399 , n20402 );
and ( n20493 , n18122 , n18576 );
and ( n20494 , n20492 , n20493 );
and ( n20495 , n20491 , n20494 );
or ( n20496 , n20490 , n20495 );
and ( n20497 , n20487 , n20496 );
or ( n20498 , n20486 , n20497 );
and ( n20499 , n20483 , n20498 );
or ( n20500 , n20482 , n20499 );
and ( n20501 , n20479 , n20500 );
or ( n20502 , n20478 , n20501 );
and ( n20503 , n20475 , n20502 );
or ( n20504 , n20474 , n20503 );
and ( n20505 , n20471 , n20504 );
or ( n20506 , n20470 , n20505 );
and ( n20507 , n20467 , n20506 );
or ( n20508 , n20466 , n20507 );
and ( n20509 , n20463 , n20508 );
or ( n20510 , n20462 , n20509 );
and ( n20511 , n20459 , n20510 );
or ( n20512 , n20458 , n20511 );
and ( n20513 , n20455 , n20512 );
or ( n20514 , n20454 , n20513 );
and ( n20515 , n20451 , n20514 );
or ( n20516 , n20450 , n20515 );
and ( n20517 , n20447 , n20516 );
or ( n20518 , n20446 , n20517 );
and ( n20519 , n20443 , n20518 );
or ( n20520 , n20442 , n20519 );
and ( n20521 , n20439 , n20520 );
or ( n20522 , n20438 , n20521 );
and ( n20523 , n20435 , n20522 );
or ( n20524 , n20434 , n20523 );
and ( n20525 , n18107 , n18572 );
and ( n20526 , n20524 , n20525 );
xor ( n20527 , n20524 , n20525 );
xor ( n20528 , n20435 , n20522 );
and ( n20529 , n18108 , n18572 );
and ( n20530 , n20528 , n20529 );
xor ( n20531 , n20528 , n20529 );
xor ( n20532 , n20439 , n20520 );
and ( n20533 , n18109 , n18572 );
and ( n20534 , n20532 , n20533 );
xor ( n20535 , n20532 , n20533 );
xor ( n20536 , n20443 , n20518 );
and ( n20537 , n18110 , n18572 );
and ( n20538 , n20536 , n20537 );
xor ( n20539 , n20536 , n20537 );
xor ( n20540 , n20447 , n20516 );
and ( n20541 , n18111 , n18572 );
and ( n20542 , n20540 , n20541 );
xor ( n20543 , n20540 , n20541 );
xor ( n20544 , n20451 , n20514 );
and ( n20545 , n18112 , n18572 );
and ( n20546 , n20544 , n20545 );
xor ( n20547 , n20544 , n20545 );
xor ( n20548 , n20455 , n20512 );
and ( n20549 , n18113 , n18572 );
and ( n20550 , n20548 , n20549 );
xor ( n20551 , n20548 , n20549 );
xor ( n20552 , n20459 , n20510 );
and ( n20553 , n18114 , n18572 );
and ( n20554 , n20552 , n20553 );
xor ( n20555 , n20552 , n20553 );
xor ( n20556 , n20463 , n20508 );
and ( n20557 , n18115 , n18572 );
and ( n20558 , n20556 , n20557 );
xor ( n20559 , n20556 , n20557 );
xor ( n20560 , n20467 , n20506 );
and ( n20561 , n18116 , n18572 );
and ( n20562 , n20560 , n20561 );
xor ( n20563 , n20560 , n20561 );
xor ( n20564 , n20471 , n20504 );
and ( n20565 , n18117 , n18572 );
and ( n20566 , n20564 , n20565 );
xor ( n20567 , n20564 , n20565 );
xor ( n20568 , n20475 , n20502 );
and ( n20569 , n18118 , n18572 );
and ( n20570 , n20568 , n20569 );
xor ( n20571 , n20568 , n20569 );
xor ( n20572 , n20479 , n20500 );
and ( n20573 , n18119 , n18572 );
and ( n20574 , n20572 , n20573 );
xor ( n20575 , n20572 , n20573 );
xor ( n20576 , n20483 , n20498 );
and ( n20577 , n18120 , n18572 );
and ( n20578 , n20576 , n20577 );
xor ( n20579 , n20576 , n20577 );
xor ( n20580 , n20487 , n20496 );
and ( n20581 , n18121 , n18572 );
and ( n20582 , n20580 , n20581 );
xor ( n20583 , n20580 , n20581 );
xor ( n20584 , n20491 , n20494 );
and ( n20585 , n18122 , n18572 );
and ( n20586 , n20584 , n20585 );
and ( n20587 , n20583 , n20586 );
or ( n20588 , n20582 , n20587 );
and ( n20589 , n20579 , n20588 );
or ( n20590 , n20578 , n20589 );
and ( n20591 , n20575 , n20590 );
or ( n20592 , n20574 , n20591 );
and ( n20593 , n20571 , n20592 );
or ( n20594 , n20570 , n20593 );
and ( n20595 , n20567 , n20594 );
or ( n20596 , n20566 , n20595 );
and ( n20597 , n20563 , n20596 );
or ( n20598 , n20562 , n20597 );
and ( n20599 , n20559 , n20598 );
or ( n20600 , n20558 , n20599 );
and ( n20601 , n20555 , n20600 );
or ( n20602 , n20554 , n20601 );
and ( n20603 , n20551 , n20602 );
or ( n20604 , n20550 , n20603 );
and ( n20605 , n20547 , n20604 );
or ( n20606 , n20546 , n20605 );
and ( n20607 , n20543 , n20606 );
or ( n20608 , n20542 , n20607 );
and ( n20609 , n20539 , n20608 );
or ( n20610 , n20538 , n20609 );
and ( n20611 , n20535 , n20610 );
or ( n20612 , n20534 , n20611 );
and ( n20613 , n20531 , n20612 );
or ( n20614 , n20530 , n20613 );
and ( n20615 , n20527 , n20614 );
or ( n20616 , n20526 , n20615 );
and ( n20617 , n18107 , n18568 );
and ( n20618 , n20616 , n20617 );
xor ( n20619 , n20616 , n20617 );
xor ( n20620 , n20527 , n20614 );
and ( n20621 , n18108 , n18568 );
and ( n20622 , n20620 , n20621 );
xor ( n20623 , n20620 , n20621 );
xor ( n20624 , n20531 , n20612 );
and ( n20625 , n18109 , n18568 );
and ( n20626 , n20624 , n20625 );
xor ( n20627 , n20624 , n20625 );
xor ( n20628 , n20535 , n20610 );
and ( n20629 , n18110 , n18568 );
and ( n20630 , n20628 , n20629 );
xor ( n20631 , n20628 , n20629 );
xor ( n20632 , n20539 , n20608 );
and ( n20633 , n18111 , n18568 );
and ( n20634 , n20632 , n20633 );
xor ( n20635 , n20632 , n20633 );
xor ( n20636 , n20543 , n20606 );
and ( n20637 , n18112 , n18568 );
and ( n20638 , n20636 , n20637 );
xor ( n20639 , n20636 , n20637 );
xor ( n20640 , n20547 , n20604 );
and ( n20641 , n18113 , n18568 );
and ( n20642 , n20640 , n20641 );
xor ( n20643 , n20640 , n20641 );
xor ( n20644 , n20551 , n20602 );
and ( n20645 , n18114 , n18568 );
and ( n20646 , n20644 , n20645 );
xor ( n20647 , n20644 , n20645 );
xor ( n20648 , n20555 , n20600 );
and ( n20649 , n18115 , n18568 );
and ( n20650 , n20648 , n20649 );
xor ( n20651 , n20648 , n20649 );
xor ( n20652 , n20559 , n20598 );
and ( n20653 , n18116 , n18568 );
and ( n20654 , n20652 , n20653 );
xor ( n20655 , n20652 , n20653 );
xor ( n20656 , n20563 , n20596 );
and ( n20657 , n18117 , n18568 );
and ( n20658 , n20656 , n20657 );
xor ( n20659 , n20656 , n20657 );
xor ( n20660 , n20567 , n20594 );
and ( n20661 , n18118 , n18568 );
and ( n20662 , n20660 , n20661 );
xor ( n20663 , n20660 , n20661 );
xor ( n20664 , n20571 , n20592 );
and ( n20665 , n18119 , n18568 );
and ( n20666 , n20664 , n20665 );
xor ( n20667 , n20664 , n20665 );
xor ( n20668 , n20575 , n20590 );
and ( n20669 , n18120 , n18568 );
and ( n20670 , n20668 , n20669 );
xor ( n20671 , n20668 , n20669 );
xor ( n20672 , n20579 , n20588 );
and ( n20673 , n18121 , n18568 );
and ( n20674 , n20672 , n20673 );
xor ( n20675 , n20672 , n20673 );
xor ( n20676 , n20583 , n20586 );
and ( n20677 , n18122 , n18568 );
and ( n20678 , n20676 , n20677 );
and ( n20679 , n20675 , n20678 );
or ( n20680 , n20674 , n20679 );
and ( n20681 , n20671 , n20680 );
or ( n20682 , n20670 , n20681 );
and ( n20683 , n20667 , n20682 );
or ( n20684 , n20666 , n20683 );
and ( n20685 , n20663 , n20684 );
or ( n20686 , n20662 , n20685 );
and ( n20687 , n20659 , n20686 );
or ( n20688 , n20658 , n20687 );
and ( n20689 , n20655 , n20688 );
or ( n20690 , n20654 , n20689 );
and ( n20691 , n20651 , n20690 );
or ( n20692 , n20650 , n20691 );
and ( n20693 , n20647 , n20692 );
or ( n20694 , n20646 , n20693 );
and ( n20695 , n20643 , n20694 );
or ( n20696 , n20642 , n20695 );
and ( n20697 , n20639 , n20696 );
or ( n20698 , n20638 , n20697 );
and ( n20699 , n20635 , n20698 );
or ( n20700 , n20634 , n20699 );
and ( n20701 , n20631 , n20700 );
or ( n20702 , n20630 , n20701 );
and ( n20703 , n20627 , n20702 );
or ( n20704 , n20626 , n20703 );
and ( n20705 , n20623 , n20704 );
or ( n20706 , n20622 , n20705 );
and ( n20707 , n20619 , n20706 );
or ( n20708 , n20618 , n20707 );
and ( n20709 , n18107 , n18564 );
and ( n20710 , n20708 , n20709 );
xor ( n20711 , n20708 , n20709 );
xor ( n20712 , n20619 , n20706 );
and ( n20713 , n18108 , n18564 );
and ( n20714 , n20712 , n20713 );
xor ( n20715 , n20712 , n20713 );
xor ( n20716 , n20623 , n20704 );
and ( n20717 , n18109 , n18564 );
and ( n20718 , n20716 , n20717 );
xor ( n20719 , n20716 , n20717 );
xor ( n20720 , n20627 , n20702 );
and ( n20721 , n18110 , n18564 );
and ( n20722 , n20720 , n20721 );
xor ( n20723 , n20720 , n20721 );
xor ( n20724 , n20631 , n20700 );
and ( n20725 , n18111 , n18564 );
and ( n20726 , n20724 , n20725 );
xor ( n20727 , n20724 , n20725 );
xor ( n20728 , n20635 , n20698 );
and ( n20729 , n18112 , n18564 );
and ( n20730 , n20728 , n20729 );
xor ( n20731 , n20728 , n20729 );
xor ( n20732 , n20639 , n20696 );
and ( n20733 , n18113 , n18564 );
and ( n20734 , n20732 , n20733 );
xor ( n20735 , n20732 , n20733 );
xor ( n20736 , n20643 , n20694 );
and ( n20737 , n18114 , n18564 );
and ( n20738 , n20736 , n20737 );
xor ( n20739 , n20736 , n20737 );
xor ( n20740 , n20647 , n20692 );
and ( n20741 , n18115 , n18564 );
and ( n20742 , n20740 , n20741 );
xor ( n20743 , n20740 , n20741 );
xor ( n20744 , n20651 , n20690 );
and ( n20745 , n18116 , n18564 );
and ( n20746 , n20744 , n20745 );
xor ( n20747 , n20744 , n20745 );
xor ( n20748 , n20655 , n20688 );
and ( n20749 , n18117 , n18564 );
and ( n20750 , n20748 , n20749 );
xor ( n20751 , n20748 , n20749 );
xor ( n20752 , n20659 , n20686 );
and ( n20753 , n18118 , n18564 );
and ( n20754 , n20752 , n20753 );
xor ( n20755 , n20752 , n20753 );
xor ( n20756 , n20663 , n20684 );
and ( n20757 , n18119 , n18564 );
and ( n20758 , n20756 , n20757 );
xor ( n20759 , n20756 , n20757 );
xor ( n20760 , n20667 , n20682 );
and ( n20761 , n18120 , n18564 );
and ( n20762 , n20760 , n20761 );
xor ( n20763 , n20760 , n20761 );
xor ( n20764 , n20671 , n20680 );
and ( n20765 , n18121 , n18564 );
and ( n20766 , n20764 , n20765 );
xor ( n20767 , n20764 , n20765 );
xor ( n20768 , n20675 , n20678 );
and ( n20769 , n18122 , n18564 );
and ( n20770 , n20768 , n20769 );
and ( n20771 , n20767 , n20770 );
or ( n20772 , n20766 , n20771 );
and ( n20773 , n20763 , n20772 );
or ( n20774 , n20762 , n20773 );
and ( n20775 , n20759 , n20774 );
or ( n20776 , n20758 , n20775 );
and ( n20777 , n20755 , n20776 );
or ( n20778 , n20754 , n20777 );
and ( n20779 , n20751 , n20778 );
or ( n20780 , n20750 , n20779 );
and ( n20781 , n20747 , n20780 );
or ( n20782 , n20746 , n20781 );
and ( n20783 , n20743 , n20782 );
or ( n20784 , n20742 , n20783 );
and ( n20785 , n20739 , n20784 );
or ( n20786 , n20738 , n20785 );
and ( n20787 , n20735 , n20786 );
or ( n20788 , n20734 , n20787 );
and ( n20789 , n20731 , n20788 );
or ( n20790 , n20730 , n20789 );
and ( n20791 , n20727 , n20790 );
or ( n20792 , n20726 , n20791 );
and ( n20793 , n20723 , n20792 );
or ( n20794 , n20722 , n20793 );
and ( n20795 , n20719 , n20794 );
or ( n20796 , n20718 , n20795 );
and ( n20797 , n20715 , n20796 );
or ( n20798 , n20714 , n20797 );
and ( n20799 , n20711 , n20798 );
or ( n20800 , n20710 , n20799 );
and ( n20801 , n18107 , n18560 );
and ( n20802 , n20800 , n20801 );
xor ( n20803 , n20800 , n20801 );
xor ( n20804 , n20711 , n20798 );
and ( n20805 , n18108 , n18560 );
and ( n20806 , n20804 , n20805 );
xor ( n20807 , n20804 , n20805 );
xor ( n20808 , n20715 , n20796 );
and ( n20809 , n18109 , n18560 );
and ( n20810 , n20808 , n20809 );
xor ( n20811 , n20808 , n20809 );
xor ( n20812 , n20719 , n20794 );
and ( n20813 , n18110 , n18560 );
and ( n20814 , n20812 , n20813 );
xor ( n20815 , n20812 , n20813 );
xor ( n20816 , n20723 , n20792 );
and ( n20817 , n18111 , n18560 );
and ( n20818 , n20816 , n20817 );
xor ( n20819 , n20816 , n20817 );
xor ( n20820 , n20727 , n20790 );
and ( n20821 , n18112 , n18560 );
and ( n20822 , n20820 , n20821 );
xor ( n20823 , n20820 , n20821 );
xor ( n20824 , n20731 , n20788 );
and ( n20825 , n18113 , n18560 );
and ( n20826 , n20824 , n20825 );
xor ( n20827 , n20824 , n20825 );
xor ( n20828 , n20735 , n20786 );
and ( n20829 , n18114 , n18560 );
and ( n20830 , n20828 , n20829 );
xor ( n20831 , n20828 , n20829 );
xor ( n20832 , n20739 , n20784 );
and ( n20833 , n18115 , n18560 );
and ( n20834 , n20832 , n20833 );
xor ( n20835 , n20832 , n20833 );
xor ( n20836 , n20743 , n20782 );
and ( n20837 , n18116 , n18560 );
and ( n20838 , n20836 , n20837 );
xor ( n20839 , n20836 , n20837 );
xor ( n20840 , n20747 , n20780 );
and ( n20841 , n18117 , n18560 );
and ( n20842 , n20840 , n20841 );
xor ( n20843 , n20840 , n20841 );
xor ( n20844 , n20751 , n20778 );
and ( n20845 , n18118 , n18560 );
and ( n20846 , n20844 , n20845 );
xor ( n20847 , n20844 , n20845 );
xor ( n20848 , n20755 , n20776 );
and ( n20849 , n18119 , n18560 );
and ( n20850 , n20848 , n20849 );
xor ( n20851 , n20848 , n20849 );
xor ( n20852 , n20759 , n20774 );
and ( n20853 , n18120 , n18560 );
and ( n20854 , n20852 , n20853 );
xor ( n20855 , n20852 , n20853 );
xor ( n20856 , n20763 , n20772 );
and ( n20857 , n18121 , n18560 );
and ( n20858 , n20856 , n20857 );
xor ( n20859 , n20856 , n20857 );
xor ( n20860 , n20767 , n20770 );
and ( n20861 , n18122 , n18560 );
and ( n20862 , n20860 , n20861 );
and ( n20863 , n20859 , n20862 );
or ( n20864 , n20858 , n20863 );
and ( n20865 , n20855 , n20864 );
or ( n20866 , n20854 , n20865 );
and ( n20867 , n20851 , n20866 );
or ( n20868 , n20850 , n20867 );
and ( n20869 , n20847 , n20868 );
or ( n20870 , n20846 , n20869 );
and ( n20871 , n20843 , n20870 );
or ( n20872 , n20842 , n20871 );
and ( n20873 , n20839 , n20872 );
or ( n20874 , n20838 , n20873 );
and ( n20875 , n20835 , n20874 );
or ( n20876 , n20834 , n20875 );
and ( n20877 , n20831 , n20876 );
or ( n20878 , n20830 , n20877 );
and ( n20879 , n20827 , n20878 );
or ( n20880 , n20826 , n20879 );
and ( n20881 , n20823 , n20880 );
or ( n20882 , n20822 , n20881 );
and ( n20883 , n20819 , n20882 );
or ( n20884 , n20818 , n20883 );
and ( n20885 , n20815 , n20884 );
or ( n20886 , n20814 , n20885 );
and ( n20887 , n20811 , n20886 );
or ( n20888 , n20810 , n20887 );
and ( n20889 , n20807 , n20888 );
or ( n20890 , n20806 , n20889 );
and ( n20891 , n20803 , n20890 );
or ( n20892 , n20802 , n20891 );
and ( n20893 , n18107 , n18556 );
and ( n20894 , n20892 , n20893 );
xor ( n20895 , n20892 , n20893 );
xor ( n20896 , n20803 , n20890 );
and ( n20897 , n18108 , n18556 );
and ( n20898 , n20896 , n20897 );
xor ( n20899 , n20896 , n20897 );
xor ( n20900 , n20807 , n20888 );
and ( n20901 , n18109 , n18556 );
and ( n20902 , n20900 , n20901 );
xor ( n20903 , n20900 , n20901 );
xor ( n20904 , n20811 , n20886 );
and ( n20905 , n18110 , n18556 );
and ( n20906 , n20904 , n20905 );
xor ( n20907 , n20904 , n20905 );
xor ( n20908 , n20815 , n20884 );
and ( n20909 , n18111 , n18556 );
and ( n20910 , n20908 , n20909 );
xor ( n20911 , n20908 , n20909 );
xor ( n20912 , n20819 , n20882 );
and ( n20913 , n18112 , n18556 );
and ( n20914 , n20912 , n20913 );
xor ( n20915 , n20912 , n20913 );
xor ( n20916 , n20823 , n20880 );
and ( n20917 , n18113 , n18556 );
and ( n20918 , n20916 , n20917 );
xor ( n20919 , n20916 , n20917 );
xor ( n20920 , n20827 , n20878 );
and ( n20921 , n18114 , n18556 );
and ( n20922 , n20920 , n20921 );
xor ( n20923 , n20920 , n20921 );
xor ( n20924 , n20831 , n20876 );
and ( n20925 , n18115 , n18556 );
and ( n20926 , n20924 , n20925 );
xor ( n20927 , n20924 , n20925 );
xor ( n20928 , n20835 , n20874 );
and ( n20929 , n18116 , n18556 );
and ( n20930 , n20928 , n20929 );
xor ( n20931 , n20928 , n20929 );
xor ( n20932 , n20839 , n20872 );
and ( n20933 , n18117 , n18556 );
and ( n20934 , n20932 , n20933 );
xor ( n20935 , n20932 , n20933 );
xor ( n20936 , n20843 , n20870 );
and ( n20937 , n18118 , n18556 );
and ( n20938 , n20936 , n20937 );
xor ( n20939 , n20936 , n20937 );
xor ( n20940 , n20847 , n20868 );
and ( n20941 , n18119 , n18556 );
and ( n20942 , n20940 , n20941 );
xor ( n20943 , n20940 , n20941 );
xor ( n20944 , n20851 , n20866 );
and ( n20945 , n18120 , n18556 );
and ( n20946 , n20944 , n20945 );
xor ( n20947 , n20944 , n20945 );
xor ( n20948 , n20855 , n20864 );
and ( n20949 , n18121 , n18556 );
and ( n20950 , n20948 , n20949 );
xor ( n20951 , n20948 , n20949 );
xor ( n20952 , n20859 , n20862 );
and ( n20953 , n18122 , n18556 );
and ( n20954 , n20952 , n20953 );
and ( n20955 , n20951 , n20954 );
or ( n20956 , n20950 , n20955 );
and ( n20957 , n20947 , n20956 );
or ( n20958 , n20946 , n20957 );
and ( n20959 , n20943 , n20958 );
or ( n20960 , n20942 , n20959 );
and ( n20961 , n20939 , n20960 );
or ( n20962 , n20938 , n20961 );
and ( n20963 , n20935 , n20962 );
or ( n20964 , n20934 , n20963 );
and ( n20965 , n20931 , n20964 );
or ( n20966 , n20930 , n20965 );
and ( n20967 , n20927 , n20966 );
or ( n20968 , n20926 , n20967 );
and ( n20969 , n20923 , n20968 );
or ( n20970 , n20922 , n20969 );
and ( n20971 , n20919 , n20970 );
or ( n20972 , n20918 , n20971 );
and ( n20973 , n20915 , n20972 );
or ( n20974 , n20914 , n20973 );
and ( n20975 , n20911 , n20974 );
or ( n20976 , n20910 , n20975 );
and ( n20977 , n20907 , n20976 );
or ( n20978 , n20906 , n20977 );
and ( n20979 , n20903 , n20978 );
or ( n20980 , n20902 , n20979 );
and ( n20981 , n20899 , n20980 );
or ( n20982 , n20898 , n20981 );
and ( n20983 , n20895 , n20982 );
or ( n20984 , n20894 , n20983 );
and ( n20985 , n18107 , n18552 );
and ( n20986 , n20984 , n20985 );
xor ( n20987 , n20984 , n20985 );
xor ( n20988 , n20895 , n20982 );
and ( n20989 , n18108 , n18552 );
and ( n20990 , n20988 , n20989 );
xor ( n20991 , n20988 , n20989 );
xor ( n20992 , n20899 , n20980 );
and ( n20993 , n18109 , n18552 );
and ( n20994 , n20992 , n20993 );
xor ( n20995 , n20992 , n20993 );
xor ( n20996 , n20903 , n20978 );
and ( n20997 , n18110 , n18552 );
and ( n20998 , n20996 , n20997 );
xor ( n20999 , n20996 , n20997 );
xor ( n21000 , n20907 , n20976 );
and ( n21001 , n18111 , n18552 );
and ( n21002 , n21000 , n21001 );
xor ( n21003 , n21000 , n21001 );
xor ( n21004 , n20911 , n20974 );
and ( n21005 , n18112 , n18552 );
and ( n21006 , n21004 , n21005 );
xor ( n21007 , n21004 , n21005 );
xor ( n21008 , n20915 , n20972 );
and ( n21009 , n18113 , n18552 );
and ( n21010 , n21008 , n21009 );
xor ( n21011 , n21008 , n21009 );
xor ( n21012 , n20919 , n20970 );
and ( n21013 , n18114 , n18552 );
and ( n21014 , n21012 , n21013 );
xor ( n21015 , n21012 , n21013 );
xor ( n21016 , n20923 , n20968 );
and ( n21017 , n18115 , n18552 );
and ( n21018 , n21016 , n21017 );
xor ( n21019 , n21016 , n21017 );
xor ( n21020 , n20927 , n20966 );
and ( n21021 , n18116 , n18552 );
and ( n21022 , n21020 , n21021 );
xor ( n21023 , n21020 , n21021 );
xor ( n21024 , n20931 , n20964 );
and ( n21025 , n18117 , n18552 );
and ( n21026 , n21024 , n21025 );
xor ( n21027 , n21024 , n21025 );
xor ( n21028 , n20935 , n20962 );
and ( n21029 , n18118 , n18552 );
and ( n21030 , n21028 , n21029 );
xor ( n21031 , n21028 , n21029 );
xor ( n21032 , n20939 , n20960 );
and ( n21033 , n18119 , n18552 );
and ( n21034 , n21032 , n21033 );
xor ( n21035 , n21032 , n21033 );
xor ( n21036 , n20943 , n20958 );
and ( n21037 , n18120 , n18552 );
and ( n21038 , n21036 , n21037 );
xor ( n21039 , n21036 , n21037 );
xor ( n21040 , n20947 , n20956 );
and ( n21041 , n18121 , n18552 );
and ( n21042 , n21040 , n21041 );
xor ( n21043 , n21040 , n21041 );
xor ( n21044 , n20951 , n20954 );
and ( n21045 , n18122 , n18552 );
and ( n21046 , n21044 , n21045 );
and ( n21047 , n21043 , n21046 );
or ( n21048 , n21042 , n21047 );
and ( n21049 , n21039 , n21048 );
or ( n21050 , n21038 , n21049 );
and ( n21051 , n21035 , n21050 );
or ( n21052 , n21034 , n21051 );
and ( n21053 , n21031 , n21052 );
or ( n21054 , n21030 , n21053 );
and ( n21055 , n21027 , n21054 );
or ( n21056 , n21026 , n21055 );
and ( n21057 , n21023 , n21056 );
or ( n21058 , n21022 , n21057 );
and ( n21059 , n21019 , n21058 );
or ( n21060 , n21018 , n21059 );
and ( n21061 , n21015 , n21060 );
or ( n21062 , n21014 , n21061 );
and ( n21063 , n21011 , n21062 );
or ( n21064 , n21010 , n21063 );
and ( n21065 , n21007 , n21064 );
or ( n21066 , n21006 , n21065 );
and ( n21067 , n21003 , n21066 );
or ( n21068 , n21002 , n21067 );
and ( n21069 , n20999 , n21068 );
or ( n21070 , n20998 , n21069 );
and ( n21071 , n20995 , n21070 );
or ( n21072 , n20994 , n21071 );
and ( n21073 , n20991 , n21072 );
or ( n21074 , n20990 , n21073 );
and ( n21075 , n20987 , n21074 );
or ( n21076 , n20986 , n21075 );
and ( n21077 , n18107 , n18548 );
and ( n21078 , n21076 , n21077 );
xor ( n21079 , n21076 , n21077 );
xor ( n21080 , n20987 , n21074 );
and ( n21081 , n18108 , n18548 );
and ( n21082 , n21080 , n21081 );
xor ( n21083 , n21080 , n21081 );
xor ( n21084 , n20991 , n21072 );
and ( n21085 , n18109 , n18548 );
and ( n21086 , n21084 , n21085 );
xor ( n21087 , n21084 , n21085 );
xor ( n21088 , n20995 , n21070 );
and ( n21089 , n18110 , n18548 );
and ( n21090 , n21088 , n21089 );
xor ( n21091 , n21088 , n21089 );
xor ( n21092 , n20999 , n21068 );
and ( n21093 , n18111 , n18548 );
and ( n21094 , n21092 , n21093 );
xor ( n21095 , n21092 , n21093 );
xor ( n21096 , n21003 , n21066 );
and ( n21097 , n18112 , n18548 );
and ( n21098 , n21096 , n21097 );
xor ( n21099 , n21096 , n21097 );
xor ( n21100 , n21007 , n21064 );
and ( n21101 , n18113 , n18548 );
and ( n21102 , n21100 , n21101 );
xor ( n21103 , n21100 , n21101 );
xor ( n21104 , n21011 , n21062 );
and ( n21105 , n18114 , n18548 );
and ( n21106 , n21104 , n21105 );
xor ( n21107 , n21104 , n21105 );
xor ( n21108 , n21015 , n21060 );
and ( n21109 , n18115 , n18548 );
and ( n21110 , n21108 , n21109 );
xor ( n21111 , n21108 , n21109 );
xor ( n21112 , n21019 , n21058 );
and ( n21113 , n18116 , n18548 );
and ( n21114 , n21112 , n21113 );
xor ( n21115 , n21112 , n21113 );
xor ( n21116 , n21023 , n21056 );
and ( n21117 , n18117 , n18548 );
and ( n21118 , n21116 , n21117 );
xor ( n21119 , n21116 , n21117 );
xor ( n21120 , n21027 , n21054 );
and ( n21121 , n18118 , n18548 );
and ( n21122 , n21120 , n21121 );
xor ( n21123 , n21120 , n21121 );
xor ( n21124 , n21031 , n21052 );
and ( n21125 , n18119 , n18548 );
and ( n21126 , n21124 , n21125 );
xor ( n21127 , n21124 , n21125 );
xor ( n21128 , n21035 , n21050 );
and ( n21129 , n18120 , n18548 );
and ( n21130 , n21128 , n21129 );
xor ( n21131 , n21128 , n21129 );
xor ( n21132 , n21039 , n21048 );
and ( n21133 , n18121 , n18548 );
and ( n21134 , n21132 , n21133 );
xor ( n21135 , n21132 , n21133 );
xor ( n21136 , n21043 , n21046 );
and ( n21137 , n18122 , n18548 );
and ( n21138 , n21136 , n21137 );
and ( n21139 , n21135 , n21138 );
or ( n21140 , n21134 , n21139 );
and ( n21141 , n21131 , n21140 );
or ( n21142 , n21130 , n21141 );
and ( n21143 , n21127 , n21142 );
or ( n21144 , n21126 , n21143 );
and ( n21145 , n21123 , n21144 );
or ( n21146 , n21122 , n21145 );
and ( n21147 , n21119 , n21146 );
or ( n21148 , n21118 , n21147 );
and ( n21149 , n21115 , n21148 );
or ( n21150 , n21114 , n21149 );
and ( n21151 , n21111 , n21150 );
or ( n21152 , n21110 , n21151 );
and ( n21153 , n21107 , n21152 );
or ( n21154 , n21106 , n21153 );
and ( n21155 , n21103 , n21154 );
or ( n21156 , n21102 , n21155 );
and ( n21157 , n21099 , n21156 );
or ( n21158 , n21098 , n21157 );
and ( n21159 , n21095 , n21158 );
or ( n21160 , n21094 , n21159 );
and ( n21161 , n21091 , n21160 );
or ( n21162 , n21090 , n21161 );
and ( n21163 , n21087 , n21162 );
or ( n21164 , n21086 , n21163 );
and ( n21165 , n21083 , n21164 );
or ( n21166 , n21082 , n21165 );
and ( n21167 , n21079 , n21166 );
or ( n21168 , n21078 , n21167 );
and ( n21169 , n18107 , n18544 );
and ( n21170 , n21168 , n21169 );
xor ( n21171 , n21168 , n21169 );
xor ( n21172 , n21079 , n21166 );
and ( n21173 , n18108 , n18544 );
and ( n21174 , n21172 , n21173 );
xor ( n21175 , n21172 , n21173 );
xor ( n21176 , n21083 , n21164 );
and ( n21177 , n18109 , n18544 );
and ( n21178 , n21176 , n21177 );
xor ( n21179 , n21176 , n21177 );
xor ( n21180 , n21087 , n21162 );
and ( n21181 , n18110 , n18544 );
and ( n21182 , n21180 , n21181 );
xor ( n21183 , n21180 , n21181 );
xor ( n21184 , n21091 , n21160 );
and ( n21185 , n18111 , n18544 );
and ( n21186 , n21184 , n21185 );
xor ( n21187 , n21184 , n21185 );
xor ( n21188 , n21095 , n21158 );
and ( n21189 , n18112 , n18544 );
and ( n21190 , n21188 , n21189 );
xor ( n21191 , n21188 , n21189 );
xor ( n21192 , n21099 , n21156 );
and ( n21193 , n18113 , n18544 );
and ( n21194 , n21192 , n21193 );
xor ( n21195 , n21192 , n21193 );
xor ( n21196 , n21103 , n21154 );
and ( n21197 , n18114 , n18544 );
and ( n21198 , n21196 , n21197 );
xor ( n21199 , n21196 , n21197 );
xor ( n21200 , n21107 , n21152 );
and ( n21201 , n18115 , n18544 );
and ( n21202 , n21200 , n21201 );
xor ( n21203 , n21200 , n21201 );
xor ( n21204 , n21111 , n21150 );
and ( n21205 , n18116 , n18544 );
and ( n21206 , n21204 , n21205 );
xor ( n21207 , n21204 , n21205 );
xor ( n21208 , n21115 , n21148 );
and ( n21209 , n18117 , n18544 );
and ( n21210 , n21208 , n21209 );
xor ( n21211 , n21208 , n21209 );
xor ( n21212 , n21119 , n21146 );
and ( n21213 , n18118 , n18544 );
and ( n21214 , n21212 , n21213 );
xor ( n21215 , n21212 , n21213 );
xor ( n21216 , n21123 , n21144 );
and ( n21217 , n18119 , n18544 );
and ( n21218 , n21216 , n21217 );
xor ( n21219 , n21216 , n21217 );
xor ( n21220 , n21127 , n21142 );
and ( n21221 , n18120 , n18544 );
and ( n21222 , n21220 , n21221 );
xor ( n21223 , n21220 , n21221 );
xor ( n21224 , n21131 , n21140 );
and ( n21225 , n18121 , n18544 );
and ( n21226 , n21224 , n21225 );
xor ( n21227 , n21224 , n21225 );
xor ( n21228 , n21135 , n21138 );
and ( n21229 , n18122 , n18544 );
and ( n21230 , n21228 , n21229 );
and ( n21231 , n21227 , n21230 );
or ( n21232 , n21226 , n21231 );
and ( n21233 , n21223 , n21232 );
or ( n21234 , n21222 , n21233 );
and ( n21235 , n21219 , n21234 );
or ( n21236 , n21218 , n21235 );
and ( n21237 , n21215 , n21236 );
or ( n21238 , n21214 , n21237 );
and ( n21239 , n21211 , n21238 );
or ( n21240 , n21210 , n21239 );
and ( n21241 , n21207 , n21240 );
or ( n21242 , n21206 , n21241 );
and ( n21243 , n21203 , n21242 );
or ( n21244 , n21202 , n21243 );
and ( n21245 , n21199 , n21244 );
or ( n21246 , n21198 , n21245 );
and ( n21247 , n21195 , n21246 );
or ( n21248 , n21194 , n21247 );
and ( n21249 , n21191 , n21248 );
or ( n21250 , n21190 , n21249 );
and ( n21251 , n21187 , n21250 );
or ( n21252 , n21186 , n21251 );
and ( n21253 , n21183 , n21252 );
or ( n21254 , n21182 , n21253 );
and ( n21255 , n21179 , n21254 );
or ( n21256 , n21178 , n21255 );
and ( n21257 , n21175 , n21256 );
or ( n21258 , n21174 , n21257 );
and ( n21259 , n21171 , n21258 );
or ( n21260 , n21170 , n21259 );
and ( n21261 , n18107 , n18540 );
and ( n21262 , n21260 , n21261 );
xor ( n21263 , n21260 , n21261 );
xor ( n21264 , n21171 , n21258 );
and ( n21265 , n18108 , n18540 );
and ( n21266 , n21264 , n21265 );
xor ( n21267 , n21264 , n21265 );
xor ( n21268 , n21175 , n21256 );
and ( n21269 , n18109 , n18540 );
and ( n21270 , n21268 , n21269 );
xor ( n21271 , n21268 , n21269 );
xor ( n21272 , n21179 , n21254 );
and ( n21273 , n18110 , n18540 );
and ( n21274 , n21272 , n21273 );
xor ( n21275 , n21272 , n21273 );
xor ( n21276 , n21183 , n21252 );
and ( n21277 , n18111 , n18540 );
and ( n21278 , n21276 , n21277 );
xor ( n21279 , n21276 , n21277 );
xor ( n21280 , n21187 , n21250 );
and ( n21281 , n18112 , n18540 );
and ( n21282 , n21280 , n21281 );
xor ( n21283 , n21280 , n21281 );
xor ( n21284 , n21191 , n21248 );
and ( n21285 , n18113 , n18540 );
and ( n21286 , n21284 , n21285 );
xor ( n21287 , n21284 , n21285 );
xor ( n21288 , n21195 , n21246 );
and ( n21289 , n18114 , n18540 );
and ( n21290 , n21288 , n21289 );
xor ( n21291 , n21288 , n21289 );
xor ( n21292 , n21199 , n21244 );
and ( n21293 , n18115 , n18540 );
and ( n21294 , n21292 , n21293 );
xor ( n21295 , n21292 , n21293 );
xor ( n21296 , n21203 , n21242 );
and ( n21297 , n18116 , n18540 );
and ( n21298 , n21296 , n21297 );
xor ( n21299 , n21296 , n21297 );
xor ( n21300 , n21207 , n21240 );
and ( n21301 , n18117 , n18540 );
and ( n21302 , n21300 , n21301 );
xor ( n21303 , n21300 , n21301 );
xor ( n21304 , n21211 , n21238 );
and ( n21305 , n18118 , n18540 );
and ( n21306 , n21304 , n21305 );
xor ( n21307 , n21304 , n21305 );
xor ( n21308 , n21215 , n21236 );
and ( n21309 , n18119 , n18540 );
and ( n21310 , n21308 , n21309 );
xor ( n21311 , n21308 , n21309 );
xor ( n21312 , n21219 , n21234 );
and ( n21313 , n18120 , n18540 );
and ( n21314 , n21312 , n21313 );
xor ( n21315 , n21312 , n21313 );
xor ( n21316 , n21223 , n21232 );
and ( n21317 , n18121 , n18540 );
and ( n21318 , n21316 , n21317 );
xor ( n21319 , n21316 , n21317 );
xor ( n21320 , n21227 , n21230 );
and ( n21321 , n18122 , n18540 );
and ( n21322 , n21320 , n21321 );
and ( n21323 , n21319 , n21322 );
or ( n21324 , n21318 , n21323 );
and ( n21325 , n21315 , n21324 );
or ( n21326 , n21314 , n21325 );
and ( n21327 , n21311 , n21326 );
or ( n21328 , n21310 , n21327 );
and ( n21329 , n21307 , n21328 );
or ( n21330 , n21306 , n21329 );
and ( n21331 , n21303 , n21330 );
or ( n21332 , n21302 , n21331 );
and ( n21333 , n21299 , n21332 );
or ( n21334 , n21298 , n21333 );
and ( n21335 , n21295 , n21334 );
or ( n21336 , n21294 , n21335 );
and ( n21337 , n21291 , n21336 );
or ( n21338 , n21290 , n21337 );
and ( n21339 , n21287 , n21338 );
or ( n21340 , n21286 , n21339 );
and ( n21341 , n21283 , n21340 );
or ( n21342 , n21282 , n21341 );
and ( n21343 , n21279 , n21342 );
or ( n21344 , n21278 , n21343 );
and ( n21345 , n21275 , n21344 );
or ( n21346 , n21274 , n21345 );
and ( n21347 , n21271 , n21346 );
or ( n21348 , n21270 , n21347 );
and ( n21349 , n21267 , n21348 );
or ( n21350 , n21266 , n21349 );
and ( n21351 , n21263 , n21350 );
or ( n21352 , n21262 , n21351 );
and ( n21353 , n18107 , n18536 );
and ( n21354 , n21352 , n21353 );
xor ( n21355 , n21352 , n21353 );
xor ( n21356 , n21263 , n21350 );
and ( n21357 , n18108 , n18536 );
and ( n21358 , n21356 , n21357 );
xor ( n21359 , n21356 , n21357 );
xor ( n21360 , n21267 , n21348 );
and ( n21361 , n18109 , n18536 );
and ( n21362 , n21360 , n21361 );
xor ( n21363 , n21360 , n21361 );
xor ( n21364 , n21271 , n21346 );
and ( n21365 , n18110 , n18536 );
and ( n21366 , n21364 , n21365 );
xor ( n21367 , n21364 , n21365 );
xor ( n21368 , n21275 , n21344 );
and ( n21369 , n18111 , n18536 );
and ( n21370 , n21368 , n21369 );
xor ( n21371 , n21368 , n21369 );
xor ( n21372 , n21279 , n21342 );
and ( n21373 , n18112 , n18536 );
and ( n21374 , n21372 , n21373 );
xor ( n21375 , n21372 , n21373 );
xor ( n21376 , n21283 , n21340 );
and ( n21377 , n18113 , n18536 );
and ( n21378 , n21376 , n21377 );
xor ( n21379 , n21376 , n21377 );
xor ( n21380 , n21287 , n21338 );
and ( n21381 , n18114 , n18536 );
and ( n21382 , n21380 , n21381 );
xor ( n21383 , n21380 , n21381 );
xor ( n21384 , n21291 , n21336 );
and ( n21385 , n18115 , n18536 );
and ( n21386 , n21384 , n21385 );
xor ( n21387 , n21384 , n21385 );
xor ( n21388 , n21295 , n21334 );
and ( n21389 , n18116 , n18536 );
and ( n21390 , n21388 , n21389 );
xor ( n21391 , n21388 , n21389 );
xor ( n21392 , n21299 , n21332 );
and ( n21393 , n18117 , n18536 );
and ( n21394 , n21392 , n21393 );
xor ( n21395 , n21392 , n21393 );
xor ( n21396 , n21303 , n21330 );
and ( n21397 , n18118 , n18536 );
and ( n21398 , n21396 , n21397 );
xor ( n21399 , n21396 , n21397 );
xor ( n21400 , n21307 , n21328 );
and ( n21401 , n18119 , n18536 );
and ( n21402 , n21400 , n21401 );
xor ( n21403 , n21400 , n21401 );
xor ( n21404 , n21311 , n21326 );
and ( n21405 , n18120 , n18536 );
and ( n21406 , n21404 , n21405 );
xor ( n21407 , n21404 , n21405 );
xor ( n21408 , n21315 , n21324 );
and ( n21409 , n18121 , n18536 );
and ( n21410 , n21408 , n21409 );
xor ( n21411 , n21408 , n21409 );
xor ( n21412 , n21319 , n21322 );
and ( n21413 , n18122 , n18536 );
and ( n21414 , n21412 , n21413 );
and ( n21415 , n21411 , n21414 );
or ( n21416 , n21410 , n21415 );
and ( n21417 , n21407 , n21416 );
or ( n21418 , n21406 , n21417 );
and ( n21419 , n21403 , n21418 );
or ( n21420 , n21402 , n21419 );
and ( n21421 , n21399 , n21420 );
or ( n21422 , n21398 , n21421 );
and ( n21423 , n21395 , n21422 );
or ( n21424 , n21394 , n21423 );
and ( n21425 , n21391 , n21424 );
or ( n21426 , n21390 , n21425 );
and ( n21427 , n21387 , n21426 );
or ( n21428 , n21386 , n21427 );
and ( n21429 , n21383 , n21428 );
or ( n21430 , n21382 , n21429 );
and ( n21431 , n21379 , n21430 );
or ( n21432 , n21378 , n21431 );
and ( n21433 , n21375 , n21432 );
or ( n21434 , n21374 , n21433 );
and ( n21435 , n21371 , n21434 );
or ( n21436 , n21370 , n21435 );
and ( n21437 , n21367 , n21436 );
or ( n21438 , n21366 , n21437 );
and ( n21439 , n21363 , n21438 );
or ( n21440 , n21362 , n21439 );
and ( n21441 , n21359 , n21440 );
or ( n21442 , n21358 , n21441 );
and ( n21443 , n21355 , n21442 );
or ( n21444 , n21354 , n21443 );
and ( n21445 , n18107 , n18532 );
and ( n21446 , n21444 , n21445 );
xor ( n21447 , n21444 , n21445 );
xor ( n21448 , n21355 , n21442 );
and ( n21449 , n18108 , n18532 );
and ( n21450 , n21448 , n21449 );
xor ( n21451 , n21448 , n21449 );
xor ( n21452 , n21359 , n21440 );
and ( n21453 , n18109 , n18532 );
and ( n21454 , n21452 , n21453 );
xor ( n21455 , n21452 , n21453 );
xor ( n21456 , n21363 , n21438 );
and ( n21457 , n18110 , n18532 );
and ( n21458 , n21456 , n21457 );
xor ( n21459 , n21456 , n21457 );
xor ( n21460 , n21367 , n21436 );
and ( n21461 , n18111 , n18532 );
and ( n21462 , n21460 , n21461 );
xor ( n21463 , n21460 , n21461 );
xor ( n21464 , n21371 , n21434 );
and ( n21465 , n18112 , n18532 );
and ( n21466 , n21464 , n21465 );
xor ( n21467 , n21464 , n21465 );
xor ( n21468 , n21375 , n21432 );
and ( n21469 , n18113 , n18532 );
and ( n21470 , n21468 , n21469 );
xor ( n21471 , n21468 , n21469 );
xor ( n21472 , n21379 , n21430 );
and ( n21473 , n18114 , n18532 );
and ( n21474 , n21472 , n21473 );
xor ( n21475 , n21472 , n21473 );
xor ( n21476 , n21383 , n21428 );
and ( n21477 , n18115 , n18532 );
and ( n21478 , n21476 , n21477 );
xor ( n21479 , n21476 , n21477 );
xor ( n21480 , n21387 , n21426 );
and ( n21481 , n18116 , n18532 );
and ( n21482 , n21480 , n21481 );
xor ( n21483 , n21480 , n21481 );
xor ( n21484 , n21391 , n21424 );
and ( n21485 , n18117 , n18532 );
and ( n21486 , n21484 , n21485 );
xor ( n21487 , n21484 , n21485 );
xor ( n21488 , n21395 , n21422 );
and ( n21489 , n18118 , n18532 );
and ( n21490 , n21488 , n21489 );
xor ( n21491 , n21488 , n21489 );
xor ( n21492 , n21399 , n21420 );
and ( n21493 , n18119 , n18532 );
and ( n21494 , n21492 , n21493 );
xor ( n21495 , n21492 , n21493 );
xor ( n21496 , n21403 , n21418 );
and ( n21497 , n18120 , n18532 );
and ( n21498 , n21496 , n21497 );
xor ( n21499 , n21496 , n21497 );
xor ( n21500 , n21407 , n21416 );
and ( n21501 , n18121 , n18532 );
and ( n21502 , n21500 , n21501 );
xor ( n21503 , n21500 , n21501 );
xor ( n21504 , n21411 , n21414 );
and ( n21505 , n18122 , n18532 );
and ( n21506 , n21504 , n21505 );
and ( n21507 , n21503 , n21506 );
or ( n21508 , n21502 , n21507 );
and ( n21509 , n21499 , n21508 );
or ( n21510 , n21498 , n21509 );
and ( n21511 , n21495 , n21510 );
or ( n21512 , n21494 , n21511 );
and ( n21513 , n21491 , n21512 );
or ( n21514 , n21490 , n21513 );
and ( n21515 , n21487 , n21514 );
or ( n21516 , n21486 , n21515 );
and ( n21517 , n21483 , n21516 );
or ( n21518 , n21482 , n21517 );
and ( n21519 , n21479 , n21518 );
or ( n21520 , n21478 , n21519 );
and ( n21521 , n21475 , n21520 );
or ( n21522 , n21474 , n21521 );
and ( n21523 , n21471 , n21522 );
or ( n21524 , n21470 , n21523 );
and ( n21525 , n21467 , n21524 );
or ( n21526 , n21466 , n21525 );
and ( n21527 , n21463 , n21526 );
or ( n21528 , n21462 , n21527 );
and ( n21529 , n21459 , n21528 );
or ( n21530 , n21458 , n21529 );
and ( n21531 , n21455 , n21530 );
or ( n21532 , n21454 , n21531 );
and ( n21533 , n21451 , n21532 );
or ( n21534 , n21450 , n21533 );
and ( n21535 , n21447 , n21534 );
or ( n21536 , n21446 , n21535 );
and ( n21537 , n18107 , n18530 );
and ( n21538 , n21536 , n21537 );
xor ( n21539 , n21536 , n21537 );
xor ( n21540 , n21447 , n21534 );
and ( n21541 , n18108 , n18530 );
and ( n21542 , n21540 , n21541 );
xor ( n21543 , n21540 , n21541 );
xor ( n21544 , n21451 , n21532 );
and ( n21545 , n18109 , n18530 );
and ( n21546 , n21544 , n21545 );
xor ( n21547 , n21544 , n21545 );
xor ( n21548 , n21455 , n21530 );
and ( n21549 , n18110 , n18530 );
and ( n21550 , n21548 , n21549 );
xor ( n21551 , n21548 , n21549 );
xor ( n21552 , n21459 , n21528 );
and ( n21553 , n18111 , n18530 );
and ( n21554 , n21552 , n21553 );
xor ( n21555 , n21552 , n21553 );
xor ( n21556 , n21463 , n21526 );
and ( n21557 , n18112 , n18530 );
and ( n21558 , n21556 , n21557 );
xor ( n21559 , n21556 , n21557 );
xor ( n21560 , n21467 , n21524 );
and ( n21561 , n18113 , n18530 );
and ( n21562 , n21560 , n21561 );
xor ( n21563 , n21560 , n21561 );
xor ( n21564 , n21471 , n21522 );
and ( n21565 , n18114 , n18530 );
and ( n21566 , n21564 , n21565 );
xor ( n21567 , n21564 , n21565 );
xor ( n21568 , n21475 , n21520 );
and ( n21569 , n18115 , n18530 );
and ( n21570 , n21568 , n21569 );
xor ( n21571 , n21568 , n21569 );
xor ( n21572 , n21479 , n21518 );
and ( n21573 , n18116 , n18530 );
and ( n21574 , n21572 , n21573 );
xor ( n21575 , n21572 , n21573 );
xor ( n21576 , n21483 , n21516 );
and ( n21577 , n18117 , n18530 );
and ( n21578 , n21576 , n21577 );
xor ( n21579 , n21576 , n21577 );
xor ( n21580 , n21487 , n21514 );
and ( n21581 , n18118 , n18530 );
and ( n21582 , n21580 , n21581 );
xor ( n21583 , n21580 , n21581 );
xor ( n21584 , n21491 , n21512 );
and ( n21585 , n18119 , n18530 );
and ( n21586 , n21584 , n21585 );
xor ( n21587 , n21584 , n21585 );
xor ( n21588 , n21495 , n21510 );
and ( n21589 , n18120 , n18530 );
and ( n21590 , n21588 , n21589 );
xor ( n21591 , n21588 , n21589 );
xor ( n21592 , n21499 , n21508 );
and ( n21593 , n18121 , n18530 );
and ( n21594 , n21592 , n21593 );
xor ( n21595 , n21592 , n21593 );
xor ( n21596 , n21503 , n21506 );
and ( n21597 , n18122 , n18530 );
and ( n21598 , n21596 , n21597 );
and ( n21599 , n21595 , n21598 );
or ( n21600 , n21594 , n21599 );
and ( n21601 , n21591 , n21600 );
or ( n21602 , n21590 , n21601 );
and ( n21603 , n21587 , n21602 );
or ( n21604 , n21586 , n21603 );
and ( n21605 , n21583 , n21604 );
or ( n21606 , n21582 , n21605 );
and ( n21607 , n21579 , n21606 );
or ( n21608 , n21578 , n21607 );
and ( n21609 , n21575 , n21608 );
or ( n21610 , n21574 , n21609 );
and ( n21611 , n21571 , n21610 );
or ( n21612 , n21570 , n21611 );
and ( n21613 , n21567 , n21612 );
or ( n21614 , n21566 , n21613 );
and ( n21615 , n21563 , n21614 );
or ( n21616 , n21562 , n21615 );
and ( n21617 , n21559 , n21616 );
or ( n21618 , n21558 , n21617 );
and ( n21619 , n21555 , n21618 );
or ( n21620 , n21554 , n21619 );
and ( n21621 , n21551 , n21620 );
or ( n21622 , n21550 , n21621 );
and ( n21623 , n21547 , n21622 );
or ( n21624 , n21546 , n21623 );
and ( n21625 , n21543 , n21624 );
or ( n21626 , n21542 , n21625 );
and ( n21627 , n21539 , n21626 );
or ( n21628 , n21538 , n21627 );
and ( n21629 , n18107 , n18528 );
and ( n21630 , n21628 , n21629 );
xor ( n21631 , n21628 , n21629 );
xor ( n21632 , n21539 , n21626 );
and ( n21633 , n18108 , n18528 );
and ( n21634 , n21632 , n21633 );
xor ( n21635 , n21632 , n21633 );
xor ( n21636 , n21543 , n21624 );
and ( n21637 , n18109 , n18528 );
and ( n21638 , n21636 , n21637 );
xor ( n21639 , n21636 , n21637 );
xor ( n21640 , n21547 , n21622 );
and ( n21641 , n18110 , n18528 );
and ( n21642 , n21640 , n21641 );
xor ( n21643 , n21640 , n21641 );
xor ( n21644 , n21551 , n21620 );
and ( n21645 , n18111 , n18528 );
and ( n21646 , n21644 , n21645 );
xor ( n21647 , n21644 , n21645 );
xor ( n21648 , n21555 , n21618 );
and ( n21649 , n18112 , n18528 );
and ( n21650 , n21648 , n21649 );
xor ( n21651 , n21648 , n21649 );
xor ( n21652 , n21559 , n21616 );
and ( n21653 , n18113 , n18528 );
and ( n21654 , n21652 , n21653 );
xor ( n21655 , n21652 , n21653 );
xor ( n21656 , n21563 , n21614 );
and ( n21657 , n18114 , n18528 );
and ( n21658 , n21656 , n21657 );
xor ( n21659 , n21656 , n21657 );
xor ( n21660 , n21567 , n21612 );
and ( n21661 , n18115 , n18528 );
and ( n21662 , n21660 , n21661 );
xor ( n21663 , n21660 , n21661 );
xor ( n21664 , n21571 , n21610 );
and ( n21665 , n18116 , n18528 );
and ( n21666 , n21664 , n21665 );
xor ( n21667 , n21664 , n21665 );
xor ( n21668 , n21575 , n21608 );
and ( n21669 , n18117 , n18528 );
and ( n21670 , n21668 , n21669 );
xor ( n21671 , n21668 , n21669 );
xor ( n21672 , n21579 , n21606 );
and ( n21673 , n18118 , n18528 );
and ( n21674 , n21672 , n21673 );
xor ( n21675 , n21672 , n21673 );
xor ( n21676 , n21583 , n21604 );
and ( n21677 , n18119 , n18528 );
and ( n21678 , n21676 , n21677 );
xor ( n21679 , n21676 , n21677 );
xor ( n21680 , n21587 , n21602 );
and ( n21681 , n18120 , n18528 );
and ( n21682 , n21680 , n21681 );
xor ( n21683 , n21680 , n21681 );
xor ( n21684 , n21591 , n21600 );
and ( n21685 , n18121 , n18528 );
and ( n21686 , n21684 , n21685 );
xor ( n21687 , n21684 , n21685 );
xor ( n21688 , n21595 , n21598 );
and ( n21689 , n18122 , n18528 );
and ( n21690 , n21688 , n21689 );
and ( n21691 , n21687 , n21690 );
or ( n21692 , n21686 , n21691 );
and ( n21693 , n21683 , n21692 );
or ( n21694 , n21682 , n21693 );
and ( n21695 , n21679 , n21694 );
or ( n21696 , n21678 , n21695 );
and ( n21697 , n21675 , n21696 );
or ( n21698 , n21674 , n21697 );
and ( n21699 , n21671 , n21698 );
or ( n21700 , n21670 , n21699 );
and ( n21701 , n21667 , n21700 );
or ( n21702 , n21666 , n21701 );
and ( n21703 , n21663 , n21702 );
or ( n21704 , n21662 , n21703 );
and ( n21705 , n21659 , n21704 );
or ( n21706 , n21658 , n21705 );
and ( n21707 , n21655 , n21706 );
or ( n21708 , n21654 , n21707 );
and ( n21709 , n21651 , n21708 );
or ( n21710 , n21650 , n21709 );
and ( n21711 , n21647 , n21710 );
or ( n21712 , n21646 , n21711 );
and ( n21713 , n21643 , n21712 );
or ( n21714 , n21642 , n21713 );
and ( n21715 , n21639 , n21714 );
or ( n21716 , n21638 , n21715 );
and ( n21717 , n21635 , n21716 );
or ( n21718 , n21634 , n21717 );
and ( n21719 , n21631 , n21718 );
or ( n21720 , n21630 , n21719 );
and ( n21721 , n18107 , n18526 );
and ( n21722 , n21720 , n21721 );
xor ( n21723 , n21720 , n21721 );
xor ( n21724 , n21631 , n21718 );
and ( n21725 , n18108 , n18526 );
and ( n21726 , n21724 , n21725 );
xor ( n21727 , n21724 , n21725 );
xor ( n21728 , n21635 , n21716 );
and ( n21729 , n18109 , n18526 );
and ( n21730 , n21728 , n21729 );
xor ( n21731 , n21728 , n21729 );
xor ( n21732 , n21639 , n21714 );
and ( n21733 , n18110 , n18526 );
and ( n21734 , n21732 , n21733 );
xor ( n21735 , n21732 , n21733 );
xor ( n21736 , n21643 , n21712 );
and ( n21737 , n18111 , n18526 );
and ( n21738 , n21736 , n21737 );
xor ( n21739 , n21736 , n21737 );
xor ( n21740 , n21647 , n21710 );
and ( n21741 , n18112 , n18526 );
and ( n21742 , n21740 , n21741 );
xor ( n21743 , n21740 , n21741 );
xor ( n21744 , n21651 , n21708 );
and ( n21745 , n18113 , n18526 );
and ( n21746 , n21744 , n21745 );
xor ( n21747 , n21744 , n21745 );
xor ( n21748 , n21655 , n21706 );
and ( n21749 , n18114 , n18526 );
and ( n21750 , n21748 , n21749 );
xor ( n21751 , n21748 , n21749 );
xor ( n21752 , n21659 , n21704 );
and ( n21753 , n18115 , n18526 );
and ( n21754 , n21752 , n21753 );
xor ( n21755 , n21752 , n21753 );
xor ( n21756 , n21663 , n21702 );
and ( n21757 , n18116 , n18526 );
and ( n21758 , n21756 , n21757 );
xor ( n21759 , n21756 , n21757 );
xor ( n21760 , n21667 , n21700 );
and ( n21761 , n18117 , n18526 );
and ( n21762 , n21760 , n21761 );
xor ( n21763 , n21760 , n21761 );
xor ( n21764 , n21671 , n21698 );
and ( n21765 , n18118 , n18526 );
and ( n21766 , n21764 , n21765 );
xor ( n21767 , n21764 , n21765 );
xor ( n21768 , n21675 , n21696 );
and ( n21769 , n18119 , n18526 );
and ( n21770 , n21768 , n21769 );
xor ( n21771 , n21768 , n21769 );
xor ( n21772 , n21679 , n21694 );
and ( n21773 , n18120 , n18526 );
and ( n21774 , n21772 , n21773 );
xor ( n21775 , n21772 , n21773 );
xor ( n21776 , n21683 , n21692 );
and ( n21777 , n18121 , n18526 );
and ( n21778 , n21776 , n21777 );
xor ( n21779 , n21776 , n21777 );
xor ( n21780 , n21687 , n21690 );
and ( n21781 , n18122 , n18526 );
and ( n21782 , n21780 , n21781 );
and ( n21783 , n21779 , n21782 );
or ( n21784 , n21778 , n21783 );
and ( n21785 , n21775 , n21784 );
or ( n21786 , n21774 , n21785 );
and ( n21787 , n21771 , n21786 );
or ( n21788 , n21770 , n21787 );
and ( n21789 , n21767 , n21788 );
or ( n21790 , n21766 , n21789 );
and ( n21791 , n21763 , n21790 );
or ( n21792 , n21762 , n21791 );
and ( n21793 , n21759 , n21792 );
or ( n21794 , n21758 , n21793 );
and ( n21795 , n21755 , n21794 );
or ( n21796 , n21754 , n21795 );
and ( n21797 , n21751 , n21796 );
or ( n21798 , n21750 , n21797 );
and ( n21799 , n21747 , n21798 );
or ( n21800 , n21746 , n21799 );
and ( n21801 , n21743 , n21800 );
or ( n21802 , n21742 , n21801 );
and ( n21803 , n21739 , n21802 );
or ( n21804 , n21738 , n21803 );
and ( n21805 , n21735 , n21804 );
or ( n21806 , n21734 , n21805 );
and ( n21807 , n21731 , n21806 );
or ( n21808 , n21730 , n21807 );
and ( n21809 , n21727 , n21808 );
or ( n21810 , n21726 , n21809 );
and ( n21811 , n21723 , n21810 );
or ( n21812 , n21722 , n21811 );
and ( n21813 , n18107 , n18524 );
and ( n21814 , n21812 , n21813 );
xor ( n21815 , n21812 , n21813 );
xor ( n21816 , n21723 , n21810 );
and ( n21817 , n18108 , n18524 );
and ( n21818 , n21816 , n21817 );
xor ( n21819 , n21816 , n21817 );
xor ( n21820 , n21727 , n21808 );
and ( n21821 , n18109 , n18524 );
and ( n21822 , n21820 , n21821 );
xor ( n21823 , n21820 , n21821 );
xor ( n21824 , n21731 , n21806 );
and ( n21825 , n18110 , n18524 );
and ( n21826 , n21824 , n21825 );
xor ( n21827 , n21824 , n21825 );
xor ( n21828 , n21735 , n21804 );
and ( n21829 , n18111 , n18524 );
and ( n21830 , n21828 , n21829 );
xor ( n21831 , n21828 , n21829 );
xor ( n21832 , n21739 , n21802 );
and ( n21833 , n18112 , n18524 );
and ( n21834 , n21832 , n21833 );
xor ( n21835 , n21832 , n21833 );
xor ( n21836 , n21743 , n21800 );
and ( n21837 , n18113 , n18524 );
and ( n21838 , n21836 , n21837 );
xor ( n21839 , n21836 , n21837 );
xor ( n21840 , n21747 , n21798 );
and ( n21841 , n18114 , n18524 );
and ( n21842 , n21840 , n21841 );
xor ( n21843 , n21840 , n21841 );
xor ( n21844 , n21751 , n21796 );
and ( n21845 , n18115 , n18524 );
and ( n21846 , n21844 , n21845 );
xor ( n21847 , n21844 , n21845 );
xor ( n21848 , n21755 , n21794 );
and ( n21849 , n18116 , n18524 );
and ( n21850 , n21848 , n21849 );
xor ( n21851 , n21848 , n21849 );
xor ( n21852 , n21759 , n21792 );
and ( n21853 , n18117 , n18524 );
and ( n21854 , n21852 , n21853 );
xor ( n21855 , n21852 , n21853 );
xor ( n21856 , n21763 , n21790 );
and ( n21857 , n18118 , n18524 );
and ( n21858 , n21856 , n21857 );
xor ( n21859 , n21856 , n21857 );
xor ( n21860 , n21767 , n21788 );
and ( n21861 , n18119 , n18524 );
and ( n21862 , n21860 , n21861 );
xor ( n21863 , n21860 , n21861 );
xor ( n21864 , n21771 , n21786 );
and ( n21865 , n18120 , n18524 );
and ( n21866 , n21864 , n21865 );
xor ( n21867 , n21864 , n21865 );
xor ( n21868 , n21775 , n21784 );
and ( n21869 , n18121 , n18524 );
and ( n21870 , n21868 , n21869 );
xor ( n21871 , n21868 , n21869 );
xor ( n21872 , n21779 , n21782 );
and ( n21873 , n18122 , n18524 );
and ( n21874 , n21872 , n21873 );
and ( n21875 , n21871 , n21874 );
or ( n21876 , n21870 , n21875 );
and ( n21877 , n21867 , n21876 );
or ( n21878 , n21866 , n21877 );
and ( n21879 , n21863 , n21878 );
or ( n21880 , n21862 , n21879 );
and ( n21881 , n21859 , n21880 );
or ( n21882 , n21858 , n21881 );
and ( n21883 , n21855 , n21882 );
or ( n21884 , n21854 , n21883 );
and ( n21885 , n21851 , n21884 );
or ( n21886 , n21850 , n21885 );
and ( n21887 , n21847 , n21886 );
or ( n21888 , n21846 , n21887 );
and ( n21889 , n21843 , n21888 );
or ( n21890 , n21842 , n21889 );
and ( n21891 , n21839 , n21890 );
or ( n21892 , n21838 , n21891 );
and ( n21893 , n21835 , n21892 );
or ( n21894 , n21834 , n21893 );
and ( n21895 , n21831 , n21894 );
or ( n21896 , n21830 , n21895 );
and ( n21897 , n21827 , n21896 );
or ( n21898 , n21826 , n21897 );
and ( n21899 , n21823 , n21898 );
or ( n21900 , n21822 , n21899 );
and ( n21901 , n21819 , n21900 );
or ( n21902 , n21818 , n21901 );
and ( n21903 , n21815 , n21902 );
or ( n21904 , n21814 , n21903 );
and ( n21905 , n18107 , n18522 );
and ( n21906 , n21904 , n21905 );
xor ( n21907 , n21904 , n21905 );
xor ( n21908 , n21815 , n21902 );
and ( n21909 , n18108 , n18522 );
and ( n21910 , n21908 , n21909 );
xor ( n21911 , n21908 , n21909 );
xor ( n21912 , n21819 , n21900 );
and ( n21913 , n18109 , n18522 );
and ( n21914 , n21912 , n21913 );
xor ( n21915 , n21912 , n21913 );
xor ( n21916 , n21823 , n21898 );
and ( n21917 , n18110 , n18522 );
and ( n21918 , n21916 , n21917 );
xor ( n21919 , n21916 , n21917 );
xor ( n21920 , n21827 , n21896 );
and ( n21921 , n18111 , n18522 );
and ( n21922 , n21920 , n21921 );
xor ( n21923 , n21920 , n21921 );
xor ( n21924 , n21831 , n21894 );
and ( n21925 , n18112 , n18522 );
and ( n21926 , n21924 , n21925 );
xor ( n21927 , n21924 , n21925 );
xor ( n21928 , n21835 , n21892 );
and ( n21929 , n18113 , n18522 );
and ( n21930 , n21928 , n21929 );
xor ( n21931 , n21928 , n21929 );
xor ( n21932 , n21839 , n21890 );
and ( n21933 , n18114 , n18522 );
and ( n21934 , n21932 , n21933 );
xor ( n21935 , n21932 , n21933 );
xor ( n21936 , n21843 , n21888 );
and ( n21937 , n18115 , n18522 );
and ( n21938 , n21936 , n21937 );
xor ( n21939 , n21936 , n21937 );
xor ( n21940 , n21847 , n21886 );
and ( n21941 , n18116 , n18522 );
and ( n21942 , n21940 , n21941 );
xor ( n21943 , n21940 , n21941 );
xor ( n21944 , n21851 , n21884 );
and ( n21945 , n18117 , n18522 );
and ( n21946 , n21944 , n21945 );
xor ( n21947 , n21944 , n21945 );
xor ( n21948 , n21855 , n21882 );
and ( n21949 , n18118 , n18522 );
and ( n21950 , n21948 , n21949 );
xor ( n21951 , n21948 , n21949 );
xor ( n21952 , n21859 , n21880 );
and ( n21953 , n18119 , n18522 );
and ( n21954 , n21952 , n21953 );
xor ( n21955 , n21952 , n21953 );
xor ( n21956 , n21863 , n21878 );
and ( n21957 , n18120 , n18522 );
and ( n21958 , n21956 , n21957 );
xor ( n21959 , n21956 , n21957 );
xor ( n21960 , n21867 , n21876 );
and ( n21961 , n18121 , n18522 );
and ( n21962 , n21960 , n21961 );
xor ( n21963 , n21960 , n21961 );
xor ( n21964 , n21871 , n21874 );
and ( n21965 , n18122 , n18522 );
and ( n21966 , n21964 , n21965 );
and ( n21967 , n21963 , n21966 );
or ( n21968 , n21962 , n21967 );
and ( n21969 , n21959 , n21968 );
or ( n21970 , n21958 , n21969 );
and ( n21971 , n21955 , n21970 );
or ( n21972 , n21954 , n21971 );
and ( n21973 , n21951 , n21972 );
or ( n21974 , n21950 , n21973 );
and ( n21975 , n21947 , n21974 );
or ( n21976 , n21946 , n21975 );
and ( n21977 , n21943 , n21976 );
or ( n21978 , n21942 , n21977 );
and ( n21979 , n21939 , n21978 );
or ( n21980 , n21938 , n21979 );
and ( n21981 , n21935 , n21980 );
or ( n21982 , n21934 , n21981 );
and ( n21983 , n21931 , n21982 );
or ( n21984 , n21930 , n21983 );
and ( n21985 , n21927 , n21984 );
or ( n21986 , n21926 , n21985 );
and ( n21987 , n21923 , n21986 );
or ( n21988 , n21922 , n21987 );
and ( n21989 , n21919 , n21988 );
or ( n21990 , n21918 , n21989 );
and ( n21991 , n21915 , n21990 );
or ( n21992 , n21914 , n21991 );
and ( n21993 , n21911 , n21992 );
or ( n21994 , n21910 , n21993 );
and ( n21995 , n21907 , n21994 );
or ( n21996 , n21906 , n21995 );
and ( n21997 , n18107 , n18520 );
and ( n21998 , n21996 , n21997 );
xor ( n21999 , n21996 , n21997 );
xor ( n22000 , n21907 , n21994 );
and ( n22001 , n18108 , n18520 );
and ( n22002 , n22000 , n22001 );
xor ( n22003 , n22000 , n22001 );
xor ( n22004 , n21911 , n21992 );
and ( n22005 , n18109 , n18520 );
and ( n22006 , n22004 , n22005 );
xor ( n22007 , n22004 , n22005 );
xor ( n22008 , n21915 , n21990 );
and ( n22009 , n18110 , n18520 );
and ( n22010 , n22008 , n22009 );
xor ( n22011 , n22008 , n22009 );
xor ( n22012 , n21919 , n21988 );
and ( n22013 , n18111 , n18520 );
and ( n22014 , n22012 , n22013 );
xor ( n22015 , n22012 , n22013 );
xor ( n22016 , n21923 , n21986 );
and ( n22017 , n18112 , n18520 );
and ( n22018 , n22016 , n22017 );
xor ( n22019 , n22016 , n22017 );
xor ( n22020 , n21927 , n21984 );
and ( n22021 , n18113 , n18520 );
and ( n22022 , n22020 , n22021 );
xor ( n22023 , n22020 , n22021 );
xor ( n22024 , n21931 , n21982 );
and ( n22025 , n18114 , n18520 );
and ( n22026 , n22024 , n22025 );
xor ( n22027 , n22024 , n22025 );
xor ( n22028 , n21935 , n21980 );
and ( n22029 , n18115 , n18520 );
and ( n22030 , n22028 , n22029 );
xor ( n22031 , n22028 , n22029 );
xor ( n22032 , n21939 , n21978 );
and ( n22033 , n18116 , n18520 );
and ( n22034 , n22032 , n22033 );
xor ( n22035 , n22032 , n22033 );
xor ( n22036 , n21943 , n21976 );
and ( n22037 , n18117 , n18520 );
and ( n22038 , n22036 , n22037 );
xor ( n22039 , n22036 , n22037 );
xor ( n22040 , n21947 , n21974 );
and ( n22041 , n18118 , n18520 );
and ( n22042 , n22040 , n22041 );
xor ( n22043 , n22040 , n22041 );
xor ( n22044 , n21951 , n21972 );
and ( n22045 , n18119 , n18520 );
and ( n22046 , n22044 , n22045 );
xor ( n22047 , n22044 , n22045 );
xor ( n22048 , n21955 , n21970 );
and ( n22049 , n18120 , n18520 );
and ( n22050 , n22048 , n22049 );
xor ( n22051 , n22048 , n22049 );
xor ( n22052 , n21959 , n21968 );
and ( n22053 , n18121 , n18520 );
and ( n22054 , n22052 , n22053 );
xor ( n22055 , n22052 , n22053 );
xor ( n22056 , n21963 , n21966 );
and ( n22057 , n18122 , n18520 );
and ( n22058 , n22056 , n22057 );
and ( n22059 , n22055 , n22058 );
or ( n22060 , n22054 , n22059 );
and ( n22061 , n22051 , n22060 );
or ( n22062 , n22050 , n22061 );
and ( n22063 , n22047 , n22062 );
or ( n22064 , n22046 , n22063 );
and ( n22065 , n22043 , n22064 );
or ( n22066 , n22042 , n22065 );
and ( n22067 , n22039 , n22066 );
or ( n22068 , n22038 , n22067 );
and ( n22069 , n22035 , n22068 );
or ( n22070 , n22034 , n22069 );
and ( n22071 , n22031 , n22070 );
or ( n22072 , n22030 , n22071 );
and ( n22073 , n22027 , n22072 );
or ( n22074 , n22026 , n22073 );
and ( n22075 , n22023 , n22074 );
or ( n22076 , n22022 , n22075 );
and ( n22077 , n22019 , n22076 );
or ( n22078 , n22018 , n22077 );
and ( n22079 , n22015 , n22078 );
or ( n22080 , n22014 , n22079 );
and ( n22081 , n22011 , n22080 );
or ( n22082 , n22010 , n22081 );
and ( n22083 , n22007 , n22082 );
or ( n22084 , n22006 , n22083 );
and ( n22085 , n22003 , n22084 );
or ( n22086 , n22002 , n22085 );
and ( n22087 , n21999 , n22086 );
or ( n22088 , n21998 , n22087 );
and ( n22089 , n18107 , n18518 );
and ( n22090 , n22088 , n22089 );
xor ( n22091 , n22088 , n22089 );
xor ( n22092 , n21999 , n22086 );
and ( n22093 , n18108 , n18518 );
and ( n22094 , n22092 , n22093 );
xor ( n22095 , n22092 , n22093 );
xor ( n22096 , n22003 , n22084 );
and ( n22097 , n18109 , n18518 );
and ( n22098 , n22096 , n22097 );
xor ( n22099 , n22096 , n22097 );
xor ( n22100 , n22007 , n22082 );
and ( n22101 , n18110 , n18518 );
and ( n22102 , n22100 , n22101 );
xor ( n22103 , n22100 , n22101 );
xor ( n22104 , n22011 , n22080 );
and ( n22105 , n18111 , n18518 );
and ( n22106 , n22104 , n22105 );
xor ( n22107 , n22104 , n22105 );
xor ( n22108 , n22015 , n22078 );
and ( n22109 , n18112 , n18518 );
and ( n22110 , n22108 , n22109 );
xor ( n22111 , n22108 , n22109 );
xor ( n22112 , n22019 , n22076 );
and ( n22113 , n18113 , n18518 );
and ( n22114 , n22112 , n22113 );
xor ( n22115 , n22112 , n22113 );
xor ( n22116 , n22023 , n22074 );
and ( n22117 , n18114 , n18518 );
and ( n22118 , n22116 , n22117 );
xor ( n22119 , n22116 , n22117 );
xor ( n22120 , n22027 , n22072 );
and ( n22121 , n18115 , n18518 );
and ( n22122 , n22120 , n22121 );
xor ( n22123 , n22120 , n22121 );
xor ( n22124 , n22031 , n22070 );
and ( n22125 , n18116 , n18518 );
and ( n22126 , n22124 , n22125 );
xor ( n22127 , n22124 , n22125 );
xor ( n22128 , n22035 , n22068 );
and ( n22129 , n18117 , n18518 );
and ( n22130 , n22128 , n22129 );
xor ( n22131 , n22128 , n22129 );
xor ( n22132 , n22039 , n22066 );
and ( n22133 , n18118 , n18518 );
and ( n22134 , n22132 , n22133 );
xor ( n22135 , n22132 , n22133 );
xor ( n22136 , n22043 , n22064 );
and ( n22137 , n18119 , n18518 );
and ( n22138 , n22136 , n22137 );
xor ( n22139 , n22136 , n22137 );
xor ( n22140 , n22047 , n22062 );
and ( n22141 , n18120 , n18518 );
and ( n22142 , n22140 , n22141 );
xor ( n22143 , n22140 , n22141 );
xor ( n22144 , n22051 , n22060 );
and ( n22145 , n18121 , n18518 );
and ( n22146 , n22144 , n22145 );
xor ( n22147 , n22144 , n22145 );
xor ( n22148 , n22055 , n22058 );
and ( n22149 , n18122 , n18518 );
and ( n22150 , n22148 , n22149 );
and ( n22151 , n22147 , n22150 );
or ( n22152 , n22146 , n22151 );
and ( n22153 , n22143 , n22152 );
or ( n22154 , n22142 , n22153 );
and ( n22155 , n22139 , n22154 );
or ( n22156 , n22138 , n22155 );
and ( n22157 , n22135 , n22156 );
or ( n22158 , n22134 , n22157 );
and ( n22159 , n22131 , n22158 );
or ( n22160 , n22130 , n22159 );
and ( n22161 , n22127 , n22160 );
or ( n22162 , n22126 , n22161 );
and ( n22163 , n22123 , n22162 );
or ( n22164 , n22122 , n22163 );
and ( n22165 , n22119 , n22164 );
or ( n22166 , n22118 , n22165 );
and ( n22167 , n22115 , n22166 );
or ( n22168 , n22114 , n22167 );
and ( n22169 , n22111 , n22168 );
or ( n22170 , n22110 , n22169 );
and ( n22171 , n22107 , n22170 );
or ( n22172 , n22106 , n22171 );
and ( n22173 , n22103 , n22172 );
or ( n22174 , n22102 , n22173 );
and ( n22175 , n22099 , n22174 );
or ( n22176 , n22098 , n22175 );
and ( n22177 , n22095 , n22176 );
or ( n22178 , n22094 , n22177 );
and ( n22179 , n22091 , n22178 );
or ( n22180 , n22090 , n22179 );
and ( n22181 , n18107 , n18516 );
and ( n22182 , n22180 , n22181 );
xor ( n22183 , n22180 , n22181 );
xor ( n22184 , n22091 , n22178 );
and ( n22185 , n18108 , n18516 );
and ( n22186 , n22184 , n22185 );
xor ( n22187 , n22184 , n22185 );
xor ( n22188 , n22095 , n22176 );
and ( n22189 , n18109 , n18516 );
and ( n22190 , n22188 , n22189 );
xor ( n22191 , n22188 , n22189 );
xor ( n22192 , n22099 , n22174 );
and ( n22193 , n18110 , n18516 );
and ( n22194 , n22192 , n22193 );
xor ( n22195 , n22192 , n22193 );
xor ( n22196 , n22103 , n22172 );
and ( n22197 , n18111 , n18516 );
and ( n22198 , n22196 , n22197 );
xor ( n22199 , n22196 , n22197 );
xor ( n22200 , n22107 , n22170 );
and ( n22201 , n18112 , n18516 );
and ( n22202 , n22200 , n22201 );
xor ( n22203 , n22200 , n22201 );
xor ( n22204 , n22111 , n22168 );
and ( n22205 , n18113 , n18516 );
and ( n22206 , n22204 , n22205 );
xor ( n22207 , n22204 , n22205 );
xor ( n22208 , n22115 , n22166 );
and ( n22209 , n18114 , n18516 );
and ( n22210 , n22208 , n22209 );
xor ( n22211 , n22208 , n22209 );
xor ( n22212 , n22119 , n22164 );
and ( n22213 , n18115 , n18516 );
and ( n22214 , n22212 , n22213 );
xor ( n22215 , n22212 , n22213 );
xor ( n22216 , n22123 , n22162 );
and ( n22217 , n18116 , n18516 );
and ( n22218 , n22216 , n22217 );
xor ( n22219 , n22216 , n22217 );
xor ( n22220 , n22127 , n22160 );
and ( n22221 , n18117 , n18516 );
and ( n22222 , n22220 , n22221 );
xor ( n22223 , n22220 , n22221 );
xor ( n22224 , n22131 , n22158 );
and ( n22225 , n18118 , n18516 );
and ( n22226 , n22224 , n22225 );
xor ( n22227 , n22224 , n22225 );
xor ( n22228 , n22135 , n22156 );
and ( n22229 , n18119 , n18516 );
and ( n22230 , n22228 , n22229 );
xor ( n22231 , n22228 , n22229 );
xor ( n22232 , n22139 , n22154 );
and ( n22233 , n18120 , n18516 );
and ( n22234 , n22232 , n22233 );
xor ( n22235 , n22232 , n22233 );
xor ( n22236 , n22143 , n22152 );
and ( n22237 , n18121 , n18516 );
and ( n22238 , n22236 , n22237 );
xor ( n22239 , n22236 , n22237 );
xor ( n22240 , n22147 , n22150 );
and ( n22241 , n18122 , n18516 );
and ( n22242 , n22240 , n22241 );
and ( n22243 , n22239 , n22242 );
or ( n22244 , n22238 , n22243 );
and ( n22245 , n22235 , n22244 );
or ( n22246 , n22234 , n22245 );
and ( n22247 , n22231 , n22246 );
or ( n22248 , n22230 , n22247 );
and ( n22249 , n22227 , n22248 );
or ( n22250 , n22226 , n22249 );
and ( n22251 , n22223 , n22250 );
or ( n22252 , n22222 , n22251 );
and ( n22253 , n22219 , n22252 );
or ( n22254 , n22218 , n22253 );
and ( n22255 , n22215 , n22254 );
or ( n22256 , n22214 , n22255 );
and ( n22257 , n22211 , n22256 );
or ( n22258 , n22210 , n22257 );
and ( n22259 , n22207 , n22258 );
or ( n22260 , n22206 , n22259 );
and ( n22261 , n22203 , n22260 );
or ( n22262 , n22202 , n22261 );
and ( n22263 , n22199 , n22262 );
or ( n22264 , n22198 , n22263 );
and ( n22265 , n22195 , n22264 );
or ( n22266 , n22194 , n22265 );
and ( n22267 , n22191 , n22266 );
or ( n22268 , n22190 , n22267 );
and ( n22269 , n22187 , n22268 );
or ( n22270 , n22186 , n22269 );
and ( n22271 , n22183 , n22270 );
or ( n22272 , n22182 , n22271 );
and ( n22273 , n18107 , n18514 );
and ( n22274 , n22272 , n22273 );
xor ( n22275 , n22272 , n22273 );
xor ( n22276 , n22183 , n22270 );
and ( n22277 , n18108 , n18514 );
and ( n22278 , n22276 , n22277 );
xor ( n22279 , n22276 , n22277 );
xor ( n22280 , n22187 , n22268 );
and ( n22281 , n18109 , n18514 );
and ( n22282 , n22280 , n22281 );
xor ( n22283 , n22280 , n22281 );
xor ( n22284 , n22191 , n22266 );
and ( n22285 , n18110 , n18514 );
and ( n22286 , n22284 , n22285 );
xor ( n22287 , n22284 , n22285 );
xor ( n22288 , n22195 , n22264 );
and ( n22289 , n18111 , n18514 );
and ( n22290 , n22288 , n22289 );
xor ( n22291 , n22288 , n22289 );
xor ( n22292 , n22199 , n22262 );
and ( n22293 , n18112 , n18514 );
and ( n22294 , n22292 , n22293 );
xor ( n22295 , n22292 , n22293 );
xor ( n22296 , n22203 , n22260 );
and ( n22297 , n18113 , n18514 );
and ( n22298 , n22296 , n22297 );
xor ( n22299 , n22296 , n22297 );
xor ( n22300 , n22207 , n22258 );
and ( n22301 , n18114 , n18514 );
and ( n22302 , n22300 , n22301 );
xor ( n22303 , n22300 , n22301 );
xor ( n22304 , n22211 , n22256 );
and ( n22305 , n18115 , n18514 );
and ( n22306 , n22304 , n22305 );
xor ( n22307 , n22304 , n22305 );
xor ( n22308 , n22215 , n22254 );
and ( n22309 , n18116 , n18514 );
and ( n22310 , n22308 , n22309 );
xor ( n22311 , n22308 , n22309 );
xor ( n22312 , n22219 , n22252 );
and ( n22313 , n18117 , n18514 );
and ( n22314 , n22312 , n22313 );
xor ( n22315 , n22312 , n22313 );
xor ( n22316 , n22223 , n22250 );
and ( n22317 , n18118 , n18514 );
and ( n22318 , n22316 , n22317 );
xor ( n22319 , n22316 , n22317 );
xor ( n22320 , n22227 , n22248 );
and ( n22321 , n18119 , n18514 );
and ( n22322 , n22320 , n22321 );
xor ( n22323 , n22320 , n22321 );
xor ( n22324 , n22231 , n22246 );
and ( n22325 , n18120 , n18514 );
and ( n22326 , n22324 , n22325 );
xor ( n22327 , n22324 , n22325 );
xor ( n22328 , n22235 , n22244 );
and ( n22329 , n18121 , n18514 );
and ( n22330 , n22328 , n22329 );
xor ( n22331 , n22328 , n22329 );
xor ( n22332 , n22239 , n22242 );
and ( n22333 , n18122 , n18514 );
and ( n22334 , n22332 , n22333 );
and ( n22335 , n22331 , n22334 );
or ( n22336 , n22330 , n22335 );
and ( n22337 , n22327 , n22336 );
or ( n22338 , n22326 , n22337 );
and ( n22339 , n22323 , n22338 );
or ( n22340 , n22322 , n22339 );
and ( n22341 , n22319 , n22340 );
or ( n22342 , n22318 , n22341 );
and ( n22343 , n22315 , n22342 );
or ( n22344 , n22314 , n22343 );
and ( n22345 , n22311 , n22344 );
or ( n22346 , n22310 , n22345 );
and ( n22347 , n22307 , n22346 );
or ( n22348 , n22306 , n22347 );
and ( n22349 , n22303 , n22348 );
or ( n22350 , n22302 , n22349 );
and ( n22351 , n22299 , n22350 );
or ( n22352 , n22298 , n22351 );
and ( n22353 , n22295 , n22352 );
or ( n22354 , n22294 , n22353 );
and ( n22355 , n22291 , n22354 );
or ( n22356 , n22290 , n22355 );
and ( n22357 , n22287 , n22356 );
or ( n22358 , n22286 , n22357 );
and ( n22359 , n22283 , n22358 );
or ( n22360 , n22282 , n22359 );
and ( n22361 , n22279 , n22360 );
or ( n22362 , n22278 , n22361 );
and ( n22363 , n22275 , n22362 );
or ( n22364 , n22274 , n22363 );
and ( n22365 , n18107 , n18512 );
and ( n22366 , n22364 , n22365 );
xor ( n22367 , n22364 , n22365 );
xor ( n22368 , n22275 , n22362 );
and ( n22369 , n18108 , n18512 );
and ( n22370 , n22368 , n22369 );
xor ( n22371 , n22368 , n22369 );
xor ( n22372 , n22279 , n22360 );
and ( n22373 , n18109 , n18512 );
and ( n22374 , n22372 , n22373 );
xor ( n22375 , n22372 , n22373 );
xor ( n22376 , n22283 , n22358 );
and ( n22377 , n18110 , n18512 );
and ( n22378 , n22376 , n22377 );
xor ( n22379 , n22376 , n22377 );
xor ( n22380 , n22287 , n22356 );
and ( n22381 , n18111 , n18512 );
and ( n22382 , n22380 , n22381 );
xor ( n22383 , n22380 , n22381 );
xor ( n22384 , n22291 , n22354 );
and ( n22385 , n18112 , n18512 );
and ( n22386 , n22384 , n22385 );
xor ( n22387 , n22384 , n22385 );
xor ( n22388 , n22295 , n22352 );
and ( n22389 , n18113 , n18512 );
and ( n22390 , n22388 , n22389 );
xor ( n22391 , n22388 , n22389 );
xor ( n22392 , n22299 , n22350 );
and ( n22393 , n18114 , n18512 );
and ( n22394 , n22392 , n22393 );
xor ( n22395 , n22392 , n22393 );
xor ( n22396 , n22303 , n22348 );
and ( n22397 , n18115 , n18512 );
and ( n22398 , n22396 , n22397 );
xor ( n22399 , n22396 , n22397 );
xor ( n22400 , n22307 , n22346 );
and ( n22401 , n18116 , n18512 );
and ( n22402 , n22400 , n22401 );
xor ( n22403 , n22400 , n22401 );
xor ( n22404 , n22311 , n22344 );
and ( n22405 , n18117 , n18512 );
and ( n22406 , n22404 , n22405 );
xor ( n22407 , n22404 , n22405 );
xor ( n22408 , n22315 , n22342 );
and ( n22409 , n18118 , n18512 );
and ( n22410 , n22408 , n22409 );
xor ( n22411 , n22408 , n22409 );
xor ( n22412 , n22319 , n22340 );
and ( n22413 , n18119 , n18512 );
and ( n22414 , n22412 , n22413 );
xor ( n22415 , n22412 , n22413 );
xor ( n22416 , n22323 , n22338 );
and ( n22417 , n18120 , n18512 );
and ( n22418 , n22416 , n22417 );
xor ( n22419 , n22416 , n22417 );
xor ( n22420 , n22327 , n22336 );
and ( n22421 , n18121 , n18512 );
and ( n22422 , n22420 , n22421 );
xor ( n22423 , n22420 , n22421 );
xor ( n22424 , n22331 , n22334 );
and ( n22425 , n18122 , n18512 );
and ( n22426 , n22424 , n22425 );
and ( n22427 , n22423 , n22426 );
or ( n22428 , n22422 , n22427 );
and ( n22429 , n22419 , n22428 );
or ( n22430 , n22418 , n22429 );
and ( n22431 , n22415 , n22430 );
or ( n22432 , n22414 , n22431 );
and ( n22433 , n22411 , n22432 );
or ( n22434 , n22410 , n22433 );
and ( n22435 , n22407 , n22434 );
or ( n22436 , n22406 , n22435 );
and ( n22437 , n22403 , n22436 );
or ( n22438 , n22402 , n22437 );
and ( n22439 , n22399 , n22438 );
or ( n22440 , n22398 , n22439 );
and ( n22441 , n22395 , n22440 );
or ( n22442 , n22394 , n22441 );
and ( n22443 , n22391 , n22442 );
or ( n22444 , n22390 , n22443 );
and ( n22445 , n22387 , n22444 );
or ( n22446 , n22386 , n22445 );
and ( n22447 , n22383 , n22446 );
or ( n22448 , n22382 , n22447 );
and ( n22449 , n22379 , n22448 );
or ( n22450 , n22378 , n22449 );
and ( n22451 , n22375 , n22450 );
or ( n22452 , n22374 , n22451 );
and ( n22453 , n22371 , n22452 );
or ( n22454 , n22370 , n22453 );
and ( n22455 , n22367 , n22454 );
or ( n22456 , n22366 , n22455 );
and ( n22457 , n18107 , n18510 );
and ( n22458 , n22456 , n22457 );
xor ( n22459 , n22456 , n22457 );
xor ( n22460 , n22367 , n22454 );
and ( n22461 , n18108 , n18510 );
and ( n22462 , n22460 , n22461 );
xor ( n22463 , n22460 , n22461 );
xor ( n22464 , n22371 , n22452 );
and ( n22465 , n18109 , n18510 );
and ( n22466 , n22464 , n22465 );
xor ( n22467 , n22464 , n22465 );
xor ( n22468 , n22375 , n22450 );
and ( n22469 , n18110 , n18510 );
and ( n22470 , n22468 , n22469 );
xor ( n22471 , n22468 , n22469 );
xor ( n22472 , n22379 , n22448 );
and ( n22473 , n18111 , n18510 );
and ( n22474 , n22472 , n22473 );
xor ( n22475 , n22472 , n22473 );
xor ( n22476 , n22383 , n22446 );
and ( n22477 , n18112 , n18510 );
and ( n22478 , n22476 , n22477 );
xor ( n22479 , n22476 , n22477 );
xor ( n22480 , n22387 , n22444 );
and ( n22481 , n18113 , n18510 );
and ( n22482 , n22480 , n22481 );
xor ( n22483 , n22480 , n22481 );
xor ( n22484 , n22391 , n22442 );
and ( n22485 , n18114 , n18510 );
and ( n22486 , n22484 , n22485 );
xor ( n22487 , n22484 , n22485 );
xor ( n22488 , n22395 , n22440 );
and ( n22489 , n18115 , n18510 );
and ( n22490 , n22488 , n22489 );
xor ( n22491 , n22488 , n22489 );
xor ( n22492 , n22399 , n22438 );
and ( n22493 , n18116 , n18510 );
and ( n22494 , n22492 , n22493 );
xor ( n22495 , n22492 , n22493 );
xor ( n22496 , n22403 , n22436 );
and ( n22497 , n18117 , n18510 );
and ( n22498 , n22496 , n22497 );
xor ( n22499 , n22496 , n22497 );
xor ( n22500 , n22407 , n22434 );
and ( n22501 , n18118 , n18510 );
and ( n22502 , n22500 , n22501 );
xor ( n22503 , n22500 , n22501 );
xor ( n22504 , n22411 , n22432 );
and ( n22505 , n18119 , n18510 );
and ( n22506 , n22504 , n22505 );
xor ( n22507 , n22504 , n22505 );
xor ( n22508 , n22415 , n22430 );
and ( n22509 , n18120 , n18510 );
and ( n22510 , n22508 , n22509 );
xor ( n22511 , n22508 , n22509 );
xor ( n22512 , n22419 , n22428 );
and ( n22513 , n18121 , n18510 );
and ( n22514 , n22512 , n22513 );
xor ( n22515 , n22512 , n22513 );
xor ( n22516 , n22423 , n22426 );
and ( n22517 , n18122 , n18510 );
and ( n22518 , n22516 , n22517 );
and ( n22519 , n22515 , n22518 );
or ( n22520 , n22514 , n22519 );
and ( n22521 , n22511 , n22520 );
or ( n22522 , n22510 , n22521 );
and ( n22523 , n22507 , n22522 );
or ( n22524 , n22506 , n22523 );
and ( n22525 , n22503 , n22524 );
or ( n22526 , n22502 , n22525 );
and ( n22527 , n22499 , n22526 );
or ( n22528 , n22498 , n22527 );
and ( n22529 , n22495 , n22528 );
or ( n22530 , n22494 , n22529 );
and ( n22531 , n22491 , n22530 );
or ( n22532 , n22490 , n22531 );
and ( n22533 , n22487 , n22532 );
or ( n22534 , n22486 , n22533 );
and ( n22535 , n22483 , n22534 );
or ( n22536 , n22482 , n22535 );
and ( n22537 , n22479 , n22536 );
or ( n22538 , n22478 , n22537 );
and ( n22539 , n22475 , n22538 );
or ( n22540 , n22474 , n22539 );
and ( n22541 , n22471 , n22540 );
or ( n22542 , n22470 , n22541 );
and ( n22543 , n22467 , n22542 );
or ( n22544 , n22466 , n22543 );
and ( n22545 , n22463 , n22544 );
or ( n22546 , n22462 , n22545 );
and ( n22547 , n22459 , n22546 );
or ( n22548 , n22458 , n22547 );
and ( n22549 , n18107 , n18508 );
and ( n22550 , n22548 , n22549 );
xor ( n22551 , n22548 , n22549 );
xor ( n22552 , n22459 , n22546 );
and ( n22553 , n18108 , n18508 );
and ( n22554 , n22552 , n22553 );
xor ( n22555 , n22552 , n22553 );
xor ( n22556 , n22463 , n22544 );
and ( n22557 , n18109 , n18508 );
and ( n22558 , n22556 , n22557 );
xor ( n22559 , n22556 , n22557 );
xor ( n22560 , n22467 , n22542 );
and ( n22561 , n18110 , n18508 );
and ( n22562 , n22560 , n22561 );
xor ( n22563 , n22560 , n22561 );
xor ( n22564 , n22471 , n22540 );
and ( n22565 , n18111 , n18508 );
and ( n22566 , n22564 , n22565 );
xor ( n22567 , n22564 , n22565 );
xor ( n22568 , n22475 , n22538 );
and ( n22569 , n18112 , n18508 );
and ( n22570 , n22568 , n22569 );
xor ( n22571 , n22568 , n22569 );
xor ( n22572 , n22479 , n22536 );
and ( n22573 , n18113 , n18508 );
and ( n22574 , n22572 , n22573 );
xor ( n22575 , n22572 , n22573 );
xor ( n22576 , n22483 , n22534 );
and ( n22577 , n18114 , n18508 );
and ( n22578 , n22576 , n22577 );
xor ( n22579 , n22576 , n22577 );
xor ( n22580 , n22487 , n22532 );
and ( n22581 , n18115 , n18508 );
and ( n22582 , n22580 , n22581 );
xor ( n22583 , n22580 , n22581 );
xor ( n22584 , n22491 , n22530 );
and ( n22585 , n18116 , n18508 );
and ( n22586 , n22584 , n22585 );
xor ( n22587 , n22584 , n22585 );
xor ( n22588 , n22495 , n22528 );
and ( n22589 , n18117 , n18508 );
and ( n22590 , n22588 , n22589 );
xor ( n22591 , n22588 , n22589 );
xor ( n22592 , n22499 , n22526 );
and ( n22593 , n18118 , n18508 );
and ( n22594 , n22592 , n22593 );
xor ( n22595 , n22592 , n22593 );
xor ( n22596 , n22503 , n22524 );
and ( n22597 , n18119 , n18508 );
and ( n22598 , n22596 , n22597 );
xor ( n22599 , n22596 , n22597 );
xor ( n22600 , n22507 , n22522 );
and ( n22601 , n18120 , n18508 );
and ( n22602 , n22600 , n22601 );
xor ( n22603 , n22600 , n22601 );
xor ( n22604 , n22511 , n22520 );
and ( n22605 , n18121 , n18508 );
and ( n22606 , n22604 , n22605 );
xor ( n22607 , n22604 , n22605 );
xor ( n22608 , n22515 , n22518 );
and ( n22609 , n18122 , n18508 );
and ( n22610 , n22608 , n22609 );
and ( n22611 , n22607 , n22610 );
or ( n22612 , n22606 , n22611 );
and ( n22613 , n22603 , n22612 );
or ( n22614 , n22602 , n22613 );
and ( n22615 , n22599 , n22614 );
or ( n22616 , n22598 , n22615 );
and ( n22617 , n22595 , n22616 );
or ( n22618 , n22594 , n22617 );
and ( n22619 , n22591 , n22618 );
or ( n22620 , n22590 , n22619 );
and ( n22621 , n22587 , n22620 );
or ( n22622 , n22586 , n22621 );
and ( n22623 , n22583 , n22622 );
or ( n22624 , n22582 , n22623 );
and ( n22625 , n22579 , n22624 );
or ( n22626 , n22578 , n22625 );
and ( n22627 , n22575 , n22626 );
or ( n22628 , n22574 , n22627 );
and ( n22629 , n22571 , n22628 );
or ( n22630 , n22570 , n22629 );
and ( n22631 , n22567 , n22630 );
or ( n22632 , n22566 , n22631 );
and ( n22633 , n22563 , n22632 );
or ( n22634 , n22562 , n22633 );
and ( n22635 , n22559 , n22634 );
or ( n22636 , n22558 , n22635 );
and ( n22637 , n22555 , n22636 );
or ( n22638 , n22554 , n22637 );
and ( n22639 , n22551 , n22638 );
or ( n22640 , n22550 , n22639 );
and ( n22641 , n18107 , n18506 );
and ( n22642 , n22640 , n22641 );
xor ( n22643 , n22640 , n22641 );
xor ( n22644 , n22551 , n22638 );
and ( n22645 , n18108 , n18506 );
and ( n22646 , n22644 , n22645 );
xor ( n22647 , n22644 , n22645 );
xor ( n22648 , n22555 , n22636 );
and ( n22649 , n18109 , n18506 );
and ( n22650 , n22648 , n22649 );
xor ( n22651 , n22648 , n22649 );
xor ( n22652 , n22559 , n22634 );
and ( n22653 , n18110 , n18506 );
and ( n22654 , n22652 , n22653 );
xor ( n22655 , n22652 , n22653 );
xor ( n22656 , n22563 , n22632 );
and ( n22657 , n18111 , n18506 );
and ( n22658 , n22656 , n22657 );
xor ( n22659 , n22656 , n22657 );
xor ( n22660 , n22567 , n22630 );
and ( n22661 , n18112 , n18506 );
and ( n22662 , n22660 , n22661 );
xor ( n22663 , n22660 , n22661 );
xor ( n22664 , n22571 , n22628 );
and ( n22665 , n18113 , n18506 );
and ( n22666 , n22664 , n22665 );
xor ( n22667 , n22664 , n22665 );
xor ( n22668 , n22575 , n22626 );
and ( n22669 , n18114 , n18506 );
and ( n22670 , n22668 , n22669 );
xor ( n22671 , n22668 , n22669 );
xor ( n22672 , n22579 , n22624 );
and ( n22673 , n18115 , n18506 );
and ( n22674 , n22672 , n22673 );
xor ( n22675 , n22672 , n22673 );
xor ( n22676 , n22583 , n22622 );
and ( n22677 , n18116 , n18506 );
and ( n22678 , n22676 , n22677 );
xor ( n22679 , n22676 , n22677 );
xor ( n22680 , n22587 , n22620 );
and ( n22681 , n18117 , n18506 );
and ( n22682 , n22680 , n22681 );
xor ( n22683 , n22680 , n22681 );
xor ( n22684 , n22591 , n22618 );
and ( n22685 , n18118 , n18506 );
and ( n22686 , n22684 , n22685 );
xor ( n22687 , n22684 , n22685 );
xor ( n22688 , n22595 , n22616 );
and ( n22689 , n18119 , n18506 );
and ( n22690 , n22688 , n22689 );
xor ( n22691 , n22688 , n22689 );
xor ( n22692 , n22599 , n22614 );
and ( n22693 , n18120 , n18506 );
and ( n22694 , n22692 , n22693 );
xor ( n22695 , n22692 , n22693 );
xor ( n22696 , n22603 , n22612 );
and ( n22697 , n18121 , n18506 );
and ( n22698 , n22696 , n22697 );
xor ( n22699 , n22696 , n22697 );
xor ( n22700 , n22607 , n22610 );
and ( n22701 , n18122 , n18506 );
and ( n22702 , n22700 , n22701 );
and ( n22703 , n22699 , n22702 );
or ( n22704 , n22698 , n22703 );
and ( n22705 , n22695 , n22704 );
or ( n22706 , n22694 , n22705 );
and ( n22707 , n22691 , n22706 );
or ( n22708 , n22690 , n22707 );
and ( n22709 , n22687 , n22708 );
or ( n22710 , n22686 , n22709 );
and ( n22711 , n22683 , n22710 );
or ( n22712 , n22682 , n22711 );
and ( n22713 , n22679 , n22712 );
or ( n22714 , n22678 , n22713 );
and ( n22715 , n22675 , n22714 );
or ( n22716 , n22674 , n22715 );
and ( n22717 , n22671 , n22716 );
or ( n22718 , n22670 , n22717 );
and ( n22719 , n22667 , n22718 );
or ( n22720 , n22666 , n22719 );
and ( n22721 , n22663 , n22720 );
or ( n22722 , n22662 , n22721 );
and ( n22723 , n22659 , n22722 );
or ( n22724 , n22658 , n22723 );
and ( n22725 , n22655 , n22724 );
or ( n22726 , n22654 , n22725 );
and ( n22727 , n22651 , n22726 );
or ( n22728 , n22650 , n22727 );
and ( n22729 , n22647 , n22728 );
or ( n22730 , n22646 , n22729 );
and ( n22731 , n22643 , n22730 );
or ( n22732 , n22642 , n22731 );
and ( n22733 , n18107 , n18504 );
and ( n22734 , n22732 , n22733 );
xor ( n22735 , n22732 , n22733 );
xor ( n22736 , n22643 , n22730 );
and ( n22737 , n18108 , n18504 );
and ( n22738 , n22736 , n22737 );
xor ( n22739 , n22736 , n22737 );
xor ( n22740 , n22647 , n22728 );
and ( n22741 , n18109 , n18504 );
and ( n22742 , n22740 , n22741 );
xor ( n22743 , n22740 , n22741 );
xor ( n22744 , n22651 , n22726 );
and ( n22745 , n18110 , n18504 );
and ( n22746 , n22744 , n22745 );
xor ( n22747 , n22744 , n22745 );
xor ( n22748 , n22655 , n22724 );
and ( n22749 , n18111 , n18504 );
and ( n22750 , n22748 , n22749 );
xor ( n22751 , n22748 , n22749 );
xor ( n22752 , n22659 , n22722 );
and ( n22753 , n18112 , n18504 );
and ( n22754 , n22752 , n22753 );
xor ( n22755 , n22752 , n22753 );
xor ( n22756 , n22663 , n22720 );
and ( n22757 , n18113 , n18504 );
and ( n22758 , n22756 , n22757 );
xor ( n22759 , n22756 , n22757 );
xor ( n22760 , n22667 , n22718 );
and ( n22761 , n18114 , n18504 );
and ( n22762 , n22760 , n22761 );
xor ( n22763 , n22760 , n22761 );
xor ( n22764 , n22671 , n22716 );
and ( n22765 , n18115 , n18504 );
and ( n22766 , n22764 , n22765 );
xor ( n22767 , n22764 , n22765 );
xor ( n22768 , n22675 , n22714 );
and ( n22769 , n18116 , n18504 );
and ( n22770 , n22768 , n22769 );
xor ( n22771 , n22768 , n22769 );
xor ( n22772 , n22679 , n22712 );
and ( n22773 , n18117 , n18504 );
and ( n22774 , n22772 , n22773 );
xor ( n22775 , n22772 , n22773 );
xor ( n22776 , n22683 , n22710 );
and ( n22777 , n18118 , n18504 );
and ( n22778 , n22776 , n22777 );
xor ( n22779 , n22776 , n22777 );
xor ( n22780 , n22687 , n22708 );
and ( n22781 , n18119 , n18504 );
and ( n22782 , n22780 , n22781 );
xor ( n22783 , n22780 , n22781 );
xor ( n22784 , n22691 , n22706 );
and ( n22785 , n18120 , n18504 );
and ( n22786 , n22784 , n22785 );
xor ( n22787 , n22784 , n22785 );
xor ( n22788 , n22695 , n22704 );
and ( n22789 , n18121 , n18504 );
and ( n22790 , n22788 , n22789 );
xor ( n22791 , n22788 , n22789 );
xor ( n22792 , n22699 , n22702 );
and ( n22793 , n18122 , n18504 );
and ( n22794 , n22792 , n22793 );
and ( n22795 , n22791 , n22794 );
or ( n22796 , n22790 , n22795 );
and ( n22797 , n22787 , n22796 );
or ( n22798 , n22786 , n22797 );
and ( n22799 , n22783 , n22798 );
or ( n22800 , n22782 , n22799 );
and ( n22801 , n22779 , n22800 );
or ( n22802 , n22778 , n22801 );
and ( n22803 , n22775 , n22802 );
or ( n22804 , n22774 , n22803 );
and ( n22805 , n22771 , n22804 );
or ( n22806 , n22770 , n22805 );
and ( n22807 , n22767 , n22806 );
or ( n22808 , n22766 , n22807 );
and ( n22809 , n22763 , n22808 );
or ( n22810 , n22762 , n22809 );
and ( n22811 , n22759 , n22810 );
or ( n22812 , n22758 , n22811 );
and ( n22813 , n22755 , n22812 );
or ( n22814 , n22754 , n22813 );
and ( n22815 , n22751 , n22814 );
or ( n22816 , n22750 , n22815 );
and ( n22817 , n22747 , n22816 );
or ( n22818 , n22746 , n22817 );
and ( n22819 , n22743 , n22818 );
or ( n22820 , n22742 , n22819 );
and ( n22821 , n22739 , n22820 );
or ( n22822 , n22738 , n22821 );
and ( n22823 , n22735 , n22822 );
or ( n22824 , n22734 , n22823 );
and ( n22825 , n18107 , n18502 );
and ( n22826 , n22824 , n22825 );
xor ( n22827 , n22824 , n22825 );
xor ( n22828 , n22735 , n22822 );
and ( n22829 , n18108 , n18502 );
and ( n22830 , n22828 , n22829 );
xor ( n22831 , n22828 , n22829 );
xor ( n22832 , n22739 , n22820 );
and ( n22833 , n18109 , n18502 );
and ( n22834 , n22832 , n22833 );
xor ( n22835 , n22832 , n22833 );
xor ( n22836 , n22743 , n22818 );
and ( n22837 , n18110 , n18502 );
and ( n22838 , n22836 , n22837 );
xor ( n22839 , n22836 , n22837 );
xor ( n22840 , n22747 , n22816 );
and ( n22841 , n18111 , n18502 );
and ( n22842 , n22840 , n22841 );
xor ( n22843 , n22840 , n22841 );
xor ( n22844 , n22751 , n22814 );
and ( n22845 , n18112 , n18502 );
and ( n22846 , n22844 , n22845 );
xor ( n22847 , n22844 , n22845 );
xor ( n22848 , n22755 , n22812 );
and ( n22849 , n18113 , n18502 );
and ( n22850 , n22848 , n22849 );
xor ( n22851 , n22848 , n22849 );
xor ( n22852 , n22759 , n22810 );
and ( n22853 , n18114 , n18502 );
and ( n22854 , n22852 , n22853 );
xor ( n22855 , n22852 , n22853 );
xor ( n22856 , n22763 , n22808 );
and ( n22857 , n18115 , n18502 );
and ( n22858 , n22856 , n22857 );
xor ( n22859 , n22856 , n22857 );
xor ( n22860 , n22767 , n22806 );
and ( n22861 , n18116 , n18502 );
and ( n22862 , n22860 , n22861 );
xor ( n22863 , n22860 , n22861 );
xor ( n22864 , n22771 , n22804 );
and ( n22865 , n18117 , n18502 );
and ( n22866 , n22864 , n22865 );
xor ( n22867 , n22864 , n22865 );
xor ( n22868 , n22775 , n22802 );
and ( n22869 , n18118 , n18502 );
and ( n22870 , n22868 , n22869 );
xor ( n22871 , n22868 , n22869 );
xor ( n22872 , n22779 , n22800 );
and ( n22873 , n18119 , n18502 );
and ( n22874 , n22872 , n22873 );
xor ( n22875 , n22872 , n22873 );
xor ( n22876 , n22783 , n22798 );
and ( n22877 , n18120 , n18502 );
and ( n22878 , n22876 , n22877 );
xor ( n22879 , n22876 , n22877 );
xor ( n22880 , n22787 , n22796 );
and ( n22881 , n18121 , n18502 );
and ( n22882 , n22880 , n22881 );
xor ( n22883 , n22880 , n22881 );
xor ( n22884 , n22791 , n22794 );
and ( n22885 , n18122 , n18502 );
and ( n22886 , n22884 , n22885 );
and ( n22887 , n22883 , n22886 );
or ( n22888 , n22882 , n22887 );
and ( n22889 , n22879 , n22888 );
or ( n22890 , n22878 , n22889 );
and ( n22891 , n22875 , n22890 );
or ( n22892 , n22874 , n22891 );
and ( n22893 , n22871 , n22892 );
or ( n22894 , n22870 , n22893 );
and ( n22895 , n22867 , n22894 );
or ( n22896 , n22866 , n22895 );
and ( n22897 , n22863 , n22896 );
or ( n22898 , n22862 , n22897 );
and ( n22899 , n22859 , n22898 );
or ( n22900 , n22858 , n22899 );
and ( n22901 , n22855 , n22900 );
or ( n22902 , n22854 , n22901 );
and ( n22903 , n22851 , n22902 );
or ( n22904 , n22850 , n22903 );
and ( n22905 , n22847 , n22904 );
or ( n22906 , n22846 , n22905 );
and ( n22907 , n22843 , n22906 );
or ( n22908 , n22842 , n22907 );
and ( n22909 , n22839 , n22908 );
or ( n22910 , n22838 , n22909 );
and ( n22911 , n22835 , n22910 );
or ( n22912 , n22834 , n22911 );
and ( n22913 , n22831 , n22912 );
or ( n22914 , n22830 , n22913 );
and ( n22915 , n22827 , n22914 );
or ( n22916 , n22826 , n22915 );
and ( n22917 , n18107 , n18500 );
and ( n22918 , n22916 , n22917 );
xor ( n22919 , n22916 , n22917 );
xor ( n22920 , n22827 , n22914 );
and ( n22921 , n18108 , n18500 );
and ( n22922 , n22920 , n22921 );
xor ( n22923 , n22920 , n22921 );
xor ( n22924 , n22831 , n22912 );
and ( n22925 , n18109 , n18500 );
and ( n22926 , n22924 , n22925 );
xor ( n22927 , n22924 , n22925 );
xor ( n22928 , n22835 , n22910 );
and ( n22929 , n18110 , n18500 );
and ( n22930 , n22928 , n22929 );
xor ( n22931 , n22928 , n22929 );
xor ( n22932 , n22839 , n22908 );
and ( n22933 , n18111 , n18500 );
and ( n22934 , n22932 , n22933 );
xor ( n22935 , n22932 , n22933 );
xor ( n22936 , n22843 , n22906 );
and ( n22937 , n18112 , n18500 );
and ( n22938 , n22936 , n22937 );
xor ( n22939 , n22936 , n22937 );
xor ( n22940 , n22847 , n22904 );
and ( n22941 , n18113 , n18500 );
and ( n22942 , n22940 , n22941 );
xor ( n22943 , n22940 , n22941 );
xor ( n22944 , n22851 , n22902 );
and ( n22945 , n18114 , n18500 );
and ( n22946 , n22944 , n22945 );
xor ( n22947 , n22944 , n22945 );
xor ( n22948 , n22855 , n22900 );
and ( n22949 , n18115 , n18500 );
and ( n22950 , n22948 , n22949 );
xor ( n22951 , n22948 , n22949 );
xor ( n22952 , n22859 , n22898 );
and ( n22953 , n18116 , n18500 );
and ( n22954 , n22952 , n22953 );
xor ( n22955 , n22952 , n22953 );
xor ( n22956 , n22863 , n22896 );
and ( n22957 , n18117 , n18500 );
and ( n22958 , n22956 , n22957 );
xor ( n22959 , n22956 , n22957 );
xor ( n22960 , n22867 , n22894 );
and ( n22961 , n18118 , n18500 );
and ( n22962 , n22960 , n22961 );
xor ( n22963 , n22960 , n22961 );
xor ( n22964 , n22871 , n22892 );
and ( n22965 , n18119 , n18500 );
and ( n22966 , n22964 , n22965 );
xor ( n22967 , n22964 , n22965 );
xor ( n22968 , n22875 , n22890 );
and ( n22969 , n18120 , n18500 );
and ( n22970 , n22968 , n22969 );
xor ( n22971 , n22968 , n22969 );
xor ( n22972 , n22879 , n22888 );
and ( n22973 , n18121 , n18500 );
and ( n22974 , n22972 , n22973 );
xor ( n22975 , n22972 , n22973 );
xor ( n22976 , n22883 , n22886 );
and ( n22977 , n18122 , n18500 );
and ( n22978 , n22976 , n22977 );
and ( n22979 , n22975 , n22978 );
or ( n22980 , n22974 , n22979 );
and ( n22981 , n22971 , n22980 );
or ( n22982 , n22970 , n22981 );
and ( n22983 , n22967 , n22982 );
or ( n22984 , n22966 , n22983 );
and ( n22985 , n22963 , n22984 );
or ( n22986 , n22962 , n22985 );
and ( n22987 , n22959 , n22986 );
or ( n22988 , n22958 , n22987 );
and ( n22989 , n22955 , n22988 );
or ( n22990 , n22954 , n22989 );
and ( n22991 , n22951 , n22990 );
or ( n22992 , n22950 , n22991 );
and ( n22993 , n22947 , n22992 );
or ( n22994 , n22946 , n22993 );
and ( n22995 , n22943 , n22994 );
or ( n22996 , n22942 , n22995 );
and ( n22997 , n22939 , n22996 );
or ( n22998 , n22938 , n22997 );
and ( n22999 , n22935 , n22998 );
or ( n23000 , n22934 , n22999 );
and ( n23001 , n22931 , n23000 );
or ( n23002 , n22930 , n23001 );
and ( n23003 , n22927 , n23002 );
or ( n23004 , n22926 , n23003 );
and ( n23005 , n22923 , n23004 );
or ( n23006 , n22922 , n23005 );
and ( n23007 , n22919 , n23006 );
or ( n23008 , n22918 , n23007 );
and ( n23009 , n18107 , n18498 );
and ( n23010 , n23008 , n23009 );
xor ( n23011 , n23008 , n23009 );
xor ( n23012 , n22919 , n23006 );
and ( n23013 , n18108 , n18498 );
and ( n23014 , n23012 , n23013 );
xor ( n23015 , n23012 , n23013 );
xor ( n23016 , n22923 , n23004 );
and ( n23017 , n18109 , n18498 );
and ( n23018 , n23016 , n23017 );
xor ( n23019 , n23016 , n23017 );
xor ( n23020 , n22927 , n23002 );
and ( n23021 , n18110 , n18498 );
and ( n23022 , n23020 , n23021 );
xor ( n23023 , n23020 , n23021 );
xor ( n23024 , n22931 , n23000 );
and ( n23025 , n18111 , n18498 );
and ( n23026 , n23024 , n23025 );
xor ( n23027 , n23024 , n23025 );
xor ( n23028 , n22935 , n22998 );
and ( n23029 , n18112 , n18498 );
and ( n23030 , n23028 , n23029 );
xor ( n23031 , n23028 , n23029 );
xor ( n23032 , n22939 , n22996 );
and ( n23033 , n18113 , n18498 );
and ( n23034 , n23032 , n23033 );
xor ( n23035 , n23032 , n23033 );
xor ( n23036 , n22943 , n22994 );
and ( n23037 , n18114 , n18498 );
and ( n23038 , n23036 , n23037 );
xor ( n23039 , n23036 , n23037 );
xor ( n23040 , n22947 , n22992 );
and ( n23041 , n18115 , n18498 );
and ( n23042 , n23040 , n23041 );
xor ( n23043 , n23040 , n23041 );
xor ( n23044 , n22951 , n22990 );
and ( n23045 , n18116 , n18498 );
and ( n23046 , n23044 , n23045 );
xor ( n23047 , n23044 , n23045 );
xor ( n23048 , n22955 , n22988 );
and ( n23049 , n18117 , n18498 );
and ( n23050 , n23048 , n23049 );
xor ( n23051 , n23048 , n23049 );
xor ( n23052 , n22959 , n22986 );
and ( n23053 , n18118 , n18498 );
and ( n23054 , n23052 , n23053 );
xor ( n23055 , n23052 , n23053 );
xor ( n23056 , n22963 , n22984 );
and ( n23057 , n18119 , n18498 );
and ( n23058 , n23056 , n23057 );
xor ( n23059 , n23056 , n23057 );
xor ( n23060 , n22967 , n22982 );
and ( n23061 , n18120 , n18498 );
and ( n23062 , n23060 , n23061 );
xor ( n23063 , n23060 , n23061 );
xor ( n23064 , n22971 , n22980 );
and ( n23065 , n18121 , n18498 );
and ( n23066 , n23064 , n23065 );
xor ( n23067 , n23064 , n23065 );
xor ( n23068 , n22975 , n22978 );
and ( n23069 , n18122 , n18498 );
and ( n23070 , n23068 , n23069 );
and ( n23071 , n23067 , n23070 );
or ( n23072 , n23066 , n23071 );
and ( n23073 , n23063 , n23072 );
or ( n23074 , n23062 , n23073 );
and ( n23075 , n23059 , n23074 );
or ( n23076 , n23058 , n23075 );
and ( n23077 , n23055 , n23076 );
or ( n23078 , n23054 , n23077 );
and ( n23079 , n23051 , n23078 );
or ( n23080 , n23050 , n23079 );
and ( n23081 , n23047 , n23080 );
or ( n23082 , n23046 , n23081 );
and ( n23083 , n23043 , n23082 );
or ( n23084 , n23042 , n23083 );
and ( n23085 , n23039 , n23084 );
or ( n23086 , n23038 , n23085 );
and ( n23087 , n23035 , n23086 );
or ( n23088 , n23034 , n23087 );
and ( n23089 , n23031 , n23088 );
or ( n23090 , n23030 , n23089 );
and ( n23091 , n23027 , n23090 );
or ( n23092 , n23026 , n23091 );
and ( n23093 , n23023 , n23092 );
or ( n23094 , n23022 , n23093 );
and ( n23095 , n23019 , n23094 );
or ( n23096 , n23018 , n23095 );
and ( n23097 , n23015 , n23096 );
or ( n23098 , n23014 , n23097 );
and ( n23099 , n23011 , n23098 );
or ( n23100 , n23010 , n23099 );
and ( n23101 , n18107 , n18496 );
and ( n23102 , n23100 , n23101 );
xor ( n23103 , n23100 , n23101 );
xor ( n23104 , n23011 , n23098 );
and ( n23105 , n18108 , n18496 );
and ( n23106 , n23104 , n23105 );
xor ( n23107 , n23104 , n23105 );
xor ( n23108 , n23015 , n23096 );
and ( n23109 , n18109 , n18496 );
and ( n23110 , n23108 , n23109 );
xor ( n23111 , n23108 , n23109 );
xor ( n23112 , n23019 , n23094 );
and ( n23113 , n18110 , n18496 );
and ( n23114 , n23112 , n23113 );
xor ( n23115 , n23112 , n23113 );
xor ( n23116 , n23023 , n23092 );
and ( n23117 , n18111 , n18496 );
and ( n23118 , n23116 , n23117 );
xor ( n23119 , n23116 , n23117 );
xor ( n23120 , n23027 , n23090 );
and ( n23121 , n18112 , n18496 );
and ( n23122 , n23120 , n23121 );
xor ( n23123 , n23120 , n23121 );
xor ( n23124 , n23031 , n23088 );
and ( n23125 , n18113 , n18496 );
and ( n23126 , n23124 , n23125 );
xor ( n23127 , n23124 , n23125 );
xor ( n23128 , n23035 , n23086 );
and ( n23129 , n18114 , n18496 );
and ( n23130 , n23128 , n23129 );
xor ( n23131 , n23128 , n23129 );
xor ( n23132 , n23039 , n23084 );
and ( n23133 , n18115 , n18496 );
and ( n23134 , n23132 , n23133 );
xor ( n23135 , n23132 , n23133 );
xor ( n23136 , n23043 , n23082 );
and ( n23137 , n18116 , n18496 );
and ( n23138 , n23136 , n23137 );
xor ( n23139 , n23136 , n23137 );
xor ( n23140 , n23047 , n23080 );
and ( n23141 , n18117 , n18496 );
and ( n23142 , n23140 , n23141 );
xor ( n23143 , n23140 , n23141 );
xor ( n23144 , n23051 , n23078 );
and ( n23145 , n18118 , n18496 );
and ( n23146 , n23144 , n23145 );
xor ( n23147 , n23144 , n23145 );
xor ( n23148 , n23055 , n23076 );
and ( n23149 , n18119 , n18496 );
and ( n23150 , n23148 , n23149 );
xor ( n23151 , n23148 , n23149 );
xor ( n23152 , n23059 , n23074 );
and ( n23153 , n18120 , n18496 );
and ( n23154 , n23152 , n23153 );
xor ( n23155 , n23152 , n23153 );
xor ( n23156 , n23063 , n23072 );
and ( n23157 , n18121 , n18496 );
and ( n23158 , n23156 , n23157 );
xor ( n23159 , n23156 , n23157 );
xor ( n23160 , n23067 , n23070 );
and ( n23161 , n18122 , n18496 );
and ( n23162 , n23160 , n23161 );
and ( n23163 , n23159 , n23162 );
or ( n23164 , n23158 , n23163 );
and ( n23165 , n23155 , n23164 );
or ( n23166 , n23154 , n23165 );
and ( n23167 , n23151 , n23166 );
or ( n23168 , n23150 , n23167 );
and ( n23169 , n23147 , n23168 );
or ( n23170 , n23146 , n23169 );
and ( n23171 , n23143 , n23170 );
or ( n23172 , n23142 , n23171 );
and ( n23173 , n23139 , n23172 );
or ( n23174 , n23138 , n23173 );
and ( n23175 , n23135 , n23174 );
or ( n23176 , n23134 , n23175 );
and ( n23177 , n23131 , n23176 );
or ( n23178 , n23130 , n23177 );
and ( n23179 , n23127 , n23178 );
or ( n23180 , n23126 , n23179 );
and ( n23181 , n23123 , n23180 );
or ( n23182 , n23122 , n23181 );
and ( n23183 , n23119 , n23182 );
or ( n23184 , n23118 , n23183 );
and ( n23185 , n23115 , n23184 );
or ( n23186 , n23114 , n23185 );
and ( n23187 , n23111 , n23186 );
or ( n23188 , n23110 , n23187 );
and ( n23189 , n23107 , n23188 );
or ( n23190 , n23106 , n23189 );
and ( n23191 , n23103 , n23190 );
or ( n23192 , n23102 , n23191 );
and ( n23193 , n18107 , n18494 );
and ( n23194 , n23192 , n23193 );
xor ( n23195 , n23192 , n23193 );
xor ( n23196 , n23103 , n23190 );
and ( n23197 , n18108 , n18494 );
and ( n23198 , n23196 , n23197 );
xor ( n23199 , n23196 , n23197 );
xor ( n23200 , n23107 , n23188 );
and ( n23201 , n18109 , n18494 );
and ( n23202 , n23200 , n23201 );
xor ( n23203 , n23200 , n23201 );
xor ( n23204 , n23111 , n23186 );
and ( n23205 , n18110 , n18494 );
and ( n23206 , n23204 , n23205 );
xor ( n23207 , n23204 , n23205 );
xor ( n23208 , n23115 , n23184 );
and ( n23209 , n18111 , n18494 );
and ( n23210 , n23208 , n23209 );
xor ( n23211 , n23208 , n23209 );
xor ( n23212 , n23119 , n23182 );
and ( n23213 , n18112 , n18494 );
and ( n23214 , n23212 , n23213 );
xor ( n23215 , n23212 , n23213 );
xor ( n23216 , n23123 , n23180 );
and ( n23217 , n18113 , n18494 );
and ( n23218 , n23216 , n23217 );
xor ( n23219 , n23216 , n23217 );
xor ( n23220 , n23127 , n23178 );
and ( n23221 , n18114 , n18494 );
and ( n23222 , n23220 , n23221 );
xor ( n23223 , n23220 , n23221 );
xor ( n23224 , n23131 , n23176 );
and ( n23225 , n18115 , n18494 );
and ( n23226 , n23224 , n23225 );
xor ( n23227 , n23224 , n23225 );
xor ( n23228 , n23135 , n23174 );
and ( n23229 , n18116 , n18494 );
and ( n23230 , n23228 , n23229 );
xor ( n23231 , n23228 , n23229 );
xor ( n23232 , n23139 , n23172 );
and ( n23233 , n18117 , n18494 );
and ( n23234 , n23232 , n23233 );
xor ( n23235 , n23232 , n23233 );
xor ( n23236 , n23143 , n23170 );
and ( n23237 , n18118 , n18494 );
and ( n23238 , n23236 , n23237 );
xor ( n23239 , n23236 , n23237 );
xor ( n23240 , n23147 , n23168 );
and ( n23241 , n18119 , n18494 );
and ( n23242 , n23240 , n23241 );
xor ( n23243 , n23240 , n23241 );
xor ( n23244 , n23151 , n23166 );
and ( n23245 , n18120 , n18494 );
and ( n23246 , n23244 , n23245 );
xor ( n23247 , n23244 , n23245 );
xor ( n23248 , n23155 , n23164 );
and ( n23249 , n18121 , n18494 );
and ( n23250 , n23248 , n23249 );
xor ( n23251 , n23248 , n23249 );
xor ( n23252 , n23159 , n23162 );
and ( n23253 , n18122 , n18494 );
and ( n23254 , n23252 , n23253 );
and ( n23255 , n23251 , n23254 );
or ( n23256 , n23250 , n23255 );
and ( n23257 , n23247 , n23256 );
or ( n23258 , n23246 , n23257 );
and ( n23259 , n23243 , n23258 );
or ( n23260 , n23242 , n23259 );
and ( n23261 , n23239 , n23260 );
or ( n23262 , n23238 , n23261 );
and ( n23263 , n23235 , n23262 );
or ( n23264 , n23234 , n23263 );
and ( n23265 , n23231 , n23264 );
or ( n23266 , n23230 , n23265 );
and ( n23267 , n23227 , n23266 );
or ( n23268 , n23226 , n23267 );
and ( n23269 , n23223 , n23268 );
or ( n23270 , n23222 , n23269 );
and ( n23271 , n23219 , n23270 );
or ( n23272 , n23218 , n23271 );
and ( n23273 , n23215 , n23272 );
or ( n23274 , n23214 , n23273 );
and ( n23275 , n23211 , n23274 );
or ( n23276 , n23210 , n23275 );
and ( n23277 , n23207 , n23276 );
or ( n23278 , n23206 , n23277 );
and ( n23279 , n23203 , n23278 );
or ( n23280 , n23202 , n23279 );
and ( n23281 , n23199 , n23280 );
or ( n23282 , n23198 , n23281 );
and ( n23283 , n23195 , n23282 );
or ( n23284 , n23194 , n23283 );
and ( n23285 , n18107 , n18492 );
and ( n23286 , n23284 , n23285 );
xor ( n23287 , n23284 , n23285 );
xor ( n23288 , n23195 , n23282 );
and ( n23289 , n18108 , n18492 );
and ( n23290 , n23288 , n23289 );
xor ( n23291 , n23288 , n23289 );
xor ( n23292 , n23199 , n23280 );
and ( n23293 , n18109 , n18492 );
and ( n23294 , n23292 , n23293 );
xor ( n23295 , n23292 , n23293 );
xor ( n23296 , n23203 , n23278 );
and ( n23297 , n18110 , n18492 );
and ( n23298 , n23296 , n23297 );
xor ( n23299 , n23296 , n23297 );
xor ( n23300 , n23207 , n23276 );
and ( n23301 , n18111 , n18492 );
and ( n23302 , n23300 , n23301 );
xor ( n23303 , n23300 , n23301 );
xor ( n23304 , n23211 , n23274 );
and ( n23305 , n18112 , n18492 );
and ( n23306 , n23304 , n23305 );
xor ( n23307 , n23304 , n23305 );
xor ( n23308 , n23215 , n23272 );
and ( n23309 , n18113 , n18492 );
and ( n23310 , n23308 , n23309 );
xor ( n23311 , n23308 , n23309 );
xor ( n23312 , n23219 , n23270 );
and ( n23313 , n18114 , n18492 );
and ( n23314 , n23312 , n23313 );
xor ( n23315 , n23312 , n23313 );
xor ( n23316 , n23223 , n23268 );
and ( n23317 , n18115 , n18492 );
and ( n23318 , n23316 , n23317 );
xor ( n23319 , n23316 , n23317 );
xor ( n23320 , n23227 , n23266 );
and ( n23321 , n18116 , n18492 );
and ( n23322 , n23320 , n23321 );
xor ( n23323 , n23320 , n23321 );
xor ( n23324 , n23231 , n23264 );
and ( n23325 , n18117 , n18492 );
and ( n23326 , n23324 , n23325 );
xor ( n23327 , n23324 , n23325 );
xor ( n23328 , n23235 , n23262 );
and ( n23329 , n18118 , n18492 );
and ( n23330 , n23328 , n23329 );
xor ( n23331 , n23328 , n23329 );
xor ( n23332 , n23239 , n23260 );
and ( n23333 , n18119 , n18492 );
and ( n23334 , n23332 , n23333 );
xor ( n23335 , n23332 , n23333 );
xor ( n23336 , n23243 , n23258 );
and ( n23337 , n18120 , n18492 );
and ( n23338 , n23336 , n23337 );
xor ( n23339 , n23336 , n23337 );
xor ( n23340 , n23247 , n23256 );
and ( n23341 , n18121 , n18492 );
and ( n23342 , n23340 , n23341 );
xor ( n23343 , n23340 , n23341 );
xor ( n23344 , n23251 , n23254 );
and ( n23345 , n18122 , n18492 );
and ( n23346 , n23344 , n23345 );
and ( n23347 , n23343 , n23346 );
or ( n23348 , n23342 , n23347 );
and ( n23349 , n23339 , n23348 );
or ( n23350 , n23338 , n23349 );
and ( n23351 , n23335 , n23350 );
or ( n23352 , n23334 , n23351 );
and ( n23353 , n23331 , n23352 );
or ( n23354 , n23330 , n23353 );
and ( n23355 , n23327 , n23354 );
or ( n23356 , n23326 , n23355 );
and ( n23357 , n23323 , n23356 );
or ( n23358 , n23322 , n23357 );
and ( n23359 , n23319 , n23358 );
or ( n23360 , n23318 , n23359 );
and ( n23361 , n23315 , n23360 );
or ( n23362 , n23314 , n23361 );
and ( n23363 , n23311 , n23362 );
or ( n23364 , n23310 , n23363 );
and ( n23365 , n23307 , n23364 );
or ( n23366 , n23306 , n23365 );
and ( n23367 , n23303 , n23366 );
or ( n23368 , n23302 , n23367 );
and ( n23369 , n23299 , n23368 );
or ( n23370 , n23298 , n23369 );
and ( n23371 , n23295 , n23370 );
or ( n23372 , n23294 , n23371 );
and ( n23373 , n23291 , n23372 );
or ( n23374 , n23290 , n23373 );
and ( n23375 , n23287 , n23374 );
or ( n23376 , n23286 , n23375 );
and ( n23377 , n18107 , n18490 );
and ( n23378 , n23376 , n23377 );
xor ( n23379 , n23376 , n23377 );
xor ( n23380 , n23287 , n23374 );
and ( n23381 , n18108 , n18490 );
and ( n23382 , n23380 , n23381 );
xor ( n23383 , n23380 , n23381 );
xor ( n23384 , n23291 , n23372 );
and ( n23385 , n18109 , n18490 );
and ( n23386 , n23384 , n23385 );
xor ( n23387 , n23384 , n23385 );
xor ( n23388 , n23295 , n23370 );
and ( n23389 , n18110 , n18490 );
and ( n23390 , n23388 , n23389 );
xor ( n23391 , n23388 , n23389 );
xor ( n23392 , n23299 , n23368 );
and ( n23393 , n18111 , n18490 );
and ( n23394 , n23392 , n23393 );
xor ( n23395 , n23392 , n23393 );
xor ( n23396 , n23303 , n23366 );
and ( n23397 , n18112 , n18490 );
and ( n23398 , n23396 , n23397 );
xor ( n23399 , n23396 , n23397 );
xor ( n23400 , n23307 , n23364 );
and ( n23401 , n18113 , n18490 );
and ( n23402 , n23400 , n23401 );
xor ( n23403 , n23400 , n23401 );
xor ( n23404 , n23311 , n23362 );
and ( n23405 , n18114 , n18490 );
and ( n23406 , n23404 , n23405 );
xor ( n23407 , n23404 , n23405 );
xor ( n23408 , n23315 , n23360 );
and ( n23409 , n18115 , n18490 );
and ( n23410 , n23408 , n23409 );
xor ( n23411 , n23408 , n23409 );
xor ( n23412 , n23319 , n23358 );
and ( n23413 , n18116 , n18490 );
and ( n23414 , n23412 , n23413 );
xor ( n23415 , n23412 , n23413 );
xor ( n23416 , n23323 , n23356 );
and ( n23417 , n18117 , n18490 );
and ( n23418 , n23416 , n23417 );
xor ( n23419 , n23416 , n23417 );
xor ( n23420 , n23327 , n23354 );
and ( n23421 , n18118 , n18490 );
and ( n23422 , n23420 , n23421 );
xor ( n23423 , n23420 , n23421 );
xor ( n23424 , n23331 , n23352 );
and ( n23425 , n18119 , n18490 );
and ( n23426 , n23424 , n23425 );
xor ( n23427 , n23424 , n23425 );
xor ( n23428 , n23335 , n23350 );
and ( n23429 , n18120 , n18490 );
and ( n23430 , n23428 , n23429 );
xor ( n23431 , n23428 , n23429 );
xor ( n23432 , n23339 , n23348 );
and ( n23433 , n18121 , n18490 );
and ( n23434 , n23432 , n23433 );
xor ( n23435 , n23432 , n23433 );
xor ( n23436 , n23343 , n23346 );
and ( n23437 , n18122 , n18490 );
and ( n23438 , n23436 , n23437 );
and ( n23439 , n23435 , n23438 );
or ( n23440 , n23434 , n23439 );
and ( n23441 , n23431 , n23440 );
or ( n23442 , n23430 , n23441 );
and ( n23443 , n23427 , n23442 );
or ( n23444 , n23426 , n23443 );
and ( n23445 , n23423 , n23444 );
or ( n23446 , n23422 , n23445 );
and ( n23447 , n23419 , n23446 );
or ( n23448 , n23418 , n23447 );
and ( n23449 , n23415 , n23448 );
or ( n23450 , n23414 , n23449 );
and ( n23451 , n23411 , n23450 );
or ( n23452 , n23410 , n23451 );
and ( n23453 , n23407 , n23452 );
or ( n23454 , n23406 , n23453 );
and ( n23455 , n23403 , n23454 );
or ( n23456 , n23402 , n23455 );
and ( n23457 , n23399 , n23456 );
or ( n23458 , n23398 , n23457 );
and ( n23459 , n23395 , n23458 );
or ( n23460 , n23394 , n23459 );
and ( n23461 , n23391 , n23460 );
or ( n23462 , n23390 , n23461 );
and ( n23463 , n23387 , n23462 );
or ( n23464 , n23386 , n23463 );
and ( n23465 , n23383 , n23464 );
or ( n23466 , n23382 , n23465 );
and ( n23467 , n23379 , n23466 );
or ( n23468 , n23378 , n23467 );
and ( n23469 , n18107 , n18488 );
and ( n23470 , n23468 , n23469 );
xor ( n23471 , n23468 , n23469 );
xor ( n23472 , n23379 , n23466 );
and ( n23473 , n18108 , n18488 );
and ( n23474 , n23472 , n23473 );
xor ( n23475 , n23472 , n23473 );
xor ( n23476 , n23383 , n23464 );
and ( n23477 , n18109 , n18488 );
and ( n23478 , n23476 , n23477 );
xor ( n23479 , n23476 , n23477 );
xor ( n23480 , n23387 , n23462 );
and ( n23481 , n18110 , n18488 );
and ( n23482 , n23480 , n23481 );
xor ( n23483 , n23480 , n23481 );
xor ( n23484 , n23391 , n23460 );
and ( n23485 , n18111 , n18488 );
and ( n23486 , n23484 , n23485 );
xor ( n23487 , n23484 , n23485 );
xor ( n23488 , n23395 , n23458 );
and ( n23489 , n18112 , n18488 );
and ( n23490 , n23488 , n23489 );
xor ( n23491 , n23488 , n23489 );
xor ( n23492 , n23399 , n23456 );
and ( n23493 , n18113 , n18488 );
and ( n23494 , n23492 , n23493 );
xor ( n23495 , n23492 , n23493 );
xor ( n23496 , n23403 , n23454 );
and ( n23497 , n18114 , n18488 );
and ( n23498 , n23496 , n23497 );
xor ( n23499 , n23496 , n23497 );
xor ( n23500 , n23407 , n23452 );
and ( n23501 , n18115 , n18488 );
and ( n23502 , n23500 , n23501 );
xor ( n23503 , n23500 , n23501 );
xor ( n23504 , n23411 , n23450 );
and ( n23505 , n18116 , n18488 );
and ( n23506 , n23504 , n23505 );
xor ( n23507 , n23504 , n23505 );
xor ( n23508 , n23415 , n23448 );
and ( n23509 , n18117 , n18488 );
and ( n23510 , n23508 , n23509 );
xor ( n23511 , n23508 , n23509 );
xor ( n23512 , n23419 , n23446 );
and ( n23513 , n18118 , n18488 );
and ( n23514 , n23512 , n23513 );
xor ( n23515 , n23512 , n23513 );
xor ( n23516 , n23423 , n23444 );
and ( n23517 , n18119 , n18488 );
and ( n23518 , n23516 , n23517 );
xor ( n23519 , n23516 , n23517 );
xor ( n23520 , n23427 , n23442 );
and ( n23521 , n18120 , n18488 );
and ( n23522 , n23520 , n23521 );
xor ( n23523 , n23520 , n23521 );
xor ( n23524 , n23431 , n23440 );
and ( n23525 , n18121 , n18488 );
and ( n23526 , n23524 , n23525 );
xor ( n23527 , n23524 , n23525 );
xor ( n23528 , n23435 , n23438 );
and ( n23529 , n18122 , n18488 );
and ( n23530 , n23528 , n23529 );
and ( n23531 , n23527 , n23530 );
or ( n23532 , n23526 , n23531 );
and ( n23533 , n23523 , n23532 );
or ( n23534 , n23522 , n23533 );
and ( n23535 , n23519 , n23534 );
or ( n23536 , n23518 , n23535 );
and ( n23537 , n23515 , n23536 );
or ( n23538 , n23514 , n23537 );
and ( n23539 , n23511 , n23538 );
or ( n23540 , n23510 , n23539 );
and ( n23541 , n23507 , n23540 );
or ( n23542 , n23506 , n23541 );
and ( n23543 , n23503 , n23542 );
or ( n23544 , n23502 , n23543 );
and ( n23545 , n23499 , n23544 );
or ( n23546 , n23498 , n23545 );
and ( n23547 , n23495 , n23546 );
or ( n23548 , n23494 , n23547 );
and ( n23549 , n23491 , n23548 );
or ( n23550 , n23490 , n23549 );
and ( n23551 , n23487 , n23550 );
or ( n23552 , n23486 , n23551 );
and ( n23553 , n23483 , n23552 );
or ( n23554 , n23482 , n23553 );
and ( n23555 , n23479 , n23554 );
or ( n23556 , n23478 , n23555 );
and ( n23557 , n23475 , n23556 );
or ( n23558 , n23474 , n23557 );
and ( n23559 , n23471 , n23558 );
or ( n23560 , n23470 , n23559 );
and ( n23561 , n18107 , n18486 );
and ( n23562 , n23560 , n23561 );
xor ( n23563 , n23560 , n23561 );
xor ( n23564 , n23471 , n23558 );
and ( n23565 , n18108 , n18486 );
and ( n23566 , n23564 , n23565 );
xor ( n23567 , n23564 , n23565 );
xor ( n23568 , n23475 , n23556 );
and ( n23569 , n18109 , n18486 );
and ( n23570 , n23568 , n23569 );
xor ( n23571 , n23568 , n23569 );
xor ( n23572 , n23479 , n23554 );
and ( n23573 , n18110 , n18486 );
and ( n23574 , n23572 , n23573 );
xor ( n23575 , n23572 , n23573 );
xor ( n23576 , n23483 , n23552 );
and ( n23577 , n18111 , n18486 );
and ( n23578 , n23576 , n23577 );
xor ( n23579 , n23576 , n23577 );
xor ( n23580 , n23487 , n23550 );
and ( n23581 , n18112 , n18486 );
and ( n23582 , n23580 , n23581 );
xor ( n23583 , n23580 , n23581 );
xor ( n23584 , n23491 , n23548 );
and ( n23585 , n18113 , n18486 );
and ( n23586 , n23584 , n23585 );
xor ( n23587 , n23584 , n23585 );
xor ( n23588 , n23495 , n23546 );
and ( n23589 , n18114 , n18486 );
and ( n23590 , n23588 , n23589 );
xor ( n23591 , n23588 , n23589 );
xor ( n23592 , n23499 , n23544 );
and ( n23593 , n18115 , n18486 );
and ( n23594 , n23592 , n23593 );
xor ( n23595 , n23592 , n23593 );
xor ( n23596 , n23503 , n23542 );
and ( n23597 , n18116 , n18486 );
and ( n23598 , n23596 , n23597 );
xor ( n23599 , n23596 , n23597 );
xor ( n23600 , n23507 , n23540 );
and ( n23601 , n18117 , n18486 );
and ( n23602 , n23600 , n23601 );
xor ( n23603 , n23600 , n23601 );
xor ( n23604 , n23511 , n23538 );
and ( n23605 , n18118 , n18486 );
and ( n23606 , n23604 , n23605 );
xor ( n23607 , n23604 , n23605 );
xor ( n23608 , n23515 , n23536 );
and ( n23609 , n18119 , n18486 );
and ( n23610 , n23608 , n23609 );
xor ( n23611 , n23608 , n23609 );
xor ( n23612 , n23519 , n23534 );
and ( n23613 , n18120 , n18486 );
and ( n23614 , n23612 , n23613 );
xor ( n23615 , n23612 , n23613 );
xor ( n23616 , n23523 , n23532 );
and ( n23617 , n18121 , n18486 );
and ( n23618 , n23616 , n23617 );
xor ( n23619 , n23616 , n23617 );
xor ( n23620 , n23527 , n23530 );
and ( n23621 , n18122 , n18486 );
and ( n23622 , n23620 , n23621 );
and ( n23623 , n23619 , n23622 );
or ( n23624 , n23618 , n23623 );
and ( n23625 , n23615 , n23624 );
or ( n23626 , n23614 , n23625 );
and ( n23627 , n23611 , n23626 );
or ( n23628 , n23610 , n23627 );
and ( n23629 , n23607 , n23628 );
or ( n23630 , n23606 , n23629 );
and ( n23631 , n23603 , n23630 );
or ( n23632 , n23602 , n23631 );
and ( n23633 , n23599 , n23632 );
or ( n23634 , n23598 , n23633 );
and ( n23635 , n23595 , n23634 );
or ( n23636 , n23594 , n23635 );
and ( n23637 , n23591 , n23636 );
or ( n23638 , n23590 , n23637 );
and ( n23639 , n23587 , n23638 );
or ( n23640 , n23586 , n23639 );
and ( n23641 , n23583 , n23640 );
or ( n23642 , n23582 , n23641 );
and ( n23643 , n23579 , n23642 );
or ( n23644 , n23578 , n23643 );
and ( n23645 , n23575 , n23644 );
or ( n23646 , n23574 , n23645 );
and ( n23647 , n23571 , n23646 );
or ( n23648 , n23570 , n23647 );
and ( n23649 , n23567 , n23648 );
or ( n23650 , n23566 , n23649 );
and ( n23651 , n23563 , n23650 );
or ( n23652 , n23562 , n23651 );
and ( n23653 , n18107 , n18484 );
and ( n23654 , n23652 , n23653 );
xor ( n23655 , n23652 , n23653 );
xor ( n23656 , n23563 , n23650 );
and ( n23657 , n18108 , n18484 );
and ( n23658 , n23656 , n23657 );
xor ( n23659 , n23656 , n23657 );
xor ( n23660 , n23567 , n23648 );
and ( n23661 , n18109 , n18484 );
and ( n23662 , n23660 , n23661 );
xor ( n23663 , n23660 , n23661 );
xor ( n23664 , n23571 , n23646 );
and ( n23665 , n18110 , n18484 );
and ( n23666 , n23664 , n23665 );
xor ( n23667 , n23664 , n23665 );
xor ( n23668 , n23575 , n23644 );
and ( n23669 , n18111 , n18484 );
and ( n23670 , n23668 , n23669 );
xor ( n23671 , n23668 , n23669 );
xor ( n23672 , n23579 , n23642 );
and ( n23673 , n18112 , n18484 );
and ( n23674 , n23672 , n23673 );
xor ( n23675 , n23672 , n23673 );
xor ( n23676 , n23583 , n23640 );
and ( n23677 , n18113 , n18484 );
and ( n23678 , n23676 , n23677 );
xor ( n23679 , n23676 , n23677 );
xor ( n23680 , n23587 , n23638 );
and ( n23681 , n18114 , n18484 );
and ( n23682 , n23680 , n23681 );
xor ( n23683 , n23680 , n23681 );
xor ( n23684 , n23591 , n23636 );
and ( n23685 , n18115 , n18484 );
and ( n23686 , n23684 , n23685 );
xor ( n23687 , n23684 , n23685 );
xor ( n23688 , n23595 , n23634 );
and ( n23689 , n18116 , n18484 );
and ( n23690 , n23688 , n23689 );
xor ( n23691 , n23688 , n23689 );
xor ( n23692 , n23599 , n23632 );
and ( n23693 , n18117 , n18484 );
and ( n23694 , n23692 , n23693 );
xor ( n23695 , n23692 , n23693 );
xor ( n23696 , n23603 , n23630 );
and ( n23697 , n18118 , n18484 );
and ( n23698 , n23696 , n23697 );
xor ( n23699 , n23696 , n23697 );
xor ( n23700 , n23607 , n23628 );
and ( n23701 , n18119 , n18484 );
and ( n23702 , n23700 , n23701 );
xor ( n23703 , n23700 , n23701 );
xor ( n23704 , n23611 , n23626 );
and ( n23705 , n18120 , n18484 );
and ( n23706 , n23704 , n23705 );
xor ( n23707 , n23704 , n23705 );
xor ( n23708 , n23615 , n23624 );
and ( n23709 , n18121 , n18484 );
and ( n23710 , n23708 , n23709 );
xor ( n23711 , n23708 , n23709 );
xor ( n23712 , n23619 , n23622 );
and ( n23713 , n18122 , n18484 );
and ( n23714 , n23712 , n23713 );
and ( n23715 , n23711 , n23714 );
or ( n23716 , n23710 , n23715 );
and ( n23717 , n23707 , n23716 );
or ( n23718 , n23706 , n23717 );
and ( n23719 , n23703 , n23718 );
or ( n23720 , n23702 , n23719 );
and ( n23721 , n23699 , n23720 );
or ( n23722 , n23698 , n23721 );
and ( n23723 , n23695 , n23722 );
or ( n23724 , n23694 , n23723 );
and ( n23725 , n23691 , n23724 );
or ( n23726 , n23690 , n23725 );
and ( n23727 , n23687 , n23726 );
or ( n23728 , n23686 , n23727 );
and ( n23729 , n23683 , n23728 );
or ( n23730 , n23682 , n23729 );
and ( n23731 , n23679 , n23730 );
or ( n23732 , n23678 , n23731 );
and ( n23733 , n23675 , n23732 );
or ( n23734 , n23674 , n23733 );
and ( n23735 , n23671 , n23734 );
or ( n23736 , n23670 , n23735 );
and ( n23737 , n23667 , n23736 );
or ( n23738 , n23666 , n23737 );
and ( n23739 , n23663 , n23738 );
or ( n23740 , n23662 , n23739 );
and ( n23741 , n23659 , n23740 );
or ( n23742 , n23658 , n23741 );
and ( n23743 , n23655 , n23742 );
or ( n23744 , n23654 , n23743 );
and ( n23745 , n18107 , n18482 );
and ( n23746 , n23744 , n23745 );
xor ( n23747 , n23744 , n23745 );
xor ( n23748 , n23655 , n23742 );
and ( n23749 , n18108 , n18482 );
and ( n23750 , n23748 , n23749 );
xor ( n23751 , n23748 , n23749 );
xor ( n23752 , n23659 , n23740 );
and ( n23753 , n18109 , n18482 );
and ( n23754 , n23752 , n23753 );
xor ( n23755 , n23752 , n23753 );
xor ( n23756 , n23663 , n23738 );
and ( n23757 , n18110 , n18482 );
and ( n23758 , n23756 , n23757 );
xor ( n23759 , n23756 , n23757 );
xor ( n23760 , n23667 , n23736 );
and ( n23761 , n18111 , n18482 );
and ( n23762 , n23760 , n23761 );
xor ( n23763 , n23760 , n23761 );
xor ( n23764 , n23671 , n23734 );
and ( n23765 , n18112 , n18482 );
and ( n23766 , n23764 , n23765 );
xor ( n23767 , n23764 , n23765 );
xor ( n23768 , n23675 , n23732 );
and ( n23769 , n18113 , n18482 );
and ( n23770 , n23768 , n23769 );
xor ( n23771 , n23768 , n23769 );
xor ( n23772 , n23679 , n23730 );
and ( n23773 , n18114 , n18482 );
and ( n23774 , n23772 , n23773 );
xor ( n23775 , n23772 , n23773 );
xor ( n23776 , n23683 , n23728 );
and ( n23777 , n18115 , n18482 );
and ( n23778 , n23776 , n23777 );
xor ( n23779 , n23776 , n23777 );
xor ( n23780 , n23687 , n23726 );
and ( n23781 , n18116 , n18482 );
and ( n23782 , n23780 , n23781 );
xor ( n23783 , n23780 , n23781 );
xor ( n23784 , n23691 , n23724 );
and ( n23785 , n18117 , n18482 );
and ( n23786 , n23784 , n23785 );
xor ( n23787 , n23784 , n23785 );
xor ( n23788 , n23695 , n23722 );
and ( n23789 , n18118 , n18482 );
and ( n23790 , n23788 , n23789 );
xor ( n23791 , n23788 , n23789 );
xor ( n23792 , n23699 , n23720 );
and ( n23793 , n18119 , n18482 );
and ( n23794 , n23792 , n23793 );
xor ( n23795 , n23792 , n23793 );
xor ( n23796 , n23703 , n23718 );
and ( n23797 , n18120 , n18482 );
and ( n23798 , n23796 , n23797 );
xor ( n23799 , n23796 , n23797 );
xor ( n23800 , n23707 , n23716 );
and ( n23801 , n18121 , n18482 );
and ( n23802 , n23800 , n23801 );
xor ( n23803 , n23800 , n23801 );
xor ( n23804 , n23711 , n23714 );
and ( n23805 , n18122 , n18482 );
and ( n23806 , n23804 , n23805 );
and ( n23807 , n23803 , n23806 );
or ( n23808 , n23802 , n23807 );
and ( n23809 , n23799 , n23808 );
or ( n23810 , n23798 , n23809 );
and ( n23811 , n23795 , n23810 );
or ( n23812 , n23794 , n23811 );
and ( n23813 , n23791 , n23812 );
or ( n23814 , n23790 , n23813 );
and ( n23815 , n23787 , n23814 );
or ( n23816 , n23786 , n23815 );
and ( n23817 , n23783 , n23816 );
or ( n23818 , n23782 , n23817 );
and ( n23819 , n23779 , n23818 );
or ( n23820 , n23778 , n23819 );
and ( n23821 , n23775 , n23820 );
or ( n23822 , n23774 , n23821 );
and ( n23823 , n23771 , n23822 );
or ( n23824 , n23770 , n23823 );
and ( n23825 , n23767 , n23824 );
or ( n23826 , n23766 , n23825 );
and ( n23827 , n23763 , n23826 );
or ( n23828 , n23762 , n23827 );
and ( n23829 , n23759 , n23828 );
or ( n23830 , n23758 , n23829 );
and ( n23831 , n23755 , n23830 );
or ( n23832 , n23754 , n23831 );
and ( n23833 , n23751 , n23832 );
or ( n23834 , n23750 , n23833 );
and ( n23835 , n23747 , n23834 );
or ( n23836 , n23746 , n23835 );
and ( n23837 , n18107 , n18480 );
and ( n23838 , n23836 , n23837 );
xor ( n23839 , n23836 , n23837 );
xor ( n23840 , n23747 , n23834 );
and ( n23841 , n18108 , n18480 );
and ( n23842 , n23840 , n23841 );
xor ( n23843 , n23840 , n23841 );
xor ( n23844 , n23751 , n23832 );
and ( n23845 , n18109 , n18480 );
and ( n23846 , n23844 , n23845 );
xor ( n23847 , n23844 , n23845 );
xor ( n23848 , n23755 , n23830 );
and ( n23849 , n18110 , n18480 );
and ( n23850 , n23848 , n23849 );
xor ( n23851 , n23848 , n23849 );
xor ( n23852 , n23759 , n23828 );
and ( n23853 , n18111 , n18480 );
and ( n23854 , n23852 , n23853 );
xor ( n23855 , n23852 , n23853 );
xor ( n23856 , n23763 , n23826 );
and ( n23857 , n18112 , n18480 );
and ( n23858 , n23856 , n23857 );
xor ( n23859 , n23856 , n23857 );
xor ( n23860 , n23767 , n23824 );
and ( n23861 , n18113 , n18480 );
and ( n23862 , n23860 , n23861 );
xor ( n23863 , n23860 , n23861 );
xor ( n23864 , n23771 , n23822 );
and ( n23865 , n18114 , n18480 );
and ( n23866 , n23864 , n23865 );
xor ( n23867 , n23864 , n23865 );
xor ( n23868 , n23775 , n23820 );
and ( n23869 , n18115 , n18480 );
and ( n23870 , n23868 , n23869 );
xor ( n23871 , n23868 , n23869 );
xor ( n23872 , n23779 , n23818 );
and ( n23873 , n18116 , n18480 );
and ( n23874 , n23872 , n23873 );
xor ( n23875 , n23872 , n23873 );
xor ( n23876 , n23783 , n23816 );
and ( n23877 , n18117 , n18480 );
and ( n23878 , n23876 , n23877 );
xor ( n23879 , n23876 , n23877 );
xor ( n23880 , n23787 , n23814 );
and ( n23881 , n18118 , n18480 );
and ( n23882 , n23880 , n23881 );
xor ( n23883 , n23880 , n23881 );
xor ( n23884 , n23791 , n23812 );
and ( n23885 , n18119 , n18480 );
and ( n23886 , n23884 , n23885 );
xor ( n23887 , n23884 , n23885 );
xor ( n23888 , n23795 , n23810 );
and ( n23889 , n18120 , n18480 );
and ( n23890 , n23888 , n23889 );
xor ( n23891 , n23888 , n23889 );
xor ( n23892 , n23799 , n23808 );
and ( n23893 , n18121 , n18480 );
and ( n23894 , n23892 , n23893 );
xor ( n23895 , n23892 , n23893 );
xor ( n23896 , n23803 , n23806 );
and ( n23897 , n18122 , n18480 );
and ( n23898 , n23896 , n23897 );
and ( n23899 , n23895 , n23898 );
or ( n23900 , n23894 , n23899 );
and ( n23901 , n23891 , n23900 );
or ( n23902 , n23890 , n23901 );
and ( n23903 , n23887 , n23902 );
or ( n23904 , n23886 , n23903 );
and ( n23905 , n23883 , n23904 );
or ( n23906 , n23882 , n23905 );
and ( n23907 , n23879 , n23906 );
or ( n23908 , n23878 , n23907 );
and ( n23909 , n23875 , n23908 );
or ( n23910 , n23874 , n23909 );
and ( n23911 , n23871 , n23910 );
or ( n23912 , n23870 , n23911 );
and ( n23913 , n23867 , n23912 );
or ( n23914 , n23866 , n23913 );
and ( n23915 , n23863 , n23914 );
or ( n23916 , n23862 , n23915 );
and ( n23917 , n23859 , n23916 );
or ( n23918 , n23858 , n23917 );
and ( n23919 , n23855 , n23918 );
or ( n23920 , n23854 , n23919 );
and ( n23921 , n23851 , n23920 );
or ( n23922 , n23850 , n23921 );
and ( n23923 , n23847 , n23922 );
or ( n23924 , n23846 , n23923 );
and ( n23925 , n23843 , n23924 );
or ( n23926 , n23842 , n23925 );
and ( n23927 , n23839 , n23926 );
or ( n23928 , n23838 , n23927 );
and ( n23929 , n18107 , n18478 );
and ( n23930 , n23928 , n23929 );
xor ( n23931 , n23928 , n23929 );
xor ( n23932 , n23839 , n23926 );
and ( n23933 , n18108 , n18478 );
and ( n23934 , n23932 , n23933 );
xor ( n23935 , n23932 , n23933 );
xor ( n23936 , n23843 , n23924 );
and ( n23937 , n18109 , n18478 );
and ( n23938 , n23936 , n23937 );
xor ( n23939 , n23936 , n23937 );
xor ( n23940 , n23847 , n23922 );
and ( n23941 , n18110 , n18478 );
and ( n23942 , n23940 , n23941 );
xor ( n23943 , n23940 , n23941 );
xor ( n23944 , n23851 , n23920 );
and ( n23945 , n18111 , n18478 );
and ( n23946 , n23944 , n23945 );
xor ( n23947 , n23944 , n23945 );
xor ( n23948 , n23855 , n23918 );
and ( n23949 , n18112 , n18478 );
and ( n23950 , n23948 , n23949 );
xor ( n23951 , n23948 , n23949 );
xor ( n23952 , n23859 , n23916 );
and ( n23953 , n18113 , n18478 );
and ( n23954 , n23952 , n23953 );
xor ( n23955 , n23952 , n23953 );
xor ( n23956 , n23863 , n23914 );
and ( n23957 , n18114 , n18478 );
and ( n23958 , n23956 , n23957 );
xor ( n23959 , n23956 , n23957 );
xor ( n23960 , n23867 , n23912 );
and ( n23961 , n18115 , n18478 );
and ( n23962 , n23960 , n23961 );
xor ( n23963 , n23960 , n23961 );
xor ( n23964 , n23871 , n23910 );
and ( n23965 , n18116 , n18478 );
and ( n23966 , n23964 , n23965 );
xor ( n23967 , n23964 , n23965 );
xor ( n23968 , n23875 , n23908 );
and ( n23969 , n18117 , n18478 );
and ( n23970 , n23968 , n23969 );
xor ( n23971 , n23968 , n23969 );
xor ( n23972 , n23879 , n23906 );
and ( n23973 , n18118 , n18478 );
and ( n23974 , n23972 , n23973 );
xor ( n23975 , n23972 , n23973 );
xor ( n23976 , n23883 , n23904 );
and ( n23977 , n18119 , n18478 );
and ( n23978 , n23976 , n23977 );
xor ( n23979 , n23976 , n23977 );
xor ( n23980 , n23887 , n23902 );
and ( n23981 , n18120 , n18478 );
and ( n23982 , n23980 , n23981 );
xor ( n23983 , n23980 , n23981 );
xor ( n23984 , n23891 , n23900 );
and ( n23985 , n18121 , n18478 );
and ( n23986 , n23984 , n23985 );
xor ( n23987 , n23984 , n23985 );
xor ( n23988 , n23895 , n23898 );
and ( n23989 , n18122 , n18478 );
and ( n23990 , n23988 , n23989 );
and ( n23991 , n23987 , n23990 );
or ( n23992 , n23986 , n23991 );
and ( n23993 , n23983 , n23992 );
or ( n23994 , n23982 , n23993 );
and ( n23995 , n23979 , n23994 );
or ( n23996 , n23978 , n23995 );
and ( n23997 , n23975 , n23996 );
or ( n23998 , n23974 , n23997 );
and ( n23999 , n23971 , n23998 );
or ( n24000 , n23970 , n23999 );
and ( n24001 , n23967 , n24000 );
or ( n24002 , n23966 , n24001 );
and ( n24003 , n23963 , n24002 );
or ( n24004 , n23962 , n24003 );
and ( n24005 , n23959 , n24004 );
or ( n24006 , n23958 , n24005 );
and ( n24007 , n23955 , n24006 );
or ( n24008 , n23954 , n24007 );
and ( n24009 , n23951 , n24008 );
or ( n24010 , n23950 , n24009 );
and ( n24011 , n23947 , n24010 );
or ( n24012 , n23946 , n24011 );
and ( n24013 , n23943 , n24012 );
or ( n24014 , n23942 , n24013 );
and ( n24015 , n23939 , n24014 );
or ( n24016 , n23938 , n24015 );
and ( n24017 , n23935 , n24016 );
or ( n24018 , n23934 , n24017 );
and ( n24019 , n23931 , n24018 );
or ( n24020 , n23930 , n24019 );
and ( n24021 , n18107 , n18476 );
and ( n24022 , n24020 , n24021 );
xor ( n24023 , n24020 , n24021 );
xor ( n24024 , n23931 , n24018 );
and ( n24025 , n18108 , n18476 );
and ( n24026 , n24024 , n24025 );
xor ( n24027 , n24024 , n24025 );
xor ( n24028 , n23935 , n24016 );
and ( n24029 , n18109 , n18476 );
and ( n24030 , n24028 , n24029 );
xor ( n24031 , n24028 , n24029 );
xor ( n24032 , n23939 , n24014 );
and ( n24033 , n18110 , n18476 );
and ( n24034 , n24032 , n24033 );
xor ( n24035 , n24032 , n24033 );
xor ( n24036 , n23943 , n24012 );
and ( n24037 , n18111 , n18476 );
and ( n24038 , n24036 , n24037 );
xor ( n24039 , n24036 , n24037 );
xor ( n24040 , n23947 , n24010 );
and ( n24041 , n18112 , n18476 );
and ( n24042 , n24040 , n24041 );
xor ( n24043 , n24040 , n24041 );
xor ( n24044 , n23951 , n24008 );
and ( n24045 , n18113 , n18476 );
and ( n24046 , n24044 , n24045 );
xor ( n24047 , n24044 , n24045 );
xor ( n24048 , n23955 , n24006 );
and ( n24049 , n18114 , n18476 );
and ( n24050 , n24048 , n24049 );
xor ( n24051 , n24048 , n24049 );
xor ( n24052 , n23959 , n24004 );
and ( n24053 , n18115 , n18476 );
and ( n24054 , n24052 , n24053 );
xor ( n24055 , n24052 , n24053 );
xor ( n24056 , n23963 , n24002 );
and ( n24057 , n18116 , n18476 );
and ( n24058 , n24056 , n24057 );
xor ( n24059 , n24056 , n24057 );
xor ( n24060 , n23967 , n24000 );
and ( n24061 , n18117 , n18476 );
and ( n24062 , n24060 , n24061 );
xor ( n24063 , n24060 , n24061 );
xor ( n24064 , n23971 , n23998 );
and ( n24065 , n18118 , n18476 );
and ( n24066 , n24064 , n24065 );
xor ( n24067 , n24064 , n24065 );
xor ( n24068 , n23975 , n23996 );
and ( n24069 , n18119 , n18476 );
and ( n24070 , n24068 , n24069 );
xor ( n24071 , n24068 , n24069 );
xor ( n24072 , n23979 , n23994 );
and ( n24073 , n18120 , n18476 );
and ( n24074 , n24072 , n24073 );
xor ( n24075 , n24072 , n24073 );
xor ( n24076 , n23983 , n23992 );
and ( n24077 , n18121 , n18476 );
and ( n24078 , n24076 , n24077 );
xor ( n24079 , n24076 , n24077 );
xor ( n24080 , n23987 , n23990 );
and ( n24081 , n18122 , n18476 );
and ( n24082 , n24080 , n24081 );
and ( n24083 , n24079 , n24082 );
or ( n24084 , n24078 , n24083 );
and ( n24085 , n24075 , n24084 );
or ( n24086 , n24074 , n24085 );
and ( n24087 , n24071 , n24086 );
or ( n24088 , n24070 , n24087 );
and ( n24089 , n24067 , n24088 );
or ( n24090 , n24066 , n24089 );
and ( n24091 , n24063 , n24090 );
or ( n24092 , n24062 , n24091 );
and ( n24093 , n24059 , n24092 );
or ( n24094 , n24058 , n24093 );
and ( n24095 , n24055 , n24094 );
or ( n24096 , n24054 , n24095 );
and ( n24097 , n24051 , n24096 );
or ( n24098 , n24050 , n24097 );
and ( n24099 , n24047 , n24098 );
or ( n24100 , n24046 , n24099 );
and ( n24101 , n24043 , n24100 );
or ( n24102 , n24042 , n24101 );
and ( n24103 , n24039 , n24102 );
or ( n24104 , n24038 , n24103 );
and ( n24105 , n24035 , n24104 );
or ( n24106 , n24034 , n24105 );
and ( n24107 , n24031 , n24106 );
or ( n24108 , n24030 , n24107 );
and ( n24109 , n24027 , n24108 );
or ( n24110 , n24026 , n24109 );
and ( n24111 , n24023 , n24110 );
or ( n24112 , n24022 , n24111 );
and ( n24113 , n18107 , n18474 );
and ( n24114 , n24112 , n24113 );
xor ( n24115 , n24112 , n24113 );
xor ( n24116 , n24023 , n24110 );
and ( n24117 , n18108 , n18474 );
and ( n24118 , n24116 , n24117 );
xor ( n24119 , n24116 , n24117 );
xor ( n24120 , n24027 , n24108 );
and ( n24121 , n18109 , n18474 );
and ( n24122 , n24120 , n24121 );
xor ( n24123 , n24120 , n24121 );
xor ( n24124 , n24031 , n24106 );
and ( n24125 , n18110 , n18474 );
and ( n24126 , n24124 , n24125 );
xor ( n24127 , n24124 , n24125 );
xor ( n24128 , n24035 , n24104 );
and ( n24129 , n18111 , n18474 );
and ( n24130 , n24128 , n24129 );
xor ( n24131 , n24128 , n24129 );
xor ( n24132 , n24039 , n24102 );
and ( n24133 , n18112 , n18474 );
and ( n24134 , n24132 , n24133 );
xor ( n24135 , n24132 , n24133 );
xor ( n24136 , n24043 , n24100 );
and ( n24137 , n18113 , n18474 );
and ( n24138 , n24136 , n24137 );
xor ( n24139 , n24136 , n24137 );
xor ( n24140 , n24047 , n24098 );
and ( n24141 , n18114 , n18474 );
and ( n24142 , n24140 , n24141 );
xor ( n24143 , n24140 , n24141 );
xor ( n24144 , n24051 , n24096 );
and ( n24145 , n18115 , n18474 );
and ( n24146 , n24144 , n24145 );
xor ( n24147 , n24144 , n24145 );
xor ( n24148 , n24055 , n24094 );
and ( n24149 , n18116 , n18474 );
and ( n24150 , n24148 , n24149 );
xor ( n24151 , n24148 , n24149 );
xor ( n24152 , n24059 , n24092 );
and ( n24153 , n18117 , n18474 );
and ( n24154 , n24152 , n24153 );
xor ( n24155 , n24152 , n24153 );
xor ( n24156 , n24063 , n24090 );
and ( n24157 , n18118 , n18474 );
and ( n24158 , n24156 , n24157 );
xor ( n24159 , n24156 , n24157 );
xor ( n24160 , n24067 , n24088 );
and ( n24161 , n18119 , n18474 );
and ( n24162 , n24160 , n24161 );
xor ( n24163 , n24160 , n24161 );
xor ( n24164 , n24071 , n24086 );
and ( n24165 , n18120 , n18474 );
and ( n24166 , n24164 , n24165 );
xor ( n24167 , n24164 , n24165 );
xor ( n24168 , n24075 , n24084 );
and ( n24169 , n18121 , n18474 );
and ( n24170 , n24168 , n24169 );
xor ( n24171 , n24168 , n24169 );
xor ( n24172 , n24079 , n24082 );
and ( n24173 , n18122 , n18474 );
and ( n24174 , n24172 , n24173 );
and ( n24175 , n24171 , n24174 );
or ( n24176 , n24170 , n24175 );
and ( n24177 , n24167 , n24176 );
or ( n24178 , n24166 , n24177 );
and ( n24179 , n24163 , n24178 );
or ( n24180 , n24162 , n24179 );
and ( n24181 , n24159 , n24180 );
or ( n24182 , n24158 , n24181 );
and ( n24183 , n24155 , n24182 );
or ( n24184 , n24154 , n24183 );
and ( n24185 , n24151 , n24184 );
or ( n24186 , n24150 , n24185 );
and ( n24187 , n24147 , n24186 );
or ( n24188 , n24146 , n24187 );
and ( n24189 , n24143 , n24188 );
or ( n24190 , n24142 , n24189 );
and ( n24191 , n24139 , n24190 );
or ( n24192 , n24138 , n24191 );
and ( n24193 , n24135 , n24192 );
or ( n24194 , n24134 , n24193 );
and ( n24195 , n24131 , n24194 );
or ( n24196 , n24130 , n24195 );
and ( n24197 , n24127 , n24196 );
or ( n24198 , n24126 , n24197 );
and ( n24199 , n24123 , n24198 );
or ( n24200 , n24122 , n24199 );
and ( n24201 , n24119 , n24200 );
or ( n24202 , n24118 , n24201 );
and ( n24203 , n24115 , n24202 );
or ( n24204 , n24114 , n24203 );
and ( n24205 , n18107 , n18472 );
and ( n24206 , n24204 , n24205 );
xor ( n24207 , n24204 , n24205 );
xor ( n24208 , n24115 , n24202 );
and ( n24209 , n18108 , n18472 );
and ( n24210 , n24208 , n24209 );
xor ( n24211 , n24208 , n24209 );
xor ( n24212 , n24119 , n24200 );
and ( n24213 , n18109 , n18472 );
and ( n24214 , n24212 , n24213 );
xor ( n24215 , n24212 , n24213 );
xor ( n24216 , n24123 , n24198 );
and ( n24217 , n18110 , n18472 );
and ( n24218 , n24216 , n24217 );
xor ( n24219 , n24216 , n24217 );
xor ( n24220 , n24127 , n24196 );
and ( n24221 , n18111 , n18472 );
and ( n24222 , n24220 , n24221 );
xor ( n24223 , n24220 , n24221 );
xor ( n24224 , n24131 , n24194 );
and ( n24225 , n18112 , n18472 );
and ( n24226 , n24224 , n24225 );
xor ( n24227 , n24224 , n24225 );
xor ( n24228 , n24135 , n24192 );
and ( n24229 , n18113 , n18472 );
and ( n24230 , n24228 , n24229 );
xor ( n24231 , n24228 , n24229 );
xor ( n24232 , n24139 , n24190 );
and ( n24233 , n18114 , n18472 );
and ( n24234 , n24232 , n24233 );
xor ( n24235 , n24232 , n24233 );
xor ( n24236 , n24143 , n24188 );
and ( n24237 , n18115 , n18472 );
and ( n24238 , n24236 , n24237 );
xor ( n24239 , n24236 , n24237 );
xor ( n24240 , n24147 , n24186 );
and ( n24241 , n18116 , n18472 );
and ( n24242 , n24240 , n24241 );
xor ( n24243 , n24240 , n24241 );
xor ( n24244 , n24151 , n24184 );
and ( n24245 , n18117 , n18472 );
and ( n24246 , n24244 , n24245 );
xor ( n24247 , n24244 , n24245 );
xor ( n24248 , n24155 , n24182 );
and ( n24249 , n18118 , n18472 );
and ( n24250 , n24248 , n24249 );
xor ( n24251 , n24248 , n24249 );
xor ( n24252 , n24159 , n24180 );
and ( n24253 , n18119 , n18472 );
and ( n24254 , n24252 , n24253 );
xor ( n24255 , n24252 , n24253 );
xor ( n24256 , n24163 , n24178 );
and ( n24257 , n18120 , n18472 );
and ( n24258 , n24256 , n24257 );
xor ( n24259 , n24256 , n24257 );
xor ( n24260 , n24167 , n24176 );
and ( n24261 , n18121 , n18472 );
and ( n24262 , n24260 , n24261 );
xor ( n24263 , n24260 , n24261 );
xor ( n24264 , n24171 , n24174 );
and ( n24265 , n18122 , n18472 );
and ( n24266 , n24264 , n24265 );
and ( n24267 , n24263 , n24266 );
or ( n24268 , n24262 , n24267 );
and ( n24269 , n24259 , n24268 );
or ( n24270 , n24258 , n24269 );
and ( n24271 , n24255 , n24270 );
or ( n24272 , n24254 , n24271 );
and ( n24273 , n24251 , n24272 );
or ( n24274 , n24250 , n24273 );
and ( n24275 , n24247 , n24274 );
or ( n24276 , n24246 , n24275 );
and ( n24277 , n24243 , n24276 );
or ( n24278 , n24242 , n24277 );
and ( n24279 , n24239 , n24278 );
or ( n24280 , n24238 , n24279 );
and ( n24281 , n24235 , n24280 );
or ( n24282 , n24234 , n24281 );
and ( n24283 , n24231 , n24282 );
or ( n24284 , n24230 , n24283 );
and ( n24285 , n24227 , n24284 );
or ( n24286 , n24226 , n24285 );
and ( n24287 , n24223 , n24286 );
or ( n24288 , n24222 , n24287 );
and ( n24289 , n24219 , n24288 );
or ( n24290 , n24218 , n24289 );
and ( n24291 , n24215 , n24290 );
or ( n24292 , n24214 , n24291 );
and ( n24293 , n24211 , n24292 );
or ( n24294 , n24210 , n24293 );
and ( n24295 , n24207 , n24294 );
or ( n24296 , n24206 , n24295 );
and ( n24297 , n18107 , n18470 );
and ( n24298 , n24296 , n24297 );
xor ( n24299 , n24296 , n24297 );
xor ( n24300 , n24207 , n24294 );
and ( n24301 , n18108 , n18470 );
and ( n24302 , n24300 , n24301 );
xor ( n24303 , n24300 , n24301 );
xor ( n24304 , n24211 , n24292 );
and ( n24305 , n18109 , n18470 );
and ( n24306 , n24304 , n24305 );
xor ( n24307 , n24304 , n24305 );
xor ( n24308 , n24215 , n24290 );
and ( n24309 , n18110 , n18470 );
and ( n24310 , n24308 , n24309 );
xor ( n24311 , n24308 , n24309 );
xor ( n24312 , n24219 , n24288 );
and ( n24313 , n18111 , n18470 );
and ( n24314 , n24312 , n24313 );
xor ( n24315 , n24312 , n24313 );
xor ( n24316 , n24223 , n24286 );
and ( n24317 , n18112 , n18470 );
and ( n24318 , n24316 , n24317 );
xor ( n24319 , n24316 , n24317 );
xor ( n24320 , n24227 , n24284 );
and ( n24321 , n18113 , n18470 );
and ( n24322 , n24320 , n24321 );
xor ( n24323 , n24320 , n24321 );
xor ( n24324 , n24231 , n24282 );
and ( n24325 , n18114 , n18470 );
and ( n24326 , n24324 , n24325 );
xor ( n24327 , n24324 , n24325 );
xor ( n24328 , n24235 , n24280 );
and ( n24329 , n18115 , n18470 );
and ( n24330 , n24328 , n24329 );
xor ( n24331 , n24328 , n24329 );
xor ( n24332 , n24239 , n24278 );
and ( n24333 , n18116 , n18470 );
and ( n24334 , n24332 , n24333 );
xor ( n24335 , n24332 , n24333 );
xor ( n24336 , n24243 , n24276 );
and ( n24337 , n18117 , n18470 );
and ( n24338 , n24336 , n24337 );
xor ( n24339 , n24336 , n24337 );
xor ( n24340 , n24247 , n24274 );
and ( n24341 , n18118 , n18470 );
and ( n24342 , n24340 , n24341 );
xor ( n24343 , n24340 , n24341 );
xor ( n24344 , n24251 , n24272 );
and ( n24345 , n18119 , n18470 );
and ( n24346 , n24344 , n24345 );
xor ( n24347 , n24344 , n24345 );
xor ( n24348 , n24255 , n24270 );
and ( n24349 , n18120 , n18470 );
and ( n24350 , n24348 , n24349 );
xor ( n24351 , n24348 , n24349 );
xor ( n24352 , n24259 , n24268 );
and ( n24353 , n18121 , n18470 );
and ( n24354 , n24352 , n24353 );
xor ( n24355 , n24352 , n24353 );
xor ( n24356 , n24263 , n24266 );
and ( n24357 , n18122 , n18470 );
and ( n24358 , n24356 , n24357 );
and ( n24359 , n24355 , n24358 );
or ( n24360 , n24354 , n24359 );
and ( n24361 , n24351 , n24360 );
or ( n24362 , n24350 , n24361 );
and ( n24363 , n24347 , n24362 );
or ( n24364 , n24346 , n24363 );
and ( n24365 , n24343 , n24364 );
or ( n24366 , n24342 , n24365 );
and ( n24367 , n24339 , n24366 );
or ( n24368 , n24338 , n24367 );
and ( n24369 , n24335 , n24368 );
or ( n24370 , n24334 , n24369 );
and ( n24371 , n24331 , n24370 );
or ( n24372 , n24330 , n24371 );
and ( n24373 , n24327 , n24372 );
or ( n24374 , n24326 , n24373 );
and ( n24375 , n24323 , n24374 );
or ( n24376 , n24322 , n24375 );
and ( n24377 , n24319 , n24376 );
or ( n24378 , n24318 , n24377 );
and ( n24379 , n24315 , n24378 );
or ( n24380 , n24314 , n24379 );
and ( n24381 , n24311 , n24380 );
or ( n24382 , n24310 , n24381 );
and ( n24383 , n24307 , n24382 );
or ( n24384 , n24306 , n24383 );
and ( n24385 , n24303 , n24384 );
or ( n24386 , n24302 , n24385 );
and ( n24387 , n24299 , n24386 );
or ( n24388 , n24298 , n24387 );
and ( n24389 , n18107 , n18468 );
and ( n24390 , n24388 , n24389 );
xor ( n24391 , n24388 , n24389 );
xor ( n24392 , n24299 , n24386 );
and ( n24393 , n18108 , n18468 );
and ( n24394 , n24392 , n24393 );
xor ( n24395 , n24392 , n24393 );
xor ( n24396 , n24303 , n24384 );
and ( n24397 , n18109 , n18468 );
and ( n24398 , n24396 , n24397 );
xor ( n24399 , n24396 , n24397 );
xor ( n24400 , n24307 , n24382 );
and ( n24401 , n18110 , n18468 );
and ( n24402 , n24400 , n24401 );
xor ( n24403 , n24400 , n24401 );
xor ( n24404 , n24311 , n24380 );
and ( n24405 , n18111 , n18468 );
and ( n24406 , n24404 , n24405 );
xor ( n24407 , n24404 , n24405 );
xor ( n24408 , n24315 , n24378 );
and ( n24409 , n18112 , n18468 );
and ( n24410 , n24408 , n24409 );
xor ( n24411 , n24408 , n24409 );
xor ( n24412 , n24319 , n24376 );
and ( n24413 , n18113 , n18468 );
and ( n24414 , n24412 , n24413 );
xor ( n24415 , n24412 , n24413 );
xor ( n24416 , n24323 , n24374 );
and ( n24417 , n18114 , n18468 );
and ( n24418 , n24416 , n24417 );
xor ( n24419 , n24416 , n24417 );
xor ( n24420 , n24327 , n24372 );
and ( n24421 , n18115 , n18468 );
and ( n24422 , n24420 , n24421 );
xor ( n24423 , n24420 , n24421 );
xor ( n24424 , n24331 , n24370 );
and ( n24425 , n18116 , n18468 );
and ( n24426 , n24424 , n24425 );
xor ( n24427 , n24424 , n24425 );
xor ( n24428 , n24335 , n24368 );
and ( n24429 , n18117 , n18468 );
and ( n24430 , n24428 , n24429 );
xor ( n24431 , n24428 , n24429 );
xor ( n24432 , n24339 , n24366 );
and ( n24433 , n18118 , n18468 );
and ( n24434 , n24432 , n24433 );
xor ( n24435 , n24432 , n24433 );
xor ( n24436 , n24343 , n24364 );
and ( n24437 , n18119 , n18468 );
and ( n24438 , n24436 , n24437 );
xor ( n24439 , n24436 , n24437 );
xor ( n24440 , n24347 , n24362 );
and ( n24441 , n18120 , n18468 );
and ( n24442 , n24440 , n24441 );
xor ( n24443 , n24440 , n24441 );
xor ( n24444 , n24351 , n24360 );
and ( n24445 , n18121 , n18468 );
and ( n24446 , n24444 , n24445 );
xor ( n24447 , n24444 , n24445 );
xor ( n24448 , n24355 , n24358 );
and ( n24449 , n18122 , n18468 );
and ( n24450 , n24448 , n24449 );
and ( n24451 , n24447 , n24450 );
or ( n24452 , n24446 , n24451 );
and ( n24453 , n24443 , n24452 );
or ( n24454 , n24442 , n24453 );
and ( n24455 , n24439 , n24454 );
or ( n24456 , n24438 , n24455 );
and ( n24457 , n24435 , n24456 );
or ( n24458 , n24434 , n24457 );
and ( n24459 , n24431 , n24458 );
or ( n24460 , n24430 , n24459 );
and ( n24461 , n24427 , n24460 );
or ( n24462 , n24426 , n24461 );
and ( n24463 , n24423 , n24462 );
or ( n24464 , n24422 , n24463 );
and ( n24465 , n24419 , n24464 );
or ( n24466 , n24418 , n24465 );
and ( n24467 , n24415 , n24466 );
or ( n24468 , n24414 , n24467 );
and ( n24469 , n24411 , n24468 );
or ( n24470 , n24410 , n24469 );
and ( n24471 , n24407 , n24470 );
or ( n24472 , n24406 , n24471 );
and ( n24473 , n24403 , n24472 );
or ( n24474 , n24402 , n24473 );
and ( n24475 , n24399 , n24474 );
or ( n24476 , n24398 , n24475 );
and ( n24477 , n24395 , n24476 );
or ( n24478 , n24394 , n24477 );
and ( n24479 , n24391 , n24478 );
or ( n24480 , n24390 , n24479 );
and ( n24481 , n18107 , n18466 );
and ( n24482 , n24480 , n24481 );
xor ( n24483 , n24480 , n24481 );
xor ( n24484 , n24391 , n24478 );
and ( n24485 , n18108 , n18466 );
and ( n24486 , n24484 , n24485 );
xor ( n24487 , n24484 , n24485 );
xor ( n24488 , n24395 , n24476 );
and ( n24489 , n18109 , n18466 );
and ( n24490 , n24488 , n24489 );
xor ( n24491 , n24488 , n24489 );
xor ( n24492 , n24399 , n24474 );
and ( n24493 , n18110 , n18466 );
and ( n24494 , n24492 , n24493 );
xor ( n24495 , n24492 , n24493 );
xor ( n24496 , n24403 , n24472 );
and ( n24497 , n18111 , n18466 );
and ( n24498 , n24496 , n24497 );
xor ( n24499 , n24496 , n24497 );
xor ( n24500 , n24407 , n24470 );
and ( n24501 , n18112 , n18466 );
and ( n24502 , n24500 , n24501 );
xor ( n24503 , n24500 , n24501 );
xor ( n24504 , n24411 , n24468 );
and ( n24505 , n18113 , n18466 );
and ( n24506 , n24504 , n24505 );
xor ( n24507 , n24504 , n24505 );
xor ( n24508 , n24415 , n24466 );
and ( n24509 , n18114 , n18466 );
and ( n24510 , n24508 , n24509 );
xor ( n24511 , n24508 , n24509 );
xor ( n24512 , n24419 , n24464 );
and ( n24513 , n18115 , n18466 );
and ( n24514 , n24512 , n24513 );
xor ( n24515 , n24512 , n24513 );
xor ( n24516 , n24423 , n24462 );
and ( n24517 , n18116 , n18466 );
and ( n24518 , n24516 , n24517 );
xor ( n24519 , n24516 , n24517 );
xor ( n24520 , n24427 , n24460 );
and ( n24521 , n18117 , n18466 );
and ( n24522 , n24520 , n24521 );
xor ( n24523 , n24520 , n24521 );
xor ( n24524 , n24431 , n24458 );
and ( n24525 , n18118 , n18466 );
and ( n24526 , n24524 , n24525 );
xor ( n24527 , n24524 , n24525 );
xor ( n24528 , n24435 , n24456 );
and ( n24529 , n18119 , n18466 );
and ( n24530 , n24528 , n24529 );
xor ( n24531 , n24528 , n24529 );
xor ( n24532 , n24439 , n24454 );
and ( n24533 , n18120 , n18466 );
and ( n24534 , n24532 , n24533 );
xor ( n24535 , n24532 , n24533 );
xor ( n24536 , n24443 , n24452 );
and ( n24537 , n18121 , n18466 );
and ( n24538 , n24536 , n24537 );
xor ( n24539 , n24536 , n24537 );
xor ( n24540 , n24447 , n24450 );
and ( n24541 , n18122 , n18466 );
and ( n24542 , n24540 , n24541 );
and ( n24543 , n24539 , n24542 );
or ( n24544 , n24538 , n24543 );
and ( n24545 , n24535 , n24544 );
or ( n24546 , n24534 , n24545 );
and ( n24547 , n24531 , n24546 );
or ( n24548 , n24530 , n24547 );
and ( n24549 , n24527 , n24548 );
or ( n24550 , n24526 , n24549 );
and ( n24551 , n24523 , n24550 );
or ( n24552 , n24522 , n24551 );
and ( n24553 , n24519 , n24552 );
or ( n24554 , n24518 , n24553 );
and ( n24555 , n24515 , n24554 );
or ( n24556 , n24514 , n24555 );
and ( n24557 , n24511 , n24556 );
or ( n24558 , n24510 , n24557 );
and ( n24559 , n24507 , n24558 );
or ( n24560 , n24506 , n24559 );
and ( n24561 , n24503 , n24560 );
or ( n24562 , n24502 , n24561 );
and ( n24563 , n24499 , n24562 );
or ( n24564 , n24498 , n24563 );
and ( n24565 , n24495 , n24564 );
or ( n24566 , n24494 , n24565 );
and ( n24567 , n24491 , n24566 );
or ( n24568 , n24490 , n24567 );
and ( n24569 , n24487 , n24568 );
or ( n24570 , n24486 , n24569 );
and ( n24571 , n24483 , n24570 );
or ( n24572 , n24482 , n24571 );
and ( n24573 , n18107 , n18464 );
and ( n24574 , n24572 , n24573 );
xor ( n24575 , n24572 , n24573 );
xor ( n24576 , n24483 , n24570 );
and ( n24577 , n18108 , n18464 );
and ( n24578 , n24576 , n24577 );
xor ( n24579 , n24576 , n24577 );
xor ( n24580 , n24487 , n24568 );
and ( n24581 , n18109 , n18464 );
and ( n24582 , n24580 , n24581 );
xor ( n24583 , n24580 , n24581 );
xor ( n24584 , n24491 , n24566 );
and ( n24585 , n18110 , n18464 );
and ( n24586 , n24584 , n24585 );
xor ( n24587 , n24584 , n24585 );
xor ( n24588 , n24495 , n24564 );
and ( n24589 , n18111 , n18464 );
and ( n24590 , n24588 , n24589 );
xor ( n24591 , n24588 , n24589 );
xor ( n24592 , n24499 , n24562 );
and ( n24593 , n18112 , n18464 );
and ( n24594 , n24592 , n24593 );
xor ( n24595 , n24592 , n24593 );
xor ( n24596 , n24503 , n24560 );
and ( n24597 , n18113 , n18464 );
and ( n24598 , n24596 , n24597 );
xor ( n24599 , n24596 , n24597 );
xor ( n24600 , n24507 , n24558 );
and ( n24601 , n18114 , n18464 );
and ( n24602 , n24600 , n24601 );
xor ( n24603 , n24600 , n24601 );
xor ( n24604 , n24511 , n24556 );
and ( n24605 , n18115 , n18464 );
and ( n24606 , n24604 , n24605 );
xor ( n24607 , n24604 , n24605 );
xor ( n24608 , n24515 , n24554 );
and ( n24609 , n18116 , n18464 );
and ( n24610 , n24608 , n24609 );
xor ( n24611 , n24608 , n24609 );
xor ( n24612 , n24519 , n24552 );
and ( n24613 , n18117 , n18464 );
and ( n24614 , n24612 , n24613 );
xor ( n24615 , n24612 , n24613 );
xor ( n24616 , n24523 , n24550 );
and ( n24617 , n18118 , n18464 );
and ( n24618 , n24616 , n24617 );
xor ( n24619 , n24616 , n24617 );
xor ( n24620 , n24527 , n24548 );
and ( n24621 , n18119 , n18464 );
and ( n24622 , n24620 , n24621 );
xor ( n24623 , n24620 , n24621 );
xor ( n24624 , n24531 , n24546 );
and ( n24625 , n18120 , n18464 );
and ( n24626 , n24624 , n24625 );
xor ( n24627 , n24624 , n24625 );
xor ( n24628 , n24535 , n24544 );
and ( n24629 , n18121 , n18464 );
and ( n24630 , n24628 , n24629 );
xor ( n24631 , n24628 , n24629 );
xor ( n24632 , n24539 , n24542 );
and ( n24633 , n18122 , n18464 );
and ( n24634 , n24632 , n24633 );
and ( n24635 , n24631 , n24634 );
or ( n24636 , n24630 , n24635 );
and ( n24637 , n24627 , n24636 );
or ( n24638 , n24626 , n24637 );
and ( n24639 , n24623 , n24638 );
or ( n24640 , n24622 , n24639 );
and ( n24641 , n24619 , n24640 );
or ( n24642 , n24618 , n24641 );
and ( n24643 , n24615 , n24642 );
or ( n24644 , n24614 , n24643 );
and ( n24645 , n24611 , n24644 );
or ( n24646 , n24610 , n24645 );
and ( n24647 , n24607 , n24646 );
or ( n24648 , n24606 , n24647 );
and ( n24649 , n24603 , n24648 );
or ( n24650 , n24602 , n24649 );
and ( n24651 , n24599 , n24650 );
or ( n24652 , n24598 , n24651 );
and ( n24653 , n24595 , n24652 );
or ( n24654 , n24594 , n24653 );
and ( n24655 , n24591 , n24654 );
or ( n24656 , n24590 , n24655 );
and ( n24657 , n24587 , n24656 );
or ( n24658 , n24586 , n24657 );
and ( n24659 , n24583 , n24658 );
or ( n24660 , n24582 , n24659 );
and ( n24661 , n24579 , n24660 );
or ( n24662 , n24578 , n24661 );
and ( n24663 , n24575 , n24662 );
or ( n24664 , n24574 , n24663 );
and ( n24665 , n18107 , n18462 );
and ( n24666 , n24664 , n24665 );
xor ( n24667 , n24664 , n24665 );
xor ( n24668 , n24575 , n24662 );
and ( n24669 , n18108 , n18462 );
and ( n24670 , n24668 , n24669 );
xor ( n24671 , n24668 , n24669 );
xor ( n24672 , n24579 , n24660 );
and ( n24673 , n18109 , n18462 );
and ( n24674 , n24672 , n24673 );
xor ( n24675 , n24672 , n24673 );
xor ( n24676 , n24583 , n24658 );
and ( n24677 , n18110 , n18462 );
and ( n24678 , n24676 , n24677 );
xor ( n24679 , n24676 , n24677 );
xor ( n24680 , n24587 , n24656 );
and ( n24681 , n18111 , n18462 );
and ( n24682 , n24680 , n24681 );
xor ( n24683 , n24680 , n24681 );
xor ( n24684 , n24591 , n24654 );
and ( n24685 , n18112 , n18462 );
and ( n24686 , n24684 , n24685 );
xor ( n24687 , n24684 , n24685 );
xor ( n24688 , n24595 , n24652 );
and ( n24689 , n18113 , n18462 );
and ( n24690 , n24688 , n24689 );
xor ( n24691 , n24688 , n24689 );
xor ( n24692 , n24599 , n24650 );
and ( n24693 , n18114 , n18462 );
and ( n24694 , n24692 , n24693 );
xor ( n24695 , n24692 , n24693 );
xor ( n24696 , n24603 , n24648 );
and ( n24697 , n18115 , n18462 );
and ( n24698 , n24696 , n24697 );
xor ( n24699 , n24696 , n24697 );
xor ( n24700 , n24607 , n24646 );
and ( n24701 , n18116 , n18462 );
and ( n24702 , n24700 , n24701 );
xor ( n24703 , n24700 , n24701 );
xor ( n24704 , n24611 , n24644 );
and ( n24705 , n18117 , n18462 );
and ( n24706 , n24704 , n24705 );
xor ( n24707 , n24704 , n24705 );
xor ( n24708 , n24615 , n24642 );
and ( n24709 , n18118 , n18462 );
and ( n24710 , n24708 , n24709 );
xor ( n24711 , n24708 , n24709 );
xor ( n24712 , n24619 , n24640 );
and ( n24713 , n18119 , n18462 );
and ( n24714 , n24712 , n24713 );
xor ( n24715 , n24712 , n24713 );
xor ( n24716 , n24623 , n24638 );
and ( n24717 , n18120 , n18462 );
and ( n24718 , n24716 , n24717 );
xor ( n24719 , n24716 , n24717 );
xor ( n24720 , n24627 , n24636 );
and ( n24721 , n18121 , n18462 );
and ( n24722 , n24720 , n24721 );
xor ( n24723 , n24720 , n24721 );
xor ( n24724 , n24631 , n24634 );
and ( n24725 , n18122 , n18462 );
and ( n24726 , n24724 , n24725 );
and ( n24727 , n24723 , n24726 );
or ( n24728 , n24722 , n24727 );
and ( n24729 , n24719 , n24728 );
or ( n24730 , n24718 , n24729 );
and ( n24731 , n24715 , n24730 );
or ( n24732 , n24714 , n24731 );
and ( n24733 , n24711 , n24732 );
or ( n24734 , n24710 , n24733 );
and ( n24735 , n24707 , n24734 );
or ( n24736 , n24706 , n24735 );
and ( n24737 , n24703 , n24736 );
or ( n24738 , n24702 , n24737 );
and ( n24739 , n24699 , n24738 );
or ( n24740 , n24698 , n24739 );
and ( n24741 , n24695 , n24740 );
or ( n24742 , n24694 , n24741 );
and ( n24743 , n24691 , n24742 );
or ( n24744 , n24690 , n24743 );
and ( n24745 , n24687 , n24744 );
or ( n24746 , n24686 , n24745 );
and ( n24747 , n24683 , n24746 );
or ( n24748 , n24682 , n24747 );
and ( n24749 , n24679 , n24748 );
or ( n24750 , n24678 , n24749 );
and ( n24751 , n24675 , n24750 );
or ( n24752 , n24674 , n24751 );
and ( n24753 , n24671 , n24752 );
or ( n24754 , n24670 , n24753 );
and ( n24755 , n24667 , n24754 );
or ( n24756 , n24666 , n24755 );
and ( n24757 , n18107 , n18460 );
and ( n24758 , n24756 , n24757 );
xor ( n24759 , n24756 , n24757 );
xor ( n24760 , n24667 , n24754 );
and ( n24761 , n18108 , n18460 );
and ( n24762 , n24760 , n24761 );
xor ( n24763 , n24760 , n24761 );
xor ( n24764 , n24671 , n24752 );
and ( n24765 , n18109 , n18460 );
and ( n24766 , n24764 , n24765 );
xor ( n24767 , n24764 , n24765 );
xor ( n24768 , n24675 , n24750 );
and ( n24769 , n18110 , n18460 );
and ( n24770 , n24768 , n24769 );
xor ( n24771 , n24768 , n24769 );
xor ( n24772 , n24679 , n24748 );
and ( n24773 , n18111 , n18460 );
and ( n24774 , n24772 , n24773 );
xor ( n24775 , n24772 , n24773 );
xor ( n24776 , n24683 , n24746 );
and ( n24777 , n18112 , n18460 );
and ( n24778 , n24776 , n24777 );
xor ( n24779 , n24776 , n24777 );
xor ( n24780 , n24687 , n24744 );
and ( n24781 , n18113 , n18460 );
and ( n24782 , n24780 , n24781 );
xor ( n24783 , n24780 , n24781 );
xor ( n24784 , n24691 , n24742 );
and ( n24785 , n18114 , n18460 );
and ( n24786 , n24784 , n24785 );
xor ( n24787 , n24784 , n24785 );
xor ( n24788 , n24695 , n24740 );
and ( n24789 , n18115 , n18460 );
and ( n24790 , n24788 , n24789 );
xor ( n24791 , n24788 , n24789 );
xor ( n24792 , n24699 , n24738 );
and ( n24793 , n18116 , n18460 );
and ( n24794 , n24792 , n24793 );
xor ( n24795 , n24792 , n24793 );
xor ( n24796 , n24703 , n24736 );
and ( n24797 , n18117 , n18460 );
and ( n24798 , n24796 , n24797 );
xor ( n24799 , n24796 , n24797 );
xor ( n24800 , n24707 , n24734 );
and ( n24801 , n18118 , n18460 );
and ( n24802 , n24800 , n24801 );
xor ( n24803 , n24800 , n24801 );
xor ( n24804 , n24711 , n24732 );
and ( n24805 , n18119 , n18460 );
and ( n24806 , n24804 , n24805 );
xor ( n24807 , n24804 , n24805 );
xor ( n24808 , n24715 , n24730 );
and ( n24809 , n18120 , n18460 );
and ( n24810 , n24808 , n24809 );
xor ( n24811 , n24808 , n24809 );
xor ( n24812 , n24719 , n24728 );
and ( n24813 , n18121 , n18460 );
and ( n24814 , n24812 , n24813 );
xor ( n24815 , n24812 , n24813 );
xor ( n24816 , n24723 , n24726 );
and ( n24817 , n18122 , n18460 );
and ( n24818 , n24816 , n24817 );
and ( n24819 , n24815 , n24818 );
or ( n24820 , n24814 , n24819 );
and ( n24821 , n24811 , n24820 );
or ( n24822 , n24810 , n24821 );
and ( n24823 , n24807 , n24822 );
or ( n24824 , n24806 , n24823 );
and ( n24825 , n24803 , n24824 );
or ( n24826 , n24802 , n24825 );
and ( n24827 , n24799 , n24826 );
or ( n24828 , n24798 , n24827 );
and ( n24829 , n24795 , n24828 );
or ( n24830 , n24794 , n24829 );
and ( n24831 , n24791 , n24830 );
or ( n24832 , n24790 , n24831 );
and ( n24833 , n24787 , n24832 );
or ( n24834 , n24786 , n24833 );
and ( n24835 , n24783 , n24834 );
or ( n24836 , n24782 , n24835 );
and ( n24837 , n24779 , n24836 );
or ( n24838 , n24778 , n24837 );
and ( n24839 , n24775 , n24838 );
or ( n24840 , n24774 , n24839 );
and ( n24841 , n24771 , n24840 );
or ( n24842 , n24770 , n24841 );
and ( n24843 , n24767 , n24842 );
or ( n24844 , n24766 , n24843 );
and ( n24845 , n24763 , n24844 );
or ( n24846 , n24762 , n24845 );
and ( n24847 , n24759 , n24846 );
or ( n24848 , n24758 , n24847 );
and ( n24849 , n18107 , n18458 );
and ( n24850 , n24848 , n24849 );
xor ( n24851 , n24848 , n24849 );
xor ( n24852 , n24759 , n24846 );
and ( n24853 , n18108 , n18458 );
and ( n24854 , n24852 , n24853 );
xor ( n24855 , n24852 , n24853 );
xor ( n24856 , n24763 , n24844 );
and ( n24857 , n18109 , n18458 );
and ( n24858 , n24856 , n24857 );
xor ( n24859 , n24856 , n24857 );
xor ( n24860 , n24767 , n24842 );
and ( n24861 , n18110 , n18458 );
and ( n24862 , n24860 , n24861 );
xor ( n24863 , n24860 , n24861 );
xor ( n24864 , n24771 , n24840 );
and ( n24865 , n18111 , n18458 );
and ( n24866 , n24864 , n24865 );
xor ( n24867 , n24864 , n24865 );
xor ( n24868 , n24775 , n24838 );
and ( n24869 , n18112 , n18458 );
and ( n24870 , n24868 , n24869 );
xor ( n24871 , n24868 , n24869 );
xor ( n24872 , n24779 , n24836 );
and ( n24873 , n18113 , n18458 );
and ( n24874 , n24872 , n24873 );
xor ( n24875 , n24872 , n24873 );
xor ( n24876 , n24783 , n24834 );
and ( n24877 , n18114 , n18458 );
and ( n24878 , n24876 , n24877 );
xor ( n24879 , n24876 , n24877 );
xor ( n24880 , n24787 , n24832 );
and ( n24881 , n18115 , n18458 );
and ( n24882 , n24880 , n24881 );
xor ( n24883 , n24880 , n24881 );
xor ( n24884 , n24791 , n24830 );
and ( n24885 , n18116 , n18458 );
and ( n24886 , n24884 , n24885 );
xor ( n24887 , n24884 , n24885 );
xor ( n24888 , n24795 , n24828 );
and ( n24889 , n18117 , n18458 );
and ( n24890 , n24888 , n24889 );
xor ( n24891 , n24888 , n24889 );
xor ( n24892 , n24799 , n24826 );
and ( n24893 , n18118 , n18458 );
and ( n24894 , n24892 , n24893 );
xor ( n24895 , n24892 , n24893 );
xor ( n24896 , n24803 , n24824 );
and ( n24897 , n18119 , n18458 );
and ( n24898 , n24896 , n24897 );
xor ( n24899 , n24896 , n24897 );
xor ( n24900 , n24807 , n24822 );
and ( n24901 , n18120 , n18458 );
and ( n24902 , n24900 , n24901 );
xor ( n24903 , n24900 , n24901 );
xor ( n24904 , n24811 , n24820 );
and ( n24905 , n18121 , n18458 );
and ( n24906 , n24904 , n24905 );
xor ( n24907 , n24904 , n24905 );
xor ( n24908 , n24815 , n24818 );
and ( n24909 , n18122 , n18458 );
and ( n24910 , n24908 , n24909 );
and ( n24911 , n24907 , n24910 );
or ( n24912 , n24906 , n24911 );
and ( n24913 , n24903 , n24912 );
or ( n24914 , n24902 , n24913 );
and ( n24915 , n24899 , n24914 );
or ( n24916 , n24898 , n24915 );
and ( n24917 , n24895 , n24916 );
or ( n24918 , n24894 , n24917 );
and ( n24919 , n24891 , n24918 );
or ( n24920 , n24890 , n24919 );
and ( n24921 , n24887 , n24920 );
or ( n24922 , n24886 , n24921 );
and ( n24923 , n24883 , n24922 );
or ( n24924 , n24882 , n24923 );
and ( n24925 , n24879 , n24924 );
or ( n24926 , n24878 , n24925 );
and ( n24927 , n24875 , n24926 );
or ( n24928 , n24874 , n24927 );
and ( n24929 , n24871 , n24928 );
or ( n24930 , n24870 , n24929 );
and ( n24931 , n24867 , n24930 );
or ( n24932 , n24866 , n24931 );
and ( n24933 , n24863 , n24932 );
or ( n24934 , n24862 , n24933 );
and ( n24935 , n24859 , n24934 );
or ( n24936 , n24858 , n24935 );
and ( n24937 , n24855 , n24936 );
or ( n24938 , n24854 , n24937 );
and ( n24939 , n24851 , n24938 );
or ( n24940 , n24850 , n24939 );
and ( n24941 , n18107 , n18456 );
and ( n24942 , n24940 , n24941 );
xor ( n24943 , n24940 , n24941 );
xor ( n24944 , n24851 , n24938 );
and ( n24945 , n18108 , n18456 );
and ( n24946 , n24944 , n24945 );
xor ( n24947 , n24944 , n24945 );
xor ( n24948 , n24855 , n24936 );
and ( n24949 , n18109 , n18456 );
and ( n24950 , n24948 , n24949 );
xor ( n24951 , n24948 , n24949 );
xor ( n24952 , n24859 , n24934 );
and ( n24953 , n18110 , n18456 );
and ( n24954 , n24952 , n24953 );
xor ( n24955 , n24952 , n24953 );
xor ( n24956 , n24863 , n24932 );
and ( n24957 , n18111 , n18456 );
and ( n24958 , n24956 , n24957 );
xor ( n24959 , n24956 , n24957 );
xor ( n24960 , n24867 , n24930 );
and ( n24961 , n18112 , n18456 );
and ( n24962 , n24960 , n24961 );
xor ( n24963 , n24960 , n24961 );
xor ( n24964 , n24871 , n24928 );
and ( n24965 , n18113 , n18456 );
and ( n24966 , n24964 , n24965 );
xor ( n24967 , n24964 , n24965 );
xor ( n24968 , n24875 , n24926 );
and ( n24969 , n18114 , n18456 );
and ( n24970 , n24968 , n24969 );
xor ( n24971 , n24968 , n24969 );
xor ( n24972 , n24879 , n24924 );
and ( n24973 , n18115 , n18456 );
and ( n24974 , n24972 , n24973 );
xor ( n24975 , n24972 , n24973 );
xor ( n24976 , n24883 , n24922 );
and ( n24977 , n18116 , n18456 );
and ( n24978 , n24976 , n24977 );
xor ( n24979 , n24976 , n24977 );
xor ( n24980 , n24887 , n24920 );
and ( n24981 , n18117 , n18456 );
and ( n24982 , n24980 , n24981 );
xor ( n24983 , n24980 , n24981 );
xor ( n24984 , n24891 , n24918 );
and ( n24985 , n18118 , n18456 );
and ( n24986 , n24984 , n24985 );
xor ( n24987 , n24984 , n24985 );
xor ( n24988 , n24895 , n24916 );
and ( n24989 , n18119 , n18456 );
and ( n24990 , n24988 , n24989 );
xor ( n24991 , n24988 , n24989 );
xor ( n24992 , n24899 , n24914 );
and ( n24993 , n18120 , n18456 );
and ( n24994 , n24992 , n24993 );
xor ( n24995 , n24992 , n24993 );
xor ( n24996 , n24903 , n24912 );
and ( n24997 , n18121 , n18456 );
and ( n24998 , n24996 , n24997 );
xor ( n24999 , n24996 , n24997 );
xor ( n25000 , n24907 , n24910 );
and ( n25001 , n18122 , n18456 );
and ( n25002 , n25000 , n25001 );
and ( n25003 , n24999 , n25002 );
or ( n25004 , n24998 , n25003 );
and ( n25005 , n24995 , n25004 );
or ( n25006 , n24994 , n25005 );
and ( n25007 , n24991 , n25006 );
or ( n25008 , n24990 , n25007 );
and ( n25009 , n24987 , n25008 );
or ( n25010 , n24986 , n25009 );
and ( n25011 , n24983 , n25010 );
or ( n25012 , n24982 , n25011 );
and ( n25013 , n24979 , n25012 );
or ( n25014 , n24978 , n25013 );
and ( n25015 , n24975 , n25014 );
or ( n25016 , n24974 , n25015 );
and ( n25017 , n24971 , n25016 );
or ( n25018 , n24970 , n25017 );
and ( n25019 , n24967 , n25018 );
or ( n25020 , n24966 , n25019 );
and ( n25021 , n24963 , n25020 );
or ( n25022 , n24962 , n25021 );
and ( n25023 , n24959 , n25022 );
or ( n25024 , n24958 , n25023 );
and ( n25025 , n24955 , n25024 );
or ( n25026 , n24954 , n25025 );
and ( n25027 , n24951 , n25026 );
or ( n25028 , n24950 , n25027 );
and ( n25029 , n24947 , n25028 );
or ( n25030 , n24946 , n25029 );
and ( n25031 , n24943 , n25030 );
or ( n25032 , n24942 , n25031 );
and ( n25033 , n18107 , n18454 );
and ( n25034 , n25032 , n25033 );
xor ( n25035 , n25032 , n25033 );
xor ( n25036 , n24943 , n25030 );
and ( n25037 , n18108 , n18454 );
and ( n25038 , n25036 , n25037 );
xor ( n25039 , n25036 , n25037 );
xor ( n25040 , n24947 , n25028 );
and ( n25041 , n18109 , n18454 );
and ( n25042 , n25040 , n25041 );
xor ( n25043 , n25040 , n25041 );
xor ( n25044 , n24951 , n25026 );
and ( n25045 , n18110 , n18454 );
and ( n25046 , n25044 , n25045 );
xor ( n25047 , n25044 , n25045 );
xor ( n25048 , n24955 , n25024 );
and ( n25049 , n18111 , n18454 );
and ( n25050 , n25048 , n25049 );
xor ( n25051 , n25048 , n25049 );
xor ( n25052 , n24959 , n25022 );
and ( n25053 , n18112 , n18454 );
and ( n25054 , n25052 , n25053 );
xor ( n25055 , n25052 , n25053 );
xor ( n25056 , n24963 , n25020 );
and ( n25057 , n18113 , n18454 );
and ( n25058 , n25056 , n25057 );
xor ( n25059 , n25056 , n25057 );
xor ( n25060 , n24967 , n25018 );
and ( n25061 , n18114 , n18454 );
and ( n25062 , n25060 , n25061 );
xor ( n25063 , n25060 , n25061 );
xor ( n25064 , n24971 , n25016 );
and ( n25065 , n18115 , n18454 );
and ( n25066 , n25064 , n25065 );
xor ( n25067 , n25064 , n25065 );
xor ( n25068 , n24975 , n25014 );
and ( n25069 , n18116 , n18454 );
and ( n25070 , n25068 , n25069 );
xor ( n25071 , n25068 , n25069 );
xor ( n25072 , n24979 , n25012 );
and ( n25073 , n18117 , n18454 );
and ( n25074 , n25072 , n25073 );
xor ( n25075 , n25072 , n25073 );
xor ( n25076 , n24983 , n25010 );
and ( n25077 , n18118 , n18454 );
and ( n25078 , n25076 , n25077 );
xor ( n25079 , n25076 , n25077 );
xor ( n25080 , n24987 , n25008 );
and ( n25081 , n18119 , n18454 );
and ( n25082 , n25080 , n25081 );
xor ( n25083 , n25080 , n25081 );
xor ( n25084 , n24991 , n25006 );
and ( n25085 , n18120 , n18454 );
and ( n25086 , n25084 , n25085 );
xor ( n25087 , n25084 , n25085 );
xor ( n25088 , n24995 , n25004 );
and ( n25089 , n18121 , n18454 );
and ( n25090 , n25088 , n25089 );
xor ( n25091 , n25088 , n25089 );
xor ( n25092 , n24999 , n25002 );
and ( n25093 , n18122 , n18454 );
and ( n25094 , n25092 , n25093 );
and ( n25095 , n25091 , n25094 );
or ( n25096 , n25090 , n25095 );
and ( n25097 , n25087 , n25096 );
or ( n25098 , n25086 , n25097 );
and ( n25099 , n25083 , n25098 );
or ( n25100 , n25082 , n25099 );
and ( n25101 , n25079 , n25100 );
or ( n25102 , n25078 , n25101 );
and ( n25103 , n25075 , n25102 );
or ( n25104 , n25074 , n25103 );
and ( n25105 , n25071 , n25104 );
or ( n25106 , n25070 , n25105 );
and ( n25107 , n25067 , n25106 );
or ( n25108 , n25066 , n25107 );
and ( n25109 , n25063 , n25108 );
or ( n25110 , n25062 , n25109 );
and ( n25111 , n25059 , n25110 );
or ( n25112 , n25058 , n25111 );
and ( n25113 , n25055 , n25112 );
or ( n25114 , n25054 , n25113 );
and ( n25115 , n25051 , n25114 );
or ( n25116 , n25050 , n25115 );
and ( n25117 , n25047 , n25116 );
or ( n25118 , n25046 , n25117 );
and ( n25119 , n25043 , n25118 );
or ( n25120 , n25042 , n25119 );
and ( n25121 , n25039 , n25120 );
or ( n25122 , n25038 , n25121 );
and ( n25123 , n25035 , n25122 );
or ( n25124 , n25034 , n25123 );
and ( n25125 , n18107 , n18452 );
and ( n25126 , n25124 , n25125 );
xor ( n25127 , n25124 , n25125 );
xor ( n25128 , n25035 , n25122 );
and ( n25129 , n18108 , n18452 );
and ( n25130 , n25128 , n25129 );
xor ( n25131 , n25128 , n25129 );
xor ( n25132 , n25039 , n25120 );
and ( n25133 , n18109 , n18452 );
and ( n25134 , n25132 , n25133 );
xor ( n25135 , n25132 , n25133 );
xor ( n25136 , n25043 , n25118 );
and ( n25137 , n18110 , n18452 );
and ( n25138 , n25136 , n25137 );
xor ( n25139 , n25136 , n25137 );
xor ( n25140 , n25047 , n25116 );
and ( n25141 , n18111 , n18452 );
and ( n25142 , n25140 , n25141 );
xor ( n25143 , n25140 , n25141 );
xor ( n25144 , n25051 , n25114 );
and ( n25145 , n18112 , n18452 );
and ( n25146 , n25144 , n25145 );
xor ( n25147 , n25144 , n25145 );
xor ( n25148 , n25055 , n25112 );
and ( n25149 , n18113 , n18452 );
and ( n25150 , n25148 , n25149 );
xor ( n25151 , n25148 , n25149 );
xor ( n25152 , n25059 , n25110 );
and ( n25153 , n18114 , n18452 );
and ( n25154 , n25152 , n25153 );
xor ( n25155 , n25152 , n25153 );
xor ( n25156 , n25063 , n25108 );
and ( n25157 , n18115 , n18452 );
and ( n25158 , n25156 , n25157 );
xor ( n25159 , n25156 , n25157 );
xor ( n25160 , n25067 , n25106 );
and ( n25161 , n18116 , n18452 );
and ( n25162 , n25160 , n25161 );
xor ( n25163 , n25160 , n25161 );
xor ( n25164 , n25071 , n25104 );
and ( n25165 , n18117 , n18452 );
and ( n25166 , n25164 , n25165 );
xor ( n25167 , n25164 , n25165 );
xor ( n25168 , n25075 , n25102 );
and ( n25169 , n18118 , n18452 );
and ( n25170 , n25168 , n25169 );
xor ( n25171 , n25168 , n25169 );
xor ( n25172 , n25079 , n25100 );
and ( n25173 , n18119 , n18452 );
and ( n25174 , n25172 , n25173 );
xor ( n25175 , n25172 , n25173 );
xor ( n25176 , n25083 , n25098 );
and ( n25177 , n18120 , n18452 );
and ( n25178 , n25176 , n25177 );
xor ( n25179 , n25176 , n25177 );
xor ( n25180 , n25087 , n25096 );
and ( n25181 , n18121 , n18452 );
and ( n25182 , n25180 , n25181 );
xor ( n25183 , n25180 , n25181 );
xor ( n25184 , n25091 , n25094 );
and ( n25185 , n18122 , n18452 );
and ( n25186 , n25184 , n25185 );
and ( n25187 , n25183 , n25186 );
or ( n25188 , n25182 , n25187 );
and ( n25189 , n25179 , n25188 );
or ( n25190 , n25178 , n25189 );
and ( n25191 , n25175 , n25190 );
or ( n25192 , n25174 , n25191 );
and ( n25193 , n25171 , n25192 );
or ( n25194 , n25170 , n25193 );
and ( n25195 , n25167 , n25194 );
or ( n25196 , n25166 , n25195 );
and ( n25197 , n25163 , n25196 );
or ( n25198 , n25162 , n25197 );
and ( n25199 , n25159 , n25198 );
or ( n25200 , n25158 , n25199 );
and ( n25201 , n25155 , n25200 );
or ( n25202 , n25154 , n25201 );
and ( n25203 , n25151 , n25202 );
or ( n25204 , n25150 , n25203 );
and ( n25205 , n25147 , n25204 );
or ( n25206 , n25146 , n25205 );
and ( n25207 , n25143 , n25206 );
or ( n25208 , n25142 , n25207 );
and ( n25209 , n25139 , n25208 );
or ( n25210 , n25138 , n25209 );
and ( n25211 , n25135 , n25210 );
or ( n25212 , n25134 , n25211 );
and ( n25213 , n25131 , n25212 );
or ( n25214 , n25130 , n25213 );
and ( n25215 , n25127 , n25214 );
or ( n25216 , n25126 , n25215 );
and ( n25217 , n18107 , n18450 );
and ( n25218 , n25216 , n25217 );
xor ( n25219 , n25216 , n25217 );
xor ( n25220 , n25127 , n25214 );
and ( n25221 , n18108 , n18450 );
and ( n25222 , n25220 , n25221 );
xor ( n25223 , n25220 , n25221 );
xor ( n25224 , n25131 , n25212 );
and ( n25225 , n18109 , n18450 );
and ( n25226 , n25224 , n25225 );
xor ( n25227 , n25224 , n25225 );
xor ( n25228 , n25135 , n25210 );
and ( n25229 , n18110 , n18450 );
and ( n25230 , n25228 , n25229 );
xor ( n25231 , n25228 , n25229 );
xor ( n25232 , n25139 , n25208 );
and ( n25233 , n18111 , n18450 );
and ( n25234 , n25232 , n25233 );
xor ( n25235 , n25232 , n25233 );
xor ( n25236 , n25143 , n25206 );
and ( n25237 , n18112 , n18450 );
and ( n25238 , n25236 , n25237 );
xor ( n25239 , n25236 , n25237 );
xor ( n25240 , n25147 , n25204 );
and ( n25241 , n18113 , n18450 );
and ( n25242 , n25240 , n25241 );
xor ( n25243 , n25240 , n25241 );
xor ( n25244 , n25151 , n25202 );
and ( n25245 , n18114 , n18450 );
and ( n25246 , n25244 , n25245 );
xor ( n25247 , n25244 , n25245 );
xor ( n25248 , n25155 , n25200 );
and ( n25249 , n18115 , n18450 );
and ( n25250 , n25248 , n25249 );
xor ( n25251 , n25248 , n25249 );
xor ( n25252 , n25159 , n25198 );
and ( n25253 , n18116 , n18450 );
and ( n25254 , n25252 , n25253 );
xor ( n25255 , n25252 , n25253 );
xor ( n25256 , n25163 , n25196 );
and ( n25257 , n18117 , n18450 );
and ( n25258 , n25256 , n25257 );
xor ( n25259 , n25256 , n25257 );
xor ( n25260 , n25167 , n25194 );
and ( n25261 , n18118 , n18450 );
and ( n25262 , n25260 , n25261 );
xor ( n25263 , n25260 , n25261 );
xor ( n25264 , n25171 , n25192 );
and ( n25265 , n18119 , n18450 );
and ( n25266 , n25264 , n25265 );
xor ( n25267 , n25264 , n25265 );
xor ( n25268 , n25175 , n25190 );
and ( n25269 , n18120 , n18450 );
and ( n25270 , n25268 , n25269 );
xor ( n25271 , n25268 , n25269 );
xor ( n25272 , n25179 , n25188 );
and ( n25273 , n18121 , n18450 );
and ( n25274 , n25272 , n25273 );
xor ( n25275 , n25272 , n25273 );
xor ( n25276 , n25183 , n25186 );
and ( n25277 , n18122 , n18450 );
and ( n25278 , n25276 , n25277 );
and ( n25279 , n25275 , n25278 );
or ( n25280 , n25274 , n25279 );
and ( n25281 , n25271 , n25280 );
or ( n25282 , n25270 , n25281 );
and ( n25283 , n25267 , n25282 );
or ( n25284 , n25266 , n25283 );
and ( n25285 , n25263 , n25284 );
or ( n25286 , n25262 , n25285 );
and ( n25287 , n25259 , n25286 );
or ( n25288 , n25258 , n25287 );
and ( n25289 , n25255 , n25288 );
or ( n25290 , n25254 , n25289 );
and ( n25291 , n25251 , n25290 );
or ( n25292 , n25250 , n25291 );
and ( n25293 , n25247 , n25292 );
or ( n25294 , n25246 , n25293 );
and ( n25295 , n25243 , n25294 );
or ( n25296 , n25242 , n25295 );
and ( n25297 , n25239 , n25296 );
or ( n25298 , n25238 , n25297 );
and ( n25299 , n25235 , n25298 );
or ( n25300 , n25234 , n25299 );
and ( n25301 , n25231 , n25300 );
or ( n25302 , n25230 , n25301 );
and ( n25303 , n25227 , n25302 );
or ( n25304 , n25226 , n25303 );
and ( n25305 , n25223 , n25304 );
or ( n25306 , n25222 , n25305 );
and ( n25307 , n25219 , n25306 );
or ( n25308 , n25218 , n25307 );
and ( n25309 , n18107 , n18448 );
and ( n25310 , n25308 , n25309 );
xor ( n25311 , n25308 , n25309 );
xor ( n25312 , n25219 , n25306 );
and ( n25313 , n18108 , n18448 );
and ( n25314 , n25312 , n25313 );
xor ( n25315 , n25312 , n25313 );
xor ( n25316 , n25223 , n25304 );
and ( n25317 , n18109 , n18448 );
and ( n25318 , n25316 , n25317 );
xor ( n25319 , n25316 , n25317 );
xor ( n25320 , n25227 , n25302 );
and ( n25321 , n18110 , n18448 );
and ( n25322 , n25320 , n25321 );
xor ( n25323 , n25320 , n25321 );
xor ( n25324 , n25231 , n25300 );
and ( n25325 , n18111 , n18448 );
and ( n25326 , n25324 , n25325 );
xor ( n25327 , n25324 , n25325 );
xor ( n25328 , n25235 , n25298 );
and ( n25329 , n18112 , n18448 );
and ( n25330 , n25328 , n25329 );
xor ( n25331 , n25328 , n25329 );
xor ( n25332 , n25239 , n25296 );
and ( n25333 , n18113 , n18448 );
and ( n25334 , n25332 , n25333 );
xor ( n25335 , n25332 , n25333 );
xor ( n25336 , n25243 , n25294 );
and ( n25337 , n18114 , n18448 );
and ( n25338 , n25336 , n25337 );
xor ( n25339 , n25336 , n25337 );
xor ( n25340 , n25247 , n25292 );
and ( n25341 , n18115 , n18448 );
and ( n25342 , n25340 , n25341 );
xor ( n25343 , n25340 , n25341 );
xor ( n25344 , n25251 , n25290 );
and ( n25345 , n18116 , n18448 );
and ( n25346 , n25344 , n25345 );
xor ( n25347 , n25344 , n25345 );
xor ( n25348 , n25255 , n25288 );
and ( n25349 , n18117 , n18448 );
and ( n25350 , n25348 , n25349 );
xor ( n25351 , n25348 , n25349 );
xor ( n25352 , n25259 , n25286 );
and ( n25353 , n18118 , n18448 );
and ( n25354 , n25352 , n25353 );
xor ( n25355 , n25352 , n25353 );
xor ( n25356 , n25263 , n25284 );
and ( n25357 , n18119 , n18448 );
and ( n25358 , n25356 , n25357 );
xor ( n25359 , n25356 , n25357 );
xor ( n25360 , n25267 , n25282 );
and ( n25361 , n18120 , n18448 );
and ( n25362 , n25360 , n25361 );
xor ( n25363 , n25360 , n25361 );
xor ( n25364 , n25271 , n25280 );
and ( n25365 , n18121 , n18448 );
and ( n25366 , n25364 , n25365 );
xor ( n25367 , n25364 , n25365 );
xor ( n25368 , n25275 , n25278 );
and ( n25369 , n18122 , n18448 );
and ( n25370 , n25368 , n25369 );
and ( n25371 , n25367 , n25370 );
or ( n25372 , n25366 , n25371 );
and ( n25373 , n25363 , n25372 );
or ( n25374 , n25362 , n25373 );
and ( n25375 , n25359 , n25374 );
or ( n25376 , n25358 , n25375 );
and ( n25377 , n25355 , n25376 );
or ( n25378 , n25354 , n25377 );
and ( n25379 , n25351 , n25378 );
or ( n25380 , n25350 , n25379 );
and ( n25381 , n25347 , n25380 );
or ( n25382 , n25346 , n25381 );
and ( n25383 , n25343 , n25382 );
or ( n25384 , n25342 , n25383 );
and ( n25385 , n25339 , n25384 );
or ( n25386 , n25338 , n25385 );
and ( n25387 , n25335 , n25386 );
or ( n25388 , n25334 , n25387 );
and ( n25389 , n25331 , n25388 );
or ( n25390 , n25330 , n25389 );
and ( n25391 , n25327 , n25390 );
or ( n25392 , n25326 , n25391 );
and ( n25393 , n25323 , n25392 );
or ( n25394 , n25322 , n25393 );
and ( n25395 , n25319 , n25394 );
or ( n25396 , n25318 , n25395 );
and ( n25397 , n25315 , n25396 );
or ( n25398 , n25314 , n25397 );
and ( n25399 , n25311 , n25398 );
or ( n25400 , n25310 , n25399 );
and ( n25401 , n18107 , n18446 );
and ( n25402 , n25400 , n25401 );
xor ( n25403 , n25400 , n25401 );
xor ( n25404 , n25311 , n25398 );
and ( n25405 , n18108 , n18446 );
and ( n25406 , n25404 , n25405 );
xor ( n25407 , n25404 , n25405 );
xor ( n25408 , n25315 , n25396 );
and ( n25409 , n18109 , n18446 );
and ( n25410 , n25408 , n25409 );
xor ( n25411 , n25408 , n25409 );
xor ( n25412 , n25319 , n25394 );
and ( n25413 , n18110 , n18446 );
and ( n25414 , n25412 , n25413 );
xor ( n25415 , n25412 , n25413 );
xor ( n25416 , n25323 , n25392 );
and ( n25417 , n18111 , n18446 );
and ( n25418 , n25416 , n25417 );
xor ( n25419 , n25416 , n25417 );
xor ( n25420 , n25327 , n25390 );
and ( n25421 , n18112 , n18446 );
and ( n25422 , n25420 , n25421 );
xor ( n25423 , n25420 , n25421 );
xor ( n25424 , n25331 , n25388 );
and ( n25425 , n18113 , n18446 );
and ( n25426 , n25424 , n25425 );
xor ( n25427 , n25424 , n25425 );
xor ( n25428 , n25335 , n25386 );
and ( n25429 , n18114 , n18446 );
and ( n25430 , n25428 , n25429 );
xor ( n25431 , n25428 , n25429 );
xor ( n25432 , n25339 , n25384 );
and ( n25433 , n18115 , n18446 );
and ( n25434 , n25432 , n25433 );
xor ( n25435 , n25432 , n25433 );
xor ( n25436 , n25343 , n25382 );
and ( n25437 , n18116 , n18446 );
and ( n25438 , n25436 , n25437 );
xor ( n25439 , n25436 , n25437 );
xor ( n25440 , n25347 , n25380 );
and ( n25441 , n18117 , n18446 );
and ( n25442 , n25440 , n25441 );
xor ( n25443 , n25440 , n25441 );
xor ( n25444 , n25351 , n25378 );
and ( n25445 , n18118 , n18446 );
and ( n25446 , n25444 , n25445 );
xor ( n25447 , n25444 , n25445 );
xor ( n25448 , n25355 , n25376 );
and ( n25449 , n18119 , n18446 );
and ( n25450 , n25448 , n25449 );
xor ( n25451 , n25448 , n25449 );
xor ( n25452 , n25359 , n25374 );
and ( n25453 , n18120 , n18446 );
and ( n25454 , n25452 , n25453 );
xor ( n25455 , n25452 , n25453 );
xor ( n25456 , n25363 , n25372 );
and ( n25457 , n18121 , n18446 );
and ( n25458 , n25456 , n25457 );
xor ( n25459 , n25456 , n25457 );
xor ( n25460 , n25367 , n25370 );
and ( n25461 , n18122 , n18446 );
and ( n25462 , n25460 , n25461 );
and ( n25463 , n25459 , n25462 );
or ( n25464 , n25458 , n25463 );
and ( n25465 , n25455 , n25464 );
or ( n25466 , n25454 , n25465 );
and ( n25467 , n25451 , n25466 );
or ( n25468 , n25450 , n25467 );
and ( n25469 , n25447 , n25468 );
or ( n25470 , n25446 , n25469 );
and ( n25471 , n25443 , n25470 );
or ( n25472 , n25442 , n25471 );
and ( n25473 , n25439 , n25472 );
or ( n25474 , n25438 , n25473 );
and ( n25475 , n25435 , n25474 );
or ( n25476 , n25434 , n25475 );
and ( n25477 , n25431 , n25476 );
or ( n25478 , n25430 , n25477 );
and ( n25479 , n25427 , n25478 );
or ( n25480 , n25426 , n25479 );
and ( n25481 , n25423 , n25480 );
or ( n25482 , n25422 , n25481 );
and ( n25483 , n25419 , n25482 );
or ( n25484 , n25418 , n25483 );
and ( n25485 , n25415 , n25484 );
or ( n25486 , n25414 , n25485 );
and ( n25487 , n25411 , n25486 );
or ( n25488 , n25410 , n25487 );
and ( n25489 , n25407 , n25488 );
or ( n25490 , n25406 , n25489 );
and ( n25491 , n25403 , n25490 );
or ( n25492 , n25402 , n25491 );
and ( n25493 , n18107 , n18444 );
and ( n25494 , n25492 , n25493 );
xor ( n25495 , n25492 , n25493 );
xor ( n25496 , n25403 , n25490 );
and ( n25497 , n18108 , n18444 );
and ( n25498 , n25496 , n25497 );
xor ( n25499 , n25496 , n25497 );
xor ( n25500 , n25407 , n25488 );
and ( n25501 , n18109 , n18444 );
and ( n25502 , n25500 , n25501 );
xor ( n25503 , n25500 , n25501 );
xor ( n25504 , n25411 , n25486 );
and ( n25505 , n18110 , n18444 );
and ( n25506 , n25504 , n25505 );
xor ( n25507 , n25504 , n25505 );
xor ( n25508 , n25415 , n25484 );
and ( n25509 , n18111 , n18444 );
and ( n25510 , n25508 , n25509 );
xor ( n25511 , n25508 , n25509 );
xor ( n25512 , n25419 , n25482 );
and ( n25513 , n18112 , n18444 );
and ( n25514 , n25512 , n25513 );
xor ( n25515 , n25512 , n25513 );
xor ( n25516 , n25423 , n25480 );
and ( n25517 , n18113 , n18444 );
and ( n25518 , n25516 , n25517 );
xor ( n25519 , n25516 , n25517 );
xor ( n25520 , n25427 , n25478 );
and ( n25521 , n18114 , n18444 );
and ( n25522 , n25520 , n25521 );
xor ( n25523 , n25520 , n25521 );
xor ( n25524 , n25431 , n25476 );
and ( n25525 , n18115 , n18444 );
and ( n25526 , n25524 , n25525 );
xor ( n25527 , n25524 , n25525 );
xor ( n25528 , n25435 , n25474 );
and ( n25529 , n18116 , n18444 );
and ( n25530 , n25528 , n25529 );
xor ( n25531 , n25528 , n25529 );
xor ( n25532 , n25439 , n25472 );
and ( n25533 , n18117 , n18444 );
and ( n25534 , n25532 , n25533 );
xor ( n25535 , n25532 , n25533 );
xor ( n25536 , n25443 , n25470 );
and ( n25537 , n18118 , n18444 );
and ( n25538 , n25536 , n25537 );
xor ( n25539 , n25536 , n25537 );
xor ( n25540 , n25447 , n25468 );
and ( n25541 , n18119 , n18444 );
and ( n25542 , n25540 , n25541 );
xor ( n25543 , n25540 , n25541 );
xor ( n25544 , n25451 , n25466 );
and ( n25545 , n18120 , n18444 );
and ( n25546 , n25544 , n25545 );
xor ( n25547 , n25544 , n25545 );
xor ( n25548 , n25455 , n25464 );
and ( n25549 , n18121 , n18444 );
and ( n25550 , n25548 , n25549 );
xor ( n25551 , n25548 , n25549 );
xor ( n25552 , n25459 , n25462 );
and ( n25553 , n18122 , n18444 );
and ( n25554 , n25552 , n25553 );
and ( n25555 , n25551 , n25554 );
or ( n25556 , n25550 , n25555 );
and ( n25557 , n25547 , n25556 );
or ( n25558 , n25546 , n25557 );
and ( n25559 , n25543 , n25558 );
or ( n25560 , n25542 , n25559 );
and ( n25561 , n25539 , n25560 );
or ( n25562 , n25538 , n25561 );
and ( n25563 , n25535 , n25562 );
or ( n25564 , n25534 , n25563 );
and ( n25565 , n25531 , n25564 );
or ( n25566 , n25530 , n25565 );
and ( n25567 , n25527 , n25566 );
or ( n25568 , n25526 , n25567 );
and ( n25569 , n25523 , n25568 );
or ( n25570 , n25522 , n25569 );
and ( n25571 , n25519 , n25570 );
or ( n25572 , n25518 , n25571 );
and ( n25573 , n25515 , n25572 );
or ( n25574 , n25514 , n25573 );
and ( n25575 , n25511 , n25574 );
or ( n25576 , n25510 , n25575 );
and ( n25577 , n25507 , n25576 );
or ( n25578 , n25506 , n25577 );
and ( n25579 , n25503 , n25578 );
or ( n25580 , n25502 , n25579 );
and ( n25581 , n25499 , n25580 );
or ( n25582 , n25498 , n25581 );
and ( n25583 , n25495 , n25582 );
or ( n25584 , n25494 , n25583 );
and ( n25585 , n18107 , n18442 );
and ( n25586 , n25584 , n25585 );
xor ( n25587 , n25584 , n25585 );
xor ( n25588 , n25495 , n25582 );
and ( n25589 , n18108 , n18442 );
and ( n25590 , n25588 , n25589 );
xor ( n25591 , n25588 , n25589 );
xor ( n25592 , n25499 , n25580 );
and ( n25593 , n18109 , n18442 );
and ( n25594 , n25592 , n25593 );
xor ( n25595 , n25592 , n25593 );
xor ( n25596 , n25503 , n25578 );
and ( n25597 , n18110 , n18442 );
and ( n25598 , n25596 , n25597 );
xor ( n25599 , n25596 , n25597 );
xor ( n25600 , n25507 , n25576 );
and ( n25601 , n18111 , n18442 );
and ( n25602 , n25600 , n25601 );
xor ( n25603 , n25600 , n25601 );
xor ( n25604 , n25511 , n25574 );
and ( n25605 , n18112 , n18442 );
and ( n25606 , n25604 , n25605 );
xor ( n25607 , n25604 , n25605 );
xor ( n25608 , n25515 , n25572 );
and ( n25609 , n18113 , n18442 );
and ( n25610 , n25608 , n25609 );
xor ( n25611 , n25608 , n25609 );
xor ( n25612 , n25519 , n25570 );
and ( n25613 , n18114 , n18442 );
and ( n25614 , n25612 , n25613 );
xor ( n25615 , n25612 , n25613 );
xor ( n25616 , n25523 , n25568 );
and ( n25617 , n18115 , n18442 );
and ( n25618 , n25616 , n25617 );
xor ( n25619 , n25616 , n25617 );
xor ( n25620 , n25527 , n25566 );
and ( n25621 , n18116 , n18442 );
and ( n25622 , n25620 , n25621 );
xor ( n25623 , n25620 , n25621 );
xor ( n25624 , n25531 , n25564 );
and ( n25625 , n18117 , n18442 );
and ( n25626 , n25624 , n25625 );
xor ( n25627 , n25624 , n25625 );
xor ( n25628 , n25535 , n25562 );
and ( n25629 , n18118 , n18442 );
and ( n25630 , n25628 , n25629 );
xor ( n25631 , n25628 , n25629 );
xor ( n25632 , n25539 , n25560 );
and ( n25633 , n18119 , n18442 );
and ( n25634 , n25632 , n25633 );
xor ( n25635 , n25632 , n25633 );
xor ( n25636 , n25543 , n25558 );
and ( n25637 , n18120 , n18442 );
and ( n25638 , n25636 , n25637 );
xor ( n25639 , n25636 , n25637 );
xor ( n25640 , n25547 , n25556 );
and ( n25641 , n18121 , n18442 );
and ( n25642 , n25640 , n25641 );
xor ( n25643 , n25640 , n25641 );
xor ( n25644 , n25551 , n25554 );
and ( n25645 , n18122 , n18442 );
and ( n25646 , n25644 , n25645 );
and ( n25647 , n25643 , n25646 );
or ( n25648 , n25642 , n25647 );
and ( n25649 , n25639 , n25648 );
or ( n25650 , n25638 , n25649 );
and ( n25651 , n25635 , n25650 );
or ( n25652 , n25634 , n25651 );
and ( n25653 , n25631 , n25652 );
or ( n25654 , n25630 , n25653 );
and ( n25655 , n25627 , n25654 );
or ( n25656 , n25626 , n25655 );
and ( n25657 , n25623 , n25656 );
or ( n25658 , n25622 , n25657 );
and ( n25659 , n25619 , n25658 );
or ( n25660 , n25618 , n25659 );
and ( n25661 , n25615 , n25660 );
or ( n25662 , n25614 , n25661 );
and ( n25663 , n25611 , n25662 );
or ( n25664 , n25610 , n25663 );
and ( n25665 , n25607 , n25664 );
or ( n25666 , n25606 , n25665 );
and ( n25667 , n25603 , n25666 );
or ( n25668 , n25602 , n25667 );
and ( n25669 , n25599 , n25668 );
or ( n25670 , n25598 , n25669 );
and ( n25671 , n25595 , n25670 );
or ( n25672 , n25594 , n25671 );
and ( n25673 , n25591 , n25672 );
or ( n25674 , n25590 , n25673 );
and ( n25675 , n25587 , n25674 );
or ( n25676 , n25586 , n25675 );
and ( n25677 , n18107 , n18440 );
and ( n25678 , n25676 , n25677 );
xor ( n25679 , n25676 , n25677 );
xor ( n25680 , n25587 , n25674 );
and ( n25681 , n18108 , n18440 );
and ( n25682 , n25680 , n25681 );
xor ( n25683 , n25680 , n25681 );
xor ( n25684 , n25591 , n25672 );
and ( n25685 , n18109 , n18440 );
and ( n25686 , n25684 , n25685 );
xor ( n25687 , n25684 , n25685 );
xor ( n25688 , n25595 , n25670 );
and ( n25689 , n18110 , n18440 );
and ( n25690 , n25688 , n25689 );
xor ( n25691 , n25688 , n25689 );
xor ( n25692 , n25599 , n25668 );
and ( n25693 , n18111 , n18440 );
and ( n25694 , n25692 , n25693 );
xor ( n25695 , n25692 , n25693 );
xor ( n25696 , n25603 , n25666 );
and ( n25697 , n18112 , n18440 );
and ( n25698 , n25696 , n25697 );
xor ( n25699 , n25696 , n25697 );
xor ( n25700 , n25607 , n25664 );
and ( n25701 , n18113 , n18440 );
and ( n25702 , n25700 , n25701 );
xor ( n25703 , n25700 , n25701 );
xor ( n25704 , n25611 , n25662 );
and ( n25705 , n18114 , n18440 );
and ( n25706 , n25704 , n25705 );
xor ( n25707 , n25704 , n25705 );
xor ( n25708 , n25615 , n25660 );
and ( n25709 , n18115 , n18440 );
and ( n25710 , n25708 , n25709 );
xor ( n25711 , n25708 , n25709 );
xor ( n25712 , n25619 , n25658 );
and ( n25713 , n18116 , n18440 );
and ( n25714 , n25712 , n25713 );
xor ( n25715 , n25712 , n25713 );
xor ( n25716 , n25623 , n25656 );
and ( n25717 , n18117 , n18440 );
and ( n25718 , n25716 , n25717 );
xor ( n25719 , n25716 , n25717 );
xor ( n25720 , n25627 , n25654 );
and ( n25721 , n18118 , n18440 );
and ( n25722 , n25720 , n25721 );
xor ( n25723 , n25720 , n25721 );
xor ( n25724 , n25631 , n25652 );
and ( n25725 , n18119 , n18440 );
and ( n25726 , n25724 , n25725 );
xor ( n25727 , n25724 , n25725 );
xor ( n25728 , n25635 , n25650 );
and ( n25729 , n18120 , n18440 );
and ( n25730 , n25728 , n25729 );
xor ( n25731 , n25728 , n25729 );
xor ( n25732 , n25639 , n25648 );
and ( n25733 , n18121 , n18440 );
and ( n25734 , n25732 , n25733 );
xor ( n25735 , n25732 , n25733 );
xor ( n25736 , n25643 , n25646 );
and ( n25737 , n18122 , n18440 );
and ( n25738 , n25736 , n25737 );
and ( n25739 , n25735 , n25738 );
or ( n25740 , n25734 , n25739 );
and ( n25741 , n25731 , n25740 );
or ( n25742 , n25730 , n25741 );
and ( n25743 , n25727 , n25742 );
or ( n25744 , n25726 , n25743 );
and ( n25745 , n25723 , n25744 );
or ( n25746 , n25722 , n25745 );
and ( n25747 , n25719 , n25746 );
or ( n25748 , n25718 , n25747 );
and ( n25749 , n25715 , n25748 );
or ( n25750 , n25714 , n25749 );
and ( n25751 , n25711 , n25750 );
or ( n25752 , n25710 , n25751 );
and ( n25753 , n25707 , n25752 );
or ( n25754 , n25706 , n25753 );
and ( n25755 , n25703 , n25754 );
or ( n25756 , n25702 , n25755 );
and ( n25757 , n25699 , n25756 );
or ( n25758 , n25698 , n25757 );
and ( n25759 , n25695 , n25758 );
or ( n25760 , n25694 , n25759 );
and ( n25761 , n25691 , n25760 );
or ( n25762 , n25690 , n25761 );
and ( n25763 , n25687 , n25762 );
or ( n25764 , n25686 , n25763 );
and ( n25765 , n25683 , n25764 );
or ( n25766 , n25682 , n25765 );
and ( n25767 , n25679 , n25766 );
or ( n25768 , n25678 , n25767 );
and ( n25769 , n18107 , n18438 );
and ( n25770 , n25768 , n25769 );
xor ( n25771 , n25768 , n25769 );
xor ( n25772 , n25679 , n25766 );
and ( n25773 , n18108 , n18438 );
and ( n25774 , n25772 , n25773 );
xor ( n25775 , n25772 , n25773 );
xor ( n25776 , n25683 , n25764 );
and ( n25777 , n18109 , n18438 );
and ( n25778 , n25776 , n25777 );
xor ( n25779 , n25776 , n25777 );
xor ( n25780 , n25687 , n25762 );
and ( n25781 , n18110 , n18438 );
and ( n25782 , n25780 , n25781 );
xor ( n25783 , n25780 , n25781 );
xor ( n25784 , n25691 , n25760 );
and ( n25785 , n18111 , n18438 );
and ( n25786 , n25784 , n25785 );
xor ( n25787 , n25784 , n25785 );
xor ( n25788 , n25695 , n25758 );
and ( n25789 , n18112 , n18438 );
and ( n25790 , n25788 , n25789 );
xor ( n25791 , n25788 , n25789 );
xor ( n25792 , n25699 , n25756 );
and ( n25793 , n18113 , n18438 );
and ( n25794 , n25792 , n25793 );
xor ( n25795 , n25792 , n25793 );
xor ( n25796 , n25703 , n25754 );
and ( n25797 , n18114 , n18438 );
and ( n25798 , n25796 , n25797 );
xor ( n25799 , n25796 , n25797 );
xor ( n25800 , n25707 , n25752 );
and ( n25801 , n18115 , n18438 );
and ( n25802 , n25800 , n25801 );
xor ( n25803 , n25800 , n25801 );
xor ( n25804 , n25711 , n25750 );
and ( n25805 , n18116 , n18438 );
and ( n25806 , n25804 , n25805 );
xor ( n25807 , n25804 , n25805 );
xor ( n25808 , n25715 , n25748 );
and ( n25809 , n18117 , n18438 );
and ( n25810 , n25808 , n25809 );
xor ( n25811 , n25808 , n25809 );
xor ( n25812 , n25719 , n25746 );
and ( n25813 , n18118 , n18438 );
and ( n25814 , n25812 , n25813 );
xor ( n25815 , n25812 , n25813 );
xor ( n25816 , n25723 , n25744 );
and ( n25817 , n18119 , n18438 );
and ( n25818 , n25816 , n25817 );
xor ( n25819 , n25816 , n25817 );
xor ( n25820 , n25727 , n25742 );
and ( n25821 , n18120 , n18438 );
and ( n25822 , n25820 , n25821 );
xor ( n25823 , n25820 , n25821 );
xor ( n25824 , n25731 , n25740 );
and ( n25825 , n18121 , n18438 );
and ( n25826 , n25824 , n25825 );
xor ( n25827 , n25824 , n25825 );
xor ( n25828 , n25735 , n25738 );
and ( n25829 , n18122 , n18438 );
and ( n25830 , n25828 , n25829 );
and ( n25831 , n25827 , n25830 );
or ( n25832 , n25826 , n25831 );
and ( n25833 , n25823 , n25832 );
or ( n25834 , n25822 , n25833 );
and ( n25835 , n25819 , n25834 );
or ( n25836 , n25818 , n25835 );
and ( n25837 , n25815 , n25836 );
or ( n25838 , n25814 , n25837 );
and ( n25839 , n25811 , n25838 );
or ( n25840 , n25810 , n25839 );
and ( n25841 , n25807 , n25840 );
or ( n25842 , n25806 , n25841 );
and ( n25843 , n25803 , n25842 );
or ( n25844 , n25802 , n25843 );
and ( n25845 , n25799 , n25844 );
or ( n25846 , n25798 , n25845 );
and ( n25847 , n25795 , n25846 );
or ( n25848 , n25794 , n25847 );
and ( n25849 , n25791 , n25848 );
or ( n25850 , n25790 , n25849 );
and ( n25851 , n25787 , n25850 );
or ( n25852 , n25786 , n25851 );
and ( n25853 , n25783 , n25852 );
or ( n25854 , n25782 , n25853 );
and ( n25855 , n25779 , n25854 );
or ( n25856 , n25778 , n25855 );
and ( n25857 , n25775 , n25856 );
or ( n25858 , n25774 , n25857 );
and ( n25859 , n25771 , n25858 );
or ( n25860 , n25770 , n25859 );
and ( n25861 , n18107 , n18436 );
and ( n25862 , n25860 , n25861 );
xor ( n25863 , n25860 , n25861 );
xor ( n25864 , n25771 , n25858 );
and ( n25865 , n18108 , n18436 );
and ( n25866 , n25864 , n25865 );
xor ( n25867 , n25864 , n25865 );
xor ( n25868 , n25775 , n25856 );
and ( n25869 , n18109 , n18436 );
and ( n25870 , n25868 , n25869 );
xor ( n25871 , n25868 , n25869 );
xor ( n25872 , n25779 , n25854 );
and ( n25873 , n18110 , n18436 );
and ( n25874 , n25872 , n25873 );
xor ( n25875 , n25872 , n25873 );
xor ( n25876 , n25783 , n25852 );
and ( n25877 , n18111 , n18436 );
and ( n25878 , n25876 , n25877 );
xor ( n25879 , n25876 , n25877 );
xor ( n25880 , n25787 , n25850 );
and ( n25881 , n18112 , n18436 );
and ( n25882 , n25880 , n25881 );
xor ( n25883 , n25880 , n25881 );
xor ( n25884 , n25791 , n25848 );
and ( n25885 , n18113 , n18436 );
and ( n25886 , n25884 , n25885 );
xor ( n25887 , n25884 , n25885 );
xor ( n25888 , n25795 , n25846 );
and ( n25889 , n18114 , n18436 );
and ( n25890 , n25888 , n25889 );
xor ( n25891 , n25888 , n25889 );
xor ( n25892 , n25799 , n25844 );
and ( n25893 , n18115 , n18436 );
and ( n25894 , n25892 , n25893 );
xor ( n25895 , n25892 , n25893 );
xor ( n25896 , n25803 , n25842 );
and ( n25897 , n18116 , n18436 );
and ( n25898 , n25896 , n25897 );
xor ( n25899 , n25896 , n25897 );
xor ( n25900 , n25807 , n25840 );
and ( n25901 , n18117 , n18436 );
and ( n25902 , n25900 , n25901 );
xor ( n25903 , n25900 , n25901 );
xor ( n25904 , n25811 , n25838 );
and ( n25905 , n18118 , n18436 );
and ( n25906 , n25904 , n25905 );
xor ( n25907 , n25904 , n25905 );
xor ( n25908 , n25815 , n25836 );
and ( n25909 , n18119 , n18436 );
and ( n25910 , n25908 , n25909 );
xor ( n25911 , n25908 , n25909 );
xor ( n25912 , n25819 , n25834 );
and ( n25913 , n18120 , n18436 );
and ( n25914 , n25912 , n25913 );
xor ( n25915 , n25912 , n25913 );
xor ( n25916 , n25823 , n25832 );
and ( n25917 , n18121 , n18436 );
and ( n25918 , n25916 , n25917 );
xor ( n25919 , n25916 , n25917 );
xor ( n25920 , n25827 , n25830 );
and ( n25921 , n18122 , n18436 );
and ( n25922 , n25920 , n25921 );
and ( n25923 , n25919 , n25922 );
or ( n25924 , n25918 , n25923 );
and ( n25925 , n25915 , n25924 );
or ( n25926 , n25914 , n25925 );
and ( n25927 , n25911 , n25926 );
or ( n25928 , n25910 , n25927 );
and ( n25929 , n25907 , n25928 );
or ( n25930 , n25906 , n25929 );
and ( n25931 , n25903 , n25930 );
or ( n25932 , n25902 , n25931 );
and ( n25933 , n25899 , n25932 );
or ( n25934 , n25898 , n25933 );
and ( n25935 , n25895 , n25934 );
or ( n25936 , n25894 , n25935 );
and ( n25937 , n25891 , n25936 );
or ( n25938 , n25890 , n25937 );
and ( n25939 , n25887 , n25938 );
or ( n25940 , n25886 , n25939 );
and ( n25941 , n25883 , n25940 );
or ( n25942 , n25882 , n25941 );
and ( n25943 , n25879 , n25942 );
or ( n25944 , n25878 , n25943 );
and ( n25945 , n25875 , n25944 );
or ( n25946 , n25874 , n25945 );
and ( n25947 , n25871 , n25946 );
or ( n25948 , n25870 , n25947 );
and ( n25949 , n25867 , n25948 );
or ( n25950 , n25866 , n25949 );
and ( n25951 , n25863 , n25950 );
or ( n25952 , n25862 , n25951 );
and ( n25953 , n18107 , n18434 );
and ( n25954 , n25952 , n25953 );
xor ( n25955 , n25952 , n25953 );
xor ( n25956 , n25863 , n25950 );
and ( n25957 , n18108 , n18434 );
and ( n25958 , n25956 , n25957 );
xor ( n25959 , n25956 , n25957 );
xor ( n25960 , n25867 , n25948 );
and ( n25961 , n18109 , n18434 );
and ( n25962 , n25960 , n25961 );
xor ( n25963 , n25960 , n25961 );
xor ( n25964 , n25871 , n25946 );
and ( n25965 , n18110 , n18434 );
and ( n25966 , n25964 , n25965 );
xor ( n25967 , n25964 , n25965 );
xor ( n25968 , n25875 , n25944 );
and ( n25969 , n18111 , n18434 );
and ( n25970 , n25968 , n25969 );
xor ( n25971 , n25968 , n25969 );
xor ( n25972 , n25879 , n25942 );
and ( n25973 , n18112 , n18434 );
and ( n25974 , n25972 , n25973 );
xor ( n25975 , n25972 , n25973 );
xor ( n25976 , n25883 , n25940 );
and ( n25977 , n18113 , n18434 );
and ( n25978 , n25976 , n25977 );
xor ( n25979 , n25976 , n25977 );
xor ( n25980 , n25887 , n25938 );
and ( n25981 , n18114 , n18434 );
and ( n25982 , n25980 , n25981 );
xor ( n25983 , n25980 , n25981 );
xor ( n25984 , n25891 , n25936 );
and ( n25985 , n18115 , n18434 );
and ( n25986 , n25984 , n25985 );
xor ( n25987 , n25984 , n25985 );
xor ( n25988 , n25895 , n25934 );
and ( n25989 , n18116 , n18434 );
and ( n25990 , n25988 , n25989 );
xor ( n25991 , n25988 , n25989 );
xor ( n25992 , n25899 , n25932 );
and ( n25993 , n18117 , n18434 );
and ( n25994 , n25992 , n25993 );
xor ( n25995 , n25992 , n25993 );
xor ( n25996 , n25903 , n25930 );
and ( n25997 , n18118 , n18434 );
and ( n25998 , n25996 , n25997 );
xor ( n25999 , n25996 , n25997 );
xor ( n26000 , n25907 , n25928 );
and ( n26001 , n18119 , n18434 );
and ( n26002 , n26000 , n26001 );
xor ( n26003 , n26000 , n26001 );
xor ( n26004 , n25911 , n25926 );
and ( n26005 , n18120 , n18434 );
and ( n26006 , n26004 , n26005 );
xor ( n26007 , n26004 , n26005 );
xor ( n26008 , n25915 , n25924 );
and ( n26009 , n18121 , n18434 );
and ( n26010 , n26008 , n26009 );
xor ( n26011 , n26008 , n26009 );
xor ( n26012 , n25919 , n25922 );
and ( n26013 , n18122 , n18434 );
and ( n26014 , n26012 , n26013 );
and ( n26015 , n26011 , n26014 );
or ( n26016 , n26010 , n26015 );
and ( n26017 , n26007 , n26016 );
or ( n26018 , n26006 , n26017 );
and ( n26019 , n26003 , n26018 );
or ( n26020 , n26002 , n26019 );
and ( n26021 , n25999 , n26020 );
or ( n26022 , n25998 , n26021 );
and ( n26023 , n25995 , n26022 );
or ( n26024 , n25994 , n26023 );
and ( n26025 , n25991 , n26024 );
or ( n26026 , n25990 , n26025 );
and ( n26027 , n25987 , n26026 );
or ( n26028 , n25986 , n26027 );
and ( n26029 , n25983 , n26028 );
or ( n26030 , n25982 , n26029 );
and ( n26031 , n25979 , n26030 );
or ( n26032 , n25978 , n26031 );
and ( n26033 , n25975 , n26032 );
or ( n26034 , n25974 , n26033 );
and ( n26035 , n25971 , n26034 );
or ( n26036 , n25970 , n26035 );
and ( n26037 , n25967 , n26036 );
or ( n26038 , n25966 , n26037 );
and ( n26039 , n25963 , n26038 );
or ( n26040 , n25962 , n26039 );
and ( n26041 , n25959 , n26040 );
or ( n26042 , n25958 , n26041 );
and ( n26043 , n25955 , n26042 );
or ( n26044 , n25954 , n26043 );
and ( n26045 , n18107 , n18432 );
and ( n26046 , n26044 , n26045 );
xor ( n26047 , n26044 , n26045 );
xor ( n26048 , n25955 , n26042 );
and ( n26049 , n18108 , n18432 );
and ( n26050 , n26048 , n26049 );
xor ( n26051 , n26048 , n26049 );
xor ( n26052 , n25959 , n26040 );
and ( n26053 , n18109 , n18432 );
and ( n26054 , n26052 , n26053 );
xor ( n26055 , n26052 , n26053 );
xor ( n26056 , n25963 , n26038 );
and ( n26057 , n18110 , n18432 );
and ( n26058 , n26056 , n26057 );
xor ( n26059 , n26056 , n26057 );
xor ( n26060 , n25967 , n26036 );
and ( n26061 , n18111 , n18432 );
and ( n26062 , n26060 , n26061 );
xor ( n26063 , n26060 , n26061 );
xor ( n26064 , n25971 , n26034 );
and ( n26065 , n18112 , n18432 );
and ( n26066 , n26064 , n26065 );
xor ( n26067 , n26064 , n26065 );
xor ( n26068 , n25975 , n26032 );
and ( n26069 , n18113 , n18432 );
and ( n26070 , n26068 , n26069 );
xor ( n26071 , n26068 , n26069 );
xor ( n26072 , n25979 , n26030 );
and ( n26073 , n18114 , n18432 );
and ( n26074 , n26072 , n26073 );
xor ( n26075 , n26072 , n26073 );
xor ( n26076 , n25983 , n26028 );
and ( n26077 , n18115 , n18432 );
and ( n26078 , n26076 , n26077 );
xor ( n26079 , n26076 , n26077 );
xor ( n26080 , n25987 , n26026 );
and ( n26081 , n18116 , n18432 );
and ( n26082 , n26080 , n26081 );
xor ( n26083 , n26080 , n26081 );
xor ( n26084 , n25991 , n26024 );
and ( n26085 , n18117 , n18432 );
and ( n26086 , n26084 , n26085 );
xor ( n26087 , n26084 , n26085 );
xor ( n26088 , n25995 , n26022 );
and ( n26089 , n18118 , n18432 );
and ( n26090 , n26088 , n26089 );
xor ( n26091 , n26088 , n26089 );
xor ( n26092 , n25999 , n26020 );
and ( n26093 , n18119 , n18432 );
and ( n26094 , n26092 , n26093 );
xor ( n26095 , n26092 , n26093 );
xor ( n26096 , n26003 , n26018 );
and ( n26097 , n18120 , n18432 );
and ( n26098 , n26096 , n26097 );
xor ( n26099 , n26096 , n26097 );
xor ( n26100 , n26007 , n26016 );
and ( n26101 , n18121 , n18432 );
and ( n26102 , n26100 , n26101 );
xor ( n26103 , n26100 , n26101 );
xor ( n26104 , n26011 , n26014 );
and ( n26105 , n18122 , n18432 );
and ( n26106 , n26104 , n26105 );
and ( n26107 , n26103 , n26106 );
or ( n26108 , n26102 , n26107 );
and ( n26109 , n26099 , n26108 );
or ( n26110 , n26098 , n26109 );
and ( n26111 , n26095 , n26110 );
or ( n26112 , n26094 , n26111 );
and ( n26113 , n26091 , n26112 );
or ( n26114 , n26090 , n26113 );
and ( n26115 , n26087 , n26114 );
or ( n26116 , n26086 , n26115 );
and ( n26117 , n26083 , n26116 );
or ( n26118 , n26082 , n26117 );
and ( n26119 , n26079 , n26118 );
or ( n26120 , n26078 , n26119 );
and ( n26121 , n26075 , n26120 );
or ( n26122 , n26074 , n26121 );
and ( n26123 , n26071 , n26122 );
or ( n26124 , n26070 , n26123 );
and ( n26125 , n26067 , n26124 );
or ( n26126 , n26066 , n26125 );
and ( n26127 , n26063 , n26126 );
or ( n26128 , n26062 , n26127 );
and ( n26129 , n26059 , n26128 );
or ( n26130 , n26058 , n26129 );
and ( n26131 , n26055 , n26130 );
or ( n26132 , n26054 , n26131 );
and ( n26133 , n26051 , n26132 );
or ( n26134 , n26050 , n26133 );
and ( n26135 , n26047 , n26134 );
or ( n26136 , n26046 , n26135 );
and ( n26137 , n18107 , n18430 );
and ( n26138 , n26136 , n26137 );
xor ( n26139 , n26136 , n26137 );
xor ( n26140 , n26047 , n26134 );
and ( n26141 , n18108 , n18430 );
and ( n26142 , n26140 , n26141 );
xor ( n26143 , n26140 , n26141 );
xor ( n26144 , n26051 , n26132 );
and ( n26145 , n18109 , n18430 );
and ( n26146 , n26144 , n26145 );
xor ( n26147 , n26144 , n26145 );
xor ( n26148 , n26055 , n26130 );
and ( n26149 , n18110 , n18430 );
and ( n26150 , n26148 , n26149 );
xor ( n26151 , n26148 , n26149 );
xor ( n26152 , n26059 , n26128 );
and ( n26153 , n18111 , n18430 );
and ( n26154 , n26152 , n26153 );
xor ( n26155 , n26152 , n26153 );
xor ( n26156 , n26063 , n26126 );
and ( n26157 , n18112 , n18430 );
and ( n26158 , n26156 , n26157 );
xor ( n26159 , n26156 , n26157 );
xor ( n26160 , n26067 , n26124 );
and ( n26161 , n18113 , n18430 );
and ( n26162 , n26160 , n26161 );
xor ( n26163 , n26160 , n26161 );
xor ( n26164 , n26071 , n26122 );
and ( n26165 , n18114 , n18430 );
and ( n26166 , n26164 , n26165 );
xor ( n26167 , n26164 , n26165 );
xor ( n26168 , n26075 , n26120 );
and ( n26169 , n18115 , n18430 );
and ( n26170 , n26168 , n26169 );
xor ( n26171 , n26168 , n26169 );
xor ( n26172 , n26079 , n26118 );
and ( n26173 , n18116 , n18430 );
and ( n26174 , n26172 , n26173 );
xor ( n26175 , n26172 , n26173 );
xor ( n26176 , n26083 , n26116 );
and ( n26177 , n18117 , n18430 );
and ( n26178 , n26176 , n26177 );
xor ( n26179 , n26176 , n26177 );
xor ( n26180 , n26087 , n26114 );
and ( n26181 , n18118 , n18430 );
and ( n26182 , n26180 , n26181 );
xor ( n26183 , n26180 , n26181 );
xor ( n26184 , n26091 , n26112 );
and ( n26185 , n18119 , n18430 );
and ( n26186 , n26184 , n26185 );
xor ( n26187 , n26184 , n26185 );
xor ( n26188 , n26095 , n26110 );
and ( n26189 , n18120 , n18430 );
and ( n26190 , n26188 , n26189 );
xor ( n26191 , n26188 , n26189 );
xor ( n26192 , n26099 , n26108 );
and ( n26193 , n18121 , n18430 );
and ( n26194 , n26192 , n26193 );
xor ( n26195 , n26192 , n26193 );
xor ( n26196 , n26103 , n26106 );
and ( n26197 , n18122 , n18430 );
and ( n26198 , n26196 , n26197 );
and ( n26199 , n26195 , n26198 );
or ( n26200 , n26194 , n26199 );
and ( n26201 , n26191 , n26200 );
or ( n26202 , n26190 , n26201 );
and ( n26203 , n26187 , n26202 );
or ( n26204 , n26186 , n26203 );
and ( n26205 , n26183 , n26204 );
or ( n26206 , n26182 , n26205 );
and ( n26207 , n26179 , n26206 );
or ( n26208 , n26178 , n26207 );
and ( n26209 , n26175 , n26208 );
or ( n26210 , n26174 , n26209 );
and ( n26211 , n26171 , n26210 );
or ( n26212 , n26170 , n26211 );
and ( n26213 , n26167 , n26212 );
or ( n26214 , n26166 , n26213 );
and ( n26215 , n26163 , n26214 );
or ( n26216 , n26162 , n26215 );
and ( n26217 , n26159 , n26216 );
or ( n26218 , n26158 , n26217 );
and ( n26219 , n26155 , n26218 );
or ( n26220 , n26154 , n26219 );
and ( n26221 , n26151 , n26220 );
or ( n26222 , n26150 , n26221 );
and ( n26223 , n26147 , n26222 );
or ( n26224 , n26146 , n26223 );
and ( n26225 , n26143 , n26224 );
or ( n26226 , n26142 , n26225 );
and ( n26227 , n26139 , n26226 );
or ( n26228 , n26138 , n26227 );
and ( n26229 , n18107 , n18428 );
and ( n26230 , n26228 , n26229 );
xor ( n26231 , n26228 , n26229 );
xor ( n26232 , n26139 , n26226 );
and ( n26233 , n18108 , n18428 );
and ( n26234 , n26232 , n26233 );
xor ( n26235 , n26232 , n26233 );
xor ( n26236 , n26143 , n26224 );
and ( n26237 , n18109 , n18428 );
and ( n26238 , n26236 , n26237 );
xor ( n26239 , n26236 , n26237 );
xor ( n26240 , n26147 , n26222 );
and ( n26241 , n18110 , n18428 );
and ( n26242 , n26240 , n26241 );
xor ( n26243 , n26240 , n26241 );
xor ( n26244 , n26151 , n26220 );
and ( n26245 , n18111 , n18428 );
and ( n26246 , n26244 , n26245 );
xor ( n26247 , n26244 , n26245 );
xor ( n26248 , n26155 , n26218 );
and ( n26249 , n18112 , n18428 );
and ( n26250 , n26248 , n26249 );
xor ( n26251 , n26248 , n26249 );
xor ( n26252 , n26159 , n26216 );
and ( n26253 , n18113 , n18428 );
and ( n26254 , n26252 , n26253 );
xor ( n26255 , n26252 , n26253 );
xor ( n26256 , n26163 , n26214 );
and ( n26257 , n18114 , n18428 );
and ( n26258 , n26256 , n26257 );
xor ( n26259 , n26256 , n26257 );
xor ( n26260 , n26167 , n26212 );
and ( n26261 , n18115 , n18428 );
and ( n26262 , n26260 , n26261 );
xor ( n26263 , n26260 , n26261 );
xor ( n26264 , n26171 , n26210 );
and ( n26265 , n18116 , n18428 );
and ( n26266 , n26264 , n26265 );
xor ( n26267 , n26264 , n26265 );
xor ( n26268 , n26175 , n26208 );
and ( n26269 , n18117 , n18428 );
and ( n26270 , n26268 , n26269 );
xor ( n26271 , n26268 , n26269 );
xor ( n26272 , n26179 , n26206 );
and ( n26273 , n18118 , n18428 );
and ( n26274 , n26272 , n26273 );
xor ( n26275 , n26272 , n26273 );
xor ( n26276 , n26183 , n26204 );
and ( n26277 , n18119 , n18428 );
and ( n26278 , n26276 , n26277 );
xor ( n26279 , n26276 , n26277 );
xor ( n26280 , n26187 , n26202 );
and ( n26281 , n18120 , n18428 );
and ( n26282 , n26280 , n26281 );
xor ( n26283 , n26280 , n26281 );
xor ( n26284 , n26191 , n26200 );
and ( n26285 , n18121 , n18428 );
and ( n26286 , n26284 , n26285 );
xor ( n26287 , n26284 , n26285 );
xor ( n26288 , n26195 , n26198 );
and ( n26289 , n18122 , n18428 );
and ( n26290 , n26288 , n26289 );
and ( n26291 , n26287 , n26290 );
or ( n26292 , n26286 , n26291 );
and ( n26293 , n26283 , n26292 );
or ( n26294 , n26282 , n26293 );
and ( n26295 , n26279 , n26294 );
or ( n26296 , n26278 , n26295 );
and ( n26297 , n26275 , n26296 );
or ( n26298 , n26274 , n26297 );
and ( n26299 , n26271 , n26298 );
or ( n26300 , n26270 , n26299 );
and ( n26301 , n26267 , n26300 );
or ( n26302 , n26266 , n26301 );
and ( n26303 , n26263 , n26302 );
or ( n26304 , n26262 , n26303 );
and ( n26305 , n26259 , n26304 );
or ( n26306 , n26258 , n26305 );
and ( n26307 , n26255 , n26306 );
or ( n26308 , n26254 , n26307 );
and ( n26309 , n26251 , n26308 );
or ( n26310 , n26250 , n26309 );
and ( n26311 , n26247 , n26310 );
or ( n26312 , n26246 , n26311 );
and ( n26313 , n26243 , n26312 );
or ( n26314 , n26242 , n26313 );
and ( n26315 , n26239 , n26314 );
or ( n26316 , n26238 , n26315 );
and ( n26317 , n26235 , n26316 );
or ( n26318 , n26234 , n26317 );
and ( n26319 , n26231 , n26318 );
or ( n26320 , n26230 , n26319 );
and ( n26321 , n18107 , n18426 );
and ( n26322 , n26320 , n26321 );
xor ( n26323 , n26320 , n26321 );
xor ( n26324 , n26231 , n26318 );
and ( n26325 , n18108 , n18426 );
and ( n26326 , n26324 , n26325 );
xor ( n26327 , n26324 , n26325 );
xor ( n26328 , n26235 , n26316 );
and ( n26329 , n18109 , n18426 );
and ( n26330 , n26328 , n26329 );
xor ( n26331 , n26328 , n26329 );
xor ( n26332 , n26239 , n26314 );
and ( n26333 , n18110 , n18426 );
and ( n26334 , n26332 , n26333 );
xor ( n26335 , n26332 , n26333 );
xor ( n26336 , n26243 , n26312 );
and ( n26337 , n18111 , n18426 );
and ( n26338 , n26336 , n26337 );
xor ( n26339 , n26336 , n26337 );
xor ( n26340 , n26247 , n26310 );
and ( n26341 , n18112 , n18426 );
and ( n26342 , n26340 , n26341 );
xor ( n26343 , n26340 , n26341 );
xor ( n26344 , n26251 , n26308 );
and ( n26345 , n18113 , n18426 );
and ( n26346 , n26344 , n26345 );
xor ( n26347 , n26344 , n26345 );
xor ( n26348 , n26255 , n26306 );
and ( n26349 , n18114 , n18426 );
and ( n26350 , n26348 , n26349 );
xor ( n26351 , n26348 , n26349 );
xor ( n26352 , n26259 , n26304 );
and ( n26353 , n18115 , n18426 );
and ( n26354 , n26352 , n26353 );
xor ( n26355 , n26352 , n26353 );
xor ( n26356 , n26263 , n26302 );
and ( n26357 , n18116 , n18426 );
and ( n26358 , n26356 , n26357 );
xor ( n26359 , n26356 , n26357 );
xor ( n26360 , n26267 , n26300 );
and ( n26361 , n18117 , n18426 );
and ( n26362 , n26360 , n26361 );
xor ( n26363 , n26360 , n26361 );
xor ( n26364 , n26271 , n26298 );
and ( n26365 , n18118 , n18426 );
and ( n26366 , n26364 , n26365 );
xor ( n26367 , n26364 , n26365 );
xor ( n26368 , n26275 , n26296 );
and ( n26369 , n18119 , n18426 );
and ( n26370 , n26368 , n26369 );
xor ( n26371 , n26368 , n26369 );
xor ( n26372 , n26279 , n26294 );
and ( n26373 , n18120 , n18426 );
and ( n26374 , n26372 , n26373 );
xor ( n26375 , n26372 , n26373 );
xor ( n26376 , n26283 , n26292 );
and ( n26377 , n18121 , n18426 );
and ( n26378 , n26376 , n26377 );
xor ( n26379 , n26376 , n26377 );
xor ( n26380 , n26287 , n26290 );
and ( n26381 , n18122 , n18426 );
and ( n26382 , n26380 , n26381 );
and ( n26383 , n26379 , n26382 );
or ( n26384 , n26378 , n26383 );
and ( n26385 , n26375 , n26384 );
or ( n26386 , n26374 , n26385 );
and ( n26387 , n26371 , n26386 );
or ( n26388 , n26370 , n26387 );
and ( n26389 , n26367 , n26388 );
or ( n26390 , n26366 , n26389 );
and ( n26391 , n26363 , n26390 );
or ( n26392 , n26362 , n26391 );
and ( n26393 , n26359 , n26392 );
or ( n26394 , n26358 , n26393 );
and ( n26395 , n26355 , n26394 );
or ( n26396 , n26354 , n26395 );
and ( n26397 , n26351 , n26396 );
or ( n26398 , n26350 , n26397 );
and ( n26399 , n26347 , n26398 );
or ( n26400 , n26346 , n26399 );
and ( n26401 , n26343 , n26400 );
or ( n26402 , n26342 , n26401 );
and ( n26403 , n26339 , n26402 );
or ( n26404 , n26338 , n26403 );
and ( n26405 , n26335 , n26404 );
or ( n26406 , n26334 , n26405 );
and ( n26407 , n26331 , n26406 );
or ( n26408 , n26330 , n26407 );
and ( n26409 , n26327 , n26408 );
or ( n26410 , n26326 , n26409 );
and ( n26411 , n26323 , n26410 );
or ( n26412 , n26322 , n26411 );
and ( n26413 , n18107 , n18424 );
and ( n26414 , n26412 , n26413 );
xor ( n26415 , n26412 , n26413 );
xor ( n26416 , n26323 , n26410 );
and ( n26417 , n18108 , n18424 );
and ( n26418 , n26416 , n26417 );
xor ( n26419 , n26416 , n26417 );
xor ( n26420 , n26327 , n26408 );
and ( n26421 , n18109 , n18424 );
and ( n26422 , n26420 , n26421 );
xor ( n26423 , n26420 , n26421 );
xor ( n26424 , n26331 , n26406 );
and ( n26425 , n18110 , n18424 );
and ( n26426 , n26424 , n26425 );
xor ( n26427 , n26424 , n26425 );
xor ( n26428 , n26335 , n26404 );
and ( n26429 , n18111 , n18424 );
and ( n26430 , n26428 , n26429 );
xor ( n26431 , n26428 , n26429 );
xor ( n26432 , n26339 , n26402 );
and ( n26433 , n18112 , n18424 );
and ( n26434 , n26432 , n26433 );
xor ( n26435 , n26432 , n26433 );
xor ( n26436 , n26343 , n26400 );
and ( n26437 , n18113 , n18424 );
and ( n26438 , n26436 , n26437 );
xor ( n26439 , n26436 , n26437 );
xor ( n26440 , n26347 , n26398 );
and ( n26441 , n18114 , n18424 );
and ( n26442 , n26440 , n26441 );
xor ( n26443 , n26440 , n26441 );
xor ( n26444 , n26351 , n26396 );
and ( n26445 , n18115 , n18424 );
and ( n26446 , n26444 , n26445 );
xor ( n26447 , n26444 , n26445 );
xor ( n26448 , n26355 , n26394 );
and ( n26449 , n18116 , n18424 );
and ( n26450 , n26448 , n26449 );
xor ( n26451 , n26448 , n26449 );
xor ( n26452 , n26359 , n26392 );
and ( n26453 , n18117 , n18424 );
and ( n26454 , n26452 , n26453 );
xor ( n26455 , n26452 , n26453 );
xor ( n26456 , n26363 , n26390 );
and ( n26457 , n18118 , n18424 );
and ( n26458 , n26456 , n26457 );
xor ( n26459 , n26456 , n26457 );
xor ( n26460 , n26367 , n26388 );
and ( n26461 , n18119 , n18424 );
and ( n26462 , n26460 , n26461 );
xor ( n26463 , n26460 , n26461 );
xor ( n26464 , n26371 , n26386 );
and ( n26465 , n18120 , n18424 );
and ( n26466 , n26464 , n26465 );
xor ( n26467 , n26464 , n26465 );
xor ( n26468 , n26375 , n26384 );
and ( n26469 , n18121 , n18424 );
and ( n26470 , n26468 , n26469 );
xor ( n26471 , n26468 , n26469 );
xor ( n26472 , n26379 , n26382 );
and ( n26473 , n18122 , n18424 );
and ( n26474 , n26472 , n26473 );
and ( n26475 , n26471 , n26474 );
or ( n26476 , n26470 , n26475 );
and ( n26477 , n26467 , n26476 );
or ( n26478 , n26466 , n26477 );
and ( n26479 , n26463 , n26478 );
or ( n26480 , n26462 , n26479 );
and ( n26481 , n26459 , n26480 );
or ( n26482 , n26458 , n26481 );
and ( n26483 , n26455 , n26482 );
or ( n26484 , n26454 , n26483 );
and ( n26485 , n26451 , n26484 );
or ( n26486 , n26450 , n26485 );
and ( n26487 , n26447 , n26486 );
or ( n26488 , n26446 , n26487 );
and ( n26489 , n26443 , n26488 );
or ( n26490 , n26442 , n26489 );
and ( n26491 , n26439 , n26490 );
or ( n26492 , n26438 , n26491 );
and ( n26493 , n26435 , n26492 );
or ( n26494 , n26434 , n26493 );
and ( n26495 , n26431 , n26494 );
or ( n26496 , n26430 , n26495 );
and ( n26497 , n26427 , n26496 );
or ( n26498 , n26426 , n26497 );
and ( n26499 , n26423 , n26498 );
or ( n26500 , n26422 , n26499 );
and ( n26501 , n26419 , n26500 );
or ( n26502 , n26418 , n26501 );
and ( n26503 , n26415 , n26502 );
or ( n26504 , n26414 , n26503 );
and ( n26505 , n18107 , n18422 );
and ( n26506 , n26504 , n26505 );
xor ( n26507 , n26504 , n26505 );
xor ( n26508 , n26415 , n26502 );
and ( n26509 , n18108 , n18422 );
and ( n26510 , n26508 , n26509 );
xor ( n26511 , n26508 , n26509 );
xor ( n26512 , n26419 , n26500 );
and ( n26513 , n18109 , n18422 );
and ( n26514 , n26512 , n26513 );
xor ( n26515 , n26512 , n26513 );
xor ( n26516 , n26423 , n26498 );
and ( n26517 , n18110 , n18422 );
and ( n26518 , n26516 , n26517 );
xor ( n26519 , n26516 , n26517 );
xor ( n26520 , n26427 , n26496 );
and ( n26521 , n18111 , n18422 );
and ( n26522 , n26520 , n26521 );
xor ( n26523 , n26520 , n26521 );
xor ( n26524 , n26431 , n26494 );
and ( n26525 , n18112 , n18422 );
and ( n26526 , n26524 , n26525 );
xor ( n26527 , n26524 , n26525 );
xor ( n26528 , n26435 , n26492 );
and ( n26529 , n18113 , n18422 );
and ( n26530 , n26528 , n26529 );
xor ( n26531 , n26528 , n26529 );
xor ( n26532 , n26439 , n26490 );
and ( n26533 , n18114 , n18422 );
and ( n26534 , n26532 , n26533 );
xor ( n26535 , n26532 , n26533 );
xor ( n26536 , n26443 , n26488 );
and ( n26537 , n18115 , n18422 );
and ( n26538 , n26536 , n26537 );
xor ( n26539 , n26536 , n26537 );
xor ( n26540 , n26447 , n26486 );
and ( n26541 , n18116 , n18422 );
and ( n26542 , n26540 , n26541 );
xor ( n26543 , n26540 , n26541 );
xor ( n26544 , n26451 , n26484 );
and ( n26545 , n18117 , n18422 );
and ( n26546 , n26544 , n26545 );
xor ( n26547 , n26544 , n26545 );
xor ( n26548 , n26455 , n26482 );
and ( n26549 , n18118 , n18422 );
and ( n26550 , n26548 , n26549 );
xor ( n26551 , n26548 , n26549 );
xor ( n26552 , n26459 , n26480 );
and ( n26553 , n18119 , n18422 );
and ( n26554 , n26552 , n26553 );
xor ( n26555 , n26552 , n26553 );
xor ( n26556 , n26463 , n26478 );
and ( n26557 , n18120 , n18422 );
and ( n26558 , n26556 , n26557 );
xor ( n26559 , n26556 , n26557 );
xor ( n26560 , n26467 , n26476 );
and ( n26561 , n18121 , n18422 );
and ( n26562 , n26560 , n26561 );
xor ( n26563 , n26560 , n26561 );
xor ( n26564 , n26471 , n26474 );
and ( n26565 , n18122 , n18422 );
and ( n26566 , n26564 , n26565 );
and ( n26567 , n26563 , n26566 );
or ( n26568 , n26562 , n26567 );
and ( n26569 , n26559 , n26568 );
or ( n26570 , n26558 , n26569 );
and ( n26571 , n26555 , n26570 );
or ( n26572 , n26554 , n26571 );
and ( n26573 , n26551 , n26572 );
or ( n26574 , n26550 , n26573 );
and ( n26575 , n26547 , n26574 );
or ( n26576 , n26546 , n26575 );
and ( n26577 , n26543 , n26576 );
or ( n26578 , n26542 , n26577 );
and ( n26579 , n26539 , n26578 );
or ( n26580 , n26538 , n26579 );
and ( n26581 , n26535 , n26580 );
or ( n26582 , n26534 , n26581 );
and ( n26583 , n26531 , n26582 );
or ( n26584 , n26530 , n26583 );
and ( n26585 , n26527 , n26584 );
or ( n26586 , n26526 , n26585 );
and ( n26587 , n26523 , n26586 );
or ( n26588 , n26522 , n26587 );
and ( n26589 , n26519 , n26588 );
or ( n26590 , n26518 , n26589 );
and ( n26591 , n26515 , n26590 );
or ( n26592 , n26514 , n26591 );
and ( n26593 , n26511 , n26592 );
or ( n26594 , n26510 , n26593 );
and ( n26595 , n26507 , n26594 );
or ( n26596 , n26506 , n26595 );
and ( n26597 , n18107 , n18420 );
and ( n26598 , n26596 , n26597 );
xor ( n26599 , n26596 , n26597 );
xor ( n26600 , n26507 , n26594 );
and ( n26601 , n18108 , n18420 );
and ( n26602 , n26600 , n26601 );
xor ( n26603 , n26600 , n26601 );
xor ( n26604 , n26511 , n26592 );
and ( n26605 , n18109 , n18420 );
and ( n26606 , n26604 , n26605 );
xor ( n26607 , n26604 , n26605 );
xor ( n26608 , n26515 , n26590 );
and ( n26609 , n18110 , n18420 );
and ( n26610 , n26608 , n26609 );
xor ( n26611 , n26608 , n26609 );
xor ( n26612 , n26519 , n26588 );
and ( n26613 , n18111 , n18420 );
and ( n26614 , n26612 , n26613 );
xor ( n26615 , n26612 , n26613 );
xor ( n26616 , n26523 , n26586 );
and ( n26617 , n18112 , n18420 );
and ( n26618 , n26616 , n26617 );
xor ( n26619 , n26616 , n26617 );
xor ( n26620 , n26527 , n26584 );
and ( n26621 , n18113 , n18420 );
and ( n26622 , n26620 , n26621 );
xor ( n26623 , n26620 , n26621 );
xor ( n26624 , n26531 , n26582 );
and ( n26625 , n18114 , n18420 );
and ( n26626 , n26624 , n26625 );
xor ( n26627 , n26624 , n26625 );
xor ( n26628 , n26535 , n26580 );
and ( n26629 , n18115 , n18420 );
and ( n26630 , n26628 , n26629 );
xor ( n26631 , n26628 , n26629 );
xor ( n26632 , n26539 , n26578 );
and ( n26633 , n18116 , n18420 );
and ( n26634 , n26632 , n26633 );
xor ( n26635 , n26632 , n26633 );
xor ( n26636 , n26543 , n26576 );
and ( n26637 , n18117 , n18420 );
and ( n26638 , n26636 , n26637 );
xor ( n26639 , n26636 , n26637 );
xor ( n26640 , n26547 , n26574 );
and ( n26641 , n18118 , n18420 );
and ( n26642 , n26640 , n26641 );
xor ( n26643 , n26640 , n26641 );
xor ( n26644 , n26551 , n26572 );
and ( n26645 , n18119 , n18420 );
and ( n26646 , n26644 , n26645 );
xor ( n26647 , n26644 , n26645 );
xor ( n26648 , n26555 , n26570 );
and ( n26649 , n18120 , n18420 );
and ( n26650 , n26648 , n26649 );
xor ( n26651 , n26648 , n26649 );
xor ( n26652 , n26559 , n26568 );
and ( n26653 , n18121 , n18420 );
and ( n26654 , n26652 , n26653 );
xor ( n26655 , n26652 , n26653 );
xor ( n26656 , n26563 , n26566 );
and ( n26657 , n18122 , n18420 );
and ( n26658 , n26656 , n26657 );
and ( n26659 , n26655 , n26658 );
or ( n26660 , n26654 , n26659 );
and ( n26661 , n26651 , n26660 );
or ( n26662 , n26650 , n26661 );
and ( n26663 , n26647 , n26662 );
or ( n26664 , n26646 , n26663 );
and ( n26665 , n26643 , n26664 );
or ( n26666 , n26642 , n26665 );
and ( n26667 , n26639 , n26666 );
or ( n26668 , n26638 , n26667 );
and ( n26669 , n26635 , n26668 );
or ( n26670 , n26634 , n26669 );
and ( n26671 , n26631 , n26670 );
or ( n26672 , n26630 , n26671 );
and ( n26673 , n26627 , n26672 );
or ( n26674 , n26626 , n26673 );
and ( n26675 , n26623 , n26674 );
or ( n26676 , n26622 , n26675 );
and ( n26677 , n26619 , n26676 );
or ( n26678 , n26618 , n26677 );
and ( n26679 , n26615 , n26678 );
or ( n26680 , n26614 , n26679 );
and ( n26681 , n26611 , n26680 );
or ( n26682 , n26610 , n26681 );
and ( n26683 , n26607 , n26682 );
or ( n26684 , n26606 , n26683 );
and ( n26685 , n26603 , n26684 );
or ( n26686 , n26602 , n26685 );
and ( n26687 , n26599 , n26686 );
or ( n26688 , n26598 , n26687 );
and ( n26689 , n18107 , n18418 );
and ( n26690 , n26688 , n26689 );
xor ( n26691 , n26688 , n26689 );
xor ( n26692 , n26599 , n26686 );
and ( n26693 , n18108 , n18418 );
and ( n26694 , n26692 , n26693 );
xor ( n26695 , n26692 , n26693 );
xor ( n26696 , n26603 , n26684 );
and ( n26697 , n18109 , n18418 );
and ( n26698 , n26696 , n26697 );
xor ( n26699 , n26696 , n26697 );
xor ( n26700 , n26607 , n26682 );
and ( n26701 , n18110 , n18418 );
and ( n26702 , n26700 , n26701 );
xor ( n26703 , n26700 , n26701 );
xor ( n26704 , n26611 , n26680 );
and ( n26705 , n18111 , n18418 );
and ( n26706 , n26704 , n26705 );
xor ( n26707 , n26704 , n26705 );
xor ( n26708 , n26615 , n26678 );
and ( n26709 , n18112 , n18418 );
and ( n26710 , n26708 , n26709 );
xor ( n26711 , n26708 , n26709 );
xor ( n26712 , n26619 , n26676 );
and ( n26713 , n18113 , n18418 );
and ( n26714 , n26712 , n26713 );
xor ( n26715 , n26712 , n26713 );
xor ( n26716 , n26623 , n26674 );
and ( n26717 , n18114 , n18418 );
and ( n26718 , n26716 , n26717 );
xor ( n26719 , n26716 , n26717 );
xor ( n26720 , n26627 , n26672 );
and ( n26721 , n18115 , n18418 );
and ( n26722 , n26720 , n26721 );
xor ( n26723 , n26720 , n26721 );
xor ( n26724 , n26631 , n26670 );
and ( n26725 , n18116 , n18418 );
and ( n26726 , n26724 , n26725 );
xor ( n26727 , n26724 , n26725 );
xor ( n26728 , n26635 , n26668 );
and ( n26729 , n18117 , n18418 );
and ( n26730 , n26728 , n26729 );
xor ( n26731 , n26728 , n26729 );
xor ( n26732 , n26639 , n26666 );
and ( n26733 , n18118 , n18418 );
and ( n26734 , n26732 , n26733 );
xor ( n26735 , n26732 , n26733 );
xor ( n26736 , n26643 , n26664 );
and ( n26737 , n18119 , n18418 );
and ( n26738 , n26736 , n26737 );
xor ( n26739 , n26736 , n26737 );
xor ( n26740 , n26647 , n26662 );
and ( n26741 , n18120 , n18418 );
and ( n26742 , n26740 , n26741 );
xor ( n26743 , n26740 , n26741 );
xor ( n26744 , n26651 , n26660 );
and ( n26745 , n18121 , n18418 );
and ( n26746 , n26744 , n26745 );
xor ( n26747 , n26744 , n26745 );
xor ( n26748 , n26655 , n26658 );
and ( n26749 , n18122 , n18418 );
and ( n26750 , n26748 , n26749 );
and ( n26751 , n26747 , n26750 );
or ( n26752 , n26746 , n26751 );
and ( n26753 , n26743 , n26752 );
or ( n26754 , n26742 , n26753 );
and ( n26755 , n26739 , n26754 );
or ( n26756 , n26738 , n26755 );
and ( n26757 , n26735 , n26756 );
or ( n26758 , n26734 , n26757 );
and ( n26759 , n26731 , n26758 );
or ( n26760 , n26730 , n26759 );
and ( n26761 , n26727 , n26760 );
or ( n26762 , n26726 , n26761 );
and ( n26763 , n26723 , n26762 );
or ( n26764 , n26722 , n26763 );
and ( n26765 , n26719 , n26764 );
or ( n26766 , n26718 , n26765 );
and ( n26767 , n26715 , n26766 );
or ( n26768 , n26714 , n26767 );
and ( n26769 , n26711 , n26768 );
or ( n26770 , n26710 , n26769 );
and ( n26771 , n26707 , n26770 );
or ( n26772 , n26706 , n26771 );
and ( n26773 , n26703 , n26772 );
or ( n26774 , n26702 , n26773 );
and ( n26775 , n26699 , n26774 );
or ( n26776 , n26698 , n26775 );
and ( n26777 , n26695 , n26776 );
or ( n26778 , n26694 , n26777 );
and ( n26779 , n26691 , n26778 );
or ( n26780 , n26690 , n26779 );
and ( n26781 , n18107 , n18416 );
and ( n26782 , n26780 , n26781 );
xor ( n26783 , n26780 , n26781 );
xor ( n26784 , n26691 , n26778 );
and ( n26785 , n18108 , n18416 );
and ( n26786 , n26784 , n26785 );
xor ( n26787 , n26784 , n26785 );
xor ( n26788 , n26695 , n26776 );
and ( n26789 , n18109 , n18416 );
and ( n26790 , n26788 , n26789 );
xor ( n26791 , n26788 , n26789 );
xor ( n26792 , n26699 , n26774 );
and ( n26793 , n18110 , n18416 );
and ( n26794 , n26792 , n26793 );
xor ( n26795 , n26792 , n26793 );
xor ( n26796 , n26703 , n26772 );
and ( n26797 , n18111 , n18416 );
and ( n26798 , n26796 , n26797 );
xor ( n26799 , n26796 , n26797 );
xor ( n26800 , n26707 , n26770 );
and ( n26801 , n18112 , n18416 );
and ( n26802 , n26800 , n26801 );
xor ( n26803 , n26800 , n26801 );
xor ( n26804 , n26711 , n26768 );
and ( n26805 , n18113 , n18416 );
and ( n26806 , n26804 , n26805 );
xor ( n26807 , n26804 , n26805 );
xor ( n26808 , n26715 , n26766 );
and ( n26809 , n18114 , n18416 );
and ( n26810 , n26808 , n26809 );
xor ( n26811 , n26808 , n26809 );
xor ( n26812 , n26719 , n26764 );
and ( n26813 , n18115 , n18416 );
and ( n26814 , n26812 , n26813 );
xor ( n26815 , n26812 , n26813 );
xor ( n26816 , n26723 , n26762 );
and ( n26817 , n18116 , n18416 );
and ( n26818 , n26816 , n26817 );
xor ( n26819 , n26816 , n26817 );
xor ( n26820 , n26727 , n26760 );
and ( n26821 , n18117 , n18416 );
and ( n26822 , n26820 , n26821 );
xor ( n26823 , n26820 , n26821 );
xor ( n26824 , n26731 , n26758 );
and ( n26825 , n18118 , n18416 );
and ( n26826 , n26824 , n26825 );
xor ( n26827 , n26824 , n26825 );
xor ( n26828 , n26735 , n26756 );
and ( n26829 , n18119 , n18416 );
and ( n26830 , n26828 , n26829 );
xor ( n26831 , n26828 , n26829 );
xor ( n26832 , n26739 , n26754 );
and ( n26833 , n18120 , n18416 );
and ( n26834 , n26832 , n26833 );
xor ( n26835 , n26832 , n26833 );
xor ( n26836 , n26743 , n26752 );
and ( n26837 , n18121 , n18416 );
and ( n26838 , n26836 , n26837 );
xor ( n26839 , n26836 , n26837 );
xor ( n26840 , n26747 , n26750 );
and ( n26841 , n18122 , n18416 );
and ( n26842 , n26840 , n26841 );
and ( n26843 , n26839 , n26842 );
or ( n26844 , n26838 , n26843 );
and ( n26845 , n26835 , n26844 );
or ( n26846 , n26834 , n26845 );
and ( n26847 , n26831 , n26846 );
or ( n26848 , n26830 , n26847 );
and ( n26849 , n26827 , n26848 );
or ( n26850 , n26826 , n26849 );
and ( n26851 , n26823 , n26850 );
or ( n26852 , n26822 , n26851 );
and ( n26853 , n26819 , n26852 );
or ( n26854 , n26818 , n26853 );
and ( n26855 , n26815 , n26854 );
or ( n26856 , n26814 , n26855 );
and ( n26857 , n26811 , n26856 );
or ( n26858 , n26810 , n26857 );
and ( n26859 , n26807 , n26858 );
or ( n26860 , n26806 , n26859 );
and ( n26861 , n26803 , n26860 );
or ( n26862 , n26802 , n26861 );
and ( n26863 , n26799 , n26862 );
or ( n26864 , n26798 , n26863 );
and ( n26865 , n26795 , n26864 );
or ( n26866 , n26794 , n26865 );
and ( n26867 , n26791 , n26866 );
or ( n26868 , n26790 , n26867 );
and ( n26869 , n26787 , n26868 );
or ( n26870 , n26786 , n26869 );
and ( n26871 , n26783 , n26870 );
or ( n26872 , n26782 , n26871 );
and ( n26873 , n18107 , n18414 );
and ( n26874 , n26872 , n26873 );
xor ( n26875 , n26872 , n26873 );
xor ( n26876 , n26783 , n26870 );
and ( n26877 , n18108 , n18414 );
and ( n26878 , n26876 , n26877 );
xor ( n26879 , n26876 , n26877 );
xor ( n26880 , n26787 , n26868 );
and ( n26881 , n18109 , n18414 );
and ( n26882 , n26880 , n26881 );
xor ( n26883 , n26880 , n26881 );
xor ( n26884 , n26791 , n26866 );
and ( n26885 , n18110 , n18414 );
and ( n26886 , n26884 , n26885 );
xor ( n26887 , n26884 , n26885 );
xor ( n26888 , n26795 , n26864 );
and ( n26889 , n18111 , n18414 );
and ( n26890 , n26888 , n26889 );
xor ( n26891 , n26888 , n26889 );
xor ( n26892 , n26799 , n26862 );
and ( n26893 , n18112 , n18414 );
and ( n26894 , n26892 , n26893 );
xor ( n26895 , n26892 , n26893 );
xor ( n26896 , n26803 , n26860 );
and ( n26897 , n18113 , n18414 );
and ( n26898 , n26896 , n26897 );
xor ( n26899 , n26896 , n26897 );
xor ( n26900 , n26807 , n26858 );
and ( n26901 , n18114 , n18414 );
and ( n26902 , n26900 , n26901 );
xor ( n26903 , n26900 , n26901 );
xor ( n26904 , n26811 , n26856 );
and ( n26905 , n18115 , n18414 );
and ( n26906 , n26904 , n26905 );
xor ( n26907 , n26904 , n26905 );
xor ( n26908 , n26815 , n26854 );
and ( n26909 , n18116 , n18414 );
and ( n26910 , n26908 , n26909 );
xor ( n26911 , n26908 , n26909 );
xor ( n26912 , n26819 , n26852 );
and ( n26913 , n18117 , n18414 );
and ( n26914 , n26912 , n26913 );
xor ( n26915 , n26912 , n26913 );
xor ( n26916 , n26823 , n26850 );
and ( n26917 , n18118 , n18414 );
and ( n26918 , n26916 , n26917 );
xor ( n26919 , n26916 , n26917 );
xor ( n26920 , n26827 , n26848 );
and ( n26921 , n18119 , n18414 );
and ( n26922 , n26920 , n26921 );
xor ( n26923 , n26920 , n26921 );
xor ( n26924 , n26831 , n26846 );
and ( n26925 , n18120 , n18414 );
and ( n26926 , n26924 , n26925 );
xor ( n26927 , n26924 , n26925 );
xor ( n26928 , n26835 , n26844 );
and ( n26929 , n18121 , n18414 );
and ( n26930 , n26928 , n26929 );
xor ( n26931 , n26928 , n26929 );
xor ( n26932 , n26839 , n26842 );
and ( n26933 , n18122 , n18414 );
and ( n26934 , n26932 , n26933 );
and ( n26935 , n26931 , n26934 );
or ( n26936 , n26930 , n26935 );
and ( n26937 , n26927 , n26936 );
or ( n26938 , n26926 , n26937 );
and ( n26939 , n26923 , n26938 );
or ( n26940 , n26922 , n26939 );
and ( n26941 , n26919 , n26940 );
or ( n26942 , n26918 , n26941 );
and ( n26943 , n26915 , n26942 );
or ( n26944 , n26914 , n26943 );
and ( n26945 , n26911 , n26944 );
or ( n26946 , n26910 , n26945 );
and ( n26947 , n26907 , n26946 );
or ( n26948 , n26906 , n26947 );
and ( n26949 , n26903 , n26948 );
or ( n26950 , n26902 , n26949 );
and ( n26951 , n26899 , n26950 );
or ( n26952 , n26898 , n26951 );
and ( n26953 , n26895 , n26952 );
or ( n26954 , n26894 , n26953 );
and ( n26955 , n26891 , n26954 );
or ( n26956 , n26890 , n26955 );
and ( n26957 , n26887 , n26956 );
or ( n26958 , n26886 , n26957 );
and ( n26959 , n26883 , n26958 );
or ( n26960 , n26882 , n26959 );
and ( n26961 , n26879 , n26960 );
or ( n26962 , n26878 , n26961 );
and ( n26963 , n26875 , n26962 );
or ( n26964 , n26874 , n26963 );
and ( n26965 , n18107 , n18412 );
and ( n26966 , n26964 , n26965 );
xor ( n26967 , n26964 , n26965 );
xor ( n26968 , n26875 , n26962 );
and ( n26969 , n18108 , n18412 );
and ( n26970 , n26968 , n26969 );
xor ( n26971 , n26968 , n26969 );
xor ( n26972 , n26879 , n26960 );
and ( n26973 , n18109 , n18412 );
and ( n26974 , n26972 , n26973 );
xor ( n26975 , n26972 , n26973 );
xor ( n26976 , n26883 , n26958 );
and ( n26977 , n18110 , n18412 );
and ( n26978 , n26976 , n26977 );
xor ( n26979 , n26976 , n26977 );
xor ( n26980 , n26887 , n26956 );
and ( n26981 , n18111 , n18412 );
and ( n26982 , n26980 , n26981 );
xor ( n26983 , n26980 , n26981 );
xor ( n26984 , n26891 , n26954 );
and ( n26985 , n18112 , n18412 );
and ( n26986 , n26984 , n26985 );
xor ( n26987 , n26984 , n26985 );
xor ( n26988 , n26895 , n26952 );
and ( n26989 , n18113 , n18412 );
and ( n26990 , n26988 , n26989 );
xor ( n26991 , n26988 , n26989 );
xor ( n26992 , n26899 , n26950 );
and ( n26993 , n18114 , n18412 );
and ( n26994 , n26992 , n26993 );
xor ( n26995 , n26992 , n26993 );
xor ( n26996 , n26903 , n26948 );
and ( n26997 , n18115 , n18412 );
and ( n26998 , n26996 , n26997 );
xor ( n26999 , n26996 , n26997 );
xor ( n27000 , n26907 , n26946 );
and ( n27001 , n18116 , n18412 );
and ( n27002 , n27000 , n27001 );
xor ( n27003 , n27000 , n27001 );
xor ( n27004 , n26911 , n26944 );
and ( n27005 , n18117 , n18412 );
and ( n27006 , n27004 , n27005 );
xor ( n27007 , n27004 , n27005 );
xor ( n27008 , n26915 , n26942 );
and ( n27009 , n18118 , n18412 );
and ( n27010 , n27008 , n27009 );
xor ( n27011 , n27008 , n27009 );
xor ( n27012 , n26919 , n26940 );
and ( n27013 , n18119 , n18412 );
and ( n27014 , n27012 , n27013 );
xor ( n27015 , n27012 , n27013 );
xor ( n27016 , n26923 , n26938 );
and ( n27017 , n18120 , n18412 );
and ( n27018 , n27016 , n27017 );
xor ( n27019 , n27016 , n27017 );
xor ( n27020 , n26927 , n26936 );
and ( n27021 , n18121 , n18412 );
and ( n27022 , n27020 , n27021 );
xor ( n27023 , n27020 , n27021 );
xor ( n27024 , n26931 , n26934 );
and ( n27025 , n18122 , n18412 );
and ( n27026 , n27024 , n27025 );
and ( n27027 , n27023 , n27026 );
or ( n27028 , n27022 , n27027 );
and ( n27029 , n27019 , n27028 );
or ( n27030 , n27018 , n27029 );
and ( n27031 , n27015 , n27030 );
or ( n27032 , n27014 , n27031 );
and ( n27033 , n27011 , n27032 );
or ( n27034 , n27010 , n27033 );
and ( n27035 , n27007 , n27034 );
or ( n27036 , n27006 , n27035 );
and ( n27037 , n27003 , n27036 );
or ( n27038 , n27002 , n27037 );
and ( n27039 , n26999 , n27038 );
or ( n27040 , n26998 , n27039 );
and ( n27041 , n26995 , n27040 );
or ( n27042 , n26994 , n27041 );
and ( n27043 , n26991 , n27042 );
or ( n27044 , n26990 , n27043 );
and ( n27045 , n26987 , n27044 );
or ( n27046 , n26986 , n27045 );
and ( n27047 , n26983 , n27046 );
or ( n27048 , n26982 , n27047 );
and ( n27049 , n26979 , n27048 );
or ( n27050 , n26978 , n27049 );
and ( n27051 , n26975 , n27050 );
or ( n27052 , n26974 , n27051 );
and ( n27053 , n26971 , n27052 );
or ( n27054 , n26970 , n27053 );
and ( n27055 , n26967 , n27054 );
or ( n27056 , n26966 , n27055 );
and ( n27057 , n18107 , n18410 );
and ( n27058 , n27056 , n27057 );
xor ( n27059 , n27056 , n27057 );
xor ( n27060 , n26967 , n27054 );
and ( n27061 , n18108 , n18410 );
and ( n27062 , n27060 , n27061 );
xor ( n27063 , n27060 , n27061 );
xor ( n27064 , n26971 , n27052 );
and ( n27065 , n18109 , n18410 );
and ( n27066 , n27064 , n27065 );
xor ( n27067 , n27064 , n27065 );
xor ( n27068 , n26975 , n27050 );
and ( n27069 , n18110 , n18410 );
and ( n27070 , n27068 , n27069 );
xor ( n27071 , n27068 , n27069 );
xor ( n27072 , n26979 , n27048 );
and ( n27073 , n18111 , n18410 );
and ( n27074 , n27072 , n27073 );
xor ( n27075 , n27072 , n27073 );
xor ( n27076 , n26983 , n27046 );
and ( n27077 , n18112 , n18410 );
and ( n27078 , n27076 , n27077 );
xor ( n27079 , n27076 , n27077 );
xor ( n27080 , n26987 , n27044 );
and ( n27081 , n18113 , n18410 );
and ( n27082 , n27080 , n27081 );
xor ( n27083 , n27080 , n27081 );
xor ( n27084 , n26991 , n27042 );
and ( n27085 , n18114 , n18410 );
and ( n27086 , n27084 , n27085 );
xor ( n27087 , n27084 , n27085 );
xor ( n27088 , n26995 , n27040 );
and ( n27089 , n18115 , n18410 );
and ( n27090 , n27088 , n27089 );
xor ( n27091 , n27088 , n27089 );
xor ( n27092 , n26999 , n27038 );
and ( n27093 , n18116 , n18410 );
and ( n27094 , n27092 , n27093 );
xor ( n27095 , n27092 , n27093 );
xor ( n27096 , n27003 , n27036 );
and ( n27097 , n18117 , n18410 );
and ( n27098 , n27096 , n27097 );
xor ( n27099 , n27096 , n27097 );
xor ( n27100 , n27007 , n27034 );
and ( n27101 , n18118 , n18410 );
and ( n27102 , n27100 , n27101 );
xor ( n27103 , n27100 , n27101 );
xor ( n27104 , n27011 , n27032 );
and ( n27105 , n18119 , n18410 );
and ( n27106 , n27104 , n27105 );
xor ( n27107 , n27104 , n27105 );
xor ( n27108 , n27015 , n27030 );
and ( n27109 , n18120 , n18410 );
and ( n27110 , n27108 , n27109 );
xor ( n27111 , n27108 , n27109 );
xor ( n27112 , n27019 , n27028 );
and ( n27113 , n18121 , n18410 );
and ( n27114 , n27112 , n27113 );
xor ( n27115 , n27112 , n27113 );
xor ( n27116 , n27023 , n27026 );
and ( n27117 , n18122 , n18410 );
and ( n27118 , n27116 , n27117 );
and ( n27119 , n27115 , n27118 );
or ( n27120 , n27114 , n27119 );
and ( n27121 , n27111 , n27120 );
or ( n27122 , n27110 , n27121 );
and ( n27123 , n27107 , n27122 );
or ( n27124 , n27106 , n27123 );
and ( n27125 , n27103 , n27124 );
or ( n27126 , n27102 , n27125 );
and ( n27127 , n27099 , n27126 );
or ( n27128 , n27098 , n27127 );
and ( n27129 , n27095 , n27128 );
or ( n27130 , n27094 , n27129 );
and ( n27131 , n27091 , n27130 );
or ( n27132 , n27090 , n27131 );
and ( n27133 , n27087 , n27132 );
or ( n27134 , n27086 , n27133 );
and ( n27135 , n27083 , n27134 );
or ( n27136 , n27082 , n27135 );
and ( n27137 , n27079 , n27136 );
or ( n27138 , n27078 , n27137 );
and ( n27139 , n27075 , n27138 );
or ( n27140 , n27074 , n27139 );
and ( n27141 , n27071 , n27140 );
or ( n27142 , n27070 , n27141 );
and ( n27143 , n27067 , n27142 );
or ( n27144 , n27066 , n27143 );
and ( n27145 , n27063 , n27144 );
or ( n27146 , n27062 , n27145 );
and ( n27147 , n27059 , n27146 );
or ( n27148 , n27058 , n27147 );
and ( n27149 , n18107 , n18408 );
and ( n27150 , n27148 , n27149 );
xor ( n27151 , n27148 , n27149 );
xor ( n27152 , n27059 , n27146 );
and ( n27153 , n18108 , n18408 );
and ( n27154 , n27152 , n27153 );
xor ( n27155 , n27152 , n27153 );
xor ( n27156 , n27063 , n27144 );
and ( n27157 , n18109 , n18408 );
and ( n27158 , n27156 , n27157 );
xor ( n27159 , n27156 , n27157 );
xor ( n27160 , n27067 , n27142 );
and ( n27161 , n18110 , n18408 );
and ( n27162 , n27160 , n27161 );
xor ( n27163 , n27160 , n27161 );
xor ( n27164 , n27071 , n27140 );
and ( n27165 , n18111 , n18408 );
and ( n27166 , n27164 , n27165 );
xor ( n27167 , n27164 , n27165 );
xor ( n27168 , n27075 , n27138 );
and ( n27169 , n18112 , n18408 );
and ( n27170 , n27168 , n27169 );
xor ( n27171 , n27168 , n27169 );
xor ( n27172 , n27079 , n27136 );
and ( n27173 , n18113 , n18408 );
and ( n27174 , n27172 , n27173 );
xor ( n27175 , n27172 , n27173 );
xor ( n27176 , n27083 , n27134 );
and ( n27177 , n18114 , n18408 );
and ( n27178 , n27176 , n27177 );
xor ( n27179 , n27176 , n27177 );
xor ( n27180 , n27087 , n27132 );
and ( n27181 , n18115 , n18408 );
and ( n27182 , n27180 , n27181 );
xor ( n27183 , n27180 , n27181 );
xor ( n27184 , n27091 , n27130 );
and ( n27185 , n18116 , n18408 );
and ( n27186 , n27184 , n27185 );
xor ( n27187 , n27184 , n27185 );
xor ( n27188 , n27095 , n27128 );
and ( n27189 , n18117 , n18408 );
and ( n27190 , n27188 , n27189 );
xor ( n27191 , n27188 , n27189 );
xor ( n27192 , n27099 , n27126 );
and ( n27193 , n18118 , n18408 );
and ( n27194 , n27192 , n27193 );
xor ( n27195 , n27192 , n27193 );
xor ( n27196 , n27103 , n27124 );
and ( n27197 , n18119 , n18408 );
and ( n27198 , n27196 , n27197 );
xor ( n27199 , n27196 , n27197 );
xor ( n27200 , n27107 , n27122 );
and ( n27201 , n18120 , n18408 );
and ( n27202 , n27200 , n27201 );
xor ( n27203 , n27200 , n27201 );
xor ( n27204 , n27111 , n27120 );
and ( n27205 , n18121 , n18408 );
and ( n27206 , n27204 , n27205 );
xor ( n27207 , n27204 , n27205 );
xor ( n27208 , n27115 , n27118 );
and ( n27209 , n18122 , n18408 );
and ( n27210 , n27208 , n27209 );
and ( n27211 , n27207 , n27210 );
or ( n27212 , n27206 , n27211 );
and ( n27213 , n27203 , n27212 );
or ( n27214 , n27202 , n27213 );
and ( n27215 , n27199 , n27214 );
or ( n27216 , n27198 , n27215 );
and ( n27217 , n27195 , n27216 );
or ( n27218 , n27194 , n27217 );
and ( n27219 , n27191 , n27218 );
or ( n27220 , n27190 , n27219 );
and ( n27221 , n27187 , n27220 );
or ( n27222 , n27186 , n27221 );
and ( n27223 , n27183 , n27222 );
or ( n27224 , n27182 , n27223 );
and ( n27225 , n27179 , n27224 );
or ( n27226 , n27178 , n27225 );
and ( n27227 , n27175 , n27226 );
or ( n27228 , n27174 , n27227 );
and ( n27229 , n27171 , n27228 );
or ( n27230 , n27170 , n27229 );
and ( n27231 , n27167 , n27230 );
or ( n27232 , n27166 , n27231 );
and ( n27233 , n27163 , n27232 );
or ( n27234 , n27162 , n27233 );
and ( n27235 , n27159 , n27234 );
or ( n27236 , n27158 , n27235 );
and ( n27237 , n27155 , n27236 );
or ( n27238 , n27154 , n27237 );
and ( n27239 , n27151 , n27238 );
or ( n27240 , n27150 , n27239 );
and ( n27241 , n18107 , n18406 );
and ( n27242 , n27240 , n27241 );
xor ( n27243 , n27240 , n27241 );
xor ( n27244 , n27151 , n27238 );
and ( n27245 , n18108 , n18406 );
and ( n27246 , n27244 , n27245 );
xor ( n27247 , n27244 , n27245 );
xor ( n27248 , n27155 , n27236 );
and ( n27249 , n18109 , n18406 );
and ( n27250 , n27248 , n27249 );
xor ( n27251 , n27248 , n27249 );
xor ( n27252 , n27159 , n27234 );
and ( n27253 , n18110 , n18406 );
and ( n27254 , n27252 , n27253 );
xor ( n27255 , n27252 , n27253 );
xor ( n27256 , n27163 , n27232 );
and ( n27257 , n18111 , n18406 );
and ( n27258 , n27256 , n27257 );
xor ( n27259 , n27256 , n27257 );
xor ( n27260 , n27167 , n27230 );
and ( n27261 , n18112 , n18406 );
and ( n27262 , n27260 , n27261 );
xor ( n27263 , n27260 , n27261 );
xor ( n27264 , n27171 , n27228 );
and ( n27265 , n18113 , n18406 );
and ( n27266 , n27264 , n27265 );
xor ( n27267 , n27264 , n27265 );
xor ( n27268 , n27175 , n27226 );
and ( n27269 , n18114 , n18406 );
and ( n27270 , n27268 , n27269 );
xor ( n27271 , n27268 , n27269 );
xor ( n27272 , n27179 , n27224 );
and ( n27273 , n18115 , n18406 );
and ( n27274 , n27272 , n27273 );
xor ( n27275 , n27272 , n27273 );
xor ( n27276 , n27183 , n27222 );
and ( n27277 , n18116 , n18406 );
and ( n27278 , n27276 , n27277 );
xor ( n27279 , n27276 , n27277 );
xor ( n27280 , n27187 , n27220 );
and ( n27281 , n18117 , n18406 );
and ( n27282 , n27280 , n27281 );
xor ( n27283 , n27280 , n27281 );
xor ( n27284 , n27191 , n27218 );
and ( n27285 , n18118 , n18406 );
and ( n27286 , n27284 , n27285 );
xor ( n27287 , n27284 , n27285 );
xor ( n27288 , n27195 , n27216 );
and ( n27289 , n18119 , n18406 );
and ( n27290 , n27288 , n27289 );
xor ( n27291 , n27288 , n27289 );
xor ( n27292 , n27199 , n27214 );
and ( n27293 , n18120 , n18406 );
and ( n27294 , n27292 , n27293 );
xor ( n27295 , n27292 , n27293 );
xor ( n27296 , n27203 , n27212 );
and ( n27297 , n18121 , n18406 );
and ( n27298 , n27296 , n27297 );
xor ( n27299 , n27296 , n27297 );
xor ( n27300 , n27207 , n27210 );
and ( n27301 , n18122 , n18406 );
and ( n27302 , n27300 , n27301 );
and ( n27303 , n27299 , n27302 );
or ( n27304 , n27298 , n27303 );
and ( n27305 , n27295 , n27304 );
or ( n27306 , n27294 , n27305 );
and ( n27307 , n27291 , n27306 );
or ( n27308 , n27290 , n27307 );
and ( n27309 , n27287 , n27308 );
or ( n27310 , n27286 , n27309 );
and ( n27311 , n27283 , n27310 );
or ( n27312 , n27282 , n27311 );
and ( n27313 , n27279 , n27312 );
or ( n27314 , n27278 , n27313 );
and ( n27315 , n27275 , n27314 );
or ( n27316 , n27274 , n27315 );
and ( n27317 , n27271 , n27316 );
or ( n27318 , n27270 , n27317 );
and ( n27319 , n27267 , n27318 );
or ( n27320 , n27266 , n27319 );
and ( n27321 , n27263 , n27320 );
or ( n27322 , n27262 , n27321 );
and ( n27323 , n27259 , n27322 );
or ( n27324 , n27258 , n27323 );
and ( n27325 , n27255 , n27324 );
or ( n27326 , n27254 , n27325 );
and ( n27327 , n27251 , n27326 );
or ( n27328 , n27250 , n27327 );
and ( n27329 , n27247 , n27328 );
or ( n27330 , n27246 , n27329 );
and ( n27331 , n27243 , n27330 );
or ( n27332 , n27242 , n27331 );
and ( n27333 , n18107 , n18404 );
and ( n27334 , n27332 , n27333 );
xor ( n27335 , n27332 , n27333 );
xor ( n27336 , n27243 , n27330 );
and ( n27337 , n18108 , n18404 );
and ( n27338 , n27336 , n27337 );
xor ( n27339 , n27336 , n27337 );
xor ( n27340 , n27247 , n27328 );
and ( n27341 , n18109 , n18404 );
and ( n27342 , n27340 , n27341 );
xor ( n27343 , n27340 , n27341 );
xor ( n27344 , n27251 , n27326 );
and ( n27345 , n18110 , n18404 );
and ( n27346 , n27344 , n27345 );
xor ( n27347 , n27344 , n27345 );
xor ( n27348 , n27255 , n27324 );
and ( n27349 , n18111 , n18404 );
and ( n27350 , n27348 , n27349 );
xor ( n27351 , n27348 , n27349 );
xor ( n27352 , n27259 , n27322 );
and ( n27353 , n18112 , n18404 );
and ( n27354 , n27352 , n27353 );
xor ( n27355 , n27352 , n27353 );
xor ( n27356 , n27263 , n27320 );
and ( n27357 , n18113 , n18404 );
and ( n27358 , n27356 , n27357 );
xor ( n27359 , n27356 , n27357 );
xor ( n27360 , n27267 , n27318 );
and ( n27361 , n18114 , n18404 );
and ( n27362 , n27360 , n27361 );
xor ( n27363 , n27360 , n27361 );
xor ( n27364 , n27271 , n27316 );
and ( n27365 , n18115 , n18404 );
and ( n27366 , n27364 , n27365 );
xor ( n27367 , n27364 , n27365 );
xor ( n27368 , n27275 , n27314 );
and ( n27369 , n18116 , n18404 );
and ( n27370 , n27368 , n27369 );
xor ( n27371 , n27368 , n27369 );
xor ( n27372 , n27279 , n27312 );
and ( n27373 , n18117 , n18404 );
and ( n27374 , n27372 , n27373 );
xor ( n27375 , n27372 , n27373 );
xor ( n27376 , n27283 , n27310 );
and ( n27377 , n18118 , n18404 );
and ( n27378 , n27376 , n27377 );
xor ( n27379 , n27376 , n27377 );
xor ( n27380 , n27287 , n27308 );
and ( n27381 , n18119 , n18404 );
and ( n27382 , n27380 , n27381 );
xor ( n27383 , n27380 , n27381 );
xor ( n27384 , n27291 , n27306 );
and ( n27385 , n18120 , n18404 );
and ( n27386 , n27384 , n27385 );
xor ( n27387 , n27384 , n27385 );
xor ( n27388 , n27295 , n27304 );
and ( n27389 , n18121 , n18404 );
and ( n27390 , n27388 , n27389 );
xor ( n27391 , n27388 , n27389 );
xor ( n27392 , n27299 , n27302 );
and ( n27393 , n18122 , n18404 );
and ( n27394 , n27392 , n27393 );
and ( n27395 , n27391 , n27394 );
or ( n27396 , n27390 , n27395 );
and ( n27397 , n27387 , n27396 );
or ( n27398 , n27386 , n27397 );
and ( n27399 , n27383 , n27398 );
or ( n27400 , n27382 , n27399 );
and ( n27401 , n27379 , n27400 );
or ( n27402 , n27378 , n27401 );
and ( n27403 , n27375 , n27402 );
or ( n27404 , n27374 , n27403 );
and ( n27405 , n27371 , n27404 );
or ( n27406 , n27370 , n27405 );
and ( n27407 , n27367 , n27406 );
or ( n27408 , n27366 , n27407 );
and ( n27409 , n27363 , n27408 );
or ( n27410 , n27362 , n27409 );
and ( n27411 , n27359 , n27410 );
or ( n27412 , n27358 , n27411 );
and ( n27413 , n27355 , n27412 );
or ( n27414 , n27354 , n27413 );
and ( n27415 , n27351 , n27414 );
or ( n27416 , n27350 , n27415 );
and ( n27417 , n27347 , n27416 );
or ( n27418 , n27346 , n27417 );
and ( n27419 , n27343 , n27418 );
or ( n27420 , n27342 , n27419 );
and ( n27421 , n27339 , n27420 );
or ( n27422 , n27338 , n27421 );
and ( n27423 , n27335 , n27422 );
or ( n27424 , n27334 , n27423 );
and ( n27425 , n18107 , n18402 );
and ( n27426 , n27424 , n27425 );
xor ( n27427 , n27424 , n27425 );
xor ( n27428 , n27335 , n27422 );
and ( n27429 , n18108 , n18402 );
and ( n27430 , n27428 , n27429 );
xor ( n27431 , n27428 , n27429 );
xor ( n27432 , n27339 , n27420 );
and ( n27433 , n18109 , n18402 );
and ( n27434 , n27432 , n27433 );
xor ( n27435 , n27432 , n27433 );
xor ( n27436 , n27343 , n27418 );
and ( n27437 , n18110 , n18402 );
and ( n27438 , n27436 , n27437 );
xor ( n27439 , n27436 , n27437 );
xor ( n27440 , n27347 , n27416 );
and ( n27441 , n18111 , n18402 );
and ( n27442 , n27440 , n27441 );
xor ( n27443 , n27440 , n27441 );
xor ( n27444 , n27351 , n27414 );
and ( n27445 , n18112 , n18402 );
and ( n27446 , n27444 , n27445 );
xor ( n27447 , n27444 , n27445 );
xor ( n27448 , n27355 , n27412 );
and ( n27449 , n18113 , n18402 );
and ( n27450 , n27448 , n27449 );
xor ( n27451 , n27448 , n27449 );
xor ( n27452 , n27359 , n27410 );
and ( n27453 , n18114 , n18402 );
and ( n27454 , n27452 , n27453 );
xor ( n27455 , n27452 , n27453 );
xor ( n27456 , n27363 , n27408 );
and ( n27457 , n18115 , n18402 );
and ( n27458 , n27456 , n27457 );
xor ( n27459 , n27456 , n27457 );
xor ( n27460 , n27367 , n27406 );
and ( n27461 , n18116 , n18402 );
and ( n27462 , n27460 , n27461 );
xor ( n27463 , n27460 , n27461 );
xor ( n27464 , n27371 , n27404 );
and ( n27465 , n18117 , n18402 );
and ( n27466 , n27464 , n27465 );
xor ( n27467 , n27464 , n27465 );
xor ( n27468 , n27375 , n27402 );
and ( n27469 , n18118 , n18402 );
and ( n27470 , n27468 , n27469 );
xor ( n27471 , n27468 , n27469 );
xor ( n27472 , n27379 , n27400 );
and ( n27473 , n18119 , n18402 );
and ( n27474 , n27472 , n27473 );
xor ( n27475 , n27472 , n27473 );
xor ( n27476 , n27383 , n27398 );
and ( n27477 , n18120 , n18402 );
and ( n27478 , n27476 , n27477 );
xor ( n27479 , n27476 , n27477 );
xor ( n27480 , n27387 , n27396 );
and ( n27481 , n18121 , n18402 );
and ( n27482 , n27480 , n27481 );
xor ( n27483 , n27480 , n27481 );
xor ( n27484 , n27391 , n27394 );
and ( n27485 , n18122 , n18402 );
and ( n27486 , n27484 , n27485 );
and ( n27487 , n27483 , n27486 );
or ( n27488 , n27482 , n27487 );
and ( n27489 , n27479 , n27488 );
or ( n27490 , n27478 , n27489 );
and ( n27491 , n27475 , n27490 );
or ( n27492 , n27474 , n27491 );
and ( n27493 , n27471 , n27492 );
or ( n27494 , n27470 , n27493 );
and ( n27495 , n27467 , n27494 );
or ( n27496 , n27466 , n27495 );
and ( n27497 , n27463 , n27496 );
or ( n27498 , n27462 , n27497 );
and ( n27499 , n27459 , n27498 );
or ( n27500 , n27458 , n27499 );
and ( n27501 , n27455 , n27500 );
or ( n27502 , n27454 , n27501 );
and ( n27503 , n27451 , n27502 );
or ( n27504 , n27450 , n27503 );
and ( n27505 , n27447 , n27504 );
or ( n27506 , n27446 , n27505 );
and ( n27507 , n27443 , n27506 );
or ( n27508 , n27442 , n27507 );
and ( n27509 , n27439 , n27508 );
or ( n27510 , n27438 , n27509 );
and ( n27511 , n27435 , n27510 );
or ( n27512 , n27434 , n27511 );
and ( n27513 , n27431 , n27512 );
or ( n27514 , n27430 , n27513 );
and ( n27515 , n27427 , n27514 );
or ( n27516 , n27426 , n27515 );
and ( n27517 , n18107 , n18400 );
and ( n27518 , n27516 , n27517 );
xor ( n27519 , n27516 , n27517 );
xor ( n27520 , n27427 , n27514 );
and ( n27521 , n18108 , n18400 );
and ( n27522 , n27520 , n27521 );
xor ( n27523 , n27520 , n27521 );
xor ( n27524 , n27431 , n27512 );
and ( n27525 , n18109 , n18400 );
and ( n27526 , n27524 , n27525 );
xor ( n27527 , n27524 , n27525 );
xor ( n27528 , n27435 , n27510 );
and ( n27529 , n18110 , n18400 );
and ( n27530 , n27528 , n27529 );
xor ( n27531 , n27528 , n27529 );
xor ( n27532 , n27439 , n27508 );
and ( n27533 , n18111 , n18400 );
and ( n27534 , n27532 , n27533 );
xor ( n27535 , n27532 , n27533 );
xor ( n27536 , n27443 , n27506 );
and ( n27537 , n18112 , n18400 );
and ( n27538 , n27536 , n27537 );
xor ( n27539 , n27536 , n27537 );
xor ( n27540 , n27447 , n27504 );
and ( n27541 , n18113 , n18400 );
and ( n27542 , n27540 , n27541 );
xor ( n27543 , n27540 , n27541 );
xor ( n27544 , n27451 , n27502 );
and ( n27545 , n18114 , n18400 );
and ( n27546 , n27544 , n27545 );
xor ( n27547 , n27544 , n27545 );
xor ( n27548 , n27455 , n27500 );
and ( n27549 , n18115 , n18400 );
and ( n27550 , n27548 , n27549 );
xor ( n27551 , n27548 , n27549 );
xor ( n27552 , n27459 , n27498 );
and ( n27553 , n18116 , n18400 );
and ( n27554 , n27552 , n27553 );
xor ( n27555 , n27552 , n27553 );
xor ( n27556 , n27463 , n27496 );
and ( n27557 , n18117 , n18400 );
and ( n27558 , n27556 , n27557 );
xor ( n27559 , n27556 , n27557 );
xor ( n27560 , n27467 , n27494 );
and ( n27561 , n18118 , n18400 );
and ( n27562 , n27560 , n27561 );
xor ( n27563 , n27560 , n27561 );
xor ( n27564 , n27471 , n27492 );
and ( n27565 , n18119 , n18400 );
and ( n27566 , n27564 , n27565 );
xor ( n27567 , n27564 , n27565 );
xor ( n27568 , n27475 , n27490 );
and ( n27569 , n18120 , n18400 );
and ( n27570 , n27568 , n27569 );
xor ( n27571 , n27568 , n27569 );
xor ( n27572 , n27479 , n27488 );
and ( n27573 , n18121 , n18400 );
and ( n27574 , n27572 , n27573 );
xor ( n27575 , n27572 , n27573 );
xor ( n27576 , n27483 , n27486 );
and ( n27577 , n18122 , n18400 );
and ( n27578 , n27576 , n27577 );
and ( n27579 , n27575 , n27578 );
or ( n27580 , n27574 , n27579 );
and ( n27581 , n27571 , n27580 );
or ( n27582 , n27570 , n27581 );
and ( n27583 , n27567 , n27582 );
or ( n27584 , n27566 , n27583 );
and ( n27585 , n27563 , n27584 );
or ( n27586 , n27562 , n27585 );
and ( n27587 , n27559 , n27586 );
or ( n27588 , n27558 , n27587 );
and ( n27589 , n27555 , n27588 );
or ( n27590 , n27554 , n27589 );
and ( n27591 , n27551 , n27590 );
or ( n27592 , n27550 , n27591 );
and ( n27593 , n27547 , n27592 );
or ( n27594 , n27546 , n27593 );
and ( n27595 , n27543 , n27594 );
or ( n27596 , n27542 , n27595 );
and ( n27597 , n27539 , n27596 );
or ( n27598 , n27538 , n27597 );
and ( n27599 , n27535 , n27598 );
or ( n27600 , n27534 , n27599 );
and ( n27601 , n27531 , n27600 );
or ( n27602 , n27530 , n27601 );
and ( n27603 , n27527 , n27602 );
or ( n27604 , n27526 , n27603 );
and ( n27605 , n27523 , n27604 );
or ( n27606 , n27522 , n27605 );
and ( n27607 , n27519 , n27606 );
or ( n27608 , n27518 , n27607 );
and ( n27609 , n18107 , n18398 );
and ( n27610 , n27608 , n27609 );
xor ( n27611 , n27608 , n27609 );
xor ( n27612 , n27519 , n27606 );
and ( n27613 , n18108 , n18398 );
and ( n27614 , n27612 , n27613 );
xor ( n27615 , n27612 , n27613 );
xor ( n27616 , n27523 , n27604 );
and ( n27617 , n18109 , n18398 );
and ( n27618 , n27616 , n27617 );
xor ( n27619 , n27616 , n27617 );
xor ( n27620 , n27527 , n27602 );
and ( n27621 , n18110 , n18398 );
and ( n27622 , n27620 , n27621 );
xor ( n27623 , n27620 , n27621 );
xor ( n27624 , n27531 , n27600 );
and ( n27625 , n18111 , n18398 );
and ( n27626 , n27624 , n27625 );
xor ( n27627 , n27624 , n27625 );
xor ( n27628 , n27535 , n27598 );
and ( n27629 , n18112 , n18398 );
and ( n27630 , n27628 , n27629 );
xor ( n27631 , n27628 , n27629 );
xor ( n27632 , n27539 , n27596 );
and ( n27633 , n18113 , n18398 );
and ( n27634 , n27632 , n27633 );
xor ( n27635 , n27632 , n27633 );
xor ( n27636 , n27543 , n27594 );
and ( n27637 , n18114 , n18398 );
and ( n27638 , n27636 , n27637 );
xor ( n27639 , n27636 , n27637 );
xor ( n27640 , n27547 , n27592 );
and ( n27641 , n18115 , n18398 );
and ( n27642 , n27640 , n27641 );
xor ( n27643 , n27640 , n27641 );
xor ( n27644 , n27551 , n27590 );
and ( n27645 , n18116 , n18398 );
and ( n27646 , n27644 , n27645 );
xor ( n27647 , n27644 , n27645 );
xor ( n27648 , n27555 , n27588 );
and ( n27649 , n18117 , n18398 );
and ( n27650 , n27648 , n27649 );
xor ( n27651 , n27648 , n27649 );
xor ( n27652 , n27559 , n27586 );
and ( n27653 , n18118 , n18398 );
and ( n27654 , n27652 , n27653 );
xor ( n27655 , n27652 , n27653 );
xor ( n27656 , n27563 , n27584 );
and ( n27657 , n18119 , n18398 );
and ( n27658 , n27656 , n27657 );
xor ( n27659 , n27656 , n27657 );
xor ( n27660 , n27567 , n27582 );
and ( n27661 , n18120 , n18398 );
and ( n27662 , n27660 , n27661 );
xor ( n27663 , n27660 , n27661 );
xor ( n27664 , n27571 , n27580 );
and ( n27665 , n18121 , n18398 );
and ( n27666 , n27664 , n27665 );
xor ( n27667 , n27664 , n27665 );
xor ( n27668 , n27575 , n27578 );
and ( n27669 , n18122 , n18398 );
and ( n27670 , n27668 , n27669 );
and ( n27671 , n27667 , n27670 );
or ( n27672 , n27666 , n27671 );
and ( n27673 , n27663 , n27672 );
or ( n27674 , n27662 , n27673 );
and ( n27675 , n27659 , n27674 );
or ( n27676 , n27658 , n27675 );
and ( n27677 , n27655 , n27676 );
or ( n27678 , n27654 , n27677 );
and ( n27679 , n27651 , n27678 );
or ( n27680 , n27650 , n27679 );
and ( n27681 , n27647 , n27680 );
or ( n27682 , n27646 , n27681 );
and ( n27683 , n27643 , n27682 );
or ( n27684 , n27642 , n27683 );
and ( n27685 , n27639 , n27684 );
or ( n27686 , n27638 , n27685 );
and ( n27687 , n27635 , n27686 );
or ( n27688 , n27634 , n27687 );
and ( n27689 , n27631 , n27688 );
or ( n27690 , n27630 , n27689 );
and ( n27691 , n27627 , n27690 );
or ( n27692 , n27626 , n27691 );
and ( n27693 , n27623 , n27692 );
or ( n27694 , n27622 , n27693 );
and ( n27695 , n27619 , n27694 );
or ( n27696 , n27618 , n27695 );
and ( n27697 , n27615 , n27696 );
or ( n27698 , n27614 , n27697 );
and ( n27699 , n27611 , n27698 );
or ( n27700 , n27610 , n27699 );
and ( n27701 , n18107 , n18396 );
and ( n27702 , n27700 , n27701 );
xor ( n27703 , n27700 , n27701 );
xor ( n27704 , n27611 , n27698 );
and ( n27705 , n18108 , n18396 );
and ( n27706 , n27704 , n27705 );
xor ( n27707 , n27704 , n27705 );
xor ( n27708 , n27615 , n27696 );
and ( n27709 , n18109 , n18396 );
and ( n27710 , n27708 , n27709 );
xor ( n27711 , n27708 , n27709 );
xor ( n27712 , n27619 , n27694 );
and ( n27713 , n18110 , n18396 );
and ( n27714 , n27712 , n27713 );
xor ( n27715 , n27712 , n27713 );
xor ( n27716 , n27623 , n27692 );
and ( n27717 , n18111 , n18396 );
and ( n27718 , n27716 , n27717 );
xor ( n27719 , n27716 , n27717 );
xor ( n27720 , n27627 , n27690 );
and ( n27721 , n18112 , n18396 );
and ( n27722 , n27720 , n27721 );
xor ( n27723 , n27720 , n27721 );
xor ( n27724 , n27631 , n27688 );
and ( n27725 , n18113 , n18396 );
and ( n27726 , n27724 , n27725 );
xor ( n27727 , n27724 , n27725 );
xor ( n27728 , n27635 , n27686 );
and ( n27729 , n18114 , n18396 );
and ( n27730 , n27728 , n27729 );
xor ( n27731 , n27728 , n27729 );
xor ( n27732 , n27639 , n27684 );
and ( n27733 , n18115 , n18396 );
and ( n27734 , n27732 , n27733 );
xor ( n27735 , n27732 , n27733 );
xor ( n27736 , n27643 , n27682 );
and ( n27737 , n18116 , n18396 );
and ( n27738 , n27736 , n27737 );
xor ( n27739 , n27736 , n27737 );
xor ( n27740 , n27647 , n27680 );
and ( n27741 , n18117 , n18396 );
and ( n27742 , n27740 , n27741 );
xor ( n27743 , n27740 , n27741 );
xor ( n27744 , n27651 , n27678 );
and ( n27745 , n18118 , n18396 );
and ( n27746 , n27744 , n27745 );
xor ( n27747 , n27744 , n27745 );
xor ( n27748 , n27655 , n27676 );
and ( n27749 , n18119 , n18396 );
and ( n27750 , n27748 , n27749 );
xor ( n27751 , n27748 , n27749 );
xor ( n27752 , n27659 , n27674 );
and ( n27753 , n18120 , n18396 );
and ( n27754 , n27752 , n27753 );
xor ( n27755 , n27752 , n27753 );
xor ( n27756 , n27663 , n27672 );
and ( n27757 , n18121 , n18396 );
and ( n27758 , n27756 , n27757 );
xor ( n27759 , n27756 , n27757 );
xor ( n27760 , n27667 , n27670 );
and ( n27761 , n18122 , n18396 );
and ( n27762 , n27760 , n27761 );
and ( n27763 , n27759 , n27762 );
or ( n27764 , n27758 , n27763 );
and ( n27765 , n27755 , n27764 );
or ( n27766 , n27754 , n27765 );
and ( n27767 , n27751 , n27766 );
or ( n27768 , n27750 , n27767 );
and ( n27769 , n27747 , n27768 );
or ( n27770 , n27746 , n27769 );
and ( n27771 , n27743 , n27770 );
or ( n27772 , n27742 , n27771 );
and ( n27773 , n27739 , n27772 );
or ( n27774 , n27738 , n27773 );
and ( n27775 , n27735 , n27774 );
or ( n27776 , n27734 , n27775 );
and ( n27777 , n27731 , n27776 );
or ( n27778 , n27730 , n27777 );
and ( n27779 , n27727 , n27778 );
or ( n27780 , n27726 , n27779 );
and ( n27781 , n27723 , n27780 );
or ( n27782 , n27722 , n27781 );
and ( n27783 , n27719 , n27782 );
or ( n27784 , n27718 , n27783 );
and ( n27785 , n27715 , n27784 );
or ( n27786 , n27714 , n27785 );
and ( n27787 , n27711 , n27786 );
or ( n27788 , n27710 , n27787 );
and ( n27789 , n27707 , n27788 );
or ( n27790 , n27706 , n27789 );
and ( n27791 , n27703 , n27790 );
or ( n27792 , n27702 , n27791 );
and ( n27793 , n18107 , n18394 );
and ( n27794 , n27792 , n27793 );
xor ( n27795 , n27792 , n27793 );
xor ( n27796 , n27703 , n27790 );
and ( n27797 , n18108 , n18394 );
and ( n27798 , n27796 , n27797 );
xor ( n27799 , n27796 , n27797 );
xor ( n27800 , n27707 , n27788 );
and ( n27801 , n18109 , n18394 );
and ( n27802 , n27800 , n27801 );
xor ( n27803 , n27800 , n27801 );
xor ( n27804 , n27711 , n27786 );
and ( n27805 , n18110 , n18394 );
and ( n27806 , n27804 , n27805 );
xor ( n27807 , n27804 , n27805 );
xor ( n27808 , n27715 , n27784 );
and ( n27809 , n18111 , n18394 );
and ( n27810 , n27808 , n27809 );
xor ( n27811 , n27808 , n27809 );
xor ( n27812 , n27719 , n27782 );
and ( n27813 , n18112 , n18394 );
and ( n27814 , n27812 , n27813 );
xor ( n27815 , n27812 , n27813 );
xor ( n27816 , n27723 , n27780 );
and ( n27817 , n18113 , n18394 );
and ( n27818 , n27816 , n27817 );
xor ( n27819 , n27816 , n27817 );
xor ( n27820 , n27727 , n27778 );
and ( n27821 , n18114 , n18394 );
and ( n27822 , n27820 , n27821 );
xor ( n27823 , n27820 , n27821 );
xor ( n27824 , n27731 , n27776 );
and ( n27825 , n18115 , n18394 );
and ( n27826 , n27824 , n27825 );
xor ( n27827 , n27824 , n27825 );
xor ( n27828 , n27735 , n27774 );
and ( n27829 , n18116 , n18394 );
and ( n27830 , n27828 , n27829 );
xor ( n27831 , n27828 , n27829 );
xor ( n27832 , n27739 , n27772 );
and ( n27833 , n18117 , n18394 );
and ( n27834 , n27832 , n27833 );
xor ( n27835 , n27832 , n27833 );
xor ( n27836 , n27743 , n27770 );
and ( n27837 , n18118 , n18394 );
and ( n27838 , n27836 , n27837 );
xor ( n27839 , n27836 , n27837 );
xor ( n27840 , n27747 , n27768 );
and ( n27841 , n18119 , n18394 );
and ( n27842 , n27840 , n27841 );
xor ( n27843 , n27840 , n27841 );
xor ( n27844 , n27751 , n27766 );
and ( n27845 , n18120 , n18394 );
and ( n27846 , n27844 , n27845 );
xor ( n27847 , n27844 , n27845 );
xor ( n27848 , n27755 , n27764 );
and ( n27849 , n18121 , n18394 );
and ( n27850 , n27848 , n27849 );
xor ( n27851 , n27848 , n27849 );
xor ( n27852 , n27759 , n27762 );
and ( n27853 , n18122 , n18394 );
and ( n27854 , n27852 , n27853 );
and ( n27855 , n27851 , n27854 );
or ( n27856 , n27850 , n27855 );
and ( n27857 , n27847 , n27856 );
or ( n27858 , n27846 , n27857 );
and ( n27859 , n27843 , n27858 );
or ( n27860 , n27842 , n27859 );
and ( n27861 , n27839 , n27860 );
or ( n27862 , n27838 , n27861 );
and ( n27863 , n27835 , n27862 );
or ( n27864 , n27834 , n27863 );
and ( n27865 , n27831 , n27864 );
or ( n27866 , n27830 , n27865 );
and ( n27867 , n27827 , n27866 );
or ( n27868 , n27826 , n27867 );
and ( n27869 , n27823 , n27868 );
or ( n27870 , n27822 , n27869 );
and ( n27871 , n27819 , n27870 );
or ( n27872 , n27818 , n27871 );
and ( n27873 , n27815 , n27872 );
or ( n27874 , n27814 , n27873 );
and ( n27875 , n27811 , n27874 );
or ( n27876 , n27810 , n27875 );
and ( n27877 , n27807 , n27876 );
or ( n27878 , n27806 , n27877 );
and ( n27879 , n27803 , n27878 );
or ( n27880 , n27802 , n27879 );
and ( n27881 , n27799 , n27880 );
or ( n27882 , n27798 , n27881 );
and ( n27883 , n27795 , n27882 );
or ( n27884 , n27794 , n27883 );
and ( n27885 , n18107 , n18392 );
and ( n27886 , n27884 , n27885 );
xor ( n27887 , n27884 , n27885 );
xor ( n27888 , n27795 , n27882 );
and ( n27889 , n18108 , n18392 );
and ( n27890 , n27888 , n27889 );
xor ( n27891 , n27888 , n27889 );
xor ( n27892 , n27799 , n27880 );
and ( n27893 , n18109 , n18392 );
and ( n27894 , n27892 , n27893 );
xor ( n27895 , n27892 , n27893 );
xor ( n27896 , n27803 , n27878 );
and ( n27897 , n18110 , n18392 );
and ( n27898 , n27896 , n27897 );
xor ( n27899 , n27896 , n27897 );
xor ( n27900 , n27807 , n27876 );
and ( n27901 , n18111 , n18392 );
and ( n27902 , n27900 , n27901 );
xor ( n27903 , n27900 , n27901 );
xor ( n27904 , n27811 , n27874 );
and ( n27905 , n18112 , n18392 );
and ( n27906 , n27904 , n27905 );
xor ( n27907 , n27904 , n27905 );
xor ( n27908 , n27815 , n27872 );
and ( n27909 , n18113 , n18392 );
and ( n27910 , n27908 , n27909 );
xor ( n27911 , n27908 , n27909 );
xor ( n27912 , n27819 , n27870 );
and ( n27913 , n18114 , n18392 );
and ( n27914 , n27912 , n27913 );
xor ( n27915 , n27912 , n27913 );
xor ( n27916 , n27823 , n27868 );
and ( n27917 , n18115 , n18392 );
and ( n27918 , n27916 , n27917 );
xor ( n27919 , n27916 , n27917 );
xor ( n27920 , n27827 , n27866 );
and ( n27921 , n18116 , n18392 );
and ( n27922 , n27920 , n27921 );
xor ( n27923 , n27920 , n27921 );
xor ( n27924 , n27831 , n27864 );
and ( n27925 , n18117 , n18392 );
and ( n27926 , n27924 , n27925 );
xor ( n27927 , n27924 , n27925 );
xor ( n27928 , n27835 , n27862 );
and ( n27929 , n18118 , n18392 );
and ( n27930 , n27928 , n27929 );
xor ( n27931 , n27928 , n27929 );
xor ( n27932 , n27839 , n27860 );
and ( n27933 , n18119 , n18392 );
and ( n27934 , n27932 , n27933 );
xor ( n27935 , n27932 , n27933 );
xor ( n27936 , n27843 , n27858 );
and ( n27937 , n18120 , n18392 );
and ( n27938 , n27936 , n27937 );
xor ( n27939 , n27936 , n27937 );
xor ( n27940 , n27847 , n27856 );
and ( n27941 , n18121 , n18392 );
and ( n27942 , n27940 , n27941 );
xor ( n27943 , n27940 , n27941 );
xor ( n27944 , n27851 , n27854 );
and ( n27945 , n18122 , n18392 );
and ( n27946 , n27944 , n27945 );
and ( n27947 , n27943 , n27946 );
or ( n27948 , n27942 , n27947 );
and ( n27949 , n27939 , n27948 );
or ( n27950 , n27938 , n27949 );
and ( n27951 , n27935 , n27950 );
or ( n27952 , n27934 , n27951 );
and ( n27953 , n27931 , n27952 );
or ( n27954 , n27930 , n27953 );
and ( n27955 , n27927 , n27954 );
or ( n27956 , n27926 , n27955 );
and ( n27957 , n27923 , n27956 );
or ( n27958 , n27922 , n27957 );
and ( n27959 , n27919 , n27958 );
or ( n27960 , n27918 , n27959 );
and ( n27961 , n27915 , n27960 );
or ( n27962 , n27914 , n27961 );
and ( n27963 , n27911 , n27962 );
or ( n27964 , n27910 , n27963 );
and ( n27965 , n27907 , n27964 );
or ( n27966 , n27906 , n27965 );
and ( n27967 , n27903 , n27966 );
or ( n27968 , n27902 , n27967 );
and ( n27969 , n27899 , n27968 );
or ( n27970 , n27898 , n27969 );
and ( n27971 , n27895 , n27970 );
or ( n27972 , n27894 , n27971 );
and ( n27973 , n27891 , n27972 );
or ( n27974 , n27890 , n27973 );
and ( n27975 , n27887 , n27974 );
or ( n27976 , n27886 , n27975 );
and ( n27977 , n18107 , n18390 );
and ( n27978 , n27976 , n27977 );
xor ( n27979 , n27976 , n27977 );
xor ( n27980 , n27887 , n27974 );
and ( n27981 , n18108 , n18390 );
and ( n27982 , n27980 , n27981 );
xor ( n27983 , n27980 , n27981 );
xor ( n27984 , n27891 , n27972 );
and ( n27985 , n18109 , n18390 );
and ( n27986 , n27984 , n27985 );
xor ( n27987 , n27984 , n27985 );
xor ( n27988 , n27895 , n27970 );
and ( n27989 , n18110 , n18390 );
and ( n27990 , n27988 , n27989 );
xor ( n27991 , n27988 , n27989 );
xor ( n27992 , n27899 , n27968 );
and ( n27993 , n18111 , n18390 );
and ( n27994 , n27992 , n27993 );
xor ( n27995 , n27992 , n27993 );
xor ( n27996 , n27903 , n27966 );
and ( n27997 , n18112 , n18390 );
and ( n27998 , n27996 , n27997 );
xor ( n27999 , n27996 , n27997 );
xor ( n28000 , n27907 , n27964 );
and ( n28001 , n18113 , n18390 );
and ( n28002 , n28000 , n28001 );
xor ( n28003 , n28000 , n28001 );
xor ( n28004 , n27911 , n27962 );
and ( n28005 , n18114 , n18390 );
and ( n28006 , n28004 , n28005 );
xor ( n28007 , n28004 , n28005 );
xor ( n28008 , n27915 , n27960 );
and ( n28009 , n18115 , n18390 );
and ( n28010 , n28008 , n28009 );
xor ( n28011 , n28008 , n28009 );
xor ( n28012 , n27919 , n27958 );
and ( n28013 , n18116 , n18390 );
and ( n28014 , n28012 , n28013 );
xor ( n28015 , n28012 , n28013 );
xor ( n28016 , n27923 , n27956 );
and ( n28017 , n18117 , n18390 );
and ( n28018 , n28016 , n28017 );
xor ( n28019 , n28016 , n28017 );
xor ( n28020 , n27927 , n27954 );
and ( n28021 , n18118 , n18390 );
and ( n28022 , n28020 , n28021 );
xor ( n28023 , n28020 , n28021 );
xor ( n28024 , n27931 , n27952 );
and ( n28025 , n18119 , n18390 );
and ( n28026 , n28024 , n28025 );
xor ( n28027 , n28024 , n28025 );
xor ( n28028 , n27935 , n27950 );
and ( n28029 , n18120 , n18390 );
and ( n28030 , n28028 , n28029 );
xor ( n28031 , n28028 , n28029 );
xor ( n28032 , n27939 , n27948 );
and ( n28033 , n18121 , n18390 );
and ( n28034 , n28032 , n28033 );
xor ( n28035 , n28032 , n28033 );
xor ( n28036 , n27943 , n27946 );
and ( n28037 , n18122 , n18390 );
and ( n28038 , n28036 , n28037 );
and ( n28039 , n28035 , n28038 );
or ( n28040 , n28034 , n28039 );
and ( n28041 , n28031 , n28040 );
or ( n28042 , n28030 , n28041 );
and ( n28043 , n28027 , n28042 );
or ( n28044 , n28026 , n28043 );
and ( n28045 , n28023 , n28044 );
or ( n28046 , n28022 , n28045 );
and ( n28047 , n28019 , n28046 );
or ( n28048 , n28018 , n28047 );
and ( n28049 , n28015 , n28048 );
or ( n28050 , n28014 , n28049 );
and ( n28051 , n28011 , n28050 );
or ( n28052 , n28010 , n28051 );
and ( n28053 , n28007 , n28052 );
or ( n28054 , n28006 , n28053 );
and ( n28055 , n28003 , n28054 );
or ( n28056 , n28002 , n28055 );
and ( n28057 , n27999 , n28056 );
or ( n28058 , n27998 , n28057 );
and ( n28059 , n27995 , n28058 );
or ( n28060 , n27994 , n28059 );
and ( n28061 , n27991 , n28060 );
or ( n28062 , n27990 , n28061 );
and ( n28063 , n27987 , n28062 );
or ( n28064 , n27986 , n28063 );
and ( n28065 , n27983 , n28064 );
or ( n28066 , n27982 , n28065 );
and ( n28067 , n27979 , n28066 );
or ( n28068 , n27978 , n28067 );
and ( n28069 , n18107 , n18388 );
and ( n28070 , n28068 , n28069 );
xor ( n28071 , n28068 , n28069 );
xor ( n28072 , n27979 , n28066 );
and ( n28073 , n18108 , n18388 );
and ( n28074 , n28072 , n28073 );
xor ( n28075 , n28072 , n28073 );
xor ( n28076 , n27983 , n28064 );
and ( n28077 , n18109 , n18388 );
and ( n28078 , n28076 , n28077 );
xor ( n28079 , n28076 , n28077 );
xor ( n28080 , n27987 , n28062 );
and ( n28081 , n18110 , n18388 );
and ( n28082 , n28080 , n28081 );
xor ( n28083 , n28080 , n28081 );
xor ( n28084 , n27991 , n28060 );
and ( n28085 , n18111 , n18388 );
and ( n28086 , n28084 , n28085 );
xor ( n28087 , n28084 , n28085 );
xor ( n28088 , n27995 , n28058 );
and ( n28089 , n18112 , n18388 );
and ( n28090 , n28088 , n28089 );
xor ( n28091 , n28088 , n28089 );
xor ( n28092 , n27999 , n28056 );
and ( n28093 , n18113 , n18388 );
and ( n28094 , n28092 , n28093 );
xor ( n28095 , n28092 , n28093 );
xor ( n28096 , n28003 , n28054 );
and ( n28097 , n18114 , n18388 );
and ( n28098 , n28096 , n28097 );
xor ( n28099 , n28096 , n28097 );
xor ( n28100 , n28007 , n28052 );
and ( n28101 , n18115 , n18388 );
and ( n28102 , n28100 , n28101 );
xor ( n28103 , n28100 , n28101 );
xor ( n28104 , n28011 , n28050 );
and ( n28105 , n18116 , n18388 );
and ( n28106 , n28104 , n28105 );
xor ( n28107 , n28104 , n28105 );
xor ( n28108 , n28015 , n28048 );
and ( n28109 , n18117 , n18388 );
and ( n28110 , n28108 , n28109 );
xor ( n28111 , n28108 , n28109 );
xor ( n28112 , n28019 , n28046 );
and ( n28113 , n18118 , n18388 );
and ( n28114 , n28112 , n28113 );
xor ( n28115 , n28112 , n28113 );
xor ( n28116 , n28023 , n28044 );
and ( n28117 , n18119 , n18388 );
and ( n28118 , n28116 , n28117 );
xor ( n28119 , n28116 , n28117 );
xor ( n28120 , n28027 , n28042 );
and ( n28121 , n18120 , n18388 );
and ( n28122 , n28120 , n28121 );
xor ( n28123 , n28120 , n28121 );
xor ( n28124 , n28031 , n28040 );
and ( n28125 , n18121 , n18388 );
and ( n28126 , n28124 , n28125 );
xor ( n28127 , n28124 , n28125 );
xor ( n28128 , n28035 , n28038 );
and ( n28129 , n18122 , n18388 );
and ( n28130 , n28128 , n28129 );
and ( n28131 , n28127 , n28130 );
or ( n28132 , n28126 , n28131 );
and ( n28133 , n28123 , n28132 );
or ( n28134 , n28122 , n28133 );
and ( n28135 , n28119 , n28134 );
or ( n28136 , n28118 , n28135 );
and ( n28137 , n28115 , n28136 );
or ( n28138 , n28114 , n28137 );
and ( n28139 , n28111 , n28138 );
or ( n28140 , n28110 , n28139 );
and ( n28141 , n28107 , n28140 );
or ( n28142 , n28106 , n28141 );
and ( n28143 , n28103 , n28142 );
or ( n28144 , n28102 , n28143 );
and ( n28145 , n28099 , n28144 );
or ( n28146 , n28098 , n28145 );
and ( n28147 , n28095 , n28146 );
or ( n28148 , n28094 , n28147 );
and ( n28149 , n28091 , n28148 );
or ( n28150 , n28090 , n28149 );
and ( n28151 , n28087 , n28150 );
or ( n28152 , n28086 , n28151 );
and ( n28153 , n28083 , n28152 );
or ( n28154 , n28082 , n28153 );
and ( n28155 , n28079 , n28154 );
or ( n28156 , n28078 , n28155 );
and ( n28157 , n28075 , n28156 );
or ( n28158 , n28074 , n28157 );
and ( n28159 , n28071 , n28158 );
or ( n28160 , n28070 , n28159 );
and ( n28161 , n18107 , n18386 );
and ( n28162 , n28160 , n28161 );
xor ( n28163 , n28160 , n28161 );
xor ( n28164 , n28071 , n28158 );
and ( n28165 , n18108 , n18386 );
and ( n28166 , n28164 , n28165 );
xor ( n28167 , n28164 , n28165 );
xor ( n28168 , n28075 , n28156 );
and ( n28169 , n18109 , n18386 );
and ( n28170 , n28168 , n28169 );
xor ( n28171 , n28168 , n28169 );
xor ( n28172 , n28079 , n28154 );
and ( n28173 , n18110 , n18386 );
and ( n28174 , n28172 , n28173 );
xor ( n28175 , n28172 , n28173 );
xor ( n28176 , n28083 , n28152 );
and ( n28177 , n18111 , n18386 );
and ( n28178 , n28176 , n28177 );
xor ( n28179 , n28176 , n28177 );
xor ( n28180 , n28087 , n28150 );
and ( n28181 , n18112 , n18386 );
and ( n28182 , n28180 , n28181 );
xor ( n28183 , n28180 , n28181 );
xor ( n28184 , n28091 , n28148 );
and ( n28185 , n18113 , n18386 );
and ( n28186 , n28184 , n28185 );
xor ( n28187 , n28184 , n28185 );
xor ( n28188 , n28095 , n28146 );
and ( n28189 , n18114 , n18386 );
and ( n28190 , n28188 , n28189 );
xor ( n28191 , n28188 , n28189 );
xor ( n28192 , n28099 , n28144 );
and ( n28193 , n18115 , n18386 );
and ( n28194 , n28192 , n28193 );
xor ( n28195 , n28192 , n28193 );
xor ( n28196 , n28103 , n28142 );
and ( n28197 , n18116 , n18386 );
and ( n28198 , n28196 , n28197 );
xor ( n28199 , n28196 , n28197 );
xor ( n28200 , n28107 , n28140 );
and ( n28201 , n18117 , n18386 );
and ( n28202 , n28200 , n28201 );
xor ( n28203 , n28200 , n28201 );
xor ( n28204 , n28111 , n28138 );
and ( n28205 , n18118 , n18386 );
and ( n28206 , n28204 , n28205 );
xor ( n28207 , n28204 , n28205 );
xor ( n28208 , n28115 , n28136 );
and ( n28209 , n18119 , n18386 );
and ( n28210 , n28208 , n28209 );
xor ( n28211 , n28208 , n28209 );
xor ( n28212 , n28119 , n28134 );
and ( n28213 , n18120 , n18386 );
and ( n28214 , n28212 , n28213 );
xor ( n28215 , n28212 , n28213 );
xor ( n28216 , n28123 , n28132 );
and ( n28217 , n18121 , n18386 );
and ( n28218 , n28216 , n28217 );
xor ( n28219 , n28216 , n28217 );
xor ( n28220 , n28127 , n28130 );
and ( n28221 , n18122 , n18386 );
and ( n28222 , n28220 , n28221 );
and ( n28223 , n28219 , n28222 );
or ( n28224 , n28218 , n28223 );
and ( n28225 , n28215 , n28224 );
or ( n28226 , n28214 , n28225 );
and ( n28227 , n28211 , n28226 );
or ( n28228 , n28210 , n28227 );
and ( n28229 , n28207 , n28228 );
or ( n28230 , n28206 , n28229 );
and ( n28231 , n28203 , n28230 );
or ( n28232 , n28202 , n28231 );
and ( n28233 , n28199 , n28232 );
or ( n28234 , n28198 , n28233 );
and ( n28235 , n28195 , n28234 );
or ( n28236 , n28194 , n28235 );
and ( n28237 , n28191 , n28236 );
or ( n28238 , n28190 , n28237 );
and ( n28239 , n28187 , n28238 );
or ( n28240 , n28186 , n28239 );
and ( n28241 , n28183 , n28240 );
or ( n28242 , n28182 , n28241 );
and ( n28243 , n28179 , n28242 );
or ( n28244 , n28178 , n28243 );
and ( n28245 , n28175 , n28244 );
or ( n28246 , n28174 , n28245 );
and ( n28247 , n28171 , n28246 );
or ( n28248 , n28170 , n28247 );
and ( n28249 , n28167 , n28248 );
or ( n28250 , n28166 , n28249 );
and ( n28251 , n28163 , n28250 );
or ( n28252 , n28162 , n28251 );
and ( n28253 , n18107 , n18384 );
and ( n28254 , n28252 , n28253 );
xor ( n28255 , n28252 , n28253 );
xor ( n28256 , n28163 , n28250 );
and ( n28257 , n18108 , n18384 );
and ( n28258 , n28256 , n28257 );
xor ( n28259 , n28256 , n28257 );
xor ( n28260 , n28167 , n28248 );
and ( n28261 , n18109 , n18384 );
and ( n28262 , n28260 , n28261 );
xor ( n28263 , n28260 , n28261 );
xor ( n28264 , n28171 , n28246 );
and ( n28265 , n18110 , n18384 );
and ( n28266 , n28264 , n28265 );
xor ( n28267 , n28264 , n28265 );
xor ( n28268 , n28175 , n28244 );
and ( n28269 , n18111 , n18384 );
and ( n28270 , n28268 , n28269 );
xor ( n28271 , n28268 , n28269 );
xor ( n28272 , n28179 , n28242 );
and ( n28273 , n18112 , n18384 );
and ( n28274 , n28272 , n28273 );
xor ( n28275 , n28272 , n28273 );
xor ( n28276 , n28183 , n28240 );
and ( n28277 , n18113 , n18384 );
and ( n28278 , n28276 , n28277 );
xor ( n28279 , n28276 , n28277 );
xor ( n28280 , n28187 , n28238 );
and ( n28281 , n18114 , n18384 );
and ( n28282 , n28280 , n28281 );
xor ( n28283 , n28280 , n28281 );
xor ( n28284 , n28191 , n28236 );
and ( n28285 , n18115 , n18384 );
and ( n28286 , n28284 , n28285 );
xor ( n28287 , n28284 , n28285 );
xor ( n28288 , n28195 , n28234 );
and ( n28289 , n18116 , n18384 );
and ( n28290 , n28288 , n28289 );
xor ( n28291 , n28288 , n28289 );
xor ( n28292 , n28199 , n28232 );
and ( n28293 , n18117 , n18384 );
and ( n28294 , n28292 , n28293 );
xor ( n28295 , n28292 , n28293 );
xor ( n28296 , n28203 , n28230 );
and ( n28297 , n18118 , n18384 );
and ( n28298 , n28296 , n28297 );
xor ( n28299 , n28296 , n28297 );
xor ( n28300 , n28207 , n28228 );
and ( n28301 , n18119 , n18384 );
and ( n28302 , n28300 , n28301 );
xor ( n28303 , n28300 , n28301 );
xor ( n28304 , n28211 , n28226 );
and ( n28305 , n18120 , n18384 );
and ( n28306 , n28304 , n28305 );
xor ( n28307 , n28304 , n28305 );
xor ( n28308 , n28215 , n28224 );
and ( n28309 , n18121 , n18384 );
and ( n28310 , n28308 , n28309 );
xor ( n28311 , n28308 , n28309 );
xor ( n28312 , n28219 , n28222 );
and ( n28313 , n18122 , n18384 );
and ( n28314 , n28312 , n28313 );
and ( n28315 , n28311 , n28314 );
or ( n28316 , n28310 , n28315 );
and ( n28317 , n28307 , n28316 );
or ( n28318 , n28306 , n28317 );
and ( n28319 , n28303 , n28318 );
or ( n28320 , n28302 , n28319 );
and ( n28321 , n28299 , n28320 );
or ( n28322 , n28298 , n28321 );
and ( n28323 , n28295 , n28322 );
or ( n28324 , n28294 , n28323 );
and ( n28325 , n28291 , n28324 );
or ( n28326 , n28290 , n28325 );
and ( n28327 , n28287 , n28326 );
or ( n28328 , n28286 , n28327 );
and ( n28329 , n28283 , n28328 );
or ( n28330 , n28282 , n28329 );
and ( n28331 , n28279 , n28330 );
or ( n28332 , n28278 , n28331 );
and ( n28333 , n28275 , n28332 );
or ( n28334 , n28274 , n28333 );
and ( n28335 , n28271 , n28334 );
or ( n28336 , n28270 , n28335 );
and ( n28337 , n28267 , n28336 );
or ( n28338 , n28266 , n28337 );
and ( n28339 , n28263 , n28338 );
or ( n28340 , n28262 , n28339 );
and ( n28341 , n28259 , n28340 );
or ( n28342 , n28258 , n28341 );
and ( n28343 , n28255 , n28342 );
or ( n28344 , n28254 , n28343 );
and ( n28345 , n18107 , n18382 );
and ( n28346 , n28344 , n28345 );
xor ( n28347 , n28344 , n28345 );
xor ( n28348 , n28255 , n28342 );
and ( n28349 , n18108 , n18382 );
and ( n28350 , n28348 , n28349 );
xor ( n28351 , n28348 , n28349 );
xor ( n28352 , n28259 , n28340 );
and ( n28353 , n18109 , n18382 );
and ( n28354 , n28352 , n28353 );
xor ( n28355 , n28352 , n28353 );
xor ( n28356 , n28263 , n28338 );
and ( n28357 , n18110 , n18382 );
and ( n28358 , n28356 , n28357 );
xor ( n28359 , n28356 , n28357 );
xor ( n28360 , n28267 , n28336 );
and ( n28361 , n18111 , n18382 );
and ( n28362 , n28360 , n28361 );
xor ( n28363 , n28360 , n28361 );
xor ( n28364 , n28271 , n28334 );
and ( n28365 , n18112 , n18382 );
and ( n28366 , n28364 , n28365 );
xor ( n28367 , n28364 , n28365 );
xor ( n28368 , n28275 , n28332 );
and ( n28369 , n18113 , n18382 );
and ( n28370 , n28368 , n28369 );
xor ( n28371 , n28368 , n28369 );
xor ( n28372 , n28279 , n28330 );
and ( n28373 , n18114 , n18382 );
and ( n28374 , n28372 , n28373 );
xor ( n28375 , n28372 , n28373 );
xor ( n28376 , n28283 , n28328 );
and ( n28377 , n18115 , n18382 );
and ( n28378 , n28376 , n28377 );
xor ( n28379 , n28376 , n28377 );
xor ( n28380 , n28287 , n28326 );
and ( n28381 , n18116 , n18382 );
and ( n28382 , n28380 , n28381 );
xor ( n28383 , n28380 , n28381 );
xor ( n28384 , n28291 , n28324 );
and ( n28385 , n18117 , n18382 );
and ( n28386 , n28384 , n28385 );
xor ( n28387 , n28384 , n28385 );
xor ( n28388 , n28295 , n28322 );
and ( n28389 , n18118 , n18382 );
and ( n28390 , n28388 , n28389 );
xor ( n28391 , n28388 , n28389 );
xor ( n28392 , n28299 , n28320 );
and ( n28393 , n18119 , n18382 );
and ( n28394 , n28392 , n28393 );
xor ( n28395 , n28392 , n28393 );
xor ( n28396 , n28303 , n28318 );
and ( n28397 , n18120 , n18382 );
and ( n28398 , n28396 , n28397 );
xor ( n28399 , n28396 , n28397 );
xor ( n28400 , n28307 , n28316 );
and ( n28401 , n18121 , n18382 );
and ( n28402 , n28400 , n28401 );
xor ( n28403 , n28400 , n28401 );
xor ( n28404 , n28311 , n28314 );
and ( n28405 , n18122 , n18382 );
and ( n28406 , n28404 , n28405 );
and ( n28407 , n28403 , n28406 );
or ( n28408 , n28402 , n28407 );
and ( n28409 , n28399 , n28408 );
or ( n28410 , n28398 , n28409 );
and ( n28411 , n28395 , n28410 );
or ( n28412 , n28394 , n28411 );
and ( n28413 , n28391 , n28412 );
or ( n28414 , n28390 , n28413 );
and ( n28415 , n28387 , n28414 );
or ( n28416 , n28386 , n28415 );
and ( n28417 , n28383 , n28416 );
or ( n28418 , n28382 , n28417 );
and ( n28419 , n28379 , n28418 );
or ( n28420 , n28378 , n28419 );
and ( n28421 , n28375 , n28420 );
or ( n28422 , n28374 , n28421 );
and ( n28423 , n28371 , n28422 );
or ( n28424 , n28370 , n28423 );
and ( n28425 , n28367 , n28424 );
or ( n28426 , n28366 , n28425 );
and ( n28427 , n28363 , n28426 );
or ( n28428 , n28362 , n28427 );
and ( n28429 , n28359 , n28428 );
or ( n28430 , n28358 , n28429 );
and ( n28431 , n28355 , n28430 );
or ( n28432 , n28354 , n28431 );
and ( n28433 , n28351 , n28432 );
or ( n28434 , n28350 , n28433 );
and ( n28435 , n28347 , n28434 );
or ( n28436 , n28346 , n28435 );
and ( n28437 , n18107 , n18380 );
and ( n28438 , n28436 , n28437 );
xor ( n28439 , n28436 , n28437 );
xor ( n28440 , n28347 , n28434 );
and ( n28441 , n18108 , n18380 );
and ( n28442 , n28440 , n28441 );
xor ( n28443 , n28440 , n28441 );
xor ( n28444 , n28351 , n28432 );
and ( n28445 , n18109 , n18380 );
and ( n28446 , n28444 , n28445 );
xor ( n28447 , n28444 , n28445 );
xor ( n28448 , n28355 , n28430 );
and ( n28449 , n18110 , n18380 );
and ( n28450 , n28448 , n28449 );
xor ( n28451 , n28448 , n28449 );
xor ( n28452 , n28359 , n28428 );
and ( n28453 , n18111 , n18380 );
and ( n28454 , n28452 , n28453 );
xor ( n28455 , n28452 , n28453 );
xor ( n28456 , n28363 , n28426 );
and ( n28457 , n18112 , n18380 );
and ( n28458 , n28456 , n28457 );
xor ( n28459 , n28456 , n28457 );
xor ( n28460 , n28367 , n28424 );
and ( n28461 , n18113 , n18380 );
and ( n28462 , n28460 , n28461 );
xor ( n28463 , n28460 , n28461 );
xor ( n28464 , n28371 , n28422 );
and ( n28465 , n18114 , n18380 );
and ( n28466 , n28464 , n28465 );
xor ( n28467 , n28464 , n28465 );
xor ( n28468 , n28375 , n28420 );
and ( n28469 , n18115 , n18380 );
and ( n28470 , n28468 , n28469 );
xor ( n28471 , n28468 , n28469 );
xor ( n28472 , n28379 , n28418 );
and ( n28473 , n18116 , n18380 );
and ( n28474 , n28472 , n28473 );
xor ( n28475 , n28472 , n28473 );
xor ( n28476 , n28383 , n28416 );
and ( n28477 , n18117 , n18380 );
and ( n28478 , n28476 , n28477 );
xor ( n28479 , n28476 , n28477 );
xor ( n28480 , n28387 , n28414 );
and ( n28481 , n18118 , n18380 );
and ( n28482 , n28480 , n28481 );
xor ( n28483 , n28480 , n28481 );
xor ( n28484 , n28391 , n28412 );
and ( n28485 , n18119 , n18380 );
and ( n28486 , n28484 , n28485 );
xor ( n28487 , n28484 , n28485 );
xor ( n28488 , n28395 , n28410 );
and ( n28489 , n18120 , n18380 );
and ( n28490 , n28488 , n28489 );
xor ( n28491 , n28488 , n28489 );
xor ( n28492 , n28399 , n28408 );
and ( n28493 , n18121 , n18380 );
and ( n28494 , n28492 , n28493 );
xor ( n28495 , n28492 , n28493 );
xor ( n28496 , n28403 , n28406 );
and ( n28497 , n18122 , n18380 );
and ( n28498 , n28496 , n28497 );
and ( n28499 , n28495 , n28498 );
or ( n28500 , n28494 , n28499 );
and ( n28501 , n28491 , n28500 );
or ( n28502 , n28490 , n28501 );
and ( n28503 , n28487 , n28502 );
or ( n28504 , n28486 , n28503 );
and ( n28505 , n28483 , n28504 );
or ( n28506 , n28482 , n28505 );
and ( n28507 , n28479 , n28506 );
or ( n28508 , n28478 , n28507 );
and ( n28509 , n28475 , n28508 );
or ( n28510 , n28474 , n28509 );
and ( n28511 , n28471 , n28510 );
or ( n28512 , n28470 , n28511 );
and ( n28513 , n28467 , n28512 );
or ( n28514 , n28466 , n28513 );
and ( n28515 , n28463 , n28514 );
or ( n28516 , n28462 , n28515 );
and ( n28517 , n28459 , n28516 );
or ( n28518 , n28458 , n28517 );
and ( n28519 , n28455 , n28518 );
or ( n28520 , n28454 , n28519 );
and ( n28521 , n28451 , n28520 );
or ( n28522 , n28450 , n28521 );
and ( n28523 , n28447 , n28522 );
or ( n28524 , n28446 , n28523 );
and ( n28525 , n28443 , n28524 );
or ( n28526 , n28442 , n28525 );
and ( n28527 , n28439 , n28526 );
or ( n28528 , n28438 , n28527 );
and ( n28529 , n18107 , n18378 );
and ( n28530 , n28528 , n28529 );
xor ( n28531 , n28528 , n28529 );
xor ( n28532 , n28439 , n28526 );
and ( n28533 , n18108 , n18378 );
and ( n28534 , n28532 , n28533 );
xor ( n28535 , n28532 , n28533 );
xor ( n28536 , n28443 , n28524 );
and ( n28537 , n18109 , n18378 );
and ( n28538 , n28536 , n28537 );
xor ( n28539 , n28536 , n28537 );
xor ( n28540 , n28447 , n28522 );
and ( n28541 , n18110 , n18378 );
and ( n28542 , n28540 , n28541 );
xor ( n28543 , n28540 , n28541 );
xor ( n28544 , n28451 , n28520 );
and ( n28545 , n18111 , n18378 );
and ( n28546 , n28544 , n28545 );
xor ( n28547 , n28544 , n28545 );
xor ( n28548 , n28455 , n28518 );
and ( n28549 , n18112 , n18378 );
and ( n28550 , n28548 , n28549 );
xor ( n28551 , n28548 , n28549 );
xor ( n28552 , n28459 , n28516 );
and ( n28553 , n18113 , n18378 );
and ( n28554 , n28552 , n28553 );
xor ( n28555 , n28552 , n28553 );
xor ( n28556 , n28463 , n28514 );
and ( n28557 , n18114 , n18378 );
and ( n28558 , n28556 , n28557 );
xor ( n28559 , n28556 , n28557 );
xor ( n28560 , n28467 , n28512 );
and ( n28561 , n18115 , n18378 );
and ( n28562 , n28560 , n28561 );
xor ( n28563 , n28560 , n28561 );
xor ( n28564 , n28471 , n28510 );
and ( n28565 , n18116 , n18378 );
and ( n28566 , n28564 , n28565 );
xor ( n28567 , n28564 , n28565 );
xor ( n28568 , n28475 , n28508 );
and ( n28569 , n18117 , n18378 );
and ( n28570 , n28568 , n28569 );
xor ( n28571 , n28568 , n28569 );
xor ( n28572 , n28479 , n28506 );
and ( n28573 , n18118 , n18378 );
and ( n28574 , n28572 , n28573 );
xor ( n28575 , n28572 , n28573 );
xor ( n28576 , n28483 , n28504 );
and ( n28577 , n18119 , n18378 );
and ( n28578 , n28576 , n28577 );
xor ( n28579 , n28576 , n28577 );
xor ( n28580 , n28487 , n28502 );
and ( n28581 , n18120 , n18378 );
and ( n28582 , n28580 , n28581 );
xor ( n28583 , n28580 , n28581 );
xor ( n28584 , n28491 , n28500 );
and ( n28585 , n18121 , n18378 );
and ( n28586 , n28584 , n28585 );
xor ( n28587 , n28584 , n28585 );
xor ( n28588 , n28495 , n28498 );
and ( n28589 , n18122 , n18378 );
and ( n28590 , n28588 , n28589 );
and ( n28591 , n28587 , n28590 );
or ( n28592 , n28586 , n28591 );
and ( n28593 , n28583 , n28592 );
or ( n28594 , n28582 , n28593 );
and ( n28595 , n28579 , n28594 );
or ( n28596 , n28578 , n28595 );
and ( n28597 , n28575 , n28596 );
or ( n28598 , n28574 , n28597 );
and ( n28599 , n28571 , n28598 );
or ( n28600 , n28570 , n28599 );
and ( n28601 , n28567 , n28600 );
or ( n28602 , n28566 , n28601 );
and ( n28603 , n28563 , n28602 );
or ( n28604 , n28562 , n28603 );
and ( n28605 , n28559 , n28604 );
or ( n28606 , n28558 , n28605 );
and ( n28607 , n28555 , n28606 );
or ( n28608 , n28554 , n28607 );
and ( n28609 , n28551 , n28608 );
or ( n28610 , n28550 , n28609 );
and ( n28611 , n28547 , n28610 );
or ( n28612 , n28546 , n28611 );
and ( n28613 , n28543 , n28612 );
or ( n28614 , n28542 , n28613 );
and ( n28615 , n28539 , n28614 );
or ( n28616 , n28538 , n28615 );
and ( n28617 , n28535 , n28616 );
or ( n28618 , n28534 , n28617 );
and ( n28619 , n28531 , n28618 );
or ( n28620 , n28530 , n28619 );
and ( n28621 , n18107 , n18376 );
and ( n28622 , n28620 , n28621 );
xor ( n28623 , n28620 , n28621 );
xor ( n28624 , n28531 , n28618 );
and ( n28625 , n18108 , n18376 );
and ( n28626 , n28624 , n28625 );
xor ( n28627 , n28624 , n28625 );
xor ( n28628 , n28535 , n28616 );
and ( n28629 , n18109 , n18376 );
and ( n28630 , n28628 , n28629 );
xor ( n28631 , n28628 , n28629 );
xor ( n28632 , n28539 , n28614 );
and ( n28633 , n18110 , n18376 );
and ( n28634 , n28632 , n28633 );
xor ( n28635 , n28632 , n28633 );
xor ( n28636 , n28543 , n28612 );
and ( n28637 , n18111 , n18376 );
and ( n28638 , n28636 , n28637 );
xor ( n28639 , n28636 , n28637 );
xor ( n28640 , n28547 , n28610 );
and ( n28641 , n18112 , n18376 );
and ( n28642 , n28640 , n28641 );
xor ( n28643 , n28640 , n28641 );
xor ( n28644 , n28551 , n28608 );
and ( n28645 , n18113 , n18376 );
and ( n28646 , n28644 , n28645 );
xor ( n28647 , n28644 , n28645 );
xor ( n28648 , n28555 , n28606 );
and ( n28649 , n18114 , n18376 );
and ( n28650 , n28648 , n28649 );
xor ( n28651 , n28648 , n28649 );
xor ( n28652 , n28559 , n28604 );
and ( n28653 , n18115 , n18376 );
and ( n28654 , n28652 , n28653 );
xor ( n28655 , n28652 , n28653 );
xor ( n28656 , n28563 , n28602 );
and ( n28657 , n18116 , n18376 );
and ( n28658 , n28656 , n28657 );
xor ( n28659 , n28656 , n28657 );
xor ( n28660 , n28567 , n28600 );
and ( n28661 , n18117 , n18376 );
and ( n28662 , n28660 , n28661 );
xor ( n28663 , n28660 , n28661 );
xor ( n28664 , n28571 , n28598 );
and ( n28665 , n18118 , n18376 );
and ( n28666 , n28664 , n28665 );
xor ( n28667 , n28664 , n28665 );
xor ( n28668 , n28575 , n28596 );
and ( n28669 , n18119 , n18376 );
and ( n28670 , n28668 , n28669 );
xor ( n28671 , n28668 , n28669 );
xor ( n28672 , n28579 , n28594 );
and ( n28673 , n18120 , n18376 );
and ( n28674 , n28672 , n28673 );
xor ( n28675 , n28672 , n28673 );
xor ( n28676 , n28583 , n28592 );
and ( n28677 , n18121 , n18376 );
and ( n28678 , n28676 , n28677 );
xor ( n28679 , n28676 , n28677 );
xor ( n28680 , n28587 , n28590 );
and ( n28681 , n18122 , n18376 );
and ( n28682 , n28680 , n28681 );
and ( n28683 , n28679 , n28682 );
or ( n28684 , n28678 , n28683 );
and ( n28685 , n28675 , n28684 );
or ( n28686 , n28674 , n28685 );
and ( n28687 , n28671 , n28686 );
or ( n28688 , n28670 , n28687 );
and ( n28689 , n28667 , n28688 );
or ( n28690 , n28666 , n28689 );
and ( n28691 , n28663 , n28690 );
or ( n28692 , n28662 , n28691 );
and ( n28693 , n28659 , n28692 );
or ( n28694 , n28658 , n28693 );
and ( n28695 , n28655 , n28694 );
or ( n28696 , n28654 , n28695 );
and ( n28697 , n28651 , n28696 );
or ( n28698 , n28650 , n28697 );
and ( n28699 , n28647 , n28698 );
or ( n28700 , n28646 , n28699 );
and ( n28701 , n28643 , n28700 );
or ( n28702 , n28642 , n28701 );
and ( n28703 , n28639 , n28702 );
or ( n28704 , n28638 , n28703 );
and ( n28705 , n28635 , n28704 );
or ( n28706 , n28634 , n28705 );
and ( n28707 , n28631 , n28706 );
or ( n28708 , n28630 , n28707 );
and ( n28709 , n28627 , n28708 );
or ( n28710 , n28626 , n28709 );
and ( n28711 , n28623 , n28710 );
or ( n28712 , n28622 , n28711 );
and ( n28713 , n18107 , n18374 );
and ( n28714 , n28712 , n28713 );
xor ( n28715 , n28712 , n28713 );
xor ( n28716 , n28623 , n28710 );
and ( n28717 , n18108 , n18374 );
and ( n28718 , n28716 , n28717 );
xor ( n28719 , n28716 , n28717 );
xor ( n28720 , n28627 , n28708 );
and ( n28721 , n18109 , n18374 );
and ( n28722 , n28720 , n28721 );
xor ( n28723 , n28720 , n28721 );
xor ( n28724 , n28631 , n28706 );
and ( n28725 , n18110 , n18374 );
and ( n28726 , n28724 , n28725 );
xor ( n28727 , n28724 , n28725 );
xor ( n28728 , n28635 , n28704 );
and ( n28729 , n18111 , n18374 );
and ( n28730 , n28728 , n28729 );
xor ( n28731 , n28728 , n28729 );
xor ( n28732 , n28639 , n28702 );
and ( n28733 , n18112 , n18374 );
and ( n28734 , n28732 , n28733 );
xor ( n28735 , n28732 , n28733 );
xor ( n28736 , n28643 , n28700 );
and ( n28737 , n18113 , n18374 );
and ( n28738 , n28736 , n28737 );
xor ( n28739 , n28736 , n28737 );
xor ( n28740 , n28647 , n28698 );
and ( n28741 , n18114 , n18374 );
and ( n28742 , n28740 , n28741 );
xor ( n28743 , n28740 , n28741 );
xor ( n28744 , n28651 , n28696 );
and ( n28745 , n18115 , n18374 );
and ( n28746 , n28744 , n28745 );
xor ( n28747 , n28744 , n28745 );
xor ( n28748 , n28655 , n28694 );
and ( n28749 , n18116 , n18374 );
and ( n28750 , n28748 , n28749 );
xor ( n28751 , n28748 , n28749 );
xor ( n28752 , n28659 , n28692 );
and ( n28753 , n18117 , n18374 );
and ( n28754 , n28752 , n28753 );
xor ( n28755 , n28752 , n28753 );
xor ( n28756 , n28663 , n28690 );
and ( n28757 , n18118 , n18374 );
and ( n28758 , n28756 , n28757 );
xor ( n28759 , n28756 , n28757 );
xor ( n28760 , n28667 , n28688 );
and ( n28761 , n18119 , n18374 );
and ( n28762 , n28760 , n28761 );
xor ( n28763 , n28760 , n28761 );
xor ( n28764 , n28671 , n28686 );
and ( n28765 , n18120 , n18374 );
and ( n28766 , n28764 , n28765 );
xor ( n28767 , n28764 , n28765 );
xor ( n28768 , n28675 , n28684 );
and ( n28769 , n18121 , n18374 );
and ( n28770 , n28768 , n28769 );
xor ( n28771 , n28768 , n28769 );
xor ( n28772 , n28679 , n28682 );
and ( n28773 , n18122 , n18374 );
and ( n28774 , n28772 , n28773 );
and ( n28775 , n28771 , n28774 );
or ( n28776 , n28770 , n28775 );
and ( n28777 , n28767 , n28776 );
or ( n28778 , n28766 , n28777 );
and ( n28779 , n28763 , n28778 );
or ( n28780 , n28762 , n28779 );
and ( n28781 , n28759 , n28780 );
or ( n28782 , n28758 , n28781 );
and ( n28783 , n28755 , n28782 );
or ( n28784 , n28754 , n28783 );
and ( n28785 , n28751 , n28784 );
or ( n28786 , n28750 , n28785 );
and ( n28787 , n28747 , n28786 );
or ( n28788 , n28746 , n28787 );
and ( n28789 , n28743 , n28788 );
or ( n28790 , n28742 , n28789 );
and ( n28791 , n28739 , n28790 );
or ( n28792 , n28738 , n28791 );
and ( n28793 , n28735 , n28792 );
or ( n28794 , n28734 , n28793 );
and ( n28795 , n28731 , n28794 );
or ( n28796 , n28730 , n28795 );
and ( n28797 , n28727 , n28796 );
or ( n28798 , n28726 , n28797 );
and ( n28799 , n28723 , n28798 );
or ( n28800 , n28722 , n28799 );
and ( n28801 , n28719 , n28800 );
or ( n28802 , n28718 , n28801 );
and ( n28803 , n28715 , n28802 );
or ( n28804 , n28714 , n28803 );
and ( n28805 , n18107 , n18372 );
xor ( n28806 , n28804 , n28805 );
xor ( n28807 , n28715 , n28802 );
and ( n28808 , n18108 , n18372 );
and ( n28809 , n28807 , n28808 );
xor ( n28810 , n28807 , n28808 );
xor ( n28811 , n28719 , n28800 );
and ( n28812 , n18109 , n18372 );
and ( n28813 , n28811 , n28812 );
xor ( n28814 , n28811 , n28812 );
xor ( n28815 , n28723 , n28798 );
and ( n28816 , n18110 , n18372 );
and ( n28817 , n28815 , n28816 );
xor ( n28818 , n28815 , n28816 );
xor ( n28819 , n28727 , n28796 );
and ( n28820 , n18111 , n18372 );
and ( n28821 , n28819 , n28820 );
xor ( n28822 , n28819 , n28820 );
xor ( n28823 , n28731 , n28794 );
and ( n28824 , n18112 , n18372 );
and ( n28825 , n28823 , n28824 );
xor ( n28826 , n28823 , n28824 );
xor ( n28827 , n28735 , n28792 );
and ( n28828 , n18113 , n18372 );
and ( n28829 , n28827 , n28828 );
xor ( n28830 , n28827 , n28828 );
xor ( n28831 , n28739 , n28790 );
and ( n28832 , n18114 , n18372 );
and ( n28833 , n28831 , n28832 );
xor ( n28834 , n28831 , n28832 );
xor ( n28835 , n28743 , n28788 );
and ( n28836 , n18115 , n18372 );
and ( n28837 , n28835 , n28836 );
xor ( n28838 , n28835 , n28836 );
xor ( n28839 , n28747 , n28786 );
and ( n28840 , n18116 , n18372 );
and ( n28841 , n28839 , n28840 );
xor ( n28842 , n28839 , n28840 );
xor ( n28843 , n28751 , n28784 );
and ( n28844 , n18117 , n18372 );
and ( n28845 , n28843 , n28844 );
xor ( n28846 , n28843 , n28844 );
xor ( n28847 , n28755 , n28782 );
and ( n28848 , n18118 , n18372 );
and ( n28849 , n28847 , n28848 );
xor ( n28850 , n28847 , n28848 );
xor ( n28851 , n28759 , n28780 );
and ( n28852 , n18119 , n18372 );
and ( n28853 , n28851 , n28852 );
xor ( n28854 , n28851 , n28852 );
xor ( n28855 , n28763 , n28778 );
and ( n28856 , n18120 , n18372 );
and ( n28857 , n28855 , n28856 );
xor ( n28858 , n28855 , n28856 );
xor ( n28859 , n28767 , n28776 );
and ( n28860 , n18121 , n18372 );
and ( n28861 , n28859 , n28860 );
xor ( n28862 , n28859 , n28860 );
xor ( n28863 , n28771 , n28774 );
and ( n28864 , n18122 , n18372 );
and ( n28865 , n28863 , n28864 );
and ( n28866 , n28862 , n28865 );
or ( n28867 , n28861 , n28866 );
and ( n28868 , n28858 , n28867 );
or ( n28869 , n28857 , n28868 );
and ( n28870 , n28854 , n28869 );
or ( n28871 , n28853 , n28870 );
and ( n28872 , n28850 , n28871 );
or ( n28873 , n28849 , n28872 );
and ( n28874 , n28846 , n28873 );
or ( n28875 , n28845 , n28874 );
and ( n28876 , n28842 , n28875 );
or ( n28877 , n28841 , n28876 );
and ( n28878 , n28838 , n28877 );
or ( n28879 , n28837 , n28878 );
and ( n28880 , n28834 , n28879 );
or ( n28881 , n28833 , n28880 );
and ( n28882 , n28830 , n28881 );
or ( n28883 , n28829 , n28882 );
and ( n28884 , n28826 , n28883 );
or ( n28885 , n28825 , n28884 );
and ( n28886 , n28822 , n28885 );
or ( n28887 , n28821 , n28886 );
and ( n28888 , n28818 , n28887 );
or ( n28889 , n28817 , n28888 );
and ( n28890 , n28814 , n28889 );
or ( n28891 , n28813 , n28890 );
and ( n28892 , n28810 , n28891 );
or ( n28893 , n28809 , n28892 );
xor ( n28894 , n28806 , n28893 );
and ( n28895 , n18108 , n18370 );
xor ( n28896 , n28894 , n28895 );
xor ( n28897 , n28810 , n28891 );
and ( n28898 , n18109 , n18370 );
and ( n28899 , n28897 , n28898 );
xor ( n28900 , n28897 , n28898 );
xor ( n28901 , n28814 , n28889 );
and ( n28902 , n18110 , n18370 );
and ( n28903 , n28901 , n28902 );
xor ( n28904 , n28901 , n28902 );
xor ( n28905 , n28818 , n28887 );
and ( n28906 , n18111 , n18370 );
and ( n28907 , n28905 , n28906 );
xor ( n28908 , n28905 , n28906 );
xor ( n28909 , n28822 , n28885 );
and ( n28910 , n18112 , n18370 );
and ( n28911 , n28909 , n28910 );
xor ( n28912 , n28909 , n28910 );
xor ( n28913 , n28826 , n28883 );
and ( n28914 , n18113 , n18370 );
and ( n28915 , n28913 , n28914 );
xor ( n28916 , n28913 , n28914 );
xor ( n28917 , n28830 , n28881 );
and ( n28918 , n18114 , n18370 );
and ( n28919 , n28917 , n28918 );
xor ( n28920 , n28917 , n28918 );
xor ( n28921 , n28834 , n28879 );
and ( n28922 , n18115 , n18370 );
and ( n28923 , n28921 , n28922 );
xor ( n28924 , n28921 , n28922 );
xor ( n28925 , n28838 , n28877 );
and ( n28926 , n18116 , n18370 );
and ( n28927 , n28925 , n28926 );
xor ( n28928 , n28925 , n28926 );
xor ( n28929 , n28842 , n28875 );
and ( n28930 , n18117 , n18370 );
and ( n28931 , n28929 , n28930 );
xor ( n28932 , n28929 , n28930 );
xor ( n28933 , n28846 , n28873 );
and ( n28934 , n18118 , n18370 );
and ( n28935 , n28933 , n28934 );
xor ( n28936 , n28933 , n28934 );
xor ( n28937 , n28850 , n28871 );
and ( n28938 , n18119 , n18370 );
and ( n28939 , n28937 , n28938 );
xor ( n28940 , n28937 , n28938 );
xor ( n28941 , n28854 , n28869 );
and ( n28942 , n18120 , n18370 );
and ( n28943 , n28941 , n28942 );
xor ( n28944 , n28941 , n28942 );
xor ( n28945 , n28858 , n28867 );
and ( n28946 , n18121 , n18370 );
and ( n28947 , n28945 , n28946 );
xor ( n28948 , n28945 , n28946 );
xor ( n28949 , n28862 , n28865 );
and ( n28950 , n18122 , n18370 );
and ( n28951 , n28949 , n28950 );
and ( n28952 , n28948 , n28951 );
or ( n28953 , n28947 , n28952 );
and ( n28954 , n28944 , n28953 );
or ( n28955 , n28943 , n28954 );
and ( n28956 , n28940 , n28955 );
or ( n28957 , n28939 , n28956 );
and ( n28958 , n28936 , n28957 );
or ( n28959 , n28935 , n28958 );
and ( n28960 , n28932 , n28959 );
or ( n28961 , n28931 , n28960 );
and ( n28962 , n28928 , n28961 );
or ( n28963 , n28927 , n28962 );
and ( n28964 , n28924 , n28963 );
or ( n28965 , n28923 , n28964 );
and ( n28966 , n28920 , n28965 );
or ( n28967 , n28919 , n28966 );
and ( n28968 , n28916 , n28967 );
or ( n28969 , n28915 , n28968 );
and ( n28970 , n28912 , n28969 );
or ( n28971 , n28911 , n28970 );
and ( n28972 , n28908 , n28971 );
or ( n28973 , n28907 , n28972 );
and ( n28974 , n28904 , n28973 );
or ( n28975 , n28903 , n28974 );
and ( n28976 , n28900 , n28975 );
or ( n28977 , n28899 , n28976 );
xor ( n28978 , n28896 , n28977 );
and ( n28979 , n18109 , n18368 );
xor ( n28980 , n28978 , n28979 );
xor ( n28981 , n28900 , n28975 );
and ( n28982 , n18110 , n18368 );
and ( n28983 , n28981 , n28982 );
xor ( n28984 , n28981 , n28982 );
xor ( n28985 , n28904 , n28973 );
and ( n28986 , n18111 , n18368 );
and ( n28987 , n28985 , n28986 );
xor ( n28988 , n28985 , n28986 );
xor ( n28989 , n28908 , n28971 );
and ( n28990 , n18112 , n18368 );
and ( n28991 , n28989 , n28990 );
xor ( n28992 , n28989 , n28990 );
xor ( n28993 , n28912 , n28969 );
and ( n28994 , n18113 , n18368 );
and ( n28995 , n28993 , n28994 );
xor ( n28996 , n28993 , n28994 );
xor ( n28997 , n28916 , n28967 );
and ( n28998 , n18114 , n18368 );
and ( n28999 , n28997 , n28998 );
xor ( n29000 , n28997 , n28998 );
xor ( n29001 , n28920 , n28965 );
and ( n29002 , n18115 , n18368 );
and ( n29003 , n29001 , n29002 );
xor ( n29004 , n29001 , n29002 );
xor ( n29005 , n28924 , n28963 );
and ( n29006 , n18116 , n18368 );
and ( n29007 , n29005 , n29006 );
xor ( n29008 , n29005 , n29006 );
xor ( n29009 , n28928 , n28961 );
and ( n29010 , n18117 , n18368 );
and ( n29011 , n29009 , n29010 );
xor ( n29012 , n29009 , n29010 );
xor ( n29013 , n28932 , n28959 );
and ( n29014 , n18118 , n18368 );
and ( n29015 , n29013 , n29014 );
xor ( n29016 , n29013 , n29014 );
xor ( n29017 , n28936 , n28957 );
and ( n29018 , n18119 , n18368 );
and ( n29019 , n29017 , n29018 );
xor ( n29020 , n29017 , n29018 );
xor ( n29021 , n28940 , n28955 );
and ( n29022 , n18120 , n18368 );
and ( n29023 , n29021 , n29022 );
xor ( n29024 , n29021 , n29022 );
xor ( n29025 , n28944 , n28953 );
and ( n29026 , n18121 , n18368 );
and ( n29027 , n29025 , n29026 );
xor ( n29028 , n29025 , n29026 );
xor ( n29029 , n28948 , n28951 );
and ( n29030 , n18122 , n18368 );
and ( n29031 , n29029 , n29030 );
and ( n29032 , n29028 , n29031 );
or ( n29033 , n29027 , n29032 );
and ( n29034 , n29024 , n29033 );
or ( n29035 , n29023 , n29034 );
and ( n29036 , n29020 , n29035 );
or ( n29037 , n29019 , n29036 );
and ( n29038 , n29016 , n29037 );
or ( n29039 , n29015 , n29038 );
and ( n29040 , n29012 , n29039 );
or ( n29041 , n29011 , n29040 );
and ( n29042 , n29008 , n29041 );
or ( n29043 , n29007 , n29042 );
and ( n29044 , n29004 , n29043 );
or ( n29045 , n29003 , n29044 );
and ( n29046 , n29000 , n29045 );
or ( n29047 , n28999 , n29046 );
and ( n29048 , n28996 , n29047 );
or ( n29049 , n28995 , n29048 );
and ( n29050 , n28992 , n29049 );
or ( n29051 , n28991 , n29050 );
and ( n29052 , n28988 , n29051 );
or ( n29053 , n28987 , n29052 );
and ( n29054 , n28984 , n29053 );
or ( n29055 , n28983 , n29054 );
xor ( n29056 , n28980 , n29055 );
and ( n29057 , n18110 , n18366 );
xor ( n29058 , n29056 , n29057 );
xor ( n29059 , n28984 , n29053 );
and ( n29060 , n18111 , n18366 );
and ( n29061 , n29059 , n29060 );
xor ( n29062 , n29059 , n29060 );
xor ( n29063 , n28988 , n29051 );
and ( n29064 , n18112 , n18366 );
and ( n29065 , n29063 , n29064 );
xor ( n29066 , n29063 , n29064 );
xor ( n29067 , n28992 , n29049 );
and ( n29068 , n18113 , n18366 );
and ( n29069 , n29067 , n29068 );
xor ( n29070 , n29067 , n29068 );
xor ( n29071 , n28996 , n29047 );
and ( n29072 , n18114 , n18366 );
and ( n29073 , n29071 , n29072 );
xor ( n29074 , n29071 , n29072 );
xor ( n29075 , n29000 , n29045 );
and ( n29076 , n18115 , n18366 );
and ( n29077 , n29075 , n29076 );
xor ( n29078 , n29075 , n29076 );
xor ( n29079 , n29004 , n29043 );
and ( n29080 , n18116 , n18366 );
and ( n29081 , n29079 , n29080 );
xor ( n29082 , n29079 , n29080 );
xor ( n29083 , n29008 , n29041 );
and ( n29084 , n18117 , n18366 );
and ( n29085 , n29083 , n29084 );
xor ( n29086 , n29083 , n29084 );
xor ( n29087 , n29012 , n29039 );
and ( n29088 , n18118 , n18366 );
and ( n29089 , n29087 , n29088 );
xor ( n29090 , n29087 , n29088 );
xor ( n29091 , n29016 , n29037 );
and ( n29092 , n18119 , n18366 );
and ( n29093 , n29091 , n29092 );
xor ( n29094 , n29091 , n29092 );
xor ( n29095 , n29020 , n29035 );
and ( n29096 , n18120 , n18366 );
and ( n29097 , n29095 , n29096 );
xor ( n29098 , n29095 , n29096 );
xor ( n29099 , n29024 , n29033 );
and ( n29100 , n18121 , n18366 );
and ( n29101 , n29099 , n29100 );
xor ( n29102 , n29099 , n29100 );
xor ( n29103 , n29028 , n29031 );
and ( n29104 , n18122 , n18366 );
and ( n29105 , n29103 , n29104 );
and ( n29106 , n29102 , n29105 );
or ( n29107 , n29101 , n29106 );
and ( n29108 , n29098 , n29107 );
or ( n29109 , n29097 , n29108 );
and ( n29110 , n29094 , n29109 );
or ( n29111 , n29093 , n29110 );
and ( n29112 , n29090 , n29111 );
or ( n29113 , n29089 , n29112 );
and ( n29114 , n29086 , n29113 );
or ( n29115 , n29085 , n29114 );
and ( n29116 , n29082 , n29115 );
or ( n29117 , n29081 , n29116 );
and ( n29118 , n29078 , n29117 );
or ( n29119 , n29077 , n29118 );
and ( n29120 , n29074 , n29119 );
or ( n29121 , n29073 , n29120 );
and ( n29122 , n29070 , n29121 );
or ( n29123 , n29069 , n29122 );
and ( n29124 , n29066 , n29123 );
or ( n29125 , n29065 , n29124 );
and ( n29126 , n29062 , n29125 );
or ( n29127 , n29061 , n29126 );
xor ( n29128 , n29058 , n29127 );
and ( n29129 , n18111 , n18364 );
xor ( n29130 , n29128 , n29129 );
xor ( n29131 , n29062 , n29125 );
and ( n29132 , n18112 , n18364 );
and ( n29133 , n29131 , n29132 );
xor ( n29134 , n29131 , n29132 );
xor ( n29135 , n29066 , n29123 );
and ( n29136 , n18113 , n18364 );
and ( n29137 , n29135 , n29136 );
xor ( n29138 , n29135 , n29136 );
xor ( n29139 , n29070 , n29121 );
and ( n29140 , n18114 , n18364 );
and ( n29141 , n29139 , n29140 );
xor ( n29142 , n29139 , n29140 );
xor ( n29143 , n29074 , n29119 );
and ( n29144 , n18115 , n18364 );
and ( n29145 , n29143 , n29144 );
xor ( n29146 , n29143 , n29144 );
xor ( n29147 , n29078 , n29117 );
and ( n29148 , n18116 , n18364 );
and ( n29149 , n29147 , n29148 );
xor ( n29150 , n29147 , n29148 );
xor ( n29151 , n29082 , n29115 );
and ( n29152 , n18117 , n18364 );
and ( n29153 , n29151 , n29152 );
xor ( n29154 , n29151 , n29152 );
xor ( n29155 , n29086 , n29113 );
and ( n29156 , n18118 , n18364 );
and ( n29157 , n29155 , n29156 );
xor ( n29158 , n29155 , n29156 );
xor ( n29159 , n29090 , n29111 );
and ( n29160 , n18119 , n18364 );
and ( n29161 , n29159 , n29160 );
xor ( n29162 , n29159 , n29160 );
xor ( n29163 , n29094 , n29109 );
and ( n29164 , n18120 , n18364 );
and ( n29165 , n29163 , n29164 );
xor ( n29166 , n29163 , n29164 );
xor ( n29167 , n29098 , n29107 );
and ( n29168 , n18121 , n18364 );
and ( n29169 , n29167 , n29168 );
xor ( n29170 , n29167 , n29168 );
xor ( n29171 , n29102 , n29105 );
and ( n29172 , n18122 , n18364 );
and ( n29173 , n29171 , n29172 );
and ( n29174 , n29170 , n29173 );
or ( n29175 , n29169 , n29174 );
and ( n29176 , n29166 , n29175 );
or ( n29177 , n29165 , n29176 );
and ( n29178 , n29162 , n29177 );
or ( n29179 , n29161 , n29178 );
and ( n29180 , n29158 , n29179 );
or ( n29181 , n29157 , n29180 );
and ( n29182 , n29154 , n29181 );
or ( n29183 , n29153 , n29182 );
and ( n29184 , n29150 , n29183 );
or ( n29185 , n29149 , n29184 );
and ( n29186 , n29146 , n29185 );
or ( n29187 , n29145 , n29186 );
and ( n29188 , n29142 , n29187 );
or ( n29189 , n29141 , n29188 );
and ( n29190 , n29138 , n29189 );
or ( n29191 , n29137 , n29190 );
and ( n29192 , n29134 , n29191 );
or ( n29193 , n29133 , n29192 );
xor ( n29194 , n29130 , n29193 );
and ( n29195 , n18112 , n18362 );
xor ( n29196 , n29194 , n29195 );
xor ( n29197 , n29134 , n29191 );
and ( n29198 , n18113 , n18362 );
and ( n29199 , n29197 , n29198 );
xor ( n29200 , n29197 , n29198 );
xor ( n29201 , n29138 , n29189 );
and ( n29202 , n18114 , n18362 );
and ( n29203 , n29201 , n29202 );
xor ( n29204 , n29201 , n29202 );
xor ( n29205 , n29142 , n29187 );
and ( n29206 , n18115 , n18362 );
and ( n29207 , n29205 , n29206 );
xor ( n29208 , n29205 , n29206 );
xor ( n29209 , n29146 , n29185 );
and ( n29210 , n18116 , n18362 );
and ( n29211 , n29209 , n29210 );
xor ( n29212 , n29209 , n29210 );
xor ( n29213 , n29150 , n29183 );
and ( n29214 , n18117 , n18362 );
and ( n29215 , n29213 , n29214 );
xor ( n29216 , n29213 , n29214 );
xor ( n29217 , n29154 , n29181 );
and ( n29218 , n18118 , n18362 );
and ( n29219 , n29217 , n29218 );
xor ( n29220 , n29217 , n29218 );
xor ( n29221 , n29158 , n29179 );
and ( n29222 , n18119 , n18362 );
and ( n29223 , n29221 , n29222 );
xor ( n29224 , n29221 , n29222 );
xor ( n29225 , n29162 , n29177 );
and ( n29226 , n18120 , n18362 );
and ( n29227 , n29225 , n29226 );
xor ( n29228 , n29225 , n29226 );
xor ( n29229 , n29166 , n29175 );
and ( n29230 , n18121 , n18362 );
and ( n29231 , n29229 , n29230 );
xor ( n29232 , n29229 , n29230 );
xor ( n29233 , n29170 , n29173 );
and ( n29234 , n18122 , n18362 );
and ( n29235 , n29233 , n29234 );
and ( n29236 , n29232 , n29235 );
or ( n29237 , n29231 , n29236 );
and ( n29238 , n29228 , n29237 );
or ( n29239 , n29227 , n29238 );
and ( n29240 , n29224 , n29239 );
or ( n29241 , n29223 , n29240 );
and ( n29242 , n29220 , n29241 );
or ( n29243 , n29219 , n29242 );
and ( n29244 , n29216 , n29243 );
or ( n29245 , n29215 , n29244 );
and ( n29246 , n29212 , n29245 );
or ( n29247 , n29211 , n29246 );
and ( n29248 , n29208 , n29247 );
or ( n29249 , n29207 , n29248 );
and ( n29250 , n29204 , n29249 );
or ( n29251 , n29203 , n29250 );
and ( n29252 , n29200 , n29251 );
or ( n29253 , n29199 , n29252 );
xor ( n29254 , n29196 , n29253 );
and ( n29255 , n18113 , n18360 );
xor ( n29256 , n29254 , n29255 );
xor ( n29257 , n29200 , n29251 );
and ( n29258 , n18114 , n18360 );
and ( n29259 , n29257 , n29258 );
xor ( n29260 , n29257 , n29258 );
xor ( n29261 , n29204 , n29249 );
and ( n29262 , n18115 , n18360 );
and ( n29263 , n29261 , n29262 );
xor ( n29264 , n29261 , n29262 );
xor ( n29265 , n29208 , n29247 );
and ( n29266 , n18116 , n18360 );
and ( n29267 , n29265 , n29266 );
xor ( n29268 , n29265 , n29266 );
xor ( n29269 , n29212 , n29245 );
and ( n29270 , n18117 , n18360 );
and ( n29271 , n29269 , n29270 );
xor ( n29272 , n29269 , n29270 );
xor ( n29273 , n29216 , n29243 );
and ( n29274 , n18118 , n18360 );
and ( n29275 , n29273 , n29274 );
xor ( n29276 , n29273 , n29274 );
xor ( n29277 , n29220 , n29241 );
and ( n29278 , n18119 , n18360 );
and ( n29279 , n29277 , n29278 );
xor ( n29280 , n29277 , n29278 );
xor ( n29281 , n29224 , n29239 );
and ( n29282 , n18120 , n18360 );
and ( n29283 , n29281 , n29282 );
xor ( n29284 , n29281 , n29282 );
xor ( n29285 , n29228 , n29237 );
and ( n29286 , n18121 , n18360 );
and ( n29287 , n29285 , n29286 );
xor ( n29288 , n29285 , n29286 );
xor ( n29289 , n29232 , n29235 );
and ( n29290 , n18122 , n18360 );
and ( n29291 , n29289 , n29290 );
and ( n29292 , n29288 , n29291 );
or ( n29293 , n29287 , n29292 );
and ( n29294 , n29284 , n29293 );
or ( n29295 , n29283 , n29294 );
and ( n29296 , n29280 , n29295 );
or ( n29297 , n29279 , n29296 );
and ( n29298 , n29276 , n29297 );
or ( n29299 , n29275 , n29298 );
and ( n29300 , n29272 , n29299 );
or ( n29301 , n29271 , n29300 );
and ( n29302 , n29268 , n29301 );
or ( n29303 , n29267 , n29302 );
and ( n29304 , n29264 , n29303 );
or ( n29305 , n29263 , n29304 );
and ( n29306 , n29260 , n29305 );
or ( n29307 , n29259 , n29306 );
xor ( n29308 , n29256 , n29307 );
and ( n29309 , n18114 , n18358 );
xor ( n29310 , n29308 , n29309 );
xor ( n29311 , n29260 , n29305 );
and ( n29312 , n18115 , n18358 );
and ( n29313 , n29311 , n29312 );
xor ( n29314 , n29311 , n29312 );
xor ( n29315 , n29264 , n29303 );
and ( n29316 , n18116 , n18358 );
and ( n29317 , n29315 , n29316 );
xor ( n29318 , n29315 , n29316 );
xor ( n29319 , n29268 , n29301 );
and ( n29320 , n18117 , n18358 );
and ( n29321 , n29319 , n29320 );
xor ( n29322 , n29319 , n29320 );
xor ( n29323 , n29272 , n29299 );
and ( n29324 , n18118 , n18358 );
and ( n29325 , n29323 , n29324 );
xor ( n29326 , n29323 , n29324 );
xor ( n29327 , n29276 , n29297 );
and ( n29328 , n18119 , n18358 );
and ( n29329 , n29327 , n29328 );
xor ( n29330 , n29327 , n29328 );
xor ( n29331 , n29280 , n29295 );
and ( n29332 , n18120 , n18358 );
and ( n29333 , n29331 , n29332 );
xor ( n29334 , n29331 , n29332 );
xor ( n29335 , n29284 , n29293 );
and ( n29336 , n18121 , n18358 );
and ( n29337 , n29335 , n29336 );
xor ( n29338 , n29335 , n29336 );
xor ( n29339 , n29288 , n29291 );
and ( n29340 , n18122 , n18358 );
and ( n29341 , n29339 , n29340 );
and ( n29342 , n29338 , n29341 );
or ( n29343 , n29337 , n29342 );
and ( n29344 , n29334 , n29343 );
or ( n29345 , n29333 , n29344 );
and ( n29346 , n29330 , n29345 );
or ( n29347 , n29329 , n29346 );
and ( n29348 , n29326 , n29347 );
or ( n29349 , n29325 , n29348 );
and ( n29350 , n29322 , n29349 );
or ( n29351 , n29321 , n29350 );
and ( n29352 , n29318 , n29351 );
or ( n29353 , n29317 , n29352 );
and ( n29354 , n29314 , n29353 );
or ( n29355 , n29313 , n29354 );
xor ( n29356 , n29310 , n29355 );
and ( n29357 , n18115 , n18356 );
xor ( n29358 , n29356 , n29357 );
xor ( n29359 , n29314 , n29353 );
and ( n29360 , n18116 , n18356 );
and ( n29361 , n29359 , n29360 );
xor ( n29362 , n29359 , n29360 );
xor ( n29363 , n29318 , n29351 );
and ( n29364 , n18117 , n18356 );
and ( n29365 , n29363 , n29364 );
xor ( n29366 , n29363 , n29364 );
xor ( n29367 , n29322 , n29349 );
and ( n29368 , n18118 , n18356 );
and ( n29369 , n29367 , n29368 );
xor ( n29370 , n29367 , n29368 );
xor ( n29371 , n29326 , n29347 );
and ( n29372 , n18119 , n18356 );
and ( n29373 , n29371 , n29372 );
xor ( n29374 , n29371 , n29372 );
xor ( n29375 , n29330 , n29345 );
and ( n29376 , n18120 , n18356 );
and ( n29377 , n29375 , n29376 );
xor ( n29378 , n29375 , n29376 );
xor ( n29379 , n29334 , n29343 );
and ( n29380 , n18121 , n18356 );
and ( n29381 , n29379 , n29380 );
xor ( n29382 , n29379 , n29380 );
xor ( n29383 , n29338 , n29341 );
and ( n29384 , n18122 , n18356 );
and ( n29385 , n29383 , n29384 );
and ( n29386 , n29382 , n29385 );
or ( n29387 , n29381 , n29386 );
and ( n29388 , n29378 , n29387 );
or ( n29389 , n29377 , n29388 );
and ( n29390 , n29374 , n29389 );
or ( n29391 , n29373 , n29390 );
and ( n29392 , n29370 , n29391 );
or ( n29393 , n29369 , n29392 );
and ( n29394 , n29366 , n29393 );
or ( n29395 , n29365 , n29394 );
and ( n29396 , n29362 , n29395 );
or ( n29397 , n29361 , n29396 );
xor ( n29398 , n29358 , n29397 );
and ( n29399 , n18116 , n18354 );
xor ( n29400 , n29398 , n29399 );
xor ( n29401 , n29362 , n29395 );
and ( n29402 , n18117 , n18354 );
and ( n29403 , n29401 , n29402 );
xor ( n29404 , n29401 , n29402 );
xor ( n29405 , n29366 , n29393 );
and ( n29406 , n18118 , n18354 );
and ( n29407 , n29405 , n29406 );
xor ( n29408 , n29405 , n29406 );
xor ( n29409 , n29370 , n29391 );
and ( n29410 , n18119 , n18354 );
and ( n29411 , n29409 , n29410 );
xor ( n29412 , n29409 , n29410 );
xor ( n29413 , n29374 , n29389 );
and ( n29414 , n18120 , n18354 );
and ( n29415 , n29413 , n29414 );
xor ( n29416 , n29413 , n29414 );
xor ( n29417 , n29378 , n29387 );
and ( n29418 , n18121 , n18354 );
and ( n29419 , n29417 , n29418 );
xor ( n29420 , n29417 , n29418 );
xor ( n29421 , n29382 , n29385 );
and ( n29422 , n18122 , n18354 );
and ( n29423 , n29421 , n29422 );
and ( n29424 , n29420 , n29423 );
or ( n29425 , n29419 , n29424 );
and ( n29426 , n29416 , n29425 );
or ( n29427 , n29415 , n29426 );
and ( n29428 , n29412 , n29427 );
or ( n29429 , n29411 , n29428 );
and ( n29430 , n29408 , n29429 );
or ( n29431 , n29407 , n29430 );
and ( n29432 , n29404 , n29431 );
or ( n29433 , n29403 , n29432 );
xor ( n29434 , n29400 , n29433 );
and ( n29435 , n18117 , n18352 );
xor ( n29436 , n29434 , n29435 );
xor ( n29437 , n29404 , n29431 );
and ( n29438 , n18118 , n18352 );
and ( n29439 , n29437 , n29438 );
xor ( n29440 , n29437 , n29438 );
xor ( n29441 , n29408 , n29429 );
and ( n29442 , n18119 , n18352 );
and ( n29443 , n29441 , n29442 );
xor ( n29444 , n29441 , n29442 );
xor ( n29445 , n29412 , n29427 );
and ( n29446 , n18120 , n18352 );
and ( n29447 , n29445 , n29446 );
xor ( n29448 , n29445 , n29446 );
xor ( n29449 , n29416 , n29425 );
and ( n29450 , n18121 , n18352 );
and ( n29451 , n29449 , n29450 );
xor ( n29452 , n29449 , n29450 );
xor ( n29453 , n29420 , n29423 );
and ( n29454 , n18122 , n18352 );
and ( n29455 , n29453 , n29454 );
and ( n29456 , n29452 , n29455 );
or ( n29457 , n29451 , n29456 );
and ( n29458 , n29448 , n29457 );
or ( n29459 , n29447 , n29458 );
and ( n29460 , n29444 , n29459 );
or ( n29461 , n29443 , n29460 );
and ( n29462 , n29440 , n29461 );
or ( n29463 , n29439 , n29462 );
xor ( n29464 , n29436 , n29463 );
and ( n29465 , n18118 , n18350 );
xor ( n29466 , n29464 , n29465 );
xor ( n29467 , n29440 , n29461 );
and ( n29468 , n18119 , n18350 );
and ( n29469 , n29467 , n29468 );
xor ( n29470 , n29467 , n29468 );
xor ( n29471 , n29444 , n29459 );
and ( n29472 , n18120 , n18350 );
and ( n29473 , n29471 , n29472 );
xor ( n29474 , n29471 , n29472 );
xor ( n29475 , n29448 , n29457 );
and ( n29476 , n18121 , n18350 );
and ( n29477 , n29475 , n29476 );
xor ( n29478 , n29475 , n29476 );
xor ( n29479 , n29452 , n29455 );
and ( n29480 , n18122 , n18350 );
and ( n29481 , n29479 , n29480 );
and ( n29482 , n29478 , n29481 );
or ( n29483 , n29477 , n29482 );
and ( n29484 , n29474 , n29483 );
or ( n29485 , n29473 , n29484 );
and ( n29486 , n29470 , n29485 );
or ( n29487 , n29469 , n29486 );
xor ( n29488 , n29466 , n29487 );
and ( n29489 , n18119 , n18348 );
xor ( n29490 , n29488 , n29489 );
xor ( n29491 , n29470 , n29485 );
and ( n29492 , n18120 , n18348 );
and ( n29493 , n29491 , n29492 );
xor ( n29494 , n29491 , n29492 );
xor ( n29495 , n29474 , n29483 );
and ( n29496 , n18121 , n18348 );
and ( n29497 , n29495 , n29496 );
xor ( n29498 , n29495 , n29496 );
xor ( n29499 , n29478 , n29481 );
and ( n29500 , n18122 , n18348 );
and ( n29501 , n29499 , n29500 );
and ( n29502 , n29498 , n29501 );
or ( n29503 , n29497 , n29502 );
and ( n29504 , n29494 , n29503 );
or ( n29505 , n29493 , n29504 );
xor ( n29506 , n29490 , n29505 );
and ( n29507 , n18120 , n18346 );
xor ( n29508 , n29506 , n29507 );
xor ( n29509 , n29494 , n29503 );
and ( n29510 , n18121 , n18346 );
and ( n29511 , n29509 , n29510 );
xor ( n29512 , n29509 , n29510 );
xor ( n29513 , n29498 , n29501 );
and ( n29514 , n18122 , n18346 );
and ( n29515 , n29513 , n29514 );
and ( n29516 , n29512 , n29515 );
or ( n29517 , n29511 , n29516 );
xor ( n29518 , n29508 , n29517 );
and ( n29519 , n18121 , n18344 );
xor ( n29520 , n29518 , n29519 );
xor ( n29521 , n29512 , n29515 );
and ( n29522 , n18122 , n18344 );
and ( n29523 , n29521 , n29522 );
xor ( n29524 , n29520 , n29523 );
and ( n29525 , n18122 , n18342 );
xor ( n29526 , n29524 , n29525 );
buf ( n29527 , n29526 );
xor ( n29528 , n29521 , n29522 );
buf ( n29529 , n29528 );
xor ( n29530 , n29513 , n29514 );
buf ( n29531 , n29530 );
xor ( n29532 , n29499 , n29500 );
buf ( n29533 , n29532 );
xor ( n29534 , n29479 , n29480 );
buf ( n29535 , n29534 );
xor ( n29536 , n29453 , n29454 );
buf ( n29537 , n29536 );
xor ( n29538 , n29421 , n29422 );
buf ( n29539 , n29538 );
xor ( n29540 , n29383 , n29384 );
buf ( n29541 , n29540 );
xor ( n29542 , n29339 , n29340 );
buf ( n29543 , n29542 );
xor ( n29544 , n29289 , n29290 );
buf ( n29545 , n29544 );
xor ( n29546 , n29233 , n29234 );
buf ( n29547 , n29546 );
xor ( n29548 , n29171 , n29172 );
buf ( n29549 , n29548 );
xor ( n29550 , n29103 , n29104 );
buf ( n29551 , n29550 );
xor ( n29552 , n29029 , n29030 );
buf ( n29553 , n29552 );
xor ( n29554 , n28949 , n28950 );
buf ( n29555 , n29554 );
xor ( n29556 , n28863 , n28864 );
buf ( n29557 , n29556 );
xor ( n29558 , n28772 , n28773 );
buf ( n29559 , n29558 );
xor ( n29560 , n28680 , n28681 );
buf ( n29561 , n29560 );
xor ( n29562 , n28588 , n28589 );
buf ( n29563 , n29562 );
xor ( n29564 , n28496 , n28497 );
buf ( n29565 , n29564 );
xor ( n29566 , n28404 , n28405 );
buf ( n29567 , n29566 );
xor ( n29568 , n28312 , n28313 );
buf ( n29569 , n29568 );
xor ( n29570 , n28220 , n28221 );
buf ( n29571 , n29570 );
xor ( n29572 , n28128 , n28129 );
buf ( n29573 , n29572 );
xor ( n29574 , n28036 , n28037 );
buf ( n29575 , n29574 );
xor ( n29576 , n27944 , n27945 );
buf ( n29577 , n29576 );
xor ( n29578 , n27852 , n27853 );
buf ( n29579 , n29578 );
xor ( n29580 , n27760 , n27761 );
buf ( n29581 , n29580 );
xor ( n29582 , n27668 , n27669 );
buf ( n29583 , n29582 );
xor ( n29584 , n27576 , n27577 );
buf ( n29585 , n29584 );
xor ( n29586 , n27484 , n27485 );
buf ( n29587 , n29586 );
xor ( n29588 , n27392 , n27393 );
buf ( n29589 , n29588 );
xor ( n29590 , n27300 , n27301 );
buf ( n29591 , n29590 );
xor ( n29592 , n27208 , n27209 );
buf ( n29593 , n29592 );
xor ( n29594 , n27116 , n27117 );
buf ( n29595 , n29594 );
xor ( n29596 , n27024 , n27025 );
buf ( n29597 , n29596 );
xor ( n29598 , n26932 , n26933 );
buf ( n29599 , n29598 );
xor ( n29600 , n26840 , n26841 );
buf ( n29601 , n29600 );
xor ( n29602 , n26748 , n26749 );
buf ( n29603 , n29602 );
xor ( n29604 , n26656 , n26657 );
buf ( n29605 , n29604 );
xor ( n29606 , n26564 , n26565 );
buf ( n29607 , n29606 );
xor ( n29608 , n26472 , n26473 );
buf ( n29609 , n29608 );
xor ( n29610 , n26380 , n26381 );
buf ( n29611 , n29610 );
xor ( n29612 , n26288 , n26289 );
buf ( n29613 , n29612 );
xor ( n29614 , n26196 , n26197 );
buf ( n29615 , n29614 );
xor ( n29616 , n26104 , n26105 );
buf ( n29617 , n29616 );
xor ( n29618 , n26012 , n26013 );
buf ( n29619 , n29618 );
xor ( n29620 , n25920 , n25921 );
buf ( n29621 , n29620 );
xor ( n29622 , n25828 , n25829 );
buf ( n29623 , n29622 );
xor ( n29624 , n25736 , n25737 );
buf ( n29625 , n29624 );
xor ( n29626 , n25644 , n25645 );
buf ( n29627 , n29626 );
xor ( n29628 , n25552 , n25553 );
buf ( n29629 , n29628 );
xor ( n29630 , n25460 , n25461 );
buf ( n29631 , n29630 );
xor ( n29632 , n25368 , n25369 );
buf ( n29633 , n29632 );
xor ( n29634 , n25276 , n25277 );
buf ( n29635 , n29634 );
xor ( n29636 , n25184 , n25185 );
buf ( n29637 , n29636 );
xor ( n29638 , n25092 , n25093 );
buf ( n29639 , n29638 );
xor ( n29640 , n25000 , n25001 );
buf ( n29641 , n29640 );
xor ( n29642 , n24908 , n24909 );
buf ( n29643 , n29642 );
xor ( n29644 , n24816 , n24817 );
buf ( n29645 , n29644 );
xor ( n29646 , n24724 , n24725 );
buf ( n29647 , n29646 );
xor ( n29648 , n24632 , n24633 );
buf ( n29649 , n29648 );
xor ( n29650 , n24540 , n24541 );
buf ( n29651 , n29650 );
xor ( n29652 , n24448 , n24449 );
buf ( n29653 , n29652 );
xor ( n29654 , n24356 , n24357 );
buf ( n29655 , n29654 );
xor ( n29656 , n24264 , n24265 );
buf ( n29657 , n29656 );
xor ( n29658 , n24172 , n24173 );
buf ( n29659 , n29658 );
xor ( n29660 , n24080 , n24081 );
buf ( n29661 , n29660 );
xor ( n29662 , n23988 , n23989 );
buf ( n29663 , n29662 );
xor ( n29664 , n23896 , n23897 );
buf ( n29665 , n29664 );
xor ( n29666 , n23804 , n23805 );
buf ( n29667 , n29666 );
xor ( n29668 , n23712 , n23713 );
buf ( n29669 , n29668 );
xor ( n29670 , n23620 , n23621 );
buf ( n29671 , n29670 );
xor ( n29672 , n23528 , n23529 );
buf ( n29673 , n29672 );
xor ( n29674 , n23436 , n23437 );
buf ( n29675 , n29674 );
xor ( n29676 , n23344 , n23345 );
buf ( n29677 , n29676 );
xor ( n29678 , n23252 , n23253 );
buf ( n29679 , n29678 );
xor ( n29680 , n23160 , n23161 );
buf ( n29681 , n29680 );
xor ( n29682 , n23068 , n23069 );
buf ( n29683 , n29682 );
xor ( n29684 , n22976 , n22977 );
buf ( n29685 , n29684 );
xor ( n29686 , n22884 , n22885 );
buf ( n29687 , n29686 );
xor ( n29688 , n22792 , n22793 );
buf ( n29689 , n29688 );
xor ( n29690 , n22700 , n22701 );
buf ( n29691 , n29690 );
xor ( n29692 , n22608 , n22609 );
buf ( n29693 , n29692 );
xor ( n29694 , n22516 , n22517 );
buf ( n29695 , n29694 );
xor ( n29696 , n22424 , n22425 );
buf ( n29697 , n29696 );
xor ( n29698 , n22332 , n22333 );
buf ( n29699 , n29698 );
xor ( n29700 , n22240 , n22241 );
buf ( n29701 , n29700 );
xor ( n29702 , n22148 , n22149 );
buf ( n29703 , n29702 );
xor ( n29704 , n22056 , n22057 );
buf ( n29705 , n29704 );
xor ( n29706 , n21964 , n21965 );
buf ( n29707 , n29706 );
xor ( n29708 , n21872 , n21873 );
buf ( n29709 , n29708 );
xor ( n29710 , n21780 , n21781 );
buf ( n29711 , n29710 );
xor ( n29712 , n21688 , n21689 );
buf ( n29713 , n29712 );
xor ( n29714 , n21596 , n21597 );
buf ( n29715 , n29714 );
xor ( n29716 , n21504 , n21505 );
buf ( n29717 , n29716 );
xor ( n29718 , n21412 , n21413 );
buf ( n29719 , n29718 );
xor ( n29720 , n21320 , n21321 );
buf ( n29721 , n29720 );
xor ( n29722 , n21228 , n21229 );
buf ( n29723 , n29722 );
xor ( n29724 , n21136 , n21137 );
buf ( n29725 , n29724 );
xor ( n29726 , n21044 , n21045 );
buf ( n29727 , n29726 );
xor ( n29728 , n20952 , n20953 );
buf ( n29729 , n29728 );
xor ( n29730 , n20860 , n20861 );
buf ( n29731 , n29730 );
xor ( n29732 , n20768 , n20769 );
buf ( n29733 , n29732 );
xor ( n29734 , n20676 , n20677 );
buf ( n29735 , n29734 );
xor ( n29736 , n20584 , n20585 );
buf ( n29737 , n29736 );
xor ( n29738 , n20492 , n20493 );
buf ( n29739 , n29738 );
xor ( n29740 , n20400 , n20401 );
buf ( n29741 , n29740 );
xor ( n29742 , n20308 , n20309 );
buf ( n29743 , n29742 );
xor ( n29744 , n20216 , n20217 );
buf ( n29745 , n29744 );
xor ( n29746 , n20124 , n20125 );
buf ( n29747 , n29746 );
xor ( n29748 , n20032 , n20033 );
buf ( n29749 , n29748 );
xor ( n29750 , n19940 , n19941 );
buf ( n29751 , n29750 );
xor ( n29752 , n19848 , n19849 );
buf ( n29753 , n29752 );
xor ( n29754 , n19756 , n19757 );
buf ( n29755 , n29754 );
xor ( n29756 , n19664 , n19665 );
buf ( n29757 , n29756 );
xor ( n29758 , n19572 , n19573 );
buf ( n29759 , n29758 );
xor ( n29760 , n19480 , n19481 );
buf ( n29761 , n29760 );
xor ( n29762 , n19388 , n19389 );
buf ( n29763 , n29762 );
xor ( n29764 , n19296 , n19297 );
buf ( n29765 , n29764 );
xor ( n29766 , n19204 , n19205 );
buf ( n29767 , n29766 );
xor ( n29768 , n19112 , n19113 );
buf ( n29769 , n29768 );
xor ( n29770 , n19020 , n19021 );
buf ( n29771 , n29770 );
xor ( n29772 , n18928 , n18929 );
buf ( n29773 , n29772 );
xor ( n29774 , n18836 , n18837 );
buf ( n29775 , n29774 );
xor ( n29776 , n18744 , n18745 );
buf ( n29777 , n29776 );
and ( n29778 , n18122 , n18656 );
buf ( n29779 , n29778 );
buf ( n29780 , n29779 );
buf ( n29781 , n29527 );
buf ( n29782 , n18106 );
and ( n29783 , n29781 , n29782 );
buf ( n29784 , n29529 );
buf ( n29785 , n18104 );
and ( n29786 , n29784 , n29785 );
xor ( n29787 , n29783 , n29786 );
and ( n29788 , n29784 , n29782 );
buf ( n29789 , n29531 );
and ( n29790 , n29789 , n29785 );
and ( n29791 , n29788 , n29790 );
xor ( n29792 , n29788 , n29790 );
and ( n29793 , n29789 , n29782 );
buf ( n29794 , n29533 );
and ( n29795 , n29794 , n29785 );
and ( n29796 , n29793 , n29795 );
xor ( n29797 , n29793 , n29795 );
and ( n29798 , n29794 , n29782 );
buf ( n29799 , n29535 );
and ( n29800 , n29799 , n29785 );
and ( n29801 , n29798 , n29800 );
xor ( n29802 , n29798 , n29800 );
and ( n29803 , n29799 , n29782 );
buf ( n29804 , n29537 );
and ( n29805 , n29804 , n29785 );
and ( n29806 , n29803 , n29805 );
xor ( n29807 , n29803 , n29805 );
and ( n29808 , n29804 , n29782 );
buf ( n29809 , n29539 );
and ( n29810 , n29809 , n29785 );
and ( n29811 , n29808 , n29810 );
xor ( n29812 , n29808 , n29810 );
and ( n29813 , n29809 , n29782 );
buf ( n29814 , n29541 );
and ( n29815 , n29814 , n29785 );
and ( n29816 , n29813 , n29815 );
xor ( n29817 , n29813 , n29815 );
and ( n29818 , n29814 , n29782 );
buf ( n29819 , n29543 );
and ( n29820 , n29819 , n29785 );
and ( n29821 , n29818 , n29820 );
xor ( n29822 , n29818 , n29820 );
and ( n29823 , n29819 , n29782 );
buf ( n29824 , n29545 );
and ( n29825 , n29824 , n29785 );
and ( n29826 , n29823 , n29825 );
xor ( n29827 , n29823 , n29825 );
and ( n29828 , n29824 , n29782 );
buf ( n29829 , n29547 );
and ( n29830 , n29829 , n29785 );
and ( n29831 , n29828 , n29830 );
xor ( n29832 , n29828 , n29830 );
and ( n29833 , n29829 , n29782 );
buf ( n29834 , n29549 );
and ( n29835 , n29834 , n29785 );
and ( n29836 , n29833 , n29835 );
xor ( n29837 , n29833 , n29835 );
and ( n29838 , n29834 , n29782 );
buf ( n29839 , n29551 );
and ( n29840 , n29839 , n29785 );
and ( n29841 , n29838 , n29840 );
xor ( n29842 , n29838 , n29840 );
and ( n29843 , n29839 , n29782 );
buf ( n29844 , n29553 );
and ( n29845 , n29844 , n29785 );
and ( n29846 , n29843 , n29845 );
xor ( n29847 , n29843 , n29845 );
and ( n29848 , n29844 , n29782 );
buf ( n29849 , n29555 );
and ( n29850 , n29849 , n29785 );
and ( n29851 , n29848 , n29850 );
xor ( n29852 , n29848 , n29850 );
and ( n29853 , n29849 , n29782 );
buf ( n29854 , n29557 );
and ( n29855 , n29854 , n29785 );
and ( n29856 , n29853 , n29855 );
xor ( n29857 , n29853 , n29855 );
and ( n29858 , n29854 , n29782 );
buf ( n29859 , n29559 );
and ( n29860 , n29859 , n29785 );
and ( n29861 , n29858 , n29860 );
xor ( n29862 , n29858 , n29860 );
and ( n29863 , n29859 , n29782 );
buf ( n29864 , n29561 );
and ( n29865 , n29864 , n29785 );
and ( n29866 , n29863 , n29865 );
xor ( n29867 , n29863 , n29865 );
and ( n29868 , n29864 , n29782 );
buf ( n29869 , n29563 );
and ( n29870 , n29869 , n29785 );
and ( n29871 , n29868 , n29870 );
xor ( n29872 , n29868 , n29870 );
and ( n29873 , n29869 , n29782 );
buf ( n29874 , n29565 );
and ( n29875 , n29874 , n29785 );
and ( n29876 , n29873 , n29875 );
xor ( n29877 , n29873 , n29875 );
and ( n29878 , n29874 , n29782 );
buf ( n29879 , n29567 );
and ( n29880 , n29879 , n29785 );
and ( n29881 , n29878 , n29880 );
xor ( n29882 , n29878 , n29880 );
and ( n29883 , n29879 , n29782 );
buf ( n29884 , n29569 );
and ( n29885 , n29884 , n29785 );
and ( n29886 , n29883 , n29885 );
xor ( n29887 , n29883 , n29885 );
and ( n29888 , n29884 , n29782 );
buf ( n29889 , n29571 );
and ( n29890 , n29889 , n29785 );
and ( n29891 , n29888 , n29890 );
xor ( n29892 , n29888 , n29890 );
and ( n29893 , n29889 , n29782 );
buf ( n29894 , n29573 );
and ( n29895 , n29894 , n29785 );
and ( n29896 , n29893 , n29895 );
xor ( n29897 , n29893 , n29895 );
and ( n29898 , n29894 , n29782 );
buf ( n29899 , n29575 );
and ( n29900 , n29899 , n29785 );
and ( n29901 , n29898 , n29900 );
xor ( n29902 , n29898 , n29900 );
and ( n29903 , n29899 , n29782 );
buf ( n29904 , n29577 );
and ( n29905 , n29904 , n29785 );
and ( n29906 , n29903 , n29905 );
xor ( n29907 , n29903 , n29905 );
and ( n29908 , n29904 , n29782 );
buf ( n29909 , n29579 );
and ( n29910 , n29909 , n29785 );
and ( n29911 , n29908 , n29910 );
xor ( n29912 , n29908 , n29910 );
and ( n29913 , n29909 , n29782 );
buf ( n29914 , n29581 );
and ( n29915 , n29914 , n29785 );
and ( n29916 , n29913 , n29915 );
xor ( n29917 , n29913 , n29915 );
and ( n29918 , n29914 , n29782 );
buf ( n29919 , n29583 );
and ( n29920 , n29919 , n29785 );
and ( n29921 , n29918 , n29920 );
xor ( n29922 , n29918 , n29920 );
and ( n29923 , n29919 , n29782 );
buf ( n29924 , n29585 );
and ( n29925 , n29924 , n29785 );
and ( n29926 , n29923 , n29925 );
xor ( n29927 , n29923 , n29925 );
and ( n29928 , n29924 , n29782 );
buf ( n29929 , n29587 );
and ( n29930 , n29929 , n29785 );
and ( n29931 , n29928 , n29930 );
xor ( n29932 , n29928 , n29930 );
and ( n29933 , n29929 , n29782 );
buf ( n29934 , n29589 );
and ( n29935 , n29934 , n29785 );
and ( n29936 , n29933 , n29935 );
xor ( n29937 , n29933 , n29935 );
and ( n29938 , n29934 , n29782 );
buf ( n29939 , n29591 );
and ( n29940 , n29939 , n29785 );
and ( n29941 , n29938 , n29940 );
xor ( n29942 , n29938 , n29940 );
and ( n29943 , n29939 , n29782 );
buf ( n29944 , n29593 );
and ( n29945 , n29944 , n29785 );
and ( n29946 , n29943 , n29945 );
xor ( n29947 , n29943 , n29945 );
and ( n29948 , n29944 , n29782 );
buf ( n29949 , n29595 );
and ( n29950 , n29949 , n29785 );
and ( n29951 , n29948 , n29950 );
xor ( n29952 , n29948 , n29950 );
and ( n29953 , n29949 , n29782 );
buf ( n29954 , n29597 );
and ( n29955 , n29954 , n29785 );
and ( n29956 , n29953 , n29955 );
xor ( n29957 , n29953 , n29955 );
and ( n29958 , n29954 , n29782 );
buf ( n29959 , n29599 );
and ( n29960 , n29959 , n29785 );
and ( n29961 , n29958 , n29960 );
xor ( n29962 , n29958 , n29960 );
and ( n29963 , n29959 , n29782 );
buf ( n29964 , n29601 );
and ( n29965 , n29964 , n29785 );
and ( n29966 , n29963 , n29965 );
xor ( n29967 , n29963 , n29965 );
and ( n29968 , n29964 , n29782 );
buf ( n29969 , n29603 );
and ( n29970 , n29969 , n29785 );
and ( n29971 , n29968 , n29970 );
xor ( n29972 , n29968 , n29970 );
and ( n29973 , n29969 , n29782 );
buf ( n29974 , n29605 );
and ( n29975 , n29974 , n29785 );
and ( n29976 , n29973 , n29975 );
xor ( n29977 , n29973 , n29975 );
and ( n29978 , n29974 , n29782 );
buf ( n29979 , n29607 );
and ( n29980 , n29979 , n29785 );
and ( n29981 , n29978 , n29980 );
xor ( n29982 , n29978 , n29980 );
and ( n29983 , n29979 , n29782 );
buf ( n29984 , n29609 );
and ( n29985 , n29984 , n29785 );
and ( n29986 , n29983 , n29985 );
xor ( n29987 , n29983 , n29985 );
and ( n29988 , n29984 , n29782 );
buf ( n29989 , n29611 );
and ( n29990 , n29989 , n29785 );
and ( n29991 , n29988 , n29990 );
xor ( n29992 , n29988 , n29990 );
and ( n29993 , n29989 , n29782 );
buf ( n29994 , n29613 );
and ( n29995 , n29994 , n29785 );
and ( n29996 , n29993 , n29995 );
xor ( n29997 , n29993 , n29995 );
and ( n29998 , n29994 , n29782 );
buf ( n29999 , n29615 );
and ( n30000 , n29999 , n29785 );
and ( n30001 , n29998 , n30000 );
xor ( n30002 , n29998 , n30000 );
and ( n30003 , n29999 , n29782 );
buf ( n30004 , n29617 );
and ( n30005 , n30004 , n29785 );
and ( n30006 , n30003 , n30005 );
xor ( n30007 , n30003 , n30005 );
and ( n30008 , n30004 , n29782 );
buf ( n30009 , n29619 );
and ( n30010 , n30009 , n29785 );
and ( n30011 , n30008 , n30010 );
xor ( n30012 , n30008 , n30010 );
and ( n30013 , n30009 , n29782 );
buf ( n30014 , n29621 );
and ( n30015 , n30014 , n29785 );
and ( n30016 , n30013 , n30015 );
xor ( n30017 , n30013 , n30015 );
and ( n30018 , n30014 , n29782 );
buf ( n30019 , n29623 );
and ( n30020 , n30019 , n29785 );
and ( n30021 , n30018 , n30020 );
xor ( n30022 , n30018 , n30020 );
and ( n30023 , n30019 , n29782 );
buf ( n30024 , n29625 );
and ( n30025 , n30024 , n29785 );
and ( n30026 , n30023 , n30025 );
xor ( n30027 , n30023 , n30025 );
and ( n30028 , n30024 , n29782 );
buf ( n30029 , n29627 );
and ( n30030 , n30029 , n29785 );
and ( n30031 , n30028 , n30030 );
xor ( n30032 , n30028 , n30030 );
and ( n30033 , n30029 , n29782 );
buf ( n30034 , n29629 );
and ( n30035 , n30034 , n29785 );
and ( n30036 , n30033 , n30035 );
xor ( n30037 , n30033 , n30035 );
and ( n30038 , n30034 , n29782 );
buf ( n30039 , n29631 );
and ( n30040 , n30039 , n29785 );
and ( n30041 , n30038 , n30040 );
xor ( n30042 , n30038 , n30040 );
and ( n30043 , n30039 , n29782 );
buf ( n30044 , n29633 );
and ( n30045 , n30044 , n29785 );
and ( n30046 , n30043 , n30045 );
xor ( n30047 , n30043 , n30045 );
and ( n30048 , n30044 , n29782 );
buf ( n30049 , n29635 );
and ( n30050 , n30049 , n29785 );
and ( n30051 , n30048 , n30050 );
xor ( n30052 , n30048 , n30050 );
and ( n30053 , n30049 , n29782 );
buf ( n30054 , n29637 );
and ( n30055 , n30054 , n29785 );
and ( n30056 , n30053 , n30055 );
xor ( n30057 , n30053 , n30055 );
and ( n30058 , n30054 , n29782 );
buf ( n30059 , n29639 );
and ( n30060 , n30059 , n29785 );
and ( n30061 , n30058 , n30060 );
xor ( n30062 , n30058 , n30060 );
and ( n30063 , n30059 , n29782 );
buf ( n30064 , n29641 );
and ( n30065 , n30064 , n29785 );
and ( n30066 , n30063 , n30065 );
xor ( n30067 , n30063 , n30065 );
and ( n30068 , n30064 , n29782 );
buf ( n30069 , n29643 );
and ( n30070 , n30069 , n29785 );
and ( n30071 , n30068 , n30070 );
xor ( n30072 , n30068 , n30070 );
and ( n30073 , n30069 , n29782 );
buf ( n30074 , n29645 );
and ( n30075 , n30074 , n29785 );
and ( n30076 , n30073 , n30075 );
xor ( n30077 , n30073 , n30075 );
and ( n30078 , n30074 , n29782 );
buf ( n30079 , n29647 );
and ( n30080 , n30079 , n29785 );
and ( n30081 , n30078 , n30080 );
xor ( n30082 , n30078 , n30080 );
and ( n30083 , n30079 , n29782 );
buf ( n30084 , n29649 );
and ( n30085 , n30084 , n29785 );
and ( n30086 , n30083 , n30085 );
xor ( n30087 , n30083 , n30085 );
and ( n30088 , n30084 , n29782 );
buf ( n30089 , n29651 );
and ( n30090 , n30089 , n29785 );
and ( n30091 , n30088 , n30090 );
xor ( n30092 , n30088 , n30090 );
and ( n30093 , n30089 , n29782 );
buf ( n30094 , n29653 );
and ( n30095 , n30094 , n29785 );
and ( n30096 , n30093 , n30095 );
xor ( n30097 , n30093 , n30095 );
and ( n30098 , n30094 , n29782 );
buf ( n30099 , n29655 );
and ( n30100 , n30099 , n29785 );
and ( n30101 , n30098 , n30100 );
xor ( n30102 , n30098 , n30100 );
and ( n30103 , n30099 , n29782 );
buf ( n30104 , n29657 );
and ( n30105 , n30104 , n29785 );
and ( n30106 , n30103 , n30105 );
xor ( n30107 , n30103 , n30105 );
and ( n30108 , n30104 , n29782 );
buf ( n30109 , n29659 );
and ( n30110 , n30109 , n29785 );
and ( n30111 , n30108 , n30110 );
xor ( n30112 , n30108 , n30110 );
and ( n30113 , n30109 , n29782 );
buf ( n30114 , n29661 );
and ( n30115 , n30114 , n29785 );
and ( n30116 , n30113 , n30115 );
xor ( n30117 , n30113 , n30115 );
and ( n30118 , n30114 , n29782 );
buf ( n30119 , n29663 );
and ( n30120 , n30119 , n29785 );
and ( n30121 , n30118 , n30120 );
xor ( n30122 , n30118 , n30120 );
and ( n30123 , n30119 , n29782 );
buf ( n30124 , n29665 );
and ( n30125 , n30124 , n29785 );
and ( n30126 , n30123 , n30125 );
xor ( n30127 , n30123 , n30125 );
and ( n30128 , n30124 , n29782 );
buf ( n30129 , n29667 );
and ( n30130 , n30129 , n29785 );
and ( n30131 , n30128 , n30130 );
xor ( n30132 , n30128 , n30130 );
and ( n30133 , n30129 , n29782 );
buf ( n30134 , n29669 );
and ( n30135 , n30134 , n29785 );
and ( n30136 , n30133 , n30135 );
xor ( n30137 , n30133 , n30135 );
and ( n30138 , n30134 , n29782 );
buf ( n30139 , n29671 );
and ( n30140 , n30139 , n29785 );
and ( n30141 , n30138 , n30140 );
xor ( n30142 , n30138 , n30140 );
and ( n30143 , n30139 , n29782 );
buf ( n30144 , n29673 );
and ( n30145 , n30144 , n29785 );
and ( n30146 , n30143 , n30145 );
xor ( n30147 , n30143 , n30145 );
and ( n30148 , n30144 , n29782 );
buf ( n30149 , n29675 );
and ( n30150 , n30149 , n29785 );
and ( n30151 , n30148 , n30150 );
xor ( n30152 , n30148 , n30150 );
and ( n30153 , n30149 , n29782 );
buf ( n30154 , n29677 );
and ( n30155 , n30154 , n29785 );
and ( n30156 , n30153 , n30155 );
xor ( n30157 , n30153 , n30155 );
and ( n30158 , n30154 , n29782 );
buf ( n30159 , n29679 );
and ( n30160 , n30159 , n29785 );
and ( n30161 , n30158 , n30160 );
xor ( n30162 , n30158 , n30160 );
and ( n30163 , n30159 , n29782 );
buf ( n30164 , n29681 );
and ( n30165 , n30164 , n29785 );
and ( n30166 , n30163 , n30165 );
xor ( n30167 , n30163 , n30165 );
and ( n30168 , n30164 , n29782 );
buf ( n30169 , n29683 );
and ( n30170 , n30169 , n29785 );
and ( n30171 , n30168 , n30170 );
xor ( n30172 , n30168 , n30170 );
and ( n30173 , n30169 , n29782 );
buf ( n30174 , n29685 );
and ( n30175 , n30174 , n29785 );
and ( n30176 , n30173 , n30175 );
xor ( n30177 , n30173 , n30175 );
and ( n30178 , n30174 , n29782 );
buf ( n30179 , n29687 );
and ( n30180 , n30179 , n29785 );
and ( n30181 , n30178 , n30180 );
xor ( n30182 , n30178 , n30180 );
and ( n30183 , n30179 , n29782 );
buf ( n30184 , n29689 );
and ( n30185 , n30184 , n29785 );
and ( n30186 , n30183 , n30185 );
xor ( n30187 , n30183 , n30185 );
and ( n30188 , n30184 , n29782 );
buf ( n30189 , n29691 );
and ( n30190 , n30189 , n29785 );
and ( n30191 , n30188 , n30190 );
xor ( n30192 , n30188 , n30190 );
and ( n30193 , n30189 , n29782 );
buf ( n30194 , n29693 );
and ( n30195 , n30194 , n29785 );
and ( n30196 , n30193 , n30195 );
xor ( n30197 , n30193 , n30195 );
and ( n30198 , n30194 , n29782 );
buf ( n30199 , n29695 );
and ( n30200 , n30199 , n29785 );
and ( n30201 , n30198 , n30200 );
xor ( n30202 , n30198 , n30200 );
and ( n30203 , n30199 , n29782 );
buf ( n30204 , n29697 );
and ( n30205 , n30204 , n29785 );
and ( n30206 , n30203 , n30205 );
xor ( n30207 , n30203 , n30205 );
and ( n30208 , n30204 , n29782 );
buf ( n30209 , n29699 );
and ( n30210 , n30209 , n29785 );
and ( n30211 , n30208 , n30210 );
xor ( n30212 , n30208 , n30210 );
and ( n30213 , n30209 , n29782 );
buf ( n30214 , n29701 );
and ( n30215 , n30214 , n29785 );
and ( n30216 , n30213 , n30215 );
xor ( n30217 , n30213 , n30215 );
and ( n30218 , n30214 , n29782 );
buf ( n30219 , n29703 );
and ( n30220 , n30219 , n29785 );
and ( n30221 , n30218 , n30220 );
xor ( n30222 , n30218 , n30220 );
and ( n30223 , n30219 , n29782 );
buf ( n30224 , n29705 );
and ( n30225 , n30224 , n29785 );
and ( n30226 , n30223 , n30225 );
xor ( n30227 , n30223 , n30225 );
and ( n30228 , n30224 , n29782 );
buf ( n30229 , n29707 );
and ( n30230 , n30229 , n29785 );
and ( n30231 , n30228 , n30230 );
xor ( n30232 , n30228 , n30230 );
and ( n30233 , n30229 , n29782 );
buf ( n30234 , n29709 );
and ( n30235 , n30234 , n29785 );
and ( n30236 , n30233 , n30235 );
xor ( n30237 , n30233 , n30235 );
and ( n30238 , n30234 , n29782 );
buf ( n30239 , n29711 );
and ( n30240 , n30239 , n29785 );
and ( n30241 , n30238 , n30240 );
xor ( n30242 , n30238 , n30240 );
and ( n30243 , n30239 , n29782 );
buf ( n30244 , n29713 );
and ( n30245 , n30244 , n29785 );
and ( n30246 , n30243 , n30245 );
xor ( n30247 , n30243 , n30245 );
and ( n30248 , n30244 , n29782 );
buf ( n30249 , n29715 );
and ( n30250 , n30249 , n29785 );
and ( n30251 , n30248 , n30250 );
xor ( n30252 , n30248 , n30250 );
and ( n30253 , n30249 , n29782 );
buf ( n30254 , n29717 );
and ( n30255 , n30254 , n29785 );
and ( n30256 , n30253 , n30255 );
xor ( n30257 , n30253 , n30255 );
and ( n30258 , n30254 , n29782 );
buf ( n30259 , n29719 );
and ( n30260 , n30259 , n29785 );
and ( n30261 , n30258 , n30260 );
xor ( n30262 , n30258 , n30260 );
and ( n30263 , n30259 , n29782 );
buf ( n30264 , n29721 );
and ( n30265 , n30264 , n29785 );
and ( n30266 , n30263 , n30265 );
xor ( n30267 , n30263 , n30265 );
and ( n30268 , n30264 , n29782 );
buf ( n30269 , n29723 );
and ( n30270 , n30269 , n29785 );
and ( n30271 , n30268 , n30270 );
xor ( n30272 , n30268 , n30270 );
and ( n30273 , n30269 , n29782 );
buf ( n30274 , n29725 );
and ( n30275 , n30274 , n29785 );
and ( n30276 , n30273 , n30275 );
xor ( n30277 , n30273 , n30275 );
and ( n30278 , n30274 , n29782 );
buf ( n30279 , n29727 );
and ( n30280 , n30279 , n29785 );
and ( n30281 , n30278 , n30280 );
xor ( n30282 , n30278 , n30280 );
and ( n30283 , n30279 , n29782 );
buf ( n30284 , n29729 );
and ( n30285 , n30284 , n29785 );
and ( n30286 , n30283 , n30285 );
xor ( n30287 , n30283 , n30285 );
and ( n30288 , n30284 , n29782 );
buf ( n30289 , n29731 );
and ( n30290 , n30289 , n29785 );
and ( n30291 , n30288 , n30290 );
xor ( n30292 , n30288 , n30290 );
and ( n30293 , n30289 , n29782 );
buf ( n30294 , n29733 );
and ( n30295 , n30294 , n29785 );
and ( n30296 , n30293 , n30295 );
xor ( n30297 , n30293 , n30295 );
and ( n30298 , n30294 , n29782 );
buf ( n30299 , n29735 );
and ( n30300 , n30299 , n29785 );
and ( n30301 , n30298 , n30300 );
xor ( n30302 , n30298 , n30300 );
and ( n30303 , n30299 , n29782 );
buf ( n30304 , n29737 );
and ( n30305 , n30304 , n29785 );
and ( n30306 , n30303 , n30305 );
xor ( n30307 , n30303 , n30305 );
and ( n30308 , n30304 , n29782 );
buf ( n30309 , n29739 );
and ( n30310 , n30309 , n29785 );
and ( n30311 , n30308 , n30310 );
xor ( n30312 , n30308 , n30310 );
and ( n30313 , n30309 , n29782 );
buf ( n30314 , n29741 );
and ( n30315 , n30314 , n29785 );
and ( n30316 , n30313 , n30315 );
xor ( n30317 , n30313 , n30315 );
and ( n30318 , n30314 , n29782 );
buf ( n30319 , n29743 );
and ( n30320 , n30319 , n29785 );
and ( n30321 , n30318 , n30320 );
xor ( n30322 , n30318 , n30320 );
and ( n30323 , n30319 , n29782 );
buf ( n30324 , n29745 );
and ( n30325 , n30324 , n29785 );
and ( n30326 , n30323 , n30325 );
xor ( n30327 , n30323 , n30325 );
and ( n30328 , n30324 , n29782 );
buf ( n30329 , n29747 );
and ( n30330 , n30329 , n29785 );
and ( n30331 , n30328 , n30330 );
xor ( n30332 , n30328 , n30330 );
and ( n30333 , n30329 , n29782 );
buf ( n30334 , n29749 );
and ( n30335 , n30334 , n29785 );
and ( n30336 , n30333 , n30335 );
xor ( n30337 , n30333 , n30335 );
and ( n30338 , n30334 , n29782 );
buf ( n30339 , n29751 );
and ( n30340 , n30339 , n29785 );
and ( n30341 , n30338 , n30340 );
xor ( n30342 , n30338 , n30340 );
and ( n30343 , n30339 , n29782 );
buf ( n30344 , n29753 );
and ( n30345 , n30344 , n29785 );
and ( n30346 , n30343 , n30345 );
xor ( n30347 , n30343 , n30345 );
and ( n30348 , n30344 , n29782 );
buf ( n30349 , n29755 );
and ( n30350 , n30349 , n29785 );
and ( n30351 , n30348 , n30350 );
xor ( n30352 , n30348 , n30350 );
and ( n30353 , n30349 , n29782 );
buf ( n30354 , n29757 );
and ( n30355 , n30354 , n29785 );
and ( n30356 , n30353 , n30355 );
xor ( n30357 , n30353 , n30355 );
and ( n30358 , n30354 , n29782 );
buf ( n30359 , n29759 );
and ( n30360 , n30359 , n29785 );
and ( n30361 , n30358 , n30360 );
xor ( n30362 , n30358 , n30360 );
and ( n30363 , n30359 , n29782 );
buf ( n30364 , n29761 );
and ( n30365 , n30364 , n29785 );
and ( n30366 , n30363 , n30365 );
xor ( n30367 , n30363 , n30365 );
and ( n30368 , n30364 , n29782 );
buf ( n30369 , n29763 );
and ( n30370 , n30369 , n29785 );
and ( n30371 , n30368 , n30370 );
xor ( n30372 , n30368 , n30370 );
and ( n30373 , n30369 , n29782 );
buf ( n30374 , n29765 );
and ( n30375 , n30374 , n29785 );
and ( n30376 , n30373 , n30375 );
xor ( n30377 , n30373 , n30375 );
and ( n30378 , n30374 , n29782 );
buf ( n30379 , n29767 );
and ( n30380 , n30379 , n29785 );
and ( n30381 , n30378 , n30380 );
xor ( n30382 , n30378 , n30380 );
and ( n30383 , n30379 , n29782 );
buf ( n30384 , n29769 );
and ( n30385 , n30384 , n29785 );
and ( n30386 , n30383 , n30385 );
xor ( n30387 , n30383 , n30385 );
and ( n30388 , n30384 , n29782 );
buf ( n30389 , n29771 );
and ( n30390 , n30389 , n29785 );
and ( n30391 , n30388 , n30390 );
xor ( n30392 , n30388 , n30390 );
and ( n30393 , n30389 , n29782 );
buf ( n30394 , n29773 );
and ( n30395 , n30394 , n29785 );
and ( n30396 , n30393 , n30395 );
xor ( n30397 , n30393 , n30395 );
and ( n30398 , n30394 , n29782 );
buf ( n30399 , n29775 );
and ( n30400 , n30399 , n29785 );
and ( n30401 , n30398 , n30400 );
xor ( n30402 , n30398 , n30400 );
and ( n30403 , n30399 , n29782 );
buf ( n30404 , n29777 );
and ( n30405 , n30404 , n29785 );
and ( n30406 , n30403 , n30405 );
xor ( n30407 , n30403 , n30405 );
and ( n30408 , n30404 , n29782 );
buf ( n30409 , n29780 );
and ( n30410 , n30409 , n29785 );
and ( n30411 , n30408 , n30410 );
buf ( n30412 , n30411 );
and ( n30413 , n30407 , n30412 );
or ( n30414 , n30406 , n30413 );
and ( n30415 , n30402 , n30414 );
or ( n30416 , n30401 , n30415 );
and ( n30417 , n30397 , n30416 );
or ( n30418 , n30396 , n30417 );
and ( n30419 , n30392 , n30418 );
or ( n30420 , n30391 , n30419 );
and ( n30421 , n30387 , n30420 );
or ( n30422 , n30386 , n30421 );
and ( n30423 , n30382 , n30422 );
or ( n30424 , n30381 , n30423 );
and ( n30425 , n30377 , n30424 );
or ( n30426 , n30376 , n30425 );
and ( n30427 , n30372 , n30426 );
or ( n30428 , n30371 , n30427 );
and ( n30429 , n30367 , n30428 );
or ( n30430 , n30366 , n30429 );
and ( n30431 , n30362 , n30430 );
or ( n30432 , n30361 , n30431 );
and ( n30433 , n30357 , n30432 );
or ( n30434 , n30356 , n30433 );
and ( n30435 , n30352 , n30434 );
or ( n30436 , n30351 , n30435 );
and ( n30437 , n30347 , n30436 );
or ( n30438 , n30346 , n30437 );
and ( n30439 , n30342 , n30438 );
or ( n30440 , n30341 , n30439 );
and ( n30441 , n30337 , n30440 );
or ( n30442 , n30336 , n30441 );
and ( n30443 , n30332 , n30442 );
or ( n30444 , n30331 , n30443 );
and ( n30445 , n30327 , n30444 );
or ( n30446 , n30326 , n30445 );
and ( n30447 , n30322 , n30446 );
or ( n30448 , n30321 , n30447 );
and ( n30449 , n30317 , n30448 );
or ( n30450 , n30316 , n30449 );
and ( n30451 , n30312 , n30450 );
or ( n30452 , n30311 , n30451 );
and ( n30453 , n30307 , n30452 );
or ( n30454 , n30306 , n30453 );
and ( n30455 , n30302 , n30454 );
or ( n30456 , n30301 , n30455 );
and ( n30457 , n30297 , n30456 );
or ( n30458 , n30296 , n30457 );
and ( n30459 , n30292 , n30458 );
or ( n30460 , n30291 , n30459 );
and ( n30461 , n30287 , n30460 );
or ( n30462 , n30286 , n30461 );
and ( n30463 , n30282 , n30462 );
or ( n30464 , n30281 , n30463 );
and ( n30465 , n30277 , n30464 );
or ( n30466 , n30276 , n30465 );
and ( n30467 , n30272 , n30466 );
or ( n30468 , n30271 , n30467 );
and ( n30469 , n30267 , n30468 );
or ( n30470 , n30266 , n30469 );
and ( n30471 , n30262 , n30470 );
or ( n30472 , n30261 , n30471 );
and ( n30473 , n30257 , n30472 );
or ( n30474 , n30256 , n30473 );
and ( n30475 , n30252 , n30474 );
or ( n30476 , n30251 , n30475 );
and ( n30477 , n30247 , n30476 );
or ( n30478 , n30246 , n30477 );
and ( n30479 , n30242 , n30478 );
or ( n30480 , n30241 , n30479 );
and ( n30481 , n30237 , n30480 );
or ( n30482 , n30236 , n30481 );
and ( n30483 , n30232 , n30482 );
or ( n30484 , n30231 , n30483 );
and ( n30485 , n30227 , n30484 );
or ( n30486 , n30226 , n30485 );
and ( n30487 , n30222 , n30486 );
or ( n30488 , n30221 , n30487 );
and ( n30489 , n30217 , n30488 );
or ( n30490 , n30216 , n30489 );
and ( n30491 , n30212 , n30490 );
or ( n30492 , n30211 , n30491 );
and ( n30493 , n30207 , n30492 );
or ( n30494 , n30206 , n30493 );
and ( n30495 , n30202 , n30494 );
or ( n30496 , n30201 , n30495 );
and ( n30497 , n30197 , n30496 );
or ( n30498 , n30196 , n30497 );
and ( n30499 , n30192 , n30498 );
or ( n30500 , n30191 , n30499 );
and ( n30501 , n30187 , n30500 );
or ( n30502 , n30186 , n30501 );
and ( n30503 , n30182 , n30502 );
or ( n30504 , n30181 , n30503 );
and ( n30505 , n30177 , n30504 );
or ( n30506 , n30176 , n30505 );
and ( n30507 , n30172 , n30506 );
or ( n30508 , n30171 , n30507 );
and ( n30509 , n30167 , n30508 );
or ( n30510 , n30166 , n30509 );
and ( n30511 , n30162 , n30510 );
or ( n30512 , n30161 , n30511 );
and ( n30513 , n30157 , n30512 );
or ( n30514 , n30156 , n30513 );
and ( n30515 , n30152 , n30514 );
or ( n30516 , n30151 , n30515 );
and ( n30517 , n30147 , n30516 );
or ( n30518 , n30146 , n30517 );
and ( n30519 , n30142 , n30518 );
or ( n30520 , n30141 , n30519 );
and ( n30521 , n30137 , n30520 );
or ( n30522 , n30136 , n30521 );
and ( n30523 , n30132 , n30522 );
or ( n30524 , n30131 , n30523 );
and ( n30525 , n30127 , n30524 );
or ( n30526 , n30126 , n30525 );
and ( n30527 , n30122 , n30526 );
or ( n30528 , n30121 , n30527 );
and ( n30529 , n30117 , n30528 );
or ( n30530 , n30116 , n30529 );
and ( n30531 , n30112 , n30530 );
or ( n30532 , n30111 , n30531 );
and ( n30533 , n30107 , n30532 );
or ( n30534 , n30106 , n30533 );
and ( n30535 , n30102 , n30534 );
or ( n30536 , n30101 , n30535 );
and ( n30537 , n30097 , n30536 );
or ( n30538 , n30096 , n30537 );
and ( n30539 , n30092 , n30538 );
or ( n30540 , n30091 , n30539 );
and ( n30541 , n30087 , n30540 );
or ( n30542 , n30086 , n30541 );
and ( n30543 , n30082 , n30542 );
or ( n30544 , n30081 , n30543 );
and ( n30545 , n30077 , n30544 );
or ( n30546 , n30076 , n30545 );
and ( n30547 , n30072 , n30546 );
or ( n30548 , n30071 , n30547 );
and ( n30549 , n30067 , n30548 );
or ( n30550 , n30066 , n30549 );
and ( n30551 , n30062 , n30550 );
or ( n30552 , n30061 , n30551 );
and ( n30553 , n30057 , n30552 );
or ( n30554 , n30056 , n30553 );
and ( n30555 , n30052 , n30554 );
or ( n30556 , n30051 , n30555 );
and ( n30557 , n30047 , n30556 );
or ( n30558 , n30046 , n30557 );
and ( n30559 , n30042 , n30558 );
or ( n30560 , n30041 , n30559 );
and ( n30561 , n30037 , n30560 );
or ( n30562 , n30036 , n30561 );
and ( n30563 , n30032 , n30562 );
or ( n30564 , n30031 , n30563 );
and ( n30565 , n30027 , n30564 );
or ( n30566 , n30026 , n30565 );
and ( n30567 , n30022 , n30566 );
or ( n30568 , n30021 , n30567 );
and ( n30569 , n30017 , n30568 );
or ( n30570 , n30016 , n30569 );
and ( n30571 , n30012 , n30570 );
or ( n30572 , n30011 , n30571 );
and ( n30573 , n30007 , n30572 );
or ( n30574 , n30006 , n30573 );
and ( n30575 , n30002 , n30574 );
or ( n30576 , n30001 , n30575 );
and ( n30577 , n29997 , n30576 );
or ( n30578 , n29996 , n30577 );
and ( n30579 , n29992 , n30578 );
or ( n30580 , n29991 , n30579 );
and ( n30581 , n29987 , n30580 );
or ( n30582 , n29986 , n30581 );
and ( n30583 , n29982 , n30582 );
or ( n30584 , n29981 , n30583 );
and ( n30585 , n29977 , n30584 );
or ( n30586 , n29976 , n30585 );
and ( n30587 , n29972 , n30586 );
or ( n30588 , n29971 , n30587 );
and ( n30589 , n29967 , n30588 );
or ( n30590 , n29966 , n30589 );
and ( n30591 , n29962 , n30590 );
or ( n30592 , n29961 , n30591 );
and ( n30593 , n29957 , n30592 );
or ( n30594 , n29956 , n30593 );
and ( n30595 , n29952 , n30594 );
or ( n30596 , n29951 , n30595 );
and ( n30597 , n29947 , n30596 );
or ( n30598 , n29946 , n30597 );
and ( n30599 , n29942 , n30598 );
or ( n30600 , n29941 , n30599 );
and ( n30601 , n29937 , n30600 );
or ( n30602 , n29936 , n30601 );
and ( n30603 , n29932 , n30602 );
or ( n30604 , n29931 , n30603 );
and ( n30605 , n29927 , n30604 );
or ( n30606 , n29926 , n30605 );
and ( n30607 , n29922 , n30606 );
or ( n30608 , n29921 , n30607 );
and ( n30609 , n29917 , n30608 );
or ( n30610 , n29916 , n30609 );
and ( n30611 , n29912 , n30610 );
or ( n30612 , n29911 , n30611 );
and ( n30613 , n29907 , n30612 );
or ( n30614 , n29906 , n30613 );
and ( n30615 , n29902 , n30614 );
or ( n30616 , n29901 , n30615 );
and ( n30617 , n29897 , n30616 );
or ( n30618 , n29896 , n30617 );
and ( n30619 , n29892 , n30618 );
or ( n30620 , n29891 , n30619 );
and ( n30621 , n29887 , n30620 );
or ( n30622 , n29886 , n30621 );
and ( n30623 , n29882 , n30622 );
or ( n30624 , n29881 , n30623 );
and ( n30625 , n29877 , n30624 );
or ( n30626 , n29876 , n30625 );
and ( n30627 , n29872 , n30626 );
or ( n30628 , n29871 , n30627 );
and ( n30629 , n29867 , n30628 );
or ( n30630 , n29866 , n30629 );
and ( n30631 , n29862 , n30630 );
or ( n30632 , n29861 , n30631 );
and ( n30633 , n29857 , n30632 );
or ( n30634 , n29856 , n30633 );
and ( n30635 , n29852 , n30634 );
or ( n30636 , n29851 , n30635 );
and ( n30637 , n29847 , n30636 );
or ( n30638 , n29846 , n30637 );
and ( n30639 , n29842 , n30638 );
or ( n30640 , n29841 , n30639 );
and ( n30641 , n29837 , n30640 );
or ( n30642 , n29836 , n30641 );
and ( n30643 , n29832 , n30642 );
or ( n30644 , n29831 , n30643 );
and ( n30645 , n29827 , n30644 );
or ( n30646 , n29826 , n30645 );
and ( n30647 , n29822 , n30646 );
or ( n30648 , n29821 , n30647 );
and ( n30649 , n29817 , n30648 );
or ( n30650 , n29816 , n30649 );
and ( n30651 , n29812 , n30650 );
or ( n30652 , n29811 , n30651 );
and ( n30653 , n29807 , n30652 );
or ( n30654 , n29806 , n30653 );
and ( n30655 , n29802 , n30654 );
or ( n30656 , n29801 , n30655 );
and ( n30657 , n29797 , n30656 );
or ( n30658 , n29796 , n30657 );
and ( n30659 , n29792 , n30658 );
or ( n30660 , n29791 , n30659 );
xor ( n30661 , n29787 , n30660 );
buf ( n30662 , n18102 );
and ( n30663 , n29789 , n30662 );
xor ( n30664 , n30661 , n30663 );
xor ( n30665 , n29792 , n30658 );
and ( n30666 , n29794 , n30662 );
and ( n30667 , n30665 , n30666 );
xor ( n30668 , n30665 , n30666 );
xor ( n30669 , n29797 , n30656 );
and ( n30670 , n29799 , n30662 );
and ( n30671 , n30669 , n30670 );
xor ( n30672 , n30669 , n30670 );
xor ( n30673 , n29802 , n30654 );
and ( n30674 , n29804 , n30662 );
and ( n30675 , n30673 , n30674 );
xor ( n30676 , n30673 , n30674 );
xor ( n30677 , n29807 , n30652 );
and ( n30678 , n29809 , n30662 );
and ( n30679 , n30677 , n30678 );
xor ( n30680 , n30677 , n30678 );
xor ( n30681 , n29812 , n30650 );
and ( n30682 , n29814 , n30662 );
and ( n30683 , n30681 , n30682 );
xor ( n30684 , n30681 , n30682 );
xor ( n30685 , n29817 , n30648 );
and ( n30686 , n29819 , n30662 );
and ( n30687 , n30685 , n30686 );
xor ( n30688 , n30685 , n30686 );
xor ( n30689 , n29822 , n30646 );
and ( n30690 , n29824 , n30662 );
and ( n30691 , n30689 , n30690 );
xor ( n30692 , n30689 , n30690 );
xor ( n30693 , n29827 , n30644 );
and ( n30694 , n29829 , n30662 );
and ( n30695 , n30693 , n30694 );
xor ( n30696 , n30693 , n30694 );
xor ( n30697 , n29832 , n30642 );
and ( n30698 , n29834 , n30662 );
and ( n30699 , n30697 , n30698 );
xor ( n30700 , n30697 , n30698 );
xor ( n30701 , n29837 , n30640 );
and ( n30702 , n29839 , n30662 );
and ( n30703 , n30701 , n30702 );
xor ( n30704 , n30701 , n30702 );
xor ( n30705 , n29842 , n30638 );
and ( n30706 , n29844 , n30662 );
and ( n30707 , n30705 , n30706 );
xor ( n30708 , n30705 , n30706 );
xor ( n30709 , n29847 , n30636 );
and ( n30710 , n29849 , n30662 );
and ( n30711 , n30709 , n30710 );
xor ( n30712 , n30709 , n30710 );
xor ( n30713 , n29852 , n30634 );
and ( n30714 , n29854 , n30662 );
and ( n30715 , n30713 , n30714 );
xor ( n30716 , n30713 , n30714 );
xor ( n30717 , n29857 , n30632 );
and ( n30718 , n29859 , n30662 );
and ( n30719 , n30717 , n30718 );
xor ( n30720 , n30717 , n30718 );
xor ( n30721 , n29862 , n30630 );
and ( n30722 , n29864 , n30662 );
and ( n30723 , n30721 , n30722 );
xor ( n30724 , n30721 , n30722 );
xor ( n30725 , n29867 , n30628 );
and ( n30726 , n29869 , n30662 );
and ( n30727 , n30725 , n30726 );
xor ( n30728 , n30725 , n30726 );
xor ( n30729 , n29872 , n30626 );
and ( n30730 , n29874 , n30662 );
and ( n30731 , n30729 , n30730 );
xor ( n30732 , n30729 , n30730 );
xor ( n30733 , n29877 , n30624 );
and ( n30734 , n29879 , n30662 );
and ( n30735 , n30733 , n30734 );
xor ( n30736 , n30733 , n30734 );
xor ( n30737 , n29882 , n30622 );
and ( n30738 , n29884 , n30662 );
and ( n30739 , n30737 , n30738 );
xor ( n30740 , n30737 , n30738 );
xor ( n30741 , n29887 , n30620 );
and ( n30742 , n29889 , n30662 );
and ( n30743 , n30741 , n30742 );
xor ( n30744 , n30741 , n30742 );
xor ( n30745 , n29892 , n30618 );
and ( n30746 , n29894 , n30662 );
and ( n30747 , n30745 , n30746 );
xor ( n30748 , n30745 , n30746 );
xor ( n30749 , n29897 , n30616 );
and ( n30750 , n29899 , n30662 );
and ( n30751 , n30749 , n30750 );
xor ( n30752 , n30749 , n30750 );
xor ( n30753 , n29902 , n30614 );
and ( n30754 , n29904 , n30662 );
and ( n30755 , n30753 , n30754 );
xor ( n30756 , n30753 , n30754 );
xor ( n30757 , n29907 , n30612 );
and ( n30758 , n29909 , n30662 );
and ( n30759 , n30757 , n30758 );
xor ( n30760 , n30757 , n30758 );
xor ( n30761 , n29912 , n30610 );
and ( n30762 , n29914 , n30662 );
and ( n30763 , n30761 , n30762 );
xor ( n30764 , n30761 , n30762 );
xor ( n30765 , n29917 , n30608 );
and ( n30766 , n29919 , n30662 );
and ( n30767 , n30765 , n30766 );
xor ( n30768 , n30765 , n30766 );
xor ( n30769 , n29922 , n30606 );
and ( n30770 , n29924 , n30662 );
and ( n30771 , n30769 , n30770 );
xor ( n30772 , n30769 , n30770 );
xor ( n30773 , n29927 , n30604 );
and ( n30774 , n29929 , n30662 );
and ( n30775 , n30773 , n30774 );
xor ( n30776 , n30773 , n30774 );
xor ( n30777 , n29932 , n30602 );
and ( n30778 , n29934 , n30662 );
and ( n30779 , n30777 , n30778 );
xor ( n30780 , n30777 , n30778 );
xor ( n30781 , n29937 , n30600 );
and ( n30782 , n29939 , n30662 );
and ( n30783 , n30781 , n30782 );
xor ( n30784 , n30781 , n30782 );
xor ( n30785 , n29942 , n30598 );
and ( n30786 , n29944 , n30662 );
and ( n30787 , n30785 , n30786 );
xor ( n30788 , n30785 , n30786 );
xor ( n30789 , n29947 , n30596 );
and ( n30790 , n29949 , n30662 );
and ( n30791 , n30789 , n30790 );
xor ( n30792 , n30789 , n30790 );
xor ( n30793 , n29952 , n30594 );
and ( n30794 , n29954 , n30662 );
and ( n30795 , n30793 , n30794 );
xor ( n30796 , n30793 , n30794 );
xor ( n30797 , n29957 , n30592 );
and ( n30798 , n29959 , n30662 );
and ( n30799 , n30797 , n30798 );
xor ( n30800 , n30797 , n30798 );
xor ( n30801 , n29962 , n30590 );
and ( n30802 , n29964 , n30662 );
and ( n30803 , n30801 , n30802 );
xor ( n30804 , n30801 , n30802 );
xor ( n30805 , n29967 , n30588 );
and ( n30806 , n29969 , n30662 );
and ( n30807 , n30805 , n30806 );
xor ( n30808 , n30805 , n30806 );
xor ( n30809 , n29972 , n30586 );
and ( n30810 , n29974 , n30662 );
and ( n30811 , n30809 , n30810 );
xor ( n30812 , n30809 , n30810 );
xor ( n30813 , n29977 , n30584 );
and ( n30814 , n29979 , n30662 );
and ( n30815 , n30813 , n30814 );
xor ( n30816 , n30813 , n30814 );
xor ( n30817 , n29982 , n30582 );
and ( n30818 , n29984 , n30662 );
and ( n30819 , n30817 , n30818 );
xor ( n30820 , n30817 , n30818 );
xor ( n30821 , n29987 , n30580 );
and ( n30822 , n29989 , n30662 );
and ( n30823 , n30821 , n30822 );
xor ( n30824 , n30821 , n30822 );
xor ( n30825 , n29992 , n30578 );
and ( n30826 , n29994 , n30662 );
and ( n30827 , n30825 , n30826 );
xor ( n30828 , n30825 , n30826 );
xor ( n30829 , n29997 , n30576 );
and ( n30830 , n29999 , n30662 );
and ( n30831 , n30829 , n30830 );
xor ( n30832 , n30829 , n30830 );
xor ( n30833 , n30002 , n30574 );
and ( n30834 , n30004 , n30662 );
and ( n30835 , n30833 , n30834 );
xor ( n30836 , n30833 , n30834 );
xor ( n30837 , n30007 , n30572 );
and ( n30838 , n30009 , n30662 );
and ( n30839 , n30837 , n30838 );
xor ( n30840 , n30837 , n30838 );
xor ( n30841 , n30012 , n30570 );
and ( n30842 , n30014 , n30662 );
and ( n30843 , n30841 , n30842 );
xor ( n30844 , n30841 , n30842 );
xor ( n30845 , n30017 , n30568 );
and ( n30846 , n30019 , n30662 );
and ( n30847 , n30845 , n30846 );
xor ( n30848 , n30845 , n30846 );
xor ( n30849 , n30022 , n30566 );
and ( n30850 , n30024 , n30662 );
and ( n30851 , n30849 , n30850 );
xor ( n30852 , n30849 , n30850 );
xor ( n30853 , n30027 , n30564 );
and ( n30854 , n30029 , n30662 );
and ( n30855 , n30853 , n30854 );
xor ( n30856 , n30853 , n30854 );
xor ( n30857 , n30032 , n30562 );
and ( n30858 , n30034 , n30662 );
and ( n30859 , n30857 , n30858 );
xor ( n30860 , n30857 , n30858 );
xor ( n30861 , n30037 , n30560 );
and ( n30862 , n30039 , n30662 );
and ( n30863 , n30861 , n30862 );
xor ( n30864 , n30861 , n30862 );
xor ( n30865 , n30042 , n30558 );
and ( n30866 , n30044 , n30662 );
and ( n30867 , n30865 , n30866 );
xor ( n30868 , n30865 , n30866 );
xor ( n30869 , n30047 , n30556 );
and ( n30870 , n30049 , n30662 );
and ( n30871 , n30869 , n30870 );
xor ( n30872 , n30869 , n30870 );
xor ( n30873 , n30052 , n30554 );
and ( n30874 , n30054 , n30662 );
and ( n30875 , n30873 , n30874 );
xor ( n30876 , n30873 , n30874 );
xor ( n30877 , n30057 , n30552 );
and ( n30878 , n30059 , n30662 );
and ( n30879 , n30877 , n30878 );
xor ( n30880 , n30877 , n30878 );
xor ( n30881 , n30062 , n30550 );
and ( n30882 , n30064 , n30662 );
and ( n30883 , n30881 , n30882 );
xor ( n30884 , n30881 , n30882 );
xor ( n30885 , n30067 , n30548 );
and ( n30886 , n30069 , n30662 );
and ( n30887 , n30885 , n30886 );
xor ( n30888 , n30885 , n30886 );
xor ( n30889 , n30072 , n30546 );
and ( n30890 , n30074 , n30662 );
and ( n30891 , n30889 , n30890 );
xor ( n30892 , n30889 , n30890 );
xor ( n30893 , n30077 , n30544 );
and ( n30894 , n30079 , n30662 );
and ( n30895 , n30893 , n30894 );
xor ( n30896 , n30893 , n30894 );
xor ( n30897 , n30082 , n30542 );
and ( n30898 , n30084 , n30662 );
and ( n30899 , n30897 , n30898 );
xor ( n30900 , n30897 , n30898 );
xor ( n30901 , n30087 , n30540 );
and ( n30902 , n30089 , n30662 );
and ( n30903 , n30901 , n30902 );
xor ( n30904 , n30901 , n30902 );
xor ( n30905 , n30092 , n30538 );
and ( n30906 , n30094 , n30662 );
and ( n30907 , n30905 , n30906 );
xor ( n30908 , n30905 , n30906 );
xor ( n30909 , n30097 , n30536 );
and ( n30910 , n30099 , n30662 );
and ( n30911 , n30909 , n30910 );
xor ( n30912 , n30909 , n30910 );
xor ( n30913 , n30102 , n30534 );
and ( n30914 , n30104 , n30662 );
and ( n30915 , n30913 , n30914 );
xor ( n30916 , n30913 , n30914 );
xor ( n30917 , n30107 , n30532 );
and ( n30918 , n30109 , n30662 );
and ( n30919 , n30917 , n30918 );
xor ( n30920 , n30917 , n30918 );
xor ( n30921 , n30112 , n30530 );
and ( n30922 , n30114 , n30662 );
and ( n30923 , n30921 , n30922 );
xor ( n30924 , n30921 , n30922 );
xor ( n30925 , n30117 , n30528 );
and ( n30926 , n30119 , n30662 );
and ( n30927 , n30925 , n30926 );
xor ( n30928 , n30925 , n30926 );
xor ( n30929 , n30122 , n30526 );
and ( n30930 , n30124 , n30662 );
and ( n30931 , n30929 , n30930 );
xor ( n30932 , n30929 , n30930 );
xor ( n30933 , n30127 , n30524 );
and ( n30934 , n30129 , n30662 );
and ( n30935 , n30933 , n30934 );
xor ( n30936 , n30933 , n30934 );
xor ( n30937 , n30132 , n30522 );
and ( n30938 , n30134 , n30662 );
and ( n30939 , n30937 , n30938 );
xor ( n30940 , n30937 , n30938 );
xor ( n30941 , n30137 , n30520 );
and ( n30942 , n30139 , n30662 );
and ( n30943 , n30941 , n30942 );
xor ( n30944 , n30941 , n30942 );
xor ( n30945 , n30142 , n30518 );
and ( n30946 , n30144 , n30662 );
and ( n30947 , n30945 , n30946 );
xor ( n30948 , n30945 , n30946 );
xor ( n30949 , n30147 , n30516 );
and ( n30950 , n30149 , n30662 );
and ( n30951 , n30949 , n30950 );
xor ( n30952 , n30949 , n30950 );
xor ( n30953 , n30152 , n30514 );
and ( n30954 , n30154 , n30662 );
and ( n30955 , n30953 , n30954 );
xor ( n30956 , n30953 , n30954 );
xor ( n30957 , n30157 , n30512 );
and ( n30958 , n30159 , n30662 );
and ( n30959 , n30957 , n30958 );
xor ( n30960 , n30957 , n30958 );
xor ( n30961 , n30162 , n30510 );
and ( n30962 , n30164 , n30662 );
and ( n30963 , n30961 , n30962 );
xor ( n30964 , n30961 , n30962 );
xor ( n30965 , n30167 , n30508 );
and ( n30966 , n30169 , n30662 );
and ( n30967 , n30965 , n30966 );
xor ( n30968 , n30965 , n30966 );
xor ( n30969 , n30172 , n30506 );
and ( n30970 , n30174 , n30662 );
and ( n30971 , n30969 , n30970 );
xor ( n30972 , n30969 , n30970 );
xor ( n30973 , n30177 , n30504 );
and ( n30974 , n30179 , n30662 );
and ( n30975 , n30973 , n30974 );
xor ( n30976 , n30973 , n30974 );
xor ( n30977 , n30182 , n30502 );
and ( n30978 , n30184 , n30662 );
and ( n30979 , n30977 , n30978 );
xor ( n30980 , n30977 , n30978 );
xor ( n30981 , n30187 , n30500 );
and ( n30982 , n30189 , n30662 );
and ( n30983 , n30981 , n30982 );
xor ( n30984 , n30981 , n30982 );
xor ( n30985 , n30192 , n30498 );
and ( n30986 , n30194 , n30662 );
and ( n30987 , n30985 , n30986 );
xor ( n30988 , n30985 , n30986 );
xor ( n30989 , n30197 , n30496 );
and ( n30990 , n30199 , n30662 );
and ( n30991 , n30989 , n30990 );
xor ( n30992 , n30989 , n30990 );
xor ( n30993 , n30202 , n30494 );
and ( n30994 , n30204 , n30662 );
and ( n30995 , n30993 , n30994 );
xor ( n30996 , n30993 , n30994 );
xor ( n30997 , n30207 , n30492 );
and ( n30998 , n30209 , n30662 );
and ( n30999 , n30997 , n30998 );
xor ( n31000 , n30997 , n30998 );
xor ( n31001 , n30212 , n30490 );
and ( n31002 , n30214 , n30662 );
and ( n31003 , n31001 , n31002 );
xor ( n31004 , n31001 , n31002 );
xor ( n31005 , n30217 , n30488 );
and ( n31006 , n30219 , n30662 );
and ( n31007 , n31005 , n31006 );
xor ( n31008 , n31005 , n31006 );
xor ( n31009 , n30222 , n30486 );
and ( n31010 , n30224 , n30662 );
and ( n31011 , n31009 , n31010 );
xor ( n31012 , n31009 , n31010 );
xor ( n31013 , n30227 , n30484 );
and ( n31014 , n30229 , n30662 );
and ( n31015 , n31013 , n31014 );
xor ( n31016 , n31013 , n31014 );
xor ( n31017 , n30232 , n30482 );
and ( n31018 , n30234 , n30662 );
and ( n31019 , n31017 , n31018 );
xor ( n31020 , n31017 , n31018 );
xor ( n31021 , n30237 , n30480 );
and ( n31022 , n30239 , n30662 );
and ( n31023 , n31021 , n31022 );
xor ( n31024 , n31021 , n31022 );
xor ( n31025 , n30242 , n30478 );
and ( n31026 , n30244 , n30662 );
and ( n31027 , n31025 , n31026 );
xor ( n31028 , n31025 , n31026 );
xor ( n31029 , n30247 , n30476 );
and ( n31030 , n30249 , n30662 );
and ( n31031 , n31029 , n31030 );
xor ( n31032 , n31029 , n31030 );
xor ( n31033 , n30252 , n30474 );
and ( n31034 , n30254 , n30662 );
and ( n31035 , n31033 , n31034 );
xor ( n31036 , n31033 , n31034 );
xor ( n31037 , n30257 , n30472 );
and ( n31038 , n30259 , n30662 );
and ( n31039 , n31037 , n31038 );
xor ( n31040 , n31037 , n31038 );
xor ( n31041 , n30262 , n30470 );
and ( n31042 , n30264 , n30662 );
and ( n31043 , n31041 , n31042 );
xor ( n31044 , n31041 , n31042 );
xor ( n31045 , n30267 , n30468 );
and ( n31046 , n30269 , n30662 );
and ( n31047 , n31045 , n31046 );
xor ( n31048 , n31045 , n31046 );
xor ( n31049 , n30272 , n30466 );
and ( n31050 , n30274 , n30662 );
and ( n31051 , n31049 , n31050 );
xor ( n31052 , n31049 , n31050 );
xor ( n31053 , n30277 , n30464 );
and ( n31054 , n30279 , n30662 );
and ( n31055 , n31053 , n31054 );
xor ( n31056 , n31053 , n31054 );
xor ( n31057 , n30282 , n30462 );
and ( n31058 , n30284 , n30662 );
and ( n31059 , n31057 , n31058 );
xor ( n31060 , n31057 , n31058 );
xor ( n31061 , n30287 , n30460 );
and ( n31062 , n30289 , n30662 );
and ( n31063 , n31061 , n31062 );
xor ( n31064 , n31061 , n31062 );
xor ( n31065 , n30292 , n30458 );
and ( n31066 , n30294 , n30662 );
and ( n31067 , n31065 , n31066 );
xor ( n31068 , n31065 , n31066 );
xor ( n31069 , n30297 , n30456 );
and ( n31070 , n30299 , n30662 );
and ( n31071 , n31069 , n31070 );
xor ( n31072 , n31069 , n31070 );
xor ( n31073 , n30302 , n30454 );
and ( n31074 , n30304 , n30662 );
and ( n31075 , n31073 , n31074 );
xor ( n31076 , n31073 , n31074 );
xor ( n31077 , n30307 , n30452 );
and ( n31078 , n30309 , n30662 );
and ( n31079 , n31077 , n31078 );
xor ( n31080 , n31077 , n31078 );
xor ( n31081 , n30312 , n30450 );
and ( n31082 , n30314 , n30662 );
and ( n31083 , n31081 , n31082 );
xor ( n31084 , n31081 , n31082 );
xor ( n31085 , n30317 , n30448 );
and ( n31086 , n30319 , n30662 );
and ( n31087 , n31085 , n31086 );
xor ( n31088 , n31085 , n31086 );
xor ( n31089 , n30322 , n30446 );
and ( n31090 , n30324 , n30662 );
and ( n31091 , n31089 , n31090 );
xor ( n31092 , n31089 , n31090 );
xor ( n31093 , n30327 , n30444 );
and ( n31094 , n30329 , n30662 );
and ( n31095 , n31093 , n31094 );
xor ( n31096 , n31093 , n31094 );
xor ( n31097 , n30332 , n30442 );
and ( n31098 , n30334 , n30662 );
and ( n31099 , n31097 , n31098 );
xor ( n31100 , n31097 , n31098 );
xor ( n31101 , n30337 , n30440 );
and ( n31102 , n30339 , n30662 );
and ( n31103 , n31101 , n31102 );
xor ( n31104 , n31101 , n31102 );
xor ( n31105 , n30342 , n30438 );
and ( n31106 , n30344 , n30662 );
and ( n31107 , n31105 , n31106 );
xor ( n31108 , n31105 , n31106 );
xor ( n31109 , n30347 , n30436 );
and ( n31110 , n30349 , n30662 );
and ( n31111 , n31109 , n31110 );
xor ( n31112 , n31109 , n31110 );
xor ( n31113 , n30352 , n30434 );
and ( n31114 , n30354 , n30662 );
and ( n31115 , n31113 , n31114 );
xor ( n31116 , n31113 , n31114 );
xor ( n31117 , n30357 , n30432 );
and ( n31118 , n30359 , n30662 );
and ( n31119 , n31117 , n31118 );
xor ( n31120 , n31117 , n31118 );
xor ( n31121 , n30362 , n30430 );
and ( n31122 , n30364 , n30662 );
and ( n31123 , n31121 , n31122 );
xor ( n31124 , n31121 , n31122 );
xor ( n31125 , n30367 , n30428 );
and ( n31126 , n30369 , n30662 );
and ( n31127 , n31125 , n31126 );
xor ( n31128 , n31125 , n31126 );
xor ( n31129 , n30372 , n30426 );
and ( n31130 , n30374 , n30662 );
and ( n31131 , n31129 , n31130 );
xor ( n31132 , n31129 , n31130 );
xor ( n31133 , n30377 , n30424 );
and ( n31134 , n30379 , n30662 );
and ( n31135 , n31133 , n31134 );
xor ( n31136 , n31133 , n31134 );
xor ( n31137 , n30382 , n30422 );
and ( n31138 , n30384 , n30662 );
and ( n31139 , n31137 , n31138 );
xor ( n31140 , n31137 , n31138 );
xor ( n31141 , n30387 , n30420 );
and ( n31142 , n30389 , n30662 );
and ( n31143 , n31141 , n31142 );
xor ( n31144 , n31141 , n31142 );
xor ( n31145 , n30392 , n30418 );
and ( n31146 , n30394 , n30662 );
and ( n31147 , n31145 , n31146 );
xor ( n31148 , n31145 , n31146 );
xor ( n31149 , n30397 , n30416 );
and ( n31150 , n30399 , n30662 );
and ( n31151 , n31149 , n31150 );
xor ( n31152 , n31149 , n31150 );
xor ( n31153 , n30402 , n30414 );
and ( n31154 , n30404 , n30662 );
and ( n31155 , n31153 , n31154 );
xor ( n31156 , n31153 , n31154 );
xor ( n31157 , n30407 , n30412 );
and ( n31158 , n30409 , n30662 );
and ( n31159 , n31157 , n31158 );
buf ( n31160 , n31159 );
and ( n31161 , n31156 , n31160 );
or ( n31162 , n31155 , n31161 );
and ( n31163 , n31152 , n31162 );
or ( n31164 , n31151 , n31163 );
and ( n31165 , n31148 , n31164 );
or ( n31166 , n31147 , n31165 );
and ( n31167 , n31144 , n31166 );
or ( n31168 , n31143 , n31167 );
and ( n31169 , n31140 , n31168 );
or ( n31170 , n31139 , n31169 );
and ( n31171 , n31136 , n31170 );
or ( n31172 , n31135 , n31171 );
and ( n31173 , n31132 , n31172 );
or ( n31174 , n31131 , n31173 );
and ( n31175 , n31128 , n31174 );
or ( n31176 , n31127 , n31175 );
and ( n31177 , n31124 , n31176 );
or ( n31178 , n31123 , n31177 );
and ( n31179 , n31120 , n31178 );
or ( n31180 , n31119 , n31179 );
and ( n31181 , n31116 , n31180 );
or ( n31182 , n31115 , n31181 );
and ( n31183 , n31112 , n31182 );
or ( n31184 , n31111 , n31183 );
and ( n31185 , n31108 , n31184 );
or ( n31186 , n31107 , n31185 );
and ( n31187 , n31104 , n31186 );
or ( n31188 , n31103 , n31187 );
and ( n31189 , n31100 , n31188 );
or ( n31190 , n31099 , n31189 );
and ( n31191 , n31096 , n31190 );
or ( n31192 , n31095 , n31191 );
and ( n31193 , n31092 , n31192 );
or ( n31194 , n31091 , n31193 );
and ( n31195 , n31088 , n31194 );
or ( n31196 , n31087 , n31195 );
and ( n31197 , n31084 , n31196 );
or ( n31198 , n31083 , n31197 );
and ( n31199 , n31080 , n31198 );
or ( n31200 , n31079 , n31199 );
and ( n31201 , n31076 , n31200 );
or ( n31202 , n31075 , n31201 );
and ( n31203 , n31072 , n31202 );
or ( n31204 , n31071 , n31203 );
and ( n31205 , n31068 , n31204 );
or ( n31206 , n31067 , n31205 );
and ( n31207 , n31064 , n31206 );
or ( n31208 , n31063 , n31207 );
and ( n31209 , n31060 , n31208 );
or ( n31210 , n31059 , n31209 );
and ( n31211 , n31056 , n31210 );
or ( n31212 , n31055 , n31211 );
and ( n31213 , n31052 , n31212 );
or ( n31214 , n31051 , n31213 );
and ( n31215 , n31048 , n31214 );
or ( n31216 , n31047 , n31215 );
and ( n31217 , n31044 , n31216 );
or ( n31218 , n31043 , n31217 );
and ( n31219 , n31040 , n31218 );
or ( n31220 , n31039 , n31219 );
and ( n31221 , n31036 , n31220 );
or ( n31222 , n31035 , n31221 );
and ( n31223 , n31032 , n31222 );
or ( n31224 , n31031 , n31223 );
and ( n31225 , n31028 , n31224 );
or ( n31226 , n31027 , n31225 );
and ( n31227 , n31024 , n31226 );
or ( n31228 , n31023 , n31227 );
and ( n31229 , n31020 , n31228 );
or ( n31230 , n31019 , n31229 );
and ( n31231 , n31016 , n31230 );
or ( n31232 , n31015 , n31231 );
and ( n31233 , n31012 , n31232 );
or ( n31234 , n31011 , n31233 );
and ( n31235 , n31008 , n31234 );
or ( n31236 , n31007 , n31235 );
and ( n31237 , n31004 , n31236 );
or ( n31238 , n31003 , n31237 );
and ( n31239 , n31000 , n31238 );
or ( n31240 , n30999 , n31239 );
and ( n31241 , n30996 , n31240 );
or ( n31242 , n30995 , n31241 );
and ( n31243 , n30992 , n31242 );
or ( n31244 , n30991 , n31243 );
and ( n31245 , n30988 , n31244 );
or ( n31246 , n30987 , n31245 );
and ( n31247 , n30984 , n31246 );
or ( n31248 , n30983 , n31247 );
and ( n31249 , n30980 , n31248 );
or ( n31250 , n30979 , n31249 );
and ( n31251 , n30976 , n31250 );
or ( n31252 , n30975 , n31251 );
and ( n31253 , n30972 , n31252 );
or ( n31254 , n30971 , n31253 );
and ( n31255 , n30968 , n31254 );
or ( n31256 , n30967 , n31255 );
and ( n31257 , n30964 , n31256 );
or ( n31258 , n30963 , n31257 );
and ( n31259 , n30960 , n31258 );
or ( n31260 , n30959 , n31259 );
and ( n31261 , n30956 , n31260 );
or ( n31262 , n30955 , n31261 );
and ( n31263 , n30952 , n31262 );
or ( n31264 , n30951 , n31263 );
and ( n31265 , n30948 , n31264 );
or ( n31266 , n30947 , n31265 );
and ( n31267 , n30944 , n31266 );
or ( n31268 , n30943 , n31267 );
and ( n31269 , n30940 , n31268 );
or ( n31270 , n30939 , n31269 );
and ( n31271 , n30936 , n31270 );
or ( n31272 , n30935 , n31271 );
and ( n31273 , n30932 , n31272 );
or ( n31274 , n30931 , n31273 );
and ( n31275 , n30928 , n31274 );
or ( n31276 , n30927 , n31275 );
and ( n31277 , n30924 , n31276 );
or ( n31278 , n30923 , n31277 );
and ( n31279 , n30920 , n31278 );
or ( n31280 , n30919 , n31279 );
and ( n31281 , n30916 , n31280 );
or ( n31282 , n30915 , n31281 );
and ( n31283 , n30912 , n31282 );
or ( n31284 , n30911 , n31283 );
and ( n31285 , n30908 , n31284 );
or ( n31286 , n30907 , n31285 );
and ( n31287 , n30904 , n31286 );
or ( n31288 , n30903 , n31287 );
and ( n31289 , n30900 , n31288 );
or ( n31290 , n30899 , n31289 );
and ( n31291 , n30896 , n31290 );
or ( n31292 , n30895 , n31291 );
and ( n31293 , n30892 , n31292 );
or ( n31294 , n30891 , n31293 );
and ( n31295 , n30888 , n31294 );
or ( n31296 , n30887 , n31295 );
and ( n31297 , n30884 , n31296 );
or ( n31298 , n30883 , n31297 );
and ( n31299 , n30880 , n31298 );
or ( n31300 , n30879 , n31299 );
and ( n31301 , n30876 , n31300 );
or ( n31302 , n30875 , n31301 );
and ( n31303 , n30872 , n31302 );
or ( n31304 , n30871 , n31303 );
and ( n31305 , n30868 , n31304 );
or ( n31306 , n30867 , n31305 );
and ( n31307 , n30864 , n31306 );
or ( n31308 , n30863 , n31307 );
and ( n31309 , n30860 , n31308 );
or ( n31310 , n30859 , n31309 );
and ( n31311 , n30856 , n31310 );
or ( n31312 , n30855 , n31311 );
and ( n31313 , n30852 , n31312 );
or ( n31314 , n30851 , n31313 );
and ( n31315 , n30848 , n31314 );
or ( n31316 , n30847 , n31315 );
and ( n31317 , n30844 , n31316 );
or ( n31318 , n30843 , n31317 );
and ( n31319 , n30840 , n31318 );
or ( n31320 , n30839 , n31319 );
and ( n31321 , n30836 , n31320 );
or ( n31322 , n30835 , n31321 );
and ( n31323 , n30832 , n31322 );
or ( n31324 , n30831 , n31323 );
and ( n31325 , n30828 , n31324 );
or ( n31326 , n30827 , n31325 );
and ( n31327 , n30824 , n31326 );
or ( n31328 , n30823 , n31327 );
and ( n31329 , n30820 , n31328 );
or ( n31330 , n30819 , n31329 );
and ( n31331 , n30816 , n31330 );
or ( n31332 , n30815 , n31331 );
and ( n31333 , n30812 , n31332 );
or ( n31334 , n30811 , n31333 );
and ( n31335 , n30808 , n31334 );
or ( n31336 , n30807 , n31335 );
and ( n31337 , n30804 , n31336 );
or ( n31338 , n30803 , n31337 );
and ( n31339 , n30800 , n31338 );
or ( n31340 , n30799 , n31339 );
and ( n31341 , n30796 , n31340 );
or ( n31342 , n30795 , n31341 );
and ( n31343 , n30792 , n31342 );
or ( n31344 , n30791 , n31343 );
and ( n31345 , n30788 , n31344 );
or ( n31346 , n30787 , n31345 );
and ( n31347 , n30784 , n31346 );
or ( n31348 , n30783 , n31347 );
and ( n31349 , n30780 , n31348 );
or ( n31350 , n30779 , n31349 );
and ( n31351 , n30776 , n31350 );
or ( n31352 , n30775 , n31351 );
and ( n31353 , n30772 , n31352 );
or ( n31354 , n30771 , n31353 );
and ( n31355 , n30768 , n31354 );
or ( n31356 , n30767 , n31355 );
and ( n31357 , n30764 , n31356 );
or ( n31358 , n30763 , n31357 );
and ( n31359 , n30760 , n31358 );
or ( n31360 , n30759 , n31359 );
and ( n31361 , n30756 , n31360 );
or ( n31362 , n30755 , n31361 );
and ( n31363 , n30752 , n31362 );
or ( n31364 , n30751 , n31363 );
and ( n31365 , n30748 , n31364 );
or ( n31366 , n30747 , n31365 );
and ( n31367 , n30744 , n31366 );
or ( n31368 , n30743 , n31367 );
and ( n31369 , n30740 , n31368 );
or ( n31370 , n30739 , n31369 );
and ( n31371 , n30736 , n31370 );
or ( n31372 , n30735 , n31371 );
and ( n31373 , n30732 , n31372 );
or ( n31374 , n30731 , n31373 );
and ( n31375 , n30728 , n31374 );
or ( n31376 , n30727 , n31375 );
and ( n31377 , n30724 , n31376 );
or ( n31378 , n30723 , n31377 );
and ( n31379 , n30720 , n31378 );
or ( n31380 , n30719 , n31379 );
and ( n31381 , n30716 , n31380 );
or ( n31382 , n30715 , n31381 );
and ( n31383 , n30712 , n31382 );
or ( n31384 , n30711 , n31383 );
and ( n31385 , n30708 , n31384 );
or ( n31386 , n30707 , n31385 );
and ( n31387 , n30704 , n31386 );
or ( n31388 , n30703 , n31387 );
and ( n31389 , n30700 , n31388 );
or ( n31390 , n30699 , n31389 );
and ( n31391 , n30696 , n31390 );
or ( n31392 , n30695 , n31391 );
and ( n31393 , n30692 , n31392 );
or ( n31394 , n30691 , n31393 );
and ( n31395 , n30688 , n31394 );
or ( n31396 , n30687 , n31395 );
and ( n31397 , n30684 , n31396 );
or ( n31398 , n30683 , n31397 );
and ( n31399 , n30680 , n31398 );
or ( n31400 , n30679 , n31399 );
and ( n31401 , n30676 , n31400 );
or ( n31402 , n30675 , n31401 );
and ( n31403 , n30672 , n31402 );
or ( n31404 , n30671 , n31403 );
and ( n31405 , n30668 , n31404 );
or ( n31406 , n30667 , n31405 );
xor ( n31407 , n30664 , n31406 );
buf ( n31408 , n18100 );
and ( n31409 , n29794 , n31408 );
xor ( n31410 , n31407 , n31409 );
xor ( n31411 , n30668 , n31404 );
and ( n31412 , n29799 , n31408 );
and ( n31413 , n31411 , n31412 );
xor ( n31414 , n31411 , n31412 );
xor ( n31415 , n30672 , n31402 );
and ( n31416 , n29804 , n31408 );
and ( n31417 , n31415 , n31416 );
xor ( n31418 , n31415 , n31416 );
xor ( n31419 , n30676 , n31400 );
and ( n31420 , n29809 , n31408 );
and ( n31421 , n31419 , n31420 );
xor ( n31422 , n31419 , n31420 );
xor ( n31423 , n30680 , n31398 );
and ( n31424 , n29814 , n31408 );
and ( n31425 , n31423 , n31424 );
xor ( n31426 , n31423 , n31424 );
xor ( n31427 , n30684 , n31396 );
and ( n31428 , n29819 , n31408 );
and ( n31429 , n31427 , n31428 );
xor ( n31430 , n31427 , n31428 );
xor ( n31431 , n30688 , n31394 );
and ( n31432 , n29824 , n31408 );
and ( n31433 , n31431 , n31432 );
xor ( n31434 , n31431 , n31432 );
xor ( n31435 , n30692 , n31392 );
and ( n31436 , n29829 , n31408 );
and ( n31437 , n31435 , n31436 );
xor ( n31438 , n31435 , n31436 );
xor ( n31439 , n30696 , n31390 );
and ( n31440 , n29834 , n31408 );
and ( n31441 , n31439 , n31440 );
xor ( n31442 , n31439 , n31440 );
xor ( n31443 , n30700 , n31388 );
and ( n31444 , n29839 , n31408 );
and ( n31445 , n31443 , n31444 );
xor ( n31446 , n31443 , n31444 );
xor ( n31447 , n30704 , n31386 );
and ( n31448 , n29844 , n31408 );
and ( n31449 , n31447 , n31448 );
xor ( n31450 , n31447 , n31448 );
xor ( n31451 , n30708 , n31384 );
and ( n31452 , n29849 , n31408 );
and ( n31453 , n31451 , n31452 );
xor ( n31454 , n31451 , n31452 );
xor ( n31455 , n30712 , n31382 );
and ( n31456 , n29854 , n31408 );
and ( n31457 , n31455 , n31456 );
xor ( n31458 , n31455 , n31456 );
xor ( n31459 , n30716 , n31380 );
and ( n31460 , n29859 , n31408 );
and ( n31461 , n31459 , n31460 );
xor ( n31462 , n31459 , n31460 );
xor ( n31463 , n30720 , n31378 );
and ( n31464 , n29864 , n31408 );
and ( n31465 , n31463 , n31464 );
xor ( n31466 , n31463 , n31464 );
xor ( n31467 , n30724 , n31376 );
and ( n31468 , n29869 , n31408 );
and ( n31469 , n31467 , n31468 );
xor ( n31470 , n31467 , n31468 );
xor ( n31471 , n30728 , n31374 );
and ( n31472 , n29874 , n31408 );
and ( n31473 , n31471 , n31472 );
xor ( n31474 , n31471 , n31472 );
xor ( n31475 , n30732 , n31372 );
and ( n31476 , n29879 , n31408 );
and ( n31477 , n31475 , n31476 );
xor ( n31478 , n31475 , n31476 );
xor ( n31479 , n30736 , n31370 );
and ( n31480 , n29884 , n31408 );
and ( n31481 , n31479 , n31480 );
xor ( n31482 , n31479 , n31480 );
xor ( n31483 , n30740 , n31368 );
and ( n31484 , n29889 , n31408 );
and ( n31485 , n31483 , n31484 );
xor ( n31486 , n31483 , n31484 );
xor ( n31487 , n30744 , n31366 );
and ( n31488 , n29894 , n31408 );
and ( n31489 , n31487 , n31488 );
xor ( n31490 , n31487 , n31488 );
xor ( n31491 , n30748 , n31364 );
and ( n31492 , n29899 , n31408 );
and ( n31493 , n31491 , n31492 );
xor ( n31494 , n31491 , n31492 );
xor ( n31495 , n30752 , n31362 );
and ( n31496 , n29904 , n31408 );
and ( n31497 , n31495 , n31496 );
xor ( n31498 , n31495 , n31496 );
xor ( n31499 , n30756 , n31360 );
and ( n31500 , n29909 , n31408 );
and ( n31501 , n31499 , n31500 );
xor ( n31502 , n31499 , n31500 );
xor ( n31503 , n30760 , n31358 );
and ( n31504 , n29914 , n31408 );
and ( n31505 , n31503 , n31504 );
xor ( n31506 , n31503 , n31504 );
xor ( n31507 , n30764 , n31356 );
and ( n31508 , n29919 , n31408 );
and ( n31509 , n31507 , n31508 );
xor ( n31510 , n31507 , n31508 );
xor ( n31511 , n30768 , n31354 );
and ( n31512 , n29924 , n31408 );
and ( n31513 , n31511 , n31512 );
xor ( n31514 , n31511 , n31512 );
xor ( n31515 , n30772 , n31352 );
and ( n31516 , n29929 , n31408 );
and ( n31517 , n31515 , n31516 );
xor ( n31518 , n31515 , n31516 );
xor ( n31519 , n30776 , n31350 );
and ( n31520 , n29934 , n31408 );
and ( n31521 , n31519 , n31520 );
xor ( n31522 , n31519 , n31520 );
xor ( n31523 , n30780 , n31348 );
and ( n31524 , n29939 , n31408 );
and ( n31525 , n31523 , n31524 );
xor ( n31526 , n31523 , n31524 );
xor ( n31527 , n30784 , n31346 );
and ( n31528 , n29944 , n31408 );
and ( n31529 , n31527 , n31528 );
xor ( n31530 , n31527 , n31528 );
xor ( n31531 , n30788 , n31344 );
and ( n31532 , n29949 , n31408 );
and ( n31533 , n31531 , n31532 );
xor ( n31534 , n31531 , n31532 );
xor ( n31535 , n30792 , n31342 );
and ( n31536 , n29954 , n31408 );
and ( n31537 , n31535 , n31536 );
xor ( n31538 , n31535 , n31536 );
xor ( n31539 , n30796 , n31340 );
and ( n31540 , n29959 , n31408 );
and ( n31541 , n31539 , n31540 );
xor ( n31542 , n31539 , n31540 );
xor ( n31543 , n30800 , n31338 );
and ( n31544 , n29964 , n31408 );
and ( n31545 , n31543 , n31544 );
xor ( n31546 , n31543 , n31544 );
xor ( n31547 , n30804 , n31336 );
and ( n31548 , n29969 , n31408 );
and ( n31549 , n31547 , n31548 );
xor ( n31550 , n31547 , n31548 );
xor ( n31551 , n30808 , n31334 );
and ( n31552 , n29974 , n31408 );
and ( n31553 , n31551 , n31552 );
xor ( n31554 , n31551 , n31552 );
xor ( n31555 , n30812 , n31332 );
and ( n31556 , n29979 , n31408 );
and ( n31557 , n31555 , n31556 );
xor ( n31558 , n31555 , n31556 );
xor ( n31559 , n30816 , n31330 );
and ( n31560 , n29984 , n31408 );
and ( n31561 , n31559 , n31560 );
xor ( n31562 , n31559 , n31560 );
xor ( n31563 , n30820 , n31328 );
and ( n31564 , n29989 , n31408 );
and ( n31565 , n31563 , n31564 );
xor ( n31566 , n31563 , n31564 );
xor ( n31567 , n30824 , n31326 );
and ( n31568 , n29994 , n31408 );
and ( n31569 , n31567 , n31568 );
xor ( n31570 , n31567 , n31568 );
xor ( n31571 , n30828 , n31324 );
and ( n31572 , n29999 , n31408 );
and ( n31573 , n31571 , n31572 );
xor ( n31574 , n31571 , n31572 );
xor ( n31575 , n30832 , n31322 );
and ( n31576 , n30004 , n31408 );
and ( n31577 , n31575 , n31576 );
xor ( n31578 , n31575 , n31576 );
xor ( n31579 , n30836 , n31320 );
and ( n31580 , n30009 , n31408 );
and ( n31581 , n31579 , n31580 );
xor ( n31582 , n31579 , n31580 );
xor ( n31583 , n30840 , n31318 );
and ( n31584 , n30014 , n31408 );
and ( n31585 , n31583 , n31584 );
xor ( n31586 , n31583 , n31584 );
xor ( n31587 , n30844 , n31316 );
and ( n31588 , n30019 , n31408 );
and ( n31589 , n31587 , n31588 );
xor ( n31590 , n31587 , n31588 );
xor ( n31591 , n30848 , n31314 );
and ( n31592 , n30024 , n31408 );
and ( n31593 , n31591 , n31592 );
xor ( n31594 , n31591 , n31592 );
xor ( n31595 , n30852 , n31312 );
and ( n31596 , n30029 , n31408 );
and ( n31597 , n31595 , n31596 );
xor ( n31598 , n31595 , n31596 );
xor ( n31599 , n30856 , n31310 );
and ( n31600 , n30034 , n31408 );
and ( n31601 , n31599 , n31600 );
xor ( n31602 , n31599 , n31600 );
xor ( n31603 , n30860 , n31308 );
and ( n31604 , n30039 , n31408 );
and ( n31605 , n31603 , n31604 );
xor ( n31606 , n31603 , n31604 );
xor ( n31607 , n30864 , n31306 );
and ( n31608 , n30044 , n31408 );
and ( n31609 , n31607 , n31608 );
xor ( n31610 , n31607 , n31608 );
xor ( n31611 , n30868 , n31304 );
and ( n31612 , n30049 , n31408 );
and ( n31613 , n31611 , n31612 );
xor ( n31614 , n31611 , n31612 );
xor ( n31615 , n30872 , n31302 );
and ( n31616 , n30054 , n31408 );
and ( n31617 , n31615 , n31616 );
xor ( n31618 , n31615 , n31616 );
xor ( n31619 , n30876 , n31300 );
and ( n31620 , n30059 , n31408 );
and ( n31621 , n31619 , n31620 );
xor ( n31622 , n31619 , n31620 );
xor ( n31623 , n30880 , n31298 );
and ( n31624 , n30064 , n31408 );
and ( n31625 , n31623 , n31624 );
xor ( n31626 , n31623 , n31624 );
xor ( n31627 , n30884 , n31296 );
and ( n31628 , n30069 , n31408 );
and ( n31629 , n31627 , n31628 );
xor ( n31630 , n31627 , n31628 );
xor ( n31631 , n30888 , n31294 );
and ( n31632 , n30074 , n31408 );
and ( n31633 , n31631 , n31632 );
xor ( n31634 , n31631 , n31632 );
xor ( n31635 , n30892 , n31292 );
and ( n31636 , n30079 , n31408 );
and ( n31637 , n31635 , n31636 );
xor ( n31638 , n31635 , n31636 );
xor ( n31639 , n30896 , n31290 );
and ( n31640 , n30084 , n31408 );
and ( n31641 , n31639 , n31640 );
xor ( n31642 , n31639 , n31640 );
xor ( n31643 , n30900 , n31288 );
and ( n31644 , n30089 , n31408 );
and ( n31645 , n31643 , n31644 );
xor ( n31646 , n31643 , n31644 );
xor ( n31647 , n30904 , n31286 );
and ( n31648 , n30094 , n31408 );
and ( n31649 , n31647 , n31648 );
xor ( n31650 , n31647 , n31648 );
xor ( n31651 , n30908 , n31284 );
and ( n31652 , n30099 , n31408 );
and ( n31653 , n31651 , n31652 );
xor ( n31654 , n31651 , n31652 );
xor ( n31655 , n30912 , n31282 );
and ( n31656 , n30104 , n31408 );
and ( n31657 , n31655 , n31656 );
xor ( n31658 , n31655 , n31656 );
xor ( n31659 , n30916 , n31280 );
and ( n31660 , n30109 , n31408 );
and ( n31661 , n31659 , n31660 );
xor ( n31662 , n31659 , n31660 );
xor ( n31663 , n30920 , n31278 );
and ( n31664 , n30114 , n31408 );
and ( n31665 , n31663 , n31664 );
xor ( n31666 , n31663 , n31664 );
xor ( n31667 , n30924 , n31276 );
and ( n31668 , n30119 , n31408 );
and ( n31669 , n31667 , n31668 );
xor ( n31670 , n31667 , n31668 );
xor ( n31671 , n30928 , n31274 );
and ( n31672 , n30124 , n31408 );
and ( n31673 , n31671 , n31672 );
xor ( n31674 , n31671 , n31672 );
xor ( n31675 , n30932 , n31272 );
and ( n31676 , n30129 , n31408 );
and ( n31677 , n31675 , n31676 );
xor ( n31678 , n31675 , n31676 );
xor ( n31679 , n30936 , n31270 );
and ( n31680 , n30134 , n31408 );
and ( n31681 , n31679 , n31680 );
xor ( n31682 , n31679 , n31680 );
xor ( n31683 , n30940 , n31268 );
and ( n31684 , n30139 , n31408 );
and ( n31685 , n31683 , n31684 );
xor ( n31686 , n31683 , n31684 );
xor ( n31687 , n30944 , n31266 );
and ( n31688 , n30144 , n31408 );
and ( n31689 , n31687 , n31688 );
xor ( n31690 , n31687 , n31688 );
xor ( n31691 , n30948 , n31264 );
and ( n31692 , n30149 , n31408 );
and ( n31693 , n31691 , n31692 );
xor ( n31694 , n31691 , n31692 );
xor ( n31695 , n30952 , n31262 );
and ( n31696 , n30154 , n31408 );
and ( n31697 , n31695 , n31696 );
xor ( n31698 , n31695 , n31696 );
xor ( n31699 , n30956 , n31260 );
and ( n31700 , n30159 , n31408 );
and ( n31701 , n31699 , n31700 );
xor ( n31702 , n31699 , n31700 );
xor ( n31703 , n30960 , n31258 );
and ( n31704 , n30164 , n31408 );
and ( n31705 , n31703 , n31704 );
xor ( n31706 , n31703 , n31704 );
xor ( n31707 , n30964 , n31256 );
and ( n31708 , n30169 , n31408 );
and ( n31709 , n31707 , n31708 );
xor ( n31710 , n31707 , n31708 );
xor ( n31711 , n30968 , n31254 );
and ( n31712 , n30174 , n31408 );
and ( n31713 , n31711 , n31712 );
xor ( n31714 , n31711 , n31712 );
xor ( n31715 , n30972 , n31252 );
and ( n31716 , n30179 , n31408 );
and ( n31717 , n31715 , n31716 );
xor ( n31718 , n31715 , n31716 );
xor ( n31719 , n30976 , n31250 );
and ( n31720 , n30184 , n31408 );
and ( n31721 , n31719 , n31720 );
xor ( n31722 , n31719 , n31720 );
xor ( n31723 , n30980 , n31248 );
and ( n31724 , n30189 , n31408 );
and ( n31725 , n31723 , n31724 );
xor ( n31726 , n31723 , n31724 );
xor ( n31727 , n30984 , n31246 );
and ( n31728 , n30194 , n31408 );
and ( n31729 , n31727 , n31728 );
xor ( n31730 , n31727 , n31728 );
xor ( n31731 , n30988 , n31244 );
and ( n31732 , n30199 , n31408 );
and ( n31733 , n31731 , n31732 );
xor ( n31734 , n31731 , n31732 );
xor ( n31735 , n30992 , n31242 );
and ( n31736 , n30204 , n31408 );
and ( n31737 , n31735 , n31736 );
xor ( n31738 , n31735 , n31736 );
xor ( n31739 , n30996 , n31240 );
and ( n31740 , n30209 , n31408 );
and ( n31741 , n31739 , n31740 );
xor ( n31742 , n31739 , n31740 );
xor ( n31743 , n31000 , n31238 );
and ( n31744 , n30214 , n31408 );
and ( n31745 , n31743 , n31744 );
xor ( n31746 , n31743 , n31744 );
xor ( n31747 , n31004 , n31236 );
and ( n31748 , n30219 , n31408 );
and ( n31749 , n31747 , n31748 );
xor ( n31750 , n31747 , n31748 );
xor ( n31751 , n31008 , n31234 );
and ( n31752 , n30224 , n31408 );
and ( n31753 , n31751 , n31752 );
xor ( n31754 , n31751 , n31752 );
xor ( n31755 , n31012 , n31232 );
and ( n31756 , n30229 , n31408 );
and ( n31757 , n31755 , n31756 );
xor ( n31758 , n31755 , n31756 );
xor ( n31759 , n31016 , n31230 );
and ( n31760 , n30234 , n31408 );
and ( n31761 , n31759 , n31760 );
xor ( n31762 , n31759 , n31760 );
xor ( n31763 , n31020 , n31228 );
and ( n31764 , n30239 , n31408 );
and ( n31765 , n31763 , n31764 );
xor ( n31766 , n31763 , n31764 );
xor ( n31767 , n31024 , n31226 );
and ( n31768 , n30244 , n31408 );
and ( n31769 , n31767 , n31768 );
xor ( n31770 , n31767 , n31768 );
xor ( n31771 , n31028 , n31224 );
and ( n31772 , n30249 , n31408 );
and ( n31773 , n31771 , n31772 );
xor ( n31774 , n31771 , n31772 );
xor ( n31775 , n31032 , n31222 );
and ( n31776 , n30254 , n31408 );
and ( n31777 , n31775 , n31776 );
xor ( n31778 , n31775 , n31776 );
xor ( n31779 , n31036 , n31220 );
and ( n31780 , n30259 , n31408 );
and ( n31781 , n31779 , n31780 );
xor ( n31782 , n31779 , n31780 );
xor ( n31783 , n31040 , n31218 );
and ( n31784 , n30264 , n31408 );
and ( n31785 , n31783 , n31784 );
xor ( n31786 , n31783 , n31784 );
xor ( n31787 , n31044 , n31216 );
and ( n31788 , n30269 , n31408 );
and ( n31789 , n31787 , n31788 );
xor ( n31790 , n31787 , n31788 );
xor ( n31791 , n31048 , n31214 );
and ( n31792 , n30274 , n31408 );
and ( n31793 , n31791 , n31792 );
xor ( n31794 , n31791 , n31792 );
xor ( n31795 , n31052 , n31212 );
and ( n31796 , n30279 , n31408 );
and ( n31797 , n31795 , n31796 );
xor ( n31798 , n31795 , n31796 );
xor ( n31799 , n31056 , n31210 );
and ( n31800 , n30284 , n31408 );
and ( n31801 , n31799 , n31800 );
xor ( n31802 , n31799 , n31800 );
xor ( n31803 , n31060 , n31208 );
and ( n31804 , n30289 , n31408 );
and ( n31805 , n31803 , n31804 );
xor ( n31806 , n31803 , n31804 );
xor ( n31807 , n31064 , n31206 );
and ( n31808 , n30294 , n31408 );
and ( n31809 , n31807 , n31808 );
xor ( n31810 , n31807 , n31808 );
xor ( n31811 , n31068 , n31204 );
and ( n31812 , n30299 , n31408 );
and ( n31813 , n31811 , n31812 );
xor ( n31814 , n31811 , n31812 );
xor ( n31815 , n31072 , n31202 );
and ( n31816 , n30304 , n31408 );
and ( n31817 , n31815 , n31816 );
xor ( n31818 , n31815 , n31816 );
xor ( n31819 , n31076 , n31200 );
and ( n31820 , n30309 , n31408 );
and ( n31821 , n31819 , n31820 );
xor ( n31822 , n31819 , n31820 );
xor ( n31823 , n31080 , n31198 );
and ( n31824 , n30314 , n31408 );
and ( n31825 , n31823 , n31824 );
xor ( n31826 , n31823 , n31824 );
xor ( n31827 , n31084 , n31196 );
and ( n31828 , n30319 , n31408 );
and ( n31829 , n31827 , n31828 );
xor ( n31830 , n31827 , n31828 );
xor ( n31831 , n31088 , n31194 );
and ( n31832 , n30324 , n31408 );
and ( n31833 , n31831 , n31832 );
xor ( n31834 , n31831 , n31832 );
xor ( n31835 , n31092 , n31192 );
and ( n31836 , n30329 , n31408 );
and ( n31837 , n31835 , n31836 );
xor ( n31838 , n31835 , n31836 );
xor ( n31839 , n31096 , n31190 );
and ( n31840 , n30334 , n31408 );
and ( n31841 , n31839 , n31840 );
xor ( n31842 , n31839 , n31840 );
xor ( n31843 , n31100 , n31188 );
and ( n31844 , n30339 , n31408 );
and ( n31845 , n31843 , n31844 );
xor ( n31846 , n31843 , n31844 );
xor ( n31847 , n31104 , n31186 );
and ( n31848 , n30344 , n31408 );
and ( n31849 , n31847 , n31848 );
xor ( n31850 , n31847 , n31848 );
xor ( n31851 , n31108 , n31184 );
and ( n31852 , n30349 , n31408 );
and ( n31853 , n31851 , n31852 );
xor ( n31854 , n31851 , n31852 );
xor ( n31855 , n31112 , n31182 );
and ( n31856 , n30354 , n31408 );
and ( n31857 , n31855 , n31856 );
xor ( n31858 , n31855 , n31856 );
xor ( n31859 , n31116 , n31180 );
and ( n31860 , n30359 , n31408 );
and ( n31861 , n31859 , n31860 );
xor ( n31862 , n31859 , n31860 );
xor ( n31863 , n31120 , n31178 );
and ( n31864 , n30364 , n31408 );
and ( n31865 , n31863 , n31864 );
xor ( n31866 , n31863 , n31864 );
xor ( n31867 , n31124 , n31176 );
and ( n31868 , n30369 , n31408 );
and ( n31869 , n31867 , n31868 );
xor ( n31870 , n31867 , n31868 );
xor ( n31871 , n31128 , n31174 );
and ( n31872 , n30374 , n31408 );
and ( n31873 , n31871 , n31872 );
xor ( n31874 , n31871 , n31872 );
xor ( n31875 , n31132 , n31172 );
and ( n31876 , n30379 , n31408 );
and ( n31877 , n31875 , n31876 );
xor ( n31878 , n31875 , n31876 );
xor ( n31879 , n31136 , n31170 );
and ( n31880 , n30384 , n31408 );
and ( n31881 , n31879 , n31880 );
xor ( n31882 , n31879 , n31880 );
xor ( n31883 , n31140 , n31168 );
and ( n31884 , n30389 , n31408 );
and ( n31885 , n31883 , n31884 );
xor ( n31886 , n31883 , n31884 );
xor ( n31887 , n31144 , n31166 );
and ( n31888 , n30394 , n31408 );
and ( n31889 , n31887 , n31888 );
xor ( n31890 , n31887 , n31888 );
xor ( n31891 , n31148 , n31164 );
and ( n31892 , n30399 , n31408 );
and ( n31893 , n31891 , n31892 );
xor ( n31894 , n31891 , n31892 );
xor ( n31895 , n31152 , n31162 );
and ( n31896 , n30404 , n31408 );
and ( n31897 , n31895 , n31896 );
xor ( n31898 , n31895 , n31896 );
xor ( n31899 , n31156 , n31160 );
and ( n31900 , n30409 , n31408 );
and ( n31901 , n31899 , n31900 );
buf ( n31902 , n31901 );
and ( n31903 , n31898 , n31902 );
or ( n31904 , n31897 , n31903 );
and ( n31905 , n31894 , n31904 );
or ( n31906 , n31893 , n31905 );
and ( n31907 , n31890 , n31906 );
or ( n31908 , n31889 , n31907 );
and ( n31909 , n31886 , n31908 );
or ( n31910 , n31885 , n31909 );
and ( n31911 , n31882 , n31910 );
or ( n31912 , n31881 , n31911 );
and ( n31913 , n31878 , n31912 );
or ( n31914 , n31877 , n31913 );
and ( n31915 , n31874 , n31914 );
or ( n31916 , n31873 , n31915 );
and ( n31917 , n31870 , n31916 );
or ( n31918 , n31869 , n31917 );
and ( n31919 , n31866 , n31918 );
or ( n31920 , n31865 , n31919 );
and ( n31921 , n31862 , n31920 );
or ( n31922 , n31861 , n31921 );
and ( n31923 , n31858 , n31922 );
or ( n31924 , n31857 , n31923 );
and ( n31925 , n31854 , n31924 );
or ( n31926 , n31853 , n31925 );
and ( n31927 , n31850 , n31926 );
or ( n31928 , n31849 , n31927 );
and ( n31929 , n31846 , n31928 );
or ( n31930 , n31845 , n31929 );
and ( n31931 , n31842 , n31930 );
or ( n31932 , n31841 , n31931 );
and ( n31933 , n31838 , n31932 );
or ( n31934 , n31837 , n31933 );
and ( n31935 , n31834 , n31934 );
or ( n31936 , n31833 , n31935 );
and ( n31937 , n31830 , n31936 );
or ( n31938 , n31829 , n31937 );
and ( n31939 , n31826 , n31938 );
or ( n31940 , n31825 , n31939 );
and ( n31941 , n31822 , n31940 );
or ( n31942 , n31821 , n31941 );
and ( n31943 , n31818 , n31942 );
or ( n31944 , n31817 , n31943 );
and ( n31945 , n31814 , n31944 );
or ( n31946 , n31813 , n31945 );
and ( n31947 , n31810 , n31946 );
or ( n31948 , n31809 , n31947 );
and ( n31949 , n31806 , n31948 );
or ( n31950 , n31805 , n31949 );
and ( n31951 , n31802 , n31950 );
or ( n31952 , n31801 , n31951 );
and ( n31953 , n31798 , n31952 );
or ( n31954 , n31797 , n31953 );
and ( n31955 , n31794 , n31954 );
or ( n31956 , n31793 , n31955 );
and ( n31957 , n31790 , n31956 );
or ( n31958 , n31789 , n31957 );
and ( n31959 , n31786 , n31958 );
or ( n31960 , n31785 , n31959 );
and ( n31961 , n31782 , n31960 );
or ( n31962 , n31781 , n31961 );
and ( n31963 , n31778 , n31962 );
or ( n31964 , n31777 , n31963 );
and ( n31965 , n31774 , n31964 );
or ( n31966 , n31773 , n31965 );
and ( n31967 , n31770 , n31966 );
or ( n31968 , n31769 , n31967 );
and ( n31969 , n31766 , n31968 );
or ( n31970 , n31765 , n31969 );
and ( n31971 , n31762 , n31970 );
or ( n31972 , n31761 , n31971 );
and ( n31973 , n31758 , n31972 );
or ( n31974 , n31757 , n31973 );
and ( n31975 , n31754 , n31974 );
or ( n31976 , n31753 , n31975 );
and ( n31977 , n31750 , n31976 );
or ( n31978 , n31749 , n31977 );
and ( n31979 , n31746 , n31978 );
or ( n31980 , n31745 , n31979 );
and ( n31981 , n31742 , n31980 );
or ( n31982 , n31741 , n31981 );
and ( n31983 , n31738 , n31982 );
or ( n31984 , n31737 , n31983 );
and ( n31985 , n31734 , n31984 );
or ( n31986 , n31733 , n31985 );
and ( n31987 , n31730 , n31986 );
or ( n31988 , n31729 , n31987 );
and ( n31989 , n31726 , n31988 );
or ( n31990 , n31725 , n31989 );
and ( n31991 , n31722 , n31990 );
or ( n31992 , n31721 , n31991 );
and ( n31993 , n31718 , n31992 );
or ( n31994 , n31717 , n31993 );
and ( n31995 , n31714 , n31994 );
or ( n31996 , n31713 , n31995 );
and ( n31997 , n31710 , n31996 );
or ( n31998 , n31709 , n31997 );
and ( n31999 , n31706 , n31998 );
or ( n32000 , n31705 , n31999 );
and ( n32001 , n31702 , n32000 );
or ( n32002 , n31701 , n32001 );
and ( n32003 , n31698 , n32002 );
or ( n32004 , n31697 , n32003 );
and ( n32005 , n31694 , n32004 );
or ( n32006 , n31693 , n32005 );
and ( n32007 , n31690 , n32006 );
or ( n32008 , n31689 , n32007 );
and ( n32009 , n31686 , n32008 );
or ( n32010 , n31685 , n32009 );
and ( n32011 , n31682 , n32010 );
or ( n32012 , n31681 , n32011 );
and ( n32013 , n31678 , n32012 );
or ( n32014 , n31677 , n32013 );
and ( n32015 , n31674 , n32014 );
or ( n32016 , n31673 , n32015 );
and ( n32017 , n31670 , n32016 );
or ( n32018 , n31669 , n32017 );
and ( n32019 , n31666 , n32018 );
or ( n32020 , n31665 , n32019 );
and ( n32021 , n31662 , n32020 );
or ( n32022 , n31661 , n32021 );
and ( n32023 , n31658 , n32022 );
or ( n32024 , n31657 , n32023 );
and ( n32025 , n31654 , n32024 );
or ( n32026 , n31653 , n32025 );
and ( n32027 , n31650 , n32026 );
or ( n32028 , n31649 , n32027 );
and ( n32029 , n31646 , n32028 );
or ( n32030 , n31645 , n32029 );
and ( n32031 , n31642 , n32030 );
or ( n32032 , n31641 , n32031 );
and ( n32033 , n31638 , n32032 );
or ( n32034 , n31637 , n32033 );
and ( n32035 , n31634 , n32034 );
or ( n32036 , n31633 , n32035 );
and ( n32037 , n31630 , n32036 );
or ( n32038 , n31629 , n32037 );
and ( n32039 , n31626 , n32038 );
or ( n32040 , n31625 , n32039 );
and ( n32041 , n31622 , n32040 );
or ( n32042 , n31621 , n32041 );
and ( n32043 , n31618 , n32042 );
or ( n32044 , n31617 , n32043 );
and ( n32045 , n31614 , n32044 );
or ( n32046 , n31613 , n32045 );
and ( n32047 , n31610 , n32046 );
or ( n32048 , n31609 , n32047 );
and ( n32049 , n31606 , n32048 );
or ( n32050 , n31605 , n32049 );
and ( n32051 , n31602 , n32050 );
or ( n32052 , n31601 , n32051 );
and ( n32053 , n31598 , n32052 );
or ( n32054 , n31597 , n32053 );
and ( n32055 , n31594 , n32054 );
or ( n32056 , n31593 , n32055 );
and ( n32057 , n31590 , n32056 );
or ( n32058 , n31589 , n32057 );
and ( n32059 , n31586 , n32058 );
or ( n32060 , n31585 , n32059 );
and ( n32061 , n31582 , n32060 );
or ( n32062 , n31581 , n32061 );
and ( n32063 , n31578 , n32062 );
or ( n32064 , n31577 , n32063 );
and ( n32065 , n31574 , n32064 );
or ( n32066 , n31573 , n32065 );
and ( n32067 , n31570 , n32066 );
or ( n32068 , n31569 , n32067 );
and ( n32069 , n31566 , n32068 );
or ( n32070 , n31565 , n32069 );
and ( n32071 , n31562 , n32070 );
or ( n32072 , n31561 , n32071 );
and ( n32073 , n31558 , n32072 );
or ( n32074 , n31557 , n32073 );
and ( n32075 , n31554 , n32074 );
or ( n32076 , n31553 , n32075 );
and ( n32077 , n31550 , n32076 );
or ( n32078 , n31549 , n32077 );
and ( n32079 , n31546 , n32078 );
or ( n32080 , n31545 , n32079 );
and ( n32081 , n31542 , n32080 );
or ( n32082 , n31541 , n32081 );
and ( n32083 , n31538 , n32082 );
or ( n32084 , n31537 , n32083 );
and ( n32085 , n31534 , n32084 );
or ( n32086 , n31533 , n32085 );
and ( n32087 , n31530 , n32086 );
or ( n32088 , n31529 , n32087 );
and ( n32089 , n31526 , n32088 );
or ( n32090 , n31525 , n32089 );
and ( n32091 , n31522 , n32090 );
or ( n32092 , n31521 , n32091 );
and ( n32093 , n31518 , n32092 );
or ( n32094 , n31517 , n32093 );
and ( n32095 , n31514 , n32094 );
or ( n32096 , n31513 , n32095 );
and ( n32097 , n31510 , n32096 );
or ( n32098 , n31509 , n32097 );
and ( n32099 , n31506 , n32098 );
or ( n32100 , n31505 , n32099 );
and ( n32101 , n31502 , n32100 );
or ( n32102 , n31501 , n32101 );
and ( n32103 , n31498 , n32102 );
or ( n32104 , n31497 , n32103 );
and ( n32105 , n31494 , n32104 );
or ( n32106 , n31493 , n32105 );
and ( n32107 , n31490 , n32106 );
or ( n32108 , n31489 , n32107 );
and ( n32109 , n31486 , n32108 );
or ( n32110 , n31485 , n32109 );
and ( n32111 , n31482 , n32110 );
or ( n32112 , n31481 , n32111 );
and ( n32113 , n31478 , n32112 );
or ( n32114 , n31477 , n32113 );
and ( n32115 , n31474 , n32114 );
or ( n32116 , n31473 , n32115 );
and ( n32117 , n31470 , n32116 );
or ( n32118 , n31469 , n32117 );
and ( n32119 , n31466 , n32118 );
or ( n32120 , n31465 , n32119 );
and ( n32121 , n31462 , n32120 );
or ( n32122 , n31461 , n32121 );
and ( n32123 , n31458 , n32122 );
or ( n32124 , n31457 , n32123 );
and ( n32125 , n31454 , n32124 );
or ( n32126 , n31453 , n32125 );
and ( n32127 , n31450 , n32126 );
or ( n32128 , n31449 , n32127 );
and ( n32129 , n31446 , n32128 );
or ( n32130 , n31445 , n32129 );
and ( n32131 , n31442 , n32130 );
or ( n32132 , n31441 , n32131 );
and ( n32133 , n31438 , n32132 );
or ( n32134 , n31437 , n32133 );
and ( n32135 , n31434 , n32134 );
or ( n32136 , n31433 , n32135 );
and ( n32137 , n31430 , n32136 );
or ( n32138 , n31429 , n32137 );
and ( n32139 , n31426 , n32138 );
or ( n32140 , n31425 , n32139 );
and ( n32141 , n31422 , n32140 );
or ( n32142 , n31421 , n32141 );
and ( n32143 , n31418 , n32142 );
or ( n32144 , n31417 , n32143 );
and ( n32145 , n31414 , n32144 );
or ( n32146 , n31413 , n32145 );
xor ( n32147 , n31410 , n32146 );
buf ( n32148 , n18098 );
and ( n32149 , n29799 , n32148 );
xor ( n32150 , n32147 , n32149 );
xor ( n32151 , n31414 , n32144 );
and ( n32152 , n29804 , n32148 );
and ( n32153 , n32151 , n32152 );
xor ( n32154 , n32151 , n32152 );
xor ( n32155 , n31418 , n32142 );
and ( n32156 , n29809 , n32148 );
and ( n32157 , n32155 , n32156 );
xor ( n32158 , n32155 , n32156 );
xor ( n32159 , n31422 , n32140 );
and ( n32160 , n29814 , n32148 );
and ( n32161 , n32159 , n32160 );
xor ( n32162 , n32159 , n32160 );
xor ( n32163 , n31426 , n32138 );
and ( n32164 , n29819 , n32148 );
and ( n32165 , n32163 , n32164 );
xor ( n32166 , n32163 , n32164 );
xor ( n32167 , n31430 , n32136 );
and ( n32168 , n29824 , n32148 );
and ( n32169 , n32167 , n32168 );
xor ( n32170 , n32167 , n32168 );
xor ( n32171 , n31434 , n32134 );
and ( n32172 , n29829 , n32148 );
and ( n32173 , n32171 , n32172 );
xor ( n32174 , n32171 , n32172 );
xor ( n32175 , n31438 , n32132 );
and ( n32176 , n29834 , n32148 );
and ( n32177 , n32175 , n32176 );
xor ( n32178 , n32175 , n32176 );
xor ( n32179 , n31442 , n32130 );
and ( n32180 , n29839 , n32148 );
and ( n32181 , n32179 , n32180 );
xor ( n32182 , n32179 , n32180 );
xor ( n32183 , n31446 , n32128 );
and ( n32184 , n29844 , n32148 );
and ( n32185 , n32183 , n32184 );
xor ( n32186 , n32183 , n32184 );
xor ( n32187 , n31450 , n32126 );
and ( n32188 , n29849 , n32148 );
and ( n32189 , n32187 , n32188 );
xor ( n32190 , n32187 , n32188 );
xor ( n32191 , n31454 , n32124 );
and ( n32192 , n29854 , n32148 );
and ( n32193 , n32191 , n32192 );
xor ( n32194 , n32191 , n32192 );
xor ( n32195 , n31458 , n32122 );
and ( n32196 , n29859 , n32148 );
and ( n32197 , n32195 , n32196 );
xor ( n32198 , n32195 , n32196 );
xor ( n32199 , n31462 , n32120 );
and ( n32200 , n29864 , n32148 );
and ( n32201 , n32199 , n32200 );
xor ( n32202 , n32199 , n32200 );
xor ( n32203 , n31466 , n32118 );
and ( n32204 , n29869 , n32148 );
and ( n32205 , n32203 , n32204 );
xor ( n32206 , n32203 , n32204 );
xor ( n32207 , n31470 , n32116 );
and ( n32208 , n29874 , n32148 );
and ( n32209 , n32207 , n32208 );
xor ( n32210 , n32207 , n32208 );
xor ( n32211 , n31474 , n32114 );
and ( n32212 , n29879 , n32148 );
and ( n32213 , n32211 , n32212 );
xor ( n32214 , n32211 , n32212 );
xor ( n32215 , n31478 , n32112 );
and ( n32216 , n29884 , n32148 );
and ( n32217 , n32215 , n32216 );
xor ( n32218 , n32215 , n32216 );
xor ( n32219 , n31482 , n32110 );
and ( n32220 , n29889 , n32148 );
and ( n32221 , n32219 , n32220 );
xor ( n32222 , n32219 , n32220 );
xor ( n32223 , n31486 , n32108 );
and ( n32224 , n29894 , n32148 );
and ( n32225 , n32223 , n32224 );
xor ( n32226 , n32223 , n32224 );
xor ( n32227 , n31490 , n32106 );
and ( n32228 , n29899 , n32148 );
and ( n32229 , n32227 , n32228 );
xor ( n32230 , n32227 , n32228 );
xor ( n32231 , n31494 , n32104 );
and ( n32232 , n29904 , n32148 );
and ( n32233 , n32231 , n32232 );
xor ( n32234 , n32231 , n32232 );
xor ( n32235 , n31498 , n32102 );
and ( n32236 , n29909 , n32148 );
and ( n32237 , n32235 , n32236 );
xor ( n32238 , n32235 , n32236 );
xor ( n32239 , n31502 , n32100 );
and ( n32240 , n29914 , n32148 );
and ( n32241 , n32239 , n32240 );
xor ( n32242 , n32239 , n32240 );
xor ( n32243 , n31506 , n32098 );
and ( n32244 , n29919 , n32148 );
and ( n32245 , n32243 , n32244 );
xor ( n32246 , n32243 , n32244 );
xor ( n32247 , n31510 , n32096 );
and ( n32248 , n29924 , n32148 );
and ( n32249 , n32247 , n32248 );
xor ( n32250 , n32247 , n32248 );
xor ( n32251 , n31514 , n32094 );
and ( n32252 , n29929 , n32148 );
and ( n32253 , n32251 , n32252 );
xor ( n32254 , n32251 , n32252 );
xor ( n32255 , n31518 , n32092 );
and ( n32256 , n29934 , n32148 );
and ( n32257 , n32255 , n32256 );
xor ( n32258 , n32255 , n32256 );
xor ( n32259 , n31522 , n32090 );
and ( n32260 , n29939 , n32148 );
and ( n32261 , n32259 , n32260 );
xor ( n32262 , n32259 , n32260 );
xor ( n32263 , n31526 , n32088 );
and ( n32264 , n29944 , n32148 );
and ( n32265 , n32263 , n32264 );
xor ( n32266 , n32263 , n32264 );
xor ( n32267 , n31530 , n32086 );
and ( n32268 , n29949 , n32148 );
and ( n32269 , n32267 , n32268 );
xor ( n32270 , n32267 , n32268 );
xor ( n32271 , n31534 , n32084 );
and ( n32272 , n29954 , n32148 );
and ( n32273 , n32271 , n32272 );
xor ( n32274 , n32271 , n32272 );
xor ( n32275 , n31538 , n32082 );
and ( n32276 , n29959 , n32148 );
and ( n32277 , n32275 , n32276 );
xor ( n32278 , n32275 , n32276 );
xor ( n32279 , n31542 , n32080 );
and ( n32280 , n29964 , n32148 );
and ( n32281 , n32279 , n32280 );
xor ( n32282 , n32279 , n32280 );
xor ( n32283 , n31546 , n32078 );
and ( n32284 , n29969 , n32148 );
and ( n32285 , n32283 , n32284 );
xor ( n32286 , n32283 , n32284 );
xor ( n32287 , n31550 , n32076 );
and ( n32288 , n29974 , n32148 );
and ( n32289 , n32287 , n32288 );
xor ( n32290 , n32287 , n32288 );
xor ( n32291 , n31554 , n32074 );
and ( n32292 , n29979 , n32148 );
and ( n32293 , n32291 , n32292 );
xor ( n32294 , n32291 , n32292 );
xor ( n32295 , n31558 , n32072 );
and ( n32296 , n29984 , n32148 );
and ( n32297 , n32295 , n32296 );
xor ( n32298 , n32295 , n32296 );
xor ( n32299 , n31562 , n32070 );
and ( n32300 , n29989 , n32148 );
and ( n32301 , n32299 , n32300 );
xor ( n32302 , n32299 , n32300 );
xor ( n32303 , n31566 , n32068 );
and ( n32304 , n29994 , n32148 );
and ( n32305 , n32303 , n32304 );
xor ( n32306 , n32303 , n32304 );
xor ( n32307 , n31570 , n32066 );
and ( n32308 , n29999 , n32148 );
and ( n32309 , n32307 , n32308 );
xor ( n32310 , n32307 , n32308 );
xor ( n32311 , n31574 , n32064 );
and ( n32312 , n30004 , n32148 );
and ( n32313 , n32311 , n32312 );
xor ( n32314 , n32311 , n32312 );
xor ( n32315 , n31578 , n32062 );
and ( n32316 , n30009 , n32148 );
and ( n32317 , n32315 , n32316 );
xor ( n32318 , n32315 , n32316 );
xor ( n32319 , n31582 , n32060 );
and ( n32320 , n30014 , n32148 );
and ( n32321 , n32319 , n32320 );
xor ( n32322 , n32319 , n32320 );
xor ( n32323 , n31586 , n32058 );
and ( n32324 , n30019 , n32148 );
and ( n32325 , n32323 , n32324 );
xor ( n32326 , n32323 , n32324 );
xor ( n32327 , n31590 , n32056 );
and ( n32328 , n30024 , n32148 );
and ( n32329 , n32327 , n32328 );
xor ( n32330 , n32327 , n32328 );
xor ( n32331 , n31594 , n32054 );
and ( n32332 , n30029 , n32148 );
and ( n32333 , n32331 , n32332 );
xor ( n32334 , n32331 , n32332 );
xor ( n32335 , n31598 , n32052 );
and ( n32336 , n30034 , n32148 );
and ( n32337 , n32335 , n32336 );
xor ( n32338 , n32335 , n32336 );
xor ( n32339 , n31602 , n32050 );
and ( n32340 , n30039 , n32148 );
and ( n32341 , n32339 , n32340 );
xor ( n32342 , n32339 , n32340 );
xor ( n32343 , n31606 , n32048 );
and ( n32344 , n30044 , n32148 );
and ( n32345 , n32343 , n32344 );
xor ( n32346 , n32343 , n32344 );
xor ( n32347 , n31610 , n32046 );
and ( n32348 , n30049 , n32148 );
and ( n32349 , n32347 , n32348 );
xor ( n32350 , n32347 , n32348 );
xor ( n32351 , n31614 , n32044 );
and ( n32352 , n30054 , n32148 );
and ( n32353 , n32351 , n32352 );
xor ( n32354 , n32351 , n32352 );
xor ( n32355 , n31618 , n32042 );
and ( n32356 , n30059 , n32148 );
and ( n32357 , n32355 , n32356 );
xor ( n32358 , n32355 , n32356 );
xor ( n32359 , n31622 , n32040 );
and ( n32360 , n30064 , n32148 );
and ( n32361 , n32359 , n32360 );
xor ( n32362 , n32359 , n32360 );
xor ( n32363 , n31626 , n32038 );
and ( n32364 , n30069 , n32148 );
and ( n32365 , n32363 , n32364 );
xor ( n32366 , n32363 , n32364 );
xor ( n32367 , n31630 , n32036 );
and ( n32368 , n30074 , n32148 );
and ( n32369 , n32367 , n32368 );
xor ( n32370 , n32367 , n32368 );
xor ( n32371 , n31634 , n32034 );
and ( n32372 , n30079 , n32148 );
and ( n32373 , n32371 , n32372 );
xor ( n32374 , n32371 , n32372 );
xor ( n32375 , n31638 , n32032 );
and ( n32376 , n30084 , n32148 );
and ( n32377 , n32375 , n32376 );
xor ( n32378 , n32375 , n32376 );
xor ( n32379 , n31642 , n32030 );
and ( n32380 , n30089 , n32148 );
and ( n32381 , n32379 , n32380 );
xor ( n32382 , n32379 , n32380 );
xor ( n32383 , n31646 , n32028 );
and ( n32384 , n30094 , n32148 );
and ( n32385 , n32383 , n32384 );
xor ( n32386 , n32383 , n32384 );
xor ( n32387 , n31650 , n32026 );
and ( n32388 , n30099 , n32148 );
and ( n32389 , n32387 , n32388 );
xor ( n32390 , n32387 , n32388 );
xor ( n32391 , n31654 , n32024 );
and ( n32392 , n30104 , n32148 );
and ( n32393 , n32391 , n32392 );
xor ( n32394 , n32391 , n32392 );
xor ( n32395 , n31658 , n32022 );
and ( n32396 , n30109 , n32148 );
and ( n32397 , n32395 , n32396 );
xor ( n32398 , n32395 , n32396 );
xor ( n32399 , n31662 , n32020 );
and ( n32400 , n30114 , n32148 );
and ( n32401 , n32399 , n32400 );
xor ( n32402 , n32399 , n32400 );
xor ( n32403 , n31666 , n32018 );
and ( n32404 , n30119 , n32148 );
and ( n32405 , n32403 , n32404 );
xor ( n32406 , n32403 , n32404 );
xor ( n32407 , n31670 , n32016 );
and ( n32408 , n30124 , n32148 );
and ( n32409 , n32407 , n32408 );
xor ( n32410 , n32407 , n32408 );
xor ( n32411 , n31674 , n32014 );
and ( n32412 , n30129 , n32148 );
and ( n32413 , n32411 , n32412 );
xor ( n32414 , n32411 , n32412 );
xor ( n32415 , n31678 , n32012 );
and ( n32416 , n30134 , n32148 );
and ( n32417 , n32415 , n32416 );
xor ( n32418 , n32415 , n32416 );
xor ( n32419 , n31682 , n32010 );
and ( n32420 , n30139 , n32148 );
and ( n32421 , n32419 , n32420 );
xor ( n32422 , n32419 , n32420 );
xor ( n32423 , n31686 , n32008 );
and ( n32424 , n30144 , n32148 );
and ( n32425 , n32423 , n32424 );
xor ( n32426 , n32423 , n32424 );
xor ( n32427 , n31690 , n32006 );
and ( n32428 , n30149 , n32148 );
and ( n32429 , n32427 , n32428 );
xor ( n32430 , n32427 , n32428 );
xor ( n32431 , n31694 , n32004 );
and ( n32432 , n30154 , n32148 );
and ( n32433 , n32431 , n32432 );
xor ( n32434 , n32431 , n32432 );
xor ( n32435 , n31698 , n32002 );
and ( n32436 , n30159 , n32148 );
and ( n32437 , n32435 , n32436 );
xor ( n32438 , n32435 , n32436 );
xor ( n32439 , n31702 , n32000 );
and ( n32440 , n30164 , n32148 );
and ( n32441 , n32439 , n32440 );
xor ( n32442 , n32439 , n32440 );
xor ( n32443 , n31706 , n31998 );
and ( n32444 , n30169 , n32148 );
and ( n32445 , n32443 , n32444 );
xor ( n32446 , n32443 , n32444 );
xor ( n32447 , n31710 , n31996 );
and ( n32448 , n30174 , n32148 );
and ( n32449 , n32447 , n32448 );
xor ( n32450 , n32447 , n32448 );
xor ( n32451 , n31714 , n31994 );
and ( n32452 , n30179 , n32148 );
and ( n32453 , n32451 , n32452 );
xor ( n32454 , n32451 , n32452 );
xor ( n32455 , n31718 , n31992 );
and ( n32456 , n30184 , n32148 );
and ( n32457 , n32455 , n32456 );
xor ( n32458 , n32455 , n32456 );
xor ( n32459 , n31722 , n31990 );
and ( n32460 , n30189 , n32148 );
and ( n32461 , n32459 , n32460 );
xor ( n32462 , n32459 , n32460 );
xor ( n32463 , n31726 , n31988 );
and ( n32464 , n30194 , n32148 );
and ( n32465 , n32463 , n32464 );
xor ( n32466 , n32463 , n32464 );
xor ( n32467 , n31730 , n31986 );
and ( n32468 , n30199 , n32148 );
and ( n32469 , n32467 , n32468 );
xor ( n32470 , n32467 , n32468 );
xor ( n32471 , n31734 , n31984 );
and ( n32472 , n30204 , n32148 );
and ( n32473 , n32471 , n32472 );
xor ( n32474 , n32471 , n32472 );
xor ( n32475 , n31738 , n31982 );
and ( n32476 , n30209 , n32148 );
and ( n32477 , n32475 , n32476 );
xor ( n32478 , n32475 , n32476 );
xor ( n32479 , n31742 , n31980 );
and ( n32480 , n30214 , n32148 );
and ( n32481 , n32479 , n32480 );
xor ( n32482 , n32479 , n32480 );
xor ( n32483 , n31746 , n31978 );
and ( n32484 , n30219 , n32148 );
and ( n32485 , n32483 , n32484 );
xor ( n32486 , n32483 , n32484 );
xor ( n32487 , n31750 , n31976 );
and ( n32488 , n30224 , n32148 );
and ( n32489 , n32487 , n32488 );
xor ( n32490 , n32487 , n32488 );
xor ( n32491 , n31754 , n31974 );
and ( n32492 , n30229 , n32148 );
and ( n32493 , n32491 , n32492 );
xor ( n32494 , n32491 , n32492 );
xor ( n32495 , n31758 , n31972 );
and ( n32496 , n30234 , n32148 );
and ( n32497 , n32495 , n32496 );
xor ( n32498 , n32495 , n32496 );
xor ( n32499 , n31762 , n31970 );
and ( n32500 , n30239 , n32148 );
and ( n32501 , n32499 , n32500 );
xor ( n32502 , n32499 , n32500 );
xor ( n32503 , n31766 , n31968 );
and ( n32504 , n30244 , n32148 );
and ( n32505 , n32503 , n32504 );
xor ( n32506 , n32503 , n32504 );
xor ( n32507 , n31770 , n31966 );
and ( n32508 , n30249 , n32148 );
and ( n32509 , n32507 , n32508 );
xor ( n32510 , n32507 , n32508 );
xor ( n32511 , n31774 , n31964 );
and ( n32512 , n30254 , n32148 );
and ( n32513 , n32511 , n32512 );
xor ( n32514 , n32511 , n32512 );
xor ( n32515 , n31778 , n31962 );
and ( n32516 , n30259 , n32148 );
and ( n32517 , n32515 , n32516 );
xor ( n32518 , n32515 , n32516 );
xor ( n32519 , n31782 , n31960 );
and ( n32520 , n30264 , n32148 );
and ( n32521 , n32519 , n32520 );
xor ( n32522 , n32519 , n32520 );
xor ( n32523 , n31786 , n31958 );
and ( n32524 , n30269 , n32148 );
and ( n32525 , n32523 , n32524 );
xor ( n32526 , n32523 , n32524 );
xor ( n32527 , n31790 , n31956 );
and ( n32528 , n30274 , n32148 );
and ( n32529 , n32527 , n32528 );
xor ( n32530 , n32527 , n32528 );
xor ( n32531 , n31794 , n31954 );
and ( n32532 , n30279 , n32148 );
and ( n32533 , n32531 , n32532 );
xor ( n32534 , n32531 , n32532 );
xor ( n32535 , n31798 , n31952 );
and ( n32536 , n30284 , n32148 );
and ( n32537 , n32535 , n32536 );
xor ( n32538 , n32535 , n32536 );
xor ( n32539 , n31802 , n31950 );
and ( n32540 , n30289 , n32148 );
and ( n32541 , n32539 , n32540 );
xor ( n32542 , n32539 , n32540 );
xor ( n32543 , n31806 , n31948 );
and ( n32544 , n30294 , n32148 );
and ( n32545 , n32543 , n32544 );
xor ( n32546 , n32543 , n32544 );
xor ( n32547 , n31810 , n31946 );
and ( n32548 , n30299 , n32148 );
and ( n32549 , n32547 , n32548 );
xor ( n32550 , n32547 , n32548 );
xor ( n32551 , n31814 , n31944 );
and ( n32552 , n30304 , n32148 );
and ( n32553 , n32551 , n32552 );
xor ( n32554 , n32551 , n32552 );
xor ( n32555 , n31818 , n31942 );
and ( n32556 , n30309 , n32148 );
and ( n32557 , n32555 , n32556 );
xor ( n32558 , n32555 , n32556 );
xor ( n32559 , n31822 , n31940 );
and ( n32560 , n30314 , n32148 );
and ( n32561 , n32559 , n32560 );
xor ( n32562 , n32559 , n32560 );
xor ( n32563 , n31826 , n31938 );
and ( n32564 , n30319 , n32148 );
and ( n32565 , n32563 , n32564 );
xor ( n32566 , n32563 , n32564 );
xor ( n32567 , n31830 , n31936 );
and ( n32568 , n30324 , n32148 );
and ( n32569 , n32567 , n32568 );
xor ( n32570 , n32567 , n32568 );
xor ( n32571 , n31834 , n31934 );
and ( n32572 , n30329 , n32148 );
and ( n32573 , n32571 , n32572 );
xor ( n32574 , n32571 , n32572 );
xor ( n32575 , n31838 , n31932 );
and ( n32576 , n30334 , n32148 );
and ( n32577 , n32575 , n32576 );
xor ( n32578 , n32575 , n32576 );
xor ( n32579 , n31842 , n31930 );
and ( n32580 , n30339 , n32148 );
and ( n32581 , n32579 , n32580 );
xor ( n32582 , n32579 , n32580 );
xor ( n32583 , n31846 , n31928 );
and ( n32584 , n30344 , n32148 );
and ( n32585 , n32583 , n32584 );
xor ( n32586 , n32583 , n32584 );
xor ( n32587 , n31850 , n31926 );
and ( n32588 , n30349 , n32148 );
and ( n32589 , n32587 , n32588 );
xor ( n32590 , n32587 , n32588 );
xor ( n32591 , n31854 , n31924 );
and ( n32592 , n30354 , n32148 );
and ( n32593 , n32591 , n32592 );
xor ( n32594 , n32591 , n32592 );
xor ( n32595 , n31858 , n31922 );
and ( n32596 , n30359 , n32148 );
and ( n32597 , n32595 , n32596 );
xor ( n32598 , n32595 , n32596 );
xor ( n32599 , n31862 , n31920 );
and ( n32600 , n30364 , n32148 );
and ( n32601 , n32599 , n32600 );
xor ( n32602 , n32599 , n32600 );
xor ( n32603 , n31866 , n31918 );
and ( n32604 , n30369 , n32148 );
and ( n32605 , n32603 , n32604 );
xor ( n32606 , n32603 , n32604 );
xor ( n32607 , n31870 , n31916 );
and ( n32608 , n30374 , n32148 );
and ( n32609 , n32607 , n32608 );
xor ( n32610 , n32607 , n32608 );
xor ( n32611 , n31874 , n31914 );
and ( n32612 , n30379 , n32148 );
and ( n32613 , n32611 , n32612 );
xor ( n32614 , n32611 , n32612 );
xor ( n32615 , n31878 , n31912 );
and ( n32616 , n30384 , n32148 );
and ( n32617 , n32615 , n32616 );
xor ( n32618 , n32615 , n32616 );
xor ( n32619 , n31882 , n31910 );
and ( n32620 , n30389 , n32148 );
and ( n32621 , n32619 , n32620 );
xor ( n32622 , n32619 , n32620 );
xor ( n32623 , n31886 , n31908 );
and ( n32624 , n30394 , n32148 );
and ( n32625 , n32623 , n32624 );
xor ( n32626 , n32623 , n32624 );
xor ( n32627 , n31890 , n31906 );
and ( n32628 , n30399 , n32148 );
and ( n32629 , n32627 , n32628 );
xor ( n32630 , n32627 , n32628 );
xor ( n32631 , n31894 , n31904 );
and ( n32632 , n30404 , n32148 );
and ( n32633 , n32631 , n32632 );
xor ( n32634 , n32631 , n32632 );
xor ( n32635 , n31898 , n31902 );
and ( n32636 , n30409 , n32148 );
and ( n32637 , n32635 , n32636 );
buf ( n32638 , n32637 );
and ( n32639 , n32634 , n32638 );
or ( n32640 , n32633 , n32639 );
and ( n32641 , n32630 , n32640 );
or ( n32642 , n32629 , n32641 );
and ( n32643 , n32626 , n32642 );
or ( n32644 , n32625 , n32643 );
and ( n32645 , n32622 , n32644 );
or ( n32646 , n32621 , n32645 );
and ( n32647 , n32618 , n32646 );
or ( n32648 , n32617 , n32647 );
and ( n32649 , n32614 , n32648 );
or ( n32650 , n32613 , n32649 );
and ( n32651 , n32610 , n32650 );
or ( n32652 , n32609 , n32651 );
and ( n32653 , n32606 , n32652 );
or ( n32654 , n32605 , n32653 );
and ( n32655 , n32602 , n32654 );
or ( n32656 , n32601 , n32655 );
and ( n32657 , n32598 , n32656 );
or ( n32658 , n32597 , n32657 );
and ( n32659 , n32594 , n32658 );
or ( n32660 , n32593 , n32659 );
and ( n32661 , n32590 , n32660 );
or ( n32662 , n32589 , n32661 );
and ( n32663 , n32586 , n32662 );
or ( n32664 , n32585 , n32663 );
and ( n32665 , n32582 , n32664 );
or ( n32666 , n32581 , n32665 );
and ( n32667 , n32578 , n32666 );
or ( n32668 , n32577 , n32667 );
and ( n32669 , n32574 , n32668 );
or ( n32670 , n32573 , n32669 );
and ( n32671 , n32570 , n32670 );
or ( n32672 , n32569 , n32671 );
and ( n32673 , n32566 , n32672 );
or ( n32674 , n32565 , n32673 );
and ( n32675 , n32562 , n32674 );
or ( n32676 , n32561 , n32675 );
and ( n32677 , n32558 , n32676 );
or ( n32678 , n32557 , n32677 );
and ( n32679 , n32554 , n32678 );
or ( n32680 , n32553 , n32679 );
and ( n32681 , n32550 , n32680 );
or ( n32682 , n32549 , n32681 );
and ( n32683 , n32546 , n32682 );
or ( n32684 , n32545 , n32683 );
and ( n32685 , n32542 , n32684 );
or ( n32686 , n32541 , n32685 );
and ( n32687 , n32538 , n32686 );
or ( n32688 , n32537 , n32687 );
and ( n32689 , n32534 , n32688 );
or ( n32690 , n32533 , n32689 );
and ( n32691 , n32530 , n32690 );
or ( n32692 , n32529 , n32691 );
and ( n32693 , n32526 , n32692 );
or ( n32694 , n32525 , n32693 );
and ( n32695 , n32522 , n32694 );
or ( n32696 , n32521 , n32695 );
and ( n32697 , n32518 , n32696 );
or ( n32698 , n32517 , n32697 );
and ( n32699 , n32514 , n32698 );
or ( n32700 , n32513 , n32699 );
and ( n32701 , n32510 , n32700 );
or ( n32702 , n32509 , n32701 );
and ( n32703 , n32506 , n32702 );
or ( n32704 , n32505 , n32703 );
and ( n32705 , n32502 , n32704 );
or ( n32706 , n32501 , n32705 );
and ( n32707 , n32498 , n32706 );
or ( n32708 , n32497 , n32707 );
and ( n32709 , n32494 , n32708 );
or ( n32710 , n32493 , n32709 );
and ( n32711 , n32490 , n32710 );
or ( n32712 , n32489 , n32711 );
and ( n32713 , n32486 , n32712 );
or ( n32714 , n32485 , n32713 );
and ( n32715 , n32482 , n32714 );
or ( n32716 , n32481 , n32715 );
and ( n32717 , n32478 , n32716 );
or ( n32718 , n32477 , n32717 );
and ( n32719 , n32474 , n32718 );
or ( n32720 , n32473 , n32719 );
and ( n32721 , n32470 , n32720 );
or ( n32722 , n32469 , n32721 );
and ( n32723 , n32466 , n32722 );
or ( n32724 , n32465 , n32723 );
and ( n32725 , n32462 , n32724 );
or ( n32726 , n32461 , n32725 );
and ( n32727 , n32458 , n32726 );
or ( n32728 , n32457 , n32727 );
and ( n32729 , n32454 , n32728 );
or ( n32730 , n32453 , n32729 );
and ( n32731 , n32450 , n32730 );
or ( n32732 , n32449 , n32731 );
and ( n32733 , n32446 , n32732 );
or ( n32734 , n32445 , n32733 );
and ( n32735 , n32442 , n32734 );
or ( n32736 , n32441 , n32735 );
and ( n32737 , n32438 , n32736 );
or ( n32738 , n32437 , n32737 );
and ( n32739 , n32434 , n32738 );
or ( n32740 , n32433 , n32739 );
and ( n32741 , n32430 , n32740 );
or ( n32742 , n32429 , n32741 );
and ( n32743 , n32426 , n32742 );
or ( n32744 , n32425 , n32743 );
and ( n32745 , n32422 , n32744 );
or ( n32746 , n32421 , n32745 );
and ( n32747 , n32418 , n32746 );
or ( n32748 , n32417 , n32747 );
and ( n32749 , n32414 , n32748 );
or ( n32750 , n32413 , n32749 );
and ( n32751 , n32410 , n32750 );
or ( n32752 , n32409 , n32751 );
and ( n32753 , n32406 , n32752 );
or ( n32754 , n32405 , n32753 );
and ( n32755 , n32402 , n32754 );
or ( n32756 , n32401 , n32755 );
and ( n32757 , n32398 , n32756 );
or ( n32758 , n32397 , n32757 );
and ( n32759 , n32394 , n32758 );
or ( n32760 , n32393 , n32759 );
and ( n32761 , n32390 , n32760 );
or ( n32762 , n32389 , n32761 );
and ( n32763 , n32386 , n32762 );
or ( n32764 , n32385 , n32763 );
and ( n32765 , n32382 , n32764 );
or ( n32766 , n32381 , n32765 );
and ( n32767 , n32378 , n32766 );
or ( n32768 , n32377 , n32767 );
and ( n32769 , n32374 , n32768 );
or ( n32770 , n32373 , n32769 );
and ( n32771 , n32370 , n32770 );
or ( n32772 , n32369 , n32771 );
and ( n32773 , n32366 , n32772 );
or ( n32774 , n32365 , n32773 );
and ( n32775 , n32362 , n32774 );
or ( n32776 , n32361 , n32775 );
and ( n32777 , n32358 , n32776 );
or ( n32778 , n32357 , n32777 );
and ( n32779 , n32354 , n32778 );
or ( n32780 , n32353 , n32779 );
and ( n32781 , n32350 , n32780 );
or ( n32782 , n32349 , n32781 );
and ( n32783 , n32346 , n32782 );
or ( n32784 , n32345 , n32783 );
and ( n32785 , n32342 , n32784 );
or ( n32786 , n32341 , n32785 );
and ( n32787 , n32338 , n32786 );
or ( n32788 , n32337 , n32787 );
and ( n32789 , n32334 , n32788 );
or ( n32790 , n32333 , n32789 );
and ( n32791 , n32330 , n32790 );
or ( n32792 , n32329 , n32791 );
and ( n32793 , n32326 , n32792 );
or ( n32794 , n32325 , n32793 );
and ( n32795 , n32322 , n32794 );
or ( n32796 , n32321 , n32795 );
and ( n32797 , n32318 , n32796 );
or ( n32798 , n32317 , n32797 );
and ( n32799 , n32314 , n32798 );
or ( n32800 , n32313 , n32799 );
and ( n32801 , n32310 , n32800 );
or ( n32802 , n32309 , n32801 );
and ( n32803 , n32306 , n32802 );
or ( n32804 , n32305 , n32803 );
and ( n32805 , n32302 , n32804 );
or ( n32806 , n32301 , n32805 );
and ( n32807 , n32298 , n32806 );
or ( n32808 , n32297 , n32807 );
and ( n32809 , n32294 , n32808 );
or ( n32810 , n32293 , n32809 );
and ( n32811 , n32290 , n32810 );
or ( n32812 , n32289 , n32811 );
and ( n32813 , n32286 , n32812 );
or ( n32814 , n32285 , n32813 );
and ( n32815 , n32282 , n32814 );
or ( n32816 , n32281 , n32815 );
and ( n32817 , n32278 , n32816 );
or ( n32818 , n32277 , n32817 );
and ( n32819 , n32274 , n32818 );
or ( n32820 , n32273 , n32819 );
and ( n32821 , n32270 , n32820 );
or ( n32822 , n32269 , n32821 );
and ( n32823 , n32266 , n32822 );
or ( n32824 , n32265 , n32823 );
and ( n32825 , n32262 , n32824 );
or ( n32826 , n32261 , n32825 );
and ( n32827 , n32258 , n32826 );
or ( n32828 , n32257 , n32827 );
and ( n32829 , n32254 , n32828 );
or ( n32830 , n32253 , n32829 );
and ( n32831 , n32250 , n32830 );
or ( n32832 , n32249 , n32831 );
and ( n32833 , n32246 , n32832 );
or ( n32834 , n32245 , n32833 );
and ( n32835 , n32242 , n32834 );
or ( n32836 , n32241 , n32835 );
and ( n32837 , n32238 , n32836 );
or ( n32838 , n32237 , n32837 );
and ( n32839 , n32234 , n32838 );
or ( n32840 , n32233 , n32839 );
and ( n32841 , n32230 , n32840 );
or ( n32842 , n32229 , n32841 );
and ( n32843 , n32226 , n32842 );
or ( n32844 , n32225 , n32843 );
and ( n32845 , n32222 , n32844 );
or ( n32846 , n32221 , n32845 );
and ( n32847 , n32218 , n32846 );
or ( n32848 , n32217 , n32847 );
and ( n32849 , n32214 , n32848 );
or ( n32850 , n32213 , n32849 );
and ( n32851 , n32210 , n32850 );
or ( n32852 , n32209 , n32851 );
and ( n32853 , n32206 , n32852 );
or ( n32854 , n32205 , n32853 );
and ( n32855 , n32202 , n32854 );
or ( n32856 , n32201 , n32855 );
and ( n32857 , n32198 , n32856 );
or ( n32858 , n32197 , n32857 );
and ( n32859 , n32194 , n32858 );
or ( n32860 , n32193 , n32859 );
and ( n32861 , n32190 , n32860 );
or ( n32862 , n32189 , n32861 );
and ( n32863 , n32186 , n32862 );
or ( n32864 , n32185 , n32863 );
and ( n32865 , n32182 , n32864 );
or ( n32866 , n32181 , n32865 );
and ( n32867 , n32178 , n32866 );
or ( n32868 , n32177 , n32867 );
and ( n32869 , n32174 , n32868 );
or ( n32870 , n32173 , n32869 );
and ( n32871 , n32170 , n32870 );
or ( n32872 , n32169 , n32871 );
and ( n32873 , n32166 , n32872 );
or ( n32874 , n32165 , n32873 );
and ( n32875 , n32162 , n32874 );
or ( n32876 , n32161 , n32875 );
and ( n32877 , n32158 , n32876 );
or ( n32878 , n32157 , n32877 );
and ( n32879 , n32154 , n32878 );
or ( n32880 , n32153 , n32879 );
xor ( n32881 , n32150 , n32880 );
buf ( n32882 , n18096 );
and ( n32883 , n29804 , n32882 );
xor ( n32884 , n32881 , n32883 );
xor ( n32885 , n32154 , n32878 );
and ( n32886 , n29809 , n32882 );
and ( n32887 , n32885 , n32886 );
xor ( n32888 , n32885 , n32886 );
xor ( n32889 , n32158 , n32876 );
and ( n32890 , n29814 , n32882 );
and ( n32891 , n32889 , n32890 );
xor ( n32892 , n32889 , n32890 );
xor ( n32893 , n32162 , n32874 );
and ( n32894 , n29819 , n32882 );
and ( n32895 , n32893 , n32894 );
xor ( n32896 , n32893 , n32894 );
xor ( n32897 , n32166 , n32872 );
and ( n32898 , n29824 , n32882 );
and ( n32899 , n32897 , n32898 );
xor ( n32900 , n32897 , n32898 );
xor ( n32901 , n32170 , n32870 );
and ( n32902 , n29829 , n32882 );
and ( n32903 , n32901 , n32902 );
xor ( n32904 , n32901 , n32902 );
xor ( n32905 , n32174 , n32868 );
and ( n32906 , n29834 , n32882 );
and ( n32907 , n32905 , n32906 );
xor ( n32908 , n32905 , n32906 );
xor ( n32909 , n32178 , n32866 );
and ( n32910 , n29839 , n32882 );
and ( n32911 , n32909 , n32910 );
xor ( n32912 , n32909 , n32910 );
xor ( n32913 , n32182 , n32864 );
and ( n32914 , n29844 , n32882 );
and ( n32915 , n32913 , n32914 );
xor ( n32916 , n32913 , n32914 );
xor ( n32917 , n32186 , n32862 );
and ( n32918 , n29849 , n32882 );
and ( n32919 , n32917 , n32918 );
xor ( n32920 , n32917 , n32918 );
xor ( n32921 , n32190 , n32860 );
and ( n32922 , n29854 , n32882 );
and ( n32923 , n32921 , n32922 );
xor ( n32924 , n32921 , n32922 );
xor ( n32925 , n32194 , n32858 );
and ( n32926 , n29859 , n32882 );
and ( n32927 , n32925 , n32926 );
xor ( n32928 , n32925 , n32926 );
xor ( n32929 , n32198 , n32856 );
and ( n32930 , n29864 , n32882 );
and ( n32931 , n32929 , n32930 );
xor ( n32932 , n32929 , n32930 );
xor ( n32933 , n32202 , n32854 );
and ( n32934 , n29869 , n32882 );
and ( n32935 , n32933 , n32934 );
xor ( n32936 , n32933 , n32934 );
xor ( n32937 , n32206 , n32852 );
and ( n32938 , n29874 , n32882 );
and ( n32939 , n32937 , n32938 );
xor ( n32940 , n32937 , n32938 );
xor ( n32941 , n32210 , n32850 );
and ( n32942 , n29879 , n32882 );
and ( n32943 , n32941 , n32942 );
xor ( n32944 , n32941 , n32942 );
xor ( n32945 , n32214 , n32848 );
and ( n32946 , n29884 , n32882 );
and ( n32947 , n32945 , n32946 );
xor ( n32948 , n32945 , n32946 );
xor ( n32949 , n32218 , n32846 );
and ( n32950 , n29889 , n32882 );
and ( n32951 , n32949 , n32950 );
xor ( n32952 , n32949 , n32950 );
xor ( n32953 , n32222 , n32844 );
and ( n32954 , n29894 , n32882 );
and ( n32955 , n32953 , n32954 );
xor ( n32956 , n32953 , n32954 );
xor ( n32957 , n32226 , n32842 );
and ( n32958 , n29899 , n32882 );
and ( n32959 , n32957 , n32958 );
xor ( n32960 , n32957 , n32958 );
xor ( n32961 , n32230 , n32840 );
and ( n32962 , n29904 , n32882 );
and ( n32963 , n32961 , n32962 );
xor ( n32964 , n32961 , n32962 );
xor ( n32965 , n32234 , n32838 );
and ( n32966 , n29909 , n32882 );
and ( n32967 , n32965 , n32966 );
xor ( n32968 , n32965 , n32966 );
xor ( n32969 , n32238 , n32836 );
and ( n32970 , n29914 , n32882 );
and ( n32971 , n32969 , n32970 );
xor ( n32972 , n32969 , n32970 );
xor ( n32973 , n32242 , n32834 );
and ( n32974 , n29919 , n32882 );
and ( n32975 , n32973 , n32974 );
xor ( n32976 , n32973 , n32974 );
xor ( n32977 , n32246 , n32832 );
and ( n32978 , n29924 , n32882 );
and ( n32979 , n32977 , n32978 );
xor ( n32980 , n32977 , n32978 );
xor ( n32981 , n32250 , n32830 );
and ( n32982 , n29929 , n32882 );
and ( n32983 , n32981 , n32982 );
xor ( n32984 , n32981 , n32982 );
xor ( n32985 , n32254 , n32828 );
and ( n32986 , n29934 , n32882 );
and ( n32987 , n32985 , n32986 );
xor ( n32988 , n32985 , n32986 );
xor ( n32989 , n32258 , n32826 );
and ( n32990 , n29939 , n32882 );
and ( n32991 , n32989 , n32990 );
xor ( n32992 , n32989 , n32990 );
xor ( n32993 , n32262 , n32824 );
and ( n32994 , n29944 , n32882 );
and ( n32995 , n32993 , n32994 );
xor ( n32996 , n32993 , n32994 );
xor ( n32997 , n32266 , n32822 );
and ( n32998 , n29949 , n32882 );
and ( n32999 , n32997 , n32998 );
xor ( n33000 , n32997 , n32998 );
xor ( n33001 , n32270 , n32820 );
and ( n33002 , n29954 , n32882 );
and ( n33003 , n33001 , n33002 );
xor ( n33004 , n33001 , n33002 );
xor ( n33005 , n32274 , n32818 );
and ( n33006 , n29959 , n32882 );
and ( n33007 , n33005 , n33006 );
xor ( n33008 , n33005 , n33006 );
xor ( n33009 , n32278 , n32816 );
and ( n33010 , n29964 , n32882 );
and ( n33011 , n33009 , n33010 );
xor ( n33012 , n33009 , n33010 );
xor ( n33013 , n32282 , n32814 );
and ( n33014 , n29969 , n32882 );
and ( n33015 , n33013 , n33014 );
xor ( n33016 , n33013 , n33014 );
xor ( n33017 , n32286 , n32812 );
and ( n33018 , n29974 , n32882 );
and ( n33019 , n33017 , n33018 );
xor ( n33020 , n33017 , n33018 );
xor ( n33021 , n32290 , n32810 );
and ( n33022 , n29979 , n32882 );
and ( n33023 , n33021 , n33022 );
xor ( n33024 , n33021 , n33022 );
xor ( n33025 , n32294 , n32808 );
and ( n33026 , n29984 , n32882 );
and ( n33027 , n33025 , n33026 );
xor ( n33028 , n33025 , n33026 );
xor ( n33029 , n32298 , n32806 );
and ( n33030 , n29989 , n32882 );
and ( n33031 , n33029 , n33030 );
xor ( n33032 , n33029 , n33030 );
xor ( n33033 , n32302 , n32804 );
and ( n33034 , n29994 , n32882 );
and ( n33035 , n33033 , n33034 );
xor ( n33036 , n33033 , n33034 );
xor ( n33037 , n32306 , n32802 );
and ( n33038 , n29999 , n32882 );
and ( n33039 , n33037 , n33038 );
xor ( n33040 , n33037 , n33038 );
xor ( n33041 , n32310 , n32800 );
and ( n33042 , n30004 , n32882 );
and ( n33043 , n33041 , n33042 );
xor ( n33044 , n33041 , n33042 );
xor ( n33045 , n32314 , n32798 );
and ( n33046 , n30009 , n32882 );
and ( n33047 , n33045 , n33046 );
xor ( n33048 , n33045 , n33046 );
xor ( n33049 , n32318 , n32796 );
and ( n33050 , n30014 , n32882 );
and ( n33051 , n33049 , n33050 );
xor ( n33052 , n33049 , n33050 );
xor ( n33053 , n32322 , n32794 );
and ( n33054 , n30019 , n32882 );
and ( n33055 , n33053 , n33054 );
xor ( n33056 , n33053 , n33054 );
xor ( n33057 , n32326 , n32792 );
and ( n33058 , n30024 , n32882 );
and ( n33059 , n33057 , n33058 );
xor ( n33060 , n33057 , n33058 );
xor ( n33061 , n32330 , n32790 );
and ( n33062 , n30029 , n32882 );
and ( n33063 , n33061 , n33062 );
xor ( n33064 , n33061 , n33062 );
xor ( n33065 , n32334 , n32788 );
and ( n33066 , n30034 , n32882 );
and ( n33067 , n33065 , n33066 );
xor ( n33068 , n33065 , n33066 );
xor ( n33069 , n32338 , n32786 );
and ( n33070 , n30039 , n32882 );
and ( n33071 , n33069 , n33070 );
xor ( n33072 , n33069 , n33070 );
xor ( n33073 , n32342 , n32784 );
and ( n33074 , n30044 , n32882 );
and ( n33075 , n33073 , n33074 );
xor ( n33076 , n33073 , n33074 );
xor ( n33077 , n32346 , n32782 );
and ( n33078 , n30049 , n32882 );
and ( n33079 , n33077 , n33078 );
xor ( n33080 , n33077 , n33078 );
xor ( n33081 , n32350 , n32780 );
and ( n33082 , n30054 , n32882 );
and ( n33083 , n33081 , n33082 );
xor ( n33084 , n33081 , n33082 );
xor ( n33085 , n32354 , n32778 );
and ( n33086 , n30059 , n32882 );
and ( n33087 , n33085 , n33086 );
xor ( n33088 , n33085 , n33086 );
xor ( n33089 , n32358 , n32776 );
and ( n33090 , n30064 , n32882 );
and ( n33091 , n33089 , n33090 );
xor ( n33092 , n33089 , n33090 );
xor ( n33093 , n32362 , n32774 );
and ( n33094 , n30069 , n32882 );
and ( n33095 , n33093 , n33094 );
xor ( n33096 , n33093 , n33094 );
xor ( n33097 , n32366 , n32772 );
and ( n33098 , n30074 , n32882 );
and ( n33099 , n33097 , n33098 );
xor ( n33100 , n33097 , n33098 );
xor ( n33101 , n32370 , n32770 );
and ( n33102 , n30079 , n32882 );
and ( n33103 , n33101 , n33102 );
xor ( n33104 , n33101 , n33102 );
xor ( n33105 , n32374 , n32768 );
and ( n33106 , n30084 , n32882 );
and ( n33107 , n33105 , n33106 );
xor ( n33108 , n33105 , n33106 );
xor ( n33109 , n32378 , n32766 );
and ( n33110 , n30089 , n32882 );
and ( n33111 , n33109 , n33110 );
xor ( n33112 , n33109 , n33110 );
xor ( n33113 , n32382 , n32764 );
and ( n33114 , n30094 , n32882 );
and ( n33115 , n33113 , n33114 );
xor ( n33116 , n33113 , n33114 );
xor ( n33117 , n32386 , n32762 );
and ( n33118 , n30099 , n32882 );
and ( n33119 , n33117 , n33118 );
xor ( n33120 , n33117 , n33118 );
xor ( n33121 , n32390 , n32760 );
and ( n33122 , n30104 , n32882 );
and ( n33123 , n33121 , n33122 );
xor ( n33124 , n33121 , n33122 );
xor ( n33125 , n32394 , n32758 );
and ( n33126 , n30109 , n32882 );
and ( n33127 , n33125 , n33126 );
xor ( n33128 , n33125 , n33126 );
xor ( n33129 , n32398 , n32756 );
and ( n33130 , n30114 , n32882 );
and ( n33131 , n33129 , n33130 );
xor ( n33132 , n33129 , n33130 );
xor ( n33133 , n32402 , n32754 );
and ( n33134 , n30119 , n32882 );
and ( n33135 , n33133 , n33134 );
xor ( n33136 , n33133 , n33134 );
xor ( n33137 , n32406 , n32752 );
and ( n33138 , n30124 , n32882 );
and ( n33139 , n33137 , n33138 );
xor ( n33140 , n33137 , n33138 );
xor ( n33141 , n32410 , n32750 );
and ( n33142 , n30129 , n32882 );
and ( n33143 , n33141 , n33142 );
xor ( n33144 , n33141 , n33142 );
xor ( n33145 , n32414 , n32748 );
and ( n33146 , n30134 , n32882 );
and ( n33147 , n33145 , n33146 );
xor ( n33148 , n33145 , n33146 );
xor ( n33149 , n32418 , n32746 );
and ( n33150 , n30139 , n32882 );
and ( n33151 , n33149 , n33150 );
xor ( n33152 , n33149 , n33150 );
xor ( n33153 , n32422 , n32744 );
and ( n33154 , n30144 , n32882 );
and ( n33155 , n33153 , n33154 );
xor ( n33156 , n33153 , n33154 );
xor ( n33157 , n32426 , n32742 );
and ( n33158 , n30149 , n32882 );
and ( n33159 , n33157 , n33158 );
xor ( n33160 , n33157 , n33158 );
xor ( n33161 , n32430 , n32740 );
and ( n33162 , n30154 , n32882 );
and ( n33163 , n33161 , n33162 );
xor ( n33164 , n33161 , n33162 );
xor ( n33165 , n32434 , n32738 );
and ( n33166 , n30159 , n32882 );
and ( n33167 , n33165 , n33166 );
xor ( n33168 , n33165 , n33166 );
xor ( n33169 , n32438 , n32736 );
and ( n33170 , n30164 , n32882 );
and ( n33171 , n33169 , n33170 );
xor ( n33172 , n33169 , n33170 );
xor ( n33173 , n32442 , n32734 );
and ( n33174 , n30169 , n32882 );
and ( n33175 , n33173 , n33174 );
xor ( n33176 , n33173 , n33174 );
xor ( n33177 , n32446 , n32732 );
and ( n33178 , n30174 , n32882 );
and ( n33179 , n33177 , n33178 );
xor ( n33180 , n33177 , n33178 );
xor ( n33181 , n32450 , n32730 );
and ( n33182 , n30179 , n32882 );
and ( n33183 , n33181 , n33182 );
xor ( n33184 , n33181 , n33182 );
xor ( n33185 , n32454 , n32728 );
and ( n33186 , n30184 , n32882 );
and ( n33187 , n33185 , n33186 );
xor ( n33188 , n33185 , n33186 );
xor ( n33189 , n32458 , n32726 );
and ( n33190 , n30189 , n32882 );
and ( n33191 , n33189 , n33190 );
xor ( n33192 , n33189 , n33190 );
xor ( n33193 , n32462 , n32724 );
and ( n33194 , n30194 , n32882 );
and ( n33195 , n33193 , n33194 );
xor ( n33196 , n33193 , n33194 );
xor ( n33197 , n32466 , n32722 );
and ( n33198 , n30199 , n32882 );
and ( n33199 , n33197 , n33198 );
xor ( n33200 , n33197 , n33198 );
xor ( n33201 , n32470 , n32720 );
and ( n33202 , n30204 , n32882 );
and ( n33203 , n33201 , n33202 );
xor ( n33204 , n33201 , n33202 );
xor ( n33205 , n32474 , n32718 );
and ( n33206 , n30209 , n32882 );
and ( n33207 , n33205 , n33206 );
xor ( n33208 , n33205 , n33206 );
xor ( n33209 , n32478 , n32716 );
and ( n33210 , n30214 , n32882 );
and ( n33211 , n33209 , n33210 );
xor ( n33212 , n33209 , n33210 );
xor ( n33213 , n32482 , n32714 );
and ( n33214 , n30219 , n32882 );
and ( n33215 , n33213 , n33214 );
xor ( n33216 , n33213 , n33214 );
xor ( n33217 , n32486 , n32712 );
and ( n33218 , n30224 , n32882 );
and ( n33219 , n33217 , n33218 );
xor ( n33220 , n33217 , n33218 );
xor ( n33221 , n32490 , n32710 );
and ( n33222 , n30229 , n32882 );
and ( n33223 , n33221 , n33222 );
xor ( n33224 , n33221 , n33222 );
xor ( n33225 , n32494 , n32708 );
and ( n33226 , n30234 , n32882 );
and ( n33227 , n33225 , n33226 );
xor ( n33228 , n33225 , n33226 );
xor ( n33229 , n32498 , n32706 );
and ( n33230 , n30239 , n32882 );
and ( n33231 , n33229 , n33230 );
xor ( n33232 , n33229 , n33230 );
xor ( n33233 , n32502 , n32704 );
and ( n33234 , n30244 , n32882 );
and ( n33235 , n33233 , n33234 );
xor ( n33236 , n33233 , n33234 );
xor ( n33237 , n32506 , n32702 );
and ( n33238 , n30249 , n32882 );
and ( n33239 , n33237 , n33238 );
xor ( n33240 , n33237 , n33238 );
xor ( n33241 , n32510 , n32700 );
and ( n33242 , n30254 , n32882 );
and ( n33243 , n33241 , n33242 );
xor ( n33244 , n33241 , n33242 );
xor ( n33245 , n32514 , n32698 );
and ( n33246 , n30259 , n32882 );
and ( n33247 , n33245 , n33246 );
xor ( n33248 , n33245 , n33246 );
xor ( n33249 , n32518 , n32696 );
and ( n33250 , n30264 , n32882 );
and ( n33251 , n33249 , n33250 );
xor ( n33252 , n33249 , n33250 );
xor ( n33253 , n32522 , n32694 );
and ( n33254 , n30269 , n32882 );
and ( n33255 , n33253 , n33254 );
xor ( n33256 , n33253 , n33254 );
xor ( n33257 , n32526 , n32692 );
and ( n33258 , n30274 , n32882 );
and ( n33259 , n33257 , n33258 );
xor ( n33260 , n33257 , n33258 );
xor ( n33261 , n32530 , n32690 );
and ( n33262 , n30279 , n32882 );
and ( n33263 , n33261 , n33262 );
xor ( n33264 , n33261 , n33262 );
xor ( n33265 , n32534 , n32688 );
and ( n33266 , n30284 , n32882 );
and ( n33267 , n33265 , n33266 );
xor ( n33268 , n33265 , n33266 );
xor ( n33269 , n32538 , n32686 );
and ( n33270 , n30289 , n32882 );
and ( n33271 , n33269 , n33270 );
xor ( n33272 , n33269 , n33270 );
xor ( n33273 , n32542 , n32684 );
and ( n33274 , n30294 , n32882 );
and ( n33275 , n33273 , n33274 );
xor ( n33276 , n33273 , n33274 );
xor ( n33277 , n32546 , n32682 );
and ( n33278 , n30299 , n32882 );
and ( n33279 , n33277 , n33278 );
xor ( n33280 , n33277 , n33278 );
xor ( n33281 , n32550 , n32680 );
and ( n33282 , n30304 , n32882 );
and ( n33283 , n33281 , n33282 );
xor ( n33284 , n33281 , n33282 );
xor ( n33285 , n32554 , n32678 );
and ( n33286 , n30309 , n32882 );
and ( n33287 , n33285 , n33286 );
xor ( n33288 , n33285 , n33286 );
xor ( n33289 , n32558 , n32676 );
and ( n33290 , n30314 , n32882 );
and ( n33291 , n33289 , n33290 );
xor ( n33292 , n33289 , n33290 );
xor ( n33293 , n32562 , n32674 );
and ( n33294 , n30319 , n32882 );
and ( n33295 , n33293 , n33294 );
xor ( n33296 , n33293 , n33294 );
xor ( n33297 , n32566 , n32672 );
and ( n33298 , n30324 , n32882 );
and ( n33299 , n33297 , n33298 );
xor ( n33300 , n33297 , n33298 );
xor ( n33301 , n32570 , n32670 );
and ( n33302 , n30329 , n32882 );
and ( n33303 , n33301 , n33302 );
xor ( n33304 , n33301 , n33302 );
xor ( n33305 , n32574 , n32668 );
and ( n33306 , n30334 , n32882 );
and ( n33307 , n33305 , n33306 );
xor ( n33308 , n33305 , n33306 );
xor ( n33309 , n32578 , n32666 );
and ( n33310 , n30339 , n32882 );
and ( n33311 , n33309 , n33310 );
xor ( n33312 , n33309 , n33310 );
xor ( n33313 , n32582 , n32664 );
and ( n33314 , n30344 , n32882 );
and ( n33315 , n33313 , n33314 );
xor ( n33316 , n33313 , n33314 );
xor ( n33317 , n32586 , n32662 );
and ( n33318 , n30349 , n32882 );
and ( n33319 , n33317 , n33318 );
xor ( n33320 , n33317 , n33318 );
xor ( n33321 , n32590 , n32660 );
and ( n33322 , n30354 , n32882 );
and ( n33323 , n33321 , n33322 );
xor ( n33324 , n33321 , n33322 );
xor ( n33325 , n32594 , n32658 );
and ( n33326 , n30359 , n32882 );
and ( n33327 , n33325 , n33326 );
xor ( n33328 , n33325 , n33326 );
xor ( n33329 , n32598 , n32656 );
and ( n33330 , n30364 , n32882 );
and ( n33331 , n33329 , n33330 );
xor ( n33332 , n33329 , n33330 );
xor ( n33333 , n32602 , n32654 );
and ( n33334 , n30369 , n32882 );
and ( n33335 , n33333 , n33334 );
xor ( n33336 , n33333 , n33334 );
xor ( n33337 , n32606 , n32652 );
and ( n33338 , n30374 , n32882 );
and ( n33339 , n33337 , n33338 );
xor ( n33340 , n33337 , n33338 );
xor ( n33341 , n32610 , n32650 );
and ( n33342 , n30379 , n32882 );
and ( n33343 , n33341 , n33342 );
xor ( n33344 , n33341 , n33342 );
xor ( n33345 , n32614 , n32648 );
and ( n33346 , n30384 , n32882 );
and ( n33347 , n33345 , n33346 );
xor ( n33348 , n33345 , n33346 );
xor ( n33349 , n32618 , n32646 );
and ( n33350 , n30389 , n32882 );
and ( n33351 , n33349 , n33350 );
xor ( n33352 , n33349 , n33350 );
xor ( n33353 , n32622 , n32644 );
and ( n33354 , n30394 , n32882 );
and ( n33355 , n33353 , n33354 );
xor ( n33356 , n33353 , n33354 );
xor ( n33357 , n32626 , n32642 );
and ( n33358 , n30399 , n32882 );
and ( n33359 , n33357 , n33358 );
xor ( n33360 , n33357 , n33358 );
xor ( n33361 , n32630 , n32640 );
and ( n33362 , n30404 , n32882 );
and ( n33363 , n33361 , n33362 );
xor ( n33364 , n33361 , n33362 );
xor ( n33365 , n32634 , n32638 );
and ( n33366 , n30409 , n32882 );
and ( n33367 , n33365 , n33366 );
buf ( n33368 , n33367 );
and ( n33369 , n33364 , n33368 );
or ( n33370 , n33363 , n33369 );
and ( n33371 , n33360 , n33370 );
or ( n33372 , n33359 , n33371 );
and ( n33373 , n33356 , n33372 );
or ( n33374 , n33355 , n33373 );
and ( n33375 , n33352 , n33374 );
or ( n33376 , n33351 , n33375 );
and ( n33377 , n33348 , n33376 );
or ( n33378 , n33347 , n33377 );
and ( n33379 , n33344 , n33378 );
or ( n33380 , n33343 , n33379 );
and ( n33381 , n33340 , n33380 );
or ( n33382 , n33339 , n33381 );
and ( n33383 , n33336 , n33382 );
or ( n33384 , n33335 , n33383 );
and ( n33385 , n33332 , n33384 );
or ( n33386 , n33331 , n33385 );
and ( n33387 , n33328 , n33386 );
or ( n33388 , n33327 , n33387 );
and ( n33389 , n33324 , n33388 );
or ( n33390 , n33323 , n33389 );
and ( n33391 , n33320 , n33390 );
or ( n33392 , n33319 , n33391 );
and ( n33393 , n33316 , n33392 );
or ( n33394 , n33315 , n33393 );
and ( n33395 , n33312 , n33394 );
or ( n33396 , n33311 , n33395 );
and ( n33397 , n33308 , n33396 );
or ( n33398 , n33307 , n33397 );
and ( n33399 , n33304 , n33398 );
or ( n33400 , n33303 , n33399 );
and ( n33401 , n33300 , n33400 );
or ( n33402 , n33299 , n33401 );
and ( n33403 , n33296 , n33402 );
or ( n33404 , n33295 , n33403 );
and ( n33405 , n33292 , n33404 );
or ( n33406 , n33291 , n33405 );
and ( n33407 , n33288 , n33406 );
or ( n33408 , n33287 , n33407 );
and ( n33409 , n33284 , n33408 );
or ( n33410 , n33283 , n33409 );
and ( n33411 , n33280 , n33410 );
or ( n33412 , n33279 , n33411 );
and ( n33413 , n33276 , n33412 );
or ( n33414 , n33275 , n33413 );
and ( n33415 , n33272 , n33414 );
or ( n33416 , n33271 , n33415 );
and ( n33417 , n33268 , n33416 );
or ( n33418 , n33267 , n33417 );
and ( n33419 , n33264 , n33418 );
or ( n33420 , n33263 , n33419 );
and ( n33421 , n33260 , n33420 );
or ( n33422 , n33259 , n33421 );
and ( n33423 , n33256 , n33422 );
or ( n33424 , n33255 , n33423 );
and ( n33425 , n33252 , n33424 );
or ( n33426 , n33251 , n33425 );
and ( n33427 , n33248 , n33426 );
or ( n33428 , n33247 , n33427 );
and ( n33429 , n33244 , n33428 );
or ( n33430 , n33243 , n33429 );
and ( n33431 , n33240 , n33430 );
or ( n33432 , n33239 , n33431 );
and ( n33433 , n33236 , n33432 );
or ( n33434 , n33235 , n33433 );
and ( n33435 , n33232 , n33434 );
or ( n33436 , n33231 , n33435 );
and ( n33437 , n33228 , n33436 );
or ( n33438 , n33227 , n33437 );
and ( n33439 , n33224 , n33438 );
or ( n33440 , n33223 , n33439 );
and ( n33441 , n33220 , n33440 );
or ( n33442 , n33219 , n33441 );
and ( n33443 , n33216 , n33442 );
or ( n33444 , n33215 , n33443 );
and ( n33445 , n33212 , n33444 );
or ( n33446 , n33211 , n33445 );
and ( n33447 , n33208 , n33446 );
or ( n33448 , n33207 , n33447 );
and ( n33449 , n33204 , n33448 );
or ( n33450 , n33203 , n33449 );
and ( n33451 , n33200 , n33450 );
or ( n33452 , n33199 , n33451 );
and ( n33453 , n33196 , n33452 );
or ( n33454 , n33195 , n33453 );
and ( n33455 , n33192 , n33454 );
or ( n33456 , n33191 , n33455 );
and ( n33457 , n33188 , n33456 );
or ( n33458 , n33187 , n33457 );
and ( n33459 , n33184 , n33458 );
or ( n33460 , n33183 , n33459 );
and ( n33461 , n33180 , n33460 );
or ( n33462 , n33179 , n33461 );
and ( n33463 , n33176 , n33462 );
or ( n33464 , n33175 , n33463 );
and ( n33465 , n33172 , n33464 );
or ( n33466 , n33171 , n33465 );
and ( n33467 , n33168 , n33466 );
or ( n33468 , n33167 , n33467 );
and ( n33469 , n33164 , n33468 );
or ( n33470 , n33163 , n33469 );
and ( n33471 , n33160 , n33470 );
or ( n33472 , n33159 , n33471 );
and ( n33473 , n33156 , n33472 );
or ( n33474 , n33155 , n33473 );
and ( n33475 , n33152 , n33474 );
or ( n33476 , n33151 , n33475 );
and ( n33477 , n33148 , n33476 );
or ( n33478 , n33147 , n33477 );
and ( n33479 , n33144 , n33478 );
or ( n33480 , n33143 , n33479 );
and ( n33481 , n33140 , n33480 );
or ( n33482 , n33139 , n33481 );
and ( n33483 , n33136 , n33482 );
or ( n33484 , n33135 , n33483 );
and ( n33485 , n33132 , n33484 );
or ( n33486 , n33131 , n33485 );
and ( n33487 , n33128 , n33486 );
or ( n33488 , n33127 , n33487 );
and ( n33489 , n33124 , n33488 );
or ( n33490 , n33123 , n33489 );
and ( n33491 , n33120 , n33490 );
or ( n33492 , n33119 , n33491 );
and ( n33493 , n33116 , n33492 );
or ( n33494 , n33115 , n33493 );
and ( n33495 , n33112 , n33494 );
or ( n33496 , n33111 , n33495 );
and ( n33497 , n33108 , n33496 );
or ( n33498 , n33107 , n33497 );
and ( n33499 , n33104 , n33498 );
or ( n33500 , n33103 , n33499 );
and ( n33501 , n33100 , n33500 );
or ( n33502 , n33099 , n33501 );
and ( n33503 , n33096 , n33502 );
or ( n33504 , n33095 , n33503 );
and ( n33505 , n33092 , n33504 );
or ( n33506 , n33091 , n33505 );
and ( n33507 , n33088 , n33506 );
or ( n33508 , n33087 , n33507 );
and ( n33509 , n33084 , n33508 );
or ( n33510 , n33083 , n33509 );
and ( n33511 , n33080 , n33510 );
or ( n33512 , n33079 , n33511 );
and ( n33513 , n33076 , n33512 );
or ( n33514 , n33075 , n33513 );
and ( n33515 , n33072 , n33514 );
or ( n33516 , n33071 , n33515 );
and ( n33517 , n33068 , n33516 );
or ( n33518 , n33067 , n33517 );
and ( n33519 , n33064 , n33518 );
or ( n33520 , n33063 , n33519 );
and ( n33521 , n33060 , n33520 );
or ( n33522 , n33059 , n33521 );
and ( n33523 , n33056 , n33522 );
or ( n33524 , n33055 , n33523 );
and ( n33525 , n33052 , n33524 );
or ( n33526 , n33051 , n33525 );
and ( n33527 , n33048 , n33526 );
or ( n33528 , n33047 , n33527 );
and ( n33529 , n33044 , n33528 );
or ( n33530 , n33043 , n33529 );
and ( n33531 , n33040 , n33530 );
or ( n33532 , n33039 , n33531 );
and ( n33533 , n33036 , n33532 );
or ( n33534 , n33035 , n33533 );
and ( n33535 , n33032 , n33534 );
or ( n33536 , n33031 , n33535 );
and ( n33537 , n33028 , n33536 );
or ( n33538 , n33027 , n33537 );
and ( n33539 , n33024 , n33538 );
or ( n33540 , n33023 , n33539 );
and ( n33541 , n33020 , n33540 );
or ( n33542 , n33019 , n33541 );
and ( n33543 , n33016 , n33542 );
or ( n33544 , n33015 , n33543 );
and ( n33545 , n33012 , n33544 );
or ( n33546 , n33011 , n33545 );
and ( n33547 , n33008 , n33546 );
or ( n33548 , n33007 , n33547 );
and ( n33549 , n33004 , n33548 );
or ( n33550 , n33003 , n33549 );
and ( n33551 , n33000 , n33550 );
or ( n33552 , n32999 , n33551 );
and ( n33553 , n32996 , n33552 );
or ( n33554 , n32995 , n33553 );
and ( n33555 , n32992 , n33554 );
or ( n33556 , n32991 , n33555 );
and ( n33557 , n32988 , n33556 );
or ( n33558 , n32987 , n33557 );
and ( n33559 , n32984 , n33558 );
or ( n33560 , n32983 , n33559 );
and ( n33561 , n32980 , n33560 );
or ( n33562 , n32979 , n33561 );
and ( n33563 , n32976 , n33562 );
or ( n33564 , n32975 , n33563 );
and ( n33565 , n32972 , n33564 );
or ( n33566 , n32971 , n33565 );
and ( n33567 , n32968 , n33566 );
or ( n33568 , n32967 , n33567 );
and ( n33569 , n32964 , n33568 );
or ( n33570 , n32963 , n33569 );
and ( n33571 , n32960 , n33570 );
or ( n33572 , n32959 , n33571 );
and ( n33573 , n32956 , n33572 );
or ( n33574 , n32955 , n33573 );
and ( n33575 , n32952 , n33574 );
or ( n33576 , n32951 , n33575 );
and ( n33577 , n32948 , n33576 );
or ( n33578 , n32947 , n33577 );
and ( n33579 , n32944 , n33578 );
or ( n33580 , n32943 , n33579 );
and ( n33581 , n32940 , n33580 );
or ( n33582 , n32939 , n33581 );
and ( n33583 , n32936 , n33582 );
or ( n33584 , n32935 , n33583 );
and ( n33585 , n32932 , n33584 );
or ( n33586 , n32931 , n33585 );
and ( n33587 , n32928 , n33586 );
or ( n33588 , n32927 , n33587 );
and ( n33589 , n32924 , n33588 );
or ( n33590 , n32923 , n33589 );
and ( n33591 , n32920 , n33590 );
or ( n33592 , n32919 , n33591 );
and ( n33593 , n32916 , n33592 );
or ( n33594 , n32915 , n33593 );
and ( n33595 , n32912 , n33594 );
or ( n33596 , n32911 , n33595 );
and ( n33597 , n32908 , n33596 );
or ( n33598 , n32907 , n33597 );
and ( n33599 , n32904 , n33598 );
or ( n33600 , n32903 , n33599 );
and ( n33601 , n32900 , n33600 );
or ( n33602 , n32899 , n33601 );
and ( n33603 , n32896 , n33602 );
or ( n33604 , n32895 , n33603 );
and ( n33605 , n32892 , n33604 );
or ( n33606 , n32891 , n33605 );
and ( n33607 , n32888 , n33606 );
or ( n33608 , n32887 , n33607 );
xor ( n33609 , n32884 , n33608 );
buf ( n33610 , n18094 );
and ( n33611 , n29809 , n33610 );
xor ( n33612 , n33609 , n33611 );
xor ( n33613 , n32888 , n33606 );
and ( n33614 , n29814 , n33610 );
and ( n33615 , n33613 , n33614 );
xor ( n33616 , n33613 , n33614 );
xor ( n33617 , n32892 , n33604 );
and ( n33618 , n29819 , n33610 );
and ( n33619 , n33617 , n33618 );
xor ( n33620 , n33617 , n33618 );
xor ( n33621 , n32896 , n33602 );
and ( n33622 , n29824 , n33610 );
and ( n33623 , n33621 , n33622 );
xor ( n33624 , n33621 , n33622 );
xor ( n33625 , n32900 , n33600 );
and ( n33626 , n29829 , n33610 );
and ( n33627 , n33625 , n33626 );
xor ( n33628 , n33625 , n33626 );
xor ( n33629 , n32904 , n33598 );
and ( n33630 , n29834 , n33610 );
and ( n33631 , n33629 , n33630 );
xor ( n33632 , n33629 , n33630 );
xor ( n33633 , n32908 , n33596 );
and ( n33634 , n29839 , n33610 );
and ( n33635 , n33633 , n33634 );
xor ( n33636 , n33633 , n33634 );
xor ( n33637 , n32912 , n33594 );
and ( n33638 , n29844 , n33610 );
and ( n33639 , n33637 , n33638 );
xor ( n33640 , n33637 , n33638 );
xor ( n33641 , n32916 , n33592 );
and ( n33642 , n29849 , n33610 );
and ( n33643 , n33641 , n33642 );
xor ( n33644 , n33641 , n33642 );
xor ( n33645 , n32920 , n33590 );
and ( n33646 , n29854 , n33610 );
and ( n33647 , n33645 , n33646 );
xor ( n33648 , n33645 , n33646 );
xor ( n33649 , n32924 , n33588 );
and ( n33650 , n29859 , n33610 );
and ( n33651 , n33649 , n33650 );
xor ( n33652 , n33649 , n33650 );
xor ( n33653 , n32928 , n33586 );
and ( n33654 , n29864 , n33610 );
and ( n33655 , n33653 , n33654 );
xor ( n33656 , n33653 , n33654 );
xor ( n33657 , n32932 , n33584 );
and ( n33658 , n29869 , n33610 );
and ( n33659 , n33657 , n33658 );
xor ( n33660 , n33657 , n33658 );
xor ( n33661 , n32936 , n33582 );
and ( n33662 , n29874 , n33610 );
and ( n33663 , n33661 , n33662 );
xor ( n33664 , n33661 , n33662 );
xor ( n33665 , n32940 , n33580 );
and ( n33666 , n29879 , n33610 );
and ( n33667 , n33665 , n33666 );
xor ( n33668 , n33665 , n33666 );
xor ( n33669 , n32944 , n33578 );
and ( n33670 , n29884 , n33610 );
and ( n33671 , n33669 , n33670 );
xor ( n33672 , n33669 , n33670 );
xor ( n33673 , n32948 , n33576 );
and ( n33674 , n29889 , n33610 );
and ( n33675 , n33673 , n33674 );
xor ( n33676 , n33673 , n33674 );
xor ( n33677 , n32952 , n33574 );
and ( n33678 , n29894 , n33610 );
and ( n33679 , n33677 , n33678 );
xor ( n33680 , n33677 , n33678 );
xor ( n33681 , n32956 , n33572 );
and ( n33682 , n29899 , n33610 );
and ( n33683 , n33681 , n33682 );
xor ( n33684 , n33681 , n33682 );
xor ( n33685 , n32960 , n33570 );
and ( n33686 , n29904 , n33610 );
and ( n33687 , n33685 , n33686 );
xor ( n33688 , n33685 , n33686 );
xor ( n33689 , n32964 , n33568 );
and ( n33690 , n29909 , n33610 );
and ( n33691 , n33689 , n33690 );
xor ( n33692 , n33689 , n33690 );
xor ( n33693 , n32968 , n33566 );
and ( n33694 , n29914 , n33610 );
and ( n33695 , n33693 , n33694 );
xor ( n33696 , n33693 , n33694 );
xor ( n33697 , n32972 , n33564 );
and ( n33698 , n29919 , n33610 );
and ( n33699 , n33697 , n33698 );
xor ( n33700 , n33697 , n33698 );
xor ( n33701 , n32976 , n33562 );
and ( n33702 , n29924 , n33610 );
and ( n33703 , n33701 , n33702 );
xor ( n33704 , n33701 , n33702 );
xor ( n33705 , n32980 , n33560 );
and ( n33706 , n29929 , n33610 );
and ( n33707 , n33705 , n33706 );
xor ( n33708 , n33705 , n33706 );
xor ( n33709 , n32984 , n33558 );
and ( n33710 , n29934 , n33610 );
and ( n33711 , n33709 , n33710 );
xor ( n33712 , n33709 , n33710 );
xor ( n33713 , n32988 , n33556 );
and ( n33714 , n29939 , n33610 );
and ( n33715 , n33713 , n33714 );
xor ( n33716 , n33713 , n33714 );
xor ( n33717 , n32992 , n33554 );
and ( n33718 , n29944 , n33610 );
and ( n33719 , n33717 , n33718 );
xor ( n33720 , n33717 , n33718 );
xor ( n33721 , n32996 , n33552 );
and ( n33722 , n29949 , n33610 );
and ( n33723 , n33721 , n33722 );
xor ( n33724 , n33721 , n33722 );
xor ( n33725 , n33000 , n33550 );
and ( n33726 , n29954 , n33610 );
and ( n33727 , n33725 , n33726 );
xor ( n33728 , n33725 , n33726 );
xor ( n33729 , n33004 , n33548 );
and ( n33730 , n29959 , n33610 );
and ( n33731 , n33729 , n33730 );
xor ( n33732 , n33729 , n33730 );
xor ( n33733 , n33008 , n33546 );
and ( n33734 , n29964 , n33610 );
and ( n33735 , n33733 , n33734 );
xor ( n33736 , n33733 , n33734 );
xor ( n33737 , n33012 , n33544 );
and ( n33738 , n29969 , n33610 );
and ( n33739 , n33737 , n33738 );
xor ( n33740 , n33737 , n33738 );
xor ( n33741 , n33016 , n33542 );
and ( n33742 , n29974 , n33610 );
and ( n33743 , n33741 , n33742 );
xor ( n33744 , n33741 , n33742 );
xor ( n33745 , n33020 , n33540 );
and ( n33746 , n29979 , n33610 );
and ( n33747 , n33745 , n33746 );
xor ( n33748 , n33745 , n33746 );
xor ( n33749 , n33024 , n33538 );
and ( n33750 , n29984 , n33610 );
and ( n33751 , n33749 , n33750 );
xor ( n33752 , n33749 , n33750 );
xor ( n33753 , n33028 , n33536 );
and ( n33754 , n29989 , n33610 );
and ( n33755 , n33753 , n33754 );
xor ( n33756 , n33753 , n33754 );
xor ( n33757 , n33032 , n33534 );
and ( n33758 , n29994 , n33610 );
and ( n33759 , n33757 , n33758 );
xor ( n33760 , n33757 , n33758 );
xor ( n33761 , n33036 , n33532 );
and ( n33762 , n29999 , n33610 );
and ( n33763 , n33761 , n33762 );
xor ( n33764 , n33761 , n33762 );
xor ( n33765 , n33040 , n33530 );
and ( n33766 , n30004 , n33610 );
and ( n33767 , n33765 , n33766 );
xor ( n33768 , n33765 , n33766 );
xor ( n33769 , n33044 , n33528 );
and ( n33770 , n30009 , n33610 );
and ( n33771 , n33769 , n33770 );
xor ( n33772 , n33769 , n33770 );
xor ( n33773 , n33048 , n33526 );
and ( n33774 , n30014 , n33610 );
and ( n33775 , n33773 , n33774 );
xor ( n33776 , n33773 , n33774 );
xor ( n33777 , n33052 , n33524 );
and ( n33778 , n30019 , n33610 );
and ( n33779 , n33777 , n33778 );
xor ( n33780 , n33777 , n33778 );
xor ( n33781 , n33056 , n33522 );
and ( n33782 , n30024 , n33610 );
and ( n33783 , n33781 , n33782 );
xor ( n33784 , n33781 , n33782 );
xor ( n33785 , n33060 , n33520 );
and ( n33786 , n30029 , n33610 );
and ( n33787 , n33785 , n33786 );
xor ( n33788 , n33785 , n33786 );
xor ( n33789 , n33064 , n33518 );
and ( n33790 , n30034 , n33610 );
and ( n33791 , n33789 , n33790 );
xor ( n33792 , n33789 , n33790 );
xor ( n33793 , n33068 , n33516 );
and ( n33794 , n30039 , n33610 );
and ( n33795 , n33793 , n33794 );
xor ( n33796 , n33793 , n33794 );
xor ( n33797 , n33072 , n33514 );
and ( n33798 , n30044 , n33610 );
and ( n33799 , n33797 , n33798 );
xor ( n33800 , n33797 , n33798 );
xor ( n33801 , n33076 , n33512 );
and ( n33802 , n30049 , n33610 );
and ( n33803 , n33801 , n33802 );
xor ( n33804 , n33801 , n33802 );
xor ( n33805 , n33080 , n33510 );
and ( n33806 , n30054 , n33610 );
and ( n33807 , n33805 , n33806 );
xor ( n33808 , n33805 , n33806 );
xor ( n33809 , n33084 , n33508 );
and ( n33810 , n30059 , n33610 );
and ( n33811 , n33809 , n33810 );
xor ( n33812 , n33809 , n33810 );
xor ( n33813 , n33088 , n33506 );
and ( n33814 , n30064 , n33610 );
and ( n33815 , n33813 , n33814 );
xor ( n33816 , n33813 , n33814 );
xor ( n33817 , n33092 , n33504 );
and ( n33818 , n30069 , n33610 );
and ( n33819 , n33817 , n33818 );
xor ( n33820 , n33817 , n33818 );
xor ( n33821 , n33096 , n33502 );
and ( n33822 , n30074 , n33610 );
and ( n33823 , n33821 , n33822 );
xor ( n33824 , n33821 , n33822 );
xor ( n33825 , n33100 , n33500 );
and ( n33826 , n30079 , n33610 );
and ( n33827 , n33825 , n33826 );
xor ( n33828 , n33825 , n33826 );
xor ( n33829 , n33104 , n33498 );
and ( n33830 , n30084 , n33610 );
and ( n33831 , n33829 , n33830 );
xor ( n33832 , n33829 , n33830 );
xor ( n33833 , n33108 , n33496 );
and ( n33834 , n30089 , n33610 );
and ( n33835 , n33833 , n33834 );
xor ( n33836 , n33833 , n33834 );
xor ( n33837 , n33112 , n33494 );
and ( n33838 , n30094 , n33610 );
and ( n33839 , n33837 , n33838 );
xor ( n33840 , n33837 , n33838 );
xor ( n33841 , n33116 , n33492 );
and ( n33842 , n30099 , n33610 );
and ( n33843 , n33841 , n33842 );
xor ( n33844 , n33841 , n33842 );
xor ( n33845 , n33120 , n33490 );
and ( n33846 , n30104 , n33610 );
and ( n33847 , n33845 , n33846 );
xor ( n33848 , n33845 , n33846 );
xor ( n33849 , n33124 , n33488 );
and ( n33850 , n30109 , n33610 );
and ( n33851 , n33849 , n33850 );
xor ( n33852 , n33849 , n33850 );
xor ( n33853 , n33128 , n33486 );
and ( n33854 , n30114 , n33610 );
and ( n33855 , n33853 , n33854 );
xor ( n33856 , n33853 , n33854 );
xor ( n33857 , n33132 , n33484 );
and ( n33858 , n30119 , n33610 );
and ( n33859 , n33857 , n33858 );
xor ( n33860 , n33857 , n33858 );
xor ( n33861 , n33136 , n33482 );
and ( n33862 , n30124 , n33610 );
and ( n33863 , n33861 , n33862 );
xor ( n33864 , n33861 , n33862 );
xor ( n33865 , n33140 , n33480 );
and ( n33866 , n30129 , n33610 );
and ( n33867 , n33865 , n33866 );
xor ( n33868 , n33865 , n33866 );
xor ( n33869 , n33144 , n33478 );
and ( n33870 , n30134 , n33610 );
and ( n33871 , n33869 , n33870 );
xor ( n33872 , n33869 , n33870 );
xor ( n33873 , n33148 , n33476 );
and ( n33874 , n30139 , n33610 );
and ( n33875 , n33873 , n33874 );
xor ( n33876 , n33873 , n33874 );
xor ( n33877 , n33152 , n33474 );
and ( n33878 , n30144 , n33610 );
and ( n33879 , n33877 , n33878 );
xor ( n33880 , n33877 , n33878 );
xor ( n33881 , n33156 , n33472 );
and ( n33882 , n30149 , n33610 );
and ( n33883 , n33881 , n33882 );
xor ( n33884 , n33881 , n33882 );
xor ( n33885 , n33160 , n33470 );
and ( n33886 , n30154 , n33610 );
and ( n33887 , n33885 , n33886 );
xor ( n33888 , n33885 , n33886 );
xor ( n33889 , n33164 , n33468 );
and ( n33890 , n30159 , n33610 );
and ( n33891 , n33889 , n33890 );
xor ( n33892 , n33889 , n33890 );
xor ( n33893 , n33168 , n33466 );
and ( n33894 , n30164 , n33610 );
and ( n33895 , n33893 , n33894 );
xor ( n33896 , n33893 , n33894 );
xor ( n33897 , n33172 , n33464 );
and ( n33898 , n30169 , n33610 );
and ( n33899 , n33897 , n33898 );
xor ( n33900 , n33897 , n33898 );
xor ( n33901 , n33176 , n33462 );
and ( n33902 , n30174 , n33610 );
and ( n33903 , n33901 , n33902 );
xor ( n33904 , n33901 , n33902 );
xor ( n33905 , n33180 , n33460 );
and ( n33906 , n30179 , n33610 );
and ( n33907 , n33905 , n33906 );
xor ( n33908 , n33905 , n33906 );
xor ( n33909 , n33184 , n33458 );
and ( n33910 , n30184 , n33610 );
and ( n33911 , n33909 , n33910 );
xor ( n33912 , n33909 , n33910 );
xor ( n33913 , n33188 , n33456 );
and ( n33914 , n30189 , n33610 );
and ( n33915 , n33913 , n33914 );
xor ( n33916 , n33913 , n33914 );
xor ( n33917 , n33192 , n33454 );
and ( n33918 , n30194 , n33610 );
and ( n33919 , n33917 , n33918 );
xor ( n33920 , n33917 , n33918 );
xor ( n33921 , n33196 , n33452 );
and ( n33922 , n30199 , n33610 );
and ( n33923 , n33921 , n33922 );
xor ( n33924 , n33921 , n33922 );
xor ( n33925 , n33200 , n33450 );
and ( n33926 , n30204 , n33610 );
and ( n33927 , n33925 , n33926 );
xor ( n33928 , n33925 , n33926 );
xor ( n33929 , n33204 , n33448 );
and ( n33930 , n30209 , n33610 );
and ( n33931 , n33929 , n33930 );
xor ( n33932 , n33929 , n33930 );
xor ( n33933 , n33208 , n33446 );
and ( n33934 , n30214 , n33610 );
and ( n33935 , n33933 , n33934 );
xor ( n33936 , n33933 , n33934 );
xor ( n33937 , n33212 , n33444 );
and ( n33938 , n30219 , n33610 );
and ( n33939 , n33937 , n33938 );
xor ( n33940 , n33937 , n33938 );
xor ( n33941 , n33216 , n33442 );
and ( n33942 , n30224 , n33610 );
and ( n33943 , n33941 , n33942 );
xor ( n33944 , n33941 , n33942 );
xor ( n33945 , n33220 , n33440 );
and ( n33946 , n30229 , n33610 );
and ( n33947 , n33945 , n33946 );
xor ( n33948 , n33945 , n33946 );
xor ( n33949 , n33224 , n33438 );
and ( n33950 , n30234 , n33610 );
and ( n33951 , n33949 , n33950 );
xor ( n33952 , n33949 , n33950 );
xor ( n33953 , n33228 , n33436 );
and ( n33954 , n30239 , n33610 );
and ( n33955 , n33953 , n33954 );
xor ( n33956 , n33953 , n33954 );
xor ( n33957 , n33232 , n33434 );
and ( n33958 , n30244 , n33610 );
and ( n33959 , n33957 , n33958 );
xor ( n33960 , n33957 , n33958 );
xor ( n33961 , n33236 , n33432 );
and ( n33962 , n30249 , n33610 );
and ( n33963 , n33961 , n33962 );
xor ( n33964 , n33961 , n33962 );
xor ( n33965 , n33240 , n33430 );
and ( n33966 , n30254 , n33610 );
and ( n33967 , n33965 , n33966 );
xor ( n33968 , n33965 , n33966 );
xor ( n33969 , n33244 , n33428 );
and ( n33970 , n30259 , n33610 );
and ( n33971 , n33969 , n33970 );
xor ( n33972 , n33969 , n33970 );
xor ( n33973 , n33248 , n33426 );
and ( n33974 , n30264 , n33610 );
and ( n33975 , n33973 , n33974 );
xor ( n33976 , n33973 , n33974 );
xor ( n33977 , n33252 , n33424 );
and ( n33978 , n30269 , n33610 );
and ( n33979 , n33977 , n33978 );
xor ( n33980 , n33977 , n33978 );
xor ( n33981 , n33256 , n33422 );
and ( n33982 , n30274 , n33610 );
and ( n33983 , n33981 , n33982 );
xor ( n33984 , n33981 , n33982 );
xor ( n33985 , n33260 , n33420 );
and ( n33986 , n30279 , n33610 );
and ( n33987 , n33985 , n33986 );
xor ( n33988 , n33985 , n33986 );
xor ( n33989 , n33264 , n33418 );
and ( n33990 , n30284 , n33610 );
and ( n33991 , n33989 , n33990 );
xor ( n33992 , n33989 , n33990 );
xor ( n33993 , n33268 , n33416 );
and ( n33994 , n30289 , n33610 );
and ( n33995 , n33993 , n33994 );
xor ( n33996 , n33993 , n33994 );
xor ( n33997 , n33272 , n33414 );
and ( n33998 , n30294 , n33610 );
and ( n33999 , n33997 , n33998 );
xor ( n34000 , n33997 , n33998 );
xor ( n34001 , n33276 , n33412 );
and ( n34002 , n30299 , n33610 );
and ( n34003 , n34001 , n34002 );
xor ( n34004 , n34001 , n34002 );
xor ( n34005 , n33280 , n33410 );
and ( n34006 , n30304 , n33610 );
and ( n34007 , n34005 , n34006 );
xor ( n34008 , n34005 , n34006 );
xor ( n34009 , n33284 , n33408 );
and ( n34010 , n30309 , n33610 );
and ( n34011 , n34009 , n34010 );
xor ( n34012 , n34009 , n34010 );
xor ( n34013 , n33288 , n33406 );
and ( n34014 , n30314 , n33610 );
and ( n34015 , n34013 , n34014 );
xor ( n34016 , n34013 , n34014 );
xor ( n34017 , n33292 , n33404 );
and ( n34018 , n30319 , n33610 );
and ( n34019 , n34017 , n34018 );
xor ( n34020 , n34017 , n34018 );
xor ( n34021 , n33296 , n33402 );
and ( n34022 , n30324 , n33610 );
and ( n34023 , n34021 , n34022 );
xor ( n34024 , n34021 , n34022 );
xor ( n34025 , n33300 , n33400 );
and ( n34026 , n30329 , n33610 );
and ( n34027 , n34025 , n34026 );
xor ( n34028 , n34025 , n34026 );
xor ( n34029 , n33304 , n33398 );
and ( n34030 , n30334 , n33610 );
and ( n34031 , n34029 , n34030 );
xor ( n34032 , n34029 , n34030 );
xor ( n34033 , n33308 , n33396 );
and ( n34034 , n30339 , n33610 );
and ( n34035 , n34033 , n34034 );
xor ( n34036 , n34033 , n34034 );
xor ( n34037 , n33312 , n33394 );
and ( n34038 , n30344 , n33610 );
and ( n34039 , n34037 , n34038 );
xor ( n34040 , n34037 , n34038 );
xor ( n34041 , n33316 , n33392 );
and ( n34042 , n30349 , n33610 );
and ( n34043 , n34041 , n34042 );
xor ( n34044 , n34041 , n34042 );
xor ( n34045 , n33320 , n33390 );
and ( n34046 , n30354 , n33610 );
and ( n34047 , n34045 , n34046 );
xor ( n34048 , n34045 , n34046 );
xor ( n34049 , n33324 , n33388 );
and ( n34050 , n30359 , n33610 );
and ( n34051 , n34049 , n34050 );
xor ( n34052 , n34049 , n34050 );
xor ( n34053 , n33328 , n33386 );
and ( n34054 , n30364 , n33610 );
and ( n34055 , n34053 , n34054 );
xor ( n34056 , n34053 , n34054 );
xor ( n34057 , n33332 , n33384 );
and ( n34058 , n30369 , n33610 );
and ( n34059 , n34057 , n34058 );
xor ( n34060 , n34057 , n34058 );
xor ( n34061 , n33336 , n33382 );
and ( n34062 , n30374 , n33610 );
and ( n34063 , n34061 , n34062 );
xor ( n34064 , n34061 , n34062 );
xor ( n34065 , n33340 , n33380 );
and ( n34066 , n30379 , n33610 );
and ( n34067 , n34065 , n34066 );
xor ( n34068 , n34065 , n34066 );
xor ( n34069 , n33344 , n33378 );
and ( n34070 , n30384 , n33610 );
and ( n34071 , n34069 , n34070 );
xor ( n34072 , n34069 , n34070 );
xor ( n34073 , n33348 , n33376 );
and ( n34074 , n30389 , n33610 );
and ( n34075 , n34073 , n34074 );
xor ( n34076 , n34073 , n34074 );
xor ( n34077 , n33352 , n33374 );
and ( n34078 , n30394 , n33610 );
and ( n34079 , n34077 , n34078 );
xor ( n34080 , n34077 , n34078 );
xor ( n34081 , n33356 , n33372 );
and ( n34082 , n30399 , n33610 );
and ( n34083 , n34081 , n34082 );
xor ( n34084 , n34081 , n34082 );
xor ( n34085 , n33360 , n33370 );
and ( n34086 , n30404 , n33610 );
and ( n34087 , n34085 , n34086 );
xor ( n34088 , n34085 , n34086 );
xor ( n34089 , n33364 , n33368 );
and ( n34090 , n30409 , n33610 );
and ( n34091 , n34089 , n34090 );
buf ( n34092 , n34091 );
and ( n34093 , n34088 , n34092 );
or ( n34094 , n34087 , n34093 );
and ( n34095 , n34084 , n34094 );
or ( n34096 , n34083 , n34095 );
and ( n34097 , n34080 , n34096 );
or ( n34098 , n34079 , n34097 );
and ( n34099 , n34076 , n34098 );
or ( n34100 , n34075 , n34099 );
and ( n34101 , n34072 , n34100 );
or ( n34102 , n34071 , n34101 );
and ( n34103 , n34068 , n34102 );
or ( n34104 , n34067 , n34103 );
and ( n34105 , n34064 , n34104 );
or ( n34106 , n34063 , n34105 );
and ( n34107 , n34060 , n34106 );
or ( n34108 , n34059 , n34107 );
and ( n34109 , n34056 , n34108 );
or ( n34110 , n34055 , n34109 );
and ( n34111 , n34052 , n34110 );
or ( n34112 , n34051 , n34111 );
and ( n34113 , n34048 , n34112 );
or ( n34114 , n34047 , n34113 );
and ( n34115 , n34044 , n34114 );
or ( n34116 , n34043 , n34115 );
and ( n34117 , n34040 , n34116 );
or ( n34118 , n34039 , n34117 );
and ( n34119 , n34036 , n34118 );
or ( n34120 , n34035 , n34119 );
and ( n34121 , n34032 , n34120 );
or ( n34122 , n34031 , n34121 );
and ( n34123 , n34028 , n34122 );
or ( n34124 , n34027 , n34123 );
and ( n34125 , n34024 , n34124 );
or ( n34126 , n34023 , n34125 );
and ( n34127 , n34020 , n34126 );
or ( n34128 , n34019 , n34127 );
and ( n34129 , n34016 , n34128 );
or ( n34130 , n34015 , n34129 );
and ( n34131 , n34012 , n34130 );
or ( n34132 , n34011 , n34131 );
and ( n34133 , n34008 , n34132 );
or ( n34134 , n34007 , n34133 );
and ( n34135 , n34004 , n34134 );
or ( n34136 , n34003 , n34135 );
and ( n34137 , n34000 , n34136 );
or ( n34138 , n33999 , n34137 );
and ( n34139 , n33996 , n34138 );
or ( n34140 , n33995 , n34139 );
and ( n34141 , n33992 , n34140 );
or ( n34142 , n33991 , n34141 );
and ( n34143 , n33988 , n34142 );
or ( n34144 , n33987 , n34143 );
and ( n34145 , n33984 , n34144 );
or ( n34146 , n33983 , n34145 );
and ( n34147 , n33980 , n34146 );
or ( n34148 , n33979 , n34147 );
and ( n34149 , n33976 , n34148 );
or ( n34150 , n33975 , n34149 );
and ( n34151 , n33972 , n34150 );
or ( n34152 , n33971 , n34151 );
and ( n34153 , n33968 , n34152 );
or ( n34154 , n33967 , n34153 );
and ( n34155 , n33964 , n34154 );
or ( n34156 , n33963 , n34155 );
and ( n34157 , n33960 , n34156 );
or ( n34158 , n33959 , n34157 );
and ( n34159 , n33956 , n34158 );
or ( n34160 , n33955 , n34159 );
and ( n34161 , n33952 , n34160 );
or ( n34162 , n33951 , n34161 );
and ( n34163 , n33948 , n34162 );
or ( n34164 , n33947 , n34163 );
and ( n34165 , n33944 , n34164 );
or ( n34166 , n33943 , n34165 );
and ( n34167 , n33940 , n34166 );
or ( n34168 , n33939 , n34167 );
and ( n34169 , n33936 , n34168 );
or ( n34170 , n33935 , n34169 );
and ( n34171 , n33932 , n34170 );
or ( n34172 , n33931 , n34171 );
and ( n34173 , n33928 , n34172 );
or ( n34174 , n33927 , n34173 );
and ( n34175 , n33924 , n34174 );
or ( n34176 , n33923 , n34175 );
and ( n34177 , n33920 , n34176 );
or ( n34178 , n33919 , n34177 );
and ( n34179 , n33916 , n34178 );
or ( n34180 , n33915 , n34179 );
and ( n34181 , n33912 , n34180 );
or ( n34182 , n33911 , n34181 );
and ( n34183 , n33908 , n34182 );
or ( n34184 , n33907 , n34183 );
and ( n34185 , n33904 , n34184 );
or ( n34186 , n33903 , n34185 );
and ( n34187 , n33900 , n34186 );
or ( n34188 , n33899 , n34187 );
and ( n34189 , n33896 , n34188 );
or ( n34190 , n33895 , n34189 );
and ( n34191 , n33892 , n34190 );
or ( n34192 , n33891 , n34191 );
and ( n34193 , n33888 , n34192 );
or ( n34194 , n33887 , n34193 );
and ( n34195 , n33884 , n34194 );
or ( n34196 , n33883 , n34195 );
and ( n34197 , n33880 , n34196 );
or ( n34198 , n33879 , n34197 );
and ( n34199 , n33876 , n34198 );
or ( n34200 , n33875 , n34199 );
and ( n34201 , n33872 , n34200 );
or ( n34202 , n33871 , n34201 );
and ( n34203 , n33868 , n34202 );
or ( n34204 , n33867 , n34203 );
and ( n34205 , n33864 , n34204 );
or ( n34206 , n33863 , n34205 );
and ( n34207 , n33860 , n34206 );
or ( n34208 , n33859 , n34207 );
and ( n34209 , n33856 , n34208 );
or ( n34210 , n33855 , n34209 );
and ( n34211 , n33852 , n34210 );
or ( n34212 , n33851 , n34211 );
and ( n34213 , n33848 , n34212 );
or ( n34214 , n33847 , n34213 );
and ( n34215 , n33844 , n34214 );
or ( n34216 , n33843 , n34215 );
and ( n34217 , n33840 , n34216 );
or ( n34218 , n33839 , n34217 );
and ( n34219 , n33836 , n34218 );
or ( n34220 , n33835 , n34219 );
and ( n34221 , n33832 , n34220 );
or ( n34222 , n33831 , n34221 );
and ( n34223 , n33828 , n34222 );
or ( n34224 , n33827 , n34223 );
and ( n34225 , n33824 , n34224 );
or ( n34226 , n33823 , n34225 );
and ( n34227 , n33820 , n34226 );
or ( n34228 , n33819 , n34227 );
and ( n34229 , n33816 , n34228 );
or ( n34230 , n33815 , n34229 );
and ( n34231 , n33812 , n34230 );
or ( n34232 , n33811 , n34231 );
and ( n34233 , n33808 , n34232 );
or ( n34234 , n33807 , n34233 );
and ( n34235 , n33804 , n34234 );
or ( n34236 , n33803 , n34235 );
and ( n34237 , n33800 , n34236 );
or ( n34238 , n33799 , n34237 );
and ( n34239 , n33796 , n34238 );
or ( n34240 , n33795 , n34239 );
and ( n34241 , n33792 , n34240 );
or ( n34242 , n33791 , n34241 );
and ( n34243 , n33788 , n34242 );
or ( n34244 , n33787 , n34243 );
and ( n34245 , n33784 , n34244 );
or ( n34246 , n33783 , n34245 );
and ( n34247 , n33780 , n34246 );
or ( n34248 , n33779 , n34247 );
and ( n34249 , n33776 , n34248 );
or ( n34250 , n33775 , n34249 );
and ( n34251 , n33772 , n34250 );
or ( n34252 , n33771 , n34251 );
and ( n34253 , n33768 , n34252 );
or ( n34254 , n33767 , n34253 );
and ( n34255 , n33764 , n34254 );
or ( n34256 , n33763 , n34255 );
and ( n34257 , n33760 , n34256 );
or ( n34258 , n33759 , n34257 );
and ( n34259 , n33756 , n34258 );
or ( n34260 , n33755 , n34259 );
and ( n34261 , n33752 , n34260 );
or ( n34262 , n33751 , n34261 );
and ( n34263 , n33748 , n34262 );
or ( n34264 , n33747 , n34263 );
and ( n34265 , n33744 , n34264 );
or ( n34266 , n33743 , n34265 );
and ( n34267 , n33740 , n34266 );
or ( n34268 , n33739 , n34267 );
and ( n34269 , n33736 , n34268 );
or ( n34270 , n33735 , n34269 );
and ( n34271 , n33732 , n34270 );
or ( n34272 , n33731 , n34271 );
and ( n34273 , n33728 , n34272 );
or ( n34274 , n33727 , n34273 );
and ( n34275 , n33724 , n34274 );
or ( n34276 , n33723 , n34275 );
and ( n34277 , n33720 , n34276 );
or ( n34278 , n33719 , n34277 );
and ( n34279 , n33716 , n34278 );
or ( n34280 , n33715 , n34279 );
and ( n34281 , n33712 , n34280 );
or ( n34282 , n33711 , n34281 );
and ( n34283 , n33708 , n34282 );
or ( n34284 , n33707 , n34283 );
and ( n34285 , n33704 , n34284 );
or ( n34286 , n33703 , n34285 );
and ( n34287 , n33700 , n34286 );
or ( n34288 , n33699 , n34287 );
and ( n34289 , n33696 , n34288 );
or ( n34290 , n33695 , n34289 );
and ( n34291 , n33692 , n34290 );
or ( n34292 , n33691 , n34291 );
and ( n34293 , n33688 , n34292 );
or ( n34294 , n33687 , n34293 );
and ( n34295 , n33684 , n34294 );
or ( n34296 , n33683 , n34295 );
and ( n34297 , n33680 , n34296 );
or ( n34298 , n33679 , n34297 );
and ( n34299 , n33676 , n34298 );
or ( n34300 , n33675 , n34299 );
and ( n34301 , n33672 , n34300 );
or ( n34302 , n33671 , n34301 );
and ( n34303 , n33668 , n34302 );
or ( n34304 , n33667 , n34303 );
and ( n34305 , n33664 , n34304 );
or ( n34306 , n33663 , n34305 );
and ( n34307 , n33660 , n34306 );
or ( n34308 , n33659 , n34307 );
and ( n34309 , n33656 , n34308 );
or ( n34310 , n33655 , n34309 );
and ( n34311 , n33652 , n34310 );
or ( n34312 , n33651 , n34311 );
and ( n34313 , n33648 , n34312 );
or ( n34314 , n33647 , n34313 );
and ( n34315 , n33644 , n34314 );
or ( n34316 , n33643 , n34315 );
and ( n34317 , n33640 , n34316 );
or ( n34318 , n33639 , n34317 );
and ( n34319 , n33636 , n34318 );
or ( n34320 , n33635 , n34319 );
and ( n34321 , n33632 , n34320 );
or ( n34322 , n33631 , n34321 );
and ( n34323 , n33628 , n34322 );
or ( n34324 , n33627 , n34323 );
and ( n34325 , n33624 , n34324 );
or ( n34326 , n33623 , n34325 );
and ( n34327 , n33620 , n34326 );
or ( n34328 , n33619 , n34327 );
and ( n34329 , n33616 , n34328 );
or ( n34330 , n33615 , n34329 );
xor ( n34331 , n33612 , n34330 );
buf ( n34332 , n18092 );
and ( n34333 , n29814 , n34332 );
xor ( n34334 , n34331 , n34333 );
xor ( n34335 , n33616 , n34328 );
and ( n34336 , n29819 , n34332 );
and ( n34337 , n34335 , n34336 );
xor ( n34338 , n34335 , n34336 );
xor ( n34339 , n33620 , n34326 );
and ( n34340 , n29824 , n34332 );
and ( n34341 , n34339 , n34340 );
xor ( n34342 , n34339 , n34340 );
xor ( n34343 , n33624 , n34324 );
and ( n34344 , n29829 , n34332 );
and ( n34345 , n34343 , n34344 );
xor ( n34346 , n34343 , n34344 );
xor ( n34347 , n33628 , n34322 );
and ( n34348 , n29834 , n34332 );
and ( n34349 , n34347 , n34348 );
xor ( n34350 , n34347 , n34348 );
xor ( n34351 , n33632 , n34320 );
and ( n34352 , n29839 , n34332 );
and ( n34353 , n34351 , n34352 );
xor ( n34354 , n34351 , n34352 );
xor ( n34355 , n33636 , n34318 );
and ( n34356 , n29844 , n34332 );
and ( n34357 , n34355 , n34356 );
xor ( n34358 , n34355 , n34356 );
xor ( n34359 , n33640 , n34316 );
and ( n34360 , n29849 , n34332 );
and ( n34361 , n34359 , n34360 );
xor ( n34362 , n34359 , n34360 );
xor ( n34363 , n33644 , n34314 );
and ( n34364 , n29854 , n34332 );
and ( n34365 , n34363 , n34364 );
xor ( n34366 , n34363 , n34364 );
xor ( n34367 , n33648 , n34312 );
and ( n34368 , n29859 , n34332 );
and ( n34369 , n34367 , n34368 );
xor ( n34370 , n34367 , n34368 );
xor ( n34371 , n33652 , n34310 );
and ( n34372 , n29864 , n34332 );
and ( n34373 , n34371 , n34372 );
xor ( n34374 , n34371 , n34372 );
xor ( n34375 , n33656 , n34308 );
and ( n34376 , n29869 , n34332 );
and ( n34377 , n34375 , n34376 );
xor ( n34378 , n34375 , n34376 );
xor ( n34379 , n33660 , n34306 );
and ( n34380 , n29874 , n34332 );
and ( n34381 , n34379 , n34380 );
xor ( n34382 , n34379 , n34380 );
xor ( n34383 , n33664 , n34304 );
and ( n34384 , n29879 , n34332 );
and ( n34385 , n34383 , n34384 );
xor ( n34386 , n34383 , n34384 );
xor ( n34387 , n33668 , n34302 );
and ( n34388 , n29884 , n34332 );
and ( n34389 , n34387 , n34388 );
xor ( n34390 , n34387 , n34388 );
xor ( n34391 , n33672 , n34300 );
and ( n34392 , n29889 , n34332 );
and ( n34393 , n34391 , n34392 );
xor ( n34394 , n34391 , n34392 );
xor ( n34395 , n33676 , n34298 );
and ( n34396 , n29894 , n34332 );
and ( n34397 , n34395 , n34396 );
xor ( n34398 , n34395 , n34396 );
xor ( n34399 , n33680 , n34296 );
and ( n34400 , n29899 , n34332 );
and ( n34401 , n34399 , n34400 );
xor ( n34402 , n34399 , n34400 );
xor ( n34403 , n33684 , n34294 );
and ( n34404 , n29904 , n34332 );
and ( n34405 , n34403 , n34404 );
xor ( n34406 , n34403 , n34404 );
xor ( n34407 , n33688 , n34292 );
and ( n34408 , n29909 , n34332 );
and ( n34409 , n34407 , n34408 );
xor ( n34410 , n34407 , n34408 );
xor ( n34411 , n33692 , n34290 );
and ( n34412 , n29914 , n34332 );
and ( n34413 , n34411 , n34412 );
xor ( n34414 , n34411 , n34412 );
xor ( n34415 , n33696 , n34288 );
and ( n34416 , n29919 , n34332 );
and ( n34417 , n34415 , n34416 );
xor ( n34418 , n34415 , n34416 );
xor ( n34419 , n33700 , n34286 );
and ( n34420 , n29924 , n34332 );
and ( n34421 , n34419 , n34420 );
xor ( n34422 , n34419 , n34420 );
xor ( n34423 , n33704 , n34284 );
and ( n34424 , n29929 , n34332 );
and ( n34425 , n34423 , n34424 );
xor ( n34426 , n34423 , n34424 );
xor ( n34427 , n33708 , n34282 );
and ( n34428 , n29934 , n34332 );
and ( n34429 , n34427 , n34428 );
xor ( n34430 , n34427 , n34428 );
xor ( n34431 , n33712 , n34280 );
and ( n34432 , n29939 , n34332 );
and ( n34433 , n34431 , n34432 );
xor ( n34434 , n34431 , n34432 );
xor ( n34435 , n33716 , n34278 );
and ( n34436 , n29944 , n34332 );
and ( n34437 , n34435 , n34436 );
xor ( n34438 , n34435 , n34436 );
xor ( n34439 , n33720 , n34276 );
and ( n34440 , n29949 , n34332 );
and ( n34441 , n34439 , n34440 );
xor ( n34442 , n34439 , n34440 );
xor ( n34443 , n33724 , n34274 );
and ( n34444 , n29954 , n34332 );
and ( n34445 , n34443 , n34444 );
xor ( n34446 , n34443 , n34444 );
xor ( n34447 , n33728 , n34272 );
and ( n34448 , n29959 , n34332 );
and ( n34449 , n34447 , n34448 );
xor ( n34450 , n34447 , n34448 );
xor ( n34451 , n33732 , n34270 );
and ( n34452 , n29964 , n34332 );
and ( n34453 , n34451 , n34452 );
xor ( n34454 , n34451 , n34452 );
xor ( n34455 , n33736 , n34268 );
and ( n34456 , n29969 , n34332 );
and ( n34457 , n34455 , n34456 );
xor ( n34458 , n34455 , n34456 );
xor ( n34459 , n33740 , n34266 );
and ( n34460 , n29974 , n34332 );
and ( n34461 , n34459 , n34460 );
xor ( n34462 , n34459 , n34460 );
xor ( n34463 , n33744 , n34264 );
and ( n34464 , n29979 , n34332 );
and ( n34465 , n34463 , n34464 );
xor ( n34466 , n34463 , n34464 );
xor ( n34467 , n33748 , n34262 );
and ( n34468 , n29984 , n34332 );
and ( n34469 , n34467 , n34468 );
xor ( n34470 , n34467 , n34468 );
xor ( n34471 , n33752 , n34260 );
and ( n34472 , n29989 , n34332 );
and ( n34473 , n34471 , n34472 );
xor ( n34474 , n34471 , n34472 );
xor ( n34475 , n33756 , n34258 );
and ( n34476 , n29994 , n34332 );
and ( n34477 , n34475 , n34476 );
xor ( n34478 , n34475 , n34476 );
xor ( n34479 , n33760 , n34256 );
and ( n34480 , n29999 , n34332 );
and ( n34481 , n34479 , n34480 );
xor ( n34482 , n34479 , n34480 );
xor ( n34483 , n33764 , n34254 );
and ( n34484 , n30004 , n34332 );
and ( n34485 , n34483 , n34484 );
xor ( n34486 , n34483 , n34484 );
xor ( n34487 , n33768 , n34252 );
and ( n34488 , n30009 , n34332 );
and ( n34489 , n34487 , n34488 );
xor ( n34490 , n34487 , n34488 );
xor ( n34491 , n33772 , n34250 );
and ( n34492 , n30014 , n34332 );
and ( n34493 , n34491 , n34492 );
xor ( n34494 , n34491 , n34492 );
xor ( n34495 , n33776 , n34248 );
and ( n34496 , n30019 , n34332 );
and ( n34497 , n34495 , n34496 );
xor ( n34498 , n34495 , n34496 );
xor ( n34499 , n33780 , n34246 );
and ( n34500 , n30024 , n34332 );
and ( n34501 , n34499 , n34500 );
xor ( n34502 , n34499 , n34500 );
xor ( n34503 , n33784 , n34244 );
and ( n34504 , n30029 , n34332 );
and ( n34505 , n34503 , n34504 );
xor ( n34506 , n34503 , n34504 );
xor ( n34507 , n33788 , n34242 );
and ( n34508 , n30034 , n34332 );
and ( n34509 , n34507 , n34508 );
xor ( n34510 , n34507 , n34508 );
xor ( n34511 , n33792 , n34240 );
and ( n34512 , n30039 , n34332 );
and ( n34513 , n34511 , n34512 );
xor ( n34514 , n34511 , n34512 );
xor ( n34515 , n33796 , n34238 );
and ( n34516 , n30044 , n34332 );
and ( n34517 , n34515 , n34516 );
xor ( n34518 , n34515 , n34516 );
xor ( n34519 , n33800 , n34236 );
and ( n34520 , n30049 , n34332 );
and ( n34521 , n34519 , n34520 );
xor ( n34522 , n34519 , n34520 );
xor ( n34523 , n33804 , n34234 );
and ( n34524 , n30054 , n34332 );
and ( n34525 , n34523 , n34524 );
xor ( n34526 , n34523 , n34524 );
xor ( n34527 , n33808 , n34232 );
and ( n34528 , n30059 , n34332 );
and ( n34529 , n34527 , n34528 );
xor ( n34530 , n34527 , n34528 );
xor ( n34531 , n33812 , n34230 );
and ( n34532 , n30064 , n34332 );
and ( n34533 , n34531 , n34532 );
xor ( n34534 , n34531 , n34532 );
xor ( n34535 , n33816 , n34228 );
and ( n34536 , n30069 , n34332 );
and ( n34537 , n34535 , n34536 );
xor ( n34538 , n34535 , n34536 );
xor ( n34539 , n33820 , n34226 );
and ( n34540 , n30074 , n34332 );
and ( n34541 , n34539 , n34540 );
xor ( n34542 , n34539 , n34540 );
xor ( n34543 , n33824 , n34224 );
and ( n34544 , n30079 , n34332 );
and ( n34545 , n34543 , n34544 );
xor ( n34546 , n34543 , n34544 );
xor ( n34547 , n33828 , n34222 );
and ( n34548 , n30084 , n34332 );
and ( n34549 , n34547 , n34548 );
xor ( n34550 , n34547 , n34548 );
xor ( n34551 , n33832 , n34220 );
and ( n34552 , n30089 , n34332 );
and ( n34553 , n34551 , n34552 );
xor ( n34554 , n34551 , n34552 );
xor ( n34555 , n33836 , n34218 );
and ( n34556 , n30094 , n34332 );
and ( n34557 , n34555 , n34556 );
xor ( n34558 , n34555 , n34556 );
xor ( n34559 , n33840 , n34216 );
and ( n34560 , n30099 , n34332 );
and ( n34561 , n34559 , n34560 );
xor ( n34562 , n34559 , n34560 );
xor ( n34563 , n33844 , n34214 );
and ( n34564 , n30104 , n34332 );
and ( n34565 , n34563 , n34564 );
xor ( n34566 , n34563 , n34564 );
xor ( n34567 , n33848 , n34212 );
and ( n34568 , n30109 , n34332 );
and ( n34569 , n34567 , n34568 );
xor ( n34570 , n34567 , n34568 );
xor ( n34571 , n33852 , n34210 );
and ( n34572 , n30114 , n34332 );
and ( n34573 , n34571 , n34572 );
xor ( n34574 , n34571 , n34572 );
xor ( n34575 , n33856 , n34208 );
and ( n34576 , n30119 , n34332 );
and ( n34577 , n34575 , n34576 );
xor ( n34578 , n34575 , n34576 );
xor ( n34579 , n33860 , n34206 );
and ( n34580 , n30124 , n34332 );
and ( n34581 , n34579 , n34580 );
xor ( n34582 , n34579 , n34580 );
xor ( n34583 , n33864 , n34204 );
and ( n34584 , n30129 , n34332 );
and ( n34585 , n34583 , n34584 );
xor ( n34586 , n34583 , n34584 );
xor ( n34587 , n33868 , n34202 );
and ( n34588 , n30134 , n34332 );
and ( n34589 , n34587 , n34588 );
xor ( n34590 , n34587 , n34588 );
xor ( n34591 , n33872 , n34200 );
and ( n34592 , n30139 , n34332 );
and ( n34593 , n34591 , n34592 );
xor ( n34594 , n34591 , n34592 );
xor ( n34595 , n33876 , n34198 );
and ( n34596 , n30144 , n34332 );
and ( n34597 , n34595 , n34596 );
xor ( n34598 , n34595 , n34596 );
xor ( n34599 , n33880 , n34196 );
and ( n34600 , n30149 , n34332 );
and ( n34601 , n34599 , n34600 );
xor ( n34602 , n34599 , n34600 );
xor ( n34603 , n33884 , n34194 );
and ( n34604 , n30154 , n34332 );
and ( n34605 , n34603 , n34604 );
xor ( n34606 , n34603 , n34604 );
xor ( n34607 , n33888 , n34192 );
and ( n34608 , n30159 , n34332 );
and ( n34609 , n34607 , n34608 );
xor ( n34610 , n34607 , n34608 );
xor ( n34611 , n33892 , n34190 );
and ( n34612 , n30164 , n34332 );
and ( n34613 , n34611 , n34612 );
xor ( n34614 , n34611 , n34612 );
xor ( n34615 , n33896 , n34188 );
and ( n34616 , n30169 , n34332 );
and ( n34617 , n34615 , n34616 );
xor ( n34618 , n34615 , n34616 );
xor ( n34619 , n33900 , n34186 );
and ( n34620 , n30174 , n34332 );
and ( n34621 , n34619 , n34620 );
xor ( n34622 , n34619 , n34620 );
xor ( n34623 , n33904 , n34184 );
and ( n34624 , n30179 , n34332 );
and ( n34625 , n34623 , n34624 );
xor ( n34626 , n34623 , n34624 );
xor ( n34627 , n33908 , n34182 );
and ( n34628 , n30184 , n34332 );
and ( n34629 , n34627 , n34628 );
xor ( n34630 , n34627 , n34628 );
xor ( n34631 , n33912 , n34180 );
and ( n34632 , n30189 , n34332 );
and ( n34633 , n34631 , n34632 );
xor ( n34634 , n34631 , n34632 );
xor ( n34635 , n33916 , n34178 );
and ( n34636 , n30194 , n34332 );
and ( n34637 , n34635 , n34636 );
xor ( n34638 , n34635 , n34636 );
xor ( n34639 , n33920 , n34176 );
and ( n34640 , n30199 , n34332 );
and ( n34641 , n34639 , n34640 );
xor ( n34642 , n34639 , n34640 );
xor ( n34643 , n33924 , n34174 );
and ( n34644 , n30204 , n34332 );
and ( n34645 , n34643 , n34644 );
xor ( n34646 , n34643 , n34644 );
xor ( n34647 , n33928 , n34172 );
and ( n34648 , n30209 , n34332 );
and ( n34649 , n34647 , n34648 );
xor ( n34650 , n34647 , n34648 );
xor ( n34651 , n33932 , n34170 );
and ( n34652 , n30214 , n34332 );
and ( n34653 , n34651 , n34652 );
xor ( n34654 , n34651 , n34652 );
xor ( n34655 , n33936 , n34168 );
and ( n34656 , n30219 , n34332 );
and ( n34657 , n34655 , n34656 );
xor ( n34658 , n34655 , n34656 );
xor ( n34659 , n33940 , n34166 );
and ( n34660 , n30224 , n34332 );
and ( n34661 , n34659 , n34660 );
xor ( n34662 , n34659 , n34660 );
xor ( n34663 , n33944 , n34164 );
and ( n34664 , n30229 , n34332 );
and ( n34665 , n34663 , n34664 );
xor ( n34666 , n34663 , n34664 );
xor ( n34667 , n33948 , n34162 );
and ( n34668 , n30234 , n34332 );
and ( n34669 , n34667 , n34668 );
xor ( n34670 , n34667 , n34668 );
xor ( n34671 , n33952 , n34160 );
and ( n34672 , n30239 , n34332 );
and ( n34673 , n34671 , n34672 );
xor ( n34674 , n34671 , n34672 );
xor ( n34675 , n33956 , n34158 );
and ( n34676 , n30244 , n34332 );
and ( n34677 , n34675 , n34676 );
xor ( n34678 , n34675 , n34676 );
xor ( n34679 , n33960 , n34156 );
and ( n34680 , n30249 , n34332 );
and ( n34681 , n34679 , n34680 );
xor ( n34682 , n34679 , n34680 );
xor ( n34683 , n33964 , n34154 );
and ( n34684 , n30254 , n34332 );
and ( n34685 , n34683 , n34684 );
xor ( n34686 , n34683 , n34684 );
xor ( n34687 , n33968 , n34152 );
and ( n34688 , n30259 , n34332 );
and ( n34689 , n34687 , n34688 );
xor ( n34690 , n34687 , n34688 );
xor ( n34691 , n33972 , n34150 );
and ( n34692 , n30264 , n34332 );
and ( n34693 , n34691 , n34692 );
xor ( n34694 , n34691 , n34692 );
xor ( n34695 , n33976 , n34148 );
and ( n34696 , n30269 , n34332 );
and ( n34697 , n34695 , n34696 );
xor ( n34698 , n34695 , n34696 );
xor ( n34699 , n33980 , n34146 );
and ( n34700 , n30274 , n34332 );
and ( n34701 , n34699 , n34700 );
xor ( n34702 , n34699 , n34700 );
xor ( n34703 , n33984 , n34144 );
and ( n34704 , n30279 , n34332 );
and ( n34705 , n34703 , n34704 );
xor ( n34706 , n34703 , n34704 );
xor ( n34707 , n33988 , n34142 );
and ( n34708 , n30284 , n34332 );
and ( n34709 , n34707 , n34708 );
xor ( n34710 , n34707 , n34708 );
xor ( n34711 , n33992 , n34140 );
and ( n34712 , n30289 , n34332 );
and ( n34713 , n34711 , n34712 );
xor ( n34714 , n34711 , n34712 );
xor ( n34715 , n33996 , n34138 );
and ( n34716 , n30294 , n34332 );
and ( n34717 , n34715 , n34716 );
xor ( n34718 , n34715 , n34716 );
xor ( n34719 , n34000 , n34136 );
and ( n34720 , n30299 , n34332 );
and ( n34721 , n34719 , n34720 );
xor ( n34722 , n34719 , n34720 );
xor ( n34723 , n34004 , n34134 );
and ( n34724 , n30304 , n34332 );
and ( n34725 , n34723 , n34724 );
xor ( n34726 , n34723 , n34724 );
xor ( n34727 , n34008 , n34132 );
and ( n34728 , n30309 , n34332 );
and ( n34729 , n34727 , n34728 );
xor ( n34730 , n34727 , n34728 );
xor ( n34731 , n34012 , n34130 );
and ( n34732 , n30314 , n34332 );
and ( n34733 , n34731 , n34732 );
xor ( n34734 , n34731 , n34732 );
xor ( n34735 , n34016 , n34128 );
and ( n34736 , n30319 , n34332 );
and ( n34737 , n34735 , n34736 );
xor ( n34738 , n34735 , n34736 );
xor ( n34739 , n34020 , n34126 );
and ( n34740 , n30324 , n34332 );
and ( n34741 , n34739 , n34740 );
xor ( n34742 , n34739 , n34740 );
xor ( n34743 , n34024 , n34124 );
and ( n34744 , n30329 , n34332 );
and ( n34745 , n34743 , n34744 );
xor ( n34746 , n34743 , n34744 );
xor ( n34747 , n34028 , n34122 );
and ( n34748 , n30334 , n34332 );
and ( n34749 , n34747 , n34748 );
xor ( n34750 , n34747 , n34748 );
xor ( n34751 , n34032 , n34120 );
and ( n34752 , n30339 , n34332 );
and ( n34753 , n34751 , n34752 );
xor ( n34754 , n34751 , n34752 );
xor ( n34755 , n34036 , n34118 );
and ( n34756 , n30344 , n34332 );
and ( n34757 , n34755 , n34756 );
xor ( n34758 , n34755 , n34756 );
xor ( n34759 , n34040 , n34116 );
and ( n34760 , n30349 , n34332 );
and ( n34761 , n34759 , n34760 );
xor ( n34762 , n34759 , n34760 );
xor ( n34763 , n34044 , n34114 );
and ( n34764 , n30354 , n34332 );
and ( n34765 , n34763 , n34764 );
xor ( n34766 , n34763 , n34764 );
xor ( n34767 , n34048 , n34112 );
and ( n34768 , n30359 , n34332 );
and ( n34769 , n34767 , n34768 );
xor ( n34770 , n34767 , n34768 );
xor ( n34771 , n34052 , n34110 );
and ( n34772 , n30364 , n34332 );
and ( n34773 , n34771 , n34772 );
xor ( n34774 , n34771 , n34772 );
xor ( n34775 , n34056 , n34108 );
and ( n34776 , n30369 , n34332 );
and ( n34777 , n34775 , n34776 );
xor ( n34778 , n34775 , n34776 );
xor ( n34779 , n34060 , n34106 );
and ( n34780 , n30374 , n34332 );
and ( n34781 , n34779 , n34780 );
xor ( n34782 , n34779 , n34780 );
xor ( n34783 , n34064 , n34104 );
and ( n34784 , n30379 , n34332 );
and ( n34785 , n34783 , n34784 );
xor ( n34786 , n34783 , n34784 );
xor ( n34787 , n34068 , n34102 );
and ( n34788 , n30384 , n34332 );
and ( n34789 , n34787 , n34788 );
xor ( n34790 , n34787 , n34788 );
xor ( n34791 , n34072 , n34100 );
and ( n34792 , n30389 , n34332 );
and ( n34793 , n34791 , n34792 );
xor ( n34794 , n34791 , n34792 );
xor ( n34795 , n34076 , n34098 );
and ( n34796 , n30394 , n34332 );
and ( n34797 , n34795 , n34796 );
xor ( n34798 , n34795 , n34796 );
xor ( n34799 , n34080 , n34096 );
and ( n34800 , n30399 , n34332 );
and ( n34801 , n34799 , n34800 );
xor ( n34802 , n34799 , n34800 );
xor ( n34803 , n34084 , n34094 );
and ( n34804 , n30404 , n34332 );
and ( n34805 , n34803 , n34804 );
xor ( n34806 , n34803 , n34804 );
xor ( n34807 , n34088 , n34092 );
and ( n34808 , n30409 , n34332 );
and ( n34809 , n34807 , n34808 );
buf ( n34810 , n34809 );
and ( n34811 , n34806 , n34810 );
or ( n34812 , n34805 , n34811 );
and ( n34813 , n34802 , n34812 );
or ( n34814 , n34801 , n34813 );
and ( n34815 , n34798 , n34814 );
or ( n34816 , n34797 , n34815 );
and ( n34817 , n34794 , n34816 );
or ( n34818 , n34793 , n34817 );
and ( n34819 , n34790 , n34818 );
or ( n34820 , n34789 , n34819 );
and ( n34821 , n34786 , n34820 );
or ( n34822 , n34785 , n34821 );
and ( n34823 , n34782 , n34822 );
or ( n34824 , n34781 , n34823 );
and ( n34825 , n34778 , n34824 );
or ( n34826 , n34777 , n34825 );
and ( n34827 , n34774 , n34826 );
or ( n34828 , n34773 , n34827 );
and ( n34829 , n34770 , n34828 );
or ( n34830 , n34769 , n34829 );
and ( n34831 , n34766 , n34830 );
or ( n34832 , n34765 , n34831 );
and ( n34833 , n34762 , n34832 );
or ( n34834 , n34761 , n34833 );
and ( n34835 , n34758 , n34834 );
or ( n34836 , n34757 , n34835 );
and ( n34837 , n34754 , n34836 );
or ( n34838 , n34753 , n34837 );
and ( n34839 , n34750 , n34838 );
or ( n34840 , n34749 , n34839 );
and ( n34841 , n34746 , n34840 );
or ( n34842 , n34745 , n34841 );
and ( n34843 , n34742 , n34842 );
or ( n34844 , n34741 , n34843 );
and ( n34845 , n34738 , n34844 );
or ( n34846 , n34737 , n34845 );
and ( n34847 , n34734 , n34846 );
or ( n34848 , n34733 , n34847 );
and ( n34849 , n34730 , n34848 );
or ( n34850 , n34729 , n34849 );
and ( n34851 , n34726 , n34850 );
or ( n34852 , n34725 , n34851 );
and ( n34853 , n34722 , n34852 );
or ( n34854 , n34721 , n34853 );
and ( n34855 , n34718 , n34854 );
or ( n34856 , n34717 , n34855 );
and ( n34857 , n34714 , n34856 );
or ( n34858 , n34713 , n34857 );
and ( n34859 , n34710 , n34858 );
or ( n34860 , n34709 , n34859 );
and ( n34861 , n34706 , n34860 );
or ( n34862 , n34705 , n34861 );
and ( n34863 , n34702 , n34862 );
or ( n34864 , n34701 , n34863 );
and ( n34865 , n34698 , n34864 );
or ( n34866 , n34697 , n34865 );
and ( n34867 , n34694 , n34866 );
or ( n34868 , n34693 , n34867 );
and ( n34869 , n34690 , n34868 );
or ( n34870 , n34689 , n34869 );
and ( n34871 , n34686 , n34870 );
or ( n34872 , n34685 , n34871 );
and ( n34873 , n34682 , n34872 );
or ( n34874 , n34681 , n34873 );
and ( n34875 , n34678 , n34874 );
or ( n34876 , n34677 , n34875 );
and ( n34877 , n34674 , n34876 );
or ( n34878 , n34673 , n34877 );
and ( n34879 , n34670 , n34878 );
or ( n34880 , n34669 , n34879 );
and ( n34881 , n34666 , n34880 );
or ( n34882 , n34665 , n34881 );
and ( n34883 , n34662 , n34882 );
or ( n34884 , n34661 , n34883 );
and ( n34885 , n34658 , n34884 );
or ( n34886 , n34657 , n34885 );
and ( n34887 , n34654 , n34886 );
or ( n34888 , n34653 , n34887 );
and ( n34889 , n34650 , n34888 );
or ( n34890 , n34649 , n34889 );
and ( n34891 , n34646 , n34890 );
or ( n34892 , n34645 , n34891 );
and ( n34893 , n34642 , n34892 );
or ( n34894 , n34641 , n34893 );
and ( n34895 , n34638 , n34894 );
or ( n34896 , n34637 , n34895 );
and ( n34897 , n34634 , n34896 );
or ( n34898 , n34633 , n34897 );
and ( n34899 , n34630 , n34898 );
or ( n34900 , n34629 , n34899 );
and ( n34901 , n34626 , n34900 );
or ( n34902 , n34625 , n34901 );
and ( n34903 , n34622 , n34902 );
or ( n34904 , n34621 , n34903 );
and ( n34905 , n34618 , n34904 );
or ( n34906 , n34617 , n34905 );
and ( n34907 , n34614 , n34906 );
or ( n34908 , n34613 , n34907 );
and ( n34909 , n34610 , n34908 );
or ( n34910 , n34609 , n34909 );
and ( n34911 , n34606 , n34910 );
or ( n34912 , n34605 , n34911 );
and ( n34913 , n34602 , n34912 );
or ( n34914 , n34601 , n34913 );
and ( n34915 , n34598 , n34914 );
or ( n34916 , n34597 , n34915 );
and ( n34917 , n34594 , n34916 );
or ( n34918 , n34593 , n34917 );
and ( n34919 , n34590 , n34918 );
or ( n34920 , n34589 , n34919 );
and ( n34921 , n34586 , n34920 );
or ( n34922 , n34585 , n34921 );
and ( n34923 , n34582 , n34922 );
or ( n34924 , n34581 , n34923 );
and ( n34925 , n34578 , n34924 );
or ( n34926 , n34577 , n34925 );
and ( n34927 , n34574 , n34926 );
or ( n34928 , n34573 , n34927 );
and ( n34929 , n34570 , n34928 );
or ( n34930 , n34569 , n34929 );
and ( n34931 , n34566 , n34930 );
or ( n34932 , n34565 , n34931 );
and ( n34933 , n34562 , n34932 );
or ( n34934 , n34561 , n34933 );
and ( n34935 , n34558 , n34934 );
or ( n34936 , n34557 , n34935 );
and ( n34937 , n34554 , n34936 );
or ( n34938 , n34553 , n34937 );
and ( n34939 , n34550 , n34938 );
or ( n34940 , n34549 , n34939 );
and ( n34941 , n34546 , n34940 );
or ( n34942 , n34545 , n34941 );
and ( n34943 , n34542 , n34942 );
or ( n34944 , n34541 , n34943 );
and ( n34945 , n34538 , n34944 );
or ( n34946 , n34537 , n34945 );
and ( n34947 , n34534 , n34946 );
or ( n34948 , n34533 , n34947 );
and ( n34949 , n34530 , n34948 );
or ( n34950 , n34529 , n34949 );
and ( n34951 , n34526 , n34950 );
or ( n34952 , n34525 , n34951 );
and ( n34953 , n34522 , n34952 );
or ( n34954 , n34521 , n34953 );
and ( n34955 , n34518 , n34954 );
or ( n34956 , n34517 , n34955 );
and ( n34957 , n34514 , n34956 );
or ( n34958 , n34513 , n34957 );
and ( n34959 , n34510 , n34958 );
or ( n34960 , n34509 , n34959 );
and ( n34961 , n34506 , n34960 );
or ( n34962 , n34505 , n34961 );
and ( n34963 , n34502 , n34962 );
or ( n34964 , n34501 , n34963 );
and ( n34965 , n34498 , n34964 );
or ( n34966 , n34497 , n34965 );
and ( n34967 , n34494 , n34966 );
or ( n34968 , n34493 , n34967 );
and ( n34969 , n34490 , n34968 );
or ( n34970 , n34489 , n34969 );
and ( n34971 , n34486 , n34970 );
or ( n34972 , n34485 , n34971 );
and ( n34973 , n34482 , n34972 );
or ( n34974 , n34481 , n34973 );
and ( n34975 , n34478 , n34974 );
or ( n34976 , n34477 , n34975 );
and ( n34977 , n34474 , n34976 );
or ( n34978 , n34473 , n34977 );
and ( n34979 , n34470 , n34978 );
or ( n34980 , n34469 , n34979 );
and ( n34981 , n34466 , n34980 );
or ( n34982 , n34465 , n34981 );
and ( n34983 , n34462 , n34982 );
or ( n34984 , n34461 , n34983 );
and ( n34985 , n34458 , n34984 );
or ( n34986 , n34457 , n34985 );
and ( n34987 , n34454 , n34986 );
or ( n34988 , n34453 , n34987 );
and ( n34989 , n34450 , n34988 );
or ( n34990 , n34449 , n34989 );
and ( n34991 , n34446 , n34990 );
or ( n34992 , n34445 , n34991 );
and ( n34993 , n34442 , n34992 );
or ( n34994 , n34441 , n34993 );
and ( n34995 , n34438 , n34994 );
or ( n34996 , n34437 , n34995 );
and ( n34997 , n34434 , n34996 );
or ( n34998 , n34433 , n34997 );
and ( n34999 , n34430 , n34998 );
or ( n35000 , n34429 , n34999 );
and ( n35001 , n34426 , n35000 );
or ( n35002 , n34425 , n35001 );
and ( n35003 , n34422 , n35002 );
or ( n35004 , n34421 , n35003 );
and ( n35005 , n34418 , n35004 );
or ( n35006 , n34417 , n35005 );
and ( n35007 , n34414 , n35006 );
or ( n35008 , n34413 , n35007 );
and ( n35009 , n34410 , n35008 );
or ( n35010 , n34409 , n35009 );
and ( n35011 , n34406 , n35010 );
or ( n35012 , n34405 , n35011 );
and ( n35013 , n34402 , n35012 );
or ( n35014 , n34401 , n35013 );
and ( n35015 , n34398 , n35014 );
or ( n35016 , n34397 , n35015 );
and ( n35017 , n34394 , n35016 );
or ( n35018 , n34393 , n35017 );
and ( n35019 , n34390 , n35018 );
or ( n35020 , n34389 , n35019 );
and ( n35021 , n34386 , n35020 );
or ( n35022 , n34385 , n35021 );
and ( n35023 , n34382 , n35022 );
or ( n35024 , n34381 , n35023 );
and ( n35025 , n34378 , n35024 );
or ( n35026 , n34377 , n35025 );
and ( n35027 , n34374 , n35026 );
or ( n35028 , n34373 , n35027 );
and ( n35029 , n34370 , n35028 );
or ( n35030 , n34369 , n35029 );
and ( n35031 , n34366 , n35030 );
or ( n35032 , n34365 , n35031 );
and ( n35033 , n34362 , n35032 );
or ( n35034 , n34361 , n35033 );
and ( n35035 , n34358 , n35034 );
or ( n35036 , n34357 , n35035 );
and ( n35037 , n34354 , n35036 );
or ( n35038 , n34353 , n35037 );
and ( n35039 , n34350 , n35038 );
or ( n35040 , n34349 , n35039 );
and ( n35041 , n34346 , n35040 );
or ( n35042 , n34345 , n35041 );
and ( n35043 , n34342 , n35042 );
or ( n35044 , n34341 , n35043 );
and ( n35045 , n34338 , n35044 );
or ( n35046 , n34337 , n35045 );
xor ( n35047 , n34334 , n35046 );
buf ( n35048 , n18090 );
and ( n35049 , n29819 , n35048 );
xor ( n35050 , n35047 , n35049 );
xor ( n35051 , n34338 , n35044 );
and ( n35052 , n29824 , n35048 );
and ( n35053 , n35051 , n35052 );
xor ( n35054 , n35051 , n35052 );
xor ( n35055 , n34342 , n35042 );
and ( n35056 , n29829 , n35048 );
and ( n35057 , n35055 , n35056 );
xor ( n35058 , n35055 , n35056 );
xor ( n35059 , n34346 , n35040 );
and ( n35060 , n29834 , n35048 );
and ( n35061 , n35059 , n35060 );
xor ( n35062 , n35059 , n35060 );
xor ( n35063 , n34350 , n35038 );
and ( n35064 , n29839 , n35048 );
and ( n35065 , n35063 , n35064 );
xor ( n35066 , n35063 , n35064 );
xor ( n35067 , n34354 , n35036 );
and ( n35068 , n29844 , n35048 );
and ( n35069 , n35067 , n35068 );
xor ( n35070 , n35067 , n35068 );
xor ( n35071 , n34358 , n35034 );
and ( n35072 , n29849 , n35048 );
and ( n35073 , n35071 , n35072 );
xor ( n35074 , n35071 , n35072 );
xor ( n35075 , n34362 , n35032 );
and ( n35076 , n29854 , n35048 );
and ( n35077 , n35075 , n35076 );
xor ( n35078 , n35075 , n35076 );
xor ( n35079 , n34366 , n35030 );
and ( n35080 , n29859 , n35048 );
and ( n35081 , n35079 , n35080 );
xor ( n35082 , n35079 , n35080 );
xor ( n35083 , n34370 , n35028 );
and ( n35084 , n29864 , n35048 );
and ( n35085 , n35083 , n35084 );
xor ( n35086 , n35083 , n35084 );
xor ( n35087 , n34374 , n35026 );
and ( n35088 , n29869 , n35048 );
and ( n35089 , n35087 , n35088 );
xor ( n35090 , n35087 , n35088 );
xor ( n35091 , n34378 , n35024 );
and ( n35092 , n29874 , n35048 );
and ( n35093 , n35091 , n35092 );
xor ( n35094 , n35091 , n35092 );
xor ( n35095 , n34382 , n35022 );
and ( n35096 , n29879 , n35048 );
and ( n35097 , n35095 , n35096 );
xor ( n35098 , n35095 , n35096 );
xor ( n35099 , n34386 , n35020 );
and ( n35100 , n29884 , n35048 );
and ( n35101 , n35099 , n35100 );
xor ( n35102 , n35099 , n35100 );
xor ( n35103 , n34390 , n35018 );
and ( n35104 , n29889 , n35048 );
and ( n35105 , n35103 , n35104 );
xor ( n35106 , n35103 , n35104 );
xor ( n35107 , n34394 , n35016 );
and ( n35108 , n29894 , n35048 );
and ( n35109 , n35107 , n35108 );
xor ( n35110 , n35107 , n35108 );
xor ( n35111 , n34398 , n35014 );
and ( n35112 , n29899 , n35048 );
and ( n35113 , n35111 , n35112 );
xor ( n35114 , n35111 , n35112 );
xor ( n35115 , n34402 , n35012 );
and ( n35116 , n29904 , n35048 );
and ( n35117 , n35115 , n35116 );
xor ( n35118 , n35115 , n35116 );
xor ( n35119 , n34406 , n35010 );
and ( n35120 , n29909 , n35048 );
and ( n35121 , n35119 , n35120 );
xor ( n35122 , n35119 , n35120 );
xor ( n35123 , n34410 , n35008 );
and ( n35124 , n29914 , n35048 );
and ( n35125 , n35123 , n35124 );
xor ( n35126 , n35123 , n35124 );
xor ( n35127 , n34414 , n35006 );
and ( n35128 , n29919 , n35048 );
and ( n35129 , n35127 , n35128 );
xor ( n35130 , n35127 , n35128 );
xor ( n35131 , n34418 , n35004 );
and ( n35132 , n29924 , n35048 );
and ( n35133 , n35131 , n35132 );
xor ( n35134 , n35131 , n35132 );
xor ( n35135 , n34422 , n35002 );
and ( n35136 , n29929 , n35048 );
and ( n35137 , n35135 , n35136 );
xor ( n35138 , n35135 , n35136 );
xor ( n35139 , n34426 , n35000 );
and ( n35140 , n29934 , n35048 );
and ( n35141 , n35139 , n35140 );
xor ( n35142 , n35139 , n35140 );
xor ( n35143 , n34430 , n34998 );
and ( n35144 , n29939 , n35048 );
and ( n35145 , n35143 , n35144 );
xor ( n35146 , n35143 , n35144 );
xor ( n35147 , n34434 , n34996 );
and ( n35148 , n29944 , n35048 );
and ( n35149 , n35147 , n35148 );
xor ( n35150 , n35147 , n35148 );
xor ( n35151 , n34438 , n34994 );
and ( n35152 , n29949 , n35048 );
and ( n35153 , n35151 , n35152 );
xor ( n35154 , n35151 , n35152 );
xor ( n35155 , n34442 , n34992 );
and ( n35156 , n29954 , n35048 );
and ( n35157 , n35155 , n35156 );
xor ( n35158 , n35155 , n35156 );
xor ( n35159 , n34446 , n34990 );
and ( n35160 , n29959 , n35048 );
and ( n35161 , n35159 , n35160 );
xor ( n35162 , n35159 , n35160 );
xor ( n35163 , n34450 , n34988 );
and ( n35164 , n29964 , n35048 );
and ( n35165 , n35163 , n35164 );
xor ( n35166 , n35163 , n35164 );
xor ( n35167 , n34454 , n34986 );
and ( n35168 , n29969 , n35048 );
and ( n35169 , n35167 , n35168 );
xor ( n35170 , n35167 , n35168 );
xor ( n35171 , n34458 , n34984 );
and ( n35172 , n29974 , n35048 );
and ( n35173 , n35171 , n35172 );
xor ( n35174 , n35171 , n35172 );
xor ( n35175 , n34462 , n34982 );
and ( n35176 , n29979 , n35048 );
and ( n35177 , n35175 , n35176 );
xor ( n35178 , n35175 , n35176 );
xor ( n35179 , n34466 , n34980 );
and ( n35180 , n29984 , n35048 );
and ( n35181 , n35179 , n35180 );
xor ( n35182 , n35179 , n35180 );
xor ( n35183 , n34470 , n34978 );
and ( n35184 , n29989 , n35048 );
and ( n35185 , n35183 , n35184 );
xor ( n35186 , n35183 , n35184 );
xor ( n35187 , n34474 , n34976 );
and ( n35188 , n29994 , n35048 );
and ( n35189 , n35187 , n35188 );
xor ( n35190 , n35187 , n35188 );
xor ( n35191 , n34478 , n34974 );
and ( n35192 , n29999 , n35048 );
and ( n35193 , n35191 , n35192 );
xor ( n35194 , n35191 , n35192 );
xor ( n35195 , n34482 , n34972 );
and ( n35196 , n30004 , n35048 );
and ( n35197 , n35195 , n35196 );
xor ( n35198 , n35195 , n35196 );
xor ( n35199 , n34486 , n34970 );
and ( n35200 , n30009 , n35048 );
and ( n35201 , n35199 , n35200 );
xor ( n35202 , n35199 , n35200 );
xor ( n35203 , n34490 , n34968 );
and ( n35204 , n30014 , n35048 );
and ( n35205 , n35203 , n35204 );
xor ( n35206 , n35203 , n35204 );
xor ( n35207 , n34494 , n34966 );
and ( n35208 , n30019 , n35048 );
and ( n35209 , n35207 , n35208 );
xor ( n35210 , n35207 , n35208 );
xor ( n35211 , n34498 , n34964 );
and ( n35212 , n30024 , n35048 );
and ( n35213 , n35211 , n35212 );
xor ( n35214 , n35211 , n35212 );
xor ( n35215 , n34502 , n34962 );
and ( n35216 , n30029 , n35048 );
and ( n35217 , n35215 , n35216 );
xor ( n35218 , n35215 , n35216 );
xor ( n35219 , n34506 , n34960 );
and ( n35220 , n30034 , n35048 );
and ( n35221 , n35219 , n35220 );
xor ( n35222 , n35219 , n35220 );
xor ( n35223 , n34510 , n34958 );
and ( n35224 , n30039 , n35048 );
and ( n35225 , n35223 , n35224 );
xor ( n35226 , n35223 , n35224 );
xor ( n35227 , n34514 , n34956 );
and ( n35228 , n30044 , n35048 );
and ( n35229 , n35227 , n35228 );
xor ( n35230 , n35227 , n35228 );
xor ( n35231 , n34518 , n34954 );
and ( n35232 , n30049 , n35048 );
and ( n35233 , n35231 , n35232 );
xor ( n35234 , n35231 , n35232 );
xor ( n35235 , n34522 , n34952 );
and ( n35236 , n30054 , n35048 );
and ( n35237 , n35235 , n35236 );
xor ( n35238 , n35235 , n35236 );
xor ( n35239 , n34526 , n34950 );
and ( n35240 , n30059 , n35048 );
and ( n35241 , n35239 , n35240 );
xor ( n35242 , n35239 , n35240 );
xor ( n35243 , n34530 , n34948 );
and ( n35244 , n30064 , n35048 );
and ( n35245 , n35243 , n35244 );
xor ( n35246 , n35243 , n35244 );
xor ( n35247 , n34534 , n34946 );
and ( n35248 , n30069 , n35048 );
and ( n35249 , n35247 , n35248 );
xor ( n35250 , n35247 , n35248 );
xor ( n35251 , n34538 , n34944 );
and ( n35252 , n30074 , n35048 );
and ( n35253 , n35251 , n35252 );
xor ( n35254 , n35251 , n35252 );
xor ( n35255 , n34542 , n34942 );
and ( n35256 , n30079 , n35048 );
and ( n35257 , n35255 , n35256 );
xor ( n35258 , n35255 , n35256 );
xor ( n35259 , n34546 , n34940 );
and ( n35260 , n30084 , n35048 );
and ( n35261 , n35259 , n35260 );
xor ( n35262 , n35259 , n35260 );
xor ( n35263 , n34550 , n34938 );
and ( n35264 , n30089 , n35048 );
and ( n35265 , n35263 , n35264 );
xor ( n35266 , n35263 , n35264 );
xor ( n35267 , n34554 , n34936 );
and ( n35268 , n30094 , n35048 );
and ( n35269 , n35267 , n35268 );
xor ( n35270 , n35267 , n35268 );
xor ( n35271 , n34558 , n34934 );
and ( n35272 , n30099 , n35048 );
and ( n35273 , n35271 , n35272 );
xor ( n35274 , n35271 , n35272 );
xor ( n35275 , n34562 , n34932 );
and ( n35276 , n30104 , n35048 );
and ( n35277 , n35275 , n35276 );
xor ( n35278 , n35275 , n35276 );
xor ( n35279 , n34566 , n34930 );
and ( n35280 , n30109 , n35048 );
and ( n35281 , n35279 , n35280 );
xor ( n35282 , n35279 , n35280 );
xor ( n35283 , n34570 , n34928 );
and ( n35284 , n30114 , n35048 );
and ( n35285 , n35283 , n35284 );
xor ( n35286 , n35283 , n35284 );
xor ( n35287 , n34574 , n34926 );
and ( n35288 , n30119 , n35048 );
and ( n35289 , n35287 , n35288 );
xor ( n35290 , n35287 , n35288 );
xor ( n35291 , n34578 , n34924 );
and ( n35292 , n30124 , n35048 );
and ( n35293 , n35291 , n35292 );
xor ( n35294 , n35291 , n35292 );
xor ( n35295 , n34582 , n34922 );
and ( n35296 , n30129 , n35048 );
and ( n35297 , n35295 , n35296 );
xor ( n35298 , n35295 , n35296 );
xor ( n35299 , n34586 , n34920 );
and ( n35300 , n30134 , n35048 );
and ( n35301 , n35299 , n35300 );
xor ( n35302 , n35299 , n35300 );
xor ( n35303 , n34590 , n34918 );
and ( n35304 , n30139 , n35048 );
and ( n35305 , n35303 , n35304 );
xor ( n35306 , n35303 , n35304 );
xor ( n35307 , n34594 , n34916 );
and ( n35308 , n30144 , n35048 );
and ( n35309 , n35307 , n35308 );
xor ( n35310 , n35307 , n35308 );
xor ( n35311 , n34598 , n34914 );
and ( n35312 , n30149 , n35048 );
and ( n35313 , n35311 , n35312 );
xor ( n35314 , n35311 , n35312 );
xor ( n35315 , n34602 , n34912 );
and ( n35316 , n30154 , n35048 );
and ( n35317 , n35315 , n35316 );
xor ( n35318 , n35315 , n35316 );
xor ( n35319 , n34606 , n34910 );
and ( n35320 , n30159 , n35048 );
and ( n35321 , n35319 , n35320 );
xor ( n35322 , n35319 , n35320 );
xor ( n35323 , n34610 , n34908 );
and ( n35324 , n30164 , n35048 );
and ( n35325 , n35323 , n35324 );
xor ( n35326 , n35323 , n35324 );
xor ( n35327 , n34614 , n34906 );
and ( n35328 , n30169 , n35048 );
and ( n35329 , n35327 , n35328 );
xor ( n35330 , n35327 , n35328 );
xor ( n35331 , n34618 , n34904 );
and ( n35332 , n30174 , n35048 );
and ( n35333 , n35331 , n35332 );
xor ( n35334 , n35331 , n35332 );
xor ( n35335 , n34622 , n34902 );
and ( n35336 , n30179 , n35048 );
and ( n35337 , n35335 , n35336 );
xor ( n35338 , n35335 , n35336 );
xor ( n35339 , n34626 , n34900 );
and ( n35340 , n30184 , n35048 );
and ( n35341 , n35339 , n35340 );
xor ( n35342 , n35339 , n35340 );
xor ( n35343 , n34630 , n34898 );
and ( n35344 , n30189 , n35048 );
and ( n35345 , n35343 , n35344 );
xor ( n35346 , n35343 , n35344 );
xor ( n35347 , n34634 , n34896 );
and ( n35348 , n30194 , n35048 );
and ( n35349 , n35347 , n35348 );
xor ( n35350 , n35347 , n35348 );
xor ( n35351 , n34638 , n34894 );
and ( n35352 , n30199 , n35048 );
and ( n35353 , n35351 , n35352 );
xor ( n35354 , n35351 , n35352 );
xor ( n35355 , n34642 , n34892 );
and ( n35356 , n30204 , n35048 );
and ( n35357 , n35355 , n35356 );
xor ( n35358 , n35355 , n35356 );
xor ( n35359 , n34646 , n34890 );
and ( n35360 , n30209 , n35048 );
and ( n35361 , n35359 , n35360 );
xor ( n35362 , n35359 , n35360 );
xor ( n35363 , n34650 , n34888 );
and ( n35364 , n30214 , n35048 );
and ( n35365 , n35363 , n35364 );
xor ( n35366 , n35363 , n35364 );
xor ( n35367 , n34654 , n34886 );
and ( n35368 , n30219 , n35048 );
and ( n35369 , n35367 , n35368 );
xor ( n35370 , n35367 , n35368 );
xor ( n35371 , n34658 , n34884 );
and ( n35372 , n30224 , n35048 );
and ( n35373 , n35371 , n35372 );
xor ( n35374 , n35371 , n35372 );
xor ( n35375 , n34662 , n34882 );
and ( n35376 , n30229 , n35048 );
and ( n35377 , n35375 , n35376 );
xor ( n35378 , n35375 , n35376 );
xor ( n35379 , n34666 , n34880 );
and ( n35380 , n30234 , n35048 );
and ( n35381 , n35379 , n35380 );
xor ( n35382 , n35379 , n35380 );
xor ( n35383 , n34670 , n34878 );
and ( n35384 , n30239 , n35048 );
and ( n35385 , n35383 , n35384 );
xor ( n35386 , n35383 , n35384 );
xor ( n35387 , n34674 , n34876 );
and ( n35388 , n30244 , n35048 );
and ( n35389 , n35387 , n35388 );
xor ( n35390 , n35387 , n35388 );
xor ( n35391 , n34678 , n34874 );
and ( n35392 , n30249 , n35048 );
and ( n35393 , n35391 , n35392 );
xor ( n35394 , n35391 , n35392 );
xor ( n35395 , n34682 , n34872 );
and ( n35396 , n30254 , n35048 );
and ( n35397 , n35395 , n35396 );
xor ( n35398 , n35395 , n35396 );
xor ( n35399 , n34686 , n34870 );
and ( n35400 , n30259 , n35048 );
and ( n35401 , n35399 , n35400 );
xor ( n35402 , n35399 , n35400 );
xor ( n35403 , n34690 , n34868 );
and ( n35404 , n30264 , n35048 );
and ( n35405 , n35403 , n35404 );
xor ( n35406 , n35403 , n35404 );
xor ( n35407 , n34694 , n34866 );
and ( n35408 , n30269 , n35048 );
and ( n35409 , n35407 , n35408 );
xor ( n35410 , n35407 , n35408 );
xor ( n35411 , n34698 , n34864 );
and ( n35412 , n30274 , n35048 );
and ( n35413 , n35411 , n35412 );
xor ( n35414 , n35411 , n35412 );
xor ( n35415 , n34702 , n34862 );
and ( n35416 , n30279 , n35048 );
and ( n35417 , n35415 , n35416 );
xor ( n35418 , n35415 , n35416 );
xor ( n35419 , n34706 , n34860 );
and ( n35420 , n30284 , n35048 );
and ( n35421 , n35419 , n35420 );
xor ( n35422 , n35419 , n35420 );
xor ( n35423 , n34710 , n34858 );
and ( n35424 , n30289 , n35048 );
and ( n35425 , n35423 , n35424 );
xor ( n35426 , n35423 , n35424 );
xor ( n35427 , n34714 , n34856 );
and ( n35428 , n30294 , n35048 );
and ( n35429 , n35427 , n35428 );
xor ( n35430 , n35427 , n35428 );
xor ( n35431 , n34718 , n34854 );
and ( n35432 , n30299 , n35048 );
and ( n35433 , n35431 , n35432 );
xor ( n35434 , n35431 , n35432 );
xor ( n35435 , n34722 , n34852 );
and ( n35436 , n30304 , n35048 );
and ( n35437 , n35435 , n35436 );
xor ( n35438 , n35435 , n35436 );
xor ( n35439 , n34726 , n34850 );
and ( n35440 , n30309 , n35048 );
and ( n35441 , n35439 , n35440 );
xor ( n35442 , n35439 , n35440 );
xor ( n35443 , n34730 , n34848 );
and ( n35444 , n30314 , n35048 );
and ( n35445 , n35443 , n35444 );
xor ( n35446 , n35443 , n35444 );
xor ( n35447 , n34734 , n34846 );
and ( n35448 , n30319 , n35048 );
and ( n35449 , n35447 , n35448 );
xor ( n35450 , n35447 , n35448 );
xor ( n35451 , n34738 , n34844 );
and ( n35452 , n30324 , n35048 );
and ( n35453 , n35451 , n35452 );
xor ( n35454 , n35451 , n35452 );
xor ( n35455 , n34742 , n34842 );
and ( n35456 , n30329 , n35048 );
and ( n35457 , n35455 , n35456 );
xor ( n35458 , n35455 , n35456 );
xor ( n35459 , n34746 , n34840 );
and ( n35460 , n30334 , n35048 );
and ( n35461 , n35459 , n35460 );
xor ( n35462 , n35459 , n35460 );
xor ( n35463 , n34750 , n34838 );
and ( n35464 , n30339 , n35048 );
and ( n35465 , n35463 , n35464 );
xor ( n35466 , n35463 , n35464 );
xor ( n35467 , n34754 , n34836 );
and ( n35468 , n30344 , n35048 );
and ( n35469 , n35467 , n35468 );
xor ( n35470 , n35467 , n35468 );
xor ( n35471 , n34758 , n34834 );
and ( n35472 , n30349 , n35048 );
and ( n35473 , n35471 , n35472 );
xor ( n35474 , n35471 , n35472 );
xor ( n35475 , n34762 , n34832 );
and ( n35476 , n30354 , n35048 );
and ( n35477 , n35475 , n35476 );
xor ( n35478 , n35475 , n35476 );
xor ( n35479 , n34766 , n34830 );
and ( n35480 , n30359 , n35048 );
and ( n35481 , n35479 , n35480 );
xor ( n35482 , n35479 , n35480 );
xor ( n35483 , n34770 , n34828 );
and ( n35484 , n30364 , n35048 );
and ( n35485 , n35483 , n35484 );
xor ( n35486 , n35483 , n35484 );
xor ( n35487 , n34774 , n34826 );
and ( n35488 , n30369 , n35048 );
and ( n35489 , n35487 , n35488 );
xor ( n35490 , n35487 , n35488 );
xor ( n35491 , n34778 , n34824 );
and ( n35492 , n30374 , n35048 );
and ( n35493 , n35491 , n35492 );
xor ( n35494 , n35491 , n35492 );
xor ( n35495 , n34782 , n34822 );
and ( n35496 , n30379 , n35048 );
and ( n35497 , n35495 , n35496 );
xor ( n35498 , n35495 , n35496 );
xor ( n35499 , n34786 , n34820 );
and ( n35500 , n30384 , n35048 );
and ( n35501 , n35499 , n35500 );
xor ( n35502 , n35499 , n35500 );
xor ( n35503 , n34790 , n34818 );
and ( n35504 , n30389 , n35048 );
and ( n35505 , n35503 , n35504 );
xor ( n35506 , n35503 , n35504 );
xor ( n35507 , n34794 , n34816 );
and ( n35508 , n30394 , n35048 );
and ( n35509 , n35507 , n35508 );
xor ( n35510 , n35507 , n35508 );
xor ( n35511 , n34798 , n34814 );
and ( n35512 , n30399 , n35048 );
and ( n35513 , n35511 , n35512 );
xor ( n35514 , n35511 , n35512 );
xor ( n35515 , n34802 , n34812 );
and ( n35516 , n30404 , n35048 );
and ( n35517 , n35515 , n35516 );
xor ( n35518 , n35515 , n35516 );
xor ( n35519 , n34806 , n34810 );
and ( n35520 , n30409 , n35048 );
and ( n35521 , n35519 , n35520 );
buf ( n35522 , n35521 );
and ( n35523 , n35518 , n35522 );
or ( n35524 , n35517 , n35523 );
and ( n35525 , n35514 , n35524 );
or ( n35526 , n35513 , n35525 );
and ( n35527 , n35510 , n35526 );
or ( n35528 , n35509 , n35527 );
and ( n35529 , n35506 , n35528 );
or ( n35530 , n35505 , n35529 );
and ( n35531 , n35502 , n35530 );
or ( n35532 , n35501 , n35531 );
and ( n35533 , n35498 , n35532 );
or ( n35534 , n35497 , n35533 );
and ( n35535 , n35494 , n35534 );
or ( n35536 , n35493 , n35535 );
and ( n35537 , n35490 , n35536 );
or ( n35538 , n35489 , n35537 );
and ( n35539 , n35486 , n35538 );
or ( n35540 , n35485 , n35539 );
and ( n35541 , n35482 , n35540 );
or ( n35542 , n35481 , n35541 );
and ( n35543 , n35478 , n35542 );
or ( n35544 , n35477 , n35543 );
and ( n35545 , n35474 , n35544 );
or ( n35546 , n35473 , n35545 );
and ( n35547 , n35470 , n35546 );
or ( n35548 , n35469 , n35547 );
and ( n35549 , n35466 , n35548 );
or ( n35550 , n35465 , n35549 );
and ( n35551 , n35462 , n35550 );
or ( n35552 , n35461 , n35551 );
and ( n35553 , n35458 , n35552 );
or ( n35554 , n35457 , n35553 );
and ( n35555 , n35454 , n35554 );
or ( n35556 , n35453 , n35555 );
and ( n35557 , n35450 , n35556 );
or ( n35558 , n35449 , n35557 );
and ( n35559 , n35446 , n35558 );
or ( n35560 , n35445 , n35559 );
and ( n35561 , n35442 , n35560 );
or ( n35562 , n35441 , n35561 );
and ( n35563 , n35438 , n35562 );
or ( n35564 , n35437 , n35563 );
and ( n35565 , n35434 , n35564 );
or ( n35566 , n35433 , n35565 );
and ( n35567 , n35430 , n35566 );
or ( n35568 , n35429 , n35567 );
and ( n35569 , n35426 , n35568 );
or ( n35570 , n35425 , n35569 );
and ( n35571 , n35422 , n35570 );
or ( n35572 , n35421 , n35571 );
and ( n35573 , n35418 , n35572 );
or ( n35574 , n35417 , n35573 );
and ( n35575 , n35414 , n35574 );
or ( n35576 , n35413 , n35575 );
and ( n35577 , n35410 , n35576 );
or ( n35578 , n35409 , n35577 );
and ( n35579 , n35406 , n35578 );
or ( n35580 , n35405 , n35579 );
and ( n35581 , n35402 , n35580 );
or ( n35582 , n35401 , n35581 );
and ( n35583 , n35398 , n35582 );
or ( n35584 , n35397 , n35583 );
and ( n35585 , n35394 , n35584 );
or ( n35586 , n35393 , n35585 );
and ( n35587 , n35390 , n35586 );
or ( n35588 , n35389 , n35587 );
and ( n35589 , n35386 , n35588 );
or ( n35590 , n35385 , n35589 );
and ( n35591 , n35382 , n35590 );
or ( n35592 , n35381 , n35591 );
and ( n35593 , n35378 , n35592 );
or ( n35594 , n35377 , n35593 );
and ( n35595 , n35374 , n35594 );
or ( n35596 , n35373 , n35595 );
and ( n35597 , n35370 , n35596 );
or ( n35598 , n35369 , n35597 );
and ( n35599 , n35366 , n35598 );
or ( n35600 , n35365 , n35599 );
and ( n35601 , n35362 , n35600 );
or ( n35602 , n35361 , n35601 );
and ( n35603 , n35358 , n35602 );
or ( n35604 , n35357 , n35603 );
and ( n35605 , n35354 , n35604 );
or ( n35606 , n35353 , n35605 );
and ( n35607 , n35350 , n35606 );
or ( n35608 , n35349 , n35607 );
and ( n35609 , n35346 , n35608 );
or ( n35610 , n35345 , n35609 );
and ( n35611 , n35342 , n35610 );
or ( n35612 , n35341 , n35611 );
and ( n35613 , n35338 , n35612 );
or ( n35614 , n35337 , n35613 );
and ( n35615 , n35334 , n35614 );
or ( n35616 , n35333 , n35615 );
and ( n35617 , n35330 , n35616 );
or ( n35618 , n35329 , n35617 );
and ( n35619 , n35326 , n35618 );
or ( n35620 , n35325 , n35619 );
and ( n35621 , n35322 , n35620 );
or ( n35622 , n35321 , n35621 );
and ( n35623 , n35318 , n35622 );
or ( n35624 , n35317 , n35623 );
and ( n35625 , n35314 , n35624 );
or ( n35626 , n35313 , n35625 );
and ( n35627 , n35310 , n35626 );
or ( n35628 , n35309 , n35627 );
and ( n35629 , n35306 , n35628 );
or ( n35630 , n35305 , n35629 );
and ( n35631 , n35302 , n35630 );
or ( n35632 , n35301 , n35631 );
and ( n35633 , n35298 , n35632 );
or ( n35634 , n35297 , n35633 );
and ( n35635 , n35294 , n35634 );
or ( n35636 , n35293 , n35635 );
and ( n35637 , n35290 , n35636 );
or ( n35638 , n35289 , n35637 );
and ( n35639 , n35286 , n35638 );
or ( n35640 , n35285 , n35639 );
and ( n35641 , n35282 , n35640 );
or ( n35642 , n35281 , n35641 );
and ( n35643 , n35278 , n35642 );
or ( n35644 , n35277 , n35643 );
and ( n35645 , n35274 , n35644 );
or ( n35646 , n35273 , n35645 );
and ( n35647 , n35270 , n35646 );
or ( n35648 , n35269 , n35647 );
and ( n35649 , n35266 , n35648 );
or ( n35650 , n35265 , n35649 );
and ( n35651 , n35262 , n35650 );
or ( n35652 , n35261 , n35651 );
and ( n35653 , n35258 , n35652 );
or ( n35654 , n35257 , n35653 );
and ( n35655 , n35254 , n35654 );
or ( n35656 , n35253 , n35655 );
and ( n35657 , n35250 , n35656 );
or ( n35658 , n35249 , n35657 );
and ( n35659 , n35246 , n35658 );
or ( n35660 , n35245 , n35659 );
and ( n35661 , n35242 , n35660 );
or ( n35662 , n35241 , n35661 );
and ( n35663 , n35238 , n35662 );
or ( n35664 , n35237 , n35663 );
and ( n35665 , n35234 , n35664 );
or ( n35666 , n35233 , n35665 );
and ( n35667 , n35230 , n35666 );
or ( n35668 , n35229 , n35667 );
and ( n35669 , n35226 , n35668 );
or ( n35670 , n35225 , n35669 );
and ( n35671 , n35222 , n35670 );
or ( n35672 , n35221 , n35671 );
and ( n35673 , n35218 , n35672 );
or ( n35674 , n35217 , n35673 );
and ( n35675 , n35214 , n35674 );
or ( n35676 , n35213 , n35675 );
and ( n35677 , n35210 , n35676 );
or ( n35678 , n35209 , n35677 );
and ( n35679 , n35206 , n35678 );
or ( n35680 , n35205 , n35679 );
and ( n35681 , n35202 , n35680 );
or ( n35682 , n35201 , n35681 );
and ( n35683 , n35198 , n35682 );
or ( n35684 , n35197 , n35683 );
and ( n35685 , n35194 , n35684 );
or ( n35686 , n35193 , n35685 );
and ( n35687 , n35190 , n35686 );
or ( n35688 , n35189 , n35687 );
and ( n35689 , n35186 , n35688 );
or ( n35690 , n35185 , n35689 );
and ( n35691 , n35182 , n35690 );
or ( n35692 , n35181 , n35691 );
and ( n35693 , n35178 , n35692 );
or ( n35694 , n35177 , n35693 );
and ( n35695 , n35174 , n35694 );
or ( n35696 , n35173 , n35695 );
and ( n35697 , n35170 , n35696 );
or ( n35698 , n35169 , n35697 );
and ( n35699 , n35166 , n35698 );
or ( n35700 , n35165 , n35699 );
and ( n35701 , n35162 , n35700 );
or ( n35702 , n35161 , n35701 );
and ( n35703 , n35158 , n35702 );
or ( n35704 , n35157 , n35703 );
and ( n35705 , n35154 , n35704 );
or ( n35706 , n35153 , n35705 );
and ( n35707 , n35150 , n35706 );
or ( n35708 , n35149 , n35707 );
and ( n35709 , n35146 , n35708 );
or ( n35710 , n35145 , n35709 );
and ( n35711 , n35142 , n35710 );
or ( n35712 , n35141 , n35711 );
and ( n35713 , n35138 , n35712 );
or ( n35714 , n35137 , n35713 );
and ( n35715 , n35134 , n35714 );
or ( n35716 , n35133 , n35715 );
and ( n35717 , n35130 , n35716 );
or ( n35718 , n35129 , n35717 );
and ( n35719 , n35126 , n35718 );
or ( n35720 , n35125 , n35719 );
and ( n35721 , n35122 , n35720 );
or ( n35722 , n35121 , n35721 );
and ( n35723 , n35118 , n35722 );
or ( n35724 , n35117 , n35723 );
and ( n35725 , n35114 , n35724 );
or ( n35726 , n35113 , n35725 );
and ( n35727 , n35110 , n35726 );
or ( n35728 , n35109 , n35727 );
and ( n35729 , n35106 , n35728 );
or ( n35730 , n35105 , n35729 );
and ( n35731 , n35102 , n35730 );
or ( n35732 , n35101 , n35731 );
and ( n35733 , n35098 , n35732 );
or ( n35734 , n35097 , n35733 );
and ( n35735 , n35094 , n35734 );
or ( n35736 , n35093 , n35735 );
and ( n35737 , n35090 , n35736 );
or ( n35738 , n35089 , n35737 );
and ( n35739 , n35086 , n35738 );
or ( n35740 , n35085 , n35739 );
and ( n35741 , n35082 , n35740 );
or ( n35742 , n35081 , n35741 );
and ( n35743 , n35078 , n35742 );
or ( n35744 , n35077 , n35743 );
and ( n35745 , n35074 , n35744 );
or ( n35746 , n35073 , n35745 );
and ( n35747 , n35070 , n35746 );
or ( n35748 , n35069 , n35747 );
and ( n35749 , n35066 , n35748 );
or ( n35750 , n35065 , n35749 );
and ( n35751 , n35062 , n35750 );
or ( n35752 , n35061 , n35751 );
and ( n35753 , n35058 , n35752 );
or ( n35754 , n35057 , n35753 );
and ( n35755 , n35054 , n35754 );
or ( n35756 , n35053 , n35755 );
xor ( n35757 , n35050 , n35756 );
buf ( n35758 , n18088 );
and ( n35759 , n29824 , n35758 );
xor ( n35760 , n35757 , n35759 );
xor ( n35761 , n35054 , n35754 );
and ( n35762 , n29829 , n35758 );
and ( n35763 , n35761 , n35762 );
xor ( n35764 , n35761 , n35762 );
xor ( n35765 , n35058 , n35752 );
and ( n35766 , n29834 , n35758 );
and ( n35767 , n35765 , n35766 );
xor ( n35768 , n35765 , n35766 );
xor ( n35769 , n35062 , n35750 );
and ( n35770 , n29839 , n35758 );
and ( n35771 , n35769 , n35770 );
xor ( n35772 , n35769 , n35770 );
xor ( n35773 , n35066 , n35748 );
and ( n35774 , n29844 , n35758 );
and ( n35775 , n35773 , n35774 );
xor ( n35776 , n35773 , n35774 );
xor ( n35777 , n35070 , n35746 );
and ( n35778 , n29849 , n35758 );
and ( n35779 , n35777 , n35778 );
xor ( n35780 , n35777 , n35778 );
xor ( n35781 , n35074 , n35744 );
and ( n35782 , n29854 , n35758 );
and ( n35783 , n35781 , n35782 );
xor ( n35784 , n35781 , n35782 );
xor ( n35785 , n35078 , n35742 );
and ( n35786 , n29859 , n35758 );
and ( n35787 , n35785 , n35786 );
xor ( n35788 , n35785 , n35786 );
xor ( n35789 , n35082 , n35740 );
and ( n35790 , n29864 , n35758 );
and ( n35791 , n35789 , n35790 );
xor ( n35792 , n35789 , n35790 );
xor ( n35793 , n35086 , n35738 );
and ( n35794 , n29869 , n35758 );
and ( n35795 , n35793 , n35794 );
xor ( n35796 , n35793 , n35794 );
xor ( n35797 , n35090 , n35736 );
and ( n35798 , n29874 , n35758 );
and ( n35799 , n35797 , n35798 );
xor ( n35800 , n35797 , n35798 );
xor ( n35801 , n35094 , n35734 );
and ( n35802 , n29879 , n35758 );
and ( n35803 , n35801 , n35802 );
xor ( n35804 , n35801 , n35802 );
xor ( n35805 , n35098 , n35732 );
and ( n35806 , n29884 , n35758 );
and ( n35807 , n35805 , n35806 );
xor ( n35808 , n35805 , n35806 );
xor ( n35809 , n35102 , n35730 );
and ( n35810 , n29889 , n35758 );
and ( n35811 , n35809 , n35810 );
xor ( n35812 , n35809 , n35810 );
xor ( n35813 , n35106 , n35728 );
and ( n35814 , n29894 , n35758 );
and ( n35815 , n35813 , n35814 );
xor ( n35816 , n35813 , n35814 );
xor ( n35817 , n35110 , n35726 );
and ( n35818 , n29899 , n35758 );
and ( n35819 , n35817 , n35818 );
xor ( n35820 , n35817 , n35818 );
xor ( n35821 , n35114 , n35724 );
and ( n35822 , n29904 , n35758 );
and ( n35823 , n35821 , n35822 );
xor ( n35824 , n35821 , n35822 );
xor ( n35825 , n35118 , n35722 );
and ( n35826 , n29909 , n35758 );
and ( n35827 , n35825 , n35826 );
xor ( n35828 , n35825 , n35826 );
xor ( n35829 , n35122 , n35720 );
and ( n35830 , n29914 , n35758 );
and ( n35831 , n35829 , n35830 );
xor ( n35832 , n35829 , n35830 );
xor ( n35833 , n35126 , n35718 );
and ( n35834 , n29919 , n35758 );
and ( n35835 , n35833 , n35834 );
xor ( n35836 , n35833 , n35834 );
xor ( n35837 , n35130 , n35716 );
and ( n35838 , n29924 , n35758 );
and ( n35839 , n35837 , n35838 );
xor ( n35840 , n35837 , n35838 );
xor ( n35841 , n35134 , n35714 );
and ( n35842 , n29929 , n35758 );
and ( n35843 , n35841 , n35842 );
xor ( n35844 , n35841 , n35842 );
xor ( n35845 , n35138 , n35712 );
and ( n35846 , n29934 , n35758 );
and ( n35847 , n35845 , n35846 );
xor ( n35848 , n35845 , n35846 );
xor ( n35849 , n35142 , n35710 );
and ( n35850 , n29939 , n35758 );
and ( n35851 , n35849 , n35850 );
xor ( n35852 , n35849 , n35850 );
xor ( n35853 , n35146 , n35708 );
and ( n35854 , n29944 , n35758 );
and ( n35855 , n35853 , n35854 );
xor ( n35856 , n35853 , n35854 );
xor ( n35857 , n35150 , n35706 );
and ( n35858 , n29949 , n35758 );
and ( n35859 , n35857 , n35858 );
xor ( n35860 , n35857 , n35858 );
xor ( n35861 , n35154 , n35704 );
and ( n35862 , n29954 , n35758 );
and ( n35863 , n35861 , n35862 );
xor ( n35864 , n35861 , n35862 );
xor ( n35865 , n35158 , n35702 );
and ( n35866 , n29959 , n35758 );
and ( n35867 , n35865 , n35866 );
xor ( n35868 , n35865 , n35866 );
xor ( n35869 , n35162 , n35700 );
and ( n35870 , n29964 , n35758 );
and ( n35871 , n35869 , n35870 );
xor ( n35872 , n35869 , n35870 );
xor ( n35873 , n35166 , n35698 );
and ( n35874 , n29969 , n35758 );
and ( n35875 , n35873 , n35874 );
xor ( n35876 , n35873 , n35874 );
xor ( n35877 , n35170 , n35696 );
and ( n35878 , n29974 , n35758 );
and ( n35879 , n35877 , n35878 );
xor ( n35880 , n35877 , n35878 );
xor ( n35881 , n35174 , n35694 );
and ( n35882 , n29979 , n35758 );
and ( n35883 , n35881 , n35882 );
xor ( n35884 , n35881 , n35882 );
xor ( n35885 , n35178 , n35692 );
and ( n35886 , n29984 , n35758 );
and ( n35887 , n35885 , n35886 );
xor ( n35888 , n35885 , n35886 );
xor ( n35889 , n35182 , n35690 );
and ( n35890 , n29989 , n35758 );
and ( n35891 , n35889 , n35890 );
xor ( n35892 , n35889 , n35890 );
xor ( n35893 , n35186 , n35688 );
and ( n35894 , n29994 , n35758 );
and ( n35895 , n35893 , n35894 );
xor ( n35896 , n35893 , n35894 );
xor ( n35897 , n35190 , n35686 );
and ( n35898 , n29999 , n35758 );
and ( n35899 , n35897 , n35898 );
xor ( n35900 , n35897 , n35898 );
xor ( n35901 , n35194 , n35684 );
and ( n35902 , n30004 , n35758 );
and ( n35903 , n35901 , n35902 );
xor ( n35904 , n35901 , n35902 );
xor ( n35905 , n35198 , n35682 );
and ( n35906 , n30009 , n35758 );
and ( n35907 , n35905 , n35906 );
xor ( n35908 , n35905 , n35906 );
xor ( n35909 , n35202 , n35680 );
and ( n35910 , n30014 , n35758 );
and ( n35911 , n35909 , n35910 );
xor ( n35912 , n35909 , n35910 );
xor ( n35913 , n35206 , n35678 );
and ( n35914 , n30019 , n35758 );
and ( n35915 , n35913 , n35914 );
xor ( n35916 , n35913 , n35914 );
xor ( n35917 , n35210 , n35676 );
and ( n35918 , n30024 , n35758 );
and ( n35919 , n35917 , n35918 );
xor ( n35920 , n35917 , n35918 );
xor ( n35921 , n35214 , n35674 );
and ( n35922 , n30029 , n35758 );
and ( n35923 , n35921 , n35922 );
xor ( n35924 , n35921 , n35922 );
xor ( n35925 , n35218 , n35672 );
and ( n35926 , n30034 , n35758 );
and ( n35927 , n35925 , n35926 );
xor ( n35928 , n35925 , n35926 );
xor ( n35929 , n35222 , n35670 );
and ( n35930 , n30039 , n35758 );
and ( n35931 , n35929 , n35930 );
xor ( n35932 , n35929 , n35930 );
xor ( n35933 , n35226 , n35668 );
and ( n35934 , n30044 , n35758 );
and ( n35935 , n35933 , n35934 );
xor ( n35936 , n35933 , n35934 );
xor ( n35937 , n35230 , n35666 );
and ( n35938 , n30049 , n35758 );
and ( n35939 , n35937 , n35938 );
xor ( n35940 , n35937 , n35938 );
xor ( n35941 , n35234 , n35664 );
and ( n35942 , n30054 , n35758 );
and ( n35943 , n35941 , n35942 );
xor ( n35944 , n35941 , n35942 );
xor ( n35945 , n35238 , n35662 );
and ( n35946 , n30059 , n35758 );
and ( n35947 , n35945 , n35946 );
xor ( n35948 , n35945 , n35946 );
xor ( n35949 , n35242 , n35660 );
and ( n35950 , n30064 , n35758 );
and ( n35951 , n35949 , n35950 );
xor ( n35952 , n35949 , n35950 );
xor ( n35953 , n35246 , n35658 );
and ( n35954 , n30069 , n35758 );
and ( n35955 , n35953 , n35954 );
xor ( n35956 , n35953 , n35954 );
xor ( n35957 , n35250 , n35656 );
and ( n35958 , n30074 , n35758 );
and ( n35959 , n35957 , n35958 );
xor ( n35960 , n35957 , n35958 );
xor ( n35961 , n35254 , n35654 );
and ( n35962 , n30079 , n35758 );
and ( n35963 , n35961 , n35962 );
xor ( n35964 , n35961 , n35962 );
xor ( n35965 , n35258 , n35652 );
and ( n35966 , n30084 , n35758 );
and ( n35967 , n35965 , n35966 );
xor ( n35968 , n35965 , n35966 );
xor ( n35969 , n35262 , n35650 );
and ( n35970 , n30089 , n35758 );
and ( n35971 , n35969 , n35970 );
xor ( n35972 , n35969 , n35970 );
xor ( n35973 , n35266 , n35648 );
and ( n35974 , n30094 , n35758 );
and ( n35975 , n35973 , n35974 );
xor ( n35976 , n35973 , n35974 );
xor ( n35977 , n35270 , n35646 );
and ( n35978 , n30099 , n35758 );
and ( n35979 , n35977 , n35978 );
xor ( n35980 , n35977 , n35978 );
xor ( n35981 , n35274 , n35644 );
and ( n35982 , n30104 , n35758 );
and ( n35983 , n35981 , n35982 );
xor ( n35984 , n35981 , n35982 );
xor ( n35985 , n35278 , n35642 );
and ( n35986 , n30109 , n35758 );
and ( n35987 , n35985 , n35986 );
xor ( n35988 , n35985 , n35986 );
xor ( n35989 , n35282 , n35640 );
and ( n35990 , n30114 , n35758 );
and ( n35991 , n35989 , n35990 );
xor ( n35992 , n35989 , n35990 );
xor ( n35993 , n35286 , n35638 );
and ( n35994 , n30119 , n35758 );
and ( n35995 , n35993 , n35994 );
xor ( n35996 , n35993 , n35994 );
xor ( n35997 , n35290 , n35636 );
and ( n35998 , n30124 , n35758 );
and ( n35999 , n35997 , n35998 );
xor ( n36000 , n35997 , n35998 );
xor ( n36001 , n35294 , n35634 );
and ( n36002 , n30129 , n35758 );
and ( n36003 , n36001 , n36002 );
xor ( n36004 , n36001 , n36002 );
xor ( n36005 , n35298 , n35632 );
and ( n36006 , n30134 , n35758 );
and ( n36007 , n36005 , n36006 );
xor ( n36008 , n36005 , n36006 );
xor ( n36009 , n35302 , n35630 );
and ( n36010 , n30139 , n35758 );
and ( n36011 , n36009 , n36010 );
xor ( n36012 , n36009 , n36010 );
xor ( n36013 , n35306 , n35628 );
and ( n36014 , n30144 , n35758 );
and ( n36015 , n36013 , n36014 );
xor ( n36016 , n36013 , n36014 );
xor ( n36017 , n35310 , n35626 );
and ( n36018 , n30149 , n35758 );
and ( n36019 , n36017 , n36018 );
xor ( n36020 , n36017 , n36018 );
xor ( n36021 , n35314 , n35624 );
and ( n36022 , n30154 , n35758 );
and ( n36023 , n36021 , n36022 );
xor ( n36024 , n36021 , n36022 );
xor ( n36025 , n35318 , n35622 );
and ( n36026 , n30159 , n35758 );
and ( n36027 , n36025 , n36026 );
xor ( n36028 , n36025 , n36026 );
xor ( n36029 , n35322 , n35620 );
and ( n36030 , n30164 , n35758 );
and ( n36031 , n36029 , n36030 );
xor ( n36032 , n36029 , n36030 );
xor ( n36033 , n35326 , n35618 );
and ( n36034 , n30169 , n35758 );
and ( n36035 , n36033 , n36034 );
xor ( n36036 , n36033 , n36034 );
xor ( n36037 , n35330 , n35616 );
and ( n36038 , n30174 , n35758 );
and ( n36039 , n36037 , n36038 );
xor ( n36040 , n36037 , n36038 );
xor ( n36041 , n35334 , n35614 );
and ( n36042 , n30179 , n35758 );
and ( n36043 , n36041 , n36042 );
xor ( n36044 , n36041 , n36042 );
xor ( n36045 , n35338 , n35612 );
and ( n36046 , n30184 , n35758 );
and ( n36047 , n36045 , n36046 );
xor ( n36048 , n36045 , n36046 );
xor ( n36049 , n35342 , n35610 );
and ( n36050 , n30189 , n35758 );
and ( n36051 , n36049 , n36050 );
xor ( n36052 , n36049 , n36050 );
xor ( n36053 , n35346 , n35608 );
and ( n36054 , n30194 , n35758 );
and ( n36055 , n36053 , n36054 );
xor ( n36056 , n36053 , n36054 );
xor ( n36057 , n35350 , n35606 );
and ( n36058 , n30199 , n35758 );
and ( n36059 , n36057 , n36058 );
xor ( n36060 , n36057 , n36058 );
xor ( n36061 , n35354 , n35604 );
and ( n36062 , n30204 , n35758 );
and ( n36063 , n36061 , n36062 );
xor ( n36064 , n36061 , n36062 );
xor ( n36065 , n35358 , n35602 );
and ( n36066 , n30209 , n35758 );
and ( n36067 , n36065 , n36066 );
xor ( n36068 , n36065 , n36066 );
xor ( n36069 , n35362 , n35600 );
and ( n36070 , n30214 , n35758 );
and ( n36071 , n36069 , n36070 );
xor ( n36072 , n36069 , n36070 );
xor ( n36073 , n35366 , n35598 );
and ( n36074 , n30219 , n35758 );
and ( n36075 , n36073 , n36074 );
xor ( n36076 , n36073 , n36074 );
xor ( n36077 , n35370 , n35596 );
and ( n36078 , n30224 , n35758 );
and ( n36079 , n36077 , n36078 );
xor ( n36080 , n36077 , n36078 );
xor ( n36081 , n35374 , n35594 );
and ( n36082 , n30229 , n35758 );
and ( n36083 , n36081 , n36082 );
xor ( n36084 , n36081 , n36082 );
xor ( n36085 , n35378 , n35592 );
and ( n36086 , n30234 , n35758 );
and ( n36087 , n36085 , n36086 );
xor ( n36088 , n36085 , n36086 );
xor ( n36089 , n35382 , n35590 );
and ( n36090 , n30239 , n35758 );
and ( n36091 , n36089 , n36090 );
xor ( n36092 , n36089 , n36090 );
xor ( n36093 , n35386 , n35588 );
and ( n36094 , n30244 , n35758 );
and ( n36095 , n36093 , n36094 );
xor ( n36096 , n36093 , n36094 );
xor ( n36097 , n35390 , n35586 );
and ( n36098 , n30249 , n35758 );
and ( n36099 , n36097 , n36098 );
xor ( n36100 , n36097 , n36098 );
xor ( n36101 , n35394 , n35584 );
and ( n36102 , n30254 , n35758 );
and ( n36103 , n36101 , n36102 );
xor ( n36104 , n36101 , n36102 );
xor ( n36105 , n35398 , n35582 );
and ( n36106 , n30259 , n35758 );
and ( n36107 , n36105 , n36106 );
xor ( n36108 , n36105 , n36106 );
xor ( n36109 , n35402 , n35580 );
and ( n36110 , n30264 , n35758 );
and ( n36111 , n36109 , n36110 );
xor ( n36112 , n36109 , n36110 );
xor ( n36113 , n35406 , n35578 );
and ( n36114 , n30269 , n35758 );
and ( n36115 , n36113 , n36114 );
xor ( n36116 , n36113 , n36114 );
xor ( n36117 , n35410 , n35576 );
and ( n36118 , n30274 , n35758 );
and ( n36119 , n36117 , n36118 );
xor ( n36120 , n36117 , n36118 );
xor ( n36121 , n35414 , n35574 );
and ( n36122 , n30279 , n35758 );
and ( n36123 , n36121 , n36122 );
xor ( n36124 , n36121 , n36122 );
xor ( n36125 , n35418 , n35572 );
and ( n36126 , n30284 , n35758 );
and ( n36127 , n36125 , n36126 );
xor ( n36128 , n36125 , n36126 );
xor ( n36129 , n35422 , n35570 );
and ( n36130 , n30289 , n35758 );
and ( n36131 , n36129 , n36130 );
xor ( n36132 , n36129 , n36130 );
xor ( n36133 , n35426 , n35568 );
and ( n36134 , n30294 , n35758 );
and ( n36135 , n36133 , n36134 );
xor ( n36136 , n36133 , n36134 );
xor ( n36137 , n35430 , n35566 );
and ( n36138 , n30299 , n35758 );
and ( n36139 , n36137 , n36138 );
xor ( n36140 , n36137 , n36138 );
xor ( n36141 , n35434 , n35564 );
and ( n36142 , n30304 , n35758 );
and ( n36143 , n36141 , n36142 );
xor ( n36144 , n36141 , n36142 );
xor ( n36145 , n35438 , n35562 );
and ( n36146 , n30309 , n35758 );
and ( n36147 , n36145 , n36146 );
xor ( n36148 , n36145 , n36146 );
xor ( n36149 , n35442 , n35560 );
and ( n36150 , n30314 , n35758 );
and ( n36151 , n36149 , n36150 );
xor ( n36152 , n36149 , n36150 );
xor ( n36153 , n35446 , n35558 );
and ( n36154 , n30319 , n35758 );
and ( n36155 , n36153 , n36154 );
xor ( n36156 , n36153 , n36154 );
xor ( n36157 , n35450 , n35556 );
and ( n36158 , n30324 , n35758 );
and ( n36159 , n36157 , n36158 );
xor ( n36160 , n36157 , n36158 );
xor ( n36161 , n35454 , n35554 );
and ( n36162 , n30329 , n35758 );
and ( n36163 , n36161 , n36162 );
xor ( n36164 , n36161 , n36162 );
xor ( n36165 , n35458 , n35552 );
and ( n36166 , n30334 , n35758 );
and ( n36167 , n36165 , n36166 );
xor ( n36168 , n36165 , n36166 );
xor ( n36169 , n35462 , n35550 );
and ( n36170 , n30339 , n35758 );
and ( n36171 , n36169 , n36170 );
xor ( n36172 , n36169 , n36170 );
xor ( n36173 , n35466 , n35548 );
and ( n36174 , n30344 , n35758 );
and ( n36175 , n36173 , n36174 );
xor ( n36176 , n36173 , n36174 );
xor ( n36177 , n35470 , n35546 );
and ( n36178 , n30349 , n35758 );
and ( n36179 , n36177 , n36178 );
xor ( n36180 , n36177 , n36178 );
xor ( n36181 , n35474 , n35544 );
and ( n36182 , n30354 , n35758 );
and ( n36183 , n36181 , n36182 );
xor ( n36184 , n36181 , n36182 );
xor ( n36185 , n35478 , n35542 );
and ( n36186 , n30359 , n35758 );
and ( n36187 , n36185 , n36186 );
xor ( n36188 , n36185 , n36186 );
xor ( n36189 , n35482 , n35540 );
and ( n36190 , n30364 , n35758 );
and ( n36191 , n36189 , n36190 );
xor ( n36192 , n36189 , n36190 );
xor ( n36193 , n35486 , n35538 );
and ( n36194 , n30369 , n35758 );
and ( n36195 , n36193 , n36194 );
xor ( n36196 , n36193 , n36194 );
xor ( n36197 , n35490 , n35536 );
and ( n36198 , n30374 , n35758 );
and ( n36199 , n36197 , n36198 );
xor ( n36200 , n36197 , n36198 );
xor ( n36201 , n35494 , n35534 );
and ( n36202 , n30379 , n35758 );
and ( n36203 , n36201 , n36202 );
xor ( n36204 , n36201 , n36202 );
xor ( n36205 , n35498 , n35532 );
and ( n36206 , n30384 , n35758 );
and ( n36207 , n36205 , n36206 );
xor ( n36208 , n36205 , n36206 );
xor ( n36209 , n35502 , n35530 );
and ( n36210 , n30389 , n35758 );
and ( n36211 , n36209 , n36210 );
xor ( n36212 , n36209 , n36210 );
xor ( n36213 , n35506 , n35528 );
and ( n36214 , n30394 , n35758 );
and ( n36215 , n36213 , n36214 );
xor ( n36216 , n36213 , n36214 );
xor ( n36217 , n35510 , n35526 );
and ( n36218 , n30399 , n35758 );
and ( n36219 , n36217 , n36218 );
xor ( n36220 , n36217 , n36218 );
xor ( n36221 , n35514 , n35524 );
and ( n36222 , n30404 , n35758 );
and ( n36223 , n36221 , n36222 );
xor ( n36224 , n36221 , n36222 );
xor ( n36225 , n35518 , n35522 );
and ( n36226 , n30409 , n35758 );
and ( n36227 , n36225 , n36226 );
buf ( n36228 , n36227 );
and ( n36229 , n36224 , n36228 );
or ( n36230 , n36223 , n36229 );
and ( n36231 , n36220 , n36230 );
or ( n36232 , n36219 , n36231 );
and ( n36233 , n36216 , n36232 );
or ( n36234 , n36215 , n36233 );
and ( n36235 , n36212 , n36234 );
or ( n36236 , n36211 , n36235 );
and ( n36237 , n36208 , n36236 );
or ( n36238 , n36207 , n36237 );
and ( n36239 , n36204 , n36238 );
or ( n36240 , n36203 , n36239 );
and ( n36241 , n36200 , n36240 );
or ( n36242 , n36199 , n36241 );
and ( n36243 , n36196 , n36242 );
or ( n36244 , n36195 , n36243 );
and ( n36245 , n36192 , n36244 );
or ( n36246 , n36191 , n36245 );
and ( n36247 , n36188 , n36246 );
or ( n36248 , n36187 , n36247 );
and ( n36249 , n36184 , n36248 );
or ( n36250 , n36183 , n36249 );
and ( n36251 , n36180 , n36250 );
or ( n36252 , n36179 , n36251 );
and ( n36253 , n36176 , n36252 );
or ( n36254 , n36175 , n36253 );
and ( n36255 , n36172 , n36254 );
or ( n36256 , n36171 , n36255 );
and ( n36257 , n36168 , n36256 );
or ( n36258 , n36167 , n36257 );
and ( n36259 , n36164 , n36258 );
or ( n36260 , n36163 , n36259 );
and ( n36261 , n36160 , n36260 );
or ( n36262 , n36159 , n36261 );
and ( n36263 , n36156 , n36262 );
or ( n36264 , n36155 , n36263 );
and ( n36265 , n36152 , n36264 );
or ( n36266 , n36151 , n36265 );
and ( n36267 , n36148 , n36266 );
or ( n36268 , n36147 , n36267 );
and ( n36269 , n36144 , n36268 );
or ( n36270 , n36143 , n36269 );
and ( n36271 , n36140 , n36270 );
or ( n36272 , n36139 , n36271 );
and ( n36273 , n36136 , n36272 );
or ( n36274 , n36135 , n36273 );
and ( n36275 , n36132 , n36274 );
or ( n36276 , n36131 , n36275 );
and ( n36277 , n36128 , n36276 );
or ( n36278 , n36127 , n36277 );
and ( n36279 , n36124 , n36278 );
or ( n36280 , n36123 , n36279 );
and ( n36281 , n36120 , n36280 );
or ( n36282 , n36119 , n36281 );
and ( n36283 , n36116 , n36282 );
or ( n36284 , n36115 , n36283 );
and ( n36285 , n36112 , n36284 );
or ( n36286 , n36111 , n36285 );
and ( n36287 , n36108 , n36286 );
or ( n36288 , n36107 , n36287 );
and ( n36289 , n36104 , n36288 );
or ( n36290 , n36103 , n36289 );
and ( n36291 , n36100 , n36290 );
or ( n36292 , n36099 , n36291 );
and ( n36293 , n36096 , n36292 );
or ( n36294 , n36095 , n36293 );
and ( n36295 , n36092 , n36294 );
or ( n36296 , n36091 , n36295 );
and ( n36297 , n36088 , n36296 );
or ( n36298 , n36087 , n36297 );
and ( n36299 , n36084 , n36298 );
or ( n36300 , n36083 , n36299 );
and ( n36301 , n36080 , n36300 );
or ( n36302 , n36079 , n36301 );
and ( n36303 , n36076 , n36302 );
or ( n36304 , n36075 , n36303 );
and ( n36305 , n36072 , n36304 );
or ( n36306 , n36071 , n36305 );
and ( n36307 , n36068 , n36306 );
or ( n36308 , n36067 , n36307 );
and ( n36309 , n36064 , n36308 );
or ( n36310 , n36063 , n36309 );
and ( n36311 , n36060 , n36310 );
or ( n36312 , n36059 , n36311 );
and ( n36313 , n36056 , n36312 );
or ( n36314 , n36055 , n36313 );
and ( n36315 , n36052 , n36314 );
or ( n36316 , n36051 , n36315 );
and ( n36317 , n36048 , n36316 );
or ( n36318 , n36047 , n36317 );
and ( n36319 , n36044 , n36318 );
or ( n36320 , n36043 , n36319 );
and ( n36321 , n36040 , n36320 );
or ( n36322 , n36039 , n36321 );
and ( n36323 , n36036 , n36322 );
or ( n36324 , n36035 , n36323 );
and ( n36325 , n36032 , n36324 );
or ( n36326 , n36031 , n36325 );
and ( n36327 , n36028 , n36326 );
or ( n36328 , n36027 , n36327 );
and ( n36329 , n36024 , n36328 );
or ( n36330 , n36023 , n36329 );
and ( n36331 , n36020 , n36330 );
or ( n36332 , n36019 , n36331 );
and ( n36333 , n36016 , n36332 );
or ( n36334 , n36015 , n36333 );
and ( n36335 , n36012 , n36334 );
or ( n36336 , n36011 , n36335 );
and ( n36337 , n36008 , n36336 );
or ( n36338 , n36007 , n36337 );
and ( n36339 , n36004 , n36338 );
or ( n36340 , n36003 , n36339 );
and ( n36341 , n36000 , n36340 );
or ( n36342 , n35999 , n36341 );
and ( n36343 , n35996 , n36342 );
or ( n36344 , n35995 , n36343 );
and ( n36345 , n35992 , n36344 );
or ( n36346 , n35991 , n36345 );
and ( n36347 , n35988 , n36346 );
or ( n36348 , n35987 , n36347 );
and ( n36349 , n35984 , n36348 );
or ( n36350 , n35983 , n36349 );
and ( n36351 , n35980 , n36350 );
or ( n36352 , n35979 , n36351 );
and ( n36353 , n35976 , n36352 );
or ( n36354 , n35975 , n36353 );
and ( n36355 , n35972 , n36354 );
or ( n36356 , n35971 , n36355 );
and ( n36357 , n35968 , n36356 );
or ( n36358 , n35967 , n36357 );
and ( n36359 , n35964 , n36358 );
or ( n36360 , n35963 , n36359 );
and ( n36361 , n35960 , n36360 );
or ( n36362 , n35959 , n36361 );
and ( n36363 , n35956 , n36362 );
or ( n36364 , n35955 , n36363 );
and ( n36365 , n35952 , n36364 );
or ( n36366 , n35951 , n36365 );
and ( n36367 , n35948 , n36366 );
or ( n36368 , n35947 , n36367 );
and ( n36369 , n35944 , n36368 );
or ( n36370 , n35943 , n36369 );
and ( n36371 , n35940 , n36370 );
or ( n36372 , n35939 , n36371 );
and ( n36373 , n35936 , n36372 );
or ( n36374 , n35935 , n36373 );
and ( n36375 , n35932 , n36374 );
or ( n36376 , n35931 , n36375 );
and ( n36377 , n35928 , n36376 );
or ( n36378 , n35927 , n36377 );
and ( n36379 , n35924 , n36378 );
or ( n36380 , n35923 , n36379 );
and ( n36381 , n35920 , n36380 );
or ( n36382 , n35919 , n36381 );
and ( n36383 , n35916 , n36382 );
or ( n36384 , n35915 , n36383 );
and ( n36385 , n35912 , n36384 );
or ( n36386 , n35911 , n36385 );
and ( n36387 , n35908 , n36386 );
or ( n36388 , n35907 , n36387 );
and ( n36389 , n35904 , n36388 );
or ( n36390 , n35903 , n36389 );
and ( n36391 , n35900 , n36390 );
or ( n36392 , n35899 , n36391 );
and ( n36393 , n35896 , n36392 );
or ( n36394 , n35895 , n36393 );
and ( n36395 , n35892 , n36394 );
or ( n36396 , n35891 , n36395 );
and ( n36397 , n35888 , n36396 );
or ( n36398 , n35887 , n36397 );
and ( n36399 , n35884 , n36398 );
or ( n36400 , n35883 , n36399 );
and ( n36401 , n35880 , n36400 );
or ( n36402 , n35879 , n36401 );
and ( n36403 , n35876 , n36402 );
or ( n36404 , n35875 , n36403 );
and ( n36405 , n35872 , n36404 );
or ( n36406 , n35871 , n36405 );
and ( n36407 , n35868 , n36406 );
or ( n36408 , n35867 , n36407 );
and ( n36409 , n35864 , n36408 );
or ( n36410 , n35863 , n36409 );
and ( n36411 , n35860 , n36410 );
or ( n36412 , n35859 , n36411 );
and ( n36413 , n35856 , n36412 );
or ( n36414 , n35855 , n36413 );
and ( n36415 , n35852 , n36414 );
or ( n36416 , n35851 , n36415 );
and ( n36417 , n35848 , n36416 );
or ( n36418 , n35847 , n36417 );
and ( n36419 , n35844 , n36418 );
or ( n36420 , n35843 , n36419 );
and ( n36421 , n35840 , n36420 );
or ( n36422 , n35839 , n36421 );
and ( n36423 , n35836 , n36422 );
or ( n36424 , n35835 , n36423 );
and ( n36425 , n35832 , n36424 );
or ( n36426 , n35831 , n36425 );
and ( n36427 , n35828 , n36426 );
or ( n36428 , n35827 , n36427 );
and ( n36429 , n35824 , n36428 );
or ( n36430 , n35823 , n36429 );
and ( n36431 , n35820 , n36430 );
or ( n36432 , n35819 , n36431 );
and ( n36433 , n35816 , n36432 );
or ( n36434 , n35815 , n36433 );
and ( n36435 , n35812 , n36434 );
or ( n36436 , n35811 , n36435 );
and ( n36437 , n35808 , n36436 );
or ( n36438 , n35807 , n36437 );
and ( n36439 , n35804 , n36438 );
or ( n36440 , n35803 , n36439 );
and ( n36441 , n35800 , n36440 );
or ( n36442 , n35799 , n36441 );
and ( n36443 , n35796 , n36442 );
or ( n36444 , n35795 , n36443 );
and ( n36445 , n35792 , n36444 );
or ( n36446 , n35791 , n36445 );
and ( n36447 , n35788 , n36446 );
or ( n36448 , n35787 , n36447 );
and ( n36449 , n35784 , n36448 );
or ( n36450 , n35783 , n36449 );
and ( n36451 , n35780 , n36450 );
or ( n36452 , n35779 , n36451 );
and ( n36453 , n35776 , n36452 );
or ( n36454 , n35775 , n36453 );
and ( n36455 , n35772 , n36454 );
or ( n36456 , n35771 , n36455 );
and ( n36457 , n35768 , n36456 );
or ( n36458 , n35767 , n36457 );
and ( n36459 , n35764 , n36458 );
or ( n36460 , n35763 , n36459 );
xor ( n36461 , n35760 , n36460 );
buf ( n36462 , n18086 );
and ( n36463 , n29829 , n36462 );
xor ( n36464 , n36461 , n36463 );
xor ( n36465 , n35764 , n36458 );
and ( n36466 , n29834 , n36462 );
and ( n36467 , n36465 , n36466 );
xor ( n36468 , n36465 , n36466 );
xor ( n36469 , n35768 , n36456 );
and ( n36470 , n29839 , n36462 );
and ( n36471 , n36469 , n36470 );
xor ( n36472 , n36469 , n36470 );
xor ( n36473 , n35772 , n36454 );
and ( n36474 , n29844 , n36462 );
and ( n36475 , n36473 , n36474 );
xor ( n36476 , n36473 , n36474 );
xor ( n36477 , n35776 , n36452 );
and ( n36478 , n29849 , n36462 );
and ( n36479 , n36477 , n36478 );
xor ( n36480 , n36477 , n36478 );
xor ( n36481 , n35780 , n36450 );
and ( n36482 , n29854 , n36462 );
and ( n36483 , n36481 , n36482 );
xor ( n36484 , n36481 , n36482 );
xor ( n36485 , n35784 , n36448 );
and ( n36486 , n29859 , n36462 );
and ( n36487 , n36485 , n36486 );
xor ( n36488 , n36485 , n36486 );
xor ( n36489 , n35788 , n36446 );
and ( n36490 , n29864 , n36462 );
and ( n36491 , n36489 , n36490 );
xor ( n36492 , n36489 , n36490 );
xor ( n36493 , n35792 , n36444 );
and ( n36494 , n29869 , n36462 );
and ( n36495 , n36493 , n36494 );
xor ( n36496 , n36493 , n36494 );
xor ( n36497 , n35796 , n36442 );
and ( n36498 , n29874 , n36462 );
and ( n36499 , n36497 , n36498 );
xor ( n36500 , n36497 , n36498 );
xor ( n36501 , n35800 , n36440 );
and ( n36502 , n29879 , n36462 );
and ( n36503 , n36501 , n36502 );
xor ( n36504 , n36501 , n36502 );
xor ( n36505 , n35804 , n36438 );
and ( n36506 , n29884 , n36462 );
and ( n36507 , n36505 , n36506 );
xor ( n36508 , n36505 , n36506 );
xor ( n36509 , n35808 , n36436 );
and ( n36510 , n29889 , n36462 );
and ( n36511 , n36509 , n36510 );
xor ( n36512 , n36509 , n36510 );
xor ( n36513 , n35812 , n36434 );
and ( n36514 , n29894 , n36462 );
and ( n36515 , n36513 , n36514 );
xor ( n36516 , n36513 , n36514 );
xor ( n36517 , n35816 , n36432 );
and ( n36518 , n29899 , n36462 );
and ( n36519 , n36517 , n36518 );
xor ( n36520 , n36517 , n36518 );
xor ( n36521 , n35820 , n36430 );
and ( n36522 , n29904 , n36462 );
and ( n36523 , n36521 , n36522 );
xor ( n36524 , n36521 , n36522 );
xor ( n36525 , n35824 , n36428 );
and ( n36526 , n29909 , n36462 );
and ( n36527 , n36525 , n36526 );
xor ( n36528 , n36525 , n36526 );
xor ( n36529 , n35828 , n36426 );
and ( n36530 , n29914 , n36462 );
and ( n36531 , n36529 , n36530 );
xor ( n36532 , n36529 , n36530 );
xor ( n36533 , n35832 , n36424 );
and ( n36534 , n29919 , n36462 );
and ( n36535 , n36533 , n36534 );
xor ( n36536 , n36533 , n36534 );
xor ( n36537 , n35836 , n36422 );
and ( n36538 , n29924 , n36462 );
and ( n36539 , n36537 , n36538 );
xor ( n36540 , n36537 , n36538 );
xor ( n36541 , n35840 , n36420 );
and ( n36542 , n29929 , n36462 );
and ( n36543 , n36541 , n36542 );
xor ( n36544 , n36541 , n36542 );
xor ( n36545 , n35844 , n36418 );
and ( n36546 , n29934 , n36462 );
and ( n36547 , n36545 , n36546 );
xor ( n36548 , n36545 , n36546 );
xor ( n36549 , n35848 , n36416 );
and ( n36550 , n29939 , n36462 );
and ( n36551 , n36549 , n36550 );
xor ( n36552 , n36549 , n36550 );
xor ( n36553 , n35852 , n36414 );
and ( n36554 , n29944 , n36462 );
and ( n36555 , n36553 , n36554 );
xor ( n36556 , n36553 , n36554 );
xor ( n36557 , n35856 , n36412 );
and ( n36558 , n29949 , n36462 );
and ( n36559 , n36557 , n36558 );
xor ( n36560 , n36557 , n36558 );
xor ( n36561 , n35860 , n36410 );
and ( n36562 , n29954 , n36462 );
and ( n36563 , n36561 , n36562 );
xor ( n36564 , n36561 , n36562 );
xor ( n36565 , n35864 , n36408 );
and ( n36566 , n29959 , n36462 );
and ( n36567 , n36565 , n36566 );
xor ( n36568 , n36565 , n36566 );
xor ( n36569 , n35868 , n36406 );
and ( n36570 , n29964 , n36462 );
and ( n36571 , n36569 , n36570 );
xor ( n36572 , n36569 , n36570 );
xor ( n36573 , n35872 , n36404 );
and ( n36574 , n29969 , n36462 );
and ( n36575 , n36573 , n36574 );
xor ( n36576 , n36573 , n36574 );
xor ( n36577 , n35876 , n36402 );
and ( n36578 , n29974 , n36462 );
and ( n36579 , n36577 , n36578 );
xor ( n36580 , n36577 , n36578 );
xor ( n36581 , n35880 , n36400 );
and ( n36582 , n29979 , n36462 );
and ( n36583 , n36581 , n36582 );
xor ( n36584 , n36581 , n36582 );
xor ( n36585 , n35884 , n36398 );
and ( n36586 , n29984 , n36462 );
and ( n36587 , n36585 , n36586 );
xor ( n36588 , n36585 , n36586 );
xor ( n36589 , n35888 , n36396 );
and ( n36590 , n29989 , n36462 );
and ( n36591 , n36589 , n36590 );
xor ( n36592 , n36589 , n36590 );
xor ( n36593 , n35892 , n36394 );
and ( n36594 , n29994 , n36462 );
and ( n36595 , n36593 , n36594 );
xor ( n36596 , n36593 , n36594 );
xor ( n36597 , n35896 , n36392 );
and ( n36598 , n29999 , n36462 );
and ( n36599 , n36597 , n36598 );
xor ( n36600 , n36597 , n36598 );
xor ( n36601 , n35900 , n36390 );
and ( n36602 , n30004 , n36462 );
and ( n36603 , n36601 , n36602 );
xor ( n36604 , n36601 , n36602 );
xor ( n36605 , n35904 , n36388 );
and ( n36606 , n30009 , n36462 );
and ( n36607 , n36605 , n36606 );
xor ( n36608 , n36605 , n36606 );
xor ( n36609 , n35908 , n36386 );
and ( n36610 , n30014 , n36462 );
and ( n36611 , n36609 , n36610 );
xor ( n36612 , n36609 , n36610 );
xor ( n36613 , n35912 , n36384 );
and ( n36614 , n30019 , n36462 );
and ( n36615 , n36613 , n36614 );
xor ( n36616 , n36613 , n36614 );
xor ( n36617 , n35916 , n36382 );
and ( n36618 , n30024 , n36462 );
and ( n36619 , n36617 , n36618 );
xor ( n36620 , n36617 , n36618 );
xor ( n36621 , n35920 , n36380 );
and ( n36622 , n30029 , n36462 );
and ( n36623 , n36621 , n36622 );
xor ( n36624 , n36621 , n36622 );
xor ( n36625 , n35924 , n36378 );
and ( n36626 , n30034 , n36462 );
and ( n36627 , n36625 , n36626 );
xor ( n36628 , n36625 , n36626 );
xor ( n36629 , n35928 , n36376 );
and ( n36630 , n30039 , n36462 );
and ( n36631 , n36629 , n36630 );
xor ( n36632 , n36629 , n36630 );
xor ( n36633 , n35932 , n36374 );
and ( n36634 , n30044 , n36462 );
and ( n36635 , n36633 , n36634 );
xor ( n36636 , n36633 , n36634 );
xor ( n36637 , n35936 , n36372 );
and ( n36638 , n30049 , n36462 );
and ( n36639 , n36637 , n36638 );
xor ( n36640 , n36637 , n36638 );
xor ( n36641 , n35940 , n36370 );
and ( n36642 , n30054 , n36462 );
and ( n36643 , n36641 , n36642 );
xor ( n36644 , n36641 , n36642 );
xor ( n36645 , n35944 , n36368 );
and ( n36646 , n30059 , n36462 );
and ( n36647 , n36645 , n36646 );
xor ( n36648 , n36645 , n36646 );
xor ( n36649 , n35948 , n36366 );
and ( n36650 , n30064 , n36462 );
and ( n36651 , n36649 , n36650 );
xor ( n36652 , n36649 , n36650 );
xor ( n36653 , n35952 , n36364 );
and ( n36654 , n30069 , n36462 );
and ( n36655 , n36653 , n36654 );
xor ( n36656 , n36653 , n36654 );
xor ( n36657 , n35956 , n36362 );
and ( n36658 , n30074 , n36462 );
and ( n36659 , n36657 , n36658 );
xor ( n36660 , n36657 , n36658 );
xor ( n36661 , n35960 , n36360 );
and ( n36662 , n30079 , n36462 );
and ( n36663 , n36661 , n36662 );
xor ( n36664 , n36661 , n36662 );
xor ( n36665 , n35964 , n36358 );
and ( n36666 , n30084 , n36462 );
and ( n36667 , n36665 , n36666 );
xor ( n36668 , n36665 , n36666 );
xor ( n36669 , n35968 , n36356 );
and ( n36670 , n30089 , n36462 );
and ( n36671 , n36669 , n36670 );
xor ( n36672 , n36669 , n36670 );
xor ( n36673 , n35972 , n36354 );
and ( n36674 , n30094 , n36462 );
and ( n36675 , n36673 , n36674 );
xor ( n36676 , n36673 , n36674 );
xor ( n36677 , n35976 , n36352 );
and ( n36678 , n30099 , n36462 );
and ( n36679 , n36677 , n36678 );
xor ( n36680 , n36677 , n36678 );
xor ( n36681 , n35980 , n36350 );
and ( n36682 , n30104 , n36462 );
and ( n36683 , n36681 , n36682 );
xor ( n36684 , n36681 , n36682 );
xor ( n36685 , n35984 , n36348 );
and ( n36686 , n30109 , n36462 );
and ( n36687 , n36685 , n36686 );
xor ( n36688 , n36685 , n36686 );
xor ( n36689 , n35988 , n36346 );
and ( n36690 , n30114 , n36462 );
and ( n36691 , n36689 , n36690 );
xor ( n36692 , n36689 , n36690 );
xor ( n36693 , n35992 , n36344 );
and ( n36694 , n30119 , n36462 );
and ( n36695 , n36693 , n36694 );
xor ( n36696 , n36693 , n36694 );
xor ( n36697 , n35996 , n36342 );
and ( n36698 , n30124 , n36462 );
and ( n36699 , n36697 , n36698 );
xor ( n36700 , n36697 , n36698 );
xor ( n36701 , n36000 , n36340 );
and ( n36702 , n30129 , n36462 );
and ( n36703 , n36701 , n36702 );
xor ( n36704 , n36701 , n36702 );
xor ( n36705 , n36004 , n36338 );
and ( n36706 , n30134 , n36462 );
and ( n36707 , n36705 , n36706 );
xor ( n36708 , n36705 , n36706 );
xor ( n36709 , n36008 , n36336 );
and ( n36710 , n30139 , n36462 );
and ( n36711 , n36709 , n36710 );
xor ( n36712 , n36709 , n36710 );
xor ( n36713 , n36012 , n36334 );
and ( n36714 , n30144 , n36462 );
and ( n36715 , n36713 , n36714 );
xor ( n36716 , n36713 , n36714 );
xor ( n36717 , n36016 , n36332 );
and ( n36718 , n30149 , n36462 );
and ( n36719 , n36717 , n36718 );
xor ( n36720 , n36717 , n36718 );
xor ( n36721 , n36020 , n36330 );
and ( n36722 , n30154 , n36462 );
and ( n36723 , n36721 , n36722 );
xor ( n36724 , n36721 , n36722 );
xor ( n36725 , n36024 , n36328 );
and ( n36726 , n30159 , n36462 );
and ( n36727 , n36725 , n36726 );
xor ( n36728 , n36725 , n36726 );
xor ( n36729 , n36028 , n36326 );
and ( n36730 , n30164 , n36462 );
and ( n36731 , n36729 , n36730 );
xor ( n36732 , n36729 , n36730 );
xor ( n36733 , n36032 , n36324 );
and ( n36734 , n30169 , n36462 );
and ( n36735 , n36733 , n36734 );
xor ( n36736 , n36733 , n36734 );
xor ( n36737 , n36036 , n36322 );
and ( n36738 , n30174 , n36462 );
and ( n36739 , n36737 , n36738 );
xor ( n36740 , n36737 , n36738 );
xor ( n36741 , n36040 , n36320 );
and ( n36742 , n30179 , n36462 );
and ( n36743 , n36741 , n36742 );
xor ( n36744 , n36741 , n36742 );
xor ( n36745 , n36044 , n36318 );
and ( n36746 , n30184 , n36462 );
and ( n36747 , n36745 , n36746 );
xor ( n36748 , n36745 , n36746 );
xor ( n36749 , n36048 , n36316 );
and ( n36750 , n30189 , n36462 );
and ( n36751 , n36749 , n36750 );
xor ( n36752 , n36749 , n36750 );
xor ( n36753 , n36052 , n36314 );
and ( n36754 , n30194 , n36462 );
and ( n36755 , n36753 , n36754 );
xor ( n36756 , n36753 , n36754 );
xor ( n36757 , n36056 , n36312 );
and ( n36758 , n30199 , n36462 );
and ( n36759 , n36757 , n36758 );
xor ( n36760 , n36757 , n36758 );
xor ( n36761 , n36060 , n36310 );
and ( n36762 , n30204 , n36462 );
and ( n36763 , n36761 , n36762 );
xor ( n36764 , n36761 , n36762 );
xor ( n36765 , n36064 , n36308 );
and ( n36766 , n30209 , n36462 );
and ( n36767 , n36765 , n36766 );
xor ( n36768 , n36765 , n36766 );
xor ( n36769 , n36068 , n36306 );
and ( n36770 , n30214 , n36462 );
and ( n36771 , n36769 , n36770 );
xor ( n36772 , n36769 , n36770 );
xor ( n36773 , n36072 , n36304 );
and ( n36774 , n30219 , n36462 );
and ( n36775 , n36773 , n36774 );
xor ( n36776 , n36773 , n36774 );
xor ( n36777 , n36076 , n36302 );
and ( n36778 , n30224 , n36462 );
and ( n36779 , n36777 , n36778 );
xor ( n36780 , n36777 , n36778 );
xor ( n36781 , n36080 , n36300 );
and ( n36782 , n30229 , n36462 );
and ( n36783 , n36781 , n36782 );
xor ( n36784 , n36781 , n36782 );
xor ( n36785 , n36084 , n36298 );
and ( n36786 , n30234 , n36462 );
and ( n36787 , n36785 , n36786 );
xor ( n36788 , n36785 , n36786 );
xor ( n36789 , n36088 , n36296 );
and ( n36790 , n30239 , n36462 );
and ( n36791 , n36789 , n36790 );
xor ( n36792 , n36789 , n36790 );
xor ( n36793 , n36092 , n36294 );
and ( n36794 , n30244 , n36462 );
and ( n36795 , n36793 , n36794 );
xor ( n36796 , n36793 , n36794 );
xor ( n36797 , n36096 , n36292 );
and ( n36798 , n30249 , n36462 );
and ( n36799 , n36797 , n36798 );
xor ( n36800 , n36797 , n36798 );
xor ( n36801 , n36100 , n36290 );
and ( n36802 , n30254 , n36462 );
and ( n36803 , n36801 , n36802 );
xor ( n36804 , n36801 , n36802 );
xor ( n36805 , n36104 , n36288 );
and ( n36806 , n30259 , n36462 );
and ( n36807 , n36805 , n36806 );
xor ( n36808 , n36805 , n36806 );
xor ( n36809 , n36108 , n36286 );
and ( n36810 , n30264 , n36462 );
and ( n36811 , n36809 , n36810 );
xor ( n36812 , n36809 , n36810 );
xor ( n36813 , n36112 , n36284 );
and ( n36814 , n30269 , n36462 );
and ( n36815 , n36813 , n36814 );
xor ( n36816 , n36813 , n36814 );
xor ( n36817 , n36116 , n36282 );
and ( n36818 , n30274 , n36462 );
and ( n36819 , n36817 , n36818 );
xor ( n36820 , n36817 , n36818 );
xor ( n36821 , n36120 , n36280 );
and ( n36822 , n30279 , n36462 );
and ( n36823 , n36821 , n36822 );
xor ( n36824 , n36821 , n36822 );
xor ( n36825 , n36124 , n36278 );
and ( n36826 , n30284 , n36462 );
and ( n36827 , n36825 , n36826 );
xor ( n36828 , n36825 , n36826 );
xor ( n36829 , n36128 , n36276 );
and ( n36830 , n30289 , n36462 );
and ( n36831 , n36829 , n36830 );
xor ( n36832 , n36829 , n36830 );
xor ( n36833 , n36132 , n36274 );
and ( n36834 , n30294 , n36462 );
and ( n36835 , n36833 , n36834 );
xor ( n36836 , n36833 , n36834 );
xor ( n36837 , n36136 , n36272 );
and ( n36838 , n30299 , n36462 );
and ( n36839 , n36837 , n36838 );
xor ( n36840 , n36837 , n36838 );
xor ( n36841 , n36140 , n36270 );
and ( n36842 , n30304 , n36462 );
and ( n36843 , n36841 , n36842 );
xor ( n36844 , n36841 , n36842 );
xor ( n36845 , n36144 , n36268 );
and ( n36846 , n30309 , n36462 );
and ( n36847 , n36845 , n36846 );
xor ( n36848 , n36845 , n36846 );
xor ( n36849 , n36148 , n36266 );
and ( n36850 , n30314 , n36462 );
and ( n36851 , n36849 , n36850 );
xor ( n36852 , n36849 , n36850 );
xor ( n36853 , n36152 , n36264 );
and ( n36854 , n30319 , n36462 );
and ( n36855 , n36853 , n36854 );
xor ( n36856 , n36853 , n36854 );
xor ( n36857 , n36156 , n36262 );
and ( n36858 , n30324 , n36462 );
and ( n36859 , n36857 , n36858 );
xor ( n36860 , n36857 , n36858 );
xor ( n36861 , n36160 , n36260 );
and ( n36862 , n30329 , n36462 );
and ( n36863 , n36861 , n36862 );
xor ( n36864 , n36861 , n36862 );
xor ( n36865 , n36164 , n36258 );
and ( n36866 , n30334 , n36462 );
and ( n36867 , n36865 , n36866 );
xor ( n36868 , n36865 , n36866 );
xor ( n36869 , n36168 , n36256 );
and ( n36870 , n30339 , n36462 );
and ( n36871 , n36869 , n36870 );
xor ( n36872 , n36869 , n36870 );
xor ( n36873 , n36172 , n36254 );
and ( n36874 , n30344 , n36462 );
and ( n36875 , n36873 , n36874 );
xor ( n36876 , n36873 , n36874 );
xor ( n36877 , n36176 , n36252 );
and ( n36878 , n30349 , n36462 );
and ( n36879 , n36877 , n36878 );
xor ( n36880 , n36877 , n36878 );
xor ( n36881 , n36180 , n36250 );
and ( n36882 , n30354 , n36462 );
and ( n36883 , n36881 , n36882 );
xor ( n36884 , n36881 , n36882 );
xor ( n36885 , n36184 , n36248 );
and ( n36886 , n30359 , n36462 );
and ( n36887 , n36885 , n36886 );
xor ( n36888 , n36885 , n36886 );
xor ( n36889 , n36188 , n36246 );
and ( n36890 , n30364 , n36462 );
and ( n36891 , n36889 , n36890 );
xor ( n36892 , n36889 , n36890 );
xor ( n36893 , n36192 , n36244 );
and ( n36894 , n30369 , n36462 );
and ( n36895 , n36893 , n36894 );
xor ( n36896 , n36893 , n36894 );
xor ( n36897 , n36196 , n36242 );
and ( n36898 , n30374 , n36462 );
and ( n36899 , n36897 , n36898 );
xor ( n36900 , n36897 , n36898 );
xor ( n36901 , n36200 , n36240 );
and ( n36902 , n30379 , n36462 );
and ( n36903 , n36901 , n36902 );
xor ( n36904 , n36901 , n36902 );
xor ( n36905 , n36204 , n36238 );
and ( n36906 , n30384 , n36462 );
and ( n36907 , n36905 , n36906 );
xor ( n36908 , n36905 , n36906 );
xor ( n36909 , n36208 , n36236 );
and ( n36910 , n30389 , n36462 );
and ( n36911 , n36909 , n36910 );
xor ( n36912 , n36909 , n36910 );
xor ( n36913 , n36212 , n36234 );
and ( n36914 , n30394 , n36462 );
and ( n36915 , n36913 , n36914 );
xor ( n36916 , n36913 , n36914 );
xor ( n36917 , n36216 , n36232 );
and ( n36918 , n30399 , n36462 );
and ( n36919 , n36917 , n36918 );
xor ( n36920 , n36917 , n36918 );
xor ( n36921 , n36220 , n36230 );
and ( n36922 , n30404 , n36462 );
and ( n36923 , n36921 , n36922 );
xor ( n36924 , n36921 , n36922 );
xor ( n36925 , n36224 , n36228 );
and ( n36926 , n30409 , n36462 );
and ( n36927 , n36925 , n36926 );
buf ( n36928 , n36927 );
and ( n36929 , n36924 , n36928 );
or ( n36930 , n36923 , n36929 );
and ( n36931 , n36920 , n36930 );
or ( n36932 , n36919 , n36931 );
and ( n36933 , n36916 , n36932 );
or ( n36934 , n36915 , n36933 );
and ( n36935 , n36912 , n36934 );
or ( n36936 , n36911 , n36935 );
and ( n36937 , n36908 , n36936 );
or ( n36938 , n36907 , n36937 );
and ( n36939 , n36904 , n36938 );
or ( n36940 , n36903 , n36939 );
and ( n36941 , n36900 , n36940 );
or ( n36942 , n36899 , n36941 );
and ( n36943 , n36896 , n36942 );
or ( n36944 , n36895 , n36943 );
and ( n36945 , n36892 , n36944 );
or ( n36946 , n36891 , n36945 );
and ( n36947 , n36888 , n36946 );
or ( n36948 , n36887 , n36947 );
and ( n36949 , n36884 , n36948 );
or ( n36950 , n36883 , n36949 );
and ( n36951 , n36880 , n36950 );
or ( n36952 , n36879 , n36951 );
and ( n36953 , n36876 , n36952 );
or ( n36954 , n36875 , n36953 );
and ( n36955 , n36872 , n36954 );
or ( n36956 , n36871 , n36955 );
and ( n36957 , n36868 , n36956 );
or ( n36958 , n36867 , n36957 );
and ( n36959 , n36864 , n36958 );
or ( n36960 , n36863 , n36959 );
and ( n36961 , n36860 , n36960 );
or ( n36962 , n36859 , n36961 );
and ( n36963 , n36856 , n36962 );
or ( n36964 , n36855 , n36963 );
and ( n36965 , n36852 , n36964 );
or ( n36966 , n36851 , n36965 );
and ( n36967 , n36848 , n36966 );
or ( n36968 , n36847 , n36967 );
and ( n36969 , n36844 , n36968 );
or ( n36970 , n36843 , n36969 );
and ( n36971 , n36840 , n36970 );
or ( n36972 , n36839 , n36971 );
and ( n36973 , n36836 , n36972 );
or ( n36974 , n36835 , n36973 );
and ( n36975 , n36832 , n36974 );
or ( n36976 , n36831 , n36975 );
and ( n36977 , n36828 , n36976 );
or ( n36978 , n36827 , n36977 );
and ( n36979 , n36824 , n36978 );
or ( n36980 , n36823 , n36979 );
and ( n36981 , n36820 , n36980 );
or ( n36982 , n36819 , n36981 );
and ( n36983 , n36816 , n36982 );
or ( n36984 , n36815 , n36983 );
and ( n36985 , n36812 , n36984 );
or ( n36986 , n36811 , n36985 );
and ( n36987 , n36808 , n36986 );
or ( n36988 , n36807 , n36987 );
and ( n36989 , n36804 , n36988 );
or ( n36990 , n36803 , n36989 );
and ( n36991 , n36800 , n36990 );
or ( n36992 , n36799 , n36991 );
and ( n36993 , n36796 , n36992 );
or ( n36994 , n36795 , n36993 );
and ( n36995 , n36792 , n36994 );
or ( n36996 , n36791 , n36995 );
and ( n36997 , n36788 , n36996 );
or ( n36998 , n36787 , n36997 );
and ( n36999 , n36784 , n36998 );
or ( n37000 , n36783 , n36999 );
and ( n37001 , n36780 , n37000 );
or ( n37002 , n36779 , n37001 );
and ( n37003 , n36776 , n37002 );
or ( n37004 , n36775 , n37003 );
and ( n37005 , n36772 , n37004 );
or ( n37006 , n36771 , n37005 );
and ( n37007 , n36768 , n37006 );
or ( n37008 , n36767 , n37007 );
and ( n37009 , n36764 , n37008 );
or ( n37010 , n36763 , n37009 );
and ( n37011 , n36760 , n37010 );
or ( n37012 , n36759 , n37011 );
and ( n37013 , n36756 , n37012 );
or ( n37014 , n36755 , n37013 );
and ( n37015 , n36752 , n37014 );
or ( n37016 , n36751 , n37015 );
and ( n37017 , n36748 , n37016 );
or ( n37018 , n36747 , n37017 );
and ( n37019 , n36744 , n37018 );
or ( n37020 , n36743 , n37019 );
and ( n37021 , n36740 , n37020 );
or ( n37022 , n36739 , n37021 );
and ( n37023 , n36736 , n37022 );
or ( n37024 , n36735 , n37023 );
and ( n37025 , n36732 , n37024 );
or ( n37026 , n36731 , n37025 );
and ( n37027 , n36728 , n37026 );
or ( n37028 , n36727 , n37027 );
and ( n37029 , n36724 , n37028 );
or ( n37030 , n36723 , n37029 );
and ( n37031 , n36720 , n37030 );
or ( n37032 , n36719 , n37031 );
and ( n37033 , n36716 , n37032 );
or ( n37034 , n36715 , n37033 );
and ( n37035 , n36712 , n37034 );
or ( n37036 , n36711 , n37035 );
and ( n37037 , n36708 , n37036 );
or ( n37038 , n36707 , n37037 );
and ( n37039 , n36704 , n37038 );
or ( n37040 , n36703 , n37039 );
and ( n37041 , n36700 , n37040 );
or ( n37042 , n36699 , n37041 );
and ( n37043 , n36696 , n37042 );
or ( n37044 , n36695 , n37043 );
and ( n37045 , n36692 , n37044 );
or ( n37046 , n36691 , n37045 );
and ( n37047 , n36688 , n37046 );
or ( n37048 , n36687 , n37047 );
and ( n37049 , n36684 , n37048 );
or ( n37050 , n36683 , n37049 );
and ( n37051 , n36680 , n37050 );
or ( n37052 , n36679 , n37051 );
and ( n37053 , n36676 , n37052 );
or ( n37054 , n36675 , n37053 );
and ( n37055 , n36672 , n37054 );
or ( n37056 , n36671 , n37055 );
and ( n37057 , n36668 , n37056 );
or ( n37058 , n36667 , n37057 );
and ( n37059 , n36664 , n37058 );
or ( n37060 , n36663 , n37059 );
and ( n37061 , n36660 , n37060 );
or ( n37062 , n36659 , n37061 );
and ( n37063 , n36656 , n37062 );
or ( n37064 , n36655 , n37063 );
and ( n37065 , n36652 , n37064 );
or ( n37066 , n36651 , n37065 );
and ( n37067 , n36648 , n37066 );
or ( n37068 , n36647 , n37067 );
and ( n37069 , n36644 , n37068 );
or ( n37070 , n36643 , n37069 );
and ( n37071 , n36640 , n37070 );
or ( n37072 , n36639 , n37071 );
and ( n37073 , n36636 , n37072 );
or ( n37074 , n36635 , n37073 );
and ( n37075 , n36632 , n37074 );
or ( n37076 , n36631 , n37075 );
and ( n37077 , n36628 , n37076 );
or ( n37078 , n36627 , n37077 );
and ( n37079 , n36624 , n37078 );
or ( n37080 , n36623 , n37079 );
and ( n37081 , n36620 , n37080 );
or ( n37082 , n36619 , n37081 );
and ( n37083 , n36616 , n37082 );
or ( n37084 , n36615 , n37083 );
and ( n37085 , n36612 , n37084 );
or ( n37086 , n36611 , n37085 );
and ( n37087 , n36608 , n37086 );
or ( n37088 , n36607 , n37087 );
and ( n37089 , n36604 , n37088 );
or ( n37090 , n36603 , n37089 );
and ( n37091 , n36600 , n37090 );
or ( n37092 , n36599 , n37091 );
and ( n37093 , n36596 , n37092 );
or ( n37094 , n36595 , n37093 );
and ( n37095 , n36592 , n37094 );
or ( n37096 , n36591 , n37095 );
and ( n37097 , n36588 , n37096 );
or ( n37098 , n36587 , n37097 );
and ( n37099 , n36584 , n37098 );
or ( n37100 , n36583 , n37099 );
and ( n37101 , n36580 , n37100 );
or ( n37102 , n36579 , n37101 );
and ( n37103 , n36576 , n37102 );
or ( n37104 , n36575 , n37103 );
and ( n37105 , n36572 , n37104 );
or ( n37106 , n36571 , n37105 );
and ( n37107 , n36568 , n37106 );
or ( n37108 , n36567 , n37107 );
and ( n37109 , n36564 , n37108 );
or ( n37110 , n36563 , n37109 );
and ( n37111 , n36560 , n37110 );
or ( n37112 , n36559 , n37111 );
and ( n37113 , n36556 , n37112 );
or ( n37114 , n36555 , n37113 );
and ( n37115 , n36552 , n37114 );
or ( n37116 , n36551 , n37115 );
and ( n37117 , n36548 , n37116 );
or ( n37118 , n36547 , n37117 );
and ( n37119 , n36544 , n37118 );
or ( n37120 , n36543 , n37119 );
and ( n37121 , n36540 , n37120 );
or ( n37122 , n36539 , n37121 );
and ( n37123 , n36536 , n37122 );
or ( n37124 , n36535 , n37123 );
and ( n37125 , n36532 , n37124 );
or ( n37126 , n36531 , n37125 );
and ( n37127 , n36528 , n37126 );
or ( n37128 , n36527 , n37127 );
and ( n37129 , n36524 , n37128 );
or ( n37130 , n36523 , n37129 );
and ( n37131 , n36520 , n37130 );
or ( n37132 , n36519 , n37131 );
and ( n37133 , n36516 , n37132 );
or ( n37134 , n36515 , n37133 );
and ( n37135 , n36512 , n37134 );
or ( n37136 , n36511 , n37135 );
and ( n37137 , n36508 , n37136 );
or ( n37138 , n36507 , n37137 );
and ( n37139 , n36504 , n37138 );
or ( n37140 , n36503 , n37139 );
and ( n37141 , n36500 , n37140 );
or ( n37142 , n36499 , n37141 );
and ( n37143 , n36496 , n37142 );
or ( n37144 , n36495 , n37143 );
and ( n37145 , n36492 , n37144 );
or ( n37146 , n36491 , n37145 );
and ( n37147 , n36488 , n37146 );
or ( n37148 , n36487 , n37147 );
and ( n37149 , n36484 , n37148 );
or ( n37150 , n36483 , n37149 );
and ( n37151 , n36480 , n37150 );
or ( n37152 , n36479 , n37151 );
and ( n37153 , n36476 , n37152 );
or ( n37154 , n36475 , n37153 );
and ( n37155 , n36472 , n37154 );
or ( n37156 , n36471 , n37155 );
and ( n37157 , n36468 , n37156 );
or ( n37158 , n36467 , n37157 );
xor ( n37159 , n36464 , n37158 );
buf ( n37160 , n18084 );
and ( n37161 , n29834 , n37160 );
xor ( n37162 , n37159 , n37161 );
xor ( n37163 , n36468 , n37156 );
and ( n37164 , n29839 , n37160 );
and ( n37165 , n37163 , n37164 );
xor ( n37166 , n37163 , n37164 );
xor ( n37167 , n36472 , n37154 );
and ( n37168 , n29844 , n37160 );
and ( n37169 , n37167 , n37168 );
xor ( n37170 , n37167 , n37168 );
xor ( n37171 , n36476 , n37152 );
and ( n37172 , n29849 , n37160 );
and ( n37173 , n37171 , n37172 );
xor ( n37174 , n37171 , n37172 );
xor ( n37175 , n36480 , n37150 );
and ( n37176 , n29854 , n37160 );
and ( n37177 , n37175 , n37176 );
xor ( n37178 , n37175 , n37176 );
xor ( n37179 , n36484 , n37148 );
and ( n37180 , n29859 , n37160 );
and ( n37181 , n37179 , n37180 );
xor ( n37182 , n37179 , n37180 );
xor ( n37183 , n36488 , n37146 );
and ( n37184 , n29864 , n37160 );
and ( n37185 , n37183 , n37184 );
xor ( n37186 , n37183 , n37184 );
xor ( n37187 , n36492 , n37144 );
and ( n37188 , n29869 , n37160 );
and ( n37189 , n37187 , n37188 );
xor ( n37190 , n37187 , n37188 );
xor ( n37191 , n36496 , n37142 );
and ( n37192 , n29874 , n37160 );
and ( n37193 , n37191 , n37192 );
xor ( n37194 , n37191 , n37192 );
xor ( n37195 , n36500 , n37140 );
and ( n37196 , n29879 , n37160 );
and ( n37197 , n37195 , n37196 );
xor ( n37198 , n37195 , n37196 );
xor ( n37199 , n36504 , n37138 );
and ( n37200 , n29884 , n37160 );
and ( n37201 , n37199 , n37200 );
xor ( n37202 , n37199 , n37200 );
xor ( n37203 , n36508 , n37136 );
and ( n37204 , n29889 , n37160 );
and ( n37205 , n37203 , n37204 );
xor ( n37206 , n37203 , n37204 );
xor ( n37207 , n36512 , n37134 );
and ( n37208 , n29894 , n37160 );
and ( n37209 , n37207 , n37208 );
xor ( n37210 , n37207 , n37208 );
xor ( n37211 , n36516 , n37132 );
and ( n37212 , n29899 , n37160 );
and ( n37213 , n37211 , n37212 );
xor ( n37214 , n37211 , n37212 );
xor ( n37215 , n36520 , n37130 );
and ( n37216 , n29904 , n37160 );
and ( n37217 , n37215 , n37216 );
xor ( n37218 , n37215 , n37216 );
xor ( n37219 , n36524 , n37128 );
and ( n37220 , n29909 , n37160 );
and ( n37221 , n37219 , n37220 );
xor ( n37222 , n37219 , n37220 );
xor ( n37223 , n36528 , n37126 );
and ( n37224 , n29914 , n37160 );
and ( n37225 , n37223 , n37224 );
xor ( n37226 , n37223 , n37224 );
xor ( n37227 , n36532 , n37124 );
and ( n37228 , n29919 , n37160 );
and ( n37229 , n37227 , n37228 );
xor ( n37230 , n37227 , n37228 );
xor ( n37231 , n36536 , n37122 );
and ( n37232 , n29924 , n37160 );
and ( n37233 , n37231 , n37232 );
xor ( n37234 , n37231 , n37232 );
xor ( n37235 , n36540 , n37120 );
and ( n37236 , n29929 , n37160 );
and ( n37237 , n37235 , n37236 );
xor ( n37238 , n37235 , n37236 );
xor ( n37239 , n36544 , n37118 );
and ( n37240 , n29934 , n37160 );
and ( n37241 , n37239 , n37240 );
xor ( n37242 , n37239 , n37240 );
xor ( n37243 , n36548 , n37116 );
and ( n37244 , n29939 , n37160 );
and ( n37245 , n37243 , n37244 );
xor ( n37246 , n37243 , n37244 );
xor ( n37247 , n36552 , n37114 );
and ( n37248 , n29944 , n37160 );
and ( n37249 , n37247 , n37248 );
xor ( n37250 , n37247 , n37248 );
xor ( n37251 , n36556 , n37112 );
and ( n37252 , n29949 , n37160 );
and ( n37253 , n37251 , n37252 );
xor ( n37254 , n37251 , n37252 );
xor ( n37255 , n36560 , n37110 );
and ( n37256 , n29954 , n37160 );
and ( n37257 , n37255 , n37256 );
xor ( n37258 , n37255 , n37256 );
xor ( n37259 , n36564 , n37108 );
and ( n37260 , n29959 , n37160 );
and ( n37261 , n37259 , n37260 );
xor ( n37262 , n37259 , n37260 );
xor ( n37263 , n36568 , n37106 );
and ( n37264 , n29964 , n37160 );
and ( n37265 , n37263 , n37264 );
xor ( n37266 , n37263 , n37264 );
xor ( n37267 , n36572 , n37104 );
and ( n37268 , n29969 , n37160 );
and ( n37269 , n37267 , n37268 );
xor ( n37270 , n37267 , n37268 );
xor ( n37271 , n36576 , n37102 );
and ( n37272 , n29974 , n37160 );
and ( n37273 , n37271 , n37272 );
xor ( n37274 , n37271 , n37272 );
xor ( n37275 , n36580 , n37100 );
and ( n37276 , n29979 , n37160 );
and ( n37277 , n37275 , n37276 );
xor ( n37278 , n37275 , n37276 );
xor ( n37279 , n36584 , n37098 );
and ( n37280 , n29984 , n37160 );
and ( n37281 , n37279 , n37280 );
xor ( n37282 , n37279 , n37280 );
xor ( n37283 , n36588 , n37096 );
and ( n37284 , n29989 , n37160 );
and ( n37285 , n37283 , n37284 );
xor ( n37286 , n37283 , n37284 );
xor ( n37287 , n36592 , n37094 );
and ( n37288 , n29994 , n37160 );
and ( n37289 , n37287 , n37288 );
xor ( n37290 , n37287 , n37288 );
xor ( n37291 , n36596 , n37092 );
and ( n37292 , n29999 , n37160 );
and ( n37293 , n37291 , n37292 );
xor ( n37294 , n37291 , n37292 );
xor ( n37295 , n36600 , n37090 );
and ( n37296 , n30004 , n37160 );
and ( n37297 , n37295 , n37296 );
xor ( n37298 , n37295 , n37296 );
xor ( n37299 , n36604 , n37088 );
and ( n37300 , n30009 , n37160 );
and ( n37301 , n37299 , n37300 );
xor ( n37302 , n37299 , n37300 );
xor ( n37303 , n36608 , n37086 );
and ( n37304 , n30014 , n37160 );
and ( n37305 , n37303 , n37304 );
xor ( n37306 , n37303 , n37304 );
xor ( n37307 , n36612 , n37084 );
and ( n37308 , n30019 , n37160 );
and ( n37309 , n37307 , n37308 );
xor ( n37310 , n37307 , n37308 );
xor ( n37311 , n36616 , n37082 );
and ( n37312 , n30024 , n37160 );
and ( n37313 , n37311 , n37312 );
xor ( n37314 , n37311 , n37312 );
xor ( n37315 , n36620 , n37080 );
and ( n37316 , n30029 , n37160 );
and ( n37317 , n37315 , n37316 );
xor ( n37318 , n37315 , n37316 );
xor ( n37319 , n36624 , n37078 );
and ( n37320 , n30034 , n37160 );
and ( n37321 , n37319 , n37320 );
xor ( n37322 , n37319 , n37320 );
xor ( n37323 , n36628 , n37076 );
and ( n37324 , n30039 , n37160 );
and ( n37325 , n37323 , n37324 );
xor ( n37326 , n37323 , n37324 );
xor ( n37327 , n36632 , n37074 );
and ( n37328 , n30044 , n37160 );
and ( n37329 , n37327 , n37328 );
xor ( n37330 , n37327 , n37328 );
xor ( n37331 , n36636 , n37072 );
and ( n37332 , n30049 , n37160 );
and ( n37333 , n37331 , n37332 );
xor ( n37334 , n37331 , n37332 );
xor ( n37335 , n36640 , n37070 );
and ( n37336 , n30054 , n37160 );
and ( n37337 , n37335 , n37336 );
xor ( n37338 , n37335 , n37336 );
xor ( n37339 , n36644 , n37068 );
and ( n37340 , n30059 , n37160 );
and ( n37341 , n37339 , n37340 );
xor ( n37342 , n37339 , n37340 );
xor ( n37343 , n36648 , n37066 );
and ( n37344 , n30064 , n37160 );
and ( n37345 , n37343 , n37344 );
xor ( n37346 , n37343 , n37344 );
xor ( n37347 , n36652 , n37064 );
and ( n37348 , n30069 , n37160 );
and ( n37349 , n37347 , n37348 );
xor ( n37350 , n37347 , n37348 );
xor ( n37351 , n36656 , n37062 );
and ( n37352 , n30074 , n37160 );
and ( n37353 , n37351 , n37352 );
xor ( n37354 , n37351 , n37352 );
xor ( n37355 , n36660 , n37060 );
and ( n37356 , n30079 , n37160 );
and ( n37357 , n37355 , n37356 );
xor ( n37358 , n37355 , n37356 );
xor ( n37359 , n36664 , n37058 );
and ( n37360 , n30084 , n37160 );
and ( n37361 , n37359 , n37360 );
xor ( n37362 , n37359 , n37360 );
xor ( n37363 , n36668 , n37056 );
and ( n37364 , n30089 , n37160 );
and ( n37365 , n37363 , n37364 );
xor ( n37366 , n37363 , n37364 );
xor ( n37367 , n36672 , n37054 );
and ( n37368 , n30094 , n37160 );
and ( n37369 , n37367 , n37368 );
xor ( n37370 , n37367 , n37368 );
xor ( n37371 , n36676 , n37052 );
and ( n37372 , n30099 , n37160 );
and ( n37373 , n37371 , n37372 );
xor ( n37374 , n37371 , n37372 );
xor ( n37375 , n36680 , n37050 );
and ( n37376 , n30104 , n37160 );
and ( n37377 , n37375 , n37376 );
xor ( n37378 , n37375 , n37376 );
xor ( n37379 , n36684 , n37048 );
and ( n37380 , n30109 , n37160 );
and ( n37381 , n37379 , n37380 );
xor ( n37382 , n37379 , n37380 );
xor ( n37383 , n36688 , n37046 );
and ( n37384 , n30114 , n37160 );
and ( n37385 , n37383 , n37384 );
xor ( n37386 , n37383 , n37384 );
xor ( n37387 , n36692 , n37044 );
and ( n37388 , n30119 , n37160 );
and ( n37389 , n37387 , n37388 );
xor ( n37390 , n37387 , n37388 );
xor ( n37391 , n36696 , n37042 );
and ( n37392 , n30124 , n37160 );
and ( n37393 , n37391 , n37392 );
xor ( n37394 , n37391 , n37392 );
xor ( n37395 , n36700 , n37040 );
and ( n37396 , n30129 , n37160 );
and ( n37397 , n37395 , n37396 );
xor ( n37398 , n37395 , n37396 );
xor ( n37399 , n36704 , n37038 );
and ( n37400 , n30134 , n37160 );
and ( n37401 , n37399 , n37400 );
xor ( n37402 , n37399 , n37400 );
xor ( n37403 , n36708 , n37036 );
and ( n37404 , n30139 , n37160 );
and ( n37405 , n37403 , n37404 );
xor ( n37406 , n37403 , n37404 );
xor ( n37407 , n36712 , n37034 );
and ( n37408 , n30144 , n37160 );
and ( n37409 , n37407 , n37408 );
xor ( n37410 , n37407 , n37408 );
xor ( n37411 , n36716 , n37032 );
and ( n37412 , n30149 , n37160 );
and ( n37413 , n37411 , n37412 );
xor ( n37414 , n37411 , n37412 );
xor ( n37415 , n36720 , n37030 );
and ( n37416 , n30154 , n37160 );
and ( n37417 , n37415 , n37416 );
xor ( n37418 , n37415 , n37416 );
xor ( n37419 , n36724 , n37028 );
and ( n37420 , n30159 , n37160 );
and ( n37421 , n37419 , n37420 );
xor ( n37422 , n37419 , n37420 );
xor ( n37423 , n36728 , n37026 );
and ( n37424 , n30164 , n37160 );
and ( n37425 , n37423 , n37424 );
xor ( n37426 , n37423 , n37424 );
xor ( n37427 , n36732 , n37024 );
and ( n37428 , n30169 , n37160 );
and ( n37429 , n37427 , n37428 );
xor ( n37430 , n37427 , n37428 );
xor ( n37431 , n36736 , n37022 );
and ( n37432 , n30174 , n37160 );
and ( n37433 , n37431 , n37432 );
xor ( n37434 , n37431 , n37432 );
xor ( n37435 , n36740 , n37020 );
and ( n37436 , n30179 , n37160 );
and ( n37437 , n37435 , n37436 );
xor ( n37438 , n37435 , n37436 );
xor ( n37439 , n36744 , n37018 );
and ( n37440 , n30184 , n37160 );
and ( n37441 , n37439 , n37440 );
xor ( n37442 , n37439 , n37440 );
xor ( n37443 , n36748 , n37016 );
and ( n37444 , n30189 , n37160 );
and ( n37445 , n37443 , n37444 );
xor ( n37446 , n37443 , n37444 );
xor ( n37447 , n36752 , n37014 );
and ( n37448 , n30194 , n37160 );
and ( n37449 , n37447 , n37448 );
xor ( n37450 , n37447 , n37448 );
xor ( n37451 , n36756 , n37012 );
and ( n37452 , n30199 , n37160 );
and ( n37453 , n37451 , n37452 );
xor ( n37454 , n37451 , n37452 );
xor ( n37455 , n36760 , n37010 );
and ( n37456 , n30204 , n37160 );
and ( n37457 , n37455 , n37456 );
xor ( n37458 , n37455 , n37456 );
xor ( n37459 , n36764 , n37008 );
and ( n37460 , n30209 , n37160 );
and ( n37461 , n37459 , n37460 );
xor ( n37462 , n37459 , n37460 );
xor ( n37463 , n36768 , n37006 );
and ( n37464 , n30214 , n37160 );
and ( n37465 , n37463 , n37464 );
xor ( n37466 , n37463 , n37464 );
xor ( n37467 , n36772 , n37004 );
and ( n37468 , n30219 , n37160 );
and ( n37469 , n37467 , n37468 );
xor ( n37470 , n37467 , n37468 );
xor ( n37471 , n36776 , n37002 );
and ( n37472 , n30224 , n37160 );
and ( n37473 , n37471 , n37472 );
xor ( n37474 , n37471 , n37472 );
xor ( n37475 , n36780 , n37000 );
and ( n37476 , n30229 , n37160 );
and ( n37477 , n37475 , n37476 );
xor ( n37478 , n37475 , n37476 );
xor ( n37479 , n36784 , n36998 );
and ( n37480 , n30234 , n37160 );
and ( n37481 , n37479 , n37480 );
xor ( n37482 , n37479 , n37480 );
xor ( n37483 , n36788 , n36996 );
and ( n37484 , n30239 , n37160 );
and ( n37485 , n37483 , n37484 );
xor ( n37486 , n37483 , n37484 );
xor ( n37487 , n36792 , n36994 );
and ( n37488 , n30244 , n37160 );
and ( n37489 , n37487 , n37488 );
xor ( n37490 , n37487 , n37488 );
xor ( n37491 , n36796 , n36992 );
and ( n37492 , n30249 , n37160 );
and ( n37493 , n37491 , n37492 );
xor ( n37494 , n37491 , n37492 );
xor ( n37495 , n36800 , n36990 );
and ( n37496 , n30254 , n37160 );
and ( n37497 , n37495 , n37496 );
xor ( n37498 , n37495 , n37496 );
xor ( n37499 , n36804 , n36988 );
and ( n37500 , n30259 , n37160 );
and ( n37501 , n37499 , n37500 );
xor ( n37502 , n37499 , n37500 );
xor ( n37503 , n36808 , n36986 );
and ( n37504 , n30264 , n37160 );
and ( n37505 , n37503 , n37504 );
xor ( n37506 , n37503 , n37504 );
xor ( n37507 , n36812 , n36984 );
and ( n37508 , n30269 , n37160 );
and ( n37509 , n37507 , n37508 );
xor ( n37510 , n37507 , n37508 );
xor ( n37511 , n36816 , n36982 );
and ( n37512 , n30274 , n37160 );
and ( n37513 , n37511 , n37512 );
xor ( n37514 , n37511 , n37512 );
xor ( n37515 , n36820 , n36980 );
and ( n37516 , n30279 , n37160 );
and ( n37517 , n37515 , n37516 );
xor ( n37518 , n37515 , n37516 );
xor ( n37519 , n36824 , n36978 );
and ( n37520 , n30284 , n37160 );
and ( n37521 , n37519 , n37520 );
xor ( n37522 , n37519 , n37520 );
xor ( n37523 , n36828 , n36976 );
and ( n37524 , n30289 , n37160 );
and ( n37525 , n37523 , n37524 );
xor ( n37526 , n37523 , n37524 );
xor ( n37527 , n36832 , n36974 );
and ( n37528 , n30294 , n37160 );
and ( n37529 , n37527 , n37528 );
xor ( n37530 , n37527 , n37528 );
xor ( n37531 , n36836 , n36972 );
and ( n37532 , n30299 , n37160 );
and ( n37533 , n37531 , n37532 );
xor ( n37534 , n37531 , n37532 );
xor ( n37535 , n36840 , n36970 );
and ( n37536 , n30304 , n37160 );
and ( n37537 , n37535 , n37536 );
xor ( n37538 , n37535 , n37536 );
xor ( n37539 , n36844 , n36968 );
and ( n37540 , n30309 , n37160 );
and ( n37541 , n37539 , n37540 );
xor ( n37542 , n37539 , n37540 );
xor ( n37543 , n36848 , n36966 );
and ( n37544 , n30314 , n37160 );
and ( n37545 , n37543 , n37544 );
xor ( n37546 , n37543 , n37544 );
xor ( n37547 , n36852 , n36964 );
and ( n37548 , n30319 , n37160 );
and ( n37549 , n37547 , n37548 );
xor ( n37550 , n37547 , n37548 );
xor ( n37551 , n36856 , n36962 );
and ( n37552 , n30324 , n37160 );
and ( n37553 , n37551 , n37552 );
xor ( n37554 , n37551 , n37552 );
xor ( n37555 , n36860 , n36960 );
and ( n37556 , n30329 , n37160 );
and ( n37557 , n37555 , n37556 );
xor ( n37558 , n37555 , n37556 );
xor ( n37559 , n36864 , n36958 );
and ( n37560 , n30334 , n37160 );
and ( n37561 , n37559 , n37560 );
xor ( n37562 , n37559 , n37560 );
xor ( n37563 , n36868 , n36956 );
and ( n37564 , n30339 , n37160 );
and ( n37565 , n37563 , n37564 );
xor ( n37566 , n37563 , n37564 );
xor ( n37567 , n36872 , n36954 );
and ( n37568 , n30344 , n37160 );
and ( n37569 , n37567 , n37568 );
xor ( n37570 , n37567 , n37568 );
xor ( n37571 , n36876 , n36952 );
and ( n37572 , n30349 , n37160 );
and ( n37573 , n37571 , n37572 );
xor ( n37574 , n37571 , n37572 );
xor ( n37575 , n36880 , n36950 );
and ( n37576 , n30354 , n37160 );
and ( n37577 , n37575 , n37576 );
xor ( n37578 , n37575 , n37576 );
xor ( n37579 , n36884 , n36948 );
and ( n37580 , n30359 , n37160 );
and ( n37581 , n37579 , n37580 );
xor ( n37582 , n37579 , n37580 );
xor ( n37583 , n36888 , n36946 );
and ( n37584 , n30364 , n37160 );
and ( n37585 , n37583 , n37584 );
xor ( n37586 , n37583 , n37584 );
xor ( n37587 , n36892 , n36944 );
and ( n37588 , n30369 , n37160 );
and ( n37589 , n37587 , n37588 );
xor ( n37590 , n37587 , n37588 );
xor ( n37591 , n36896 , n36942 );
and ( n37592 , n30374 , n37160 );
and ( n37593 , n37591 , n37592 );
xor ( n37594 , n37591 , n37592 );
xor ( n37595 , n36900 , n36940 );
and ( n37596 , n30379 , n37160 );
and ( n37597 , n37595 , n37596 );
xor ( n37598 , n37595 , n37596 );
xor ( n37599 , n36904 , n36938 );
and ( n37600 , n30384 , n37160 );
and ( n37601 , n37599 , n37600 );
xor ( n37602 , n37599 , n37600 );
xor ( n37603 , n36908 , n36936 );
and ( n37604 , n30389 , n37160 );
and ( n37605 , n37603 , n37604 );
xor ( n37606 , n37603 , n37604 );
xor ( n37607 , n36912 , n36934 );
and ( n37608 , n30394 , n37160 );
and ( n37609 , n37607 , n37608 );
xor ( n37610 , n37607 , n37608 );
xor ( n37611 , n36916 , n36932 );
and ( n37612 , n30399 , n37160 );
and ( n37613 , n37611 , n37612 );
xor ( n37614 , n37611 , n37612 );
xor ( n37615 , n36920 , n36930 );
and ( n37616 , n30404 , n37160 );
and ( n37617 , n37615 , n37616 );
xor ( n37618 , n37615 , n37616 );
xor ( n37619 , n36924 , n36928 );
and ( n37620 , n30409 , n37160 );
and ( n37621 , n37619 , n37620 );
buf ( n37622 , n37621 );
and ( n37623 , n37618 , n37622 );
or ( n37624 , n37617 , n37623 );
and ( n37625 , n37614 , n37624 );
or ( n37626 , n37613 , n37625 );
and ( n37627 , n37610 , n37626 );
or ( n37628 , n37609 , n37627 );
and ( n37629 , n37606 , n37628 );
or ( n37630 , n37605 , n37629 );
and ( n37631 , n37602 , n37630 );
or ( n37632 , n37601 , n37631 );
and ( n37633 , n37598 , n37632 );
or ( n37634 , n37597 , n37633 );
and ( n37635 , n37594 , n37634 );
or ( n37636 , n37593 , n37635 );
and ( n37637 , n37590 , n37636 );
or ( n37638 , n37589 , n37637 );
and ( n37639 , n37586 , n37638 );
or ( n37640 , n37585 , n37639 );
and ( n37641 , n37582 , n37640 );
or ( n37642 , n37581 , n37641 );
and ( n37643 , n37578 , n37642 );
or ( n37644 , n37577 , n37643 );
and ( n37645 , n37574 , n37644 );
or ( n37646 , n37573 , n37645 );
and ( n37647 , n37570 , n37646 );
or ( n37648 , n37569 , n37647 );
and ( n37649 , n37566 , n37648 );
or ( n37650 , n37565 , n37649 );
and ( n37651 , n37562 , n37650 );
or ( n37652 , n37561 , n37651 );
and ( n37653 , n37558 , n37652 );
or ( n37654 , n37557 , n37653 );
and ( n37655 , n37554 , n37654 );
or ( n37656 , n37553 , n37655 );
and ( n37657 , n37550 , n37656 );
or ( n37658 , n37549 , n37657 );
and ( n37659 , n37546 , n37658 );
or ( n37660 , n37545 , n37659 );
and ( n37661 , n37542 , n37660 );
or ( n37662 , n37541 , n37661 );
and ( n37663 , n37538 , n37662 );
or ( n37664 , n37537 , n37663 );
and ( n37665 , n37534 , n37664 );
or ( n37666 , n37533 , n37665 );
and ( n37667 , n37530 , n37666 );
or ( n37668 , n37529 , n37667 );
and ( n37669 , n37526 , n37668 );
or ( n37670 , n37525 , n37669 );
and ( n37671 , n37522 , n37670 );
or ( n37672 , n37521 , n37671 );
and ( n37673 , n37518 , n37672 );
or ( n37674 , n37517 , n37673 );
and ( n37675 , n37514 , n37674 );
or ( n37676 , n37513 , n37675 );
and ( n37677 , n37510 , n37676 );
or ( n37678 , n37509 , n37677 );
and ( n37679 , n37506 , n37678 );
or ( n37680 , n37505 , n37679 );
and ( n37681 , n37502 , n37680 );
or ( n37682 , n37501 , n37681 );
and ( n37683 , n37498 , n37682 );
or ( n37684 , n37497 , n37683 );
and ( n37685 , n37494 , n37684 );
or ( n37686 , n37493 , n37685 );
and ( n37687 , n37490 , n37686 );
or ( n37688 , n37489 , n37687 );
and ( n37689 , n37486 , n37688 );
or ( n37690 , n37485 , n37689 );
and ( n37691 , n37482 , n37690 );
or ( n37692 , n37481 , n37691 );
and ( n37693 , n37478 , n37692 );
or ( n37694 , n37477 , n37693 );
and ( n37695 , n37474 , n37694 );
or ( n37696 , n37473 , n37695 );
and ( n37697 , n37470 , n37696 );
or ( n37698 , n37469 , n37697 );
and ( n37699 , n37466 , n37698 );
or ( n37700 , n37465 , n37699 );
and ( n37701 , n37462 , n37700 );
or ( n37702 , n37461 , n37701 );
and ( n37703 , n37458 , n37702 );
or ( n37704 , n37457 , n37703 );
and ( n37705 , n37454 , n37704 );
or ( n37706 , n37453 , n37705 );
and ( n37707 , n37450 , n37706 );
or ( n37708 , n37449 , n37707 );
and ( n37709 , n37446 , n37708 );
or ( n37710 , n37445 , n37709 );
and ( n37711 , n37442 , n37710 );
or ( n37712 , n37441 , n37711 );
and ( n37713 , n37438 , n37712 );
or ( n37714 , n37437 , n37713 );
and ( n37715 , n37434 , n37714 );
or ( n37716 , n37433 , n37715 );
and ( n37717 , n37430 , n37716 );
or ( n37718 , n37429 , n37717 );
and ( n37719 , n37426 , n37718 );
or ( n37720 , n37425 , n37719 );
and ( n37721 , n37422 , n37720 );
or ( n37722 , n37421 , n37721 );
and ( n37723 , n37418 , n37722 );
or ( n37724 , n37417 , n37723 );
and ( n37725 , n37414 , n37724 );
or ( n37726 , n37413 , n37725 );
and ( n37727 , n37410 , n37726 );
or ( n37728 , n37409 , n37727 );
and ( n37729 , n37406 , n37728 );
or ( n37730 , n37405 , n37729 );
and ( n37731 , n37402 , n37730 );
or ( n37732 , n37401 , n37731 );
and ( n37733 , n37398 , n37732 );
or ( n37734 , n37397 , n37733 );
and ( n37735 , n37394 , n37734 );
or ( n37736 , n37393 , n37735 );
and ( n37737 , n37390 , n37736 );
or ( n37738 , n37389 , n37737 );
and ( n37739 , n37386 , n37738 );
or ( n37740 , n37385 , n37739 );
and ( n37741 , n37382 , n37740 );
or ( n37742 , n37381 , n37741 );
and ( n37743 , n37378 , n37742 );
or ( n37744 , n37377 , n37743 );
and ( n37745 , n37374 , n37744 );
or ( n37746 , n37373 , n37745 );
and ( n37747 , n37370 , n37746 );
or ( n37748 , n37369 , n37747 );
and ( n37749 , n37366 , n37748 );
or ( n37750 , n37365 , n37749 );
and ( n37751 , n37362 , n37750 );
or ( n37752 , n37361 , n37751 );
and ( n37753 , n37358 , n37752 );
or ( n37754 , n37357 , n37753 );
and ( n37755 , n37354 , n37754 );
or ( n37756 , n37353 , n37755 );
and ( n37757 , n37350 , n37756 );
or ( n37758 , n37349 , n37757 );
and ( n37759 , n37346 , n37758 );
or ( n37760 , n37345 , n37759 );
and ( n37761 , n37342 , n37760 );
or ( n37762 , n37341 , n37761 );
and ( n37763 , n37338 , n37762 );
or ( n37764 , n37337 , n37763 );
and ( n37765 , n37334 , n37764 );
or ( n37766 , n37333 , n37765 );
and ( n37767 , n37330 , n37766 );
or ( n37768 , n37329 , n37767 );
and ( n37769 , n37326 , n37768 );
or ( n37770 , n37325 , n37769 );
and ( n37771 , n37322 , n37770 );
or ( n37772 , n37321 , n37771 );
and ( n37773 , n37318 , n37772 );
or ( n37774 , n37317 , n37773 );
and ( n37775 , n37314 , n37774 );
or ( n37776 , n37313 , n37775 );
and ( n37777 , n37310 , n37776 );
or ( n37778 , n37309 , n37777 );
and ( n37779 , n37306 , n37778 );
or ( n37780 , n37305 , n37779 );
and ( n37781 , n37302 , n37780 );
or ( n37782 , n37301 , n37781 );
and ( n37783 , n37298 , n37782 );
or ( n37784 , n37297 , n37783 );
and ( n37785 , n37294 , n37784 );
or ( n37786 , n37293 , n37785 );
and ( n37787 , n37290 , n37786 );
or ( n37788 , n37289 , n37787 );
and ( n37789 , n37286 , n37788 );
or ( n37790 , n37285 , n37789 );
and ( n37791 , n37282 , n37790 );
or ( n37792 , n37281 , n37791 );
and ( n37793 , n37278 , n37792 );
or ( n37794 , n37277 , n37793 );
and ( n37795 , n37274 , n37794 );
or ( n37796 , n37273 , n37795 );
and ( n37797 , n37270 , n37796 );
or ( n37798 , n37269 , n37797 );
and ( n37799 , n37266 , n37798 );
or ( n37800 , n37265 , n37799 );
and ( n37801 , n37262 , n37800 );
or ( n37802 , n37261 , n37801 );
and ( n37803 , n37258 , n37802 );
or ( n37804 , n37257 , n37803 );
and ( n37805 , n37254 , n37804 );
or ( n37806 , n37253 , n37805 );
and ( n37807 , n37250 , n37806 );
or ( n37808 , n37249 , n37807 );
and ( n37809 , n37246 , n37808 );
or ( n37810 , n37245 , n37809 );
and ( n37811 , n37242 , n37810 );
or ( n37812 , n37241 , n37811 );
and ( n37813 , n37238 , n37812 );
or ( n37814 , n37237 , n37813 );
and ( n37815 , n37234 , n37814 );
or ( n37816 , n37233 , n37815 );
and ( n37817 , n37230 , n37816 );
or ( n37818 , n37229 , n37817 );
and ( n37819 , n37226 , n37818 );
or ( n37820 , n37225 , n37819 );
and ( n37821 , n37222 , n37820 );
or ( n37822 , n37221 , n37821 );
and ( n37823 , n37218 , n37822 );
or ( n37824 , n37217 , n37823 );
and ( n37825 , n37214 , n37824 );
or ( n37826 , n37213 , n37825 );
and ( n37827 , n37210 , n37826 );
or ( n37828 , n37209 , n37827 );
and ( n37829 , n37206 , n37828 );
or ( n37830 , n37205 , n37829 );
and ( n37831 , n37202 , n37830 );
or ( n37832 , n37201 , n37831 );
and ( n37833 , n37198 , n37832 );
or ( n37834 , n37197 , n37833 );
and ( n37835 , n37194 , n37834 );
or ( n37836 , n37193 , n37835 );
and ( n37837 , n37190 , n37836 );
or ( n37838 , n37189 , n37837 );
and ( n37839 , n37186 , n37838 );
or ( n37840 , n37185 , n37839 );
and ( n37841 , n37182 , n37840 );
or ( n37842 , n37181 , n37841 );
and ( n37843 , n37178 , n37842 );
or ( n37844 , n37177 , n37843 );
and ( n37845 , n37174 , n37844 );
or ( n37846 , n37173 , n37845 );
and ( n37847 , n37170 , n37846 );
or ( n37848 , n37169 , n37847 );
and ( n37849 , n37166 , n37848 );
or ( n37850 , n37165 , n37849 );
xor ( n37851 , n37162 , n37850 );
buf ( n37852 , n18082 );
and ( n37853 , n29839 , n37852 );
xor ( n37854 , n37851 , n37853 );
xor ( n37855 , n37166 , n37848 );
and ( n37856 , n29844 , n37852 );
and ( n37857 , n37855 , n37856 );
xor ( n37858 , n37855 , n37856 );
xor ( n37859 , n37170 , n37846 );
and ( n37860 , n29849 , n37852 );
and ( n37861 , n37859 , n37860 );
xor ( n37862 , n37859 , n37860 );
xor ( n37863 , n37174 , n37844 );
and ( n37864 , n29854 , n37852 );
and ( n37865 , n37863 , n37864 );
xor ( n37866 , n37863 , n37864 );
xor ( n37867 , n37178 , n37842 );
and ( n37868 , n29859 , n37852 );
and ( n37869 , n37867 , n37868 );
xor ( n37870 , n37867 , n37868 );
xor ( n37871 , n37182 , n37840 );
and ( n37872 , n29864 , n37852 );
and ( n37873 , n37871 , n37872 );
xor ( n37874 , n37871 , n37872 );
xor ( n37875 , n37186 , n37838 );
and ( n37876 , n29869 , n37852 );
and ( n37877 , n37875 , n37876 );
xor ( n37878 , n37875 , n37876 );
xor ( n37879 , n37190 , n37836 );
and ( n37880 , n29874 , n37852 );
and ( n37881 , n37879 , n37880 );
xor ( n37882 , n37879 , n37880 );
xor ( n37883 , n37194 , n37834 );
and ( n37884 , n29879 , n37852 );
and ( n37885 , n37883 , n37884 );
xor ( n37886 , n37883 , n37884 );
xor ( n37887 , n37198 , n37832 );
and ( n37888 , n29884 , n37852 );
and ( n37889 , n37887 , n37888 );
xor ( n37890 , n37887 , n37888 );
xor ( n37891 , n37202 , n37830 );
and ( n37892 , n29889 , n37852 );
and ( n37893 , n37891 , n37892 );
xor ( n37894 , n37891 , n37892 );
xor ( n37895 , n37206 , n37828 );
and ( n37896 , n29894 , n37852 );
and ( n37897 , n37895 , n37896 );
xor ( n37898 , n37895 , n37896 );
xor ( n37899 , n37210 , n37826 );
and ( n37900 , n29899 , n37852 );
and ( n37901 , n37899 , n37900 );
xor ( n37902 , n37899 , n37900 );
xor ( n37903 , n37214 , n37824 );
and ( n37904 , n29904 , n37852 );
and ( n37905 , n37903 , n37904 );
xor ( n37906 , n37903 , n37904 );
xor ( n37907 , n37218 , n37822 );
and ( n37908 , n29909 , n37852 );
and ( n37909 , n37907 , n37908 );
xor ( n37910 , n37907 , n37908 );
xor ( n37911 , n37222 , n37820 );
and ( n37912 , n29914 , n37852 );
and ( n37913 , n37911 , n37912 );
xor ( n37914 , n37911 , n37912 );
xor ( n37915 , n37226 , n37818 );
and ( n37916 , n29919 , n37852 );
and ( n37917 , n37915 , n37916 );
xor ( n37918 , n37915 , n37916 );
xor ( n37919 , n37230 , n37816 );
and ( n37920 , n29924 , n37852 );
and ( n37921 , n37919 , n37920 );
xor ( n37922 , n37919 , n37920 );
xor ( n37923 , n37234 , n37814 );
and ( n37924 , n29929 , n37852 );
and ( n37925 , n37923 , n37924 );
xor ( n37926 , n37923 , n37924 );
xor ( n37927 , n37238 , n37812 );
and ( n37928 , n29934 , n37852 );
and ( n37929 , n37927 , n37928 );
xor ( n37930 , n37927 , n37928 );
xor ( n37931 , n37242 , n37810 );
and ( n37932 , n29939 , n37852 );
and ( n37933 , n37931 , n37932 );
xor ( n37934 , n37931 , n37932 );
xor ( n37935 , n37246 , n37808 );
and ( n37936 , n29944 , n37852 );
and ( n37937 , n37935 , n37936 );
xor ( n37938 , n37935 , n37936 );
xor ( n37939 , n37250 , n37806 );
and ( n37940 , n29949 , n37852 );
and ( n37941 , n37939 , n37940 );
xor ( n37942 , n37939 , n37940 );
xor ( n37943 , n37254 , n37804 );
and ( n37944 , n29954 , n37852 );
and ( n37945 , n37943 , n37944 );
xor ( n37946 , n37943 , n37944 );
xor ( n37947 , n37258 , n37802 );
and ( n37948 , n29959 , n37852 );
and ( n37949 , n37947 , n37948 );
xor ( n37950 , n37947 , n37948 );
xor ( n37951 , n37262 , n37800 );
and ( n37952 , n29964 , n37852 );
and ( n37953 , n37951 , n37952 );
xor ( n37954 , n37951 , n37952 );
xor ( n37955 , n37266 , n37798 );
and ( n37956 , n29969 , n37852 );
and ( n37957 , n37955 , n37956 );
xor ( n37958 , n37955 , n37956 );
xor ( n37959 , n37270 , n37796 );
and ( n37960 , n29974 , n37852 );
and ( n37961 , n37959 , n37960 );
xor ( n37962 , n37959 , n37960 );
xor ( n37963 , n37274 , n37794 );
and ( n37964 , n29979 , n37852 );
and ( n37965 , n37963 , n37964 );
xor ( n37966 , n37963 , n37964 );
xor ( n37967 , n37278 , n37792 );
and ( n37968 , n29984 , n37852 );
and ( n37969 , n37967 , n37968 );
xor ( n37970 , n37967 , n37968 );
xor ( n37971 , n37282 , n37790 );
and ( n37972 , n29989 , n37852 );
and ( n37973 , n37971 , n37972 );
xor ( n37974 , n37971 , n37972 );
xor ( n37975 , n37286 , n37788 );
and ( n37976 , n29994 , n37852 );
and ( n37977 , n37975 , n37976 );
xor ( n37978 , n37975 , n37976 );
xor ( n37979 , n37290 , n37786 );
and ( n37980 , n29999 , n37852 );
and ( n37981 , n37979 , n37980 );
xor ( n37982 , n37979 , n37980 );
xor ( n37983 , n37294 , n37784 );
and ( n37984 , n30004 , n37852 );
and ( n37985 , n37983 , n37984 );
xor ( n37986 , n37983 , n37984 );
xor ( n37987 , n37298 , n37782 );
and ( n37988 , n30009 , n37852 );
and ( n37989 , n37987 , n37988 );
xor ( n37990 , n37987 , n37988 );
xor ( n37991 , n37302 , n37780 );
and ( n37992 , n30014 , n37852 );
and ( n37993 , n37991 , n37992 );
xor ( n37994 , n37991 , n37992 );
xor ( n37995 , n37306 , n37778 );
and ( n37996 , n30019 , n37852 );
and ( n37997 , n37995 , n37996 );
xor ( n37998 , n37995 , n37996 );
xor ( n37999 , n37310 , n37776 );
and ( n38000 , n30024 , n37852 );
and ( n38001 , n37999 , n38000 );
xor ( n38002 , n37999 , n38000 );
xor ( n38003 , n37314 , n37774 );
and ( n38004 , n30029 , n37852 );
and ( n38005 , n38003 , n38004 );
xor ( n38006 , n38003 , n38004 );
xor ( n38007 , n37318 , n37772 );
and ( n38008 , n30034 , n37852 );
and ( n38009 , n38007 , n38008 );
xor ( n38010 , n38007 , n38008 );
xor ( n38011 , n37322 , n37770 );
and ( n38012 , n30039 , n37852 );
and ( n38013 , n38011 , n38012 );
xor ( n38014 , n38011 , n38012 );
xor ( n38015 , n37326 , n37768 );
and ( n38016 , n30044 , n37852 );
and ( n38017 , n38015 , n38016 );
xor ( n38018 , n38015 , n38016 );
xor ( n38019 , n37330 , n37766 );
and ( n38020 , n30049 , n37852 );
and ( n38021 , n38019 , n38020 );
xor ( n38022 , n38019 , n38020 );
xor ( n38023 , n37334 , n37764 );
and ( n38024 , n30054 , n37852 );
and ( n38025 , n38023 , n38024 );
xor ( n38026 , n38023 , n38024 );
xor ( n38027 , n37338 , n37762 );
and ( n38028 , n30059 , n37852 );
and ( n38029 , n38027 , n38028 );
xor ( n38030 , n38027 , n38028 );
xor ( n38031 , n37342 , n37760 );
and ( n38032 , n30064 , n37852 );
and ( n38033 , n38031 , n38032 );
xor ( n38034 , n38031 , n38032 );
xor ( n38035 , n37346 , n37758 );
and ( n38036 , n30069 , n37852 );
and ( n38037 , n38035 , n38036 );
xor ( n38038 , n38035 , n38036 );
xor ( n38039 , n37350 , n37756 );
and ( n38040 , n30074 , n37852 );
and ( n38041 , n38039 , n38040 );
xor ( n38042 , n38039 , n38040 );
xor ( n38043 , n37354 , n37754 );
and ( n38044 , n30079 , n37852 );
and ( n38045 , n38043 , n38044 );
xor ( n38046 , n38043 , n38044 );
xor ( n38047 , n37358 , n37752 );
and ( n38048 , n30084 , n37852 );
and ( n38049 , n38047 , n38048 );
xor ( n38050 , n38047 , n38048 );
xor ( n38051 , n37362 , n37750 );
and ( n38052 , n30089 , n37852 );
and ( n38053 , n38051 , n38052 );
xor ( n38054 , n38051 , n38052 );
xor ( n38055 , n37366 , n37748 );
and ( n38056 , n30094 , n37852 );
and ( n38057 , n38055 , n38056 );
xor ( n38058 , n38055 , n38056 );
xor ( n38059 , n37370 , n37746 );
and ( n38060 , n30099 , n37852 );
and ( n38061 , n38059 , n38060 );
xor ( n38062 , n38059 , n38060 );
xor ( n38063 , n37374 , n37744 );
and ( n38064 , n30104 , n37852 );
and ( n38065 , n38063 , n38064 );
xor ( n38066 , n38063 , n38064 );
xor ( n38067 , n37378 , n37742 );
and ( n38068 , n30109 , n37852 );
and ( n38069 , n38067 , n38068 );
xor ( n38070 , n38067 , n38068 );
xor ( n38071 , n37382 , n37740 );
and ( n38072 , n30114 , n37852 );
and ( n38073 , n38071 , n38072 );
xor ( n38074 , n38071 , n38072 );
xor ( n38075 , n37386 , n37738 );
and ( n38076 , n30119 , n37852 );
and ( n38077 , n38075 , n38076 );
xor ( n38078 , n38075 , n38076 );
xor ( n38079 , n37390 , n37736 );
and ( n38080 , n30124 , n37852 );
and ( n38081 , n38079 , n38080 );
xor ( n38082 , n38079 , n38080 );
xor ( n38083 , n37394 , n37734 );
and ( n38084 , n30129 , n37852 );
and ( n38085 , n38083 , n38084 );
xor ( n38086 , n38083 , n38084 );
xor ( n38087 , n37398 , n37732 );
and ( n38088 , n30134 , n37852 );
and ( n38089 , n38087 , n38088 );
xor ( n38090 , n38087 , n38088 );
xor ( n38091 , n37402 , n37730 );
and ( n38092 , n30139 , n37852 );
and ( n38093 , n38091 , n38092 );
xor ( n38094 , n38091 , n38092 );
xor ( n38095 , n37406 , n37728 );
and ( n38096 , n30144 , n37852 );
and ( n38097 , n38095 , n38096 );
xor ( n38098 , n38095 , n38096 );
xor ( n38099 , n37410 , n37726 );
and ( n38100 , n30149 , n37852 );
and ( n38101 , n38099 , n38100 );
xor ( n38102 , n38099 , n38100 );
xor ( n38103 , n37414 , n37724 );
and ( n38104 , n30154 , n37852 );
and ( n38105 , n38103 , n38104 );
xor ( n38106 , n38103 , n38104 );
xor ( n38107 , n37418 , n37722 );
and ( n38108 , n30159 , n37852 );
and ( n38109 , n38107 , n38108 );
xor ( n38110 , n38107 , n38108 );
xor ( n38111 , n37422 , n37720 );
and ( n38112 , n30164 , n37852 );
and ( n38113 , n38111 , n38112 );
xor ( n38114 , n38111 , n38112 );
xor ( n38115 , n37426 , n37718 );
and ( n38116 , n30169 , n37852 );
and ( n38117 , n38115 , n38116 );
xor ( n38118 , n38115 , n38116 );
xor ( n38119 , n37430 , n37716 );
and ( n38120 , n30174 , n37852 );
and ( n38121 , n38119 , n38120 );
xor ( n38122 , n38119 , n38120 );
xor ( n38123 , n37434 , n37714 );
and ( n38124 , n30179 , n37852 );
and ( n38125 , n38123 , n38124 );
xor ( n38126 , n38123 , n38124 );
xor ( n38127 , n37438 , n37712 );
and ( n38128 , n30184 , n37852 );
and ( n38129 , n38127 , n38128 );
xor ( n38130 , n38127 , n38128 );
xor ( n38131 , n37442 , n37710 );
and ( n38132 , n30189 , n37852 );
and ( n38133 , n38131 , n38132 );
xor ( n38134 , n38131 , n38132 );
xor ( n38135 , n37446 , n37708 );
and ( n38136 , n30194 , n37852 );
and ( n38137 , n38135 , n38136 );
xor ( n38138 , n38135 , n38136 );
xor ( n38139 , n37450 , n37706 );
and ( n38140 , n30199 , n37852 );
and ( n38141 , n38139 , n38140 );
xor ( n38142 , n38139 , n38140 );
xor ( n38143 , n37454 , n37704 );
and ( n38144 , n30204 , n37852 );
and ( n38145 , n38143 , n38144 );
xor ( n38146 , n38143 , n38144 );
xor ( n38147 , n37458 , n37702 );
and ( n38148 , n30209 , n37852 );
and ( n38149 , n38147 , n38148 );
xor ( n38150 , n38147 , n38148 );
xor ( n38151 , n37462 , n37700 );
and ( n38152 , n30214 , n37852 );
and ( n38153 , n38151 , n38152 );
xor ( n38154 , n38151 , n38152 );
xor ( n38155 , n37466 , n37698 );
and ( n38156 , n30219 , n37852 );
and ( n38157 , n38155 , n38156 );
xor ( n38158 , n38155 , n38156 );
xor ( n38159 , n37470 , n37696 );
and ( n38160 , n30224 , n37852 );
and ( n38161 , n38159 , n38160 );
xor ( n38162 , n38159 , n38160 );
xor ( n38163 , n37474 , n37694 );
and ( n38164 , n30229 , n37852 );
and ( n38165 , n38163 , n38164 );
xor ( n38166 , n38163 , n38164 );
xor ( n38167 , n37478 , n37692 );
and ( n38168 , n30234 , n37852 );
and ( n38169 , n38167 , n38168 );
xor ( n38170 , n38167 , n38168 );
xor ( n38171 , n37482 , n37690 );
and ( n38172 , n30239 , n37852 );
and ( n38173 , n38171 , n38172 );
xor ( n38174 , n38171 , n38172 );
xor ( n38175 , n37486 , n37688 );
and ( n38176 , n30244 , n37852 );
and ( n38177 , n38175 , n38176 );
xor ( n38178 , n38175 , n38176 );
xor ( n38179 , n37490 , n37686 );
and ( n38180 , n30249 , n37852 );
and ( n38181 , n38179 , n38180 );
xor ( n38182 , n38179 , n38180 );
xor ( n38183 , n37494 , n37684 );
and ( n38184 , n30254 , n37852 );
and ( n38185 , n38183 , n38184 );
xor ( n38186 , n38183 , n38184 );
xor ( n38187 , n37498 , n37682 );
and ( n38188 , n30259 , n37852 );
and ( n38189 , n38187 , n38188 );
xor ( n38190 , n38187 , n38188 );
xor ( n38191 , n37502 , n37680 );
and ( n38192 , n30264 , n37852 );
and ( n38193 , n38191 , n38192 );
xor ( n38194 , n38191 , n38192 );
xor ( n38195 , n37506 , n37678 );
and ( n38196 , n30269 , n37852 );
and ( n38197 , n38195 , n38196 );
xor ( n38198 , n38195 , n38196 );
xor ( n38199 , n37510 , n37676 );
and ( n38200 , n30274 , n37852 );
and ( n38201 , n38199 , n38200 );
xor ( n38202 , n38199 , n38200 );
xor ( n38203 , n37514 , n37674 );
and ( n38204 , n30279 , n37852 );
and ( n38205 , n38203 , n38204 );
xor ( n38206 , n38203 , n38204 );
xor ( n38207 , n37518 , n37672 );
and ( n38208 , n30284 , n37852 );
and ( n38209 , n38207 , n38208 );
xor ( n38210 , n38207 , n38208 );
xor ( n38211 , n37522 , n37670 );
and ( n38212 , n30289 , n37852 );
and ( n38213 , n38211 , n38212 );
xor ( n38214 , n38211 , n38212 );
xor ( n38215 , n37526 , n37668 );
and ( n38216 , n30294 , n37852 );
and ( n38217 , n38215 , n38216 );
xor ( n38218 , n38215 , n38216 );
xor ( n38219 , n37530 , n37666 );
and ( n38220 , n30299 , n37852 );
and ( n38221 , n38219 , n38220 );
xor ( n38222 , n38219 , n38220 );
xor ( n38223 , n37534 , n37664 );
and ( n38224 , n30304 , n37852 );
and ( n38225 , n38223 , n38224 );
xor ( n38226 , n38223 , n38224 );
xor ( n38227 , n37538 , n37662 );
and ( n38228 , n30309 , n37852 );
and ( n38229 , n38227 , n38228 );
xor ( n38230 , n38227 , n38228 );
xor ( n38231 , n37542 , n37660 );
and ( n38232 , n30314 , n37852 );
and ( n38233 , n38231 , n38232 );
xor ( n38234 , n38231 , n38232 );
xor ( n38235 , n37546 , n37658 );
and ( n38236 , n30319 , n37852 );
and ( n38237 , n38235 , n38236 );
xor ( n38238 , n38235 , n38236 );
xor ( n38239 , n37550 , n37656 );
and ( n38240 , n30324 , n37852 );
and ( n38241 , n38239 , n38240 );
xor ( n38242 , n38239 , n38240 );
xor ( n38243 , n37554 , n37654 );
and ( n38244 , n30329 , n37852 );
and ( n38245 , n38243 , n38244 );
xor ( n38246 , n38243 , n38244 );
xor ( n38247 , n37558 , n37652 );
and ( n38248 , n30334 , n37852 );
and ( n38249 , n38247 , n38248 );
xor ( n38250 , n38247 , n38248 );
xor ( n38251 , n37562 , n37650 );
and ( n38252 , n30339 , n37852 );
and ( n38253 , n38251 , n38252 );
xor ( n38254 , n38251 , n38252 );
xor ( n38255 , n37566 , n37648 );
and ( n38256 , n30344 , n37852 );
and ( n38257 , n38255 , n38256 );
xor ( n38258 , n38255 , n38256 );
xor ( n38259 , n37570 , n37646 );
and ( n38260 , n30349 , n37852 );
and ( n38261 , n38259 , n38260 );
xor ( n38262 , n38259 , n38260 );
xor ( n38263 , n37574 , n37644 );
and ( n38264 , n30354 , n37852 );
and ( n38265 , n38263 , n38264 );
xor ( n38266 , n38263 , n38264 );
xor ( n38267 , n37578 , n37642 );
and ( n38268 , n30359 , n37852 );
and ( n38269 , n38267 , n38268 );
xor ( n38270 , n38267 , n38268 );
xor ( n38271 , n37582 , n37640 );
and ( n38272 , n30364 , n37852 );
and ( n38273 , n38271 , n38272 );
xor ( n38274 , n38271 , n38272 );
xor ( n38275 , n37586 , n37638 );
and ( n38276 , n30369 , n37852 );
and ( n38277 , n38275 , n38276 );
xor ( n38278 , n38275 , n38276 );
xor ( n38279 , n37590 , n37636 );
and ( n38280 , n30374 , n37852 );
and ( n38281 , n38279 , n38280 );
xor ( n38282 , n38279 , n38280 );
xor ( n38283 , n37594 , n37634 );
and ( n38284 , n30379 , n37852 );
and ( n38285 , n38283 , n38284 );
xor ( n38286 , n38283 , n38284 );
xor ( n38287 , n37598 , n37632 );
and ( n38288 , n30384 , n37852 );
and ( n38289 , n38287 , n38288 );
xor ( n38290 , n38287 , n38288 );
xor ( n38291 , n37602 , n37630 );
and ( n38292 , n30389 , n37852 );
and ( n38293 , n38291 , n38292 );
xor ( n38294 , n38291 , n38292 );
xor ( n38295 , n37606 , n37628 );
and ( n38296 , n30394 , n37852 );
and ( n38297 , n38295 , n38296 );
xor ( n38298 , n38295 , n38296 );
xor ( n38299 , n37610 , n37626 );
and ( n38300 , n30399 , n37852 );
and ( n38301 , n38299 , n38300 );
xor ( n38302 , n38299 , n38300 );
xor ( n38303 , n37614 , n37624 );
and ( n38304 , n30404 , n37852 );
and ( n38305 , n38303 , n38304 );
xor ( n38306 , n38303 , n38304 );
xor ( n38307 , n37618 , n37622 );
and ( n38308 , n30409 , n37852 );
and ( n38309 , n38307 , n38308 );
buf ( n38310 , n38309 );
and ( n38311 , n38306 , n38310 );
or ( n38312 , n38305 , n38311 );
and ( n38313 , n38302 , n38312 );
or ( n38314 , n38301 , n38313 );
and ( n38315 , n38298 , n38314 );
or ( n38316 , n38297 , n38315 );
and ( n38317 , n38294 , n38316 );
or ( n38318 , n38293 , n38317 );
and ( n38319 , n38290 , n38318 );
or ( n38320 , n38289 , n38319 );
and ( n38321 , n38286 , n38320 );
or ( n38322 , n38285 , n38321 );
and ( n38323 , n38282 , n38322 );
or ( n38324 , n38281 , n38323 );
and ( n38325 , n38278 , n38324 );
or ( n38326 , n38277 , n38325 );
and ( n38327 , n38274 , n38326 );
or ( n38328 , n38273 , n38327 );
and ( n38329 , n38270 , n38328 );
or ( n38330 , n38269 , n38329 );
and ( n38331 , n38266 , n38330 );
or ( n38332 , n38265 , n38331 );
and ( n38333 , n38262 , n38332 );
or ( n38334 , n38261 , n38333 );
and ( n38335 , n38258 , n38334 );
or ( n38336 , n38257 , n38335 );
and ( n38337 , n38254 , n38336 );
or ( n38338 , n38253 , n38337 );
and ( n38339 , n38250 , n38338 );
or ( n38340 , n38249 , n38339 );
and ( n38341 , n38246 , n38340 );
or ( n38342 , n38245 , n38341 );
and ( n38343 , n38242 , n38342 );
or ( n38344 , n38241 , n38343 );
and ( n38345 , n38238 , n38344 );
or ( n38346 , n38237 , n38345 );
and ( n38347 , n38234 , n38346 );
or ( n38348 , n38233 , n38347 );
and ( n38349 , n38230 , n38348 );
or ( n38350 , n38229 , n38349 );
and ( n38351 , n38226 , n38350 );
or ( n38352 , n38225 , n38351 );
and ( n38353 , n38222 , n38352 );
or ( n38354 , n38221 , n38353 );
and ( n38355 , n38218 , n38354 );
or ( n38356 , n38217 , n38355 );
and ( n38357 , n38214 , n38356 );
or ( n38358 , n38213 , n38357 );
and ( n38359 , n38210 , n38358 );
or ( n38360 , n38209 , n38359 );
and ( n38361 , n38206 , n38360 );
or ( n38362 , n38205 , n38361 );
and ( n38363 , n38202 , n38362 );
or ( n38364 , n38201 , n38363 );
and ( n38365 , n38198 , n38364 );
or ( n38366 , n38197 , n38365 );
and ( n38367 , n38194 , n38366 );
or ( n38368 , n38193 , n38367 );
and ( n38369 , n38190 , n38368 );
or ( n38370 , n38189 , n38369 );
and ( n38371 , n38186 , n38370 );
or ( n38372 , n38185 , n38371 );
and ( n38373 , n38182 , n38372 );
or ( n38374 , n38181 , n38373 );
and ( n38375 , n38178 , n38374 );
or ( n38376 , n38177 , n38375 );
and ( n38377 , n38174 , n38376 );
or ( n38378 , n38173 , n38377 );
and ( n38379 , n38170 , n38378 );
or ( n38380 , n38169 , n38379 );
and ( n38381 , n38166 , n38380 );
or ( n38382 , n38165 , n38381 );
and ( n38383 , n38162 , n38382 );
or ( n38384 , n38161 , n38383 );
and ( n38385 , n38158 , n38384 );
or ( n38386 , n38157 , n38385 );
and ( n38387 , n38154 , n38386 );
or ( n38388 , n38153 , n38387 );
and ( n38389 , n38150 , n38388 );
or ( n38390 , n38149 , n38389 );
and ( n38391 , n38146 , n38390 );
or ( n38392 , n38145 , n38391 );
and ( n38393 , n38142 , n38392 );
or ( n38394 , n38141 , n38393 );
and ( n38395 , n38138 , n38394 );
or ( n38396 , n38137 , n38395 );
and ( n38397 , n38134 , n38396 );
or ( n38398 , n38133 , n38397 );
and ( n38399 , n38130 , n38398 );
or ( n38400 , n38129 , n38399 );
and ( n38401 , n38126 , n38400 );
or ( n38402 , n38125 , n38401 );
and ( n38403 , n38122 , n38402 );
or ( n38404 , n38121 , n38403 );
and ( n38405 , n38118 , n38404 );
or ( n38406 , n38117 , n38405 );
and ( n38407 , n38114 , n38406 );
or ( n38408 , n38113 , n38407 );
and ( n38409 , n38110 , n38408 );
or ( n38410 , n38109 , n38409 );
and ( n38411 , n38106 , n38410 );
or ( n38412 , n38105 , n38411 );
and ( n38413 , n38102 , n38412 );
or ( n38414 , n38101 , n38413 );
and ( n38415 , n38098 , n38414 );
or ( n38416 , n38097 , n38415 );
and ( n38417 , n38094 , n38416 );
or ( n38418 , n38093 , n38417 );
and ( n38419 , n38090 , n38418 );
or ( n38420 , n38089 , n38419 );
and ( n38421 , n38086 , n38420 );
or ( n38422 , n38085 , n38421 );
and ( n38423 , n38082 , n38422 );
or ( n38424 , n38081 , n38423 );
and ( n38425 , n38078 , n38424 );
or ( n38426 , n38077 , n38425 );
and ( n38427 , n38074 , n38426 );
or ( n38428 , n38073 , n38427 );
and ( n38429 , n38070 , n38428 );
or ( n38430 , n38069 , n38429 );
and ( n38431 , n38066 , n38430 );
or ( n38432 , n38065 , n38431 );
and ( n38433 , n38062 , n38432 );
or ( n38434 , n38061 , n38433 );
and ( n38435 , n38058 , n38434 );
or ( n38436 , n38057 , n38435 );
and ( n38437 , n38054 , n38436 );
or ( n38438 , n38053 , n38437 );
and ( n38439 , n38050 , n38438 );
or ( n38440 , n38049 , n38439 );
and ( n38441 , n38046 , n38440 );
or ( n38442 , n38045 , n38441 );
and ( n38443 , n38042 , n38442 );
or ( n38444 , n38041 , n38443 );
and ( n38445 , n38038 , n38444 );
or ( n38446 , n38037 , n38445 );
and ( n38447 , n38034 , n38446 );
or ( n38448 , n38033 , n38447 );
and ( n38449 , n38030 , n38448 );
or ( n38450 , n38029 , n38449 );
and ( n38451 , n38026 , n38450 );
or ( n38452 , n38025 , n38451 );
and ( n38453 , n38022 , n38452 );
or ( n38454 , n38021 , n38453 );
and ( n38455 , n38018 , n38454 );
or ( n38456 , n38017 , n38455 );
and ( n38457 , n38014 , n38456 );
or ( n38458 , n38013 , n38457 );
and ( n38459 , n38010 , n38458 );
or ( n38460 , n38009 , n38459 );
and ( n38461 , n38006 , n38460 );
or ( n38462 , n38005 , n38461 );
and ( n38463 , n38002 , n38462 );
or ( n38464 , n38001 , n38463 );
and ( n38465 , n37998 , n38464 );
or ( n38466 , n37997 , n38465 );
and ( n38467 , n37994 , n38466 );
or ( n38468 , n37993 , n38467 );
and ( n38469 , n37990 , n38468 );
or ( n38470 , n37989 , n38469 );
and ( n38471 , n37986 , n38470 );
or ( n38472 , n37985 , n38471 );
and ( n38473 , n37982 , n38472 );
or ( n38474 , n37981 , n38473 );
and ( n38475 , n37978 , n38474 );
or ( n38476 , n37977 , n38475 );
and ( n38477 , n37974 , n38476 );
or ( n38478 , n37973 , n38477 );
and ( n38479 , n37970 , n38478 );
or ( n38480 , n37969 , n38479 );
and ( n38481 , n37966 , n38480 );
or ( n38482 , n37965 , n38481 );
and ( n38483 , n37962 , n38482 );
or ( n38484 , n37961 , n38483 );
and ( n38485 , n37958 , n38484 );
or ( n38486 , n37957 , n38485 );
and ( n38487 , n37954 , n38486 );
or ( n38488 , n37953 , n38487 );
and ( n38489 , n37950 , n38488 );
or ( n38490 , n37949 , n38489 );
and ( n38491 , n37946 , n38490 );
or ( n38492 , n37945 , n38491 );
and ( n38493 , n37942 , n38492 );
or ( n38494 , n37941 , n38493 );
and ( n38495 , n37938 , n38494 );
or ( n38496 , n37937 , n38495 );
and ( n38497 , n37934 , n38496 );
or ( n38498 , n37933 , n38497 );
and ( n38499 , n37930 , n38498 );
or ( n38500 , n37929 , n38499 );
and ( n38501 , n37926 , n38500 );
or ( n38502 , n37925 , n38501 );
and ( n38503 , n37922 , n38502 );
or ( n38504 , n37921 , n38503 );
and ( n38505 , n37918 , n38504 );
or ( n38506 , n37917 , n38505 );
and ( n38507 , n37914 , n38506 );
or ( n38508 , n37913 , n38507 );
and ( n38509 , n37910 , n38508 );
or ( n38510 , n37909 , n38509 );
and ( n38511 , n37906 , n38510 );
or ( n38512 , n37905 , n38511 );
and ( n38513 , n37902 , n38512 );
or ( n38514 , n37901 , n38513 );
and ( n38515 , n37898 , n38514 );
or ( n38516 , n37897 , n38515 );
and ( n38517 , n37894 , n38516 );
or ( n38518 , n37893 , n38517 );
and ( n38519 , n37890 , n38518 );
or ( n38520 , n37889 , n38519 );
and ( n38521 , n37886 , n38520 );
or ( n38522 , n37885 , n38521 );
and ( n38523 , n37882 , n38522 );
or ( n38524 , n37881 , n38523 );
and ( n38525 , n37878 , n38524 );
or ( n38526 , n37877 , n38525 );
and ( n38527 , n37874 , n38526 );
or ( n38528 , n37873 , n38527 );
and ( n38529 , n37870 , n38528 );
or ( n38530 , n37869 , n38529 );
and ( n38531 , n37866 , n38530 );
or ( n38532 , n37865 , n38531 );
and ( n38533 , n37862 , n38532 );
or ( n38534 , n37861 , n38533 );
and ( n38535 , n37858 , n38534 );
or ( n38536 , n37857 , n38535 );
xor ( n38537 , n37854 , n38536 );
buf ( n38538 , n18080 );
and ( n38539 , n29844 , n38538 );
xor ( n38540 , n38537 , n38539 );
xor ( n38541 , n37858 , n38534 );
and ( n38542 , n29849 , n38538 );
and ( n38543 , n38541 , n38542 );
xor ( n38544 , n38541 , n38542 );
xor ( n38545 , n37862 , n38532 );
and ( n38546 , n29854 , n38538 );
and ( n38547 , n38545 , n38546 );
xor ( n38548 , n38545 , n38546 );
xor ( n38549 , n37866 , n38530 );
and ( n38550 , n29859 , n38538 );
and ( n38551 , n38549 , n38550 );
xor ( n38552 , n38549 , n38550 );
xor ( n38553 , n37870 , n38528 );
and ( n38554 , n29864 , n38538 );
and ( n38555 , n38553 , n38554 );
xor ( n38556 , n38553 , n38554 );
xor ( n38557 , n37874 , n38526 );
and ( n38558 , n29869 , n38538 );
and ( n38559 , n38557 , n38558 );
xor ( n38560 , n38557 , n38558 );
xor ( n38561 , n37878 , n38524 );
and ( n38562 , n29874 , n38538 );
and ( n38563 , n38561 , n38562 );
xor ( n38564 , n38561 , n38562 );
xor ( n38565 , n37882 , n38522 );
and ( n38566 , n29879 , n38538 );
and ( n38567 , n38565 , n38566 );
xor ( n38568 , n38565 , n38566 );
xor ( n38569 , n37886 , n38520 );
and ( n38570 , n29884 , n38538 );
and ( n38571 , n38569 , n38570 );
xor ( n38572 , n38569 , n38570 );
xor ( n38573 , n37890 , n38518 );
and ( n38574 , n29889 , n38538 );
and ( n38575 , n38573 , n38574 );
xor ( n38576 , n38573 , n38574 );
xor ( n38577 , n37894 , n38516 );
and ( n38578 , n29894 , n38538 );
and ( n38579 , n38577 , n38578 );
xor ( n38580 , n38577 , n38578 );
xor ( n38581 , n37898 , n38514 );
and ( n38582 , n29899 , n38538 );
and ( n38583 , n38581 , n38582 );
xor ( n38584 , n38581 , n38582 );
xor ( n38585 , n37902 , n38512 );
and ( n38586 , n29904 , n38538 );
and ( n38587 , n38585 , n38586 );
xor ( n38588 , n38585 , n38586 );
xor ( n38589 , n37906 , n38510 );
and ( n38590 , n29909 , n38538 );
and ( n38591 , n38589 , n38590 );
xor ( n38592 , n38589 , n38590 );
xor ( n38593 , n37910 , n38508 );
and ( n38594 , n29914 , n38538 );
and ( n38595 , n38593 , n38594 );
xor ( n38596 , n38593 , n38594 );
xor ( n38597 , n37914 , n38506 );
and ( n38598 , n29919 , n38538 );
and ( n38599 , n38597 , n38598 );
xor ( n38600 , n38597 , n38598 );
xor ( n38601 , n37918 , n38504 );
and ( n38602 , n29924 , n38538 );
and ( n38603 , n38601 , n38602 );
xor ( n38604 , n38601 , n38602 );
xor ( n38605 , n37922 , n38502 );
and ( n38606 , n29929 , n38538 );
and ( n38607 , n38605 , n38606 );
xor ( n38608 , n38605 , n38606 );
xor ( n38609 , n37926 , n38500 );
and ( n38610 , n29934 , n38538 );
and ( n38611 , n38609 , n38610 );
xor ( n38612 , n38609 , n38610 );
xor ( n38613 , n37930 , n38498 );
and ( n38614 , n29939 , n38538 );
and ( n38615 , n38613 , n38614 );
xor ( n38616 , n38613 , n38614 );
xor ( n38617 , n37934 , n38496 );
and ( n38618 , n29944 , n38538 );
and ( n38619 , n38617 , n38618 );
xor ( n38620 , n38617 , n38618 );
xor ( n38621 , n37938 , n38494 );
and ( n38622 , n29949 , n38538 );
and ( n38623 , n38621 , n38622 );
xor ( n38624 , n38621 , n38622 );
xor ( n38625 , n37942 , n38492 );
and ( n38626 , n29954 , n38538 );
and ( n38627 , n38625 , n38626 );
xor ( n38628 , n38625 , n38626 );
xor ( n38629 , n37946 , n38490 );
and ( n38630 , n29959 , n38538 );
and ( n38631 , n38629 , n38630 );
xor ( n38632 , n38629 , n38630 );
xor ( n38633 , n37950 , n38488 );
and ( n38634 , n29964 , n38538 );
and ( n38635 , n38633 , n38634 );
xor ( n38636 , n38633 , n38634 );
xor ( n38637 , n37954 , n38486 );
and ( n38638 , n29969 , n38538 );
and ( n38639 , n38637 , n38638 );
xor ( n38640 , n38637 , n38638 );
xor ( n38641 , n37958 , n38484 );
and ( n38642 , n29974 , n38538 );
and ( n38643 , n38641 , n38642 );
xor ( n38644 , n38641 , n38642 );
xor ( n38645 , n37962 , n38482 );
and ( n38646 , n29979 , n38538 );
and ( n38647 , n38645 , n38646 );
xor ( n38648 , n38645 , n38646 );
xor ( n38649 , n37966 , n38480 );
and ( n38650 , n29984 , n38538 );
and ( n38651 , n38649 , n38650 );
xor ( n38652 , n38649 , n38650 );
xor ( n38653 , n37970 , n38478 );
and ( n38654 , n29989 , n38538 );
and ( n38655 , n38653 , n38654 );
xor ( n38656 , n38653 , n38654 );
xor ( n38657 , n37974 , n38476 );
and ( n38658 , n29994 , n38538 );
and ( n38659 , n38657 , n38658 );
xor ( n38660 , n38657 , n38658 );
xor ( n38661 , n37978 , n38474 );
and ( n38662 , n29999 , n38538 );
and ( n38663 , n38661 , n38662 );
xor ( n38664 , n38661 , n38662 );
xor ( n38665 , n37982 , n38472 );
and ( n38666 , n30004 , n38538 );
and ( n38667 , n38665 , n38666 );
xor ( n38668 , n38665 , n38666 );
xor ( n38669 , n37986 , n38470 );
and ( n38670 , n30009 , n38538 );
and ( n38671 , n38669 , n38670 );
xor ( n38672 , n38669 , n38670 );
xor ( n38673 , n37990 , n38468 );
and ( n38674 , n30014 , n38538 );
and ( n38675 , n38673 , n38674 );
xor ( n38676 , n38673 , n38674 );
xor ( n38677 , n37994 , n38466 );
and ( n38678 , n30019 , n38538 );
and ( n38679 , n38677 , n38678 );
xor ( n38680 , n38677 , n38678 );
xor ( n38681 , n37998 , n38464 );
and ( n38682 , n30024 , n38538 );
and ( n38683 , n38681 , n38682 );
xor ( n38684 , n38681 , n38682 );
xor ( n38685 , n38002 , n38462 );
and ( n38686 , n30029 , n38538 );
and ( n38687 , n38685 , n38686 );
xor ( n38688 , n38685 , n38686 );
xor ( n38689 , n38006 , n38460 );
and ( n38690 , n30034 , n38538 );
and ( n38691 , n38689 , n38690 );
xor ( n38692 , n38689 , n38690 );
xor ( n38693 , n38010 , n38458 );
and ( n38694 , n30039 , n38538 );
and ( n38695 , n38693 , n38694 );
xor ( n38696 , n38693 , n38694 );
xor ( n38697 , n38014 , n38456 );
and ( n38698 , n30044 , n38538 );
and ( n38699 , n38697 , n38698 );
xor ( n38700 , n38697 , n38698 );
xor ( n38701 , n38018 , n38454 );
and ( n38702 , n30049 , n38538 );
and ( n38703 , n38701 , n38702 );
xor ( n38704 , n38701 , n38702 );
xor ( n38705 , n38022 , n38452 );
and ( n38706 , n30054 , n38538 );
and ( n38707 , n38705 , n38706 );
xor ( n38708 , n38705 , n38706 );
xor ( n38709 , n38026 , n38450 );
and ( n38710 , n30059 , n38538 );
and ( n38711 , n38709 , n38710 );
xor ( n38712 , n38709 , n38710 );
xor ( n38713 , n38030 , n38448 );
and ( n38714 , n30064 , n38538 );
and ( n38715 , n38713 , n38714 );
xor ( n38716 , n38713 , n38714 );
xor ( n38717 , n38034 , n38446 );
and ( n38718 , n30069 , n38538 );
and ( n38719 , n38717 , n38718 );
xor ( n38720 , n38717 , n38718 );
xor ( n38721 , n38038 , n38444 );
and ( n38722 , n30074 , n38538 );
and ( n38723 , n38721 , n38722 );
xor ( n38724 , n38721 , n38722 );
xor ( n38725 , n38042 , n38442 );
and ( n38726 , n30079 , n38538 );
and ( n38727 , n38725 , n38726 );
xor ( n38728 , n38725 , n38726 );
xor ( n38729 , n38046 , n38440 );
and ( n38730 , n30084 , n38538 );
and ( n38731 , n38729 , n38730 );
xor ( n38732 , n38729 , n38730 );
xor ( n38733 , n38050 , n38438 );
and ( n38734 , n30089 , n38538 );
and ( n38735 , n38733 , n38734 );
xor ( n38736 , n38733 , n38734 );
xor ( n38737 , n38054 , n38436 );
and ( n38738 , n30094 , n38538 );
and ( n38739 , n38737 , n38738 );
xor ( n38740 , n38737 , n38738 );
xor ( n38741 , n38058 , n38434 );
and ( n38742 , n30099 , n38538 );
and ( n38743 , n38741 , n38742 );
xor ( n38744 , n38741 , n38742 );
xor ( n38745 , n38062 , n38432 );
and ( n38746 , n30104 , n38538 );
and ( n38747 , n38745 , n38746 );
xor ( n38748 , n38745 , n38746 );
xor ( n38749 , n38066 , n38430 );
and ( n38750 , n30109 , n38538 );
and ( n38751 , n38749 , n38750 );
xor ( n38752 , n38749 , n38750 );
xor ( n38753 , n38070 , n38428 );
and ( n38754 , n30114 , n38538 );
and ( n38755 , n38753 , n38754 );
xor ( n38756 , n38753 , n38754 );
xor ( n38757 , n38074 , n38426 );
and ( n38758 , n30119 , n38538 );
and ( n38759 , n38757 , n38758 );
xor ( n38760 , n38757 , n38758 );
xor ( n38761 , n38078 , n38424 );
and ( n38762 , n30124 , n38538 );
and ( n38763 , n38761 , n38762 );
xor ( n38764 , n38761 , n38762 );
xor ( n38765 , n38082 , n38422 );
and ( n38766 , n30129 , n38538 );
and ( n38767 , n38765 , n38766 );
xor ( n38768 , n38765 , n38766 );
xor ( n38769 , n38086 , n38420 );
and ( n38770 , n30134 , n38538 );
and ( n38771 , n38769 , n38770 );
xor ( n38772 , n38769 , n38770 );
xor ( n38773 , n38090 , n38418 );
and ( n38774 , n30139 , n38538 );
and ( n38775 , n38773 , n38774 );
xor ( n38776 , n38773 , n38774 );
xor ( n38777 , n38094 , n38416 );
and ( n38778 , n30144 , n38538 );
and ( n38779 , n38777 , n38778 );
xor ( n38780 , n38777 , n38778 );
xor ( n38781 , n38098 , n38414 );
and ( n38782 , n30149 , n38538 );
and ( n38783 , n38781 , n38782 );
xor ( n38784 , n38781 , n38782 );
xor ( n38785 , n38102 , n38412 );
and ( n38786 , n30154 , n38538 );
and ( n38787 , n38785 , n38786 );
xor ( n38788 , n38785 , n38786 );
xor ( n38789 , n38106 , n38410 );
and ( n38790 , n30159 , n38538 );
and ( n38791 , n38789 , n38790 );
xor ( n38792 , n38789 , n38790 );
xor ( n38793 , n38110 , n38408 );
and ( n38794 , n30164 , n38538 );
and ( n38795 , n38793 , n38794 );
xor ( n38796 , n38793 , n38794 );
xor ( n38797 , n38114 , n38406 );
and ( n38798 , n30169 , n38538 );
and ( n38799 , n38797 , n38798 );
xor ( n38800 , n38797 , n38798 );
xor ( n38801 , n38118 , n38404 );
and ( n38802 , n30174 , n38538 );
and ( n38803 , n38801 , n38802 );
xor ( n38804 , n38801 , n38802 );
xor ( n38805 , n38122 , n38402 );
and ( n38806 , n30179 , n38538 );
and ( n38807 , n38805 , n38806 );
xor ( n38808 , n38805 , n38806 );
xor ( n38809 , n38126 , n38400 );
and ( n38810 , n30184 , n38538 );
and ( n38811 , n38809 , n38810 );
xor ( n38812 , n38809 , n38810 );
xor ( n38813 , n38130 , n38398 );
and ( n38814 , n30189 , n38538 );
and ( n38815 , n38813 , n38814 );
xor ( n38816 , n38813 , n38814 );
xor ( n38817 , n38134 , n38396 );
and ( n38818 , n30194 , n38538 );
and ( n38819 , n38817 , n38818 );
xor ( n38820 , n38817 , n38818 );
xor ( n38821 , n38138 , n38394 );
and ( n38822 , n30199 , n38538 );
and ( n38823 , n38821 , n38822 );
xor ( n38824 , n38821 , n38822 );
xor ( n38825 , n38142 , n38392 );
and ( n38826 , n30204 , n38538 );
and ( n38827 , n38825 , n38826 );
xor ( n38828 , n38825 , n38826 );
xor ( n38829 , n38146 , n38390 );
and ( n38830 , n30209 , n38538 );
and ( n38831 , n38829 , n38830 );
xor ( n38832 , n38829 , n38830 );
xor ( n38833 , n38150 , n38388 );
and ( n38834 , n30214 , n38538 );
and ( n38835 , n38833 , n38834 );
xor ( n38836 , n38833 , n38834 );
xor ( n38837 , n38154 , n38386 );
and ( n38838 , n30219 , n38538 );
and ( n38839 , n38837 , n38838 );
xor ( n38840 , n38837 , n38838 );
xor ( n38841 , n38158 , n38384 );
and ( n38842 , n30224 , n38538 );
and ( n38843 , n38841 , n38842 );
xor ( n38844 , n38841 , n38842 );
xor ( n38845 , n38162 , n38382 );
and ( n38846 , n30229 , n38538 );
and ( n38847 , n38845 , n38846 );
xor ( n38848 , n38845 , n38846 );
xor ( n38849 , n38166 , n38380 );
and ( n38850 , n30234 , n38538 );
and ( n38851 , n38849 , n38850 );
xor ( n38852 , n38849 , n38850 );
xor ( n38853 , n38170 , n38378 );
and ( n38854 , n30239 , n38538 );
and ( n38855 , n38853 , n38854 );
xor ( n38856 , n38853 , n38854 );
xor ( n38857 , n38174 , n38376 );
and ( n38858 , n30244 , n38538 );
and ( n38859 , n38857 , n38858 );
xor ( n38860 , n38857 , n38858 );
xor ( n38861 , n38178 , n38374 );
and ( n38862 , n30249 , n38538 );
and ( n38863 , n38861 , n38862 );
xor ( n38864 , n38861 , n38862 );
xor ( n38865 , n38182 , n38372 );
and ( n38866 , n30254 , n38538 );
and ( n38867 , n38865 , n38866 );
xor ( n38868 , n38865 , n38866 );
xor ( n38869 , n38186 , n38370 );
and ( n38870 , n30259 , n38538 );
and ( n38871 , n38869 , n38870 );
xor ( n38872 , n38869 , n38870 );
xor ( n38873 , n38190 , n38368 );
and ( n38874 , n30264 , n38538 );
and ( n38875 , n38873 , n38874 );
xor ( n38876 , n38873 , n38874 );
xor ( n38877 , n38194 , n38366 );
and ( n38878 , n30269 , n38538 );
and ( n38879 , n38877 , n38878 );
xor ( n38880 , n38877 , n38878 );
xor ( n38881 , n38198 , n38364 );
and ( n38882 , n30274 , n38538 );
and ( n38883 , n38881 , n38882 );
xor ( n38884 , n38881 , n38882 );
xor ( n38885 , n38202 , n38362 );
and ( n38886 , n30279 , n38538 );
and ( n38887 , n38885 , n38886 );
xor ( n38888 , n38885 , n38886 );
xor ( n38889 , n38206 , n38360 );
and ( n38890 , n30284 , n38538 );
and ( n38891 , n38889 , n38890 );
xor ( n38892 , n38889 , n38890 );
xor ( n38893 , n38210 , n38358 );
and ( n38894 , n30289 , n38538 );
and ( n38895 , n38893 , n38894 );
xor ( n38896 , n38893 , n38894 );
xor ( n38897 , n38214 , n38356 );
and ( n38898 , n30294 , n38538 );
and ( n38899 , n38897 , n38898 );
xor ( n38900 , n38897 , n38898 );
xor ( n38901 , n38218 , n38354 );
and ( n38902 , n30299 , n38538 );
and ( n38903 , n38901 , n38902 );
xor ( n38904 , n38901 , n38902 );
xor ( n38905 , n38222 , n38352 );
and ( n38906 , n30304 , n38538 );
and ( n38907 , n38905 , n38906 );
xor ( n38908 , n38905 , n38906 );
xor ( n38909 , n38226 , n38350 );
and ( n38910 , n30309 , n38538 );
and ( n38911 , n38909 , n38910 );
xor ( n38912 , n38909 , n38910 );
xor ( n38913 , n38230 , n38348 );
and ( n38914 , n30314 , n38538 );
and ( n38915 , n38913 , n38914 );
xor ( n38916 , n38913 , n38914 );
xor ( n38917 , n38234 , n38346 );
and ( n38918 , n30319 , n38538 );
and ( n38919 , n38917 , n38918 );
xor ( n38920 , n38917 , n38918 );
xor ( n38921 , n38238 , n38344 );
and ( n38922 , n30324 , n38538 );
and ( n38923 , n38921 , n38922 );
xor ( n38924 , n38921 , n38922 );
xor ( n38925 , n38242 , n38342 );
and ( n38926 , n30329 , n38538 );
and ( n38927 , n38925 , n38926 );
xor ( n38928 , n38925 , n38926 );
xor ( n38929 , n38246 , n38340 );
and ( n38930 , n30334 , n38538 );
and ( n38931 , n38929 , n38930 );
xor ( n38932 , n38929 , n38930 );
xor ( n38933 , n38250 , n38338 );
and ( n38934 , n30339 , n38538 );
and ( n38935 , n38933 , n38934 );
xor ( n38936 , n38933 , n38934 );
xor ( n38937 , n38254 , n38336 );
and ( n38938 , n30344 , n38538 );
and ( n38939 , n38937 , n38938 );
xor ( n38940 , n38937 , n38938 );
xor ( n38941 , n38258 , n38334 );
and ( n38942 , n30349 , n38538 );
and ( n38943 , n38941 , n38942 );
xor ( n38944 , n38941 , n38942 );
xor ( n38945 , n38262 , n38332 );
and ( n38946 , n30354 , n38538 );
and ( n38947 , n38945 , n38946 );
xor ( n38948 , n38945 , n38946 );
xor ( n38949 , n38266 , n38330 );
and ( n38950 , n30359 , n38538 );
and ( n38951 , n38949 , n38950 );
xor ( n38952 , n38949 , n38950 );
xor ( n38953 , n38270 , n38328 );
and ( n38954 , n30364 , n38538 );
and ( n38955 , n38953 , n38954 );
xor ( n38956 , n38953 , n38954 );
xor ( n38957 , n38274 , n38326 );
and ( n38958 , n30369 , n38538 );
and ( n38959 , n38957 , n38958 );
xor ( n38960 , n38957 , n38958 );
xor ( n38961 , n38278 , n38324 );
and ( n38962 , n30374 , n38538 );
and ( n38963 , n38961 , n38962 );
xor ( n38964 , n38961 , n38962 );
xor ( n38965 , n38282 , n38322 );
and ( n38966 , n30379 , n38538 );
and ( n38967 , n38965 , n38966 );
xor ( n38968 , n38965 , n38966 );
xor ( n38969 , n38286 , n38320 );
and ( n38970 , n30384 , n38538 );
and ( n38971 , n38969 , n38970 );
xor ( n38972 , n38969 , n38970 );
xor ( n38973 , n38290 , n38318 );
and ( n38974 , n30389 , n38538 );
and ( n38975 , n38973 , n38974 );
xor ( n38976 , n38973 , n38974 );
xor ( n38977 , n38294 , n38316 );
and ( n38978 , n30394 , n38538 );
and ( n38979 , n38977 , n38978 );
xor ( n38980 , n38977 , n38978 );
xor ( n38981 , n38298 , n38314 );
and ( n38982 , n30399 , n38538 );
and ( n38983 , n38981 , n38982 );
xor ( n38984 , n38981 , n38982 );
xor ( n38985 , n38302 , n38312 );
and ( n38986 , n30404 , n38538 );
and ( n38987 , n38985 , n38986 );
xor ( n38988 , n38985 , n38986 );
xor ( n38989 , n38306 , n38310 );
and ( n38990 , n30409 , n38538 );
and ( n38991 , n38989 , n38990 );
buf ( n38992 , n38991 );
and ( n38993 , n38988 , n38992 );
or ( n38994 , n38987 , n38993 );
and ( n38995 , n38984 , n38994 );
or ( n38996 , n38983 , n38995 );
and ( n38997 , n38980 , n38996 );
or ( n38998 , n38979 , n38997 );
and ( n38999 , n38976 , n38998 );
or ( n39000 , n38975 , n38999 );
and ( n39001 , n38972 , n39000 );
or ( n39002 , n38971 , n39001 );
and ( n39003 , n38968 , n39002 );
or ( n39004 , n38967 , n39003 );
and ( n39005 , n38964 , n39004 );
or ( n39006 , n38963 , n39005 );
and ( n39007 , n38960 , n39006 );
or ( n39008 , n38959 , n39007 );
and ( n39009 , n38956 , n39008 );
or ( n39010 , n38955 , n39009 );
and ( n39011 , n38952 , n39010 );
or ( n39012 , n38951 , n39011 );
and ( n39013 , n38948 , n39012 );
or ( n39014 , n38947 , n39013 );
and ( n39015 , n38944 , n39014 );
or ( n39016 , n38943 , n39015 );
and ( n39017 , n38940 , n39016 );
or ( n39018 , n38939 , n39017 );
and ( n39019 , n38936 , n39018 );
or ( n39020 , n38935 , n39019 );
and ( n39021 , n38932 , n39020 );
or ( n39022 , n38931 , n39021 );
and ( n39023 , n38928 , n39022 );
or ( n39024 , n38927 , n39023 );
and ( n39025 , n38924 , n39024 );
or ( n39026 , n38923 , n39025 );
and ( n39027 , n38920 , n39026 );
or ( n39028 , n38919 , n39027 );
and ( n39029 , n38916 , n39028 );
or ( n39030 , n38915 , n39029 );
and ( n39031 , n38912 , n39030 );
or ( n39032 , n38911 , n39031 );
and ( n39033 , n38908 , n39032 );
or ( n39034 , n38907 , n39033 );
and ( n39035 , n38904 , n39034 );
or ( n39036 , n38903 , n39035 );
and ( n39037 , n38900 , n39036 );
or ( n39038 , n38899 , n39037 );
and ( n39039 , n38896 , n39038 );
or ( n39040 , n38895 , n39039 );
and ( n39041 , n38892 , n39040 );
or ( n39042 , n38891 , n39041 );
and ( n39043 , n38888 , n39042 );
or ( n39044 , n38887 , n39043 );
and ( n39045 , n38884 , n39044 );
or ( n39046 , n38883 , n39045 );
and ( n39047 , n38880 , n39046 );
or ( n39048 , n38879 , n39047 );
and ( n39049 , n38876 , n39048 );
or ( n39050 , n38875 , n39049 );
and ( n39051 , n38872 , n39050 );
or ( n39052 , n38871 , n39051 );
and ( n39053 , n38868 , n39052 );
or ( n39054 , n38867 , n39053 );
and ( n39055 , n38864 , n39054 );
or ( n39056 , n38863 , n39055 );
and ( n39057 , n38860 , n39056 );
or ( n39058 , n38859 , n39057 );
and ( n39059 , n38856 , n39058 );
or ( n39060 , n38855 , n39059 );
and ( n39061 , n38852 , n39060 );
or ( n39062 , n38851 , n39061 );
and ( n39063 , n38848 , n39062 );
or ( n39064 , n38847 , n39063 );
and ( n39065 , n38844 , n39064 );
or ( n39066 , n38843 , n39065 );
and ( n39067 , n38840 , n39066 );
or ( n39068 , n38839 , n39067 );
and ( n39069 , n38836 , n39068 );
or ( n39070 , n38835 , n39069 );
and ( n39071 , n38832 , n39070 );
or ( n39072 , n38831 , n39071 );
and ( n39073 , n38828 , n39072 );
or ( n39074 , n38827 , n39073 );
and ( n39075 , n38824 , n39074 );
or ( n39076 , n38823 , n39075 );
and ( n39077 , n38820 , n39076 );
or ( n39078 , n38819 , n39077 );
and ( n39079 , n38816 , n39078 );
or ( n39080 , n38815 , n39079 );
and ( n39081 , n38812 , n39080 );
or ( n39082 , n38811 , n39081 );
and ( n39083 , n38808 , n39082 );
or ( n39084 , n38807 , n39083 );
and ( n39085 , n38804 , n39084 );
or ( n39086 , n38803 , n39085 );
and ( n39087 , n38800 , n39086 );
or ( n39088 , n38799 , n39087 );
and ( n39089 , n38796 , n39088 );
or ( n39090 , n38795 , n39089 );
and ( n39091 , n38792 , n39090 );
or ( n39092 , n38791 , n39091 );
and ( n39093 , n38788 , n39092 );
or ( n39094 , n38787 , n39093 );
and ( n39095 , n38784 , n39094 );
or ( n39096 , n38783 , n39095 );
and ( n39097 , n38780 , n39096 );
or ( n39098 , n38779 , n39097 );
and ( n39099 , n38776 , n39098 );
or ( n39100 , n38775 , n39099 );
and ( n39101 , n38772 , n39100 );
or ( n39102 , n38771 , n39101 );
and ( n39103 , n38768 , n39102 );
or ( n39104 , n38767 , n39103 );
and ( n39105 , n38764 , n39104 );
or ( n39106 , n38763 , n39105 );
and ( n39107 , n38760 , n39106 );
or ( n39108 , n38759 , n39107 );
and ( n39109 , n38756 , n39108 );
or ( n39110 , n38755 , n39109 );
and ( n39111 , n38752 , n39110 );
or ( n39112 , n38751 , n39111 );
and ( n39113 , n38748 , n39112 );
or ( n39114 , n38747 , n39113 );
and ( n39115 , n38744 , n39114 );
or ( n39116 , n38743 , n39115 );
and ( n39117 , n38740 , n39116 );
or ( n39118 , n38739 , n39117 );
and ( n39119 , n38736 , n39118 );
or ( n39120 , n38735 , n39119 );
and ( n39121 , n38732 , n39120 );
or ( n39122 , n38731 , n39121 );
and ( n39123 , n38728 , n39122 );
or ( n39124 , n38727 , n39123 );
and ( n39125 , n38724 , n39124 );
or ( n39126 , n38723 , n39125 );
and ( n39127 , n38720 , n39126 );
or ( n39128 , n38719 , n39127 );
and ( n39129 , n38716 , n39128 );
or ( n39130 , n38715 , n39129 );
and ( n39131 , n38712 , n39130 );
or ( n39132 , n38711 , n39131 );
and ( n39133 , n38708 , n39132 );
or ( n39134 , n38707 , n39133 );
and ( n39135 , n38704 , n39134 );
or ( n39136 , n38703 , n39135 );
and ( n39137 , n38700 , n39136 );
or ( n39138 , n38699 , n39137 );
and ( n39139 , n38696 , n39138 );
or ( n39140 , n38695 , n39139 );
and ( n39141 , n38692 , n39140 );
or ( n39142 , n38691 , n39141 );
and ( n39143 , n38688 , n39142 );
or ( n39144 , n38687 , n39143 );
and ( n39145 , n38684 , n39144 );
or ( n39146 , n38683 , n39145 );
and ( n39147 , n38680 , n39146 );
or ( n39148 , n38679 , n39147 );
and ( n39149 , n38676 , n39148 );
or ( n39150 , n38675 , n39149 );
and ( n39151 , n38672 , n39150 );
or ( n39152 , n38671 , n39151 );
and ( n39153 , n38668 , n39152 );
or ( n39154 , n38667 , n39153 );
and ( n39155 , n38664 , n39154 );
or ( n39156 , n38663 , n39155 );
and ( n39157 , n38660 , n39156 );
or ( n39158 , n38659 , n39157 );
and ( n39159 , n38656 , n39158 );
or ( n39160 , n38655 , n39159 );
and ( n39161 , n38652 , n39160 );
or ( n39162 , n38651 , n39161 );
and ( n39163 , n38648 , n39162 );
or ( n39164 , n38647 , n39163 );
and ( n39165 , n38644 , n39164 );
or ( n39166 , n38643 , n39165 );
and ( n39167 , n38640 , n39166 );
or ( n39168 , n38639 , n39167 );
and ( n39169 , n38636 , n39168 );
or ( n39170 , n38635 , n39169 );
and ( n39171 , n38632 , n39170 );
or ( n39172 , n38631 , n39171 );
and ( n39173 , n38628 , n39172 );
or ( n39174 , n38627 , n39173 );
and ( n39175 , n38624 , n39174 );
or ( n39176 , n38623 , n39175 );
and ( n39177 , n38620 , n39176 );
or ( n39178 , n38619 , n39177 );
and ( n39179 , n38616 , n39178 );
or ( n39180 , n38615 , n39179 );
and ( n39181 , n38612 , n39180 );
or ( n39182 , n38611 , n39181 );
and ( n39183 , n38608 , n39182 );
or ( n39184 , n38607 , n39183 );
and ( n39185 , n38604 , n39184 );
or ( n39186 , n38603 , n39185 );
and ( n39187 , n38600 , n39186 );
or ( n39188 , n38599 , n39187 );
and ( n39189 , n38596 , n39188 );
or ( n39190 , n38595 , n39189 );
and ( n39191 , n38592 , n39190 );
or ( n39192 , n38591 , n39191 );
and ( n39193 , n38588 , n39192 );
or ( n39194 , n38587 , n39193 );
and ( n39195 , n38584 , n39194 );
or ( n39196 , n38583 , n39195 );
and ( n39197 , n38580 , n39196 );
or ( n39198 , n38579 , n39197 );
and ( n39199 , n38576 , n39198 );
or ( n39200 , n38575 , n39199 );
and ( n39201 , n38572 , n39200 );
or ( n39202 , n38571 , n39201 );
and ( n39203 , n38568 , n39202 );
or ( n39204 , n38567 , n39203 );
and ( n39205 , n38564 , n39204 );
or ( n39206 , n38563 , n39205 );
and ( n39207 , n38560 , n39206 );
or ( n39208 , n38559 , n39207 );
and ( n39209 , n38556 , n39208 );
or ( n39210 , n38555 , n39209 );
and ( n39211 , n38552 , n39210 );
or ( n39212 , n38551 , n39211 );
and ( n39213 , n38548 , n39212 );
or ( n39214 , n38547 , n39213 );
and ( n39215 , n38544 , n39214 );
or ( n39216 , n38543 , n39215 );
xor ( n39217 , n38540 , n39216 );
buf ( n39218 , n18078 );
and ( n39219 , n29849 , n39218 );
xor ( n39220 , n39217 , n39219 );
xor ( n39221 , n38544 , n39214 );
and ( n39222 , n29854 , n39218 );
and ( n39223 , n39221 , n39222 );
xor ( n39224 , n39221 , n39222 );
xor ( n39225 , n38548 , n39212 );
and ( n39226 , n29859 , n39218 );
and ( n39227 , n39225 , n39226 );
xor ( n39228 , n39225 , n39226 );
xor ( n39229 , n38552 , n39210 );
and ( n39230 , n29864 , n39218 );
and ( n39231 , n39229 , n39230 );
xor ( n39232 , n39229 , n39230 );
xor ( n39233 , n38556 , n39208 );
and ( n39234 , n29869 , n39218 );
and ( n39235 , n39233 , n39234 );
xor ( n39236 , n39233 , n39234 );
xor ( n39237 , n38560 , n39206 );
and ( n39238 , n29874 , n39218 );
and ( n39239 , n39237 , n39238 );
xor ( n39240 , n39237 , n39238 );
xor ( n39241 , n38564 , n39204 );
and ( n39242 , n29879 , n39218 );
and ( n39243 , n39241 , n39242 );
xor ( n39244 , n39241 , n39242 );
xor ( n39245 , n38568 , n39202 );
and ( n39246 , n29884 , n39218 );
and ( n39247 , n39245 , n39246 );
xor ( n39248 , n39245 , n39246 );
xor ( n39249 , n38572 , n39200 );
and ( n39250 , n29889 , n39218 );
and ( n39251 , n39249 , n39250 );
xor ( n39252 , n39249 , n39250 );
xor ( n39253 , n38576 , n39198 );
and ( n39254 , n29894 , n39218 );
and ( n39255 , n39253 , n39254 );
xor ( n39256 , n39253 , n39254 );
xor ( n39257 , n38580 , n39196 );
and ( n39258 , n29899 , n39218 );
and ( n39259 , n39257 , n39258 );
xor ( n39260 , n39257 , n39258 );
xor ( n39261 , n38584 , n39194 );
and ( n39262 , n29904 , n39218 );
and ( n39263 , n39261 , n39262 );
xor ( n39264 , n39261 , n39262 );
xor ( n39265 , n38588 , n39192 );
and ( n39266 , n29909 , n39218 );
and ( n39267 , n39265 , n39266 );
xor ( n39268 , n39265 , n39266 );
xor ( n39269 , n38592 , n39190 );
and ( n39270 , n29914 , n39218 );
and ( n39271 , n39269 , n39270 );
xor ( n39272 , n39269 , n39270 );
xor ( n39273 , n38596 , n39188 );
and ( n39274 , n29919 , n39218 );
and ( n39275 , n39273 , n39274 );
xor ( n39276 , n39273 , n39274 );
xor ( n39277 , n38600 , n39186 );
and ( n39278 , n29924 , n39218 );
and ( n39279 , n39277 , n39278 );
xor ( n39280 , n39277 , n39278 );
xor ( n39281 , n38604 , n39184 );
and ( n39282 , n29929 , n39218 );
and ( n39283 , n39281 , n39282 );
xor ( n39284 , n39281 , n39282 );
xor ( n39285 , n38608 , n39182 );
and ( n39286 , n29934 , n39218 );
and ( n39287 , n39285 , n39286 );
xor ( n39288 , n39285 , n39286 );
xor ( n39289 , n38612 , n39180 );
and ( n39290 , n29939 , n39218 );
and ( n39291 , n39289 , n39290 );
xor ( n39292 , n39289 , n39290 );
xor ( n39293 , n38616 , n39178 );
and ( n39294 , n29944 , n39218 );
and ( n39295 , n39293 , n39294 );
xor ( n39296 , n39293 , n39294 );
xor ( n39297 , n38620 , n39176 );
and ( n39298 , n29949 , n39218 );
and ( n39299 , n39297 , n39298 );
xor ( n39300 , n39297 , n39298 );
xor ( n39301 , n38624 , n39174 );
and ( n39302 , n29954 , n39218 );
and ( n39303 , n39301 , n39302 );
xor ( n39304 , n39301 , n39302 );
xor ( n39305 , n38628 , n39172 );
and ( n39306 , n29959 , n39218 );
and ( n39307 , n39305 , n39306 );
xor ( n39308 , n39305 , n39306 );
xor ( n39309 , n38632 , n39170 );
and ( n39310 , n29964 , n39218 );
and ( n39311 , n39309 , n39310 );
xor ( n39312 , n39309 , n39310 );
xor ( n39313 , n38636 , n39168 );
and ( n39314 , n29969 , n39218 );
and ( n39315 , n39313 , n39314 );
xor ( n39316 , n39313 , n39314 );
xor ( n39317 , n38640 , n39166 );
and ( n39318 , n29974 , n39218 );
and ( n39319 , n39317 , n39318 );
xor ( n39320 , n39317 , n39318 );
xor ( n39321 , n38644 , n39164 );
and ( n39322 , n29979 , n39218 );
and ( n39323 , n39321 , n39322 );
xor ( n39324 , n39321 , n39322 );
xor ( n39325 , n38648 , n39162 );
and ( n39326 , n29984 , n39218 );
and ( n39327 , n39325 , n39326 );
xor ( n39328 , n39325 , n39326 );
xor ( n39329 , n38652 , n39160 );
and ( n39330 , n29989 , n39218 );
and ( n39331 , n39329 , n39330 );
xor ( n39332 , n39329 , n39330 );
xor ( n39333 , n38656 , n39158 );
and ( n39334 , n29994 , n39218 );
and ( n39335 , n39333 , n39334 );
xor ( n39336 , n39333 , n39334 );
xor ( n39337 , n38660 , n39156 );
and ( n39338 , n29999 , n39218 );
and ( n39339 , n39337 , n39338 );
xor ( n39340 , n39337 , n39338 );
xor ( n39341 , n38664 , n39154 );
and ( n39342 , n30004 , n39218 );
and ( n39343 , n39341 , n39342 );
xor ( n39344 , n39341 , n39342 );
xor ( n39345 , n38668 , n39152 );
and ( n39346 , n30009 , n39218 );
and ( n39347 , n39345 , n39346 );
xor ( n39348 , n39345 , n39346 );
xor ( n39349 , n38672 , n39150 );
and ( n39350 , n30014 , n39218 );
and ( n39351 , n39349 , n39350 );
xor ( n39352 , n39349 , n39350 );
xor ( n39353 , n38676 , n39148 );
and ( n39354 , n30019 , n39218 );
and ( n39355 , n39353 , n39354 );
xor ( n39356 , n39353 , n39354 );
xor ( n39357 , n38680 , n39146 );
and ( n39358 , n30024 , n39218 );
and ( n39359 , n39357 , n39358 );
xor ( n39360 , n39357 , n39358 );
xor ( n39361 , n38684 , n39144 );
and ( n39362 , n30029 , n39218 );
and ( n39363 , n39361 , n39362 );
xor ( n39364 , n39361 , n39362 );
xor ( n39365 , n38688 , n39142 );
and ( n39366 , n30034 , n39218 );
and ( n39367 , n39365 , n39366 );
xor ( n39368 , n39365 , n39366 );
xor ( n39369 , n38692 , n39140 );
and ( n39370 , n30039 , n39218 );
and ( n39371 , n39369 , n39370 );
xor ( n39372 , n39369 , n39370 );
xor ( n39373 , n38696 , n39138 );
and ( n39374 , n30044 , n39218 );
and ( n39375 , n39373 , n39374 );
xor ( n39376 , n39373 , n39374 );
xor ( n39377 , n38700 , n39136 );
and ( n39378 , n30049 , n39218 );
and ( n39379 , n39377 , n39378 );
xor ( n39380 , n39377 , n39378 );
xor ( n39381 , n38704 , n39134 );
and ( n39382 , n30054 , n39218 );
and ( n39383 , n39381 , n39382 );
xor ( n39384 , n39381 , n39382 );
xor ( n39385 , n38708 , n39132 );
and ( n39386 , n30059 , n39218 );
and ( n39387 , n39385 , n39386 );
xor ( n39388 , n39385 , n39386 );
xor ( n39389 , n38712 , n39130 );
and ( n39390 , n30064 , n39218 );
and ( n39391 , n39389 , n39390 );
xor ( n39392 , n39389 , n39390 );
xor ( n39393 , n38716 , n39128 );
and ( n39394 , n30069 , n39218 );
and ( n39395 , n39393 , n39394 );
xor ( n39396 , n39393 , n39394 );
xor ( n39397 , n38720 , n39126 );
and ( n39398 , n30074 , n39218 );
and ( n39399 , n39397 , n39398 );
xor ( n39400 , n39397 , n39398 );
xor ( n39401 , n38724 , n39124 );
and ( n39402 , n30079 , n39218 );
and ( n39403 , n39401 , n39402 );
xor ( n39404 , n39401 , n39402 );
xor ( n39405 , n38728 , n39122 );
and ( n39406 , n30084 , n39218 );
and ( n39407 , n39405 , n39406 );
xor ( n39408 , n39405 , n39406 );
xor ( n39409 , n38732 , n39120 );
and ( n39410 , n30089 , n39218 );
and ( n39411 , n39409 , n39410 );
xor ( n39412 , n39409 , n39410 );
xor ( n39413 , n38736 , n39118 );
and ( n39414 , n30094 , n39218 );
and ( n39415 , n39413 , n39414 );
xor ( n39416 , n39413 , n39414 );
xor ( n39417 , n38740 , n39116 );
and ( n39418 , n30099 , n39218 );
and ( n39419 , n39417 , n39418 );
xor ( n39420 , n39417 , n39418 );
xor ( n39421 , n38744 , n39114 );
and ( n39422 , n30104 , n39218 );
and ( n39423 , n39421 , n39422 );
xor ( n39424 , n39421 , n39422 );
xor ( n39425 , n38748 , n39112 );
and ( n39426 , n30109 , n39218 );
and ( n39427 , n39425 , n39426 );
xor ( n39428 , n39425 , n39426 );
xor ( n39429 , n38752 , n39110 );
and ( n39430 , n30114 , n39218 );
and ( n39431 , n39429 , n39430 );
xor ( n39432 , n39429 , n39430 );
xor ( n39433 , n38756 , n39108 );
and ( n39434 , n30119 , n39218 );
and ( n39435 , n39433 , n39434 );
xor ( n39436 , n39433 , n39434 );
xor ( n39437 , n38760 , n39106 );
and ( n39438 , n30124 , n39218 );
and ( n39439 , n39437 , n39438 );
xor ( n39440 , n39437 , n39438 );
xor ( n39441 , n38764 , n39104 );
and ( n39442 , n30129 , n39218 );
and ( n39443 , n39441 , n39442 );
xor ( n39444 , n39441 , n39442 );
xor ( n39445 , n38768 , n39102 );
and ( n39446 , n30134 , n39218 );
and ( n39447 , n39445 , n39446 );
xor ( n39448 , n39445 , n39446 );
xor ( n39449 , n38772 , n39100 );
and ( n39450 , n30139 , n39218 );
and ( n39451 , n39449 , n39450 );
xor ( n39452 , n39449 , n39450 );
xor ( n39453 , n38776 , n39098 );
and ( n39454 , n30144 , n39218 );
and ( n39455 , n39453 , n39454 );
xor ( n39456 , n39453 , n39454 );
xor ( n39457 , n38780 , n39096 );
and ( n39458 , n30149 , n39218 );
and ( n39459 , n39457 , n39458 );
xor ( n39460 , n39457 , n39458 );
xor ( n39461 , n38784 , n39094 );
and ( n39462 , n30154 , n39218 );
and ( n39463 , n39461 , n39462 );
xor ( n39464 , n39461 , n39462 );
xor ( n39465 , n38788 , n39092 );
and ( n39466 , n30159 , n39218 );
and ( n39467 , n39465 , n39466 );
xor ( n39468 , n39465 , n39466 );
xor ( n39469 , n38792 , n39090 );
and ( n39470 , n30164 , n39218 );
and ( n39471 , n39469 , n39470 );
xor ( n39472 , n39469 , n39470 );
xor ( n39473 , n38796 , n39088 );
and ( n39474 , n30169 , n39218 );
and ( n39475 , n39473 , n39474 );
xor ( n39476 , n39473 , n39474 );
xor ( n39477 , n38800 , n39086 );
and ( n39478 , n30174 , n39218 );
and ( n39479 , n39477 , n39478 );
xor ( n39480 , n39477 , n39478 );
xor ( n39481 , n38804 , n39084 );
and ( n39482 , n30179 , n39218 );
and ( n39483 , n39481 , n39482 );
xor ( n39484 , n39481 , n39482 );
xor ( n39485 , n38808 , n39082 );
and ( n39486 , n30184 , n39218 );
and ( n39487 , n39485 , n39486 );
xor ( n39488 , n39485 , n39486 );
xor ( n39489 , n38812 , n39080 );
and ( n39490 , n30189 , n39218 );
and ( n39491 , n39489 , n39490 );
xor ( n39492 , n39489 , n39490 );
xor ( n39493 , n38816 , n39078 );
and ( n39494 , n30194 , n39218 );
and ( n39495 , n39493 , n39494 );
xor ( n39496 , n39493 , n39494 );
xor ( n39497 , n38820 , n39076 );
and ( n39498 , n30199 , n39218 );
and ( n39499 , n39497 , n39498 );
xor ( n39500 , n39497 , n39498 );
xor ( n39501 , n38824 , n39074 );
and ( n39502 , n30204 , n39218 );
and ( n39503 , n39501 , n39502 );
xor ( n39504 , n39501 , n39502 );
xor ( n39505 , n38828 , n39072 );
and ( n39506 , n30209 , n39218 );
and ( n39507 , n39505 , n39506 );
xor ( n39508 , n39505 , n39506 );
xor ( n39509 , n38832 , n39070 );
and ( n39510 , n30214 , n39218 );
and ( n39511 , n39509 , n39510 );
xor ( n39512 , n39509 , n39510 );
xor ( n39513 , n38836 , n39068 );
and ( n39514 , n30219 , n39218 );
and ( n39515 , n39513 , n39514 );
xor ( n39516 , n39513 , n39514 );
xor ( n39517 , n38840 , n39066 );
and ( n39518 , n30224 , n39218 );
and ( n39519 , n39517 , n39518 );
xor ( n39520 , n39517 , n39518 );
xor ( n39521 , n38844 , n39064 );
and ( n39522 , n30229 , n39218 );
and ( n39523 , n39521 , n39522 );
xor ( n39524 , n39521 , n39522 );
xor ( n39525 , n38848 , n39062 );
and ( n39526 , n30234 , n39218 );
and ( n39527 , n39525 , n39526 );
xor ( n39528 , n39525 , n39526 );
xor ( n39529 , n38852 , n39060 );
and ( n39530 , n30239 , n39218 );
and ( n39531 , n39529 , n39530 );
xor ( n39532 , n39529 , n39530 );
xor ( n39533 , n38856 , n39058 );
and ( n39534 , n30244 , n39218 );
and ( n39535 , n39533 , n39534 );
xor ( n39536 , n39533 , n39534 );
xor ( n39537 , n38860 , n39056 );
and ( n39538 , n30249 , n39218 );
and ( n39539 , n39537 , n39538 );
xor ( n39540 , n39537 , n39538 );
xor ( n39541 , n38864 , n39054 );
and ( n39542 , n30254 , n39218 );
and ( n39543 , n39541 , n39542 );
xor ( n39544 , n39541 , n39542 );
xor ( n39545 , n38868 , n39052 );
and ( n39546 , n30259 , n39218 );
and ( n39547 , n39545 , n39546 );
xor ( n39548 , n39545 , n39546 );
xor ( n39549 , n38872 , n39050 );
and ( n39550 , n30264 , n39218 );
and ( n39551 , n39549 , n39550 );
xor ( n39552 , n39549 , n39550 );
xor ( n39553 , n38876 , n39048 );
and ( n39554 , n30269 , n39218 );
and ( n39555 , n39553 , n39554 );
xor ( n39556 , n39553 , n39554 );
xor ( n39557 , n38880 , n39046 );
and ( n39558 , n30274 , n39218 );
and ( n39559 , n39557 , n39558 );
xor ( n39560 , n39557 , n39558 );
xor ( n39561 , n38884 , n39044 );
and ( n39562 , n30279 , n39218 );
and ( n39563 , n39561 , n39562 );
xor ( n39564 , n39561 , n39562 );
xor ( n39565 , n38888 , n39042 );
and ( n39566 , n30284 , n39218 );
and ( n39567 , n39565 , n39566 );
xor ( n39568 , n39565 , n39566 );
xor ( n39569 , n38892 , n39040 );
and ( n39570 , n30289 , n39218 );
and ( n39571 , n39569 , n39570 );
xor ( n39572 , n39569 , n39570 );
xor ( n39573 , n38896 , n39038 );
and ( n39574 , n30294 , n39218 );
and ( n39575 , n39573 , n39574 );
xor ( n39576 , n39573 , n39574 );
xor ( n39577 , n38900 , n39036 );
and ( n39578 , n30299 , n39218 );
and ( n39579 , n39577 , n39578 );
xor ( n39580 , n39577 , n39578 );
xor ( n39581 , n38904 , n39034 );
and ( n39582 , n30304 , n39218 );
and ( n39583 , n39581 , n39582 );
xor ( n39584 , n39581 , n39582 );
xor ( n39585 , n38908 , n39032 );
and ( n39586 , n30309 , n39218 );
and ( n39587 , n39585 , n39586 );
xor ( n39588 , n39585 , n39586 );
xor ( n39589 , n38912 , n39030 );
and ( n39590 , n30314 , n39218 );
and ( n39591 , n39589 , n39590 );
xor ( n39592 , n39589 , n39590 );
xor ( n39593 , n38916 , n39028 );
and ( n39594 , n30319 , n39218 );
and ( n39595 , n39593 , n39594 );
xor ( n39596 , n39593 , n39594 );
xor ( n39597 , n38920 , n39026 );
and ( n39598 , n30324 , n39218 );
and ( n39599 , n39597 , n39598 );
xor ( n39600 , n39597 , n39598 );
xor ( n39601 , n38924 , n39024 );
and ( n39602 , n30329 , n39218 );
and ( n39603 , n39601 , n39602 );
xor ( n39604 , n39601 , n39602 );
xor ( n39605 , n38928 , n39022 );
and ( n39606 , n30334 , n39218 );
and ( n39607 , n39605 , n39606 );
xor ( n39608 , n39605 , n39606 );
xor ( n39609 , n38932 , n39020 );
and ( n39610 , n30339 , n39218 );
and ( n39611 , n39609 , n39610 );
xor ( n39612 , n39609 , n39610 );
xor ( n39613 , n38936 , n39018 );
and ( n39614 , n30344 , n39218 );
and ( n39615 , n39613 , n39614 );
xor ( n39616 , n39613 , n39614 );
xor ( n39617 , n38940 , n39016 );
and ( n39618 , n30349 , n39218 );
and ( n39619 , n39617 , n39618 );
xor ( n39620 , n39617 , n39618 );
xor ( n39621 , n38944 , n39014 );
and ( n39622 , n30354 , n39218 );
and ( n39623 , n39621 , n39622 );
xor ( n39624 , n39621 , n39622 );
xor ( n39625 , n38948 , n39012 );
and ( n39626 , n30359 , n39218 );
and ( n39627 , n39625 , n39626 );
xor ( n39628 , n39625 , n39626 );
xor ( n39629 , n38952 , n39010 );
and ( n39630 , n30364 , n39218 );
and ( n39631 , n39629 , n39630 );
xor ( n39632 , n39629 , n39630 );
xor ( n39633 , n38956 , n39008 );
and ( n39634 , n30369 , n39218 );
and ( n39635 , n39633 , n39634 );
xor ( n39636 , n39633 , n39634 );
xor ( n39637 , n38960 , n39006 );
and ( n39638 , n30374 , n39218 );
and ( n39639 , n39637 , n39638 );
xor ( n39640 , n39637 , n39638 );
xor ( n39641 , n38964 , n39004 );
and ( n39642 , n30379 , n39218 );
and ( n39643 , n39641 , n39642 );
xor ( n39644 , n39641 , n39642 );
xor ( n39645 , n38968 , n39002 );
and ( n39646 , n30384 , n39218 );
and ( n39647 , n39645 , n39646 );
xor ( n39648 , n39645 , n39646 );
xor ( n39649 , n38972 , n39000 );
and ( n39650 , n30389 , n39218 );
and ( n39651 , n39649 , n39650 );
xor ( n39652 , n39649 , n39650 );
xor ( n39653 , n38976 , n38998 );
and ( n39654 , n30394 , n39218 );
and ( n39655 , n39653 , n39654 );
xor ( n39656 , n39653 , n39654 );
xor ( n39657 , n38980 , n38996 );
and ( n39658 , n30399 , n39218 );
and ( n39659 , n39657 , n39658 );
xor ( n39660 , n39657 , n39658 );
xor ( n39661 , n38984 , n38994 );
and ( n39662 , n30404 , n39218 );
and ( n39663 , n39661 , n39662 );
xor ( n39664 , n39661 , n39662 );
xor ( n39665 , n38988 , n38992 );
and ( n39666 , n30409 , n39218 );
and ( n39667 , n39665 , n39666 );
buf ( n39668 , n39667 );
and ( n39669 , n39664 , n39668 );
or ( n39670 , n39663 , n39669 );
and ( n39671 , n39660 , n39670 );
or ( n39672 , n39659 , n39671 );
and ( n39673 , n39656 , n39672 );
or ( n39674 , n39655 , n39673 );
and ( n39675 , n39652 , n39674 );
or ( n39676 , n39651 , n39675 );
and ( n39677 , n39648 , n39676 );
or ( n39678 , n39647 , n39677 );
and ( n39679 , n39644 , n39678 );
or ( n39680 , n39643 , n39679 );
and ( n39681 , n39640 , n39680 );
or ( n39682 , n39639 , n39681 );
and ( n39683 , n39636 , n39682 );
or ( n39684 , n39635 , n39683 );
and ( n39685 , n39632 , n39684 );
or ( n39686 , n39631 , n39685 );
and ( n39687 , n39628 , n39686 );
or ( n39688 , n39627 , n39687 );
and ( n39689 , n39624 , n39688 );
or ( n39690 , n39623 , n39689 );
and ( n39691 , n39620 , n39690 );
or ( n39692 , n39619 , n39691 );
and ( n39693 , n39616 , n39692 );
or ( n39694 , n39615 , n39693 );
and ( n39695 , n39612 , n39694 );
or ( n39696 , n39611 , n39695 );
and ( n39697 , n39608 , n39696 );
or ( n39698 , n39607 , n39697 );
and ( n39699 , n39604 , n39698 );
or ( n39700 , n39603 , n39699 );
and ( n39701 , n39600 , n39700 );
or ( n39702 , n39599 , n39701 );
and ( n39703 , n39596 , n39702 );
or ( n39704 , n39595 , n39703 );
and ( n39705 , n39592 , n39704 );
or ( n39706 , n39591 , n39705 );
and ( n39707 , n39588 , n39706 );
or ( n39708 , n39587 , n39707 );
and ( n39709 , n39584 , n39708 );
or ( n39710 , n39583 , n39709 );
and ( n39711 , n39580 , n39710 );
or ( n39712 , n39579 , n39711 );
and ( n39713 , n39576 , n39712 );
or ( n39714 , n39575 , n39713 );
and ( n39715 , n39572 , n39714 );
or ( n39716 , n39571 , n39715 );
and ( n39717 , n39568 , n39716 );
or ( n39718 , n39567 , n39717 );
and ( n39719 , n39564 , n39718 );
or ( n39720 , n39563 , n39719 );
and ( n39721 , n39560 , n39720 );
or ( n39722 , n39559 , n39721 );
and ( n39723 , n39556 , n39722 );
or ( n39724 , n39555 , n39723 );
and ( n39725 , n39552 , n39724 );
or ( n39726 , n39551 , n39725 );
and ( n39727 , n39548 , n39726 );
or ( n39728 , n39547 , n39727 );
and ( n39729 , n39544 , n39728 );
or ( n39730 , n39543 , n39729 );
and ( n39731 , n39540 , n39730 );
or ( n39732 , n39539 , n39731 );
and ( n39733 , n39536 , n39732 );
or ( n39734 , n39535 , n39733 );
and ( n39735 , n39532 , n39734 );
or ( n39736 , n39531 , n39735 );
and ( n39737 , n39528 , n39736 );
or ( n39738 , n39527 , n39737 );
and ( n39739 , n39524 , n39738 );
or ( n39740 , n39523 , n39739 );
and ( n39741 , n39520 , n39740 );
or ( n39742 , n39519 , n39741 );
and ( n39743 , n39516 , n39742 );
or ( n39744 , n39515 , n39743 );
and ( n39745 , n39512 , n39744 );
or ( n39746 , n39511 , n39745 );
and ( n39747 , n39508 , n39746 );
or ( n39748 , n39507 , n39747 );
and ( n39749 , n39504 , n39748 );
or ( n39750 , n39503 , n39749 );
and ( n39751 , n39500 , n39750 );
or ( n39752 , n39499 , n39751 );
and ( n39753 , n39496 , n39752 );
or ( n39754 , n39495 , n39753 );
and ( n39755 , n39492 , n39754 );
or ( n39756 , n39491 , n39755 );
and ( n39757 , n39488 , n39756 );
or ( n39758 , n39487 , n39757 );
and ( n39759 , n39484 , n39758 );
or ( n39760 , n39483 , n39759 );
and ( n39761 , n39480 , n39760 );
or ( n39762 , n39479 , n39761 );
and ( n39763 , n39476 , n39762 );
or ( n39764 , n39475 , n39763 );
and ( n39765 , n39472 , n39764 );
or ( n39766 , n39471 , n39765 );
and ( n39767 , n39468 , n39766 );
or ( n39768 , n39467 , n39767 );
and ( n39769 , n39464 , n39768 );
or ( n39770 , n39463 , n39769 );
and ( n39771 , n39460 , n39770 );
or ( n39772 , n39459 , n39771 );
and ( n39773 , n39456 , n39772 );
or ( n39774 , n39455 , n39773 );
and ( n39775 , n39452 , n39774 );
or ( n39776 , n39451 , n39775 );
and ( n39777 , n39448 , n39776 );
or ( n39778 , n39447 , n39777 );
and ( n39779 , n39444 , n39778 );
or ( n39780 , n39443 , n39779 );
and ( n39781 , n39440 , n39780 );
or ( n39782 , n39439 , n39781 );
and ( n39783 , n39436 , n39782 );
or ( n39784 , n39435 , n39783 );
and ( n39785 , n39432 , n39784 );
or ( n39786 , n39431 , n39785 );
and ( n39787 , n39428 , n39786 );
or ( n39788 , n39427 , n39787 );
and ( n39789 , n39424 , n39788 );
or ( n39790 , n39423 , n39789 );
and ( n39791 , n39420 , n39790 );
or ( n39792 , n39419 , n39791 );
and ( n39793 , n39416 , n39792 );
or ( n39794 , n39415 , n39793 );
and ( n39795 , n39412 , n39794 );
or ( n39796 , n39411 , n39795 );
and ( n39797 , n39408 , n39796 );
or ( n39798 , n39407 , n39797 );
and ( n39799 , n39404 , n39798 );
or ( n39800 , n39403 , n39799 );
and ( n39801 , n39400 , n39800 );
or ( n39802 , n39399 , n39801 );
and ( n39803 , n39396 , n39802 );
or ( n39804 , n39395 , n39803 );
and ( n39805 , n39392 , n39804 );
or ( n39806 , n39391 , n39805 );
and ( n39807 , n39388 , n39806 );
or ( n39808 , n39387 , n39807 );
and ( n39809 , n39384 , n39808 );
or ( n39810 , n39383 , n39809 );
and ( n39811 , n39380 , n39810 );
or ( n39812 , n39379 , n39811 );
and ( n39813 , n39376 , n39812 );
or ( n39814 , n39375 , n39813 );
and ( n39815 , n39372 , n39814 );
or ( n39816 , n39371 , n39815 );
and ( n39817 , n39368 , n39816 );
or ( n39818 , n39367 , n39817 );
and ( n39819 , n39364 , n39818 );
or ( n39820 , n39363 , n39819 );
and ( n39821 , n39360 , n39820 );
or ( n39822 , n39359 , n39821 );
and ( n39823 , n39356 , n39822 );
or ( n39824 , n39355 , n39823 );
and ( n39825 , n39352 , n39824 );
or ( n39826 , n39351 , n39825 );
and ( n39827 , n39348 , n39826 );
or ( n39828 , n39347 , n39827 );
and ( n39829 , n39344 , n39828 );
or ( n39830 , n39343 , n39829 );
and ( n39831 , n39340 , n39830 );
or ( n39832 , n39339 , n39831 );
and ( n39833 , n39336 , n39832 );
or ( n39834 , n39335 , n39833 );
and ( n39835 , n39332 , n39834 );
or ( n39836 , n39331 , n39835 );
and ( n39837 , n39328 , n39836 );
or ( n39838 , n39327 , n39837 );
and ( n39839 , n39324 , n39838 );
or ( n39840 , n39323 , n39839 );
and ( n39841 , n39320 , n39840 );
or ( n39842 , n39319 , n39841 );
and ( n39843 , n39316 , n39842 );
or ( n39844 , n39315 , n39843 );
and ( n39845 , n39312 , n39844 );
or ( n39846 , n39311 , n39845 );
and ( n39847 , n39308 , n39846 );
or ( n39848 , n39307 , n39847 );
and ( n39849 , n39304 , n39848 );
or ( n39850 , n39303 , n39849 );
and ( n39851 , n39300 , n39850 );
or ( n39852 , n39299 , n39851 );
and ( n39853 , n39296 , n39852 );
or ( n39854 , n39295 , n39853 );
and ( n39855 , n39292 , n39854 );
or ( n39856 , n39291 , n39855 );
and ( n39857 , n39288 , n39856 );
or ( n39858 , n39287 , n39857 );
and ( n39859 , n39284 , n39858 );
or ( n39860 , n39283 , n39859 );
and ( n39861 , n39280 , n39860 );
or ( n39862 , n39279 , n39861 );
and ( n39863 , n39276 , n39862 );
or ( n39864 , n39275 , n39863 );
and ( n39865 , n39272 , n39864 );
or ( n39866 , n39271 , n39865 );
and ( n39867 , n39268 , n39866 );
or ( n39868 , n39267 , n39867 );
and ( n39869 , n39264 , n39868 );
or ( n39870 , n39263 , n39869 );
and ( n39871 , n39260 , n39870 );
or ( n39872 , n39259 , n39871 );
and ( n39873 , n39256 , n39872 );
or ( n39874 , n39255 , n39873 );
and ( n39875 , n39252 , n39874 );
or ( n39876 , n39251 , n39875 );
and ( n39877 , n39248 , n39876 );
or ( n39878 , n39247 , n39877 );
and ( n39879 , n39244 , n39878 );
or ( n39880 , n39243 , n39879 );
and ( n39881 , n39240 , n39880 );
or ( n39882 , n39239 , n39881 );
and ( n39883 , n39236 , n39882 );
or ( n39884 , n39235 , n39883 );
and ( n39885 , n39232 , n39884 );
or ( n39886 , n39231 , n39885 );
and ( n39887 , n39228 , n39886 );
or ( n39888 , n39227 , n39887 );
and ( n39889 , n39224 , n39888 );
or ( n39890 , n39223 , n39889 );
xor ( n39891 , n39220 , n39890 );
buf ( n39892 , n18076 );
and ( n39893 , n29854 , n39892 );
xor ( n39894 , n39891 , n39893 );
xor ( n39895 , n39224 , n39888 );
and ( n39896 , n29859 , n39892 );
and ( n39897 , n39895 , n39896 );
xor ( n39898 , n39895 , n39896 );
xor ( n39899 , n39228 , n39886 );
and ( n39900 , n29864 , n39892 );
and ( n39901 , n39899 , n39900 );
xor ( n39902 , n39899 , n39900 );
xor ( n39903 , n39232 , n39884 );
and ( n39904 , n29869 , n39892 );
and ( n39905 , n39903 , n39904 );
xor ( n39906 , n39903 , n39904 );
xor ( n39907 , n39236 , n39882 );
and ( n39908 , n29874 , n39892 );
and ( n39909 , n39907 , n39908 );
xor ( n39910 , n39907 , n39908 );
xor ( n39911 , n39240 , n39880 );
and ( n39912 , n29879 , n39892 );
and ( n39913 , n39911 , n39912 );
xor ( n39914 , n39911 , n39912 );
xor ( n39915 , n39244 , n39878 );
and ( n39916 , n29884 , n39892 );
and ( n39917 , n39915 , n39916 );
xor ( n39918 , n39915 , n39916 );
xor ( n39919 , n39248 , n39876 );
and ( n39920 , n29889 , n39892 );
and ( n39921 , n39919 , n39920 );
xor ( n39922 , n39919 , n39920 );
xor ( n39923 , n39252 , n39874 );
and ( n39924 , n29894 , n39892 );
and ( n39925 , n39923 , n39924 );
xor ( n39926 , n39923 , n39924 );
xor ( n39927 , n39256 , n39872 );
and ( n39928 , n29899 , n39892 );
and ( n39929 , n39927 , n39928 );
xor ( n39930 , n39927 , n39928 );
xor ( n39931 , n39260 , n39870 );
and ( n39932 , n29904 , n39892 );
and ( n39933 , n39931 , n39932 );
xor ( n39934 , n39931 , n39932 );
xor ( n39935 , n39264 , n39868 );
and ( n39936 , n29909 , n39892 );
and ( n39937 , n39935 , n39936 );
xor ( n39938 , n39935 , n39936 );
xor ( n39939 , n39268 , n39866 );
and ( n39940 , n29914 , n39892 );
and ( n39941 , n39939 , n39940 );
xor ( n39942 , n39939 , n39940 );
xor ( n39943 , n39272 , n39864 );
and ( n39944 , n29919 , n39892 );
and ( n39945 , n39943 , n39944 );
xor ( n39946 , n39943 , n39944 );
xor ( n39947 , n39276 , n39862 );
and ( n39948 , n29924 , n39892 );
and ( n39949 , n39947 , n39948 );
xor ( n39950 , n39947 , n39948 );
xor ( n39951 , n39280 , n39860 );
and ( n39952 , n29929 , n39892 );
and ( n39953 , n39951 , n39952 );
xor ( n39954 , n39951 , n39952 );
xor ( n39955 , n39284 , n39858 );
and ( n39956 , n29934 , n39892 );
and ( n39957 , n39955 , n39956 );
xor ( n39958 , n39955 , n39956 );
xor ( n39959 , n39288 , n39856 );
and ( n39960 , n29939 , n39892 );
and ( n39961 , n39959 , n39960 );
xor ( n39962 , n39959 , n39960 );
xor ( n39963 , n39292 , n39854 );
and ( n39964 , n29944 , n39892 );
and ( n39965 , n39963 , n39964 );
xor ( n39966 , n39963 , n39964 );
xor ( n39967 , n39296 , n39852 );
and ( n39968 , n29949 , n39892 );
and ( n39969 , n39967 , n39968 );
xor ( n39970 , n39967 , n39968 );
xor ( n39971 , n39300 , n39850 );
and ( n39972 , n29954 , n39892 );
and ( n39973 , n39971 , n39972 );
xor ( n39974 , n39971 , n39972 );
xor ( n39975 , n39304 , n39848 );
and ( n39976 , n29959 , n39892 );
and ( n39977 , n39975 , n39976 );
xor ( n39978 , n39975 , n39976 );
xor ( n39979 , n39308 , n39846 );
and ( n39980 , n29964 , n39892 );
and ( n39981 , n39979 , n39980 );
xor ( n39982 , n39979 , n39980 );
xor ( n39983 , n39312 , n39844 );
and ( n39984 , n29969 , n39892 );
and ( n39985 , n39983 , n39984 );
xor ( n39986 , n39983 , n39984 );
xor ( n39987 , n39316 , n39842 );
and ( n39988 , n29974 , n39892 );
and ( n39989 , n39987 , n39988 );
xor ( n39990 , n39987 , n39988 );
xor ( n39991 , n39320 , n39840 );
and ( n39992 , n29979 , n39892 );
and ( n39993 , n39991 , n39992 );
xor ( n39994 , n39991 , n39992 );
xor ( n39995 , n39324 , n39838 );
and ( n39996 , n29984 , n39892 );
and ( n39997 , n39995 , n39996 );
xor ( n39998 , n39995 , n39996 );
xor ( n39999 , n39328 , n39836 );
and ( n40000 , n29989 , n39892 );
and ( n40001 , n39999 , n40000 );
xor ( n40002 , n39999 , n40000 );
xor ( n40003 , n39332 , n39834 );
and ( n40004 , n29994 , n39892 );
and ( n40005 , n40003 , n40004 );
xor ( n40006 , n40003 , n40004 );
xor ( n40007 , n39336 , n39832 );
and ( n40008 , n29999 , n39892 );
and ( n40009 , n40007 , n40008 );
xor ( n40010 , n40007 , n40008 );
xor ( n40011 , n39340 , n39830 );
and ( n40012 , n30004 , n39892 );
and ( n40013 , n40011 , n40012 );
xor ( n40014 , n40011 , n40012 );
xor ( n40015 , n39344 , n39828 );
and ( n40016 , n30009 , n39892 );
and ( n40017 , n40015 , n40016 );
xor ( n40018 , n40015 , n40016 );
xor ( n40019 , n39348 , n39826 );
and ( n40020 , n30014 , n39892 );
and ( n40021 , n40019 , n40020 );
xor ( n40022 , n40019 , n40020 );
xor ( n40023 , n39352 , n39824 );
and ( n40024 , n30019 , n39892 );
and ( n40025 , n40023 , n40024 );
xor ( n40026 , n40023 , n40024 );
xor ( n40027 , n39356 , n39822 );
and ( n40028 , n30024 , n39892 );
and ( n40029 , n40027 , n40028 );
xor ( n40030 , n40027 , n40028 );
xor ( n40031 , n39360 , n39820 );
and ( n40032 , n30029 , n39892 );
and ( n40033 , n40031 , n40032 );
xor ( n40034 , n40031 , n40032 );
xor ( n40035 , n39364 , n39818 );
and ( n40036 , n30034 , n39892 );
and ( n40037 , n40035 , n40036 );
xor ( n40038 , n40035 , n40036 );
xor ( n40039 , n39368 , n39816 );
and ( n40040 , n30039 , n39892 );
and ( n40041 , n40039 , n40040 );
xor ( n40042 , n40039 , n40040 );
xor ( n40043 , n39372 , n39814 );
and ( n40044 , n30044 , n39892 );
and ( n40045 , n40043 , n40044 );
xor ( n40046 , n40043 , n40044 );
xor ( n40047 , n39376 , n39812 );
and ( n40048 , n30049 , n39892 );
and ( n40049 , n40047 , n40048 );
xor ( n40050 , n40047 , n40048 );
xor ( n40051 , n39380 , n39810 );
and ( n40052 , n30054 , n39892 );
and ( n40053 , n40051 , n40052 );
xor ( n40054 , n40051 , n40052 );
xor ( n40055 , n39384 , n39808 );
and ( n40056 , n30059 , n39892 );
and ( n40057 , n40055 , n40056 );
xor ( n40058 , n40055 , n40056 );
xor ( n40059 , n39388 , n39806 );
and ( n40060 , n30064 , n39892 );
and ( n40061 , n40059 , n40060 );
xor ( n40062 , n40059 , n40060 );
xor ( n40063 , n39392 , n39804 );
and ( n40064 , n30069 , n39892 );
and ( n40065 , n40063 , n40064 );
xor ( n40066 , n40063 , n40064 );
xor ( n40067 , n39396 , n39802 );
and ( n40068 , n30074 , n39892 );
and ( n40069 , n40067 , n40068 );
xor ( n40070 , n40067 , n40068 );
xor ( n40071 , n39400 , n39800 );
and ( n40072 , n30079 , n39892 );
and ( n40073 , n40071 , n40072 );
xor ( n40074 , n40071 , n40072 );
xor ( n40075 , n39404 , n39798 );
and ( n40076 , n30084 , n39892 );
and ( n40077 , n40075 , n40076 );
xor ( n40078 , n40075 , n40076 );
xor ( n40079 , n39408 , n39796 );
and ( n40080 , n30089 , n39892 );
and ( n40081 , n40079 , n40080 );
xor ( n40082 , n40079 , n40080 );
xor ( n40083 , n39412 , n39794 );
and ( n40084 , n30094 , n39892 );
and ( n40085 , n40083 , n40084 );
xor ( n40086 , n40083 , n40084 );
xor ( n40087 , n39416 , n39792 );
and ( n40088 , n30099 , n39892 );
and ( n40089 , n40087 , n40088 );
xor ( n40090 , n40087 , n40088 );
xor ( n40091 , n39420 , n39790 );
and ( n40092 , n30104 , n39892 );
and ( n40093 , n40091 , n40092 );
xor ( n40094 , n40091 , n40092 );
xor ( n40095 , n39424 , n39788 );
and ( n40096 , n30109 , n39892 );
and ( n40097 , n40095 , n40096 );
xor ( n40098 , n40095 , n40096 );
xor ( n40099 , n39428 , n39786 );
and ( n40100 , n30114 , n39892 );
and ( n40101 , n40099 , n40100 );
xor ( n40102 , n40099 , n40100 );
xor ( n40103 , n39432 , n39784 );
and ( n40104 , n30119 , n39892 );
and ( n40105 , n40103 , n40104 );
xor ( n40106 , n40103 , n40104 );
xor ( n40107 , n39436 , n39782 );
and ( n40108 , n30124 , n39892 );
and ( n40109 , n40107 , n40108 );
xor ( n40110 , n40107 , n40108 );
xor ( n40111 , n39440 , n39780 );
and ( n40112 , n30129 , n39892 );
and ( n40113 , n40111 , n40112 );
xor ( n40114 , n40111 , n40112 );
xor ( n40115 , n39444 , n39778 );
and ( n40116 , n30134 , n39892 );
and ( n40117 , n40115 , n40116 );
xor ( n40118 , n40115 , n40116 );
xor ( n40119 , n39448 , n39776 );
and ( n40120 , n30139 , n39892 );
and ( n40121 , n40119 , n40120 );
xor ( n40122 , n40119 , n40120 );
xor ( n40123 , n39452 , n39774 );
and ( n40124 , n30144 , n39892 );
and ( n40125 , n40123 , n40124 );
xor ( n40126 , n40123 , n40124 );
xor ( n40127 , n39456 , n39772 );
and ( n40128 , n30149 , n39892 );
and ( n40129 , n40127 , n40128 );
xor ( n40130 , n40127 , n40128 );
xor ( n40131 , n39460 , n39770 );
and ( n40132 , n30154 , n39892 );
and ( n40133 , n40131 , n40132 );
xor ( n40134 , n40131 , n40132 );
xor ( n40135 , n39464 , n39768 );
and ( n40136 , n30159 , n39892 );
and ( n40137 , n40135 , n40136 );
xor ( n40138 , n40135 , n40136 );
xor ( n40139 , n39468 , n39766 );
and ( n40140 , n30164 , n39892 );
and ( n40141 , n40139 , n40140 );
xor ( n40142 , n40139 , n40140 );
xor ( n40143 , n39472 , n39764 );
and ( n40144 , n30169 , n39892 );
and ( n40145 , n40143 , n40144 );
xor ( n40146 , n40143 , n40144 );
xor ( n40147 , n39476 , n39762 );
and ( n40148 , n30174 , n39892 );
and ( n40149 , n40147 , n40148 );
xor ( n40150 , n40147 , n40148 );
xor ( n40151 , n39480 , n39760 );
and ( n40152 , n30179 , n39892 );
and ( n40153 , n40151 , n40152 );
xor ( n40154 , n40151 , n40152 );
xor ( n40155 , n39484 , n39758 );
and ( n40156 , n30184 , n39892 );
and ( n40157 , n40155 , n40156 );
xor ( n40158 , n40155 , n40156 );
xor ( n40159 , n39488 , n39756 );
and ( n40160 , n30189 , n39892 );
and ( n40161 , n40159 , n40160 );
xor ( n40162 , n40159 , n40160 );
xor ( n40163 , n39492 , n39754 );
and ( n40164 , n30194 , n39892 );
and ( n40165 , n40163 , n40164 );
xor ( n40166 , n40163 , n40164 );
xor ( n40167 , n39496 , n39752 );
and ( n40168 , n30199 , n39892 );
and ( n40169 , n40167 , n40168 );
xor ( n40170 , n40167 , n40168 );
xor ( n40171 , n39500 , n39750 );
and ( n40172 , n30204 , n39892 );
and ( n40173 , n40171 , n40172 );
xor ( n40174 , n40171 , n40172 );
xor ( n40175 , n39504 , n39748 );
and ( n40176 , n30209 , n39892 );
and ( n40177 , n40175 , n40176 );
xor ( n40178 , n40175 , n40176 );
xor ( n40179 , n39508 , n39746 );
and ( n40180 , n30214 , n39892 );
and ( n40181 , n40179 , n40180 );
xor ( n40182 , n40179 , n40180 );
xor ( n40183 , n39512 , n39744 );
and ( n40184 , n30219 , n39892 );
and ( n40185 , n40183 , n40184 );
xor ( n40186 , n40183 , n40184 );
xor ( n40187 , n39516 , n39742 );
and ( n40188 , n30224 , n39892 );
and ( n40189 , n40187 , n40188 );
xor ( n40190 , n40187 , n40188 );
xor ( n40191 , n39520 , n39740 );
and ( n40192 , n30229 , n39892 );
and ( n40193 , n40191 , n40192 );
xor ( n40194 , n40191 , n40192 );
xor ( n40195 , n39524 , n39738 );
and ( n40196 , n30234 , n39892 );
and ( n40197 , n40195 , n40196 );
xor ( n40198 , n40195 , n40196 );
xor ( n40199 , n39528 , n39736 );
and ( n40200 , n30239 , n39892 );
and ( n40201 , n40199 , n40200 );
xor ( n40202 , n40199 , n40200 );
xor ( n40203 , n39532 , n39734 );
and ( n40204 , n30244 , n39892 );
and ( n40205 , n40203 , n40204 );
xor ( n40206 , n40203 , n40204 );
xor ( n40207 , n39536 , n39732 );
and ( n40208 , n30249 , n39892 );
and ( n40209 , n40207 , n40208 );
xor ( n40210 , n40207 , n40208 );
xor ( n40211 , n39540 , n39730 );
and ( n40212 , n30254 , n39892 );
and ( n40213 , n40211 , n40212 );
xor ( n40214 , n40211 , n40212 );
xor ( n40215 , n39544 , n39728 );
and ( n40216 , n30259 , n39892 );
and ( n40217 , n40215 , n40216 );
xor ( n40218 , n40215 , n40216 );
xor ( n40219 , n39548 , n39726 );
and ( n40220 , n30264 , n39892 );
and ( n40221 , n40219 , n40220 );
xor ( n40222 , n40219 , n40220 );
xor ( n40223 , n39552 , n39724 );
and ( n40224 , n30269 , n39892 );
and ( n40225 , n40223 , n40224 );
xor ( n40226 , n40223 , n40224 );
xor ( n40227 , n39556 , n39722 );
and ( n40228 , n30274 , n39892 );
and ( n40229 , n40227 , n40228 );
xor ( n40230 , n40227 , n40228 );
xor ( n40231 , n39560 , n39720 );
and ( n40232 , n30279 , n39892 );
and ( n40233 , n40231 , n40232 );
xor ( n40234 , n40231 , n40232 );
xor ( n40235 , n39564 , n39718 );
and ( n40236 , n30284 , n39892 );
and ( n40237 , n40235 , n40236 );
xor ( n40238 , n40235 , n40236 );
xor ( n40239 , n39568 , n39716 );
and ( n40240 , n30289 , n39892 );
and ( n40241 , n40239 , n40240 );
xor ( n40242 , n40239 , n40240 );
xor ( n40243 , n39572 , n39714 );
and ( n40244 , n30294 , n39892 );
and ( n40245 , n40243 , n40244 );
xor ( n40246 , n40243 , n40244 );
xor ( n40247 , n39576 , n39712 );
and ( n40248 , n30299 , n39892 );
and ( n40249 , n40247 , n40248 );
xor ( n40250 , n40247 , n40248 );
xor ( n40251 , n39580 , n39710 );
and ( n40252 , n30304 , n39892 );
and ( n40253 , n40251 , n40252 );
xor ( n40254 , n40251 , n40252 );
xor ( n40255 , n39584 , n39708 );
and ( n40256 , n30309 , n39892 );
and ( n40257 , n40255 , n40256 );
xor ( n40258 , n40255 , n40256 );
xor ( n40259 , n39588 , n39706 );
and ( n40260 , n30314 , n39892 );
and ( n40261 , n40259 , n40260 );
xor ( n40262 , n40259 , n40260 );
xor ( n40263 , n39592 , n39704 );
and ( n40264 , n30319 , n39892 );
and ( n40265 , n40263 , n40264 );
xor ( n40266 , n40263 , n40264 );
xor ( n40267 , n39596 , n39702 );
and ( n40268 , n30324 , n39892 );
and ( n40269 , n40267 , n40268 );
xor ( n40270 , n40267 , n40268 );
xor ( n40271 , n39600 , n39700 );
and ( n40272 , n30329 , n39892 );
and ( n40273 , n40271 , n40272 );
xor ( n40274 , n40271 , n40272 );
xor ( n40275 , n39604 , n39698 );
and ( n40276 , n30334 , n39892 );
and ( n40277 , n40275 , n40276 );
xor ( n40278 , n40275 , n40276 );
xor ( n40279 , n39608 , n39696 );
and ( n40280 , n30339 , n39892 );
and ( n40281 , n40279 , n40280 );
xor ( n40282 , n40279 , n40280 );
xor ( n40283 , n39612 , n39694 );
and ( n40284 , n30344 , n39892 );
and ( n40285 , n40283 , n40284 );
xor ( n40286 , n40283 , n40284 );
xor ( n40287 , n39616 , n39692 );
and ( n40288 , n30349 , n39892 );
and ( n40289 , n40287 , n40288 );
xor ( n40290 , n40287 , n40288 );
xor ( n40291 , n39620 , n39690 );
and ( n40292 , n30354 , n39892 );
and ( n40293 , n40291 , n40292 );
xor ( n40294 , n40291 , n40292 );
xor ( n40295 , n39624 , n39688 );
and ( n40296 , n30359 , n39892 );
and ( n40297 , n40295 , n40296 );
xor ( n40298 , n40295 , n40296 );
xor ( n40299 , n39628 , n39686 );
and ( n40300 , n30364 , n39892 );
and ( n40301 , n40299 , n40300 );
xor ( n40302 , n40299 , n40300 );
xor ( n40303 , n39632 , n39684 );
and ( n40304 , n30369 , n39892 );
and ( n40305 , n40303 , n40304 );
xor ( n40306 , n40303 , n40304 );
xor ( n40307 , n39636 , n39682 );
and ( n40308 , n30374 , n39892 );
and ( n40309 , n40307 , n40308 );
xor ( n40310 , n40307 , n40308 );
xor ( n40311 , n39640 , n39680 );
and ( n40312 , n30379 , n39892 );
and ( n40313 , n40311 , n40312 );
xor ( n40314 , n40311 , n40312 );
xor ( n40315 , n39644 , n39678 );
and ( n40316 , n30384 , n39892 );
and ( n40317 , n40315 , n40316 );
xor ( n40318 , n40315 , n40316 );
xor ( n40319 , n39648 , n39676 );
and ( n40320 , n30389 , n39892 );
and ( n40321 , n40319 , n40320 );
xor ( n40322 , n40319 , n40320 );
xor ( n40323 , n39652 , n39674 );
and ( n40324 , n30394 , n39892 );
and ( n40325 , n40323 , n40324 );
xor ( n40326 , n40323 , n40324 );
xor ( n40327 , n39656 , n39672 );
and ( n40328 , n30399 , n39892 );
and ( n40329 , n40327 , n40328 );
xor ( n40330 , n40327 , n40328 );
xor ( n40331 , n39660 , n39670 );
and ( n40332 , n30404 , n39892 );
and ( n40333 , n40331 , n40332 );
xor ( n40334 , n40331 , n40332 );
xor ( n40335 , n39664 , n39668 );
and ( n40336 , n30409 , n39892 );
and ( n40337 , n40335 , n40336 );
buf ( n40338 , n40337 );
and ( n40339 , n40334 , n40338 );
or ( n40340 , n40333 , n40339 );
and ( n40341 , n40330 , n40340 );
or ( n40342 , n40329 , n40341 );
and ( n40343 , n40326 , n40342 );
or ( n40344 , n40325 , n40343 );
and ( n40345 , n40322 , n40344 );
or ( n40346 , n40321 , n40345 );
and ( n40347 , n40318 , n40346 );
or ( n40348 , n40317 , n40347 );
and ( n40349 , n40314 , n40348 );
or ( n40350 , n40313 , n40349 );
and ( n40351 , n40310 , n40350 );
or ( n40352 , n40309 , n40351 );
and ( n40353 , n40306 , n40352 );
or ( n40354 , n40305 , n40353 );
and ( n40355 , n40302 , n40354 );
or ( n40356 , n40301 , n40355 );
and ( n40357 , n40298 , n40356 );
or ( n40358 , n40297 , n40357 );
and ( n40359 , n40294 , n40358 );
or ( n40360 , n40293 , n40359 );
and ( n40361 , n40290 , n40360 );
or ( n40362 , n40289 , n40361 );
and ( n40363 , n40286 , n40362 );
or ( n40364 , n40285 , n40363 );
and ( n40365 , n40282 , n40364 );
or ( n40366 , n40281 , n40365 );
and ( n40367 , n40278 , n40366 );
or ( n40368 , n40277 , n40367 );
and ( n40369 , n40274 , n40368 );
or ( n40370 , n40273 , n40369 );
and ( n40371 , n40270 , n40370 );
or ( n40372 , n40269 , n40371 );
and ( n40373 , n40266 , n40372 );
or ( n40374 , n40265 , n40373 );
and ( n40375 , n40262 , n40374 );
or ( n40376 , n40261 , n40375 );
and ( n40377 , n40258 , n40376 );
or ( n40378 , n40257 , n40377 );
and ( n40379 , n40254 , n40378 );
or ( n40380 , n40253 , n40379 );
and ( n40381 , n40250 , n40380 );
or ( n40382 , n40249 , n40381 );
and ( n40383 , n40246 , n40382 );
or ( n40384 , n40245 , n40383 );
and ( n40385 , n40242 , n40384 );
or ( n40386 , n40241 , n40385 );
and ( n40387 , n40238 , n40386 );
or ( n40388 , n40237 , n40387 );
and ( n40389 , n40234 , n40388 );
or ( n40390 , n40233 , n40389 );
and ( n40391 , n40230 , n40390 );
or ( n40392 , n40229 , n40391 );
and ( n40393 , n40226 , n40392 );
or ( n40394 , n40225 , n40393 );
and ( n40395 , n40222 , n40394 );
or ( n40396 , n40221 , n40395 );
and ( n40397 , n40218 , n40396 );
or ( n40398 , n40217 , n40397 );
and ( n40399 , n40214 , n40398 );
or ( n40400 , n40213 , n40399 );
and ( n40401 , n40210 , n40400 );
or ( n40402 , n40209 , n40401 );
and ( n40403 , n40206 , n40402 );
or ( n40404 , n40205 , n40403 );
and ( n40405 , n40202 , n40404 );
or ( n40406 , n40201 , n40405 );
and ( n40407 , n40198 , n40406 );
or ( n40408 , n40197 , n40407 );
and ( n40409 , n40194 , n40408 );
or ( n40410 , n40193 , n40409 );
and ( n40411 , n40190 , n40410 );
or ( n40412 , n40189 , n40411 );
and ( n40413 , n40186 , n40412 );
or ( n40414 , n40185 , n40413 );
and ( n40415 , n40182 , n40414 );
or ( n40416 , n40181 , n40415 );
and ( n40417 , n40178 , n40416 );
or ( n40418 , n40177 , n40417 );
and ( n40419 , n40174 , n40418 );
or ( n40420 , n40173 , n40419 );
and ( n40421 , n40170 , n40420 );
or ( n40422 , n40169 , n40421 );
and ( n40423 , n40166 , n40422 );
or ( n40424 , n40165 , n40423 );
and ( n40425 , n40162 , n40424 );
or ( n40426 , n40161 , n40425 );
and ( n40427 , n40158 , n40426 );
or ( n40428 , n40157 , n40427 );
and ( n40429 , n40154 , n40428 );
or ( n40430 , n40153 , n40429 );
and ( n40431 , n40150 , n40430 );
or ( n40432 , n40149 , n40431 );
and ( n40433 , n40146 , n40432 );
or ( n40434 , n40145 , n40433 );
and ( n40435 , n40142 , n40434 );
or ( n40436 , n40141 , n40435 );
and ( n40437 , n40138 , n40436 );
or ( n40438 , n40137 , n40437 );
and ( n40439 , n40134 , n40438 );
or ( n40440 , n40133 , n40439 );
and ( n40441 , n40130 , n40440 );
or ( n40442 , n40129 , n40441 );
and ( n40443 , n40126 , n40442 );
or ( n40444 , n40125 , n40443 );
and ( n40445 , n40122 , n40444 );
or ( n40446 , n40121 , n40445 );
and ( n40447 , n40118 , n40446 );
or ( n40448 , n40117 , n40447 );
and ( n40449 , n40114 , n40448 );
or ( n40450 , n40113 , n40449 );
and ( n40451 , n40110 , n40450 );
or ( n40452 , n40109 , n40451 );
and ( n40453 , n40106 , n40452 );
or ( n40454 , n40105 , n40453 );
and ( n40455 , n40102 , n40454 );
or ( n40456 , n40101 , n40455 );
and ( n40457 , n40098 , n40456 );
or ( n40458 , n40097 , n40457 );
and ( n40459 , n40094 , n40458 );
or ( n40460 , n40093 , n40459 );
and ( n40461 , n40090 , n40460 );
or ( n40462 , n40089 , n40461 );
and ( n40463 , n40086 , n40462 );
or ( n40464 , n40085 , n40463 );
and ( n40465 , n40082 , n40464 );
or ( n40466 , n40081 , n40465 );
and ( n40467 , n40078 , n40466 );
or ( n40468 , n40077 , n40467 );
and ( n40469 , n40074 , n40468 );
or ( n40470 , n40073 , n40469 );
and ( n40471 , n40070 , n40470 );
or ( n40472 , n40069 , n40471 );
and ( n40473 , n40066 , n40472 );
or ( n40474 , n40065 , n40473 );
and ( n40475 , n40062 , n40474 );
or ( n40476 , n40061 , n40475 );
and ( n40477 , n40058 , n40476 );
or ( n40478 , n40057 , n40477 );
and ( n40479 , n40054 , n40478 );
or ( n40480 , n40053 , n40479 );
and ( n40481 , n40050 , n40480 );
or ( n40482 , n40049 , n40481 );
and ( n40483 , n40046 , n40482 );
or ( n40484 , n40045 , n40483 );
and ( n40485 , n40042 , n40484 );
or ( n40486 , n40041 , n40485 );
and ( n40487 , n40038 , n40486 );
or ( n40488 , n40037 , n40487 );
and ( n40489 , n40034 , n40488 );
or ( n40490 , n40033 , n40489 );
and ( n40491 , n40030 , n40490 );
or ( n40492 , n40029 , n40491 );
and ( n40493 , n40026 , n40492 );
or ( n40494 , n40025 , n40493 );
and ( n40495 , n40022 , n40494 );
or ( n40496 , n40021 , n40495 );
and ( n40497 , n40018 , n40496 );
or ( n40498 , n40017 , n40497 );
and ( n40499 , n40014 , n40498 );
or ( n40500 , n40013 , n40499 );
and ( n40501 , n40010 , n40500 );
or ( n40502 , n40009 , n40501 );
and ( n40503 , n40006 , n40502 );
or ( n40504 , n40005 , n40503 );
and ( n40505 , n40002 , n40504 );
or ( n40506 , n40001 , n40505 );
and ( n40507 , n39998 , n40506 );
or ( n40508 , n39997 , n40507 );
and ( n40509 , n39994 , n40508 );
or ( n40510 , n39993 , n40509 );
and ( n40511 , n39990 , n40510 );
or ( n40512 , n39989 , n40511 );
and ( n40513 , n39986 , n40512 );
or ( n40514 , n39985 , n40513 );
and ( n40515 , n39982 , n40514 );
or ( n40516 , n39981 , n40515 );
and ( n40517 , n39978 , n40516 );
or ( n40518 , n39977 , n40517 );
and ( n40519 , n39974 , n40518 );
or ( n40520 , n39973 , n40519 );
and ( n40521 , n39970 , n40520 );
or ( n40522 , n39969 , n40521 );
and ( n40523 , n39966 , n40522 );
or ( n40524 , n39965 , n40523 );
and ( n40525 , n39962 , n40524 );
or ( n40526 , n39961 , n40525 );
and ( n40527 , n39958 , n40526 );
or ( n40528 , n39957 , n40527 );
and ( n40529 , n39954 , n40528 );
or ( n40530 , n39953 , n40529 );
and ( n40531 , n39950 , n40530 );
or ( n40532 , n39949 , n40531 );
and ( n40533 , n39946 , n40532 );
or ( n40534 , n39945 , n40533 );
and ( n40535 , n39942 , n40534 );
or ( n40536 , n39941 , n40535 );
and ( n40537 , n39938 , n40536 );
or ( n40538 , n39937 , n40537 );
and ( n40539 , n39934 , n40538 );
or ( n40540 , n39933 , n40539 );
and ( n40541 , n39930 , n40540 );
or ( n40542 , n39929 , n40541 );
and ( n40543 , n39926 , n40542 );
or ( n40544 , n39925 , n40543 );
and ( n40545 , n39922 , n40544 );
or ( n40546 , n39921 , n40545 );
and ( n40547 , n39918 , n40546 );
or ( n40548 , n39917 , n40547 );
and ( n40549 , n39914 , n40548 );
or ( n40550 , n39913 , n40549 );
and ( n40551 , n39910 , n40550 );
or ( n40552 , n39909 , n40551 );
and ( n40553 , n39906 , n40552 );
or ( n40554 , n39905 , n40553 );
and ( n40555 , n39902 , n40554 );
or ( n40556 , n39901 , n40555 );
and ( n40557 , n39898 , n40556 );
or ( n40558 , n39897 , n40557 );
xor ( n40559 , n39894 , n40558 );
buf ( n40560 , n18074 );
and ( n40561 , n29859 , n40560 );
xor ( n40562 , n40559 , n40561 );
xor ( n40563 , n39898 , n40556 );
and ( n40564 , n29864 , n40560 );
and ( n40565 , n40563 , n40564 );
xor ( n40566 , n40563 , n40564 );
xor ( n40567 , n39902 , n40554 );
and ( n40568 , n29869 , n40560 );
and ( n40569 , n40567 , n40568 );
xor ( n40570 , n40567 , n40568 );
xor ( n40571 , n39906 , n40552 );
and ( n40572 , n29874 , n40560 );
and ( n40573 , n40571 , n40572 );
xor ( n40574 , n40571 , n40572 );
xor ( n40575 , n39910 , n40550 );
and ( n40576 , n29879 , n40560 );
and ( n40577 , n40575 , n40576 );
xor ( n40578 , n40575 , n40576 );
xor ( n40579 , n39914 , n40548 );
and ( n40580 , n29884 , n40560 );
and ( n40581 , n40579 , n40580 );
xor ( n40582 , n40579 , n40580 );
xor ( n40583 , n39918 , n40546 );
and ( n40584 , n29889 , n40560 );
and ( n40585 , n40583 , n40584 );
xor ( n40586 , n40583 , n40584 );
xor ( n40587 , n39922 , n40544 );
and ( n40588 , n29894 , n40560 );
and ( n40589 , n40587 , n40588 );
xor ( n40590 , n40587 , n40588 );
xor ( n40591 , n39926 , n40542 );
and ( n40592 , n29899 , n40560 );
and ( n40593 , n40591 , n40592 );
xor ( n40594 , n40591 , n40592 );
xor ( n40595 , n39930 , n40540 );
and ( n40596 , n29904 , n40560 );
and ( n40597 , n40595 , n40596 );
xor ( n40598 , n40595 , n40596 );
xor ( n40599 , n39934 , n40538 );
and ( n40600 , n29909 , n40560 );
and ( n40601 , n40599 , n40600 );
xor ( n40602 , n40599 , n40600 );
xor ( n40603 , n39938 , n40536 );
and ( n40604 , n29914 , n40560 );
and ( n40605 , n40603 , n40604 );
xor ( n40606 , n40603 , n40604 );
xor ( n40607 , n39942 , n40534 );
and ( n40608 , n29919 , n40560 );
and ( n40609 , n40607 , n40608 );
xor ( n40610 , n40607 , n40608 );
xor ( n40611 , n39946 , n40532 );
and ( n40612 , n29924 , n40560 );
and ( n40613 , n40611 , n40612 );
xor ( n40614 , n40611 , n40612 );
xor ( n40615 , n39950 , n40530 );
and ( n40616 , n29929 , n40560 );
and ( n40617 , n40615 , n40616 );
xor ( n40618 , n40615 , n40616 );
xor ( n40619 , n39954 , n40528 );
and ( n40620 , n29934 , n40560 );
and ( n40621 , n40619 , n40620 );
xor ( n40622 , n40619 , n40620 );
xor ( n40623 , n39958 , n40526 );
and ( n40624 , n29939 , n40560 );
and ( n40625 , n40623 , n40624 );
xor ( n40626 , n40623 , n40624 );
xor ( n40627 , n39962 , n40524 );
and ( n40628 , n29944 , n40560 );
and ( n40629 , n40627 , n40628 );
xor ( n40630 , n40627 , n40628 );
xor ( n40631 , n39966 , n40522 );
and ( n40632 , n29949 , n40560 );
and ( n40633 , n40631 , n40632 );
xor ( n40634 , n40631 , n40632 );
xor ( n40635 , n39970 , n40520 );
and ( n40636 , n29954 , n40560 );
and ( n40637 , n40635 , n40636 );
xor ( n40638 , n40635 , n40636 );
xor ( n40639 , n39974 , n40518 );
and ( n40640 , n29959 , n40560 );
and ( n40641 , n40639 , n40640 );
xor ( n40642 , n40639 , n40640 );
xor ( n40643 , n39978 , n40516 );
and ( n40644 , n29964 , n40560 );
and ( n40645 , n40643 , n40644 );
xor ( n40646 , n40643 , n40644 );
xor ( n40647 , n39982 , n40514 );
and ( n40648 , n29969 , n40560 );
and ( n40649 , n40647 , n40648 );
xor ( n40650 , n40647 , n40648 );
xor ( n40651 , n39986 , n40512 );
and ( n40652 , n29974 , n40560 );
and ( n40653 , n40651 , n40652 );
xor ( n40654 , n40651 , n40652 );
xor ( n40655 , n39990 , n40510 );
and ( n40656 , n29979 , n40560 );
and ( n40657 , n40655 , n40656 );
xor ( n40658 , n40655 , n40656 );
xor ( n40659 , n39994 , n40508 );
and ( n40660 , n29984 , n40560 );
and ( n40661 , n40659 , n40660 );
xor ( n40662 , n40659 , n40660 );
xor ( n40663 , n39998 , n40506 );
and ( n40664 , n29989 , n40560 );
and ( n40665 , n40663 , n40664 );
xor ( n40666 , n40663 , n40664 );
xor ( n40667 , n40002 , n40504 );
and ( n40668 , n29994 , n40560 );
and ( n40669 , n40667 , n40668 );
xor ( n40670 , n40667 , n40668 );
xor ( n40671 , n40006 , n40502 );
and ( n40672 , n29999 , n40560 );
and ( n40673 , n40671 , n40672 );
xor ( n40674 , n40671 , n40672 );
xor ( n40675 , n40010 , n40500 );
and ( n40676 , n30004 , n40560 );
and ( n40677 , n40675 , n40676 );
xor ( n40678 , n40675 , n40676 );
xor ( n40679 , n40014 , n40498 );
and ( n40680 , n30009 , n40560 );
and ( n40681 , n40679 , n40680 );
xor ( n40682 , n40679 , n40680 );
xor ( n40683 , n40018 , n40496 );
and ( n40684 , n30014 , n40560 );
and ( n40685 , n40683 , n40684 );
xor ( n40686 , n40683 , n40684 );
xor ( n40687 , n40022 , n40494 );
and ( n40688 , n30019 , n40560 );
and ( n40689 , n40687 , n40688 );
xor ( n40690 , n40687 , n40688 );
xor ( n40691 , n40026 , n40492 );
and ( n40692 , n30024 , n40560 );
and ( n40693 , n40691 , n40692 );
xor ( n40694 , n40691 , n40692 );
xor ( n40695 , n40030 , n40490 );
and ( n40696 , n30029 , n40560 );
and ( n40697 , n40695 , n40696 );
xor ( n40698 , n40695 , n40696 );
xor ( n40699 , n40034 , n40488 );
and ( n40700 , n30034 , n40560 );
and ( n40701 , n40699 , n40700 );
xor ( n40702 , n40699 , n40700 );
xor ( n40703 , n40038 , n40486 );
and ( n40704 , n30039 , n40560 );
and ( n40705 , n40703 , n40704 );
xor ( n40706 , n40703 , n40704 );
xor ( n40707 , n40042 , n40484 );
and ( n40708 , n30044 , n40560 );
and ( n40709 , n40707 , n40708 );
xor ( n40710 , n40707 , n40708 );
xor ( n40711 , n40046 , n40482 );
and ( n40712 , n30049 , n40560 );
and ( n40713 , n40711 , n40712 );
xor ( n40714 , n40711 , n40712 );
xor ( n40715 , n40050 , n40480 );
and ( n40716 , n30054 , n40560 );
and ( n40717 , n40715 , n40716 );
xor ( n40718 , n40715 , n40716 );
xor ( n40719 , n40054 , n40478 );
and ( n40720 , n30059 , n40560 );
and ( n40721 , n40719 , n40720 );
xor ( n40722 , n40719 , n40720 );
xor ( n40723 , n40058 , n40476 );
and ( n40724 , n30064 , n40560 );
and ( n40725 , n40723 , n40724 );
xor ( n40726 , n40723 , n40724 );
xor ( n40727 , n40062 , n40474 );
and ( n40728 , n30069 , n40560 );
and ( n40729 , n40727 , n40728 );
xor ( n40730 , n40727 , n40728 );
xor ( n40731 , n40066 , n40472 );
and ( n40732 , n30074 , n40560 );
and ( n40733 , n40731 , n40732 );
xor ( n40734 , n40731 , n40732 );
xor ( n40735 , n40070 , n40470 );
and ( n40736 , n30079 , n40560 );
and ( n40737 , n40735 , n40736 );
xor ( n40738 , n40735 , n40736 );
xor ( n40739 , n40074 , n40468 );
and ( n40740 , n30084 , n40560 );
and ( n40741 , n40739 , n40740 );
xor ( n40742 , n40739 , n40740 );
xor ( n40743 , n40078 , n40466 );
and ( n40744 , n30089 , n40560 );
and ( n40745 , n40743 , n40744 );
xor ( n40746 , n40743 , n40744 );
xor ( n40747 , n40082 , n40464 );
and ( n40748 , n30094 , n40560 );
and ( n40749 , n40747 , n40748 );
xor ( n40750 , n40747 , n40748 );
xor ( n40751 , n40086 , n40462 );
and ( n40752 , n30099 , n40560 );
and ( n40753 , n40751 , n40752 );
xor ( n40754 , n40751 , n40752 );
xor ( n40755 , n40090 , n40460 );
and ( n40756 , n30104 , n40560 );
and ( n40757 , n40755 , n40756 );
xor ( n40758 , n40755 , n40756 );
xor ( n40759 , n40094 , n40458 );
and ( n40760 , n30109 , n40560 );
and ( n40761 , n40759 , n40760 );
xor ( n40762 , n40759 , n40760 );
xor ( n40763 , n40098 , n40456 );
and ( n40764 , n30114 , n40560 );
and ( n40765 , n40763 , n40764 );
xor ( n40766 , n40763 , n40764 );
xor ( n40767 , n40102 , n40454 );
and ( n40768 , n30119 , n40560 );
and ( n40769 , n40767 , n40768 );
xor ( n40770 , n40767 , n40768 );
xor ( n40771 , n40106 , n40452 );
and ( n40772 , n30124 , n40560 );
and ( n40773 , n40771 , n40772 );
xor ( n40774 , n40771 , n40772 );
xor ( n40775 , n40110 , n40450 );
and ( n40776 , n30129 , n40560 );
and ( n40777 , n40775 , n40776 );
xor ( n40778 , n40775 , n40776 );
xor ( n40779 , n40114 , n40448 );
and ( n40780 , n30134 , n40560 );
and ( n40781 , n40779 , n40780 );
xor ( n40782 , n40779 , n40780 );
xor ( n40783 , n40118 , n40446 );
and ( n40784 , n30139 , n40560 );
and ( n40785 , n40783 , n40784 );
xor ( n40786 , n40783 , n40784 );
xor ( n40787 , n40122 , n40444 );
and ( n40788 , n30144 , n40560 );
and ( n40789 , n40787 , n40788 );
xor ( n40790 , n40787 , n40788 );
xor ( n40791 , n40126 , n40442 );
and ( n40792 , n30149 , n40560 );
and ( n40793 , n40791 , n40792 );
xor ( n40794 , n40791 , n40792 );
xor ( n40795 , n40130 , n40440 );
and ( n40796 , n30154 , n40560 );
and ( n40797 , n40795 , n40796 );
xor ( n40798 , n40795 , n40796 );
xor ( n40799 , n40134 , n40438 );
and ( n40800 , n30159 , n40560 );
and ( n40801 , n40799 , n40800 );
xor ( n40802 , n40799 , n40800 );
xor ( n40803 , n40138 , n40436 );
and ( n40804 , n30164 , n40560 );
and ( n40805 , n40803 , n40804 );
xor ( n40806 , n40803 , n40804 );
xor ( n40807 , n40142 , n40434 );
and ( n40808 , n30169 , n40560 );
and ( n40809 , n40807 , n40808 );
xor ( n40810 , n40807 , n40808 );
xor ( n40811 , n40146 , n40432 );
and ( n40812 , n30174 , n40560 );
and ( n40813 , n40811 , n40812 );
xor ( n40814 , n40811 , n40812 );
xor ( n40815 , n40150 , n40430 );
and ( n40816 , n30179 , n40560 );
and ( n40817 , n40815 , n40816 );
xor ( n40818 , n40815 , n40816 );
xor ( n40819 , n40154 , n40428 );
and ( n40820 , n30184 , n40560 );
and ( n40821 , n40819 , n40820 );
xor ( n40822 , n40819 , n40820 );
xor ( n40823 , n40158 , n40426 );
and ( n40824 , n30189 , n40560 );
and ( n40825 , n40823 , n40824 );
xor ( n40826 , n40823 , n40824 );
xor ( n40827 , n40162 , n40424 );
and ( n40828 , n30194 , n40560 );
and ( n40829 , n40827 , n40828 );
xor ( n40830 , n40827 , n40828 );
xor ( n40831 , n40166 , n40422 );
and ( n40832 , n30199 , n40560 );
and ( n40833 , n40831 , n40832 );
xor ( n40834 , n40831 , n40832 );
xor ( n40835 , n40170 , n40420 );
and ( n40836 , n30204 , n40560 );
and ( n40837 , n40835 , n40836 );
xor ( n40838 , n40835 , n40836 );
xor ( n40839 , n40174 , n40418 );
and ( n40840 , n30209 , n40560 );
and ( n40841 , n40839 , n40840 );
xor ( n40842 , n40839 , n40840 );
xor ( n40843 , n40178 , n40416 );
and ( n40844 , n30214 , n40560 );
and ( n40845 , n40843 , n40844 );
xor ( n40846 , n40843 , n40844 );
xor ( n40847 , n40182 , n40414 );
and ( n40848 , n30219 , n40560 );
and ( n40849 , n40847 , n40848 );
xor ( n40850 , n40847 , n40848 );
xor ( n40851 , n40186 , n40412 );
and ( n40852 , n30224 , n40560 );
and ( n40853 , n40851 , n40852 );
xor ( n40854 , n40851 , n40852 );
xor ( n40855 , n40190 , n40410 );
and ( n40856 , n30229 , n40560 );
and ( n40857 , n40855 , n40856 );
xor ( n40858 , n40855 , n40856 );
xor ( n40859 , n40194 , n40408 );
and ( n40860 , n30234 , n40560 );
and ( n40861 , n40859 , n40860 );
xor ( n40862 , n40859 , n40860 );
xor ( n40863 , n40198 , n40406 );
and ( n40864 , n30239 , n40560 );
and ( n40865 , n40863 , n40864 );
xor ( n40866 , n40863 , n40864 );
xor ( n40867 , n40202 , n40404 );
and ( n40868 , n30244 , n40560 );
and ( n40869 , n40867 , n40868 );
xor ( n40870 , n40867 , n40868 );
xor ( n40871 , n40206 , n40402 );
and ( n40872 , n30249 , n40560 );
and ( n40873 , n40871 , n40872 );
xor ( n40874 , n40871 , n40872 );
xor ( n40875 , n40210 , n40400 );
and ( n40876 , n30254 , n40560 );
and ( n40877 , n40875 , n40876 );
xor ( n40878 , n40875 , n40876 );
xor ( n40879 , n40214 , n40398 );
and ( n40880 , n30259 , n40560 );
and ( n40881 , n40879 , n40880 );
xor ( n40882 , n40879 , n40880 );
xor ( n40883 , n40218 , n40396 );
and ( n40884 , n30264 , n40560 );
and ( n40885 , n40883 , n40884 );
xor ( n40886 , n40883 , n40884 );
xor ( n40887 , n40222 , n40394 );
and ( n40888 , n30269 , n40560 );
and ( n40889 , n40887 , n40888 );
xor ( n40890 , n40887 , n40888 );
xor ( n40891 , n40226 , n40392 );
and ( n40892 , n30274 , n40560 );
and ( n40893 , n40891 , n40892 );
xor ( n40894 , n40891 , n40892 );
xor ( n40895 , n40230 , n40390 );
and ( n40896 , n30279 , n40560 );
and ( n40897 , n40895 , n40896 );
xor ( n40898 , n40895 , n40896 );
xor ( n40899 , n40234 , n40388 );
and ( n40900 , n30284 , n40560 );
and ( n40901 , n40899 , n40900 );
xor ( n40902 , n40899 , n40900 );
xor ( n40903 , n40238 , n40386 );
and ( n40904 , n30289 , n40560 );
and ( n40905 , n40903 , n40904 );
xor ( n40906 , n40903 , n40904 );
xor ( n40907 , n40242 , n40384 );
and ( n40908 , n30294 , n40560 );
and ( n40909 , n40907 , n40908 );
xor ( n40910 , n40907 , n40908 );
xor ( n40911 , n40246 , n40382 );
and ( n40912 , n30299 , n40560 );
and ( n40913 , n40911 , n40912 );
xor ( n40914 , n40911 , n40912 );
xor ( n40915 , n40250 , n40380 );
and ( n40916 , n30304 , n40560 );
and ( n40917 , n40915 , n40916 );
xor ( n40918 , n40915 , n40916 );
xor ( n40919 , n40254 , n40378 );
and ( n40920 , n30309 , n40560 );
and ( n40921 , n40919 , n40920 );
xor ( n40922 , n40919 , n40920 );
xor ( n40923 , n40258 , n40376 );
and ( n40924 , n30314 , n40560 );
and ( n40925 , n40923 , n40924 );
xor ( n40926 , n40923 , n40924 );
xor ( n40927 , n40262 , n40374 );
and ( n40928 , n30319 , n40560 );
and ( n40929 , n40927 , n40928 );
xor ( n40930 , n40927 , n40928 );
xor ( n40931 , n40266 , n40372 );
and ( n40932 , n30324 , n40560 );
and ( n40933 , n40931 , n40932 );
xor ( n40934 , n40931 , n40932 );
xor ( n40935 , n40270 , n40370 );
and ( n40936 , n30329 , n40560 );
and ( n40937 , n40935 , n40936 );
xor ( n40938 , n40935 , n40936 );
xor ( n40939 , n40274 , n40368 );
and ( n40940 , n30334 , n40560 );
and ( n40941 , n40939 , n40940 );
xor ( n40942 , n40939 , n40940 );
xor ( n40943 , n40278 , n40366 );
and ( n40944 , n30339 , n40560 );
and ( n40945 , n40943 , n40944 );
xor ( n40946 , n40943 , n40944 );
xor ( n40947 , n40282 , n40364 );
and ( n40948 , n30344 , n40560 );
and ( n40949 , n40947 , n40948 );
xor ( n40950 , n40947 , n40948 );
xor ( n40951 , n40286 , n40362 );
and ( n40952 , n30349 , n40560 );
and ( n40953 , n40951 , n40952 );
xor ( n40954 , n40951 , n40952 );
xor ( n40955 , n40290 , n40360 );
and ( n40956 , n30354 , n40560 );
and ( n40957 , n40955 , n40956 );
xor ( n40958 , n40955 , n40956 );
xor ( n40959 , n40294 , n40358 );
and ( n40960 , n30359 , n40560 );
and ( n40961 , n40959 , n40960 );
xor ( n40962 , n40959 , n40960 );
xor ( n40963 , n40298 , n40356 );
and ( n40964 , n30364 , n40560 );
and ( n40965 , n40963 , n40964 );
xor ( n40966 , n40963 , n40964 );
xor ( n40967 , n40302 , n40354 );
and ( n40968 , n30369 , n40560 );
and ( n40969 , n40967 , n40968 );
xor ( n40970 , n40967 , n40968 );
xor ( n40971 , n40306 , n40352 );
and ( n40972 , n30374 , n40560 );
and ( n40973 , n40971 , n40972 );
xor ( n40974 , n40971 , n40972 );
xor ( n40975 , n40310 , n40350 );
and ( n40976 , n30379 , n40560 );
and ( n40977 , n40975 , n40976 );
xor ( n40978 , n40975 , n40976 );
xor ( n40979 , n40314 , n40348 );
and ( n40980 , n30384 , n40560 );
and ( n40981 , n40979 , n40980 );
xor ( n40982 , n40979 , n40980 );
xor ( n40983 , n40318 , n40346 );
and ( n40984 , n30389 , n40560 );
and ( n40985 , n40983 , n40984 );
xor ( n40986 , n40983 , n40984 );
xor ( n40987 , n40322 , n40344 );
and ( n40988 , n30394 , n40560 );
and ( n40989 , n40987 , n40988 );
xor ( n40990 , n40987 , n40988 );
xor ( n40991 , n40326 , n40342 );
and ( n40992 , n30399 , n40560 );
and ( n40993 , n40991 , n40992 );
xor ( n40994 , n40991 , n40992 );
xor ( n40995 , n40330 , n40340 );
and ( n40996 , n30404 , n40560 );
and ( n40997 , n40995 , n40996 );
xor ( n40998 , n40995 , n40996 );
xor ( n40999 , n40334 , n40338 );
and ( n41000 , n30409 , n40560 );
and ( n41001 , n40999 , n41000 );
buf ( n41002 , n41001 );
and ( n41003 , n40998 , n41002 );
or ( n41004 , n40997 , n41003 );
and ( n41005 , n40994 , n41004 );
or ( n41006 , n40993 , n41005 );
and ( n41007 , n40990 , n41006 );
or ( n41008 , n40989 , n41007 );
and ( n41009 , n40986 , n41008 );
or ( n41010 , n40985 , n41009 );
and ( n41011 , n40982 , n41010 );
or ( n41012 , n40981 , n41011 );
and ( n41013 , n40978 , n41012 );
or ( n41014 , n40977 , n41013 );
and ( n41015 , n40974 , n41014 );
or ( n41016 , n40973 , n41015 );
and ( n41017 , n40970 , n41016 );
or ( n41018 , n40969 , n41017 );
and ( n41019 , n40966 , n41018 );
or ( n41020 , n40965 , n41019 );
and ( n41021 , n40962 , n41020 );
or ( n41022 , n40961 , n41021 );
and ( n41023 , n40958 , n41022 );
or ( n41024 , n40957 , n41023 );
and ( n41025 , n40954 , n41024 );
or ( n41026 , n40953 , n41025 );
and ( n41027 , n40950 , n41026 );
or ( n41028 , n40949 , n41027 );
and ( n41029 , n40946 , n41028 );
or ( n41030 , n40945 , n41029 );
and ( n41031 , n40942 , n41030 );
or ( n41032 , n40941 , n41031 );
and ( n41033 , n40938 , n41032 );
or ( n41034 , n40937 , n41033 );
and ( n41035 , n40934 , n41034 );
or ( n41036 , n40933 , n41035 );
and ( n41037 , n40930 , n41036 );
or ( n41038 , n40929 , n41037 );
and ( n41039 , n40926 , n41038 );
or ( n41040 , n40925 , n41039 );
and ( n41041 , n40922 , n41040 );
or ( n41042 , n40921 , n41041 );
and ( n41043 , n40918 , n41042 );
or ( n41044 , n40917 , n41043 );
and ( n41045 , n40914 , n41044 );
or ( n41046 , n40913 , n41045 );
and ( n41047 , n40910 , n41046 );
or ( n41048 , n40909 , n41047 );
and ( n41049 , n40906 , n41048 );
or ( n41050 , n40905 , n41049 );
and ( n41051 , n40902 , n41050 );
or ( n41052 , n40901 , n41051 );
and ( n41053 , n40898 , n41052 );
or ( n41054 , n40897 , n41053 );
and ( n41055 , n40894 , n41054 );
or ( n41056 , n40893 , n41055 );
and ( n41057 , n40890 , n41056 );
or ( n41058 , n40889 , n41057 );
and ( n41059 , n40886 , n41058 );
or ( n41060 , n40885 , n41059 );
and ( n41061 , n40882 , n41060 );
or ( n41062 , n40881 , n41061 );
and ( n41063 , n40878 , n41062 );
or ( n41064 , n40877 , n41063 );
and ( n41065 , n40874 , n41064 );
or ( n41066 , n40873 , n41065 );
and ( n41067 , n40870 , n41066 );
or ( n41068 , n40869 , n41067 );
and ( n41069 , n40866 , n41068 );
or ( n41070 , n40865 , n41069 );
and ( n41071 , n40862 , n41070 );
or ( n41072 , n40861 , n41071 );
and ( n41073 , n40858 , n41072 );
or ( n41074 , n40857 , n41073 );
and ( n41075 , n40854 , n41074 );
or ( n41076 , n40853 , n41075 );
and ( n41077 , n40850 , n41076 );
or ( n41078 , n40849 , n41077 );
and ( n41079 , n40846 , n41078 );
or ( n41080 , n40845 , n41079 );
and ( n41081 , n40842 , n41080 );
or ( n41082 , n40841 , n41081 );
and ( n41083 , n40838 , n41082 );
or ( n41084 , n40837 , n41083 );
and ( n41085 , n40834 , n41084 );
or ( n41086 , n40833 , n41085 );
and ( n41087 , n40830 , n41086 );
or ( n41088 , n40829 , n41087 );
and ( n41089 , n40826 , n41088 );
or ( n41090 , n40825 , n41089 );
and ( n41091 , n40822 , n41090 );
or ( n41092 , n40821 , n41091 );
and ( n41093 , n40818 , n41092 );
or ( n41094 , n40817 , n41093 );
and ( n41095 , n40814 , n41094 );
or ( n41096 , n40813 , n41095 );
and ( n41097 , n40810 , n41096 );
or ( n41098 , n40809 , n41097 );
and ( n41099 , n40806 , n41098 );
or ( n41100 , n40805 , n41099 );
and ( n41101 , n40802 , n41100 );
or ( n41102 , n40801 , n41101 );
and ( n41103 , n40798 , n41102 );
or ( n41104 , n40797 , n41103 );
and ( n41105 , n40794 , n41104 );
or ( n41106 , n40793 , n41105 );
and ( n41107 , n40790 , n41106 );
or ( n41108 , n40789 , n41107 );
and ( n41109 , n40786 , n41108 );
or ( n41110 , n40785 , n41109 );
and ( n41111 , n40782 , n41110 );
or ( n41112 , n40781 , n41111 );
and ( n41113 , n40778 , n41112 );
or ( n41114 , n40777 , n41113 );
and ( n41115 , n40774 , n41114 );
or ( n41116 , n40773 , n41115 );
and ( n41117 , n40770 , n41116 );
or ( n41118 , n40769 , n41117 );
and ( n41119 , n40766 , n41118 );
or ( n41120 , n40765 , n41119 );
and ( n41121 , n40762 , n41120 );
or ( n41122 , n40761 , n41121 );
and ( n41123 , n40758 , n41122 );
or ( n41124 , n40757 , n41123 );
and ( n41125 , n40754 , n41124 );
or ( n41126 , n40753 , n41125 );
and ( n41127 , n40750 , n41126 );
or ( n41128 , n40749 , n41127 );
and ( n41129 , n40746 , n41128 );
or ( n41130 , n40745 , n41129 );
and ( n41131 , n40742 , n41130 );
or ( n41132 , n40741 , n41131 );
and ( n41133 , n40738 , n41132 );
or ( n41134 , n40737 , n41133 );
and ( n41135 , n40734 , n41134 );
or ( n41136 , n40733 , n41135 );
and ( n41137 , n40730 , n41136 );
or ( n41138 , n40729 , n41137 );
and ( n41139 , n40726 , n41138 );
or ( n41140 , n40725 , n41139 );
and ( n41141 , n40722 , n41140 );
or ( n41142 , n40721 , n41141 );
and ( n41143 , n40718 , n41142 );
or ( n41144 , n40717 , n41143 );
and ( n41145 , n40714 , n41144 );
or ( n41146 , n40713 , n41145 );
and ( n41147 , n40710 , n41146 );
or ( n41148 , n40709 , n41147 );
and ( n41149 , n40706 , n41148 );
or ( n41150 , n40705 , n41149 );
and ( n41151 , n40702 , n41150 );
or ( n41152 , n40701 , n41151 );
and ( n41153 , n40698 , n41152 );
or ( n41154 , n40697 , n41153 );
and ( n41155 , n40694 , n41154 );
or ( n41156 , n40693 , n41155 );
and ( n41157 , n40690 , n41156 );
or ( n41158 , n40689 , n41157 );
and ( n41159 , n40686 , n41158 );
or ( n41160 , n40685 , n41159 );
and ( n41161 , n40682 , n41160 );
or ( n41162 , n40681 , n41161 );
and ( n41163 , n40678 , n41162 );
or ( n41164 , n40677 , n41163 );
and ( n41165 , n40674 , n41164 );
or ( n41166 , n40673 , n41165 );
and ( n41167 , n40670 , n41166 );
or ( n41168 , n40669 , n41167 );
and ( n41169 , n40666 , n41168 );
or ( n41170 , n40665 , n41169 );
and ( n41171 , n40662 , n41170 );
or ( n41172 , n40661 , n41171 );
and ( n41173 , n40658 , n41172 );
or ( n41174 , n40657 , n41173 );
and ( n41175 , n40654 , n41174 );
or ( n41176 , n40653 , n41175 );
and ( n41177 , n40650 , n41176 );
or ( n41178 , n40649 , n41177 );
and ( n41179 , n40646 , n41178 );
or ( n41180 , n40645 , n41179 );
and ( n41181 , n40642 , n41180 );
or ( n41182 , n40641 , n41181 );
and ( n41183 , n40638 , n41182 );
or ( n41184 , n40637 , n41183 );
and ( n41185 , n40634 , n41184 );
or ( n41186 , n40633 , n41185 );
and ( n41187 , n40630 , n41186 );
or ( n41188 , n40629 , n41187 );
and ( n41189 , n40626 , n41188 );
or ( n41190 , n40625 , n41189 );
and ( n41191 , n40622 , n41190 );
or ( n41192 , n40621 , n41191 );
and ( n41193 , n40618 , n41192 );
or ( n41194 , n40617 , n41193 );
and ( n41195 , n40614 , n41194 );
or ( n41196 , n40613 , n41195 );
and ( n41197 , n40610 , n41196 );
or ( n41198 , n40609 , n41197 );
and ( n41199 , n40606 , n41198 );
or ( n41200 , n40605 , n41199 );
and ( n41201 , n40602 , n41200 );
or ( n41202 , n40601 , n41201 );
and ( n41203 , n40598 , n41202 );
or ( n41204 , n40597 , n41203 );
and ( n41205 , n40594 , n41204 );
or ( n41206 , n40593 , n41205 );
and ( n41207 , n40590 , n41206 );
or ( n41208 , n40589 , n41207 );
and ( n41209 , n40586 , n41208 );
or ( n41210 , n40585 , n41209 );
and ( n41211 , n40582 , n41210 );
or ( n41212 , n40581 , n41211 );
and ( n41213 , n40578 , n41212 );
or ( n41214 , n40577 , n41213 );
and ( n41215 , n40574 , n41214 );
or ( n41216 , n40573 , n41215 );
and ( n41217 , n40570 , n41216 );
or ( n41218 , n40569 , n41217 );
and ( n41219 , n40566 , n41218 );
or ( n41220 , n40565 , n41219 );
xor ( n41221 , n40562 , n41220 );
buf ( n41222 , n18072 );
and ( n41223 , n29864 , n41222 );
xor ( n41224 , n41221 , n41223 );
xor ( n41225 , n40566 , n41218 );
and ( n41226 , n29869 , n41222 );
and ( n41227 , n41225 , n41226 );
xor ( n41228 , n41225 , n41226 );
xor ( n41229 , n40570 , n41216 );
and ( n41230 , n29874 , n41222 );
and ( n41231 , n41229 , n41230 );
xor ( n41232 , n41229 , n41230 );
xor ( n41233 , n40574 , n41214 );
and ( n41234 , n29879 , n41222 );
and ( n41235 , n41233 , n41234 );
xor ( n41236 , n41233 , n41234 );
xor ( n41237 , n40578 , n41212 );
and ( n41238 , n29884 , n41222 );
and ( n41239 , n41237 , n41238 );
xor ( n41240 , n41237 , n41238 );
xor ( n41241 , n40582 , n41210 );
and ( n41242 , n29889 , n41222 );
and ( n41243 , n41241 , n41242 );
xor ( n41244 , n41241 , n41242 );
xor ( n41245 , n40586 , n41208 );
and ( n41246 , n29894 , n41222 );
and ( n41247 , n41245 , n41246 );
xor ( n41248 , n41245 , n41246 );
xor ( n41249 , n40590 , n41206 );
and ( n41250 , n29899 , n41222 );
and ( n41251 , n41249 , n41250 );
xor ( n41252 , n41249 , n41250 );
xor ( n41253 , n40594 , n41204 );
and ( n41254 , n29904 , n41222 );
and ( n41255 , n41253 , n41254 );
xor ( n41256 , n41253 , n41254 );
xor ( n41257 , n40598 , n41202 );
and ( n41258 , n29909 , n41222 );
and ( n41259 , n41257 , n41258 );
xor ( n41260 , n41257 , n41258 );
xor ( n41261 , n40602 , n41200 );
and ( n41262 , n29914 , n41222 );
and ( n41263 , n41261 , n41262 );
xor ( n41264 , n41261 , n41262 );
xor ( n41265 , n40606 , n41198 );
and ( n41266 , n29919 , n41222 );
and ( n41267 , n41265 , n41266 );
xor ( n41268 , n41265 , n41266 );
xor ( n41269 , n40610 , n41196 );
and ( n41270 , n29924 , n41222 );
and ( n41271 , n41269 , n41270 );
xor ( n41272 , n41269 , n41270 );
xor ( n41273 , n40614 , n41194 );
and ( n41274 , n29929 , n41222 );
and ( n41275 , n41273 , n41274 );
xor ( n41276 , n41273 , n41274 );
xor ( n41277 , n40618 , n41192 );
and ( n41278 , n29934 , n41222 );
and ( n41279 , n41277 , n41278 );
xor ( n41280 , n41277 , n41278 );
xor ( n41281 , n40622 , n41190 );
and ( n41282 , n29939 , n41222 );
and ( n41283 , n41281 , n41282 );
xor ( n41284 , n41281 , n41282 );
xor ( n41285 , n40626 , n41188 );
and ( n41286 , n29944 , n41222 );
and ( n41287 , n41285 , n41286 );
xor ( n41288 , n41285 , n41286 );
xor ( n41289 , n40630 , n41186 );
and ( n41290 , n29949 , n41222 );
and ( n41291 , n41289 , n41290 );
xor ( n41292 , n41289 , n41290 );
xor ( n41293 , n40634 , n41184 );
and ( n41294 , n29954 , n41222 );
and ( n41295 , n41293 , n41294 );
xor ( n41296 , n41293 , n41294 );
xor ( n41297 , n40638 , n41182 );
and ( n41298 , n29959 , n41222 );
and ( n41299 , n41297 , n41298 );
xor ( n41300 , n41297 , n41298 );
xor ( n41301 , n40642 , n41180 );
and ( n41302 , n29964 , n41222 );
and ( n41303 , n41301 , n41302 );
xor ( n41304 , n41301 , n41302 );
xor ( n41305 , n40646 , n41178 );
and ( n41306 , n29969 , n41222 );
and ( n41307 , n41305 , n41306 );
xor ( n41308 , n41305 , n41306 );
xor ( n41309 , n40650 , n41176 );
and ( n41310 , n29974 , n41222 );
and ( n41311 , n41309 , n41310 );
xor ( n41312 , n41309 , n41310 );
xor ( n41313 , n40654 , n41174 );
and ( n41314 , n29979 , n41222 );
and ( n41315 , n41313 , n41314 );
xor ( n41316 , n41313 , n41314 );
xor ( n41317 , n40658 , n41172 );
and ( n41318 , n29984 , n41222 );
and ( n41319 , n41317 , n41318 );
xor ( n41320 , n41317 , n41318 );
xor ( n41321 , n40662 , n41170 );
and ( n41322 , n29989 , n41222 );
and ( n41323 , n41321 , n41322 );
xor ( n41324 , n41321 , n41322 );
xor ( n41325 , n40666 , n41168 );
and ( n41326 , n29994 , n41222 );
and ( n41327 , n41325 , n41326 );
xor ( n41328 , n41325 , n41326 );
xor ( n41329 , n40670 , n41166 );
and ( n41330 , n29999 , n41222 );
and ( n41331 , n41329 , n41330 );
xor ( n41332 , n41329 , n41330 );
xor ( n41333 , n40674 , n41164 );
and ( n41334 , n30004 , n41222 );
and ( n41335 , n41333 , n41334 );
xor ( n41336 , n41333 , n41334 );
xor ( n41337 , n40678 , n41162 );
and ( n41338 , n30009 , n41222 );
and ( n41339 , n41337 , n41338 );
xor ( n41340 , n41337 , n41338 );
xor ( n41341 , n40682 , n41160 );
and ( n41342 , n30014 , n41222 );
and ( n41343 , n41341 , n41342 );
xor ( n41344 , n41341 , n41342 );
xor ( n41345 , n40686 , n41158 );
and ( n41346 , n30019 , n41222 );
and ( n41347 , n41345 , n41346 );
xor ( n41348 , n41345 , n41346 );
xor ( n41349 , n40690 , n41156 );
and ( n41350 , n30024 , n41222 );
and ( n41351 , n41349 , n41350 );
xor ( n41352 , n41349 , n41350 );
xor ( n41353 , n40694 , n41154 );
and ( n41354 , n30029 , n41222 );
and ( n41355 , n41353 , n41354 );
xor ( n41356 , n41353 , n41354 );
xor ( n41357 , n40698 , n41152 );
and ( n41358 , n30034 , n41222 );
and ( n41359 , n41357 , n41358 );
xor ( n41360 , n41357 , n41358 );
xor ( n41361 , n40702 , n41150 );
and ( n41362 , n30039 , n41222 );
and ( n41363 , n41361 , n41362 );
xor ( n41364 , n41361 , n41362 );
xor ( n41365 , n40706 , n41148 );
and ( n41366 , n30044 , n41222 );
and ( n41367 , n41365 , n41366 );
xor ( n41368 , n41365 , n41366 );
xor ( n41369 , n40710 , n41146 );
and ( n41370 , n30049 , n41222 );
and ( n41371 , n41369 , n41370 );
xor ( n41372 , n41369 , n41370 );
xor ( n41373 , n40714 , n41144 );
and ( n41374 , n30054 , n41222 );
and ( n41375 , n41373 , n41374 );
xor ( n41376 , n41373 , n41374 );
xor ( n41377 , n40718 , n41142 );
and ( n41378 , n30059 , n41222 );
and ( n41379 , n41377 , n41378 );
xor ( n41380 , n41377 , n41378 );
xor ( n41381 , n40722 , n41140 );
and ( n41382 , n30064 , n41222 );
and ( n41383 , n41381 , n41382 );
xor ( n41384 , n41381 , n41382 );
xor ( n41385 , n40726 , n41138 );
and ( n41386 , n30069 , n41222 );
and ( n41387 , n41385 , n41386 );
xor ( n41388 , n41385 , n41386 );
xor ( n41389 , n40730 , n41136 );
and ( n41390 , n30074 , n41222 );
and ( n41391 , n41389 , n41390 );
xor ( n41392 , n41389 , n41390 );
xor ( n41393 , n40734 , n41134 );
and ( n41394 , n30079 , n41222 );
and ( n41395 , n41393 , n41394 );
xor ( n41396 , n41393 , n41394 );
xor ( n41397 , n40738 , n41132 );
and ( n41398 , n30084 , n41222 );
and ( n41399 , n41397 , n41398 );
xor ( n41400 , n41397 , n41398 );
xor ( n41401 , n40742 , n41130 );
and ( n41402 , n30089 , n41222 );
and ( n41403 , n41401 , n41402 );
xor ( n41404 , n41401 , n41402 );
xor ( n41405 , n40746 , n41128 );
and ( n41406 , n30094 , n41222 );
and ( n41407 , n41405 , n41406 );
xor ( n41408 , n41405 , n41406 );
xor ( n41409 , n40750 , n41126 );
and ( n41410 , n30099 , n41222 );
and ( n41411 , n41409 , n41410 );
xor ( n41412 , n41409 , n41410 );
xor ( n41413 , n40754 , n41124 );
and ( n41414 , n30104 , n41222 );
and ( n41415 , n41413 , n41414 );
xor ( n41416 , n41413 , n41414 );
xor ( n41417 , n40758 , n41122 );
and ( n41418 , n30109 , n41222 );
and ( n41419 , n41417 , n41418 );
xor ( n41420 , n41417 , n41418 );
xor ( n41421 , n40762 , n41120 );
and ( n41422 , n30114 , n41222 );
and ( n41423 , n41421 , n41422 );
xor ( n41424 , n41421 , n41422 );
xor ( n41425 , n40766 , n41118 );
and ( n41426 , n30119 , n41222 );
and ( n41427 , n41425 , n41426 );
xor ( n41428 , n41425 , n41426 );
xor ( n41429 , n40770 , n41116 );
and ( n41430 , n30124 , n41222 );
and ( n41431 , n41429 , n41430 );
xor ( n41432 , n41429 , n41430 );
xor ( n41433 , n40774 , n41114 );
and ( n41434 , n30129 , n41222 );
and ( n41435 , n41433 , n41434 );
xor ( n41436 , n41433 , n41434 );
xor ( n41437 , n40778 , n41112 );
and ( n41438 , n30134 , n41222 );
and ( n41439 , n41437 , n41438 );
xor ( n41440 , n41437 , n41438 );
xor ( n41441 , n40782 , n41110 );
and ( n41442 , n30139 , n41222 );
and ( n41443 , n41441 , n41442 );
xor ( n41444 , n41441 , n41442 );
xor ( n41445 , n40786 , n41108 );
and ( n41446 , n30144 , n41222 );
and ( n41447 , n41445 , n41446 );
xor ( n41448 , n41445 , n41446 );
xor ( n41449 , n40790 , n41106 );
and ( n41450 , n30149 , n41222 );
and ( n41451 , n41449 , n41450 );
xor ( n41452 , n41449 , n41450 );
xor ( n41453 , n40794 , n41104 );
and ( n41454 , n30154 , n41222 );
and ( n41455 , n41453 , n41454 );
xor ( n41456 , n41453 , n41454 );
xor ( n41457 , n40798 , n41102 );
and ( n41458 , n30159 , n41222 );
and ( n41459 , n41457 , n41458 );
xor ( n41460 , n41457 , n41458 );
xor ( n41461 , n40802 , n41100 );
and ( n41462 , n30164 , n41222 );
and ( n41463 , n41461 , n41462 );
xor ( n41464 , n41461 , n41462 );
xor ( n41465 , n40806 , n41098 );
and ( n41466 , n30169 , n41222 );
and ( n41467 , n41465 , n41466 );
xor ( n41468 , n41465 , n41466 );
xor ( n41469 , n40810 , n41096 );
and ( n41470 , n30174 , n41222 );
and ( n41471 , n41469 , n41470 );
xor ( n41472 , n41469 , n41470 );
xor ( n41473 , n40814 , n41094 );
and ( n41474 , n30179 , n41222 );
and ( n41475 , n41473 , n41474 );
xor ( n41476 , n41473 , n41474 );
xor ( n41477 , n40818 , n41092 );
and ( n41478 , n30184 , n41222 );
and ( n41479 , n41477 , n41478 );
xor ( n41480 , n41477 , n41478 );
xor ( n41481 , n40822 , n41090 );
and ( n41482 , n30189 , n41222 );
and ( n41483 , n41481 , n41482 );
xor ( n41484 , n41481 , n41482 );
xor ( n41485 , n40826 , n41088 );
and ( n41486 , n30194 , n41222 );
and ( n41487 , n41485 , n41486 );
xor ( n41488 , n41485 , n41486 );
xor ( n41489 , n40830 , n41086 );
and ( n41490 , n30199 , n41222 );
and ( n41491 , n41489 , n41490 );
xor ( n41492 , n41489 , n41490 );
xor ( n41493 , n40834 , n41084 );
and ( n41494 , n30204 , n41222 );
and ( n41495 , n41493 , n41494 );
xor ( n41496 , n41493 , n41494 );
xor ( n41497 , n40838 , n41082 );
and ( n41498 , n30209 , n41222 );
and ( n41499 , n41497 , n41498 );
xor ( n41500 , n41497 , n41498 );
xor ( n41501 , n40842 , n41080 );
and ( n41502 , n30214 , n41222 );
and ( n41503 , n41501 , n41502 );
xor ( n41504 , n41501 , n41502 );
xor ( n41505 , n40846 , n41078 );
and ( n41506 , n30219 , n41222 );
and ( n41507 , n41505 , n41506 );
xor ( n41508 , n41505 , n41506 );
xor ( n41509 , n40850 , n41076 );
and ( n41510 , n30224 , n41222 );
and ( n41511 , n41509 , n41510 );
xor ( n41512 , n41509 , n41510 );
xor ( n41513 , n40854 , n41074 );
and ( n41514 , n30229 , n41222 );
and ( n41515 , n41513 , n41514 );
xor ( n41516 , n41513 , n41514 );
xor ( n41517 , n40858 , n41072 );
and ( n41518 , n30234 , n41222 );
and ( n41519 , n41517 , n41518 );
xor ( n41520 , n41517 , n41518 );
xor ( n41521 , n40862 , n41070 );
and ( n41522 , n30239 , n41222 );
and ( n41523 , n41521 , n41522 );
xor ( n41524 , n41521 , n41522 );
xor ( n41525 , n40866 , n41068 );
and ( n41526 , n30244 , n41222 );
and ( n41527 , n41525 , n41526 );
xor ( n41528 , n41525 , n41526 );
xor ( n41529 , n40870 , n41066 );
and ( n41530 , n30249 , n41222 );
and ( n41531 , n41529 , n41530 );
xor ( n41532 , n41529 , n41530 );
xor ( n41533 , n40874 , n41064 );
and ( n41534 , n30254 , n41222 );
and ( n41535 , n41533 , n41534 );
xor ( n41536 , n41533 , n41534 );
xor ( n41537 , n40878 , n41062 );
and ( n41538 , n30259 , n41222 );
and ( n41539 , n41537 , n41538 );
xor ( n41540 , n41537 , n41538 );
xor ( n41541 , n40882 , n41060 );
and ( n41542 , n30264 , n41222 );
and ( n41543 , n41541 , n41542 );
xor ( n41544 , n41541 , n41542 );
xor ( n41545 , n40886 , n41058 );
and ( n41546 , n30269 , n41222 );
and ( n41547 , n41545 , n41546 );
xor ( n41548 , n41545 , n41546 );
xor ( n41549 , n40890 , n41056 );
and ( n41550 , n30274 , n41222 );
and ( n41551 , n41549 , n41550 );
xor ( n41552 , n41549 , n41550 );
xor ( n41553 , n40894 , n41054 );
and ( n41554 , n30279 , n41222 );
and ( n41555 , n41553 , n41554 );
xor ( n41556 , n41553 , n41554 );
xor ( n41557 , n40898 , n41052 );
and ( n41558 , n30284 , n41222 );
and ( n41559 , n41557 , n41558 );
xor ( n41560 , n41557 , n41558 );
xor ( n41561 , n40902 , n41050 );
and ( n41562 , n30289 , n41222 );
and ( n41563 , n41561 , n41562 );
xor ( n41564 , n41561 , n41562 );
xor ( n41565 , n40906 , n41048 );
and ( n41566 , n30294 , n41222 );
and ( n41567 , n41565 , n41566 );
xor ( n41568 , n41565 , n41566 );
xor ( n41569 , n40910 , n41046 );
and ( n41570 , n30299 , n41222 );
and ( n41571 , n41569 , n41570 );
xor ( n41572 , n41569 , n41570 );
xor ( n41573 , n40914 , n41044 );
and ( n41574 , n30304 , n41222 );
and ( n41575 , n41573 , n41574 );
xor ( n41576 , n41573 , n41574 );
xor ( n41577 , n40918 , n41042 );
and ( n41578 , n30309 , n41222 );
and ( n41579 , n41577 , n41578 );
xor ( n41580 , n41577 , n41578 );
xor ( n41581 , n40922 , n41040 );
and ( n41582 , n30314 , n41222 );
and ( n41583 , n41581 , n41582 );
xor ( n41584 , n41581 , n41582 );
xor ( n41585 , n40926 , n41038 );
and ( n41586 , n30319 , n41222 );
and ( n41587 , n41585 , n41586 );
xor ( n41588 , n41585 , n41586 );
xor ( n41589 , n40930 , n41036 );
and ( n41590 , n30324 , n41222 );
and ( n41591 , n41589 , n41590 );
xor ( n41592 , n41589 , n41590 );
xor ( n41593 , n40934 , n41034 );
and ( n41594 , n30329 , n41222 );
and ( n41595 , n41593 , n41594 );
xor ( n41596 , n41593 , n41594 );
xor ( n41597 , n40938 , n41032 );
and ( n41598 , n30334 , n41222 );
and ( n41599 , n41597 , n41598 );
xor ( n41600 , n41597 , n41598 );
xor ( n41601 , n40942 , n41030 );
and ( n41602 , n30339 , n41222 );
and ( n41603 , n41601 , n41602 );
xor ( n41604 , n41601 , n41602 );
xor ( n41605 , n40946 , n41028 );
and ( n41606 , n30344 , n41222 );
and ( n41607 , n41605 , n41606 );
xor ( n41608 , n41605 , n41606 );
xor ( n41609 , n40950 , n41026 );
and ( n41610 , n30349 , n41222 );
and ( n41611 , n41609 , n41610 );
xor ( n41612 , n41609 , n41610 );
xor ( n41613 , n40954 , n41024 );
and ( n41614 , n30354 , n41222 );
and ( n41615 , n41613 , n41614 );
xor ( n41616 , n41613 , n41614 );
xor ( n41617 , n40958 , n41022 );
and ( n41618 , n30359 , n41222 );
and ( n41619 , n41617 , n41618 );
xor ( n41620 , n41617 , n41618 );
xor ( n41621 , n40962 , n41020 );
and ( n41622 , n30364 , n41222 );
and ( n41623 , n41621 , n41622 );
xor ( n41624 , n41621 , n41622 );
xor ( n41625 , n40966 , n41018 );
and ( n41626 , n30369 , n41222 );
and ( n41627 , n41625 , n41626 );
xor ( n41628 , n41625 , n41626 );
xor ( n41629 , n40970 , n41016 );
and ( n41630 , n30374 , n41222 );
and ( n41631 , n41629 , n41630 );
xor ( n41632 , n41629 , n41630 );
xor ( n41633 , n40974 , n41014 );
and ( n41634 , n30379 , n41222 );
and ( n41635 , n41633 , n41634 );
xor ( n41636 , n41633 , n41634 );
xor ( n41637 , n40978 , n41012 );
and ( n41638 , n30384 , n41222 );
and ( n41639 , n41637 , n41638 );
xor ( n41640 , n41637 , n41638 );
xor ( n41641 , n40982 , n41010 );
and ( n41642 , n30389 , n41222 );
and ( n41643 , n41641 , n41642 );
xor ( n41644 , n41641 , n41642 );
xor ( n41645 , n40986 , n41008 );
and ( n41646 , n30394 , n41222 );
and ( n41647 , n41645 , n41646 );
xor ( n41648 , n41645 , n41646 );
xor ( n41649 , n40990 , n41006 );
and ( n41650 , n30399 , n41222 );
and ( n41651 , n41649 , n41650 );
xor ( n41652 , n41649 , n41650 );
xor ( n41653 , n40994 , n41004 );
and ( n41654 , n30404 , n41222 );
and ( n41655 , n41653 , n41654 );
xor ( n41656 , n41653 , n41654 );
xor ( n41657 , n40998 , n41002 );
and ( n41658 , n30409 , n41222 );
and ( n41659 , n41657 , n41658 );
buf ( n41660 , n41659 );
and ( n41661 , n41656 , n41660 );
or ( n41662 , n41655 , n41661 );
and ( n41663 , n41652 , n41662 );
or ( n41664 , n41651 , n41663 );
and ( n41665 , n41648 , n41664 );
or ( n41666 , n41647 , n41665 );
and ( n41667 , n41644 , n41666 );
or ( n41668 , n41643 , n41667 );
and ( n41669 , n41640 , n41668 );
or ( n41670 , n41639 , n41669 );
and ( n41671 , n41636 , n41670 );
or ( n41672 , n41635 , n41671 );
and ( n41673 , n41632 , n41672 );
or ( n41674 , n41631 , n41673 );
and ( n41675 , n41628 , n41674 );
or ( n41676 , n41627 , n41675 );
and ( n41677 , n41624 , n41676 );
or ( n41678 , n41623 , n41677 );
and ( n41679 , n41620 , n41678 );
or ( n41680 , n41619 , n41679 );
and ( n41681 , n41616 , n41680 );
or ( n41682 , n41615 , n41681 );
and ( n41683 , n41612 , n41682 );
or ( n41684 , n41611 , n41683 );
and ( n41685 , n41608 , n41684 );
or ( n41686 , n41607 , n41685 );
and ( n41687 , n41604 , n41686 );
or ( n41688 , n41603 , n41687 );
and ( n41689 , n41600 , n41688 );
or ( n41690 , n41599 , n41689 );
and ( n41691 , n41596 , n41690 );
or ( n41692 , n41595 , n41691 );
and ( n41693 , n41592 , n41692 );
or ( n41694 , n41591 , n41693 );
and ( n41695 , n41588 , n41694 );
or ( n41696 , n41587 , n41695 );
and ( n41697 , n41584 , n41696 );
or ( n41698 , n41583 , n41697 );
and ( n41699 , n41580 , n41698 );
or ( n41700 , n41579 , n41699 );
and ( n41701 , n41576 , n41700 );
or ( n41702 , n41575 , n41701 );
and ( n41703 , n41572 , n41702 );
or ( n41704 , n41571 , n41703 );
and ( n41705 , n41568 , n41704 );
or ( n41706 , n41567 , n41705 );
and ( n41707 , n41564 , n41706 );
or ( n41708 , n41563 , n41707 );
and ( n41709 , n41560 , n41708 );
or ( n41710 , n41559 , n41709 );
and ( n41711 , n41556 , n41710 );
or ( n41712 , n41555 , n41711 );
and ( n41713 , n41552 , n41712 );
or ( n41714 , n41551 , n41713 );
and ( n41715 , n41548 , n41714 );
or ( n41716 , n41547 , n41715 );
and ( n41717 , n41544 , n41716 );
or ( n41718 , n41543 , n41717 );
and ( n41719 , n41540 , n41718 );
or ( n41720 , n41539 , n41719 );
and ( n41721 , n41536 , n41720 );
or ( n41722 , n41535 , n41721 );
and ( n41723 , n41532 , n41722 );
or ( n41724 , n41531 , n41723 );
and ( n41725 , n41528 , n41724 );
or ( n41726 , n41527 , n41725 );
and ( n41727 , n41524 , n41726 );
or ( n41728 , n41523 , n41727 );
and ( n41729 , n41520 , n41728 );
or ( n41730 , n41519 , n41729 );
and ( n41731 , n41516 , n41730 );
or ( n41732 , n41515 , n41731 );
and ( n41733 , n41512 , n41732 );
or ( n41734 , n41511 , n41733 );
and ( n41735 , n41508 , n41734 );
or ( n41736 , n41507 , n41735 );
and ( n41737 , n41504 , n41736 );
or ( n41738 , n41503 , n41737 );
and ( n41739 , n41500 , n41738 );
or ( n41740 , n41499 , n41739 );
and ( n41741 , n41496 , n41740 );
or ( n41742 , n41495 , n41741 );
and ( n41743 , n41492 , n41742 );
or ( n41744 , n41491 , n41743 );
and ( n41745 , n41488 , n41744 );
or ( n41746 , n41487 , n41745 );
and ( n41747 , n41484 , n41746 );
or ( n41748 , n41483 , n41747 );
and ( n41749 , n41480 , n41748 );
or ( n41750 , n41479 , n41749 );
and ( n41751 , n41476 , n41750 );
or ( n41752 , n41475 , n41751 );
and ( n41753 , n41472 , n41752 );
or ( n41754 , n41471 , n41753 );
and ( n41755 , n41468 , n41754 );
or ( n41756 , n41467 , n41755 );
and ( n41757 , n41464 , n41756 );
or ( n41758 , n41463 , n41757 );
and ( n41759 , n41460 , n41758 );
or ( n41760 , n41459 , n41759 );
and ( n41761 , n41456 , n41760 );
or ( n41762 , n41455 , n41761 );
and ( n41763 , n41452 , n41762 );
or ( n41764 , n41451 , n41763 );
and ( n41765 , n41448 , n41764 );
or ( n41766 , n41447 , n41765 );
and ( n41767 , n41444 , n41766 );
or ( n41768 , n41443 , n41767 );
and ( n41769 , n41440 , n41768 );
or ( n41770 , n41439 , n41769 );
and ( n41771 , n41436 , n41770 );
or ( n41772 , n41435 , n41771 );
and ( n41773 , n41432 , n41772 );
or ( n41774 , n41431 , n41773 );
and ( n41775 , n41428 , n41774 );
or ( n41776 , n41427 , n41775 );
and ( n41777 , n41424 , n41776 );
or ( n41778 , n41423 , n41777 );
and ( n41779 , n41420 , n41778 );
or ( n41780 , n41419 , n41779 );
and ( n41781 , n41416 , n41780 );
or ( n41782 , n41415 , n41781 );
and ( n41783 , n41412 , n41782 );
or ( n41784 , n41411 , n41783 );
and ( n41785 , n41408 , n41784 );
or ( n41786 , n41407 , n41785 );
and ( n41787 , n41404 , n41786 );
or ( n41788 , n41403 , n41787 );
and ( n41789 , n41400 , n41788 );
or ( n41790 , n41399 , n41789 );
and ( n41791 , n41396 , n41790 );
or ( n41792 , n41395 , n41791 );
and ( n41793 , n41392 , n41792 );
or ( n41794 , n41391 , n41793 );
and ( n41795 , n41388 , n41794 );
or ( n41796 , n41387 , n41795 );
and ( n41797 , n41384 , n41796 );
or ( n41798 , n41383 , n41797 );
and ( n41799 , n41380 , n41798 );
or ( n41800 , n41379 , n41799 );
and ( n41801 , n41376 , n41800 );
or ( n41802 , n41375 , n41801 );
and ( n41803 , n41372 , n41802 );
or ( n41804 , n41371 , n41803 );
and ( n41805 , n41368 , n41804 );
or ( n41806 , n41367 , n41805 );
and ( n41807 , n41364 , n41806 );
or ( n41808 , n41363 , n41807 );
and ( n41809 , n41360 , n41808 );
or ( n41810 , n41359 , n41809 );
and ( n41811 , n41356 , n41810 );
or ( n41812 , n41355 , n41811 );
and ( n41813 , n41352 , n41812 );
or ( n41814 , n41351 , n41813 );
and ( n41815 , n41348 , n41814 );
or ( n41816 , n41347 , n41815 );
and ( n41817 , n41344 , n41816 );
or ( n41818 , n41343 , n41817 );
and ( n41819 , n41340 , n41818 );
or ( n41820 , n41339 , n41819 );
and ( n41821 , n41336 , n41820 );
or ( n41822 , n41335 , n41821 );
and ( n41823 , n41332 , n41822 );
or ( n41824 , n41331 , n41823 );
and ( n41825 , n41328 , n41824 );
or ( n41826 , n41327 , n41825 );
and ( n41827 , n41324 , n41826 );
or ( n41828 , n41323 , n41827 );
and ( n41829 , n41320 , n41828 );
or ( n41830 , n41319 , n41829 );
and ( n41831 , n41316 , n41830 );
or ( n41832 , n41315 , n41831 );
and ( n41833 , n41312 , n41832 );
or ( n41834 , n41311 , n41833 );
and ( n41835 , n41308 , n41834 );
or ( n41836 , n41307 , n41835 );
and ( n41837 , n41304 , n41836 );
or ( n41838 , n41303 , n41837 );
and ( n41839 , n41300 , n41838 );
or ( n41840 , n41299 , n41839 );
and ( n41841 , n41296 , n41840 );
or ( n41842 , n41295 , n41841 );
and ( n41843 , n41292 , n41842 );
or ( n41844 , n41291 , n41843 );
and ( n41845 , n41288 , n41844 );
or ( n41846 , n41287 , n41845 );
and ( n41847 , n41284 , n41846 );
or ( n41848 , n41283 , n41847 );
and ( n41849 , n41280 , n41848 );
or ( n41850 , n41279 , n41849 );
and ( n41851 , n41276 , n41850 );
or ( n41852 , n41275 , n41851 );
and ( n41853 , n41272 , n41852 );
or ( n41854 , n41271 , n41853 );
and ( n41855 , n41268 , n41854 );
or ( n41856 , n41267 , n41855 );
and ( n41857 , n41264 , n41856 );
or ( n41858 , n41263 , n41857 );
and ( n41859 , n41260 , n41858 );
or ( n41860 , n41259 , n41859 );
and ( n41861 , n41256 , n41860 );
or ( n41862 , n41255 , n41861 );
and ( n41863 , n41252 , n41862 );
or ( n41864 , n41251 , n41863 );
and ( n41865 , n41248 , n41864 );
or ( n41866 , n41247 , n41865 );
and ( n41867 , n41244 , n41866 );
or ( n41868 , n41243 , n41867 );
and ( n41869 , n41240 , n41868 );
or ( n41870 , n41239 , n41869 );
and ( n41871 , n41236 , n41870 );
or ( n41872 , n41235 , n41871 );
and ( n41873 , n41232 , n41872 );
or ( n41874 , n41231 , n41873 );
and ( n41875 , n41228 , n41874 );
or ( n41876 , n41227 , n41875 );
xor ( n41877 , n41224 , n41876 );
buf ( n41878 , n18070 );
and ( n41879 , n29869 , n41878 );
xor ( n41880 , n41877 , n41879 );
xor ( n41881 , n41228 , n41874 );
and ( n41882 , n29874 , n41878 );
and ( n41883 , n41881 , n41882 );
xor ( n41884 , n41881 , n41882 );
xor ( n41885 , n41232 , n41872 );
and ( n41886 , n29879 , n41878 );
and ( n41887 , n41885 , n41886 );
xor ( n41888 , n41885 , n41886 );
xor ( n41889 , n41236 , n41870 );
and ( n41890 , n29884 , n41878 );
and ( n41891 , n41889 , n41890 );
xor ( n41892 , n41889 , n41890 );
xor ( n41893 , n41240 , n41868 );
and ( n41894 , n29889 , n41878 );
and ( n41895 , n41893 , n41894 );
xor ( n41896 , n41893 , n41894 );
xor ( n41897 , n41244 , n41866 );
and ( n41898 , n29894 , n41878 );
and ( n41899 , n41897 , n41898 );
xor ( n41900 , n41897 , n41898 );
xor ( n41901 , n41248 , n41864 );
and ( n41902 , n29899 , n41878 );
and ( n41903 , n41901 , n41902 );
xor ( n41904 , n41901 , n41902 );
xor ( n41905 , n41252 , n41862 );
and ( n41906 , n29904 , n41878 );
and ( n41907 , n41905 , n41906 );
xor ( n41908 , n41905 , n41906 );
xor ( n41909 , n41256 , n41860 );
and ( n41910 , n29909 , n41878 );
and ( n41911 , n41909 , n41910 );
xor ( n41912 , n41909 , n41910 );
xor ( n41913 , n41260 , n41858 );
and ( n41914 , n29914 , n41878 );
and ( n41915 , n41913 , n41914 );
xor ( n41916 , n41913 , n41914 );
xor ( n41917 , n41264 , n41856 );
and ( n41918 , n29919 , n41878 );
and ( n41919 , n41917 , n41918 );
xor ( n41920 , n41917 , n41918 );
xor ( n41921 , n41268 , n41854 );
and ( n41922 , n29924 , n41878 );
and ( n41923 , n41921 , n41922 );
xor ( n41924 , n41921 , n41922 );
xor ( n41925 , n41272 , n41852 );
and ( n41926 , n29929 , n41878 );
and ( n41927 , n41925 , n41926 );
xor ( n41928 , n41925 , n41926 );
xor ( n41929 , n41276 , n41850 );
and ( n41930 , n29934 , n41878 );
and ( n41931 , n41929 , n41930 );
xor ( n41932 , n41929 , n41930 );
xor ( n41933 , n41280 , n41848 );
and ( n41934 , n29939 , n41878 );
and ( n41935 , n41933 , n41934 );
xor ( n41936 , n41933 , n41934 );
xor ( n41937 , n41284 , n41846 );
and ( n41938 , n29944 , n41878 );
and ( n41939 , n41937 , n41938 );
xor ( n41940 , n41937 , n41938 );
xor ( n41941 , n41288 , n41844 );
and ( n41942 , n29949 , n41878 );
and ( n41943 , n41941 , n41942 );
xor ( n41944 , n41941 , n41942 );
xor ( n41945 , n41292 , n41842 );
and ( n41946 , n29954 , n41878 );
and ( n41947 , n41945 , n41946 );
xor ( n41948 , n41945 , n41946 );
xor ( n41949 , n41296 , n41840 );
and ( n41950 , n29959 , n41878 );
and ( n41951 , n41949 , n41950 );
xor ( n41952 , n41949 , n41950 );
xor ( n41953 , n41300 , n41838 );
and ( n41954 , n29964 , n41878 );
and ( n41955 , n41953 , n41954 );
xor ( n41956 , n41953 , n41954 );
xor ( n41957 , n41304 , n41836 );
and ( n41958 , n29969 , n41878 );
and ( n41959 , n41957 , n41958 );
xor ( n41960 , n41957 , n41958 );
xor ( n41961 , n41308 , n41834 );
and ( n41962 , n29974 , n41878 );
and ( n41963 , n41961 , n41962 );
xor ( n41964 , n41961 , n41962 );
xor ( n41965 , n41312 , n41832 );
and ( n41966 , n29979 , n41878 );
and ( n41967 , n41965 , n41966 );
xor ( n41968 , n41965 , n41966 );
xor ( n41969 , n41316 , n41830 );
and ( n41970 , n29984 , n41878 );
and ( n41971 , n41969 , n41970 );
xor ( n41972 , n41969 , n41970 );
xor ( n41973 , n41320 , n41828 );
and ( n41974 , n29989 , n41878 );
and ( n41975 , n41973 , n41974 );
xor ( n41976 , n41973 , n41974 );
xor ( n41977 , n41324 , n41826 );
and ( n41978 , n29994 , n41878 );
and ( n41979 , n41977 , n41978 );
xor ( n41980 , n41977 , n41978 );
xor ( n41981 , n41328 , n41824 );
and ( n41982 , n29999 , n41878 );
and ( n41983 , n41981 , n41982 );
xor ( n41984 , n41981 , n41982 );
xor ( n41985 , n41332 , n41822 );
and ( n41986 , n30004 , n41878 );
and ( n41987 , n41985 , n41986 );
xor ( n41988 , n41985 , n41986 );
xor ( n41989 , n41336 , n41820 );
and ( n41990 , n30009 , n41878 );
and ( n41991 , n41989 , n41990 );
xor ( n41992 , n41989 , n41990 );
xor ( n41993 , n41340 , n41818 );
and ( n41994 , n30014 , n41878 );
and ( n41995 , n41993 , n41994 );
xor ( n41996 , n41993 , n41994 );
xor ( n41997 , n41344 , n41816 );
and ( n41998 , n30019 , n41878 );
and ( n41999 , n41997 , n41998 );
xor ( n42000 , n41997 , n41998 );
xor ( n42001 , n41348 , n41814 );
and ( n42002 , n30024 , n41878 );
and ( n42003 , n42001 , n42002 );
xor ( n42004 , n42001 , n42002 );
xor ( n42005 , n41352 , n41812 );
and ( n42006 , n30029 , n41878 );
and ( n42007 , n42005 , n42006 );
xor ( n42008 , n42005 , n42006 );
xor ( n42009 , n41356 , n41810 );
and ( n42010 , n30034 , n41878 );
and ( n42011 , n42009 , n42010 );
xor ( n42012 , n42009 , n42010 );
xor ( n42013 , n41360 , n41808 );
and ( n42014 , n30039 , n41878 );
and ( n42015 , n42013 , n42014 );
xor ( n42016 , n42013 , n42014 );
xor ( n42017 , n41364 , n41806 );
and ( n42018 , n30044 , n41878 );
and ( n42019 , n42017 , n42018 );
xor ( n42020 , n42017 , n42018 );
xor ( n42021 , n41368 , n41804 );
and ( n42022 , n30049 , n41878 );
and ( n42023 , n42021 , n42022 );
xor ( n42024 , n42021 , n42022 );
xor ( n42025 , n41372 , n41802 );
and ( n42026 , n30054 , n41878 );
and ( n42027 , n42025 , n42026 );
xor ( n42028 , n42025 , n42026 );
xor ( n42029 , n41376 , n41800 );
and ( n42030 , n30059 , n41878 );
and ( n42031 , n42029 , n42030 );
xor ( n42032 , n42029 , n42030 );
xor ( n42033 , n41380 , n41798 );
and ( n42034 , n30064 , n41878 );
and ( n42035 , n42033 , n42034 );
xor ( n42036 , n42033 , n42034 );
xor ( n42037 , n41384 , n41796 );
and ( n42038 , n30069 , n41878 );
and ( n42039 , n42037 , n42038 );
xor ( n42040 , n42037 , n42038 );
xor ( n42041 , n41388 , n41794 );
and ( n42042 , n30074 , n41878 );
and ( n42043 , n42041 , n42042 );
xor ( n42044 , n42041 , n42042 );
xor ( n42045 , n41392 , n41792 );
and ( n42046 , n30079 , n41878 );
and ( n42047 , n42045 , n42046 );
xor ( n42048 , n42045 , n42046 );
xor ( n42049 , n41396 , n41790 );
and ( n42050 , n30084 , n41878 );
and ( n42051 , n42049 , n42050 );
xor ( n42052 , n42049 , n42050 );
xor ( n42053 , n41400 , n41788 );
and ( n42054 , n30089 , n41878 );
and ( n42055 , n42053 , n42054 );
xor ( n42056 , n42053 , n42054 );
xor ( n42057 , n41404 , n41786 );
and ( n42058 , n30094 , n41878 );
and ( n42059 , n42057 , n42058 );
xor ( n42060 , n42057 , n42058 );
xor ( n42061 , n41408 , n41784 );
and ( n42062 , n30099 , n41878 );
and ( n42063 , n42061 , n42062 );
xor ( n42064 , n42061 , n42062 );
xor ( n42065 , n41412 , n41782 );
and ( n42066 , n30104 , n41878 );
and ( n42067 , n42065 , n42066 );
xor ( n42068 , n42065 , n42066 );
xor ( n42069 , n41416 , n41780 );
and ( n42070 , n30109 , n41878 );
and ( n42071 , n42069 , n42070 );
xor ( n42072 , n42069 , n42070 );
xor ( n42073 , n41420 , n41778 );
and ( n42074 , n30114 , n41878 );
and ( n42075 , n42073 , n42074 );
xor ( n42076 , n42073 , n42074 );
xor ( n42077 , n41424 , n41776 );
and ( n42078 , n30119 , n41878 );
and ( n42079 , n42077 , n42078 );
xor ( n42080 , n42077 , n42078 );
xor ( n42081 , n41428 , n41774 );
and ( n42082 , n30124 , n41878 );
and ( n42083 , n42081 , n42082 );
xor ( n42084 , n42081 , n42082 );
xor ( n42085 , n41432 , n41772 );
and ( n42086 , n30129 , n41878 );
and ( n42087 , n42085 , n42086 );
xor ( n42088 , n42085 , n42086 );
xor ( n42089 , n41436 , n41770 );
and ( n42090 , n30134 , n41878 );
and ( n42091 , n42089 , n42090 );
xor ( n42092 , n42089 , n42090 );
xor ( n42093 , n41440 , n41768 );
and ( n42094 , n30139 , n41878 );
and ( n42095 , n42093 , n42094 );
xor ( n42096 , n42093 , n42094 );
xor ( n42097 , n41444 , n41766 );
and ( n42098 , n30144 , n41878 );
and ( n42099 , n42097 , n42098 );
xor ( n42100 , n42097 , n42098 );
xor ( n42101 , n41448 , n41764 );
and ( n42102 , n30149 , n41878 );
and ( n42103 , n42101 , n42102 );
xor ( n42104 , n42101 , n42102 );
xor ( n42105 , n41452 , n41762 );
and ( n42106 , n30154 , n41878 );
and ( n42107 , n42105 , n42106 );
xor ( n42108 , n42105 , n42106 );
xor ( n42109 , n41456 , n41760 );
and ( n42110 , n30159 , n41878 );
and ( n42111 , n42109 , n42110 );
xor ( n42112 , n42109 , n42110 );
xor ( n42113 , n41460 , n41758 );
and ( n42114 , n30164 , n41878 );
and ( n42115 , n42113 , n42114 );
xor ( n42116 , n42113 , n42114 );
xor ( n42117 , n41464 , n41756 );
and ( n42118 , n30169 , n41878 );
and ( n42119 , n42117 , n42118 );
xor ( n42120 , n42117 , n42118 );
xor ( n42121 , n41468 , n41754 );
and ( n42122 , n30174 , n41878 );
and ( n42123 , n42121 , n42122 );
xor ( n42124 , n42121 , n42122 );
xor ( n42125 , n41472 , n41752 );
and ( n42126 , n30179 , n41878 );
and ( n42127 , n42125 , n42126 );
xor ( n42128 , n42125 , n42126 );
xor ( n42129 , n41476 , n41750 );
and ( n42130 , n30184 , n41878 );
and ( n42131 , n42129 , n42130 );
xor ( n42132 , n42129 , n42130 );
xor ( n42133 , n41480 , n41748 );
and ( n42134 , n30189 , n41878 );
and ( n42135 , n42133 , n42134 );
xor ( n42136 , n42133 , n42134 );
xor ( n42137 , n41484 , n41746 );
and ( n42138 , n30194 , n41878 );
and ( n42139 , n42137 , n42138 );
xor ( n42140 , n42137 , n42138 );
xor ( n42141 , n41488 , n41744 );
and ( n42142 , n30199 , n41878 );
and ( n42143 , n42141 , n42142 );
xor ( n42144 , n42141 , n42142 );
xor ( n42145 , n41492 , n41742 );
and ( n42146 , n30204 , n41878 );
and ( n42147 , n42145 , n42146 );
xor ( n42148 , n42145 , n42146 );
xor ( n42149 , n41496 , n41740 );
and ( n42150 , n30209 , n41878 );
and ( n42151 , n42149 , n42150 );
xor ( n42152 , n42149 , n42150 );
xor ( n42153 , n41500 , n41738 );
and ( n42154 , n30214 , n41878 );
and ( n42155 , n42153 , n42154 );
xor ( n42156 , n42153 , n42154 );
xor ( n42157 , n41504 , n41736 );
and ( n42158 , n30219 , n41878 );
and ( n42159 , n42157 , n42158 );
xor ( n42160 , n42157 , n42158 );
xor ( n42161 , n41508 , n41734 );
and ( n42162 , n30224 , n41878 );
and ( n42163 , n42161 , n42162 );
xor ( n42164 , n42161 , n42162 );
xor ( n42165 , n41512 , n41732 );
and ( n42166 , n30229 , n41878 );
and ( n42167 , n42165 , n42166 );
xor ( n42168 , n42165 , n42166 );
xor ( n42169 , n41516 , n41730 );
and ( n42170 , n30234 , n41878 );
and ( n42171 , n42169 , n42170 );
xor ( n42172 , n42169 , n42170 );
xor ( n42173 , n41520 , n41728 );
and ( n42174 , n30239 , n41878 );
and ( n42175 , n42173 , n42174 );
xor ( n42176 , n42173 , n42174 );
xor ( n42177 , n41524 , n41726 );
and ( n42178 , n30244 , n41878 );
and ( n42179 , n42177 , n42178 );
xor ( n42180 , n42177 , n42178 );
xor ( n42181 , n41528 , n41724 );
and ( n42182 , n30249 , n41878 );
and ( n42183 , n42181 , n42182 );
xor ( n42184 , n42181 , n42182 );
xor ( n42185 , n41532 , n41722 );
and ( n42186 , n30254 , n41878 );
and ( n42187 , n42185 , n42186 );
xor ( n42188 , n42185 , n42186 );
xor ( n42189 , n41536 , n41720 );
and ( n42190 , n30259 , n41878 );
and ( n42191 , n42189 , n42190 );
xor ( n42192 , n42189 , n42190 );
xor ( n42193 , n41540 , n41718 );
and ( n42194 , n30264 , n41878 );
and ( n42195 , n42193 , n42194 );
xor ( n42196 , n42193 , n42194 );
xor ( n42197 , n41544 , n41716 );
and ( n42198 , n30269 , n41878 );
and ( n42199 , n42197 , n42198 );
xor ( n42200 , n42197 , n42198 );
xor ( n42201 , n41548 , n41714 );
and ( n42202 , n30274 , n41878 );
and ( n42203 , n42201 , n42202 );
xor ( n42204 , n42201 , n42202 );
xor ( n42205 , n41552 , n41712 );
and ( n42206 , n30279 , n41878 );
and ( n42207 , n42205 , n42206 );
xor ( n42208 , n42205 , n42206 );
xor ( n42209 , n41556 , n41710 );
and ( n42210 , n30284 , n41878 );
and ( n42211 , n42209 , n42210 );
xor ( n42212 , n42209 , n42210 );
xor ( n42213 , n41560 , n41708 );
and ( n42214 , n30289 , n41878 );
and ( n42215 , n42213 , n42214 );
xor ( n42216 , n42213 , n42214 );
xor ( n42217 , n41564 , n41706 );
and ( n42218 , n30294 , n41878 );
and ( n42219 , n42217 , n42218 );
xor ( n42220 , n42217 , n42218 );
xor ( n42221 , n41568 , n41704 );
and ( n42222 , n30299 , n41878 );
and ( n42223 , n42221 , n42222 );
xor ( n42224 , n42221 , n42222 );
xor ( n42225 , n41572 , n41702 );
and ( n42226 , n30304 , n41878 );
and ( n42227 , n42225 , n42226 );
xor ( n42228 , n42225 , n42226 );
xor ( n42229 , n41576 , n41700 );
and ( n42230 , n30309 , n41878 );
and ( n42231 , n42229 , n42230 );
xor ( n42232 , n42229 , n42230 );
xor ( n42233 , n41580 , n41698 );
and ( n42234 , n30314 , n41878 );
and ( n42235 , n42233 , n42234 );
xor ( n42236 , n42233 , n42234 );
xor ( n42237 , n41584 , n41696 );
and ( n42238 , n30319 , n41878 );
and ( n42239 , n42237 , n42238 );
xor ( n42240 , n42237 , n42238 );
xor ( n42241 , n41588 , n41694 );
and ( n42242 , n30324 , n41878 );
and ( n42243 , n42241 , n42242 );
xor ( n42244 , n42241 , n42242 );
xor ( n42245 , n41592 , n41692 );
and ( n42246 , n30329 , n41878 );
and ( n42247 , n42245 , n42246 );
xor ( n42248 , n42245 , n42246 );
xor ( n42249 , n41596 , n41690 );
and ( n42250 , n30334 , n41878 );
and ( n42251 , n42249 , n42250 );
xor ( n42252 , n42249 , n42250 );
xor ( n42253 , n41600 , n41688 );
and ( n42254 , n30339 , n41878 );
and ( n42255 , n42253 , n42254 );
xor ( n42256 , n42253 , n42254 );
xor ( n42257 , n41604 , n41686 );
and ( n42258 , n30344 , n41878 );
and ( n42259 , n42257 , n42258 );
xor ( n42260 , n42257 , n42258 );
xor ( n42261 , n41608 , n41684 );
and ( n42262 , n30349 , n41878 );
and ( n42263 , n42261 , n42262 );
xor ( n42264 , n42261 , n42262 );
xor ( n42265 , n41612 , n41682 );
and ( n42266 , n30354 , n41878 );
and ( n42267 , n42265 , n42266 );
xor ( n42268 , n42265 , n42266 );
xor ( n42269 , n41616 , n41680 );
and ( n42270 , n30359 , n41878 );
and ( n42271 , n42269 , n42270 );
xor ( n42272 , n42269 , n42270 );
xor ( n42273 , n41620 , n41678 );
and ( n42274 , n30364 , n41878 );
and ( n42275 , n42273 , n42274 );
xor ( n42276 , n42273 , n42274 );
xor ( n42277 , n41624 , n41676 );
and ( n42278 , n30369 , n41878 );
and ( n42279 , n42277 , n42278 );
xor ( n42280 , n42277 , n42278 );
xor ( n42281 , n41628 , n41674 );
and ( n42282 , n30374 , n41878 );
and ( n42283 , n42281 , n42282 );
xor ( n42284 , n42281 , n42282 );
xor ( n42285 , n41632 , n41672 );
and ( n42286 , n30379 , n41878 );
and ( n42287 , n42285 , n42286 );
xor ( n42288 , n42285 , n42286 );
xor ( n42289 , n41636 , n41670 );
and ( n42290 , n30384 , n41878 );
and ( n42291 , n42289 , n42290 );
xor ( n42292 , n42289 , n42290 );
xor ( n42293 , n41640 , n41668 );
and ( n42294 , n30389 , n41878 );
and ( n42295 , n42293 , n42294 );
xor ( n42296 , n42293 , n42294 );
xor ( n42297 , n41644 , n41666 );
and ( n42298 , n30394 , n41878 );
and ( n42299 , n42297 , n42298 );
xor ( n42300 , n42297 , n42298 );
xor ( n42301 , n41648 , n41664 );
and ( n42302 , n30399 , n41878 );
and ( n42303 , n42301 , n42302 );
xor ( n42304 , n42301 , n42302 );
xor ( n42305 , n41652 , n41662 );
and ( n42306 , n30404 , n41878 );
and ( n42307 , n42305 , n42306 );
xor ( n42308 , n42305 , n42306 );
xor ( n42309 , n41656 , n41660 );
and ( n42310 , n30409 , n41878 );
and ( n42311 , n42309 , n42310 );
buf ( n42312 , n42311 );
and ( n42313 , n42308 , n42312 );
or ( n42314 , n42307 , n42313 );
and ( n42315 , n42304 , n42314 );
or ( n42316 , n42303 , n42315 );
and ( n42317 , n42300 , n42316 );
or ( n42318 , n42299 , n42317 );
and ( n42319 , n42296 , n42318 );
or ( n42320 , n42295 , n42319 );
and ( n42321 , n42292 , n42320 );
or ( n42322 , n42291 , n42321 );
and ( n42323 , n42288 , n42322 );
or ( n42324 , n42287 , n42323 );
and ( n42325 , n42284 , n42324 );
or ( n42326 , n42283 , n42325 );
and ( n42327 , n42280 , n42326 );
or ( n42328 , n42279 , n42327 );
and ( n42329 , n42276 , n42328 );
or ( n42330 , n42275 , n42329 );
and ( n42331 , n42272 , n42330 );
or ( n42332 , n42271 , n42331 );
and ( n42333 , n42268 , n42332 );
or ( n42334 , n42267 , n42333 );
and ( n42335 , n42264 , n42334 );
or ( n42336 , n42263 , n42335 );
and ( n42337 , n42260 , n42336 );
or ( n42338 , n42259 , n42337 );
and ( n42339 , n42256 , n42338 );
or ( n42340 , n42255 , n42339 );
and ( n42341 , n42252 , n42340 );
or ( n42342 , n42251 , n42341 );
and ( n42343 , n42248 , n42342 );
or ( n42344 , n42247 , n42343 );
and ( n42345 , n42244 , n42344 );
or ( n42346 , n42243 , n42345 );
and ( n42347 , n42240 , n42346 );
or ( n42348 , n42239 , n42347 );
and ( n42349 , n42236 , n42348 );
or ( n42350 , n42235 , n42349 );
and ( n42351 , n42232 , n42350 );
or ( n42352 , n42231 , n42351 );
and ( n42353 , n42228 , n42352 );
or ( n42354 , n42227 , n42353 );
and ( n42355 , n42224 , n42354 );
or ( n42356 , n42223 , n42355 );
and ( n42357 , n42220 , n42356 );
or ( n42358 , n42219 , n42357 );
and ( n42359 , n42216 , n42358 );
or ( n42360 , n42215 , n42359 );
and ( n42361 , n42212 , n42360 );
or ( n42362 , n42211 , n42361 );
and ( n42363 , n42208 , n42362 );
or ( n42364 , n42207 , n42363 );
and ( n42365 , n42204 , n42364 );
or ( n42366 , n42203 , n42365 );
and ( n42367 , n42200 , n42366 );
or ( n42368 , n42199 , n42367 );
and ( n42369 , n42196 , n42368 );
or ( n42370 , n42195 , n42369 );
and ( n42371 , n42192 , n42370 );
or ( n42372 , n42191 , n42371 );
and ( n42373 , n42188 , n42372 );
or ( n42374 , n42187 , n42373 );
and ( n42375 , n42184 , n42374 );
or ( n42376 , n42183 , n42375 );
and ( n42377 , n42180 , n42376 );
or ( n42378 , n42179 , n42377 );
and ( n42379 , n42176 , n42378 );
or ( n42380 , n42175 , n42379 );
and ( n42381 , n42172 , n42380 );
or ( n42382 , n42171 , n42381 );
and ( n42383 , n42168 , n42382 );
or ( n42384 , n42167 , n42383 );
and ( n42385 , n42164 , n42384 );
or ( n42386 , n42163 , n42385 );
and ( n42387 , n42160 , n42386 );
or ( n42388 , n42159 , n42387 );
and ( n42389 , n42156 , n42388 );
or ( n42390 , n42155 , n42389 );
and ( n42391 , n42152 , n42390 );
or ( n42392 , n42151 , n42391 );
and ( n42393 , n42148 , n42392 );
or ( n42394 , n42147 , n42393 );
and ( n42395 , n42144 , n42394 );
or ( n42396 , n42143 , n42395 );
and ( n42397 , n42140 , n42396 );
or ( n42398 , n42139 , n42397 );
and ( n42399 , n42136 , n42398 );
or ( n42400 , n42135 , n42399 );
and ( n42401 , n42132 , n42400 );
or ( n42402 , n42131 , n42401 );
and ( n42403 , n42128 , n42402 );
or ( n42404 , n42127 , n42403 );
and ( n42405 , n42124 , n42404 );
or ( n42406 , n42123 , n42405 );
and ( n42407 , n42120 , n42406 );
or ( n42408 , n42119 , n42407 );
and ( n42409 , n42116 , n42408 );
or ( n42410 , n42115 , n42409 );
and ( n42411 , n42112 , n42410 );
or ( n42412 , n42111 , n42411 );
and ( n42413 , n42108 , n42412 );
or ( n42414 , n42107 , n42413 );
and ( n42415 , n42104 , n42414 );
or ( n42416 , n42103 , n42415 );
and ( n42417 , n42100 , n42416 );
or ( n42418 , n42099 , n42417 );
and ( n42419 , n42096 , n42418 );
or ( n42420 , n42095 , n42419 );
and ( n42421 , n42092 , n42420 );
or ( n42422 , n42091 , n42421 );
and ( n42423 , n42088 , n42422 );
or ( n42424 , n42087 , n42423 );
and ( n42425 , n42084 , n42424 );
or ( n42426 , n42083 , n42425 );
and ( n42427 , n42080 , n42426 );
or ( n42428 , n42079 , n42427 );
and ( n42429 , n42076 , n42428 );
or ( n42430 , n42075 , n42429 );
and ( n42431 , n42072 , n42430 );
or ( n42432 , n42071 , n42431 );
and ( n42433 , n42068 , n42432 );
or ( n42434 , n42067 , n42433 );
and ( n42435 , n42064 , n42434 );
or ( n42436 , n42063 , n42435 );
and ( n42437 , n42060 , n42436 );
or ( n42438 , n42059 , n42437 );
and ( n42439 , n42056 , n42438 );
or ( n42440 , n42055 , n42439 );
and ( n42441 , n42052 , n42440 );
or ( n42442 , n42051 , n42441 );
and ( n42443 , n42048 , n42442 );
or ( n42444 , n42047 , n42443 );
and ( n42445 , n42044 , n42444 );
or ( n42446 , n42043 , n42445 );
and ( n42447 , n42040 , n42446 );
or ( n42448 , n42039 , n42447 );
and ( n42449 , n42036 , n42448 );
or ( n42450 , n42035 , n42449 );
and ( n42451 , n42032 , n42450 );
or ( n42452 , n42031 , n42451 );
and ( n42453 , n42028 , n42452 );
or ( n42454 , n42027 , n42453 );
and ( n42455 , n42024 , n42454 );
or ( n42456 , n42023 , n42455 );
and ( n42457 , n42020 , n42456 );
or ( n42458 , n42019 , n42457 );
and ( n42459 , n42016 , n42458 );
or ( n42460 , n42015 , n42459 );
and ( n42461 , n42012 , n42460 );
or ( n42462 , n42011 , n42461 );
and ( n42463 , n42008 , n42462 );
or ( n42464 , n42007 , n42463 );
and ( n42465 , n42004 , n42464 );
or ( n42466 , n42003 , n42465 );
and ( n42467 , n42000 , n42466 );
or ( n42468 , n41999 , n42467 );
and ( n42469 , n41996 , n42468 );
or ( n42470 , n41995 , n42469 );
and ( n42471 , n41992 , n42470 );
or ( n42472 , n41991 , n42471 );
and ( n42473 , n41988 , n42472 );
or ( n42474 , n41987 , n42473 );
and ( n42475 , n41984 , n42474 );
or ( n42476 , n41983 , n42475 );
and ( n42477 , n41980 , n42476 );
or ( n42478 , n41979 , n42477 );
and ( n42479 , n41976 , n42478 );
or ( n42480 , n41975 , n42479 );
and ( n42481 , n41972 , n42480 );
or ( n42482 , n41971 , n42481 );
and ( n42483 , n41968 , n42482 );
or ( n42484 , n41967 , n42483 );
and ( n42485 , n41964 , n42484 );
or ( n42486 , n41963 , n42485 );
and ( n42487 , n41960 , n42486 );
or ( n42488 , n41959 , n42487 );
and ( n42489 , n41956 , n42488 );
or ( n42490 , n41955 , n42489 );
and ( n42491 , n41952 , n42490 );
or ( n42492 , n41951 , n42491 );
and ( n42493 , n41948 , n42492 );
or ( n42494 , n41947 , n42493 );
and ( n42495 , n41944 , n42494 );
or ( n42496 , n41943 , n42495 );
and ( n42497 , n41940 , n42496 );
or ( n42498 , n41939 , n42497 );
and ( n42499 , n41936 , n42498 );
or ( n42500 , n41935 , n42499 );
and ( n42501 , n41932 , n42500 );
or ( n42502 , n41931 , n42501 );
and ( n42503 , n41928 , n42502 );
or ( n42504 , n41927 , n42503 );
and ( n42505 , n41924 , n42504 );
or ( n42506 , n41923 , n42505 );
and ( n42507 , n41920 , n42506 );
or ( n42508 , n41919 , n42507 );
and ( n42509 , n41916 , n42508 );
or ( n42510 , n41915 , n42509 );
and ( n42511 , n41912 , n42510 );
or ( n42512 , n41911 , n42511 );
and ( n42513 , n41908 , n42512 );
or ( n42514 , n41907 , n42513 );
and ( n42515 , n41904 , n42514 );
or ( n42516 , n41903 , n42515 );
and ( n42517 , n41900 , n42516 );
or ( n42518 , n41899 , n42517 );
and ( n42519 , n41896 , n42518 );
or ( n42520 , n41895 , n42519 );
and ( n42521 , n41892 , n42520 );
or ( n42522 , n41891 , n42521 );
and ( n42523 , n41888 , n42522 );
or ( n42524 , n41887 , n42523 );
and ( n42525 , n41884 , n42524 );
or ( n42526 , n41883 , n42525 );
xor ( n42527 , n41880 , n42526 );
buf ( n42528 , n18068 );
and ( n42529 , n29874 , n42528 );
xor ( n42530 , n42527 , n42529 );
xor ( n42531 , n41884 , n42524 );
and ( n42532 , n29879 , n42528 );
and ( n42533 , n42531 , n42532 );
xor ( n42534 , n42531 , n42532 );
xor ( n42535 , n41888 , n42522 );
and ( n42536 , n29884 , n42528 );
and ( n42537 , n42535 , n42536 );
xor ( n42538 , n42535 , n42536 );
xor ( n42539 , n41892 , n42520 );
and ( n42540 , n29889 , n42528 );
and ( n42541 , n42539 , n42540 );
xor ( n42542 , n42539 , n42540 );
xor ( n42543 , n41896 , n42518 );
and ( n42544 , n29894 , n42528 );
and ( n42545 , n42543 , n42544 );
xor ( n42546 , n42543 , n42544 );
xor ( n42547 , n41900 , n42516 );
and ( n42548 , n29899 , n42528 );
and ( n42549 , n42547 , n42548 );
xor ( n42550 , n42547 , n42548 );
xor ( n42551 , n41904 , n42514 );
and ( n42552 , n29904 , n42528 );
and ( n42553 , n42551 , n42552 );
xor ( n42554 , n42551 , n42552 );
xor ( n42555 , n41908 , n42512 );
and ( n42556 , n29909 , n42528 );
and ( n42557 , n42555 , n42556 );
xor ( n42558 , n42555 , n42556 );
xor ( n42559 , n41912 , n42510 );
and ( n42560 , n29914 , n42528 );
and ( n42561 , n42559 , n42560 );
xor ( n42562 , n42559 , n42560 );
xor ( n42563 , n41916 , n42508 );
and ( n42564 , n29919 , n42528 );
and ( n42565 , n42563 , n42564 );
xor ( n42566 , n42563 , n42564 );
xor ( n42567 , n41920 , n42506 );
and ( n42568 , n29924 , n42528 );
and ( n42569 , n42567 , n42568 );
xor ( n42570 , n42567 , n42568 );
xor ( n42571 , n41924 , n42504 );
and ( n42572 , n29929 , n42528 );
and ( n42573 , n42571 , n42572 );
xor ( n42574 , n42571 , n42572 );
xor ( n42575 , n41928 , n42502 );
and ( n42576 , n29934 , n42528 );
and ( n42577 , n42575 , n42576 );
xor ( n42578 , n42575 , n42576 );
xor ( n42579 , n41932 , n42500 );
and ( n42580 , n29939 , n42528 );
and ( n42581 , n42579 , n42580 );
xor ( n42582 , n42579 , n42580 );
xor ( n42583 , n41936 , n42498 );
and ( n42584 , n29944 , n42528 );
and ( n42585 , n42583 , n42584 );
xor ( n42586 , n42583 , n42584 );
xor ( n42587 , n41940 , n42496 );
and ( n42588 , n29949 , n42528 );
and ( n42589 , n42587 , n42588 );
xor ( n42590 , n42587 , n42588 );
xor ( n42591 , n41944 , n42494 );
and ( n42592 , n29954 , n42528 );
and ( n42593 , n42591 , n42592 );
xor ( n42594 , n42591 , n42592 );
xor ( n42595 , n41948 , n42492 );
and ( n42596 , n29959 , n42528 );
and ( n42597 , n42595 , n42596 );
xor ( n42598 , n42595 , n42596 );
xor ( n42599 , n41952 , n42490 );
and ( n42600 , n29964 , n42528 );
and ( n42601 , n42599 , n42600 );
xor ( n42602 , n42599 , n42600 );
xor ( n42603 , n41956 , n42488 );
and ( n42604 , n29969 , n42528 );
and ( n42605 , n42603 , n42604 );
xor ( n42606 , n42603 , n42604 );
xor ( n42607 , n41960 , n42486 );
and ( n42608 , n29974 , n42528 );
and ( n42609 , n42607 , n42608 );
xor ( n42610 , n42607 , n42608 );
xor ( n42611 , n41964 , n42484 );
and ( n42612 , n29979 , n42528 );
and ( n42613 , n42611 , n42612 );
xor ( n42614 , n42611 , n42612 );
xor ( n42615 , n41968 , n42482 );
and ( n42616 , n29984 , n42528 );
and ( n42617 , n42615 , n42616 );
xor ( n42618 , n42615 , n42616 );
xor ( n42619 , n41972 , n42480 );
and ( n42620 , n29989 , n42528 );
and ( n42621 , n42619 , n42620 );
xor ( n42622 , n42619 , n42620 );
xor ( n42623 , n41976 , n42478 );
and ( n42624 , n29994 , n42528 );
and ( n42625 , n42623 , n42624 );
xor ( n42626 , n42623 , n42624 );
xor ( n42627 , n41980 , n42476 );
and ( n42628 , n29999 , n42528 );
and ( n42629 , n42627 , n42628 );
xor ( n42630 , n42627 , n42628 );
xor ( n42631 , n41984 , n42474 );
and ( n42632 , n30004 , n42528 );
and ( n42633 , n42631 , n42632 );
xor ( n42634 , n42631 , n42632 );
xor ( n42635 , n41988 , n42472 );
and ( n42636 , n30009 , n42528 );
and ( n42637 , n42635 , n42636 );
xor ( n42638 , n42635 , n42636 );
xor ( n42639 , n41992 , n42470 );
and ( n42640 , n30014 , n42528 );
and ( n42641 , n42639 , n42640 );
xor ( n42642 , n42639 , n42640 );
xor ( n42643 , n41996 , n42468 );
and ( n42644 , n30019 , n42528 );
and ( n42645 , n42643 , n42644 );
xor ( n42646 , n42643 , n42644 );
xor ( n42647 , n42000 , n42466 );
and ( n42648 , n30024 , n42528 );
and ( n42649 , n42647 , n42648 );
xor ( n42650 , n42647 , n42648 );
xor ( n42651 , n42004 , n42464 );
and ( n42652 , n30029 , n42528 );
and ( n42653 , n42651 , n42652 );
xor ( n42654 , n42651 , n42652 );
xor ( n42655 , n42008 , n42462 );
and ( n42656 , n30034 , n42528 );
and ( n42657 , n42655 , n42656 );
xor ( n42658 , n42655 , n42656 );
xor ( n42659 , n42012 , n42460 );
and ( n42660 , n30039 , n42528 );
and ( n42661 , n42659 , n42660 );
xor ( n42662 , n42659 , n42660 );
xor ( n42663 , n42016 , n42458 );
and ( n42664 , n30044 , n42528 );
and ( n42665 , n42663 , n42664 );
xor ( n42666 , n42663 , n42664 );
xor ( n42667 , n42020 , n42456 );
and ( n42668 , n30049 , n42528 );
and ( n42669 , n42667 , n42668 );
xor ( n42670 , n42667 , n42668 );
xor ( n42671 , n42024 , n42454 );
and ( n42672 , n30054 , n42528 );
and ( n42673 , n42671 , n42672 );
xor ( n42674 , n42671 , n42672 );
xor ( n42675 , n42028 , n42452 );
and ( n42676 , n30059 , n42528 );
and ( n42677 , n42675 , n42676 );
xor ( n42678 , n42675 , n42676 );
xor ( n42679 , n42032 , n42450 );
and ( n42680 , n30064 , n42528 );
and ( n42681 , n42679 , n42680 );
xor ( n42682 , n42679 , n42680 );
xor ( n42683 , n42036 , n42448 );
and ( n42684 , n30069 , n42528 );
and ( n42685 , n42683 , n42684 );
xor ( n42686 , n42683 , n42684 );
xor ( n42687 , n42040 , n42446 );
and ( n42688 , n30074 , n42528 );
and ( n42689 , n42687 , n42688 );
xor ( n42690 , n42687 , n42688 );
xor ( n42691 , n42044 , n42444 );
and ( n42692 , n30079 , n42528 );
and ( n42693 , n42691 , n42692 );
xor ( n42694 , n42691 , n42692 );
xor ( n42695 , n42048 , n42442 );
and ( n42696 , n30084 , n42528 );
and ( n42697 , n42695 , n42696 );
xor ( n42698 , n42695 , n42696 );
xor ( n42699 , n42052 , n42440 );
and ( n42700 , n30089 , n42528 );
and ( n42701 , n42699 , n42700 );
xor ( n42702 , n42699 , n42700 );
xor ( n42703 , n42056 , n42438 );
and ( n42704 , n30094 , n42528 );
and ( n42705 , n42703 , n42704 );
xor ( n42706 , n42703 , n42704 );
xor ( n42707 , n42060 , n42436 );
and ( n42708 , n30099 , n42528 );
and ( n42709 , n42707 , n42708 );
xor ( n42710 , n42707 , n42708 );
xor ( n42711 , n42064 , n42434 );
and ( n42712 , n30104 , n42528 );
and ( n42713 , n42711 , n42712 );
xor ( n42714 , n42711 , n42712 );
xor ( n42715 , n42068 , n42432 );
and ( n42716 , n30109 , n42528 );
and ( n42717 , n42715 , n42716 );
xor ( n42718 , n42715 , n42716 );
xor ( n42719 , n42072 , n42430 );
and ( n42720 , n30114 , n42528 );
and ( n42721 , n42719 , n42720 );
xor ( n42722 , n42719 , n42720 );
xor ( n42723 , n42076 , n42428 );
and ( n42724 , n30119 , n42528 );
and ( n42725 , n42723 , n42724 );
xor ( n42726 , n42723 , n42724 );
xor ( n42727 , n42080 , n42426 );
and ( n42728 , n30124 , n42528 );
and ( n42729 , n42727 , n42728 );
xor ( n42730 , n42727 , n42728 );
xor ( n42731 , n42084 , n42424 );
and ( n42732 , n30129 , n42528 );
and ( n42733 , n42731 , n42732 );
xor ( n42734 , n42731 , n42732 );
xor ( n42735 , n42088 , n42422 );
and ( n42736 , n30134 , n42528 );
and ( n42737 , n42735 , n42736 );
xor ( n42738 , n42735 , n42736 );
xor ( n42739 , n42092 , n42420 );
and ( n42740 , n30139 , n42528 );
and ( n42741 , n42739 , n42740 );
xor ( n42742 , n42739 , n42740 );
xor ( n42743 , n42096 , n42418 );
and ( n42744 , n30144 , n42528 );
and ( n42745 , n42743 , n42744 );
xor ( n42746 , n42743 , n42744 );
xor ( n42747 , n42100 , n42416 );
and ( n42748 , n30149 , n42528 );
and ( n42749 , n42747 , n42748 );
xor ( n42750 , n42747 , n42748 );
xor ( n42751 , n42104 , n42414 );
and ( n42752 , n30154 , n42528 );
and ( n42753 , n42751 , n42752 );
xor ( n42754 , n42751 , n42752 );
xor ( n42755 , n42108 , n42412 );
and ( n42756 , n30159 , n42528 );
and ( n42757 , n42755 , n42756 );
xor ( n42758 , n42755 , n42756 );
xor ( n42759 , n42112 , n42410 );
and ( n42760 , n30164 , n42528 );
and ( n42761 , n42759 , n42760 );
xor ( n42762 , n42759 , n42760 );
xor ( n42763 , n42116 , n42408 );
and ( n42764 , n30169 , n42528 );
and ( n42765 , n42763 , n42764 );
xor ( n42766 , n42763 , n42764 );
xor ( n42767 , n42120 , n42406 );
and ( n42768 , n30174 , n42528 );
and ( n42769 , n42767 , n42768 );
xor ( n42770 , n42767 , n42768 );
xor ( n42771 , n42124 , n42404 );
and ( n42772 , n30179 , n42528 );
and ( n42773 , n42771 , n42772 );
xor ( n42774 , n42771 , n42772 );
xor ( n42775 , n42128 , n42402 );
and ( n42776 , n30184 , n42528 );
and ( n42777 , n42775 , n42776 );
xor ( n42778 , n42775 , n42776 );
xor ( n42779 , n42132 , n42400 );
and ( n42780 , n30189 , n42528 );
and ( n42781 , n42779 , n42780 );
xor ( n42782 , n42779 , n42780 );
xor ( n42783 , n42136 , n42398 );
and ( n42784 , n30194 , n42528 );
and ( n42785 , n42783 , n42784 );
xor ( n42786 , n42783 , n42784 );
xor ( n42787 , n42140 , n42396 );
and ( n42788 , n30199 , n42528 );
and ( n42789 , n42787 , n42788 );
xor ( n42790 , n42787 , n42788 );
xor ( n42791 , n42144 , n42394 );
and ( n42792 , n30204 , n42528 );
and ( n42793 , n42791 , n42792 );
xor ( n42794 , n42791 , n42792 );
xor ( n42795 , n42148 , n42392 );
and ( n42796 , n30209 , n42528 );
and ( n42797 , n42795 , n42796 );
xor ( n42798 , n42795 , n42796 );
xor ( n42799 , n42152 , n42390 );
and ( n42800 , n30214 , n42528 );
and ( n42801 , n42799 , n42800 );
xor ( n42802 , n42799 , n42800 );
xor ( n42803 , n42156 , n42388 );
and ( n42804 , n30219 , n42528 );
and ( n42805 , n42803 , n42804 );
xor ( n42806 , n42803 , n42804 );
xor ( n42807 , n42160 , n42386 );
and ( n42808 , n30224 , n42528 );
and ( n42809 , n42807 , n42808 );
xor ( n42810 , n42807 , n42808 );
xor ( n42811 , n42164 , n42384 );
and ( n42812 , n30229 , n42528 );
and ( n42813 , n42811 , n42812 );
xor ( n42814 , n42811 , n42812 );
xor ( n42815 , n42168 , n42382 );
and ( n42816 , n30234 , n42528 );
and ( n42817 , n42815 , n42816 );
xor ( n42818 , n42815 , n42816 );
xor ( n42819 , n42172 , n42380 );
and ( n42820 , n30239 , n42528 );
and ( n42821 , n42819 , n42820 );
xor ( n42822 , n42819 , n42820 );
xor ( n42823 , n42176 , n42378 );
and ( n42824 , n30244 , n42528 );
and ( n42825 , n42823 , n42824 );
xor ( n42826 , n42823 , n42824 );
xor ( n42827 , n42180 , n42376 );
and ( n42828 , n30249 , n42528 );
and ( n42829 , n42827 , n42828 );
xor ( n42830 , n42827 , n42828 );
xor ( n42831 , n42184 , n42374 );
and ( n42832 , n30254 , n42528 );
and ( n42833 , n42831 , n42832 );
xor ( n42834 , n42831 , n42832 );
xor ( n42835 , n42188 , n42372 );
and ( n42836 , n30259 , n42528 );
and ( n42837 , n42835 , n42836 );
xor ( n42838 , n42835 , n42836 );
xor ( n42839 , n42192 , n42370 );
and ( n42840 , n30264 , n42528 );
and ( n42841 , n42839 , n42840 );
xor ( n42842 , n42839 , n42840 );
xor ( n42843 , n42196 , n42368 );
and ( n42844 , n30269 , n42528 );
and ( n42845 , n42843 , n42844 );
xor ( n42846 , n42843 , n42844 );
xor ( n42847 , n42200 , n42366 );
and ( n42848 , n30274 , n42528 );
and ( n42849 , n42847 , n42848 );
xor ( n42850 , n42847 , n42848 );
xor ( n42851 , n42204 , n42364 );
and ( n42852 , n30279 , n42528 );
and ( n42853 , n42851 , n42852 );
xor ( n42854 , n42851 , n42852 );
xor ( n42855 , n42208 , n42362 );
and ( n42856 , n30284 , n42528 );
and ( n42857 , n42855 , n42856 );
xor ( n42858 , n42855 , n42856 );
xor ( n42859 , n42212 , n42360 );
and ( n42860 , n30289 , n42528 );
and ( n42861 , n42859 , n42860 );
xor ( n42862 , n42859 , n42860 );
xor ( n42863 , n42216 , n42358 );
and ( n42864 , n30294 , n42528 );
and ( n42865 , n42863 , n42864 );
xor ( n42866 , n42863 , n42864 );
xor ( n42867 , n42220 , n42356 );
and ( n42868 , n30299 , n42528 );
and ( n42869 , n42867 , n42868 );
xor ( n42870 , n42867 , n42868 );
xor ( n42871 , n42224 , n42354 );
and ( n42872 , n30304 , n42528 );
and ( n42873 , n42871 , n42872 );
xor ( n42874 , n42871 , n42872 );
xor ( n42875 , n42228 , n42352 );
and ( n42876 , n30309 , n42528 );
and ( n42877 , n42875 , n42876 );
xor ( n42878 , n42875 , n42876 );
xor ( n42879 , n42232 , n42350 );
and ( n42880 , n30314 , n42528 );
and ( n42881 , n42879 , n42880 );
xor ( n42882 , n42879 , n42880 );
xor ( n42883 , n42236 , n42348 );
and ( n42884 , n30319 , n42528 );
and ( n42885 , n42883 , n42884 );
xor ( n42886 , n42883 , n42884 );
xor ( n42887 , n42240 , n42346 );
and ( n42888 , n30324 , n42528 );
and ( n42889 , n42887 , n42888 );
xor ( n42890 , n42887 , n42888 );
xor ( n42891 , n42244 , n42344 );
and ( n42892 , n30329 , n42528 );
and ( n42893 , n42891 , n42892 );
xor ( n42894 , n42891 , n42892 );
xor ( n42895 , n42248 , n42342 );
and ( n42896 , n30334 , n42528 );
and ( n42897 , n42895 , n42896 );
xor ( n42898 , n42895 , n42896 );
xor ( n42899 , n42252 , n42340 );
and ( n42900 , n30339 , n42528 );
and ( n42901 , n42899 , n42900 );
xor ( n42902 , n42899 , n42900 );
xor ( n42903 , n42256 , n42338 );
and ( n42904 , n30344 , n42528 );
and ( n42905 , n42903 , n42904 );
xor ( n42906 , n42903 , n42904 );
xor ( n42907 , n42260 , n42336 );
and ( n42908 , n30349 , n42528 );
and ( n42909 , n42907 , n42908 );
xor ( n42910 , n42907 , n42908 );
xor ( n42911 , n42264 , n42334 );
and ( n42912 , n30354 , n42528 );
and ( n42913 , n42911 , n42912 );
xor ( n42914 , n42911 , n42912 );
xor ( n42915 , n42268 , n42332 );
and ( n42916 , n30359 , n42528 );
and ( n42917 , n42915 , n42916 );
xor ( n42918 , n42915 , n42916 );
xor ( n42919 , n42272 , n42330 );
and ( n42920 , n30364 , n42528 );
and ( n42921 , n42919 , n42920 );
xor ( n42922 , n42919 , n42920 );
xor ( n42923 , n42276 , n42328 );
and ( n42924 , n30369 , n42528 );
and ( n42925 , n42923 , n42924 );
xor ( n42926 , n42923 , n42924 );
xor ( n42927 , n42280 , n42326 );
and ( n42928 , n30374 , n42528 );
and ( n42929 , n42927 , n42928 );
xor ( n42930 , n42927 , n42928 );
xor ( n42931 , n42284 , n42324 );
and ( n42932 , n30379 , n42528 );
and ( n42933 , n42931 , n42932 );
xor ( n42934 , n42931 , n42932 );
xor ( n42935 , n42288 , n42322 );
and ( n42936 , n30384 , n42528 );
and ( n42937 , n42935 , n42936 );
xor ( n42938 , n42935 , n42936 );
xor ( n42939 , n42292 , n42320 );
and ( n42940 , n30389 , n42528 );
and ( n42941 , n42939 , n42940 );
xor ( n42942 , n42939 , n42940 );
xor ( n42943 , n42296 , n42318 );
and ( n42944 , n30394 , n42528 );
and ( n42945 , n42943 , n42944 );
xor ( n42946 , n42943 , n42944 );
xor ( n42947 , n42300 , n42316 );
and ( n42948 , n30399 , n42528 );
and ( n42949 , n42947 , n42948 );
xor ( n42950 , n42947 , n42948 );
xor ( n42951 , n42304 , n42314 );
and ( n42952 , n30404 , n42528 );
and ( n42953 , n42951 , n42952 );
xor ( n42954 , n42951 , n42952 );
xor ( n42955 , n42308 , n42312 );
and ( n42956 , n30409 , n42528 );
and ( n42957 , n42955 , n42956 );
buf ( n42958 , n42957 );
and ( n42959 , n42954 , n42958 );
or ( n42960 , n42953 , n42959 );
and ( n42961 , n42950 , n42960 );
or ( n42962 , n42949 , n42961 );
and ( n42963 , n42946 , n42962 );
or ( n42964 , n42945 , n42963 );
and ( n42965 , n42942 , n42964 );
or ( n42966 , n42941 , n42965 );
and ( n42967 , n42938 , n42966 );
or ( n42968 , n42937 , n42967 );
and ( n42969 , n42934 , n42968 );
or ( n42970 , n42933 , n42969 );
and ( n42971 , n42930 , n42970 );
or ( n42972 , n42929 , n42971 );
and ( n42973 , n42926 , n42972 );
or ( n42974 , n42925 , n42973 );
and ( n42975 , n42922 , n42974 );
or ( n42976 , n42921 , n42975 );
and ( n42977 , n42918 , n42976 );
or ( n42978 , n42917 , n42977 );
and ( n42979 , n42914 , n42978 );
or ( n42980 , n42913 , n42979 );
and ( n42981 , n42910 , n42980 );
or ( n42982 , n42909 , n42981 );
and ( n42983 , n42906 , n42982 );
or ( n42984 , n42905 , n42983 );
and ( n42985 , n42902 , n42984 );
or ( n42986 , n42901 , n42985 );
and ( n42987 , n42898 , n42986 );
or ( n42988 , n42897 , n42987 );
and ( n42989 , n42894 , n42988 );
or ( n42990 , n42893 , n42989 );
and ( n42991 , n42890 , n42990 );
or ( n42992 , n42889 , n42991 );
and ( n42993 , n42886 , n42992 );
or ( n42994 , n42885 , n42993 );
and ( n42995 , n42882 , n42994 );
or ( n42996 , n42881 , n42995 );
and ( n42997 , n42878 , n42996 );
or ( n42998 , n42877 , n42997 );
and ( n42999 , n42874 , n42998 );
or ( n43000 , n42873 , n42999 );
and ( n43001 , n42870 , n43000 );
or ( n43002 , n42869 , n43001 );
and ( n43003 , n42866 , n43002 );
or ( n43004 , n42865 , n43003 );
and ( n43005 , n42862 , n43004 );
or ( n43006 , n42861 , n43005 );
and ( n43007 , n42858 , n43006 );
or ( n43008 , n42857 , n43007 );
and ( n43009 , n42854 , n43008 );
or ( n43010 , n42853 , n43009 );
and ( n43011 , n42850 , n43010 );
or ( n43012 , n42849 , n43011 );
and ( n43013 , n42846 , n43012 );
or ( n43014 , n42845 , n43013 );
and ( n43015 , n42842 , n43014 );
or ( n43016 , n42841 , n43015 );
and ( n43017 , n42838 , n43016 );
or ( n43018 , n42837 , n43017 );
and ( n43019 , n42834 , n43018 );
or ( n43020 , n42833 , n43019 );
and ( n43021 , n42830 , n43020 );
or ( n43022 , n42829 , n43021 );
and ( n43023 , n42826 , n43022 );
or ( n43024 , n42825 , n43023 );
and ( n43025 , n42822 , n43024 );
or ( n43026 , n42821 , n43025 );
and ( n43027 , n42818 , n43026 );
or ( n43028 , n42817 , n43027 );
and ( n43029 , n42814 , n43028 );
or ( n43030 , n42813 , n43029 );
and ( n43031 , n42810 , n43030 );
or ( n43032 , n42809 , n43031 );
and ( n43033 , n42806 , n43032 );
or ( n43034 , n42805 , n43033 );
and ( n43035 , n42802 , n43034 );
or ( n43036 , n42801 , n43035 );
and ( n43037 , n42798 , n43036 );
or ( n43038 , n42797 , n43037 );
and ( n43039 , n42794 , n43038 );
or ( n43040 , n42793 , n43039 );
and ( n43041 , n42790 , n43040 );
or ( n43042 , n42789 , n43041 );
and ( n43043 , n42786 , n43042 );
or ( n43044 , n42785 , n43043 );
and ( n43045 , n42782 , n43044 );
or ( n43046 , n42781 , n43045 );
and ( n43047 , n42778 , n43046 );
or ( n43048 , n42777 , n43047 );
and ( n43049 , n42774 , n43048 );
or ( n43050 , n42773 , n43049 );
and ( n43051 , n42770 , n43050 );
or ( n43052 , n42769 , n43051 );
and ( n43053 , n42766 , n43052 );
or ( n43054 , n42765 , n43053 );
and ( n43055 , n42762 , n43054 );
or ( n43056 , n42761 , n43055 );
and ( n43057 , n42758 , n43056 );
or ( n43058 , n42757 , n43057 );
and ( n43059 , n42754 , n43058 );
or ( n43060 , n42753 , n43059 );
and ( n43061 , n42750 , n43060 );
or ( n43062 , n42749 , n43061 );
and ( n43063 , n42746 , n43062 );
or ( n43064 , n42745 , n43063 );
and ( n43065 , n42742 , n43064 );
or ( n43066 , n42741 , n43065 );
and ( n43067 , n42738 , n43066 );
or ( n43068 , n42737 , n43067 );
and ( n43069 , n42734 , n43068 );
or ( n43070 , n42733 , n43069 );
and ( n43071 , n42730 , n43070 );
or ( n43072 , n42729 , n43071 );
and ( n43073 , n42726 , n43072 );
or ( n43074 , n42725 , n43073 );
and ( n43075 , n42722 , n43074 );
or ( n43076 , n42721 , n43075 );
and ( n43077 , n42718 , n43076 );
or ( n43078 , n42717 , n43077 );
and ( n43079 , n42714 , n43078 );
or ( n43080 , n42713 , n43079 );
and ( n43081 , n42710 , n43080 );
or ( n43082 , n42709 , n43081 );
and ( n43083 , n42706 , n43082 );
or ( n43084 , n42705 , n43083 );
and ( n43085 , n42702 , n43084 );
or ( n43086 , n42701 , n43085 );
and ( n43087 , n42698 , n43086 );
or ( n43088 , n42697 , n43087 );
and ( n43089 , n42694 , n43088 );
or ( n43090 , n42693 , n43089 );
and ( n43091 , n42690 , n43090 );
or ( n43092 , n42689 , n43091 );
and ( n43093 , n42686 , n43092 );
or ( n43094 , n42685 , n43093 );
and ( n43095 , n42682 , n43094 );
or ( n43096 , n42681 , n43095 );
and ( n43097 , n42678 , n43096 );
or ( n43098 , n42677 , n43097 );
and ( n43099 , n42674 , n43098 );
or ( n43100 , n42673 , n43099 );
and ( n43101 , n42670 , n43100 );
or ( n43102 , n42669 , n43101 );
and ( n43103 , n42666 , n43102 );
or ( n43104 , n42665 , n43103 );
and ( n43105 , n42662 , n43104 );
or ( n43106 , n42661 , n43105 );
and ( n43107 , n42658 , n43106 );
or ( n43108 , n42657 , n43107 );
and ( n43109 , n42654 , n43108 );
or ( n43110 , n42653 , n43109 );
and ( n43111 , n42650 , n43110 );
or ( n43112 , n42649 , n43111 );
and ( n43113 , n42646 , n43112 );
or ( n43114 , n42645 , n43113 );
and ( n43115 , n42642 , n43114 );
or ( n43116 , n42641 , n43115 );
and ( n43117 , n42638 , n43116 );
or ( n43118 , n42637 , n43117 );
and ( n43119 , n42634 , n43118 );
or ( n43120 , n42633 , n43119 );
and ( n43121 , n42630 , n43120 );
or ( n43122 , n42629 , n43121 );
and ( n43123 , n42626 , n43122 );
or ( n43124 , n42625 , n43123 );
and ( n43125 , n42622 , n43124 );
or ( n43126 , n42621 , n43125 );
and ( n43127 , n42618 , n43126 );
or ( n43128 , n42617 , n43127 );
and ( n43129 , n42614 , n43128 );
or ( n43130 , n42613 , n43129 );
and ( n43131 , n42610 , n43130 );
or ( n43132 , n42609 , n43131 );
and ( n43133 , n42606 , n43132 );
or ( n43134 , n42605 , n43133 );
and ( n43135 , n42602 , n43134 );
or ( n43136 , n42601 , n43135 );
and ( n43137 , n42598 , n43136 );
or ( n43138 , n42597 , n43137 );
and ( n43139 , n42594 , n43138 );
or ( n43140 , n42593 , n43139 );
and ( n43141 , n42590 , n43140 );
or ( n43142 , n42589 , n43141 );
and ( n43143 , n42586 , n43142 );
or ( n43144 , n42585 , n43143 );
and ( n43145 , n42582 , n43144 );
or ( n43146 , n42581 , n43145 );
and ( n43147 , n42578 , n43146 );
or ( n43148 , n42577 , n43147 );
and ( n43149 , n42574 , n43148 );
or ( n43150 , n42573 , n43149 );
and ( n43151 , n42570 , n43150 );
or ( n43152 , n42569 , n43151 );
and ( n43153 , n42566 , n43152 );
or ( n43154 , n42565 , n43153 );
and ( n43155 , n42562 , n43154 );
or ( n43156 , n42561 , n43155 );
and ( n43157 , n42558 , n43156 );
or ( n43158 , n42557 , n43157 );
and ( n43159 , n42554 , n43158 );
or ( n43160 , n42553 , n43159 );
and ( n43161 , n42550 , n43160 );
or ( n43162 , n42549 , n43161 );
and ( n43163 , n42546 , n43162 );
or ( n43164 , n42545 , n43163 );
and ( n43165 , n42542 , n43164 );
or ( n43166 , n42541 , n43165 );
and ( n43167 , n42538 , n43166 );
or ( n43168 , n42537 , n43167 );
and ( n43169 , n42534 , n43168 );
or ( n43170 , n42533 , n43169 );
xor ( n43171 , n42530 , n43170 );
buf ( n43172 , n18066 );
and ( n43173 , n29879 , n43172 );
xor ( n43174 , n43171 , n43173 );
xor ( n43175 , n42534 , n43168 );
and ( n43176 , n29884 , n43172 );
and ( n43177 , n43175 , n43176 );
xor ( n43178 , n43175 , n43176 );
xor ( n43179 , n42538 , n43166 );
and ( n43180 , n29889 , n43172 );
and ( n43181 , n43179 , n43180 );
xor ( n43182 , n43179 , n43180 );
xor ( n43183 , n42542 , n43164 );
and ( n43184 , n29894 , n43172 );
and ( n43185 , n43183 , n43184 );
xor ( n43186 , n43183 , n43184 );
xor ( n43187 , n42546 , n43162 );
and ( n43188 , n29899 , n43172 );
and ( n43189 , n43187 , n43188 );
xor ( n43190 , n43187 , n43188 );
xor ( n43191 , n42550 , n43160 );
and ( n43192 , n29904 , n43172 );
and ( n43193 , n43191 , n43192 );
xor ( n43194 , n43191 , n43192 );
xor ( n43195 , n42554 , n43158 );
and ( n43196 , n29909 , n43172 );
and ( n43197 , n43195 , n43196 );
xor ( n43198 , n43195 , n43196 );
xor ( n43199 , n42558 , n43156 );
and ( n43200 , n29914 , n43172 );
and ( n43201 , n43199 , n43200 );
xor ( n43202 , n43199 , n43200 );
xor ( n43203 , n42562 , n43154 );
and ( n43204 , n29919 , n43172 );
and ( n43205 , n43203 , n43204 );
xor ( n43206 , n43203 , n43204 );
xor ( n43207 , n42566 , n43152 );
and ( n43208 , n29924 , n43172 );
and ( n43209 , n43207 , n43208 );
xor ( n43210 , n43207 , n43208 );
xor ( n43211 , n42570 , n43150 );
and ( n43212 , n29929 , n43172 );
and ( n43213 , n43211 , n43212 );
xor ( n43214 , n43211 , n43212 );
xor ( n43215 , n42574 , n43148 );
and ( n43216 , n29934 , n43172 );
and ( n43217 , n43215 , n43216 );
xor ( n43218 , n43215 , n43216 );
xor ( n43219 , n42578 , n43146 );
and ( n43220 , n29939 , n43172 );
and ( n43221 , n43219 , n43220 );
xor ( n43222 , n43219 , n43220 );
xor ( n43223 , n42582 , n43144 );
and ( n43224 , n29944 , n43172 );
and ( n43225 , n43223 , n43224 );
xor ( n43226 , n43223 , n43224 );
xor ( n43227 , n42586 , n43142 );
and ( n43228 , n29949 , n43172 );
and ( n43229 , n43227 , n43228 );
xor ( n43230 , n43227 , n43228 );
xor ( n43231 , n42590 , n43140 );
and ( n43232 , n29954 , n43172 );
and ( n43233 , n43231 , n43232 );
xor ( n43234 , n43231 , n43232 );
xor ( n43235 , n42594 , n43138 );
and ( n43236 , n29959 , n43172 );
and ( n43237 , n43235 , n43236 );
xor ( n43238 , n43235 , n43236 );
xor ( n43239 , n42598 , n43136 );
and ( n43240 , n29964 , n43172 );
and ( n43241 , n43239 , n43240 );
xor ( n43242 , n43239 , n43240 );
xor ( n43243 , n42602 , n43134 );
and ( n43244 , n29969 , n43172 );
and ( n43245 , n43243 , n43244 );
xor ( n43246 , n43243 , n43244 );
xor ( n43247 , n42606 , n43132 );
and ( n43248 , n29974 , n43172 );
and ( n43249 , n43247 , n43248 );
xor ( n43250 , n43247 , n43248 );
xor ( n43251 , n42610 , n43130 );
and ( n43252 , n29979 , n43172 );
and ( n43253 , n43251 , n43252 );
xor ( n43254 , n43251 , n43252 );
xor ( n43255 , n42614 , n43128 );
and ( n43256 , n29984 , n43172 );
and ( n43257 , n43255 , n43256 );
xor ( n43258 , n43255 , n43256 );
xor ( n43259 , n42618 , n43126 );
and ( n43260 , n29989 , n43172 );
and ( n43261 , n43259 , n43260 );
xor ( n43262 , n43259 , n43260 );
xor ( n43263 , n42622 , n43124 );
and ( n43264 , n29994 , n43172 );
and ( n43265 , n43263 , n43264 );
xor ( n43266 , n43263 , n43264 );
xor ( n43267 , n42626 , n43122 );
and ( n43268 , n29999 , n43172 );
and ( n43269 , n43267 , n43268 );
xor ( n43270 , n43267 , n43268 );
xor ( n43271 , n42630 , n43120 );
and ( n43272 , n30004 , n43172 );
and ( n43273 , n43271 , n43272 );
xor ( n43274 , n43271 , n43272 );
xor ( n43275 , n42634 , n43118 );
and ( n43276 , n30009 , n43172 );
and ( n43277 , n43275 , n43276 );
xor ( n43278 , n43275 , n43276 );
xor ( n43279 , n42638 , n43116 );
and ( n43280 , n30014 , n43172 );
and ( n43281 , n43279 , n43280 );
xor ( n43282 , n43279 , n43280 );
xor ( n43283 , n42642 , n43114 );
and ( n43284 , n30019 , n43172 );
and ( n43285 , n43283 , n43284 );
xor ( n43286 , n43283 , n43284 );
xor ( n43287 , n42646 , n43112 );
and ( n43288 , n30024 , n43172 );
and ( n43289 , n43287 , n43288 );
xor ( n43290 , n43287 , n43288 );
xor ( n43291 , n42650 , n43110 );
and ( n43292 , n30029 , n43172 );
and ( n43293 , n43291 , n43292 );
xor ( n43294 , n43291 , n43292 );
xor ( n43295 , n42654 , n43108 );
and ( n43296 , n30034 , n43172 );
and ( n43297 , n43295 , n43296 );
xor ( n43298 , n43295 , n43296 );
xor ( n43299 , n42658 , n43106 );
and ( n43300 , n30039 , n43172 );
and ( n43301 , n43299 , n43300 );
xor ( n43302 , n43299 , n43300 );
xor ( n43303 , n42662 , n43104 );
and ( n43304 , n30044 , n43172 );
and ( n43305 , n43303 , n43304 );
xor ( n43306 , n43303 , n43304 );
xor ( n43307 , n42666 , n43102 );
and ( n43308 , n30049 , n43172 );
and ( n43309 , n43307 , n43308 );
xor ( n43310 , n43307 , n43308 );
xor ( n43311 , n42670 , n43100 );
and ( n43312 , n30054 , n43172 );
and ( n43313 , n43311 , n43312 );
xor ( n43314 , n43311 , n43312 );
xor ( n43315 , n42674 , n43098 );
and ( n43316 , n30059 , n43172 );
and ( n43317 , n43315 , n43316 );
xor ( n43318 , n43315 , n43316 );
xor ( n43319 , n42678 , n43096 );
and ( n43320 , n30064 , n43172 );
and ( n43321 , n43319 , n43320 );
xor ( n43322 , n43319 , n43320 );
xor ( n43323 , n42682 , n43094 );
and ( n43324 , n30069 , n43172 );
and ( n43325 , n43323 , n43324 );
xor ( n43326 , n43323 , n43324 );
xor ( n43327 , n42686 , n43092 );
and ( n43328 , n30074 , n43172 );
and ( n43329 , n43327 , n43328 );
xor ( n43330 , n43327 , n43328 );
xor ( n43331 , n42690 , n43090 );
and ( n43332 , n30079 , n43172 );
and ( n43333 , n43331 , n43332 );
xor ( n43334 , n43331 , n43332 );
xor ( n43335 , n42694 , n43088 );
and ( n43336 , n30084 , n43172 );
and ( n43337 , n43335 , n43336 );
xor ( n43338 , n43335 , n43336 );
xor ( n43339 , n42698 , n43086 );
and ( n43340 , n30089 , n43172 );
and ( n43341 , n43339 , n43340 );
xor ( n43342 , n43339 , n43340 );
xor ( n43343 , n42702 , n43084 );
and ( n43344 , n30094 , n43172 );
and ( n43345 , n43343 , n43344 );
xor ( n43346 , n43343 , n43344 );
xor ( n43347 , n42706 , n43082 );
and ( n43348 , n30099 , n43172 );
and ( n43349 , n43347 , n43348 );
xor ( n43350 , n43347 , n43348 );
xor ( n43351 , n42710 , n43080 );
and ( n43352 , n30104 , n43172 );
and ( n43353 , n43351 , n43352 );
xor ( n43354 , n43351 , n43352 );
xor ( n43355 , n42714 , n43078 );
and ( n43356 , n30109 , n43172 );
and ( n43357 , n43355 , n43356 );
xor ( n43358 , n43355 , n43356 );
xor ( n43359 , n42718 , n43076 );
and ( n43360 , n30114 , n43172 );
and ( n43361 , n43359 , n43360 );
xor ( n43362 , n43359 , n43360 );
xor ( n43363 , n42722 , n43074 );
and ( n43364 , n30119 , n43172 );
and ( n43365 , n43363 , n43364 );
xor ( n43366 , n43363 , n43364 );
xor ( n43367 , n42726 , n43072 );
and ( n43368 , n30124 , n43172 );
and ( n43369 , n43367 , n43368 );
xor ( n43370 , n43367 , n43368 );
xor ( n43371 , n42730 , n43070 );
and ( n43372 , n30129 , n43172 );
and ( n43373 , n43371 , n43372 );
xor ( n43374 , n43371 , n43372 );
xor ( n43375 , n42734 , n43068 );
and ( n43376 , n30134 , n43172 );
and ( n43377 , n43375 , n43376 );
xor ( n43378 , n43375 , n43376 );
xor ( n43379 , n42738 , n43066 );
and ( n43380 , n30139 , n43172 );
and ( n43381 , n43379 , n43380 );
xor ( n43382 , n43379 , n43380 );
xor ( n43383 , n42742 , n43064 );
and ( n43384 , n30144 , n43172 );
and ( n43385 , n43383 , n43384 );
xor ( n43386 , n43383 , n43384 );
xor ( n43387 , n42746 , n43062 );
and ( n43388 , n30149 , n43172 );
and ( n43389 , n43387 , n43388 );
xor ( n43390 , n43387 , n43388 );
xor ( n43391 , n42750 , n43060 );
and ( n43392 , n30154 , n43172 );
and ( n43393 , n43391 , n43392 );
xor ( n43394 , n43391 , n43392 );
xor ( n43395 , n42754 , n43058 );
and ( n43396 , n30159 , n43172 );
and ( n43397 , n43395 , n43396 );
xor ( n43398 , n43395 , n43396 );
xor ( n43399 , n42758 , n43056 );
and ( n43400 , n30164 , n43172 );
and ( n43401 , n43399 , n43400 );
xor ( n43402 , n43399 , n43400 );
xor ( n43403 , n42762 , n43054 );
and ( n43404 , n30169 , n43172 );
and ( n43405 , n43403 , n43404 );
xor ( n43406 , n43403 , n43404 );
xor ( n43407 , n42766 , n43052 );
and ( n43408 , n30174 , n43172 );
and ( n43409 , n43407 , n43408 );
xor ( n43410 , n43407 , n43408 );
xor ( n43411 , n42770 , n43050 );
and ( n43412 , n30179 , n43172 );
and ( n43413 , n43411 , n43412 );
xor ( n43414 , n43411 , n43412 );
xor ( n43415 , n42774 , n43048 );
and ( n43416 , n30184 , n43172 );
and ( n43417 , n43415 , n43416 );
xor ( n43418 , n43415 , n43416 );
xor ( n43419 , n42778 , n43046 );
and ( n43420 , n30189 , n43172 );
and ( n43421 , n43419 , n43420 );
xor ( n43422 , n43419 , n43420 );
xor ( n43423 , n42782 , n43044 );
and ( n43424 , n30194 , n43172 );
and ( n43425 , n43423 , n43424 );
xor ( n43426 , n43423 , n43424 );
xor ( n43427 , n42786 , n43042 );
and ( n43428 , n30199 , n43172 );
and ( n43429 , n43427 , n43428 );
xor ( n43430 , n43427 , n43428 );
xor ( n43431 , n42790 , n43040 );
and ( n43432 , n30204 , n43172 );
and ( n43433 , n43431 , n43432 );
xor ( n43434 , n43431 , n43432 );
xor ( n43435 , n42794 , n43038 );
and ( n43436 , n30209 , n43172 );
and ( n43437 , n43435 , n43436 );
xor ( n43438 , n43435 , n43436 );
xor ( n43439 , n42798 , n43036 );
and ( n43440 , n30214 , n43172 );
and ( n43441 , n43439 , n43440 );
xor ( n43442 , n43439 , n43440 );
xor ( n43443 , n42802 , n43034 );
and ( n43444 , n30219 , n43172 );
and ( n43445 , n43443 , n43444 );
xor ( n43446 , n43443 , n43444 );
xor ( n43447 , n42806 , n43032 );
and ( n43448 , n30224 , n43172 );
and ( n43449 , n43447 , n43448 );
xor ( n43450 , n43447 , n43448 );
xor ( n43451 , n42810 , n43030 );
and ( n43452 , n30229 , n43172 );
and ( n43453 , n43451 , n43452 );
xor ( n43454 , n43451 , n43452 );
xor ( n43455 , n42814 , n43028 );
and ( n43456 , n30234 , n43172 );
and ( n43457 , n43455 , n43456 );
xor ( n43458 , n43455 , n43456 );
xor ( n43459 , n42818 , n43026 );
and ( n43460 , n30239 , n43172 );
and ( n43461 , n43459 , n43460 );
xor ( n43462 , n43459 , n43460 );
xor ( n43463 , n42822 , n43024 );
and ( n43464 , n30244 , n43172 );
and ( n43465 , n43463 , n43464 );
xor ( n43466 , n43463 , n43464 );
xor ( n43467 , n42826 , n43022 );
and ( n43468 , n30249 , n43172 );
and ( n43469 , n43467 , n43468 );
xor ( n43470 , n43467 , n43468 );
xor ( n43471 , n42830 , n43020 );
and ( n43472 , n30254 , n43172 );
and ( n43473 , n43471 , n43472 );
xor ( n43474 , n43471 , n43472 );
xor ( n43475 , n42834 , n43018 );
and ( n43476 , n30259 , n43172 );
and ( n43477 , n43475 , n43476 );
xor ( n43478 , n43475 , n43476 );
xor ( n43479 , n42838 , n43016 );
and ( n43480 , n30264 , n43172 );
and ( n43481 , n43479 , n43480 );
xor ( n43482 , n43479 , n43480 );
xor ( n43483 , n42842 , n43014 );
and ( n43484 , n30269 , n43172 );
and ( n43485 , n43483 , n43484 );
xor ( n43486 , n43483 , n43484 );
xor ( n43487 , n42846 , n43012 );
and ( n43488 , n30274 , n43172 );
and ( n43489 , n43487 , n43488 );
xor ( n43490 , n43487 , n43488 );
xor ( n43491 , n42850 , n43010 );
and ( n43492 , n30279 , n43172 );
and ( n43493 , n43491 , n43492 );
xor ( n43494 , n43491 , n43492 );
xor ( n43495 , n42854 , n43008 );
and ( n43496 , n30284 , n43172 );
and ( n43497 , n43495 , n43496 );
xor ( n43498 , n43495 , n43496 );
xor ( n43499 , n42858 , n43006 );
and ( n43500 , n30289 , n43172 );
and ( n43501 , n43499 , n43500 );
xor ( n43502 , n43499 , n43500 );
xor ( n43503 , n42862 , n43004 );
and ( n43504 , n30294 , n43172 );
and ( n43505 , n43503 , n43504 );
xor ( n43506 , n43503 , n43504 );
xor ( n43507 , n42866 , n43002 );
and ( n43508 , n30299 , n43172 );
and ( n43509 , n43507 , n43508 );
xor ( n43510 , n43507 , n43508 );
xor ( n43511 , n42870 , n43000 );
and ( n43512 , n30304 , n43172 );
and ( n43513 , n43511 , n43512 );
xor ( n43514 , n43511 , n43512 );
xor ( n43515 , n42874 , n42998 );
and ( n43516 , n30309 , n43172 );
and ( n43517 , n43515 , n43516 );
xor ( n43518 , n43515 , n43516 );
xor ( n43519 , n42878 , n42996 );
and ( n43520 , n30314 , n43172 );
and ( n43521 , n43519 , n43520 );
xor ( n43522 , n43519 , n43520 );
xor ( n43523 , n42882 , n42994 );
and ( n43524 , n30319 , n43172 );
and ( n43525 , n43523 , n43524 );
xor ( n43526 , n43523 , n43524 );
xor ( n43527 , n42886 , n42992 );
and ( n43528 , n30324 , n43172 );
and ( n43529 , n43527 , n43528 );
xor ( n43530 , n43527 , n43528 );
xor ( n43531 , n42890 , n42990 );
and ( n43532 , n30329 , n43172 );
and ( n43533 , n43531 , n43532 );
xor ( n43534 , n43531 , n43532 );
xor ( n43535 , n42894 , n42988 );
and ( n43536 , n30334 , n43172 );
and ( n43537 , n43535 , n43536 );
xor ( n43538 , n43535 , n43536 );
xor ( n43539 , n42898 , n42986 );
and ( n43540 , n30339 , n43172 );
and ( n43541 , n43539 , n43540 );
xor ( n43542 , n43539 , n43540 );
xor ( n43543 , n42902 , n42984 );
and ( n43544 , n30344 , n43172 );
and ( n43545 , n43543 , n43544 );
xor ( n43546 , n43543 , n43544 );
xor ( n43547 , n42906 , n42982 );
and ( n43548 , n30349 , n43172 );
and ( n43549 , n43547 , n43548 );
xor ( n43550 , n43547 , n43548 );
xor ( n43551 , n42910 , n42980 );
and ( n43552 , n30354 , n43172 );
and ( n43553 , n43551 , n43552 );
xor ( n43554 , n43551 , n43552 );
xor ( n43555 , n42914 , n42978 );
and ( n43556 , n30359 , n43172 );
and ( n43557 , n43555 , n43556 );
xor ( n43558 , n43555 , n43556 );
xor ( n43559 , n42918 , n42976 );
and ( n43560 , n30364 , n43172 );
and ( n43561 , n43559 , n43560 );
xor ( n43562 , n43559 , n43560 );
xor ( n43563 , n42922 , n42974 );
and ( n43564 , n30369 , n43172 );
and ( n43565 , n43563 , n43564 );
xor ( n43566 , n43563 , n43564 );
xor ( n43567 , n42926 , n42972 );
and ( n43568 , n30374 , n43172 );
and ( n43569 , n43567 , n43568 );
xor ( n43570 , n43567 , n43568 );
xor ( n43571 , n42930 , n42970 );
and ( n43572 , n30379 , n43172 );
and ( n43573 , n43571 , n43572 );
xor ( n43574 , n43571 , n43572 );
xor ( n43575 , n42934 , n42968 );
and ( n43576 , n30384 , n43172 );
and ( n43577 , n43575 , n43576 );
xor ( n43578 , n43575 , n43576 );
xor ( n43579 , n42938 , n42966 );
and ( n43580 , n30389 , n43172 );
and ( n43581 , n43579 , n43580 );
xor ( n43582 , n43579 , n43580 );
xor ( n43583 , n42942 , n42964 );
and ( n43584 , n30394 , n43172 );
and ( n43585 , n43583 , n43584 );
xor ( n43586 , n43583 , n43584 );
xor ( n43587 , n42946 , n42962 );
and ( n43588 , n30399 , n43172 );
and ( n43589 , n43587 , n43588 );
xor ( n43590 , n43587 , n43588 );
xor ( n43591 , n42950 , n42960 );
and ( n43592 , n30404 , n43172 );
and ( n43593 , n43591 , n43592 );
xor ( n43594 , n43591 , n43592 );
xor ( n43595 , n42954 , n42958 );
and ( n43596 , n30409 , n43172 );
and ( n43597 , n43595 , n43596 );
buf ( n43598 , n43597 );
and ( n43599 , n43594 , n43598 );
or ( n43600 , n43593 , n43599 );
and ( n43601 , n43590 , n43600 );
or ( n43602 , n43589 , n43601 );
and ( n43603 , n43586 , n43602 );
or ( n43604 , n43585 , n43603 );
and ( n43605 , n43582 , n43604 );
or ( n43606 , n43581 , n43605 );
and ( n43607 , n43578 , n43606 );
or ( n43608 , n43577 , n43607 );
and ( n43609 , n43574 , n43608 );
or ( n43610 , n43573 , n43609 );
and ( n43611 , n43570 , n43610 );
or ( n43612 , n43569 , n43611 );
and ( n43613 , n43566 , n43612 );
or ( n43614 , n43565 , n43613 );
and ( n43615 , n43562 , n43614 );
or ( n43616 , n43561 , n43615 );
and ( n43617 , n43558 , n43616 );
or ( n43618 , n43557 , n43617 );
and ( n43619 , n43554 , n43618 );
or ( n43620 , n43553 , n43619 );
and ( n43621 , n43550 , n43620 );
or ( n43622 , n43549 , n43621 );
and ( n43623 , n43546 , n43622 );
or ( n43624 , n43545 , n43623 );
and ( n43625 , n43542 , n43624 );
or ( n43626 , n43541 , n43625 );
and ( n43627 , n43538 , n43626 );
or ( n43628 , n43537 , n43627 );
and ( n43629 , n43534 , n43628 );
or ( n43630 , n43533 , n43629 );
and ( n43631 , n43530 , n43630 );
or ( n43632 , n43529 , n43631 );
and ( n43633 , n43526 , n43632 );
or ( n43634 , n43525 , n43633 );
and ( n43635 , n43522 , n43634 );
or ( n43636 , n43521 , n43635 );
and ( n43637 , n43518 , n43636 );
or ( n43638 , n43517 , n43637 );
and ( n43639 , n43514 , n43638 );
or ( n43640 , n43513 , n43639 );
and ( n43641 , n43510 , n43640 );
or ( n43642 , n43509 , n43641 );
and ( n43643 , n43506 , n43642 );
or ( n43644 , n43505 , n43643 );
and ( n43645 , n43502 , n43644 );
or ( n43646 , n43501 , n43645 );
and ( n43647 , n43498 , n43646 );
or ( n43648 , n43497 , n43647 );
and ( n43649 , n43494 , n43648 );
or ( n43650 , n43493 , n43649 );
and ( n43651 , n43490 , n43650 );
or ( n43652 , n43489 , n43651 );
and ( n43653 , n43486 , n43652 );
or ( n43654 , n43485 , n43653 );
and ( n43655 , n43482 , n43654 );
or ( n43656 , n43481 , n43655 );
and ( n43657 , n43478 , n43656 );
or ( n43658 , n43477 , n43657 );
and ( n43659 , n43474 , n43658 );
or ( n43660 , n43473 , n43659 );
and ( n43661 , n43470 , n43660 );
or ( n43662 , n43469 , n43661 );
and ( n43663 , n43466 , n43662 );
or ( n43664 , n43465 , n43663 );
and ( n43665 , n43462 , n43664 );
or ( n43666 , n43461 , n43665 );
and ( n43667 , n43458 , n43666 );
or ( n43668 , n43457 , n43667 );
and ( n43669 , n43454 , n43668 );
or ( n43670 , n43453 , n43669 );
and ( n43671 , n43450 , n43670 );
or ( n43672 , n43449 , n43671 );
and ( n43673 , n43446 , n43672 );
or ( n43674 , n43445 , n43673 );
and ( n43675 , n43442 , n43674 );
or ( n43676 , n43441 , n43675 );
and ( n43677 , n43438 , n43676 );
or ( n43678 , n43437 , n43677 );
and ( n43679 , n43434 , n43678 );
or ( n43680 , n43433 , n43679 );
and ( n43681 , n43430 , n43680 );
or ( n43682 , n43429 , n43681 );
and ( n43683 , n43426 , n43682 );
or ( n43684 , n43425 , n43683 );
and ( n43685 , n43422 , n43684 );
or ( n43686 , n43421 , n43685 );
and ( n43687 , n43418 , n43686 );
or ( n43688 , n43417 , n43687 );
and ( n43689 , n43414 , n43688 );
or ( n43690 , n43413 , n43689 );
and ( n43691 , n43410 , n43690 );
or ( n43692 , n43409 , n43691 );
and ( n43693 , n43406 , n43692 );
or ( n43694 , n43405 , n43693 );
and ( n43695 , n43402 , n43694 );
or ( n43696 , n43401 , n43695 );
and ( n43697 , n43398 , n43696 );
or ( n43698 , n43397 , n43697 );
and ( n43699 , n43394 , n43698 );
or ( n43700 , n43393 , n43699 );
and ( n43701 , n43390 , n43700 );
or ( n43702 , n43389 , n43701 );
and ( n43703 , n43386 , n43702 );
or ( n43704 , n43385 , n43703 );
and ( n43705 , n43382 , n43704 );
or ( n43706 , n43381 , n43705 );
and ( n43707 , n43378 , n43706 );
or ( n43708 , n43377 , n43707 );
and ( n43709 , n43374 , n43708 );
or ( n43710 , n43373 , n43709 );
and ( n43711 , n43370 , n43710 );
or ( n43712 , n43369 , n43711 );
and ( n43713 , n43366 , n43712 );
or ( n43714 , n43365 , n43713 );
and ( n43715 , n43362 , n43714 );
or ( n43716 , n43361 , n43715 );
and ( n43717 , n43358 , n43716 );
or ( n43718 , n43357 , n43717 );
and ( n43719 , n43354 , n43718 );
or ( n43720 , n43353 , n43719 );
and ( n43721 , n43350 , n43720 );
or ( n43722 , n43349 , n43721 );
and ( n43723 , n43346 , n43722 );
or ( n43724 , n43345 , n43723 );
and ( n43725 , n43342 , n43724 );
or ( n43726 , n43341 , n43725 );
and ( n43727 , n43338 , n43726 );
or ( n43728 , n43337 , n43727 );
and ( n43729 , n43334 , n43728 );
or ( n43730 , n43333 , n43729 );
and ( n43731 , n43330 , n43730 );
or ( n43732 , n43329 , n43731 );
and ( n43733 , n43326 , n43732 );
or ( n43734 , n43325 , n43733 );
and ( n43735 , n43322 , n43734 );
or ( n43736 , n43321 , n43735 );
and ( n43737 , n43318 , n43736 );
or ( n43738 , n43317 , n43737 );
and ( n43739 , n43314 , n43738 );
or ( n43740 , n43313 , n43739 );
and ( n43741 , n43310 , n43740 );
or ( n43742 , n43309 , n43741 );
and ( n43743 , n43306 , n43742 );
or ( n43744 , n43305 , n43743 );
and ( n43745 , n43302 , n43744 );
or ( n43746 , n43301 , n43745 );
and ( n43747 , n43298 , n43746 );
or ( n43748 , n43297 , n43747 );
and ( n43749 , n43294 , n43748 );
or ( n43750 , n43293 , n43749 );
and ( n43751 , n43290 , n43750 );
or ( n43752 , n43289 , n43751 );
and ( n43753 , n43286 , n43752 );
or ( n43754 , n43285 , n43753 );
and ( n43755 , n43282 , n43754 );
or ( n43756 , n43281 , n43755 );
and ( n43757 , n43278 , n43756 );
or ( n43758 , n43277 , n43757 );
and ( n43759 , n43274 , n43758 );
or ( n43760 , n43273 , n43759 );
and ( n43761 , n43270 , n43760 );
or ( n43762 , n43269 , n43761 );
and ( n43763 , n43266 , n43762 );
or ( n43764 , n43265 , n43763 );
and ( n43765 , n43262 , n43764 );
or ( n43766 , n43261 , n43765 );
and ( n43767 , n43258 , n43766 );
or ( n43768 , n43257 , n43767 );
and ( n43769 , n43254 , n43768 );
or ( n43770 , n43253 , n43769 );
and ( n43771 , n43250 , n43770 );
or ( n43772 , n43249 , n43771 );
and ( n43773 , n43246 , n43772 );
or ( n43774 , n43245 , n43773 );
and ( n43775 , n43242 , n43774 );
or ( n43776 , n43241 , n43775 );
and ( n43777 , n43238 , n43776 );
or ( n43778 , n43237 , n43777 );
and ( n43779 , n43234 , n43778 );
or ( n43780 , n43233 , n43779 );
and ( n43781 , n43230 , n43780 );
or ( n43782 , n43229 , n43781 );
and ( n43783 , n43226 , n43782 );
or ( n43784 , n43225 , n43783 );
and ( n43785 , n43222 , n43784 );
or ( n43786 , n43221 , n43785 );
and ( n43787 , n43218 , n43786 );
or ( n43788 , n43217 , n43787 );
and ( n43789 , n43214 , n43788 );
or ( n43790 , n43213 , n43789 );
and ( n43791 , n43210 , n43790 );
or ( n43792 , n43209 , n43791 );
and ( n43793 , n43206 , n43792 );
or ( n43794 , n43205 , n43793 );
and ( n43795 , n43202 , n43794 );
or ( n43796 , n43201 , n43795 );
and ( n43797 , n43198 , n43796 );
or ( n43798 , n43197 , n43797 );
and ( n43799 , n43194 , n43798 );
or ( n43800 , n43193 , n43799 );
and ( n43801 , n43190 , n43800 );
or ( n43802 , n43189 , n43801 );
and ( n43803 , n43186 , n43802 );
or ( n43804 , n43185 , n43803 );
and ( n43805 , n43182 , n43804 );
or ( n43806 , n43181 , n43805 );
and ( n43807 , n43178 , n43806 );
or ( n43808 , n43177 , n43807 );
xor ( n43809 , n43174 , n43808 );
buf ( n43810 , n18064 );
and ( n43811 , n29884 , n43810 );
xor ( n43812 , n43809 , n43811 );
xor ( n43813 , n43178 , n43806 );
and ( n43814 , n29889 , n43810 );
and ( n43815 , n43813 , n43814 );
xor ( n43816 , n43813 , n43814 );
xor ( n43817 , n43182 , n43804 );
and ( n43818 , n29894 , n43810 );
and ( n43819 , n43817 , n43818 );
xor ( n43820 , n43817 , n43818 );
xor ( n43821 , n43186 , n43802 );
and ( n43822 , n29899 , n43810 );
and ( n43823 , n43821 , n43822 );
xor ( n43824 , n43821 , n43822 );
xor ( n43825 , n43190 , n43800 );
and ( n43826 , n29904 , n43810 );
and ( n43827 , n43825 , n43826 );
xor ( n43828 , n43825 , n43826 );
xor ( n43829 , n43194 , n43798 );
and ( n43830 , n29909 , n43810 );
and ( n43831 , n43829 , n43830 );
xor ( n43832 , n43829 , n43830 );
xor ( n43833 , n43198 , n43796 );
and ( n43834 , n29914 , n43810 );
and ( n43835 , n43833 , n43834 );
xor ( n43836 , n43833 , n43834 );
xor ( n43837 , n43202 , n43794 );
and ( n43838 , n29919 , n43810 );
and ( n43839 , n43837 , n43838 );
xor ( n43840 , n43837 , n43838 );
xor ( n43841 , n43206 , n43792 );
and ( n43842 , n29924 , n43810 );
and ( n43843 , n43841 , n43842 );
xor ( n43844 , n43841 , n43842 );
xor ( n43845 , n43210 , n43790 );
and ( n43846 , n29929 , n43810 );
and ( n43847 , n43845 , n43846 );
xor ( n43848 , n43845 , n43846 );
xor ( n43849 , n43214 , n43788 );
and ( n43850 , n29934 , n43810 );
and ( n43851 , n43849 , n43850 );
xor ( n43852 , n43849 , n43850 );
xor ( n43853 , n43218 , n43786 );
and ( n43854 , n29939 , n43810 );
and ( n43855 , n43853 , n43854 );
xor ( n43856 , n43853 , n43854 );
xor ( n43857 , n43222 , n43784 );
and ( n43858 , n29944 , n43810 );
and ( n43859 , n43857 , n43858 );
xor ( n43860 , n43857 , n43858 );
xor ( n43861 , n43226 , n43782 );
and ( n43862 , n29949 , n43810 );
and ( n43863 , n43861 , n43862 );
xor ( n43864 , n43861 , n43862 );
xor ( n43865 , n43230 , n43780 );
and ( n43866 , n29954 , n43810 );
and ( n43867 , n43865 , n43866 );
xor ( n43868 , n43865 , n43866 );
xor ( n43869 , n43234 , n43778 );
and ( n43870 , n29959 , n43810 );
and ( n43871 , n43869 , n43870 );
xor ( n43872 , n43869 , n43870 );
xor ( n43873 , n43238 , n43776 );
and ( n43874 , n29964 , n43810 );
and ( n43875 , n43873 , n43874 );
xor ( n43876 , n43873 , n43874 );
xor ( n43877 , n43242 , n43774 );
and ( n43878 , n29969 , n43810 );
and ( n43879 , n43877 , n43878 );
xor ( n43880 , n43877 , n43878 );
xor ( n43881 , n43246 , n43772 );
and ( n43882 , n29974 , n43810 );
and ( n43883 , n43881 , n43882 );
xor ( n43884 , n43881 , n43882 );
xor ( n43885 , n43250 , n43770 );
and ( n43886 , n29979 , n43810 );
and ( n43887 , n43885 , n43886 );
xor ( n43888 , n43885 , n43886 );
xor ( n43889 , n43254 , n43768 );
and ( n43890 , n29984 , n43810 );
and ( n43891 , n43889 , n43890 );
xor ( n43892 , n43889 , n43890 );
xor ( n43893 , n43258 , n43766 );
and ( n43894 , n29989 , n43810 );
and ( n43895 , n43893 , n43894 );
xor ( n43896 , n43893 , n43894 );
xor ( n43897 , n43262 , n43764 );
and ( n43898 , n29994 , n43810 );
and ( n43899 , n43897 , n43898 );
xor ( n43900 , n43897 , n43898 );
xor ( n43901 , n43266 , n43762 );
and ( n43902 , n29999 , n43810 );
and ( n43903 , n43901 , n43902 );
xor ( n43904 , n43901 , n43902 );
xor ( n43905 , n43270 , n43760 );
and ( n43906 , n30004 , n43810 );
and ( n43907 , n43905 , n43906 );
xor ( n43908 , n43905 , n43906 );
xor ( n43909 , n43274 , n43758 );
and ( n43910 , n30009 , n43810 );
and ( n43911 , n43909 , n43910 );
xor ( n43912 , n43909 , n43910 );
xor ( n43913 , n43278 , n43756 );
and ( n43914 , n30014 , n43810 );
and ( n43915 , n43913 , n43914 );
xor ( n43916 , n43913 , n43914 );
xor ( n43917 , n43282 , n43754 );
and ( n43918 , n30019 , n43810 );
and ( n43919 , n43917 , n43918 );
xor ( n43920 , n43917 , n43918 );
xor ( n43921 , n43286 , n43752 );
and ( n43922 , n30024 , n43810 );
and ( n43923 , n43921 , n43922 );
xor ( n43924 , n43921 , n43922 );
xor ( n43925 , n43290 , n43750 );
and ( n43926 , n30029 , n43810 );
and ( n43927 , n43925 , n43926 );
xor ( n43928 , n43925 , n43926 );
xor ( n43929 , n43294 , n43748 );
and ( n43930 , n30034 , n43810 );
and ( n43931 , n43929 , n43930 );
xor ( n43932 , n43929 , n43930 );
xor ( n43933 , n43298 , n43746 );
and ( n43934 , n30039 , n43810 );
and ( n43935 , n43933 , n43934 );
xor ( n43936 , n43933 , n43934 );
xor ( n43937 , n43302 , n43744 );
and ( n43938 , n30044 , n43810 );
and ( n43939 , n43937 , n43938 );
xor ( n43940 , n43937 , n43938 );
xor ( n43941 , n43306 , n43742 );
and ( n43942 , n30049 , n43810 );
and ( n43943 , n43941 , n43942 );
xor ( n43944 , n43941 , n43942 );
xor ( n43945 , n43310 , n43740 );
and ( n43946 , n30054 , n43810 );
and ( n43947 , n43945 , n43946 );
xor ( n43948 , n43945 , n43946 );
xor ( n43949 , n43314 , n43738 );
and ( n43950 , n30059 , n43810 );
and ( n43951 , n43949 , n43950 );
xor ( n43952 , n43949 , n43950 );
xor ( n43953 , n43318 , n43736 );
and ( n43954 , n30064 , n43810 );
and ( n43955 , n43953 , n43954 );
xor ( n43956 , n43953 , n43954 );
xor ( n43957 , n43322 , n43734 );
and ( n43958 , n30069 , n43810 );
and ( n43959 , n43957 , n43958 );
xor ( n43960 , n43957 , n43958 );
xor ( n43961 , n43326 , n43732 );
and ( n43962 , n30074 , n43810 );
and ( n43963 , n43961 , n43962 );
xor ( n43964 , n43961 , n43962 );
xor ( n43965 , n43330 , n43730 );
and ( n43966 , n30079 , n43810 );
and ( n43967 , n43965 , n43966 );
xor ( n43968 , n43965 , n43966 );
xor ( n43969 , n43334 , n43728 );
and ( n43970 , n30084 , n43810 );
and ( n43971 , n43969 , n43970 );
xor ( n43972 , n43969 , n43970 );
xor ( n43973 , n43338 , n43726 );
and ( n43974 , n30089 , n43810 );
and ( n43975 , n43973 , n43974 );
xor ( n43976 , n43973 , n43974 );
xor ( n43977 , n43342 , n43724 );
and ( n43978 , n30094 , n43810 );
and ( n43979 , n43977 , n43978 );
xor ( n43980 , n43977 , n43978 );
xor ( n43981 , n43346 , n43722 );
and ( n43982 , n30099 , n43810 );
and ( n43983 , n43981 , n43982 );
xor ( n43984 , n43981 , n43982 );
xor ( n43985 , n43350 , n43720 );
and ( n43986 , n30104 , n43810 );
and ( n43987 , n43985 , n43986 );
xor ( n43988 , n43985 , n43986 );
xor ( n43989 , n43354 , n43718 );
and ( n43990 , n30109 , n43810 );
and ( n43991 , n43989 , n43990 );
xor ( n43992 , n43989 , n43990 );
xor ( n43993 , n43358 , n43716 );
and ( n43994 , n30114 , n43810 );
and ( n43995 , n43993 , n43994 );
xor ( n43996 , n43993 , n43994 );
xor ( n43997 , n43362 , n43714 );
and ( n43998 , n30119 , n43810 );
and ( n43999 , n43997 , n43998 );
xor ( n44000 , n43997 , n43998 );
xor ( n44001 , n43366 , n43712 );
and ( n44002 , n30124 , n43810 );
and ( n44003 , n44001 , n44002 );
xor ( n44004 , n44001 , n44002 );
xor ( n44005 , n43370 , n43710 );
and ( n44006 , n30129 , n43810 );
and ( n44007 , n44005 , n44006 );
xor ( n44008 , n44005 , n44006 );
xor ( n44009 , n43374 , n43708 );
and ( n44010 , n30134 , n43810 );
and ( n44011 , n44009 , n44010 );
xor ( n44012 , n44009 , n44010 );
xor ( n44013 , n43378 , n43706 );
and ( n44014 , n30139 , n43810 );
and ( n44015 , n44013 , n44014 );
xor ( n44016 , n44013 , n44014 );
xor ( n44017 , n43382 , n43704 );
and ( n44018 , n30144 , n43810 );
and ( n44019 , n44017 , n44018 );
xor ( n44020 , n44017 , n44018 );
xor ( n44021 , n43386 , n43702 );
and ( n44022 , n30149 , n43810 );
and ( n44023 , n44021 , n44022 );
xor ( n44024 , n44021 , n44022 );
xor ( n44025 , n43390 , n43700 );
and ( n44026 , n30154 , n43810 );
and ( n44027 , n44025 , n44026 );
xor ( n44028 , n44025 , n44026 );
xor ( n44029 , n43394 , n43698 );
and ( n44030 , n30159 , n43810 );
and ( n44031 , n44029 , n44030 );
xor ( n44032 , n44029 , n44030 );
xor ( n44033 , n43398 , n43696 );
and ( n44034 , n30164 , n43810 );
and ( n44035 , n44033 , n44034 );
xor ( n44036 , n44033 , n44034 );
xor ( n44037 , n43402 , n43694 );
and ( n44038 , n30169 , n43810 );
and ( n44039 , n44037 , n44038 );
xor ( n44040 , n44037 , n44038 );
xor ( n44041 , n43406 , n43692 );
and ( n44042 , n30174 , n43810 );
and ( n44043 , n44041 , n44042 );
xor ( n44044 , n44041 , n44042 );
xor ( n44045 , n43410 , n43690 );
and ( n44046 , n30179 , n43810 );
and ( n44047 , n44045 , n44046 );
xor ( n44048 , n44045 , n44046 );
xor ( n44049 , n43414 , n43688 );
and ( n44050 , n30184 , n43810 );
and ( n44051 , n44049 , n44050 );
xor ( n44052 , n44049 , n44050 );
xor ( n44053 , n43418 , n43686 );
and ( n44054 , n30189 , n43810 );
and ( n44055 , n44053 , n44054 );
xor ( n44056 , n44053 , n44054 );
xor ( n44057 , n43422 , n43684 );
and ( n44058 , n30194 , n43810 );
and ( n44059 , n44057 , n44058 );
xor ( n44060 , n44057 , n44058 );
xor ( n44061 , n43426 , n43682 );
and ( n44062 , n30199 , n43810 );
and ( n44063 , n44061 , n44062 );
xor ( n44064 , n44061 , n44062 );
xor ( n44065 , n43430 , n43680 );
and ( n44066 , n30204 , n43810 );
and ( n44067 , n44065 , n44066 );
xor ( n44068 , n44065 , n44066 );
xor ( n44069 , n43434 , n43678 );
and ( n44070 , n30209 , n43810 );
and ( n44071 , n44069 , n44070 );
xor ( n44072 , n44069 , n44070 );
xor ( n44073 , n43438 , n43676 );
and ( n44074 , n30214 , n43810 );
and ( n44075 , n44073 , n44074 );
xor ( n44076 , n44073 , n44074 );
xor ( n44077 , n43442 , n43674 );
and ( n44078 , n30219 , n43810 );
and ( n44079 , n44077 , n44078 );
xor ( n44080 , n44077 , n44078 );
xor ( n44081 , n43446 , n43672 );
and ( n44082 , n30224 , n43810 );
and ( n44083 , n44081 , n44082 );
xor ( n44084 , n44081 , n44082 );
xor ( n44085 , n43450 , n43670 );
and ( n44086 , n30229 , n43810 );
and ( n44087 , n44085 , n44086 );
xor ( n44088 , n44085 , n44086 );
xor ( n44089 , n43454 , n43668 );
and ( n44090 , n30234 , n43810 );
and ( n44091 , n44089 , n44090 );
xor ( n44092 , n44089 , n44090 );
xor ( n44093 , n43458 , n43666 );
and ( n44094 , n30239 , n43810 );
and ( n44095 , n44093 , n44094 );
xor ( n44096 , n44093 , n44094 );
xor ( n44097 , n43462 , n43664 );
and ( n44098 , n30244 , n43810 );
and ( n44099 , n44097 , n44098 );
xor ( n44100 , n44097 , n44098 );
xor ( n44101 , n43466 , n43662 );
and ( n44102 , n30249 , n43810 );
and ( n44103 , n44101 , n44102 );
xor ( n44104 , n44101 , n44102 );
xor ( n44105 , n43470 , n43660 );
and ( n44106 , n30254 , n43810 );
and ( n44107 , n44105 , n44106 );
xor ( n44108 , n44105 , n44106 );
xor ( n44109 , n43474 , n43658 );
and ( n44110 , n30259 , n43810 );
and ( n44111 , n44109 , n44110 );
xor ( n44112 , n44109 , n44110 );
xor ( n44113 , n43478 , n43656 );
and ( n44114 , n30264 , n43810 );
and ( n44115 , n44113 , n44114 );
xor ( n44116 , n44113 , n44114 );
xor ( n44117 , n43482 , n43654 );
and ( n44118 , n30269 , n43810 );
and ( n44119 , n44117 , n44118 );
xor ( n44120 , n44117 , n44118 );
xor ( n44121 , n43486 , n43652 );
and ( n44122 , n30274 , n43810 );
and ( n44123 , n44121 , n44122 );
xor ( n44124 , n44121 , n44122 );
xor ( n44125 , n43490 , n43650 );
and ( n44126 , n30279 , n43810 );
and ( n44127 , n44125 , n44126 );
xor ( n44128 , n44125 , n44126 );
xor ( n44129 , n43494 , n43648 );
and ( n44130 , n30284 , n43810 );
and ( n44131 , n44129 , n44130 );
xor ( n44132 , n44129 , n44130 );
xor ( n44133 , n43498 , n43646 );
and ( n44134 , n30289 , n43810 );
and ( n44135 , n44133 , n44134 );
xor ( n44136 , n44133 , n44134 );
xor ( n44137 , n43502 , n43644 );
and ( n44138 , n30294 , n43810 );
and ( n44139 , n44137 , n44138 );
xor ( n44140 , n44137 , n44138 );
xor ( n44141 , n43506 , n43642 );
and ( n44142 , n30299 , n43810 );
and ( n44143 , n44141 , n44142 );
xor ( n44144 , n44141 , n44142 );
xor ( n44145 , n43510 , n43640 );
and ( n44146 , n30304 , n43810 );
and ( n44147 , n44145 , n44146 );
xor ( n44148 , n44145 , n44146 );
xor ( n44149 , n43514 , n43638 );
and ( n44150 , n30309 , n43810 );
and ( n44151 , n44149 , n44150 );
xor ( n44152 , n44149 , n44150 );
xor ( n44153 , n43518 , n43636 );
and ( n44154 , n30314 , n43810 );
and ( n44155 , n44153 , n44154 );
xor ( n44156 , n44153 , n44154 );
xor ( n44157 , n43522 , n43634 );
and ( n44158 , n30319 , n43810 );
and ( n44159 , n44157 , n44158 );
xor ( n44160 , n44157 , n44158 );
xor ( n44161 , n43526 , n43632 );
and ( n44162 , n30324 , n43810 );
and ( n44163 , n44161 , n44162 );
xor ( n44164 , n44161 , n44162 );
xor ( n44165 , n43530 , n43630 );
and ( n44166 , n30329 , n43810 );
and ( n44167 , n44165 , n44166 );
xor ( n44168 , n44165 , n44166 );
xor ( n44169 , n43534 , n43628 );
and ( n44170 , n30334 , n43810 );
and ( n44171 , n44169 , n44170 );
xor ( n44172 , n44169 , n44170 );
xor ( n44173 , n43538 , n43626 );
and ( n44174 , n30339 , n43810 );
and ( n44175 , n44173 , n44174 );
xor ( n44176 , n44173 , n44174 );
xor ( n44177 , n43542 , n43624 );
and ( n44178 , n30344 , n43810 );
and ( n44179 , n44177 , n44178 );
xor ( n44180 , n44177 , n44178 );
xor ( n44181 , n43546 , n43622 );
and ( n44182 , n30349 , n43810 );
and ( n44183 , n44181 , n44182 );
xor ( n44184 , n44181 , n44182 );
xor ( n44185 , n43550 , n43620 );
and ( n44186 , n30354 , n43810 );
and ( n44187 , n44185 , n44186 );
xor ( n44188 , n44185 , n44186 );
xor ( n44189 , n43554 , n43618 );
and ( n44190 , n30359 , n43810 );
and ( n44191 , n44189 , n44190 );
xor ( n44192 , n44189 , n44190 );
xor ( n44193 , n43558 , n43616 );
and ( n44194 , n30364 , n43810 );
and ( n44195 , n44193 , n44194 );
xor ( n44196 , n44193 , n44194 );
xor ( n44197 , n43562 , n43614 );
and ( n44198 , n30369 , n43810 );
and ( n44199 , n44197 , n44198 );
xor ( n44200 , n44197 , n44198 );
xor ( n44201 , n43566 , n43612 );
and ( n44202 , n30374 , n43810 );
and ( n44203 , n44201 , n44202 );
xor ( n44204 , n44201 , n44202 );
xor ( n44205 , n43570 , n43610 );
and ( n44206 , n30379 , n43810 );
and ( n44207 , n44205 , n44206 );
xor ( n44208 , n44205 , n44206 );
xor ( n44209 , n43574 , n43608 );
and ( n44210 , n30384 , n43810 );
and ( n44211 , n44209 , n44210 );
xor ( n44212 , n44209 , n44210 );
xor ( n44213 , n43578 , n43606 );
and ( n44214 , n30389 , n43810 );
and ( n44215 , n44213 , n44214 );
xor ( n44216 , n44213 , n44214 );
xor ( n44217 , n43582 , n43604 );
and ( n44218 , n30394 , n43810 );
and ( n44219 , n44217 , n44218 );
xor ( n44220 , n44217 , n44218 );
xor ( n44221 , n43586 , n43602 );
and ( n44222 , n30399 , n43810 );
and ( n44223 , n44221 , n44222 );
xor ( n44224 , n44221 , n44222 );
xor ( n44225 , n43590 , n43600 );
and ( n44226 , n30404 , n43810 );
and ( n44227 , n44225 , n44226 );
xor ( n44228 , n44225 , n44226 );
xor ( n44229 , n43594 , n43598 );
and ( n44230 , n30409 , n43810 );
and ( n44231 , n44229 , n44230 );
buf ( n44232 , n44231 );
and ( n44233 , n44228 , n44232 );
or ( n44234 , n44227 , n44233 );
and ( n44235 , n44224 , n44234 );
or ( n44236 , n44223 , n44235 );
and ( n44237 , n44220 , n44236 );
or ( n44238 , n44219 , n44237 );
and ( n44239 , n44216 , n44238 );
or ( n44240 , n44215 , n44239 );
and ( n44241 , n44212 , n44240 );
or ( n44242 , n44211 , n44241 );
and ( n44243 , n44208 , n44242 );
or ( n44244 , n44207 , n44243 );
and ( n44245 , n44204 , n44244 );
or ( n44246 , n44203 , n44245 );
and ( n44247 , n44200 , n44246 );
or ( n44248 , n44199 , n44247 );
and ( n44249 , n44196 , n44248 );
or ( n44250 , n44195 , n44249 );
and ( n44251 , n44192 , n44250 );
or ( n44252 , n44191 , n44251 );
and ( n44253 , n44188 , n44252 );
or ( n44254 , n44187 , n44253 );
and ( n44255 , n44184 , n44254 );
or ( n44256 , n44183 , n44255 );
and ( n44257 , n44180 , n44256 );
or ( n44258 , n44179 , n44257 );
and ( n44259 , n44176 , n44258 );
or ( n44260 , n44175 , n44259 );
and ( n44261 , n44172 , n44260 );
or ( n44262 , n44171 , n44261 );
and ( n44263 , n44168 , n44262 );
or ( n44264 , n44167 , n44263 );
and ( n44265 , n44164 , n44264 );
or ( n44266 , n44163 , n44265 );
and ( n44267 , n44160 , n44266 );
or ( n44268 , n44159 , n44267 );
and ( n44269 , n44156 , n44268 );
or ( n44270 , n44155 , n44269 );
and ( n44271 , n44152 , n44270 );
or ( n44272 , n44151 , n44271 );
and ( n44273 , n44148 , n44272 );
or ( n44274 , n44147 , n44273 );
and ( n44275 , n44144 , n44274 );
or ( n44276 , n44143 , n44275 );
and ( n44277 , n44140 , n44276 );
or ( n44278 , n44139 , n44277 );
and ( n44279 , n44136 , n44278 );
or ( n44280 , n44135 , n44279 );
and ( n44281 , n44132 , n44280 );
or ( n44282 , n44131 , n44281 );
and ( n44283 , n44128 , n44282 );
or ( n44284 , n44127 , n44283 );
and ( n44285 , n44124 , n44284 );
or ( n44286 , n44123 , n44285 );
and ( n44287 , n44120 , n44286 );
or ( n44288 , n44119 , n44287 );
and ( n44289 , n44116 , n44288 );
or ( n44290 , n44115 , n44289 );
and ( n44291 , n44112 , n44290 );
or ( n44292 , n44111 , n44291 );
and ( n44293 , n44108 , n44292 );
or ( n44294 , n44107 , n44293 );
and ( n44295 , n44104 , n44294 );
or ( n44296 , n44103 , n44295 );
and ( n44297 , n44100 , n44296 );
or ( n44298 , n44099 , n44297 );
and ( n44299 , n44096 , n44298 );
or ( n44300 , n44095 , n44299 );
and ( n44301 , n44092 , n44300 );
or ( n44302 , n44091 , n44301 );
and ( n44303 , n44088 , n44302 );
or ( n44304 , n44087 , n44303 );
and ( n44305 , n44084 , n44304 );
or ( n44306 , n44083 , n44305 );
and ( n44307 , n44080 , n44306 );
or ( n44308 , n44079 , n44307 );
and ( n44309 , n44076 , n44308 );
or ( n44310 , n44075 , n44309 );
and ( n44311 , n44072 , n44310 );
or ( n44312 , n44071 , n44311 );
and ( n44313 , n44068 , n44312 );
or ( n44314 , n44067 , n44313 );
and ( n44315 , n44064 , n44314 );
or ( n44316 , n44063 , n44315 );
and ( n44317 , n44060 , n44316 );
or ( n44318 , n44059 , n44317 );
and ( n44319 , n44056 , n44318 );
or ( n44320 , n44055 , n44319 );
and ( n44321 , n44052 , n44320 );
or ( n44322 , n44051 , n44321 );
and ( n44323 , n44048 , n44322 );
or ( n44324 , n44047 , n44323 );
and ( n44325 , n44044 , n44324 );
or ( n44326 , n44043 , n44325 );
and ( n44327 , n44040 , n44326 );
or ( n44328 , n44039 , n44327 );
and ( n44329 , n44036 , n44328 );
or ( n44330 , n44035 , n44329 );
and ( n44331 , n44032 , n44330 );
or ( n44332 , n44031 , n44331 );
and ( n44333 , n44028 , n44332 );
or ( n44334 , n44027 , n44333 );
and ( n44335 , n44024 , n44334 );
or ( n44336 , n44023 , n44335 );
and ( n44337 , n44020 , n44336 );
or ( n44338 , n44019 , n44337 );
and ( n44339 , n44016 , n44338 );
or ( n44340 , n44015 , n44339 );
and ( n44341 , n44012 , n44340 );
or ( n44342 , n44011 , n44341 );
and ( n44343 , n44008 , n44342 );
or ( n44344 , n44007 , n44343 );
and ( n44345 , n44004 , n44344 );
or ( n44346 , n44003 , n44345 );
and ( n44347 , n44000 , n44346 );
or ( n44348 , n43999 , n44347 );
and ( n44349 , n43996 , n44348 );
or ( n44350 , n43995 , n44349 );
and ( n44351 , n43992 , n44350 );
or ( n44352 , n43991 , n44351 );
and ( n44353 , n43988 , n44352 );
or ( n44354 , n43987 , n44353 );
and ( n44355 , n43984 , n44354 );
or ( n44356 , n43983 , n44355 );
and ( n44357 , n43980 , n44356 );
or ( n44358 , n43979 , n44357 );
and ( n44359 , n43976 , n44358 );
or ( n44360 , n43975 , n44359 );
and ( n44361 , n43972 , n44360 );
or ( n44362 , n43971 , n44361 );
and ( n44363 , n43968 , n44362 );
or ( n44364 , n43967 , n44363 );
and ( n44365 , n43964 , n44364 );
or ( n44366 , n43963 , n44365 );
and ( n44367 , n43960 , n44366 );
or ( n44368 , n43959 , n44367 );
and ( n44369 , n43956 , n44368 );
or ( n44370 , n43955 , n44369 );
and ( n44371 , n43952 , n44370 );
or ( n44372 , n43951 , n44371 );
and ( n44373 , n43948 , n44372 );
or ( n44374 , n43947 , n44373 );
and ( n44375 , n43944 , n44374 );
or ( n44376 , n43943 , n44375 );
and ( n44377 , n43940 , n44376 );
or ( n44378 , n43939 , n44377 );
and ( n44379 , n43936 , n44378 );
or ( n44380 , n43935 , n44379 );
and ( n44381 , n43932 , n44380 );
or ( n44382 , n43931 , n44381 );
and ( n44383 , n43928 , n44382 );
or ( n44384 , n43927 , n44383 );
and ( n44385 , n43924 , n44384 );
or ( n44386 , n43923 , n44385 );
and ( n44387 , n43920 , n44386 );
or ( n44388 , n43919 , n44387 );
and ( n44389 , n43916 , n44388 );
or ( n44390 , n43915 , n44389 );
and ( n44391 , n43912 , n44390 );
or ( n44392 , n43911 , n44391 );
and ( n44393 , n43908 , n44392 );
or ( n44394 , n43907 , n44393 );
and ( n44395 , n43904 , n44394 );
or ( n44396 , n43903 , n44395 );
and ( n44397 , n43900 , n44396 );
or ( n44398 , n43899 , n44397 );
and ( n44399 , n43896 , n44398 );
or ( n44400 , n43895 , n44399 );
and ( n44401 , n43892 , n44400 );
or ( n44402 , n43891 , n44401 );
and ( n44403 , n43888 , n44402 );
or ( n44404 , n43887 , n44403 );
and ( n44405 , n43884 , n44404 );
or ( n44406 , n43883 , n44405 );
and ( n44407 , n43880 , n44406 );
or ( n44408 , n43879 , n44407 );
and ( n44409 , n43876 , n44408 );
or ( n44410 , n43875 , n44409 );
and ( n44411 , n43872 , n44410 );
or ( n44412 , n43871 , n44411 );
and ( n44413 , n43868 , n44412 );
or ( n44414 , n43867 , n44413 );
and ( n44415 , n43864 , n44414 );
or ( n44416 , n43863 , n44415 );
and ( n44417 , n43860 , n44416 );
or ( n44418 , n43859 , n44417 );
and ( n44419 , n43856 , n44418 );
or ( n44420 , n43855 , n44419 );
and ( n44421 , n43852 , n44420 );
or ( n44422 , n43851 , n44421 );
and ( n44423 , n43848 , n44422 );
or ( n44424 , n43847 , n44423 );
and ( n44425 , n43844 , n44424 );
or ( n44426 , n43843 , n44425 );
and ( n44427 , n43840 , n44426 );
or ( n44428 , n43839 , n44427 );
and ( n44429 , n43836 , n44428 );
or ( n44430 , n43835 , n44429 );
and ( n44431 , n43832 , n44430 );
or ( n44432 , n43831 , n44431 );
and ( n44433 , n43828 , n44432 );
or ( n44434 , n43827 , n44433 );
and ( n44435 , n43824 , n44434 );
or ( n44436 , n43823 , n44435 );
and ( n44437 , n43820 , n44436 );
or ( n44438 , n43819 , n44437 );
and ( n44439 , n43816 , n44438 );
or ( n44440 , n43815 , n44439 );
xor ( n44441 , n43812 , n44440 );
buf ( n44442 , n18062 );
and ( n44443 , n29889 , n44442 );
xor ( n44444 , n44441 , n44443 );
xor ( n44445 , n43816 , n44438 );
and ( n44446 , n29894 , n44442 );
and ( n44447 , n44445 , n44446 );
xor ( n44448 , n44445 , n44446 );
xor ( n44449 , n43820 , n44436 );
and ( n44450 , n29899 , n44442 );
and ( n44451 , n44449 , n44450 );
xor ( n44452 , n44449 , n44450 );
xor ( n44453 , n43824 , n44434 );
and ( n44454 , n29904 , n44442 );
and ( n44455 , n44453 , n44454 );
xor ( n44456 , n44453 , n44454 );
xor ( n44457 , n43828 , n44432 );
and ( n44458 , n29909 , n44442 );
and ( n44459 , n44457 , n44458 );
xor ( n44460 , n44457 , n44458 );
xor ( n44461 , n43832 , n44430 );
and ( n44462 , n29914 , n44442 );
and ( n44463 , n44461 , n44462 );
xor ( n44464 , n44461 , n44462 );
xor ( n44465 , n43836 , n44428 );
and ( n44466 , n29919 , n44442 );
and ( n44467 , n44465 , n44466 );
xor ( n44468 , n44465 , n44466 );
xor ( n44469 , n43840 , n44426 );
and ( n44470 , n29924 , n44442 );
and ( n44471 , n44469 , n44470 );
xor ( n44472 , n44469 , n44470 );
xor ( n44473 , n43844 , n44424 );
and ( n44474 , n29929 , n44442 );
and ( n44475 , n44473 , n44474 );
xor ( n44476 , n44473 , n44474 );
xor ( n44477 , n43848 , n44422 );
and ( n44478 , n29934 , n44442 );
and ( n44479 , n44477 , n44478 );
xor ( n44480 , n44477 , n44478 );
xor ( n44481 , n43852 , n44420 );
and ( n44482 , n29939 , n44442 );
and ( n44483 , n44481 , n44482 );
xor ( n44484 , n44481 , n44482 );
xor ( n44485 , n43856 , n44418 );
and ( n44486 , n29944 , n44442 );
and ( n44487 , n44485 , n44486 );
xor ( n44488 , n44485 , n44486 );
xor ( n44489 , n43860 , n44416 );
and ( n44490 , n29949 , n44442 );
and ( n44491 , n44489 , n44490 );
xor ( n44492 , n44489 , n44490 );
xor ( n44493 , n43864 , n44414 );
and ( n44494 , n29954 , n44442 );
and ( n44495 , n44493 , n44494 );
xor ( n44496 , n44493 , n44494 );
xor ( n44497 , n43868 , n44412 );
and ( n44498 , n29959 , n44442 );
and ( n44499 , n44497 , n44498 );
xor ( n44500 , n44497 , n44498 );
xor ( n44501 , n43872 , n44410 );
and ( n44502 , n29964 , n44442 );
and ( n44503 , n44501 , n44502 );
xor ( n44504 , n44501 , n44502 );
xor ( n44505 , n43876 , n44408 );
and ( n44506 , n29969 , n44442 );
and ( n44507 , n44505 , n44506 );
xor ( n44508 , n44505 , n44506 );
xor ( n44509 , n43880 , n44406 );
and ( n44510 , n29974 , n44442 );
and ( n44511 , n44509 , n44510 );
xor ( n44512 , n44509 , n44510 );
xor ( n44513 , n43884 , n44404 );
and ( n44514 , n29979 , n44442 );
and ( n44515 , n44513 , n44514 );
xor ( n44516 , n44513 , n44514 );
xor ( n44517 , n43888 , n44402 );
and ( n44518 , n29984 , n44442 );
and ( n44519 , n44517 , n44518 );
xor ( n44520 , n44517 , n44518 );
xor ( n44521 , n43892 , n44400 );
and ( n44522 , n29989 , n44442 );
and ( n44523 , n44521 , n44522 );
xor ( n44524 , n44521 , n44522 );
xor ( n44525 , n43896 , n44398 );
and ( n44526 , n29994 , n44442 );
and ( n44527 , n44525 , n44526 );
xor ( n44528 , n44525 , n44526 );
xor ( n44529 , n43900 , n44396 );
and ( n44530 , n29999 , n44442 );
and ( n44531 , n44529 , n44530 );
xor ( n44532 , n44529 , n44530 );
xor ( n44533 , n43904 , n44394 );
and ( n44534 , n30004 , n44442 );
and ( n44535 , n44533 , n44534 );
xor ( n44536 , n44533 , n44534 );
xor ( n44537 , n43908 , n44392 );
and ( n44538 , n30009 , n44442 );
and ( n44539 , n44537 , n44538 );
xor ( n44540 , n44537 , n44538 );
xor ( n44541 , n43912 , n44390 );
and ( n44542 , n30014 , n44442 );
and ( n44543 , n44541 , n44542 );
xor ( n44544 , n44541 , n44542 );
xor ( n44545 , n43916 , n44388 );
and ( n44546 , n30019 , n44442 );
and ( n44547 , n44545 , n44546 );
xor ( n44548 , n44545 , n44546 );
xor ( n44549 , n43920 , n44386 );
and ( n44550 , n30024 , n44442 );
and ( n44551 , n44549 , n44550 );
xor ( n44552 , n44549 , n44550 );
xor ( n44553 , n43924 , n44384 );
and ( n44554 , n30029 , n44442 );
and ( n44555 , n44553 , n44554 );
xor ( n44556 , n44553 , n44554 );
xor ( n44557 , n43928 , n44382 );
and ( n44558 , n30034 , n44442 );
and ( n44559 , n44557 , n44558 );
xor ( n44560 , n44557 , n44558 );
xor ( n44561 , n43932 , n44380 );
and ( n44562 , n30039 , n44442 );
and ( n44563 , n44561 , n44562 );
xor ( n44564 , n44561 , n44562 );
xor ( n44565 , n43936 , n44378 );
and ( n44566 , n30044 , n44442 );
and ( n44567 , n44565 , n44566 );
xor ( n44568 , n44565 , n44566 );
xor ( n44569 , n43940 , n44376 );
and ( n44570 , n30049 , n44442 );
and ( n44571 , n44569 , n44570 );
xor ( n44572 , n44569 , n44570 );
xor ( n44573 , n43944 , n44374 );
and ( n44574 , n30054 , n44442 );
and ( n44575 , n44573 , n44574 );
xor ( n44576 , n44573 , n44574 );
xor ( n44577 , n43948 , n44372 );
and ( n44578 , n30059 , n44442 );
and ( n44579 , n44577 , n44578 );
xor ( n44580 , n44577 , n44578 );
xor ( n44581 , n43952 , n44370 );
and ( n44582 , n30064 , n44442 );
and ( n44583 , n44581 , n44582 );
xor ( n44584 , n44581 , n44582 );
xor ( n44585 , n43956 , n44368 );
and ( n44586 , n30069 , n44442 );
and ( n44587 , n44585 , n44586 );
xor ( n44588 , n44585 , n44586 );
xor ( n44589 , n43960 , n44366 );
and ( n44590 , n30074 , n44442 );
and ( n44591 , n44589 , n44590 );
xor ( n44592 , n44589 , n44590 );
xor ( n44593 , n43964 , n44364 );
and ( n44594 , n30079 , n44442 );
and ( n44595 , n44593 , n44594 );
xor ( n44596 , n44593 , n44594 );
xor ( n44597 , n43968 , n44362 );
and ( n44598 , n30084 , n44442 );
and ( n44599 , n44597 , n44598 );
xor ( n44600 , n44597 , n44598 );
xor ( n44601 , n43972 , n44360 );
and ( n44602 , n30089 , n44442 );
and ( n44603 , n44601 , n44602 );
xor ( n44604 , n44601 , n44602 );
xor ( n44605 , n43976 , n44358 );
and ( n44606 , n30094 , n44442 );
and ( n44607 , n44605 , n44606 );
xor ( n44608 , n44605 , n44606 );
xor ( n44609 , n43980 , n44356 );
and ( n44610 , n30099 , n44442 );
and ( n44611 , n44609 , n44610 );
xor ( n44612 , n44609 , n44610 );
xor ( n44613 , n43984 , n44354 );
and ( n44614 , n30104 , n44442 );
and ( n44615 , n44613 , n44614 );
xor ( n44616 , n44613 , n44614 );
xor ( n44617 , n43988 , n44352 );
and ( n44618 , n30109 , n44442 );
and ( n44619 , n44617 , n44618 );
xor ( n44620 , n44617 , n44618 );
xor ( n44621 , n43992 , n44350 );
and ( n44622 , n30114 , n44442 );
and ( n44623 , n44621 , n44622 );
xor ( n44624 , n44621 , n44622 );
xor ( n44625 , n43996 , n44348 );
and ( n44626 , n30119 , n44442 );
and ( n44627 , n44625 , n44626 );
xor ( n44628 , n44625 , n44626 );
xor ( n44629 , n44000 , n44346 );
and ( n44630 , n30124 , n44442 );
and ( n44631 , n44629 , n44630 );
xor ( n44632 , n44629 , n44630 );
xor ( n44633 , n44004 , n44344 );
and ( n44634 , n30129 , n44442 );
and ( n44635 , n44633 , n44634 );
xor ( n44636 , n44633 , n44634 );
xor ( n44637 , n44008 , n44342 );
and ( n44638 , n30134 , n44442 );
and ( n44639 , n44637 , n44638 );
xor ( n44640 , n44637 , n44638 );
xor ( n44641 , n44012 , n44340 );
and ( n44642 , n30139 , n44442 );
and ( n44643 , n44641 , n44642 );
xor ( n44644 , n44641 , n44642 );
xor ( n44645 , n44016 , n44338 );
and ( n44646 , n30144 , n44442 );
and ( n44647 , n44645 , n44646 );
xor ( n44648 , n44645 , n44646 );
xor ( n44649 , n44020 , n44336 );
and ( n44650 , n30149 , n44442 );
and ( n44651 , n44649 , n44650 );
xor ( n44652 , n44649 , n44650 );
xor ( n44653 , n44024 , n44334 );
and ( n44654 , n30154 , n44442 );
and ( n44655 , n44653 , n44654 );
xor ( n44656 , n44653 , n44654 );
xor ( n44657 , n44028 , n44332 );
and ( n44658 , n30159 , n44442 );
and ( n44659 , n44657 , n44658 );
xor ( n44660 , n44657 , n44658 );
xor ( n44661 , n44032 , n44330 );
and ( n44662 , n30164 , n44442 );
and ( n44663 , n44661 , n44662 );
xor ( n44664 , n44661 , n44662 );
xor ( n44665 , n44036 , n44328 );
and ( n44666 , n30169 , n44442 );
and ( n44667 , n44665 , n44666 );
xor ( n44668 , n44665 , n44666 );
xor ( n44669 , n44040 , n44326 );
and ( n44670 , n30174 , n44442 );
and ( n44671 , n44669 , n44670 );
xor ( n44672 , n44669 , n44670 );
xor ( n44673 , n44044 , n44324 );
and ( n44674 , n30179 , n44442 );
and ( n44675 , n44673 , n44674 );
xor ( n44676 , n44673 , n44674 );
xor ( n44677 , n44048 , n44322 );
and ( n44678 , n30184 , n44442 );
and ( n44679 , n44677 , n44678 );
xor ( n44680 , n44677 , n44678 );
xor ( n44681 , n44052 , n44320 );
and ( n44682 , n30189 , n44442 );
and ( n44683 , n44681 , n44682 );
xor ( n44684 , n44681 , n44682 );
xor ( n44685 , n44056 , n44318 );
and ( n44686 , n30194 , n44442 );
and ( n44687 , n44685 , n44686 );
xor ( n44688 , n44685 , n44686 );
xor ( n44689 , n44060 , n44316 );
and ( n44690 , n30199 , n44442 );
and ( n44691 , n44689 , n44690 );
xor ( n44692 , n44689 , n44690 );
xor ( n44693 , n44064 , n44314 );
and ( n44694 , n30204 , n44442 );
and ( n44695 , n44693 , n44694 );
xor ( n44696 , n44693 , n44694 );
xor ( n44697 , n44068 , n44312 );
and ( n44698 , n30209 , n44442 );
and ( n44699 , n44697 , n44698 );
xor ( n44700 , n44697 , n44698 );
xor ( n44701 , n44072 , n44310 );
and ( n44702 , n30214 , n44442 );
and ( n44703 , n44701 , n44702 );
xor ( n44704 , n44701 , n44702 );
xor ( n44705 , n44076 , n44308 );
and ( n44706 , n30219 , n44442 );
and ( n44707 , n44705 , n44706 );
xor ( n44708 , n44705 , n44706 );
xor ( n44709 , n44080 , n44306 );
and ( n44710 , n30224 , n44442 );
and ( n44711 , n44709 , n44710 );
xor ( n44712 , n44709 , n44710 );
xor ( n44713 , n44084 , n44304 );
and ( n44714 , n30229 , n44442 );
and ( n44715 , n44713 , n44714 );
xor ( n44716 , n44713 , n44714 );
xor ( n44717 , n44088 , n44302 );
and ( n44718 , n30234 , n44442 );
and ( n44719 , n44717 , n44718 );
xor ( n44720 , n44717 , n44718 );
xor ( n44721 , n44092 , n44300 );
and ( n44722 , n30239 , n44442 );
and ( n44723 , n44721 , n44722 );
xor ( n44724 , n44721 , n44722 );
xor ( n44725 , n44096 , n44298 );
and ( n44726 , n30244 , n44442 );
and ( n44727 , n44725 , n44726 );
xor ( n44728 , n44725 , n44726 );
xor ( n44729 , n44100 , n44296 );
and ( n44730 , n30249 , n44442 );
and ( n44731 , n44729 , n44730 );
xor ( n44732 , n44729 , n44730 );
xor ( n44733 , n44104 , n44294 );
and ( n44734 , n30254 , n44442 );
and ( n44735 , n44733 , n44734 );
xor ( n44736 , n44733 , n44734 );
xor ( n44737 , n44108 , n44292 );
and ( n44738 , n30259 , n44442 );
and ( n44739 , n44737 , n44738 );
xor ( n44740 , n44737 , n44738 );
xor ( n44741 , n44112 , n44290 );
and ( n44742 , n30264 , n44442 );
and ( n44743 , n44741 , n44742 );
xor ( n44744 , n44741 , n44742 );
xor ( n44745 , n44116 , n44288 );
and ( n44746 , n30269 , n44442 );
and ( n44747 , n44745 , n44746 );
xor ( n44748 , n44745 , n44746 );
xor ( n44749 , n44120 , n44286 );
and ( n44750 , n30274 , n44442 );
and ( n44751 , n44749 , n44750 );
xor ( n44752 , n44749 , n44750 );
xor ( n44753 , n44124 , n44284 );
and ( n44754 , n30279 , n44442 );
and ( n44755 , n44753 , n44754 );
xor ( n44756 , n44753 , n44754 );
xor ( n44757 , n44128 , n44282 );
and ( n44758 , n30284 , n44442 );
and ( n44759 , n44757 , n44758 );
xor ( n44760 , n44757 , n44758 );
xor ( n44761 , n44132 , n44280 );
and ( n44762 , n30289 , n44442 );
and ( n44763 , n44761 , n44762 );
xor ( n44764 , n44761 , n44762 );
xor ( n44765 , n44136 , n44278 );
and ( n44766 , n30294 , n44442 );
and ( n44767 , n44765 , n44766 );
xor ( n44768 , n44765 , n44766 );
xor ( n44769 , n44140 , n44276 );
and ( n44770 , n30299 , n44442 );
and ( n44771 , n44769 , n44770 );
xor ( n44772 , n44769 , n44770 );
xor ( n44773 , n44144 , n44274 );
and ( n44774 , n30304 , n44442 );
and ( n44775 , n44773 , n44774 );
xor ( n44776 , n44773 , n44774 );
xor ( n44777 , n44148 , n44272 );
and ( n44778 , n30309 , n44442 );
and ( n44779 , n44777 , n44778 );
xor ( n44780 , n44777 , n44778 );
xor ( n44781 , n44152 , n44270 );
and ( n44782 , n30314 , n44442 );
and ( n44783 , n44781 , n44782 );
xor ( n44784 , n44781 , n44782 );
xor ( n44785 , n44156 , n44268 );
and ( n44786 , n30319 , n44442 );
and ( n44787 , n44785 , n44786 );
xor ( n44788 , n44785 , n44786 );
xor ( n44789 , n44160 , n44266 );
and ( n44790 , n30324 , n44442 );
and ( n44791 , n44789 , n44790 );
xor ( n44792 , n44789 , n44790 );
xor ( n44793 , n44164 , n44264 );
and ( n44794 , n30329 , n44442 );
and ( n44795 , n44793 , n44794 );
xor ( n44796 , n44793 , n44794 );
xor ( n44797 , n44168 , n44262 );
and ( n44798 , n30334 , n44442 );
and ( n44799 , n44797 , n44798 );
xor ( n44800 , n44797 , n44798 );
xor ( n44801 , n44172 , n44260 );
and ( n44802 , n30339 , n44442 );
and ( n44803 , n44801 , n44802 );
xor ( n44804 , n44801 , n44802 );
xor ( n44805 , n44176 , n44258 );
and ( n44806 , n30344 , n44442 );
and ( n44807 , n44805 , n44806 );
xor ( n44808 , n44805 , n44806 );
xor ( n44809 , n44180 , n44256 );
and ( n44810 , n30349 , n44442 );
and ( n44811 , n44809 , n44810 );
xor ( n44812 , n44809 , n44810 );
xor ( n44813 , n44184 , n44254 );
and ( n44814 , n30354 , n44442 );
and ( n44815 , n44813 , n44814 );
xor ( n44816 , n44813 , n44814 );
xor ( n44817 , n44188 , n44252 );
and ( n44818 , n30359 , n44442 );
and ( n44819 , n44817 , n44818 );
xor ( n44820 , n44817 , n44818 );
xor ( n44821 , n44192 , n44250 );
and ( n44822 , n30364 , n44442 );
and ( n44823 , n44821 , n44822 );
xor ( n44824 , n44821 , n44822 );
xor ( n44825 , n44196 , n44248 );
and ( n44826 , n30369 , n44442 );
and ( n44827 , n44825 , n44826 );
xor ( n44828 , n44825 , n44826 );
xor ( n44829 , n44200 , n44246 );
and ( n44830 , n30374 , n44442 );
and ( n44831 , n44829 , n44830 );
xor ( n44832 , n44829 , n44830 );
xor ( n44833 , n44204 , n44244 );
and ( n44834 , n30379 , n44442 );
and ( n44835 , n44833 , n44834 );
xor ( n44836 , n44833 , n44834 );
xor ( n44837 , n44208 , n44242 );
and ( n44838 , n30384 , n44442 );
and ( n44839 , n44837 , n44838 );
xor ( n44840 , n44837 , n44838 );
xor ( n44841 , n44212 , n44240 );
and ( n44842 , n30389 , n44442 );
and ( n44843 , n44841 , n44842 );
xor ( n44844 , n44841 , n44842 );
xor ( n44845 , n44216 , n44238 );
and ( n44846 , n30394 , n44442 );
and ( n44847 , n44845 , n44846 );
xor ( n44848 , n44845 , n44846 );
xor ( n44849 , n44220 , n44236 );
and ( n44850 , n30399 , n44442 );
and ( n44851 , n44849 , n44850 );
xor ( n44852 , n44849 , n44850 );
xor ( n44853 , n44224 , n44234 );
and ( n44854 , n30404 , n44442 );
and ( n44855 , n44853 , n44854 );
xor ( n44856 , n44853 , n44854 );
xor ( n44857 , n44228 , n44232 );
and ( n44858 , n30409 , n44442 );
and ( n44859 , n44857 , n44858 );
buf ( n44860 , n44859 );
and ( n44861 , n44856 , n44860 );
or ( n44862 , n44855 , n44861 );
and ( n44863 , n44852 , n44862 );
or ( n44864 , n44851 , n44863 );
and ( n44865 , n44848 , n44864 );
or ( n44866 , n44847 , n44865 );
and ( n44867 , n44844 , n44866 );
or ( n44868 , n44843 , n44867 );
and ( n44869 , n44840 , n44868 );
or ( n44870 , n44839 , n44869 );
and ( n44871 , n44836 , n44870 );
or ( n44872 , n44835 , n44871 );
and ( n44873 , n44832 , n44872 );
or ( n44874 , n44831 , n44873 );
and ( n44875 , n44828 , n44874 );
or ( n44876 , n44827 , n44875 );
and ( n44877 , n44824 , n44876 );
or ( n44878 , n44823 , n44877 );
and ( n44879 , n44820 , n44878 );
or ( n44880 , n44819 , n44879 );
and ( n44881 , n44816 , n44880 );
or ( n44882 , n44815 , n44881 );
and ( n44883 , n44812 , n44882 );
or ( n44884 , n44811 , n44883 );
and ( n44885 , n44808 , n44884 );
or ( n44886 , n44807 , n44885 );
and ( n44887 , n44804 , n44886 );
or ( n44888 , n44803 , n44887 );
and ( n44889 , n44800 , n44888 );
or ( n44890 , n44799 , n44889 );
and ( n44891 , n44796 , n44890 );
or ( n44892 , n44795 , n44891 );
and ( n44893 , n44792 , n44892 );
or ( n44894 , n44791 , n44893 );
and ( n44895 , n44788 , n44894 );
or ( n44896 , n44787 , n44895 );
and ( n44897 , n44784 , n44896 );
or ( n44898 , n44783 , n44897 );
and ( n44899 , n44780 , n44898 );
or ( n44900 , n44779 , n44899 );
and ( n44901 , n44776 , n44900 );
or ( n44902 , n44775 , n44901 );
and ( n44903 , n44772 , n44902 );
or ( n44904 , n44771 , n44903 );
and ( n44905 , n44768 , n44904 );
or ( n44906 , n44767 , n44905 );
and ( n44907 , n44764 , n44906 );
or ( n44908 , n44763 , n44907 );
and ( n44909 , n44760 , n44908 );
or ( n44910 , n44759 , n44909 );
and ( n44911 , n44756 , n44910 );
or ( n44912 , n44755 , n44911 );
and ( n44913 , n44752 , n44912 );
or ( n44914 , n44751 , n44913 );
and ( n44915 , n44748 , n44914 );
or ( n44916 , n44747 , n44915 );
and ( n44917 , n44744 , n44916 );
or ( n44918 , n44743 , n44917 );
and ( n44919 , n44740 , n44918 );
or ( n44920 , n44739 , n44919 );
and ( n44921 , n44736 , n44920 );
or ( n44922 , n44735 , n44921 );
and ( n44923 , n44732 , n44922 );
or ( n44924 , n44731 , n44923 );
and ( n44925 , n44728 , n44924 );
or ( n44926 , n44727 , n44925 );
and ( n44927 , n44724 , n44926 );
or ( n44928 , n44723 , n44927 );
and ( n44929 , n44720 , n44928 );
or ( n44930 , n44719 , n44929 );
and ( n44931 , n44716 , n44930 );
or ( n44932 , n44715 , n44931 );
and ( n44933 , n44712 , n44932 );
or ( n44934 , n44711 , n44933 );
and ( n44935 , n44708 , n44934 );
or ( n44936 , n44707 , n44935 );
and ( n44937 , n44704 , n44936 );
or ( n44938 , n44703 , n44937 );
and ( n44939 , n44700 , n44938 );
or ( n44940 , n44699 , n44939 );
and ( n44941 , n44696 , n44940 );
or ( n44942 , n44695 , n44941 );
and ( n44943 , n44692 , n44942 );
or ( n44944 , n44691 , n44943 );
and ( n44945 , n44688 , n44944 );
or ( n44946 , n44687 , n44945 );
and ( n44947 , n44684 , n44946 );
or ( n44948 , n44683 , n44947 );
and ( n44949 , n44680 , n44948 );
or ( n44950 , n44679 , n44949 );
and ( n44951 , n44676 , n44950 );
or ( n44952 , n44675 , n44951 );
and ( n44953 , n44672 , n44952 );
or ( n44954 , n44671 , n44953 );
and ( n44955 , n44668 , n44954 );
or ( n44956 , n44667 , n44955 );
and ( n44957 , n44664 , n44956 );
or ( n44958 , n44663 , n44957 );
and ( n44959 , n44660 , n44958 );
or ( n44960 , n44659 , n44959 );
and ( n44961 , n44656 , n44960 );
or ( n44962 , n44655 , n44961 );
and ( n44963 , n44652 , n44962 );
or ( n44964 , n44651 , n44963 );
and ( n44965 , n44648 , n44964 );
or ( n44966 , n44647 , n44965 );
and ( n44967 , n44644 , n44966 );
or ( n44968 , n44643 , n44967 );
and ( n44969 , n44640 , n44968 );
or ( n44970 , n44639 , n44969 );
and ( n44971 , n44636 , n44970 );
or ( n44972 , n44635 , n44971 );
and ( n44973 , n44632 , n44972 );
or ( n44974 , n44631 , n44973 );
and ( n44975 , n44628 , n44974 );
or ( n44976 , n44627 , n44975 );
and ( n44977 , n44624 , n44976 );
or ( n44978 , n44623 , n44977 );
and ( n44979 , n44620 , n44978 );
or ( n44980 , n44619 , n44979 );
and ( n44981 , n44616 , n44980 );
or ( n44982 , n44615 , n44981 );
and ( n44983 , n44612 , n44982 );
or ( n44984 , n44611 , n44983 );
and ( n44985 , n44608 , n44984 );
or ( n44986 , n44607 , n44985 );
and ( n44987 , n44604 , n44986 );
or ( n44988 , n44603 , n44987 );
and ( n44989 , n44600 , n44988 );
or ( n44990 , n44599 , n44989 );
and ( n44991 , n44596 , n44990 );
or ( n44992 , n44595 , n44991 );
and ( n44993 , n44592 , n44992 );
or ( n44994 , n44591 , n44993 );
and ( n44995 , n44588 , n44994 );
or ( n44996 , n44587 , n44995 );
and ( n44997 , n44584 , n44996 );
or ( n44998 , n44583 , n44997 );
and ( n44999 , n44580 , n44998 );
or ( n45000 , n44579 , n44999 );
and ( n45001 , n44576 , n45000 );
or ( n45002 , n44575 , n45001 );
and ( n45003 , n44572 , n45002 );
or ( n45004 , n44571 , n45003 );
and ( n45005 , n44568 , n45004 );
or ( n45006 , n44567 , n45005 );
and ( n45007 , n44564 , n45006 );
or ( n45008 , n44563 , n45007 );
and ( n45009 , n44560 , n45008 );
or ( n45010 , n44559 , n45009 );
and ( n45011 , n44556 , n45010 );
or ( n45012 , n44555 , n45011 );
and ( n45013 , n44552 , n45012 );
or ( n45014 , n44551 , n45013 );
and ( n45015 , n44548 , n45014 );
or ( n45016 , n44547 , n45015 );
and ( n45017 , n44544 , n45016 );
or ( n45018 , n44543 , n45017 );
and ( n45019 , n44540 , n45018 );
or ( n45020 , n44539 , n45019 );
and ( n45021 , n44536 , n45020 );
or ( n45022 , n44535 , n45021 );
and ( n45023 , n44532 , n45022 );
or ( n45024 , n44531 , n45023 );
and ( n45025 , n44528 , n45024 );
or ( n45026 , n44527 , n45025 );
and ( n45027 , n44524 , n45026 );
or ( n45028 , n44523 , n45027 );
and ( n45029 , n44520 , n45028 );
or ( n45030 , n44519 , n45029 );
and ( n45031 , n44516 , n45030 );
or ( n45032 , n44515 , n45031 );
and ( n45033 , n44512 , n45032 );
or ( n45034 , n44511 , n45033 );
and ( n45035 , n44508 , n45034 );
or ( n45036 , n44507 , n45035 );
and ( n45037 , n44504 , n45036 );
or ( n45038 , n44503 , n45037 );
and ( n45039 , n44500 , n45038 );
or ( n45040 , n44499 , n45039 );
and ( n45041 , n44496 , n45040 );
or ( n45042 , n44495 , n45041 );
and ( n45043 , n44492 , n45042 );
or ( n45044 , n44491 , n45043 );
and ( n45045 , n44488 , n45044 );
or ( n45046 , n44487 , n45045 );
and ( n45047 , n44484 , n45046 );
or ( n45048 , n44483 , n45047 );
and ( n45049 , n44480 , n45048 );
or ( n45050 , n44479 , n45049 );
and ( n45051 , n44476 , n45050 );
or ( n45052 , n44475 , n45051 );
and ( n45053 , n44472 , n45052 );
or ( n45054 , n44471 , n45053 );
and ( n45055 , n44468 , n45054 );
or ( n45056 , n44467 , n45055 );
and ( n45057 , n44464 , n45056 );
or ( n45058 , n44463 , n45057 );
and ( n45059 , n44460 , n45058 );
or ( n45060 , n44459 , n45059 );
and ( n45061 , n44456 , n45060 );
or ( n45062 , n44455 , n45061 );
and ( n45063 , n44452 , n45062 );
or ( n45064 , n44451 , n45063 );
and ( n45065 , n44448 , n45064 );
or ( n45066 , n44447 , n45065 );
xor ( n45067 , n44444 , n45066 );
buf ( n45068 , n18060 );
and ( n45069 , n29894 , n45068 );
xor ( n45070 , n45067 , n45069 );
xor ( n45071 , n44448 , n45064 );
and ( n45072 , n29899 , n45068 );
and ( n45073 , n45071 , n45072 );
xor ( n45074 , n45071 , n45072 );
xor ( n45075 , n44452 , n45062 );
and ( n45076 , n29904 , n45068 );
and ( n45077 , n45075 , n45076 );
xor ( n45078 , n45075 , n45076 );
xor ( n45079 , n44456 , n45060 );
and ( n45080 , n29909 , n45068 );
and ( n45081 , n45079 , n45080 );
xor ( n45082 , n45079 , n45080 );
xor ( n45083 , n44460 , n45058 );
and ( n45084 , n29914 , n45068 );
and ( n45085 , n45083 , n45084 );
xor ( n45086 , n45083 , n45084 );
xor ( n45087 , n44464 , n45056 );
and ( n45088 , n29919 , n45068 );
and ( n45089 , n45087 , n45088 );
xor ( n45090 , n45087 , n45088 );
xor ( n45091 , n44468 , n45054 );
and ( n45092 , n29924 , n45068 );
and ( n45093 , n45091 , n45092 );
xor ( n45094 , n45091 , n45092 );
xor ( n45095 , n44472 , n45052 );
and ( n45096 , n29929 , n45068 );
and ( n45097 , n45095 , n45096 );
xor ( n45098 , n45095 , n45096 );
xor ( n45099 , n44476 , n45050 );
and ( n45100 , n29934 , n45068 );
and ( n45101 , n45099 , n45100 );
xor ( n45102 , n45099 , n45100 );
xor ( n45103 , n44480 , n45048 );
and ( n45104 , n29939 , n45068 );
and ( n45105 , n45103 , n45104 );
xor ( n45106 , n45103 , n45104 );
xor ( n45107 , n44484 , n45046 );
and ( n45108 , n29944 , n45068 );
and ( n45109 , n45107 , n45108 );
xor ( n45110 , n45107 , n45108 );
xor ( n45111 , n44488 , n45044 );
and ( n45112 , n29949 , n45068 );
and ( n45113 , n45111 , n45112 );
xor ( n45114 , n45111 , n45112 );
xor ( n45115 , n44492 , n45042 );
and ( n45116 , n29954 , n45068 );
and ( n45117 , n45115 , n45116 );
xor ( n45118 , n45115 , n45116 );
xor ( n45119 , n44496 , n45040 );
and ( n45120 , n29959 , n45068 );
and ( n45121 , n45119 , n45120 );
xor ( n45122 , n45119 , n45120 );
xor ( n45123 , n44500 , n45038 );
and ( n45124 , n29964 , n45068 );
and ( n45125 , n45123 , n45124 );
xor ( n45126 , n45123 , n45124 );
xor ( n45127 , n44504 , n45036 );
and ( n45128 , n29969 , n45068 );
and ( n45129 , n45127 , n45128 );
xor ( n45130 , n45127 , n45128 );
xor ( n45131 , n44508 , n45034 );
and ( n45132 , n29974 , n45068 );
and ( n45133 , n45131 , n45132 );
xor ( n45134 , n45131 , n45132 );
xor ( n45135 , n44512 , n45032 );
and ( n45136 , n29979 , n45068 );
and ( n45137 , n45135 , n45136 );
xor ( n45138 , n45135 , n45136 );
xor ( n45139 , n44516 , n45030 );
and ( n45140 , n29984 , n45068 );
and ( n45141 , n45139 , n45140 );
xor ( n45142 , n45139 , n45140 );
xor ( n45143 , n44520 , n45028 );
and ( n45144 , n29989 , n45068 );
and ( n45145 , n45143 , n45144 );
xor ( n45146 , n45143 , n45144 );
xor ( n45147 , n44524 , n45026 );
and ( n45148 , n29994 , n45068 );
and ( n45149 , n45147 , n45148 );
xor ( n45150 , n45147 , n45148 );
xor ( n45151 , n44528 , n45024 );
and ( n45152 , n29999 , n45068 );
and ( n45153 , n45151 , n45152 );
xor ( n45154 , n45151 , n45152 );
xor ( n45155 , n44532 , n45022 );
and ( n45156 , n30004 , n45068 );
and ( n45157 , n45155 , n45156 );
xor ( n45158 , n45155 , n45156 );
xor ( n45159 , n44536 , n45020 );
and ( n45160 , n30009 , n45068 );
and ( n45161 , n45159 , n45160 );
xor ( n45162 , n45159 , n45160 );
xor ( n45163 , n44540 , n45018 );
and ( n45164 , n30014 , n45068 );
and ( n45165 , n45163 , n45164 );
xor ( n45166 , n45163 , n45164 );
xor ( n45167 , n44544 , n45016 );
and ( n45168 , n30019 , n45068 );
and ( n45169 , n45167 , n45168 );
xor ( n45170 , n45167 , n45168 );
xor ( n45171 , n44548 , n45014 );
and ( n45172 , n30024 , n45068 );
and ( n45173 , n45171 , n45172 );
xor ( n45174 , n45171 , n45172 );
xor ( n45175 , n44552 , n45012 );
and ( n45176 , n30029 , n45068 );
and ( n45177 , n45175 , n45176 );
xor ( n45178 , n45175 , n45176 );
xor ( n45179 , n44556 , n45010 );
and ( n45180 , n30034 , n45068 );
and ( n45181 , n45179 , n45180 );
xor ( n45182 , n45179 , n45180 );
xor ( n45183 , n44560 , n45008 );
and ( n45184 , n30039 , n45068 );
and ( n45185 , n45183 , n45184 );
xor ( n45186 , n45183 , n45184 );
xor ( n45187 , n44564 , n45006 );
and ( n45188 , n30044 , n45068 );
and ( n45189 , n45187 , n45188 );
xor ( n45190 , n45187 , n45188 );
xor ( n45191 , n44568 , n45004 );
and ( n45192 , n30049 , n45068 );
and ( n45193 , n45191 , n45192 );
xor ( n45194 , n45191 , n45192 );
xor ( n45195 , n44572 , n45002 );
and ( n45196 , n30054 , n45068 );
and ( n45197 , n45195 , n45196 );
xor ( n45198 , n45195 , n45196 );
xor ( n45199 , n44576 , n45000 );
and ( n45200 , n30059 , n45068 );
and ( n45201 , n45199 , n45200 );
xor ( n45202 , n45199 , n45200 );
xor ( n45203 , n44580 , n44998 );
and ( n45204 , n30064 , n45068 );
and ( n45205 , n45203 , n45204 );
xor ( n45206 , n45203 , n45204 );
xor ( n45207 , n44584 , n44996 );
and ( n45208 , n30069 , n45068 );
and ( n45209 , n45207 , n45208 );
xor ( n45210 , n45207 , n45208 );
xor ( n45211 , n44588 , n44994 );
and ( n45212 , n30074 , n45068 );
and ( n45213 , n45211 , n45212 );
xor ( n45214 , n45211 , n45212 );
xor ( n45215 , n44592 , n44992 );
and ( n45216 , n30079 , n45068 );
and ( n45217 , n45215 , n45216 );
xor ( n45218 , n45215 , n45216 );
xor ( n45219 , n44596 , n44990 );
and ( n45220 , n30084 , n45068 );
and ( n45221 , n45219 , n45220 );
xor ( n45222 , n45219 , n45220 );
xor ( n45223 , n44600 , n44988 );
and ( n45224 , n30089 , n45068 );
and ( n45225 , n45223 , n45224 );
xor ( n45226 , n45223 , n45224 );
xor ( n45227 , n44604 , n44986 );
and ( n45228 , n30094 , n45068 );
and ( n45229 , n45227 , n45228 );
xor ( n45230 , n45227 , n45228 );
xor ( n45231 , n44608 , n44984 );
and ( n45232 , n30099 , n45068 );
and ( n45233 , n45231 , n45232 );
xor ( n45234 , n45231 , n45232 );
xor ( n45235 , n44612 , n44982 );
and ( n45236 , n30104 , n45068 );
and ( n45237 , n45235 , n45236 );
xor ( n45238 , n45235 , n45236 );
xor ( n45239 , n44616 , n44980 );
and ( n45240 , n30109 , n45068 );
and ( n45241 , n45239 , n45240 );
xor ( n45242 , n45239 , n45240 );
xor ( n45243 , n44620 , n44978 );
and ( n45244 , n30114 , n45068 );
and ( n45245 , n45243 , n45244 );
xor ( n45246 , n45243 , n45244 );
xor ( n45247 , n44624 , n44976 );
and ( n45248 , n30119 , n45068 );
and ( n45249 , n45247 , n45248 );
xor ( n45250 , n45247 , n45248 );
xor ( n45251 , n44628 , n44974 );
and ( n45252 , n30124 , n45068 );
and ( n45253 , n45251 , n45252 );
xor ( n45254 , n45251 , n45252 );
xor ( n45255 , n44632 , n44972 );
and ( n45256 , n30129 , n45068 );
and ( n45257 , n45255 , n45256 );
xor ( n45258 , n45255 , n45256 );
xor ( n45259 , n44636 , n44970 );
and ( n45260 , n30134 , n45068 );
and ( n45261 , n45259 , n45260 );
xor ( n45262 , n45259 , n45260 );
xor ( n45263 , n44640 , n44968 );
and ( n45264 , n30139 , n45068 );
and ( n45265 , n45263 , n45264 );
xor ( n45266 , n45263 , n45264 );
xor ( n45267 , n44644 , n44966 );
and ( n45268 , n30144 , n45068 );
and ( n45269 , n45267 , n45268 );
xor ( n45270 , n45267 , n45268 );
xor ( n45271 , n44648 , n44964 );
and ( n45272 , n30149 , n45068 );
and ( n45273 , n45271 , n45272 );
xor ( n45274 , n45271 , n45272 );
xor ( n45275 , n44652 , n44962 );
and ( n45276 , n30154 , n45068 );
and ( n45277 , n45275 , n45276 );
xor ( n45278 , n45275 , n45276 );
xor ( n45279 , n44656 , n44960 );
and ( n45280 , n30159 , n45068 );
and ( n45281 , n45279 , n45280 );
xor ( n45282 , n45279 , n45280 );
xor ( n45283 , n44660 , n44958 );
and ( n45284 , n30164 , n45068 );
and ( n45285 , n45283 , n45284 );
xor ( n45286 , n45283 , n45284 );
xor ( n45287 , n44664 , n44956 );
and ( n45288 , n30169 , n45068 );
and ( n45289 , n45287 , n45288 );
xor ( n45290 , n45287 , n45288 );
xor ( n45291 , n44668 , n44954 );
and ( n45292 , n30174 , n45068 );
and ( n45293 , n45291 , n45292 );
xor ( n45294 , n45291 , n45292 );
xor ( n45295 , n44672 , n44952 );
and ( n45296 , n30179 , n45068 );
and ( n45297 , n45295 , n45296 );
xor ( n45298 , n45295 , n45296 );
xor ( n45299 , n44676 , n44950 );
and ( n45300 , n30184 , n45068 );
and ( n45301 , n45299 , n45300 );
xor ( n45302 , n45299 , n45300 );
xor ( n45303 , n44680 , n44948 );
and ( n45304 , n30189 , n45068 );
and ( n45305 , n45303 , n45304 );
xor ( n45306 , n45303 , n45304 );
xor ( n45307 , n44684 , n44946 );
and ( n45308 , n30194 , n45068 );
and ( n45309 , n45307 , n45308 );
xor ( n45310 , n45307 , n45308 );
xor ( n45311 , n44688 , n44944 );
and ( n45312 , n30199 , n45068 );
and ( n45313 , n45311 , n45312 );
xor ( n45314 , n45311 , n45312 );
xor ( n45315 , n44692 , n44942 );
and ( n45316 , n30204 , n45068 );
and ( n45317 , n45315 , n45316 );
xor ( n45318 , n45315 , n45316 );
xor ( n45319 , n44696 , n44940 );
and ( n45320 , n30209 , n45068 );
and ( n45321 , n45319 , n45320 );
xor ( n45322 , n45319 , n45320 );
xor ( n45323 , n44700 , n44938 );
and ( n45324 , n30214 , n45068 );
and ( n45325 , n45323 , n45324 );
xor ( n45326 , n45323 , n45324 );
xor ( n45327 , n44704 , n44936 );
and ( n45328 , n30219 , n45068 );
and ( n45329 , n45327 , n45328 );
xor ( n45330 , n45327 , n45328 );
xor ( n45331 , n44708 , n44934 );
and ( n45332 , n30224 , n45068 );
and ( n45333 , n45331 , n45332 );
xor ( n45334 , n45331 , n45332 );
xor ( n45335 , n44712 , n44932 );
and ( n45336 , n30229 , n45068 );
and ( n45337 , n45335 , n45336 );
xor ( n45338 , n45335 , n45336 );
xor ( n45339 , n44716 , n44930 );
and ( n45340 , n30234 , n45068 );
and ( n45341 , n45339 , n45340 );
xor ( n45342 , n45339 , n45340 );
xor ( n45343 , n44720 , n44928 );
and ( n45344 , n30239 , n45068 );
and ( n45345 , n45343 , n45344 );
xor ( n45346 , n45343 , n45344 );
xor ( n45347 , n44724 , n44926 );
and ( n45348 , n30244 , n45068 );
and ( n45349 , n45347 , n45348 );
xor ( n45350 , n45347 , n45348 );
xor ( n45351 , n44728 , n44924 );
and ( n45352 , n30249 , n45068 );
and ( n45353 , n45351 , n45352 );
xor ( n45354 , n45351 , n45352 );
xor ( n45355 , n44732 , n44922 );
and ( n45356 , n30254 , n45068 );
and ( n45357 , n45355 , n45356 );
xor ( n45358 , n45355 , n45356 );
xor ( n45359 , n44736 , n44920 );
and ( n45360 , n30259 , n45068 );
and ( n45361 , n45359 , n45360 );
xor ( n45362 , n45359 , n45360 );
xor ( n45363 , n44740 , n44918 );
and ( n45364 , n30264 , n45068 );
and ( n45365 , n45363 , n45364 );
xor ( n45366 , n45363 , n45364 );
xor ( n45367 , n44744 , n44916 );
and ( n45368 , n30269 , n45068 );
and ( n45369 , n45367 , n45368 );
xor ( n45370 , n45367 , n45368 );
xor ( n45371 , n44748 , n44914 );
and ( n45372 , n30274 , n45068 );
and ( n45373 , n45371 , n45372 );
xor ( n45374 , n45371 , n45372 );
xor ( n45375 , n44752 , n44912 );
and ( n45376 , n30279 , n45068 );
and ( n45377 , n45375 , n45376 );
xor ( n45378 , n45375 , n45376 );
xor ( n45379 , n44756 , n44910 );
and ( n45380 , n30284 , n45068 );
and ( n45381 , n45379 , n45380 );
xor ( n45382 , n45379 , n45380 );
xor ( n45383 , n44760 , n44908 );
and ( n45384 , n30289 , n45068 );
and ( n45385 , n45383 , n45384 );
xor ( n45386 , n45383 , n45384 );
xor ( n45387 , n44764 , n44906 );
and ( n45388 , n30294 , n45068 );
and ( n45389 , n45387 , n45388 );
xor ( n45390 , n45387 , n45388 );
xor ( n45391 , n44768 , n44904 );
and ( n45392 , n30299 , n45068 );
and ( n45393 , n45391 , n45392 );
xor ( n45394 , n45391 , n45392 );
xor ( n45395 , n44772 , n44902 );
and ( n45396 , n30304 , n45068 );
and ( n45397 , n45395 , n45396 );
xor ( n45398 , n45395 , n45396 );
xor ( n45399 , n44776 , n44900 );
and ( n45400 , n30309 , n45068 );
and ( n45401 , n45399 , n45400 );
xor ( n45402 , n45399 , n45400 );
xor ( n45403 , n44780 , n44898 );
and ( n45404 , n30314 , n45068 );
and ( n45405 , n45403 , n45404 );
xor ( n45406 , n45403 , n45404 );
xor ( n45407 , n44784 , n44896 );
and ( n45408 , n30319 , n45068 );
and ( n45409 , n45407 , n45408 );
xor ( n45410 , n45407 , n45408 );
xor ( n45411 , n44788 , n44894 );
and ( n45412 , n30324 , n45068 );
and ( n45413 , n45411 , n45412 );
xor ( n45414 , n45411 , n45412 );
xor ( n45415 , n44792 , n44892 );
and ( n45416 , n30329 , n45068 );
and ( n45417 , n45415 , n45416 );
xor ( n45418 , n45415 , n45416 );
xor ( n45419 , n44796 , n44890 );
and ( n45420 , n30334 , n45068 );
and ( n45421 , n45419 , n45420 );
xor ( n45422 , n45419 , n45420 );
xor ( n45423 , n44800 , n44888 );
and ( n45424 , n30339 , n45068 );
and ( n45425 , n45423 , n45424 );
xor ( n45426 , n45423 , n45424 );
xor ( n45427 , n44804 , n44886 );
and ( n45428 , n30344 , n45068 );
and ( n45429 , n45427 , n45428 );
xor ( n45430 , n45427 , n45428 );
xor ( n45431 , n44808 , n44884 );
and ( n45432 , n30349 , n45068 );
and ( n45433 , n45431 , n45432 );
xor ( n45434 , n45431 , n45432 );
xor ( n45435 , n44812 , n44882 );
and ( n45436 , n30354 , n45068 );
and ( n45437 , n45435 , n45436 );
xor ( n45438 , n45435 , n45436 );
xor ( n45439 , n44816 , n44880 );
and ( n45440 , n30359 , n45068 );
and ( n45441 , n45439 , n45440 );
xor ( n45442 , n45439 , n45440 );
xor ( n45443 , n44820 , n44878 );
and ( n45444 , n30364 , n45068 );
and ( n45445 , n45443 , n45444 );
xor ( n45446 , n45443 , n45444 );
xor ( n45447 , n44824 , n44876 );
and ( n45448 , n30369 , n45068 );
and ( n45449 , n45447 , n45448 );
xor ( n45450 , n45447 , n45448 );
xor ( n45451 , n44828 , n44874 );
and ( n45452 , n30374 , n45068 );
and ( n45453 , n45451 , n45452 );
xor ( n45454 , n45451 , n45452 );
xor ( n45455 , n44832 , n44872 );
and ( n45456 , n30379 , n45068 );
and ( n45457 , n45455 , n45456 );
xor ( n45458 , n45455 , n45456 );
xor ( n45459 , n44836 , n44870 );
and ( n45460 , n30384 , n45068 );
and ( n45461 , n45459 , n45460 );
xor ( n45462 , n45459 , n45460 );
xor ( n45463 , n44840 , n44868 );
and ( n45464 , n30389 , n45068 );
and ( n45465 , n45463 , n45464 );
xor ( n45466 , n45463 , n45464 );
xor ( n45467 , n44844 , n44866 );
and ( n45468 , n30394 , n45068 );
and ( n45469 , n45467 , n45468 );
xor ( n45470 , n45467 , n45468 );
xor ( n45471 , n44848 , n44864 );
and ( n45472 , n30399 , n45068 );
and ( n45473 , n45471 , n45472 );
xor ( n45474 , n45471 , n45472 );
xor ( n45475 , n44852 , n44862 );
and ( n45476 , n30404 , n45068 );
and ( n45477 , n45475 , n45476 );
xor ( n45478 , n45475 , n45476 );
xor ( n45479 , n44856 , n44860 );
and ( n45480 , n30409 , n45068 );
and ( n45481 , n45479 , n45480 );
buf ( n45482 , n45481 );
and ( n45483 , n45478 , n45482 );
or ( n45484 , n45477 , n45483 );
and ( n45485 , n45474 , n45484 );
or ( n45486 , n45473 , n45485 );
and ( n45487 , n45470 , n45486 );
or ( n45488 , n45469 , n45487 );
and ( n45489 , n45466 , n45488 );
or ( n45490 , n45465 , n45489 );
and ( n45491 , n45462 , n45490 );
or ( n45492 , n45461 , n45491 );
and ( n45493 , n45458 , n45492 );
or ( n45494 , n45457 , n45493 );
and ( n45495 , n45454 , n45494 );
or ( n45496 , n45453 , n45495 );
and ( n45497 , n45450 , n45496 );
or ( n45498 , n45449 , n45497 );
and ( n45499 , n45446 , n45498 );
or ( n45500 , n45445 , n45499 );
and ( n45501 , n45442 , n45500 );
or ( n45502 , n45441 , n45501 );
and ( n45503 , n45438 , n45502 );
or ( n45504 , n45437 , n45503 );
and ( n45505 , n45434 , n45504 );
or ( n45506 , n45433 , n45505 );
and ( n45507 , n45430 , n45506 );
or ( n45508 , n45429 , n45507 );
and ( n45509 , n45426 , n45508 );
or ( n45510 , n45425 , n45509 );
and ( n45511 , n45422 , n45510 );
or ( n45512 , n45421 , n45511 );
and ( n45513 , n45418 , n45512 );
or ( n45514 , n45417 , n45513 );
and ( n45515 , n45414 , n45514 );
or ( n45516 , n45413 , n45515 );
and ( n45517 , n45410 , n45516 );
or ( n45518 , n45409 , n45517 );
and ( n45519 , n45406 , n45518 );
or ( n45520 , n45405 , n45519 );
and ( n45521 , n45402 , n45520 );
or ( n45522 , n45401 , n45521 );
and ( n45523 , n45398 , n45522 );
or ( n45524 , n45397 , n45523 );
and ( n45525 , n45394 , n45524 );
or ( n45526 , n45393 , n45525 );
and ( n45527 , n45390 , n45526 );
or ( n45528 , n45389 , n45527 );
and ( n45529 , n45386 , n45528 );
or ( n45530 , n45385 , n45529 );
and ( n45531 , n45382 , n45530 );
or ( n45532 , n45381 , n45531 );
and ( n45533 , n45378 , n45532 );
or ( n45534 , n45377 , n45533 );
and ( n45535 , n45374 , n45534 );
or ( n45536 , n45373 , n45535 );
and ( n45537 , n45370 , n45536 );
or ( n45538 , n45369 , n45537 );
and ( n45539 , n45366 , n45538 );
or ( n45540 , n45365 , n45539 );
and ( n45541 , n45362 , n45540 );
or ( n45542 , n45361 , n45541 );
and ( n45543 , n45358 , n45542 );
or ( n45544 , n45357 , n45543 );
and ( n45545 , n45354 , n45544 );
or ( n45546 , n45353 , n45545 );
and ( n45547 , n45350 , n45546 );
or ( n45548 , n45349 , n45547 );
and ( n45549 , n45346 , n45548 );
or ( n45550 , n45345 , n45549 );
and ( n45551 , n45342 , n45550 );
or ( n45552 , n45341 , n45551 );
and ( n45553 , n45338 , n45552 );
or ( n45554 , n45337 , n45553 );
and ( n45555 , n45334 , n45554 );
or ( n45556 , n45333 , n45555 );
and ( n45557 , n45330 , n45556 );
or ( n45558 , n45329 , n45557 );
and ( n45559 , n45326 , n45558 );
or ( n45560 , n45325 , n45559 );
and ( n45561 , n45322 , n45560 );
or ( n45562 , n45321 , n45561 );
and ( n45563 , n45318 , n45562 );
or ( n45564 , n45317 , n45563 );
and ( n45565 , n45314 , n45564 );
or ( n45566 , n45313 , n45565 );
and ( n45567 , n45310 , n45566 );
or ( n45568 , n45309 , n45567 );
and ( n45569 , n45306 , n45568 );
or ( n45570 , n45305 , n45569 );
and ( n45571 , n45302 , n45570 );
or ( n45572 , n45301 , n45571 );
and ( n45573 , n45298 , n45572 );
or ( n45574 , n45297 , n45573 );
and ( n45575 , n45294 , n45574 );
or ( n45576 , n45293 , n45575 );
and ( n45577 , n45290 , n45576 );
or ( n45578 , n45289 , n45577 );
and ( n45579 , n45286 , n45578 );
or ( n45580 , n45285 , n45579 );
and ( n45581 , n45282 , n45580 );
or ( n45582 , n45281 , n45581 );
and ( n45583 , n45278 , n45582 );
or ( n45584 , n45277 , n45583 );
and ( n45585 , n45274 , n45584 );
or ( n45586 , n45273 , n45585 );
and ( n45587 , n45270 , n45586 );
or ( n45588 , n45269 , n45587 );
and ( n45589 , n45266 , n45588 );
or ( n45590 , n45265 , n45589 );
and ( n45591 , n45262 , n45590 );
or ( n45592 , n45261 , n45591 );
and ( n45593 , n45258 , n45592 );
or ( n45594 , n45257 , n45593 );
and ( n45595 , n45254 , n45594 );
or ( n45596 , n45253 , n45595 );
and ( n45597 , n45250 , n45596 );
or ( n45598 , n45249 , n45597 );
and ( n45599 , n45246 , n45598 );
or ( n45600 , n45245 , n45599 );
and ( n45601 , n45242 , n45600 );
or ( n45602 , n45241 , n45601 );
and ( n45603 , n45238 , n45602 );
or ( n45604 , n45237 , n45603 );
and ( n45605 , n45234 , n45604 );
or ( n45606 , n45233 , n45605 );
and ( n45607 , n45230 , n45606 );
or ( n45608 , n45229 , n45607 );
and ( n45609 , n45226 , n45608 );
or ( n45610 , n45225 , n45609 );
and ( n45611 , n45222 , n45610 );
or ( n45612 , n45221 , n45611 );
and ( n45613 , n45218 , n45612 );
or ( n45614 , n45217 , n45613 );
and ( n45615 , n45214 , n45614 );
or ( n45616 , n45213 , n45615 );
and ( n45617 , n45210 , n45616 );
or ( n45618 , n45209 , n45617 );
and ( n45619 , n45206 , n45618 );
or ( n45620 , n45205 , n45619 );
and ( n45621 , n45202 , n45620 );
or ( n45622 , n45201 , n45621 );
and ( n45623 , n45198 , n45622 );
or ( n45624 , n45197 , n45623 );
and ( n45625 , n45194 , n45624 );
or ( n45626 , n45193 , n45625 );
and ( n45627 , n45190 , n45626 );
or ( n45628 , n45189 , n45627 );
and ( n45629 , n45186 , n45628 );
or ( n45630 , n45185 , n45629 );
and ( n45631 , n45182 , n45630 );
or ( n45632 , n45181 , n45631 );
and ( n45633 , n45178 , n45632 );
or ( n45634 , n45177 , n45633 );
and ( n45635 , n45174 , n45634 );
or ( n45636 , n45173 , n45635 );
and ( n45637 , n45170 , n45636 );
or ( n45638 , n45169 , n45637 );
and ( n45639 , n45166 , n45638 );
or ( n45640 , n45165 , n45639 );
and ( n45641 , n45162 , n45640 );
or ( n45642 , n45161 , n45641 );
and ( n45643 , n45158 , n45642 );
or ( n45644 , n45157 , n45643 );
and ( n45645 , n45154 , n45644 );
or ( n45646 , n45153 , n45645 );
and ( n45647 , n45150 , n45646 );
or ( n45648 , n45149 , n45647 );
and ( n45649 , n45146 , n45648 );
or ( n45650 , n45145 , n45649 );
and ( n45651 , n45142 , n45650 );
or ( n45652 , n45141 , n45651 );
and ( n45653 , n45138 , n45652 );
or ( n45654 , n45137 , n45653 );
and ( n45655 , n45134 , n45654 );
or ( n45656 , n45133 , n45655 );
and ( n45657 , n45130 , n45656 );
or ( n45658 , n45129 , n45657 );
and ( n45659 , n45126 , n45658 );
or ( n45660 , n45125 , n45659 );
and ( n45661 , n45122 , n45660 );
or ( n45662 , n45121 , n45661 );
and ( n45663 , n45118 , n45662 );
or ( n45664 , n45117 , n45663 );
and ( n45665 , n45114 , n45664 );
or ( n45666 , n45113 , n45665 );
and ( n45667 , n45110 , n45666 );
or ( n45668 , n45109 , n45667 );
and ( n45669 , n45106 , n45668 );
or ( n45670 , n45105 , n45669 );
and ( n45671 , n45102 , n45670 );
or ( n45672 , n45101 , n45671 );
and ( n45673 , n45098 , n45672 );
or ( n45674 , n45097 , n45673 );
and ( n45675 , n45094 , n45674 );
or ( n45676 , n45093 , n45675 );
and ( n45677 , n45090 , n45676 );
or ( n45678 , n45089 , n45677 );
and ( n45679 , n45086 , n45678 );
or ( n45680 , n45085 , n45679 );
and ( n45681 , n45082 , n45680 );
or ( n45682 , n45081 , n45681 );
and ( n45683 , n45078 , n45682 );
or ( n45684 , n45077 , n45683 );
and ( n45685 , n45074 , n45684 );
or ( n45686 , n45073 , n45685 );
xor ( n45687 , n45070 , n45686 );
buf ( n45688 , n18058 );
and ( n45689 , n29899 , n45688 );
xor ( n45690 , n45687 , n45689 );
xor ( n45691 , n45074 , n45684 );
and ( n45692 , n29904 , n45688 );
and ( n45693 , n45691 , n45692 );
xor ( n45694 , n45691 , n45692 );
xor ( n45695 , n45078 , n45682 );
and ( n45696 , n29909 , n45688 );
and ( n45697 , n45695 , n45696 );
xor ( n45698 , n45695 , n45696 );
xor ( n45699 , n45082 , n45680 );
and ( n45700 , n29914 , n45688 );
and ( n45701 , n45699 , n45700 );
xor ( n45702 , n45699 , n45700 );
xor ( n45703 , n45086 , n45678 );
and ( n45704 , n29919 , n45688 );
and ( n45705 , n45703 , n45704 );
xor ( n45706 , n45703 , n45704 );
xor ( n45707 , n45090 , n45676 );
and ( n45708 , n29924 , n45688 );
and ( n45709 , n45707 , n45708 );
xor ( n45710 , n45707 , n45708 );
xor ( n45711 , n45094 , n45674 );
and ( n45712 , n29929 , n45688 );
and ( n45713 , n45711 , n45712 );
xor ( n45714 , n45711 , n45712 );
xor ( n45715 , n45098 , n45672 );
and ( n45716 , n29934 , n45688 );
and ( n45717 , n45715 , n45716 );
xor ( n45718 , n45715 , n45716 );
xor ( n45719 , n45102 , n45670 );
and ( n45720 , n29939 , n45688 );
and ( n45721 , n45719 , n45720 );
xor ( n45722 , n45719 , n45720 );
xor ( n45723 , n45106 , n45668 );
and ( n45724 , n29944 , n45688 );
and ( n45725 , n45723 , n45724 );
xor ( n45726 , n45723 , n45724 );
xor ( n45727 , n45110 , n45666 );
and ( n45728 , n29949 , n45688 );
and ( n45729 , n45727 , n45728 );
xor ( n45730 , n45727 , n45728 );
xor ( n45731 , n45114 , n45664 );
and ( n45732 , n29954 , n45688 );
and ( n45733 , n45731 , n45732 );
xor ( n45734 , n45731 , n45732 );
xor ( n45735 , n45118 , n45662 );
and ( n45736 , n29959 , n45688 );
and ( n45737 , n45735 , n45736 );
xor ( n45738 , n45735 , n45736 );
xor ( n45739 , n45122 , n45660 );
and ( n45740 , n29964 , n45688 );
and ( n45741 , n45739 , n45740 );
xor ( n45742 , n45739 , n45740 );
xor ( n45743 , n45126 , n45658 );
and ( n45744 , n29969 , n45688 );
and ( n45745 , n45743 , n45744 );
xor ( n45746 , n45743 , n45744 );
xor ( n45747 , n45130 , n45656 );
and ( n45748 , n29974 , n45688 );
and ( n45749 , n45747 , n45748 );
xor ( n45750 , n45747 , n45748 );
xor ( n45751 , n45134 , n45654 );
and ( n45752 , n29979 , n45688 );
and ( n45753 , n45751 , n45752 );
xor ( n45754 , n45751 , n45752 );
xor ( n45755 , n45138 , n45652 );
and ( n45756 , n29984 , n45688 );
and ( n45757 , n45755 , n45756 );
xor ( n45758 , n45755 , n45756 );
xor ( n45759 , n45142 , n45650 );
and ( n45760 , n29989 , n45688 );
and ( n45761 , n45759 , n45760 );
xor ( n45762 , n45759 , n45760 );
xor ( n45763 , n45146 , n45648 );
and ( n45764 , n29994 , n45688 );
and ( n45765 , n45763 , n45764 );
xor ( n45766 , n45763 , n45764 );
xor ( n45767 , n45150 , n45646 );
and ( n45768 , n29999 , n45688 );
and ( n45769 , n45767 , n45768 );
xor ( n45770 , n45767 , n45768 );
xor ( n45771 , n45154 , n45644 );
and ( n45772 , n30004 , n45688 );
and ( n45773 , n45771 , n45772 );
xor ( n45774 , n45771 , n45772 );
xor ( n45775 , n45158 , n45642 );
and ( n45776 , n30009 , n45688 );
and ( n45777 , n45775 , n45776 );
xor ( n45778 , n45775 , n45776 );
xor ( n45779 , n45162 , n45640 );
and ( n45780 , n30014 , n45688 );
and ( n45781 , n45779 , n45780 );
xor ( n45782 , n45779 , n45780 );
xor ( n45783 , n45166 , n45638 );
and ( n45784 , n30019 , n45688 );
and ( n45785 , n45783 , n45784 );
xor ( n45786 , n45783 , n45784 );
xor ( n45787 , n45170 , n45636 );
and ( n45788 , n30024 , n45688 );
and ( n45789 , n45787 , n45788 );
xor ( n45790 , n45787 , n45788 );
xor ( n45791 , n45174 , n45634 );
and ( n45792 , n30029 , n45688 );
and ( n45793 , n45791 , n45792 );
xor ( n45794 , n45791 , n45792 );
xor ( n45795 , n45178 , n45632 );
and ( n45796 , n30034 , n45688 );
and ( n45797 , n45795 , n45796 );
xor ( n45798 , n45795 , n45796 );
xor ( n45799 , n45182 , n45630 );
and ( n45800 , n30039 , n45688 );
and ( n45801 , n45799 , n45800 );
xor ( n45802 , n45799 , n45800 );
xor ( n45803 , n45186 , n45628 );
and ( n45804 , n30044 , n45688 );
and ( n45805 , n45803 , n45804 );
xor ( n45806 , n45803 , n45804 );
xor ( n45807 , n45190 , n45626 );
and ( n45808 , n30049 , n45688 );
and ( n45809 , n45807 , n45808 );
xor ( n45810 , n45807 , n45808 );
xor ( n45811 , n45194 , n45624 );
and ( n45812 , n30054 , n45688 );
and ( n45813 , n45811 , n45812 );
xor ( n45814 , n45811 , n45812 );
xor ( n45815 , n45198 , n45622 );
and ( n45816 , n30059 , n45688 );
and ( n45817 , n45815 , n45816 );
xor ( n45818 , n45815 , n45816 );
xor ( n45819 , n45202 , n45620 );
and ( n45820 , n30064 , n45688 );
and ( n45821 , n45819 , n45820 );
xor ( n45822 , n45819 , n45820 );
xor ( n45823 , n45206 , n45618 );
and ( n45824 , n30069 , n45688 );
and ( n45825 , n45823 , n45824 );
xor ( n45826 , n45823 , n45824 );
xor ( n45827 , n45210 , n45616 );
and ( n45828 , n30074 , n45688 );
and ( n45829 , n45827 , n45828 );
xor ( n45830 , n45827 , n45828 );
xor ( n45831 , n45214 , n45614 );
and ( n45832 , n30079 , n45688 );
and ( n45833 , n45831 , n45832 );
xor ( n45834 , n45831 , n45832 );
xor ( n45835 , n45218 , n45612 );
and ( n45836 , n30084 , n45688 );
and ( n45837 , n45835 , n45836 );
xor ( n45838 , n45835 , n45836 );
xor ( n45839 , n45222 , n45610 );
and ( n45840 , n30089 , n45688 );
and ( n45841 , n45839 , n45840 );
xor ( n45842 , n45839 , n45840 );
xor ( n45843 , n45226 , n45608 );
and ( n45844 , n30094 , n45688 );
and ( n45845 , n45843 , n45844 );
xor ( n45846 , n45843 , n45844 );
xor ( n45847 , n45230 , n45606 );
and ( n45848 , n30099 , n45688 );
and ( n45849 , n45847 , n45848 );
xor ( n45850 , n45847 , n45848 );
xor ( n45851 , n45234 , n45604 );
and ( n45852 , n30104 , n45688 );
and ( n45853 , n45851 , n45852 );
xor ( n45854 , n45851 , n45852 );
xor ( n45855 , n45238 , n45602 );
and ( n45856 , n30109 , n45688 );
and ( n45857 , n45855 , n45856 );
xor ( n45858 , n45855 , n45856 );
xor ( n45859 , n45242 , n45600 );
and ( n45860 , n30114 , n45688 );
and ( n45861 , n45859 , n45860 );
xor ( n45862 , n45859 , n45860 );
xor ( n45863 , n45246 , n45598 );
and ( n45864 , n30119 , n45688 );
and ( n45865 , n45863 , n45864 );
xor ( n45866 , n45863 , n45864 );
xor ( n45867 , n45250 , n45596 );
and ( n45868 , n30124 , n45688 );
and ( n45869 , n45867 , n45868 );
xor ( n45870 , n45867 , n45868 );
xor ( n45871 , n45254 , n45594 );
and ( n45872 , n30129 , n45688 );
and ( n45873 , n45871 , n45872 );
xor ( n45874 , n45871 , n45872 );
xor ( n45875 , n45258 , n45592 );
and ( n45876 , n30134 , n45688 );
and ( n45877 , n45875 , n45876 );
xor ( n45878 , n45875 , n45876 );
xor ( n45879 , n45262 , n45590 );
and ( n45880 , n30139 , n45688 );
and ( n45881 , n45879 , n45880 );
xor ( n45882 , n45879 , n45880 );
xor ( n45883 , n45266 , n45588 );
and ( n45884 , n30144 , n45688 );
and ( n45885 , n45883 , n45884 );
xor ( n45886 , n45883 , n45884 );
xor ( n45887 , n45270 , n45586 );
and ( n45888 , n30149 , n45688 );
and ( n45889 , n45887 , n45888 );
xor ( n45890 , n45887 , n45888 );
xor ( n45891 , n45274 , n45584 );
and ( n45892 , n30154 , n45688 );
and ( n45893 , n45891 , n45892 );
xor ( n45894 , n45891 , n45892 );
xor ( n45895 , n45278 , n45582 );
and ( n45896 , n30159 , n45688 );
and ( n45897 , n45895 , n45896 );
xor ( n45898 , n45895 , n45896 );
xor ( n45899 , n45282 , n45580 );
and ( n45900 , n30164 , n45688 );
and ( n45901 , n45899 , n45900 );
xor ( n45902 , n45899 , n45900 );
xor ( n45903 , n45286 , n45578 );
and ( n45904 , n30169 , n45688 );
and ( n45905 , n45903 , n45904 );
xor ( n45906 , n45903 , n45904 );
xor ( n45907 , n45290 , n45576 );
and ( n45908 , n30174 , n45688 );
and ( n45909 , n45907 , n45908 );
xor ( n45910 , n45907 , n45908 );
xor ( n45911 , n45294 , n45574 );
and ( n45912 , n30179 , n45688 );
and ( n45913 , n45911 , n45912 );
xor ( n45914 , n45911 , n45912 );
xor ( n45915 , n45298 , n45572 );
and ( n45916 , n30184 , n45688 );
and ( n45917 , n45915 , n45916 );
xor ( n45918 , n45915 , n45916 );
xor ( n45919 , n45302 , n45570 );
and ( n45920 , n30189 , n45688 );
and ( n45921 , n45919 , n45920 );
xor ( n45922 , n45919 , n45920 );
xor ( n45923 , n45306 , n45568 );
and ( n45924 , n30194 , n45688 );
and ( n45925 , n45923 , n45924 );
xor ( n45926 , n45923 , n45924 );
xor ( n45927 , n45310 , n45566 );
and ( n45928 , n30199 , n45688 );
and ( n45929 , n45927 , n45928 );
xor ( n45930 , n45927 , n45928 );
xor ( n45931 , n45314 , n45564 );
and ( n45932 , n30204 , n45688 );
and ( n45933 , n45931 , n45932 );
xor ( n45934 , n45931 , n45932 );
xor ( n45935 , n45318 , n45562 );
and ( n45936 , n30209 , n45688 );
and ( n45937 , n45935 , n45936 );
xor ( n45938 , n45935 , n45936 );
xor ( n45939 , n45322 , n45560 );
and ( n45940 , n30214 , n45688 );
and ( n45941 , n45939 , n45940 );
xor ( n45942 , n45939 , n45940 );
xor ( n45943 , n45326 , n45558 );
and ( n45944 , n30219 , n45688 );
and ( n45945 , n45943 , n45944 );
xor ( n45946 , n45943 , n45944 );
xor ( n45947 , n45330 , n45556 );
and ( n45948 , n30224 , n45688 );
and ( n45949 , n45947 , n45948 );
xor ( n45950 , n45947 , n45948 );
xor ( n45951 , n45334 , n45554 );
and ( n45952 , n30229 , n45688 );
and ( n45953 , n45951 , n45952 );
xor ( n45954 , n45951 , n45952 );
xor ( n45955 , n45338 , n45552 );
and ( n45956 , n30234 , n45688 );
and ( n45957 , n45955 , n45956 );
xor ( n45958 , n45955 , n45956 );
xor ( n45959 , n45342 , n45550 );
and ( n45960 , n30239 , n45688 );
and ( n45961 , n45959 , n45960 );
xor ( n45962 , n45959 , n45960 );
xor ( n45963 , n45346 , n45548 );
and ( n45964 , n30244 , n45688 );
and ( n45965 , n45963 , n45964 );
xor ( n45966 , n45963 , n45964 );
xor ( n45967 , n45350 , n45546 );
and ( n45968 , n30249 , n45688 );
and ( n45969 , n45967 , n45968 );
xor ( n45970 , n45967 , n45968 );
xor ( n45971 , n45354 , n45544 );
and ( n45972 , n30254 , n45688 );
and ( n45973 , n45971 , n45972 );
xor ( n45974 , n45971 , n45972 );
xor ( n45975 , n45358 , n45542 );
and ( n45976 , n30259 , n45688 );
and ( n45977 , n45975 , n45976 );
xor ( n45978 , n45975 , n45976 );
xor ( n45979 , n45362 , n45540 );
and ( n45980 , n30264 , n45688 );
and ( n45981 , n45979 , n45980 );
xor ( n45982 , n45979 , n45980 );
xor ( n45983 , n45366 , n45538 );
and ( n45984 , n30269 , n45688 );
and ( n45985 , n45983 , n45984 );
xor ( n45986 , n45983 , n45984 );
xor ( n45987 , n45370 , n45536 );
and ( n45988 , n30274 , n45688 );
and ( n45989 , n45987 , n45988 );
xor ( n45990 , n45987 , n45988 );
xor ( n45991 , n45374 , n45534 );
and ( n45992 , n30279 , n45688 );
and ( n45993 , n45991 , n45992 );
xor ( n45994 , n45991 , n45992 );
xor ( n45995 , n45378 , n45532 );
and ( n45996 , n30284 , n45688 );
and ( n45997 , n45995 , n45996 );
xor ( n45998 , n45995 , n45996 );
xor ( n45999 , n45382 , n45530 );
and ( n46000 , n30289 , n45688 );
and ( n46001 , n45999 , n46000 );
xor ( n46002 , n45999 , n46000 );
xor ( n46003 , n45386 , n45528 );
and ( n46004 , n30294 , n45688 );
and ( n46005 , n46003 , n46004 );
xor ( n46006 , n46003 , n46004 );
xor ( n46007 , n45390 , n45526 );
and ( n46008 , n30299 , n45688 );
and ( n46009 , n46007 , n46008 );
xor ( n46010 , n46007 , n46008 );
xor ( n46011 , n45394 , n45524 );
and ( n46012 , n30304 , n45688 );
and ( n46013 , n46011 , n46012 );
xor ( n46014 , n46011 , n46012 );
xor ( n46015 , n45398 , n45522 );
and ( n46016 , n30309 , n45688 );
and ( n46017 , n46015 , n46016 );
xor ( n46018 , n46015 , n46016 );
xor ( n46019 , n45402 , n45520 );
and ( n46020 , n30314 , n45688 );
and ( n46021 , n46019 , n46020 );
xor ( n46022 , n46019 , n46020 );
xor ( n46023 , n45406 , n45518 );
and ( n46024 , n30319 , n45688 );
and ( n46025 , n46023 , n46024 );
xor ( n46026 , n46023 , n46024 );
xor ( n46027 , n45410 , n45516 );
and ( n46028 , n30324 , n45688 );
and ( n46029 , n46027 , n46028 );
xor ( n46030 , n46027 , n46028 );
xor ( n46031 , n45414 , n45514 );
and ( n46032 , n30329 , n45688 );
and ( n46033 , n46031 , n46032 );
xor ( n46034 , n46031 , n46032 );
xor ( n46035 , n45418 , n45512 );
and ( n46036 , n30334 , n45688 );
and ( n46037 , n46035 , n46036 );
xor ( n46038 , n46035 , n46036 );
xor ( n46039 , n45422 , n45510 );
and ( n46040 , n30339 , n45688 );
and ( n46041 , n46039 , n46040 );
xor ( n46042 , n46039 , n46040 );
xor ( n46043 , n45426 , n45508 );
and ( n46044 , n30344 , n45688 );
and ( n46045 , n46043 , n46044 );
xor ( n46046 , n46043 , n46044 );
xor ( n46047 , n45430 , n45506 );
and ( n46048 , n30349 , n45688 );
and ( n46049 , n46047 , n46048 );
xor ( n46050 , n46047 , n46048 );
xor ( n46051 , n45434 , n45504 );
and ( n46052 , n30354 , n45688 );
and ( n46053 , n46051 , n46052 );
xor ( n46054 , n46051 , n46052 );
xor ( n46055 , n45438 , n45502 );
and ( n46056 , n30359 , n45688 );
and ( n46057 , n46055 , n46056 );
xor ( n46058 , n46055 , n46056 );
xor ( n46059 , n45442 , n45500 );
and ( n46060 , n30364 , n45688 );
and ( n46061 , n46059 , n46060 );
xor ( n46062 , n46059 , n46060 );
xor ( n46063 , n45446 , n45498 );
and ( n46064 , n30369 , n45688 );
and ( n46065 , n46063 , n46064 );
xor ( n46066 , n46063 , n46064 );
xor ( n46067 , n45450 , n45496 );
and ( n46068 , n30374 , n45688 );
and ( n46069 , n46067 , n46068 );
xor ( n46070 , n46067 , n46068 );
xor ( n46071 , n45454 , n45494 );
and ( n46072 , n30379 , n45688 );
and ( n46073 , n46071 , n46072 );
xor ( n46074 , n46071 , n46072 );
xor ( n46075 , n45458 , n45492 );
and ( n46076 , n30384 , n45688 );
and ( n46077 , n46075 , n46076 );
xor ( n46078 , n46075 , n46076 );
xor ( n46079 , n45462 , n45490 );
and ( n46080 , n30389 , n45688 );
and ( n46081 , n46079 , n46080 );
xor ( n46082 , n46079 , n46080 );
xor ( n46083 , n45466 , n45488 );
and ( n46084 , n30394 , n45688 );
and ( n46085 , n46083 , n46084 );
xor ( n46086 , n46083 , n46084 );
xor ( n46087 , n45470 , n45486 );
and ( n46088 , n30399 , n45688 );
and ( n46089 , n46087 , n46088 );
xor ( n46090 , n46087 , n46088 );
xor ( n46091 , n45474 , n45484 );
and ( n46092 , n30404 , n45688 );
and ( n46093 , n46091 , n46092 );
xor ( n46094 , n46091 , n46092 );
xor ( n46095 , n45478 , n45482 );
and ( n46096 , n30409 , n45688 );
and ( n46097 , n46095 , n46096 );
buf ( n46098 , n46097 );
and ( n46099 , n46094 , n46098 );
or ( n46100 , n46093 , n46099 );
and ( n46101 , n46090 , n46100 );
or ( n46102 , n46089 , n46101 );
and ( n46103 , n46086 , n46102 );
or ( n46104 , n46085 , n46103 );
and ( n46105 , n46082 , n46104 );
or ( n46106 , n46081 , n46105 );
and ( n46107 , n46078 , n46106 );
or ( n46108 , n46077 , n46107 );
and ( n46109 , n46074 , n46108 );
or ( n46110 , n46073 , n46109 );
and ( n46111 , n46070 , n46110 );
or ( n46112 , n46069 , n46111 );
and ( n46113 , n46066 , n46112 );
or ( n46114 , n46065 , n46113 );
and ( n46115 , n46062 , n46114 );
or ( n46116 , n46061 , n46115 );
and ( n46117 , n46058 , n46116 );
or ( n46118 , n46057 , n46117 );
and ( n46119 , n46054 , n46118 );
or ( n46120 , n46053 , n46119 );
and ( n46121 , n46050 , n46120 );
or ( n46122 , n46049 , n46121 );
and ( n46123 , n46046 , n46122 );
or ( n46124 , n46045 , n46123 );
and ( n46125 , n46042 , n46124 );
or ( n46126 , n46041 , n46125 );
and ( n46127 , n46038 , n46126 );
or ( n46128 , n46037 , n46127 );
and ( n46129 , n46034 , n46128 );
or ( n46130 , n46033 , n46129 );
and ( n46131 , n46030 , n46130 );
or ( n46132 , n46029 , n46131 );
and ( n46133 , n46026 , n46132 );
or ( n46134 , n46025 , n46133 );
and ( n46135 , n46022 , n46134 );
or ( n46136 , n46021 , n46135 );
and ( n46137 , n46018 , n46136 );
or ( n46138 , n46017 , n46137 );
and ( n46139 , n46014 , n46138 );
or ( n46140 , n46013 , n46139 );
and ( n46141 , n46010 , n46140 );
or ( n46142 , n46009 , n46141 );
and ( n46143 , n46006 , n46142 );
or ( n46144 , n46005 , n46143 );
and ( n46145 , n46002 , n46144 );
or ( n46146 , n46001 , n46145 );
and ( n46147 , n45998 , n46146 );
or ( n46148 , n45997 , n46147 );
and ( n46149 , n45994 , n46148 );
or ( n46150 , n45993 , n46149 );
and ( n46151 , n45990 , n46150 );
or ( n46152 , n45989 , n46151 );
and ( n46153 , n45986 , n46152 );
or ( n46154 , n45985 , n46153 );
and ( n46155 , n45982 , n46154 );
or ( n46156 , n45981 , n46155 );
and ( n46157 , n45978 , n46156 );
or ( n46158 , n45977 , n46157 );
and ( n46159 , n45974 , n46158 );
or ( n46160 , n45973 , n46159 );
and ( n46161 , n45970 , n46160 );
or ( n46162 , n45969 , n46161 );
and ( n46163 , n45966 , n46162 );
or ( n46164 , n45965 , n46163 );
and ( n46165 , n45962 , n46164 );
or ( n46166 , n45961 , n46165 );
and ( n46167 , n45958 , n46166 );
or ( n46168 , n45957 , n46167 );
and ( n46169 , n45954 , n46168 );
or ( n46170 , n45953 , n46169 );
and ( n46171 , n45950 , n46170 );
or ( n46172 , n45949 , n46171 );
and ( n46173 , n45946 , n46172 );
or ( n46174 , n45945 , n46173 );
and ( n46175 , n45942 , n46174 );
or ( n46176 , n45941 , n46175 );
and ( n46177 , n45938 , n46176 );
or ( n46178 , n45937 , n46177 );
and ( n46179 , n45934 , n46178 );
or ( n46180 , n45933 , n46179 );
and ( n46181 , n45930 , n46180 );
or ( n46182 , n45929 , n46181 );
and ( n46183 , n45926 , n46182 );
or ( n46184 , n45925 , n46183 );
and ( n46185 , n45922 , n46184 );
or ( n46186 , n45921 , n46185 );
and ( n46187 , n45918 , n46186 );
or ( n46188 , n45917 , n46187 );
and ( n46189 , n45914 , n46188 );
or ( n46190 , n45913 , n46189 );
and ( n46191 , n45910 , n46190 );
or ( n46192 , n45909 , n46191 );
and ( n46193 , n45906 , n46192 );
or ( n46194 , n45905 , n46193 );
and ( n46195 , n45902 , n46194 );
or ( n46196 , n45901 , n46195 );
and ( n46197 , n45898 , n46196 );
or ( n46198 , n45897 , n46197 );
and ( n46199 , n45894 , n46198 );
or ( n46200 , n45893 , n46199 );
and ( n46201 , n45890 , n46200 );
or ( n46202 , n45889 , n46201 );
and ( n46203 , n45886 , n46202 );
or ( n46204 , n45885 , n46203 );
and ( n46205 , n45882 , n46204 );
or ( n46206 , n45881 , n46205 );
and ( n46207 , n45878 , n46206 );
or ( n46208 , n45877 , n46207 );
and ( n46209 , n45874 , n46208 );
or ( n46210 , n45873 , n46209 );
and ( n46211 , n45870 , n46210 );
or ( n46212 , n45869 , n46211 );
and ( n46213 , n45866 , n46212 );
or ( n46214 , n45865 , n46213 );
and ( n46215 , n45862 , n46214 );
or ( n46216 , n45861 , n46215 );
and ( n46217 , n45858 , n46216 );
or ( n46218 , n45857 , n46217 );
and ( n46219 , n45854 , n46218 );
or ( n46220 , n45853 , n46219 );
and ( n46221 , n45850 , n46220 );
or ( n46222 , n45849 , n46221 );
and ( n46223 , n45846 , n46222 );
or ( n46224 , n45845 , n46223 );
and ( n46225 , n45842 , n46224 );
or ( n46226 , n45841 , n46225 );
and ( n46227 , n45838 , n46226 );
or ( n46228 , n45837 , n46227 );
and ( n46229 , n45834 , n46228 );
or ( n46230 , n45833 , n46229 );
and ( n46231 , n45830 , n46230 );
or ( n46232 , n45829 , n46231 );
and ( n46233 , n45826 , n46232 );
or ( n46234 , n45825 , n46233 );
and ( n46235 , n45822 , n46234 );
or ( n46236 , n45821 , n46235 );
and ( n46237 , n45818 , n46236 );
or ( n46238 , n45817 , n46237 );
and ( n46239 , n45814 , n46238 );
or ( n46240 , n45813 , n46239 );
and ( n46241 , n45810 , n46240 );
or ( n46242 , n45809 , n46241 );
and ( n46243 , n45806 , n46242 );
or ( n46244 , n45805 , n46243 );
and ( n46245 , n45802 , n46244 );
or ( n46246 , n45801 , n46245 );
and ( n46247 , n45798 , n46246 );
or ( n46248 , n45797 , n46247 );
and ( n46249 , n45794 , n46248 );
or ( n46250 , n45793 , n46249 );
and ( n46251 , n45790 , n46250 );
or ( n46252 , n45789 , n46251 );
and ( n46253 , n45786 , n46252 );
or ( n46254 , n45785 , n46253 );
and ( n46255 , n45782 , n46254 );
or ( n46256 , n45781 , n46255 );
and ( n46257 , n45778 , n46256 );
or ( n46258 , n45777 , n46257 );
and ( n46259 , n45774 , n46258 );
or ( n46260 , n45773 , n46259 );
and ( n46261 , n45770 , n46260 );
or ( n46262 , n45769 , n46261 );
and ( n46263 , n45766 , n46262 );
or ( n46264 , n45765 , n46263 );
and ( n46265 , n45762 , n46264 );
or ( n46266 , n45761 , n46265 );
and ( n46267 , n45758 , n46266 );
or ( n46268 , n45757 , n46267 );
and ( n46269 , n45754 , n46268 );
or ( n46270 , n45753 , n46269 );
and ( n46271 , n45750 , n46270 );
or ( n46272 , n45749 , n46271 );
and ( n46273 , n45746 , n46272 );
or ( n46274 , n45745 , n46273 );
and ( n46275 , n45742 , n46274 );
or ( n46276 , n45741 , n46275 );
and ( n46277 , n45738 , n46276 );
or ( n46278 , n45737 , n46277 );
and ( n46279 , n45734 , n46278 );
or ( n46280 , n45733 , n46279 );
and ( n46281 , n45730 , n46280 );
or ( n46282 , n45729 , n46281 );
and ( n46283 , n45726 , n46282 );
or ( n46284 , n45725 , n46283 );
and ( n46285 , n45722 , n46284 );
or ( n46286 , n45721 , n46285 );
and ( n46287 , n45718 , n46286 );
or ( n46288 , n45717 , n46287 );
and ( n46289 , n45714 , n46288 );
or ( n46290 , n45713 , n46289 );
and ( n46291 , n45710 , n46290 );
or ( n46292 , n45709 , n46291 );
and ( n46293 , n45706 , n46292 );
or ( n46294 , n45705 , n46293 );
and ( n46295 , n45702 , n46294 );
or ( n46296 , n45701 , n46295 );
and ( n46297 , n45698 , n46296 );
or ( n46298 , n45697 , n46297 );
and ( n46299 , n45694 , n46298 );
or ( n46300 , n45693 , n46299 );
xor ( n46301 , n45690 , n46300 );
buf ( n46302 , n18056 );
and ( n46303 , n29904 , n46302 );
xor ( n46304 , n46301 , n46303 );
xor ( n46305 , n45694 , n46298 );
and ( n46306 , n29909 , n46302 );
and ( n46307 , n46305 , n46306 );
xor ( n46308 , n46305 , n46306 );
xor ( n46309 , n45698 , n46296 );
and ( n46310 , n29914 , n46302 );
and ( n46311 , n46309 , n46310 );
xor ( n46312 , n46309 , n46310 );
xor ( n46313 , n45702 , n46294 );
and ( n46314 , n29919 , n46302 );
and ( n46315 , n46313 , n46314 );
xor ( n46316 , n46313 , n46314 );
xor ( n46317 , n45706 , n46292 );
and ( n46318 , n29924 , n46302 );
and ( n46319 , n46317 , n46318 );
xor ( n46320 , n46317 , n46318 );
xor ( n46321 , n45710 , n46290 );
and ( n46322 , n29929 , n46302 );
and ( n46323 , n46321 , n46322 );
xor ( n46324 , n46321 , n46322 );
xor ( n46325 , n45714 , n46288 );
and ( n46326 , n29934 , n46302 );
and ( n46327 , n46325 , n46326 );
xor ( n46328 , n46325 , n46326 );
xor ( n46329 , n45718 , n46286 );
and ( n46330 , n29939 , n46302 );
and ( n46331 , n46329 , n46330 );
xor ( n46332 , n46329 , n46330 );
xor ( n46333 , n45722 , n46284 );
and ( n46334 , n29944 , n46302 );
and ( n46335 , n46333 , n46334 );
xor ( n46336 , n46333 , n46334 );
xor ( n46337 , n45726 , n46282 );
and ( n46338 , n29949 , n46302 );
and ( n46339 , n46337 , n46338 );
xor ( n46340 , n46337 , n46338 );
xor ( n46341 , n45730 , n46280 );
and ( n46342 , n29954 , n46302 );
and ( n46343 , n46341 , n46342 );
xor ( n46344 , n46341 , n46342 );
xor ( n46345 , n45734 , n46278 );
and ( n46346 , n29959 , n46302 );
and ( n46347 , n46345 , n46346 );
xor ( n46348 , n46345 , n46346 );
xor ( n46349 , n45738 , n46276 );
and ( n46350 , n29964 , n46302 );
and ( n46351 , n46349 , n46350 );
xor ( n46352 , n46349 , n46350 );
xor ( n46353 , n45742 , n46274 );
and ( n46354 , n29969 , n46302 );
and ( n46355 , n46353 , n46354 );
xor ( n46356 , n46353 , n46354 );
xor ( n46357 , n45746 , n46272 );
and ( n46358 , n29974 , n46302 );
and ( n46359 , n46357 , n46358 );
xor ( n46360 , n46357 , n46358 );
xor ( n46361 , n45750 , n46270 );
and ( n46362 , n29979 , n46302 );
and ( n46363 , n46361 , n46362 );
xor ( n46364 , n46361 , n46362 );
xor ( n46365 , n45754 , n46268 );
and ( n46366 , n29984 , n46302 );
and ( n46367 , n46365 , n46366 );
xor ( n46368 , n46365 , n46366 );
xor ( n46369 , n45758 , n46266 );
and ( n46370 , n29989 , n46302 );
and ( n46371 , n46369 , n46370 );
xor ( n46372 , n46369 , n46370 );
xor ( n46373 , n45762 , n46264 );
and ( n46374 , n29994 , n46302 );
and ( n46375 , n46373 , n46374 );
xor ( n46376 , n46373 , n46374 );
xor ( n46377 , n45766 , n46262 );
and ( n46378 , n29999 , n46302 );
and ( n46379 , n46377 , n46378 );
xor ( n46380 , n46377 , n46378 );
xor ( n46381 , n45770 , n46260 );
and ( n46382 , n30004 , n46302 );
and ( n46383 , n46381 , n46382 );
xor ( n46384 , n46381 , n46382 );
xor ( n46385 , n45774 , n46258 );
and ( n46386 , n30009 , n46302 );
and ( n46387 , n46385 , n46386 );
xor ( n46388 , n46385 , n46386 );
xor ( n46389 , n45778 , n46256 );
and ( n46390 , n30014 , n46302 );
and ( n46391 , n46389 , n46390 );
xor ( n46392 , n46389 , n46390 );
xor ( n46393 , n45782 , n46254 );
and ( n46394 , n30019 , n46302 );
and ( n46395 , n46393 , n46394 );
xor ( n46396 , n46393 , n46394 );
xor ( n46397 , n45786 , n46252 );
and ( n46398 , n30024 , n46302 );
and ( n46399 , n46397 , n46398 );
xor ( n46400 , n46397 , n46398 );
xor ( n46401 , n45790 , n46250 );
and ( n46402 , n30029 , n46302 );
and ( n46403 , n46401 , n46402 );
xor ( n46404 , n46401 , n46402 );
xor ( n46405 , n45794 , n46248 );
and ( n46406 , n30034 , n46302 );
and ( n46407 , n46405 , n46406 );
xor ( n46408 , n46405 , n46406 );
xor ( n46409 , n45798 , n46246 );
and ( n46410 , n30039 , n46302 );
and ( n46411 , n46409 , n46410 );
xor ( n46412 , n46409 , n46410 );
xor ( n46413 , n45802 , n46244 );
and ( n46414 , n30044 , n46302 );
and ( n46415 , n46413 , n46414 );
xor ( n46416 , n46413 , n46414 );
xor ( n46417 , n45806 , n46242 );
and ( n46418 , n30049 , n46302 );
and ( n46419 , n46417 , n46418 );
xor ( n46420 , n46417 , n46418 );
xor ( n46421 , n45810 , n46240 );
and ( n46422 , n30054 , n46302 );
and ( n46423 , n46421 , n46422 );
xor ( n46424 , n46421 , n46422 );
xor ( n46425 , n45814 , n46238 );
and ( n46426 , n30059 , n46302 );
and ( n46427 , n46425 , n46426 );
xor ( n46428 , n46425 , n46426 );
xor ( n46429 , n45818 , n46236 );
and ( n46430 , n30064 , n46302 );
and ( n46431 , n46429 , n46430 );
xor ( n46432 , n46429 , n46430 );
xor ( n46433 , n45822 , n46234 );
and ( n46434 , n30069 , n46302 );
and ( n46435 , n46433 , n46434 );
xor ( n46436 , n46433 , n46434 );
xor ( n46437 , n45826 , n46232 );
and ( n46438 , n30074 , n46302 );
and ( n46439 , n46437 , n46438 );
xor ( n46440 , n46437 , n46438 );
xor ( n46441 , n45830 , n46230 );
and ( n46442 , n30079 , n46302 );
and ( n46443 , n46441 , n46442 );
xor ( n46444 , n46441 , n46442 );
xor ( n46445 , n45834 , n46228 );
and ( n46446 , n30084 , n46302 );
and ( n46447 , n46445 , n46446 );
xor ( n46448 , n46445 , n46446 );
xor ( n46449 , n45838 , n46226 );
and ( n46450 , n30089 , n46302 );
and ( n46451 , n46449 , n46450 );
xor ( n46452 , n46449 , n46450 );
xor ( n46453 , n45842 , n46224 );
and ( n46454 , n30094 , n46302 );
and ( n46455 , n46453 , n46454 );
xor ( n46456 , n46453 , n46454 );
xor ( n46457 , n45846 , n46222 );
and ( n46458 , n30099 , n46302 );
and ( n46459 , n46457 , n46458 );
xor ( n46460 , n46457 , n46458 );
xor ( n46461 , n45850 , n46220 );
and ( n46462 , n30104 , n46302 );
and ( n46463 , n46461 , n46462 );
xor ( n46464 , n46461 , n46462 );
xor ( n46465 , n45854 , n46218 );
and ( n46466 , n30109 , n46302 );
and ( n46467 , n46465 , n46466 );
xor ( n46468 , n46465 , n46466 );
xor ( n46469 , n45858 , n46216 );
and ( n46470 , n30114 , n46302 );
and ( n46471 , n46469 , n46470 );
xor ( n46472 , n46469 , n46470 );
xor ( n46473 , n45862 , n46214 );
and ( n46474 , n30119 , n46302 );
and ( n46475 , n46473 , n46474 );
xor ( n46476 , n46473 , n46474 );
xor ( n46477 , n45866 , n46212 );
and ( n46478 , n30124 , n46302 );
and ( n46479 , n46477 , n46478 );
xor ( n46480 , n46477 , n46478 );
xor ( n46481 , n45870 , n46210 );
and ( n46482 , n30129 , n46302 );
and ( n46483 , n46481 , n46482 );
xor ( n46484 , n46481 , n46482 );
xor ( n46485 , n45874 , n46208 );
and ( n46486 , n30134 , n46302 );
and ( n46487 , n46485 , n46486 );
xor ( n46488 , n46485 , n46486 );
xor ( n46489 , n45878 , n46206 );
and ( n46490 , n30139 , n46302 );
and ( n46491 , n46489 , n46490 );
xor ( n46492 , n46489 , n46490 );
xor ( n46493 , n45882 , n46204 );
and ( n46494 , n30144 , n46302 );
and ( n46495 , n46493 , n46494 );
xor ( n46496 , n46493 , n46494 );
xor ( n46497 , n45886 , n46202 );
and ( n46498 , n30149 , n46302 );
and ( n46499 , n46497 , n46498 );
xor ( n46500 , n46497 , n46498 );
xor ( n46501 , n45890 , n46200 );
and ( n46502 , n30154 , n46302 );
and ( n46503 , n46501 , n46502 );
xor ( n46504 , n46501 , n46502 );
xor ( n46505 , n45894 , n46198 );
and ( n46506 , n30159 , n46302 );
and ( n46507 , n46505 , n46506 );
xor ( n46508 , n46505 , n46506 );
xor ( n46509 , n45898 , n46196 );
and ( n46510 , n30164 , n46302 );
and ( n46511 , n46509 , n46510 );
xor ( n46512 , n46509 , n46510 );
xor ( n46513 , n45902 , n46194 );
and ( n46514 , n30169 , n46302 );
and ( n46515 , n46513 , n46514 );
xor ( n46516 , n46513 , n46514 );
xor ( n46517 , n45906 , n46192 );
and ( n46518 , n30174 , n46302 );
and ( n46519 , n46517 , n46518 );
xor ( n46520 , n46517 , n46518 );
xor ( n46521 , n45910 , n46190 );
and ( n46522 , n30179 , n46302 );
and ( n46523 , n46521 , n46522 );
xor ( n46524 , n46521 , n46522 );
xor ( n46525 , n45914 , n46188 );
and ( n46526 , n30184 , n46302 );
and ( n46527 , n46525 , n46526 );
xor ( n46528 , n46525 , n46526 );
xor ( n46529 , n45918 , n46186 );
and ( n46530 , n30189 , n46302 );
and ( n46531 , n46529 , n46530 );
xor ( n46532 , n46529 , n46530 );
xor ( n46533 , n45922 , n46184 );
and ( n46534 , n30194 , n46302 );
and ( n46535 , n46533 , n46534 );
xor ( n46536 , n46533 , n46534 );
xor ( n46537 , n45926 , n46182 );
and ( n46538 , n30199 , n46302 );
and ( n46539 , n46537 , n46538 );
xor ( n46540 , n46537 , n46538 );
xor ( n46541 , n45930 , n46180 );
and ( n46542 , n30204 , n46302 );
and ( n46543 , n46541 , n46542 );
xor ( n46544 , n46541 , n46542 );
xor ( n46545 , n45934 , n46178 );
and ( n46546 , n30209 , n46302 );
and ( n46547 , n46545 , n46546 );
xor ( n46548 , n46545 , n46546 );
xor ( n46549 , n45938 , n46176 );
and ( n46550 , n30214 , n46302 );
and ( n46551 , n46549 , n46550 );
xor ( n46552 , n46549 , n46550 );
xor ( n46553 , n45942 , n46174 );
and ( n46554 , n30219 , n46302 );
and ( n46555 , n46553 , n46554 );
xor ( n46556 , n46553 , n46554 );
xor ( n46557 , n45946 , n46172 );
and ( n46558 , n30224 , n46302 );
and ( n46559 , n46557 , n46558 );
xor ( n46560 , n46557 , n46558 );
xor ( n46561 , n45950 , n46170 );
and ( n46562 , n30229 , n46302 );
and ( n46563 , n46561 , n46562 );
xor ( n46564 , n46561 , n46562 );
xor ( n46565 , n45954 , n46168 );
and ( n46566 , n30234 , n46302 );
and ( n46567 , n46565 , n46566 );
xor ( n46568 , n46565 , n46566 );
xor ( n46569 , n45958 , n46166 );
and ( n46570 , n30239 , n46302 );
and ( n46571 , n46569 , n46570 );
xor ( n46572 , n46569 , n46570 );
xor ( n46573 , n45962 , n46164 );
and ( n46574 , n30244 , n46302 );
and ( n46575 , n46573 , n46574 );
xor ( n46576 , n46573 , n46574 );
xor ( n46577 , n45966 , n46162 );
and ( n46578 , n30249 , n46302 );
and ( n46579 , n46577 , n46578 );
xor ( n46580 , n46577 , n46578 );
xor ( n46581 , n45970 , n46160 );
and ( n46582 , n30254 , n46302 );
and ( n46583 , n46581 , n46582 );
xor ( n46584 , n46581 , n46582 );
xor ( n46585 , n45974 , n46158 );
and ( n46586 , n30259 , n46302 );
and ( n46587 , n46585 , n46586 );
xor ( n46588 , n46585 , n46586 );
xor ( n46589 , n45978 , n46156 );
and ( n46590 , n30264 , n46302 );
and ( n46591 , n46589 , n46590 );
xor ( n46592 , n46589 , n46590 );
xor ( n46593 , n45982 , n46154 );
and ( n46594 , n30269 , n46302 );
and ( n46595 , n46593 , n46594 );
xor ( n46596 , n46593 , n46594 );
xor ( n46597 , n45986 , n46152 );
and ( n46598 , n30274 , n46302 );
and ( n46599 , n46597 , n46598 );
xor ( n46600 , n46597 , n46598 );
xor ( n46601 , n45990 , n46150 );
and ( n46602 , n30279 , n46302 );
and ( n46603 , n46601 , n46602 );
xor ( n46604 , n46601 , n46602 );
xor ( n46605 , n45994 , n46148 );
and ( n46606 , n30284 , n46302 );
and ( n46607 , n46605 , n46606 );
xor ( n46608 , n46605 , n46606 );
xor ( n46609 , n45998 , n46146 );
and ( n46610 , n30289 , n46302 );
and ( n46611 , n46609 , n46610 );
xor ( n46612 , n46609 , n46610 );
xor ( n46613 , n46002 , n46144 );
and ( n46614 , n30294 , n46302 );
and ( n46615 , n46613 , n46614 );
xor ( n46616 , n46613 , n46614 );
xor ( n46617 , n46006 , n46142 );
and ( n46618 , n30299 , n46302 );
and ( n46619 , n46617 , n46618 );
xor ( n46620 , n46617 , n46618 );
xor ( n46621 , n46010 , n46140 );
and ( n46622 , n30304 , n46302 );
and ( n46623 , n46621 , n46622 );
xor ( n46624 , n46621 , n46622 );
xor ( n46625 , n46014 , n46138 );
and ( n46626 , n30309 , n46302 );
and ( n46627 , n46625 , n46626 );
xor ( n46628 , n46625 , n46626 );
xor ( n46629 , n46018 , n46136 );
and ( n46630 , n30314 , n46302 );
and ( n46631 , n46629 , n46630 );
xor ( n46632 , n46629 , n46630 );
xor ( n46633 , n46022 , n46134 );
and ( n46634 , n30319 , n46302 );
and ( n46635 , n46633 , n46634 );
xor ( n46636 , n46633 , n46634 );
xor ( n46637 , n46026 , n46132 );
and ( n46638 , n30324 , n46302 );
and ( n46639 , n46637 , n46638 );
xor ( n46640 , n46637 , n46638 );
xor ( n46641 , n46030 , n46130 );
and ( n46642 , n30329 , n46302 );
and ( n46643 , n46641 , n46642 );
xor ( n46644 , n46641 , n46642 );
xor ( n46645 , n46034 , n46128 );
and ( n46646 , n30334 , n46302 );
and ( n46647 , n46645 , n46646 );
xor ( n46648 , n46645 , n46646 );
xor ( n46649 , n46038 , n46126 );
and ( n46650 , n30339 , n46302 );
and ( n46651 , n46649 , n46650 );
xor ( n46652 , n46649 , n46650 );
xor ( n46653 , n46042 , n46124 );
and ( n46654 , n30344 , n46302 );
and ( n46655 , n46653 , n46654 );
xor ( n46656 , n46653 , n46654 );
xor ( n46657 , n46046 , n46122 );
and ( n46658 , n30349 , n46302 );
and ( n46659 , n46657 , n46658 );
xor ( n46660 , n46657 , n46658 );
xor ( n46661 , n46050 , n46120 );
and ( n46662 , n30354 , n46302 );
and ( n46663 , n46661 , n46662 );
xor ( n46664 , n46661 , n46662 );
xor ( n46665 , n46054 , n46118 );
and ( n46666 , n30359 , n46302 );
and ( n46667 , n46665 , n46666 );
xor ( n46668 , n46665 , n46666 );
xor ( n46669 , n46058 , n46116 );
and ( n46670 , n30364 , n46302 );
and ( n46671 , n46669 , n46670 );
xor ( n46672 , n46669 , n46670 );
xor ( n46673 , n46062 , n46114 );
and ( n46674 , n30369 , n46302 );
and ( n46675 , n46673 , n46674 );
xor ( n46676 , n46673 , n46674 );
xor ( n46677 , n46066 , n46112 );
and ( n46678 , n30374 , n46302 );
and ( n46679 , n46677 , n46678 );
xor ( n46680 , n46677 , n46678 );
xor ( n46681 , n46070 , n46110 );
and ( n46682 , n30379 , n46302 );
and ( n46683 , n46681 , n46682 );
xor ( n46684 , n46681 , n46682 );
xor ( n46685 , n46074 , n46108 );
and ( n46686 , n30384 , n46302 );
and ( n46687 , n46685 , n46686 );
xor ( n46688 , n46685 , n46686 );
xor ( n46689 , n46078 , n46106 );
and ( n46690 , n30389 , n46302 );
and ( n46691 , n46689 , n46690 );
xor ( n46692 , n46689 , n46690 );
xor ( n46693 , n46082 , n46104 );
and ( n46694 , n30394 , n46302 );
and ( n46695 , n46693 , n46694 );
xor ( n46696 , n46693 , n46694 );
xor ( n46697 , n46086 , n46102 );
and ( n46698 , n30399 , n46302 );
and ( n46699 , n46697 , n46698 );
xor ( n46700 , n46697 , n46698 );
xor ( n46701 , n46090 , n46100 );
and ( n46702 , n30404 , n46302 );
and ( n46703 , n46701 , n46702 );
xor ( n46704 , n46701 , n46702 );
xor ( n46705 , n46094 , n46098 );
and ( n46706 , n30409 , n46302 );
and ( n46707 , n46705 , n46706 );
buf ( n46708 , n46707 );
and ( n46709 , n46704 , n46708 );
or ( n46710 , n46703 , n46709 );
and ( n46711 , n46700 , n46710 );
or ( n46712 , n46699 , n46711 );
and ( n46713 , n46696 , n46712 );
or ( n46714 , n46695 , n46713 );
and ( n46715 , n46692 , n46714 );
or ( n46716 , n46691 , n46715 );
and ( n46717 , n46688 , n46716 );
or ( n46718 , n46687 , n46717 );
and ( n46719 , n46684 , n46718 );
or ( n46720 , n46683 , n46719 );
and ( n46721 , n46680 , n46720 );
or ( n46722 , n46679 , n46721 );
and ( n46723 , n46676 , n46722 );
or ( n46724 , n46675 , n46723 );
and ( n46725 , n46672 , n46724 );
or ( n46726 , n46671 , n46725 );
and ( n46727 , n46668 , n46726 );
or ( n46728 , n46667 , n46727 );
and ( n46729 , n46664 , n46728 );
or ( n46730 , n46663 , n46729 );
and ( n46731 , n46660 , n46730 );
or ( n46732 , n46659 , n46731 );
and ( n46733 , n46656 , n46732 );
or ( n46734 , n46655 , n46733 );
and ( n46735 , n46652 , n46734 );
or ( n46736 , n46651 , n46735 );
and ( n46737 , n46648 , n46736 );
or ( n46738 , n46647 , n46737 );
and ( n46739 , n46644 , n46738 );
or ( n46740 , n46643 , n46739 );
and ( n46741 , n46640 , n46740 );
or ( n46742 , n46639 , n46741 );
and ( n46743 , n46636 , n46742 );
or ( n46744 , n46635 , n46743 );
and ( n46745 , n46632 , n46744 );
or ( n46746 , n46631 , n46745 );
and ( n46747 , n46628 , n46746 );
or ( n46748 , n46627 , n46747 );
and ( n46749 , n46624 , n46748 );
or ( n46750 , n46623 , n46749 );
and ( n46751 , n46620 , n46750 );
or ( n46752 , n46619 , n46751 );
and ( n46753 , n46616 , n46752 );
or ( n46754 , n46615 , n46753 );
and ( n46755 , n46612 , n46754 );
or ( n46756 , n46611 , n46755 );
and ( n46757 , n46608 , n46756 );
or ( n46758 , n46607 , n46757 );
and ( n46759 , n46604 , n46758 );
or ( n46760 , n46603 , n46759 );
and ( n46761 , n46600 , n46760 );
or ( n46762 , n46599 , n46761 );
and ( n46763 , n46596 , n46762 );
or ( n46764 , n46595 , n46763 );
and ( n46765 , n46592 , n46764 );
or ( n46766 , n46591 , n46765 );
and ( n46767 , n46588 , n46766 );
or ( n46768 , n46587 , n46767 );
and ( n46769 , n46584 , n46768 );
or ( n46770 , n46583 , n46769 );
and ( n46771 , n46580 , n46770 );
or ( n46772 , n46579 , n46771 );
and ( n46773 , n46576 , n46772 );
or ( n46774 , n46575 , n46773 );
and ( n46775 , n46572 , n46774 );
or ( n46776 , n46571 , n46775 );
and ( n46777 , n46568 , n46776 );
or ( n46778 , n46567 , n46777 );
and ( n46779 , n46564 , n46778 );
or ( n46780 , n46563 , n46779 );
and ( n46781 , n46560 , n46780 );
or ( n46782 , n46559 , n46781 );
and ( n46783 , n46556 , n46782 );
or ( n46784 , n46555 , n46783 );
and ( n46785 , n46552 , n46784 );
or ( n46786 , n46551 , n46785 );
and ( n46787 , n46548 , n46786 );
or ( n46788 , n46547 , n46787 );
and ( n46789 , n46544 , n46788 );
or ( n46790 , n46543 , n46789 );
and ( n46791 , n46540 , n46790 );
or ( n46792 , n46539 , n46791 );
and ( n46793 , n46536 , n46792 );
or ( n46794 , n46535 , n46793 );
and ( n46795 , n46532 , n46794 );
or ( n46796 , n46531 , n46795 );
and ( n46797 , n46528 , n46796 );
or ( n46798 , n46527 , n46797 );
and ( n46799 , n46524 , n46798 );
or ( n46800 , n46523 , n46799 );
and ( n46801 , n46520 , n46800 );
or ( n46802 , n46519 , n46801 );
and ( n46803 , n46516 , n46802 );
or ( n46804 , n46515 , n46803 );
and ( n46805 , n46512 , n46804 );
or ( n46806 , n46511 , n46805 );
and ( n46807 , n46508 , n46806 );
or ( n46808 , n46507 , n46807 );
and ( n46809 , n46504 , n46808 );
or ( n46810 , n46503 , n46809 );
and ( n46811 , n46500 , n46810 );
or ( n46812 , n46499 , n46811 );
and ( n46813 , n46496 , n46812 );
or ( n46814 , n46495 , n46813 );
and ( n46815 , n46492 , n46814 );
or ( n46816 , n46491 , n46815 );
and ( n46817 , n46488 , n46816 );
or ( n46818 , n46487 , n46817 );
and ( n46819 , n46484 , n46818 );
or ( n46820 , n46483 , n46819 );
and ( n46821 , n46480 , n46820 );
or ( n46822 , n46479 , n46821 );
and ( n46823 , n46476 , n46822 );
or ( n46824 , n46475 , n46823 );
and ( n46825 , n46472 , n46824 );
or ( n46826 , n46471 , n46825 );
and ( n46827 , n46468 , n46826 );
or ( n46828 , n46467 , n46827 );
and ( n46829 , n46464 , n46828 );
or ( n46830 , n46463 , n46829 );
and ( n46831 , n46460 , n46830 );
or ( n46832 , n46459 , n46831 );
and ( n46833 , n46456 , n46832 );
or ( n46834 , n46455 , n46833 );
and ( n46835 , n46452 , n46834 );
or ( n46836 , n46451 , n46835 );
and ( n46837 , n46448 , n46836 );
or ( n46838 , n46447 , n46837 );
and ( n46839 , n46444 , n46838 );
or ( n46840 , n46443 , n46839 );
and ( n46841 , n46440 , n46840 );
or ( n46842 , n46439 , n46841 );
and ( n46843 , n46436 , n46842 );
or ( n46844 , n46435 , n46843 );
and ( n46845 , n46432 , n46844 );
or ( n46846 , n46431 , n46845 );
and ( n46847 , n46428 , n46846 );
or ( n46848 , n46427 , n46847 );
and ( n46849 , n46424 , n46848 );
or ( n46850 , n46423 , n46849 );
and ( n46851 , n46420 , n46850 );
or ( n46852 , n46419 , n46851 );
and ( n46853 , n46416 , n46852 );
or ( n46854 , n46415 , n46853 );
and ( n46855 , n46412 , n46854 );
or ( n46856 , n46411 , n46855 );
and ( n46857 , n46408 , n46856 );
or ( n46858 , n46407 , n46857 );
and ( n46859 , n46404 , n46858 );
or ( n46860 , n46403 , n46859 );
and ( n46861 , n46400 , n46860 );
or ( n46862 , n46399 , n46861 );
and ( n46863 , n46396 , n46862 );
or ( n46864 , n46395 , n46863 );
and ( n46865 , n46392 , n46864 );
or ( n46866 , n46391 , n46865 );
and ( n46867 , n46388 , n46866 );
or ( n46868 , n46387 , n46867 );
and ( n46869 , n46384 , n46868 );
or ( n46870 , n46383 , n46869 );
and ( n46871 , n46380 , n46870 );
or ( n46872 , n46379 , n46871 );
and ( n46873 , n46376 , n46872 );
or ( n46874 , n46375 , n46873 );
and ( n46875 , n46372 , n46874 );
or ( n46876 , n46371 , n46875 );
and ( n46877 , n46368 , n46876 );
or ( n46878 , n46367 , n46877 );
and ( n46879 , n46364 , n46878 );
or ( n46880 , n46363 , n46879 );
and ( n46881 , n46360 , n46880 );
or ( n46882 , n46359 , n46881 );
and ( n46883 , n46356 , n46882 );
or ( n46884 , n46355 , n46883 );
and ( n46885 , n46352 , n46884 );
or ( n46886 , n46351 , n46885 );
and ( n46887 , n46348 , n46886 );
or ( n46888 , n46347 , n46887 );
and ( n46889 , n46344 , n46888 );
or ( n46890 , n46343 , n46889 );
and ( n46891 , n46340 , n46890 );
or ( n46892 , n46339 , n46891 );
and ( n46893 , n46336 , n46892 );
or ( n46894 , n46335 , n46893 );
and ( n46895 , n46332 , n46894 );
or ( n46896 , n46331 , n46895 );
and ( n46897 , n46328 , n46896 );
or ( n46898 , n46327 , n46897 );
and ( n46899 , n46324 , n46898 );
or ( n46900 , n46323 , n46899 );
and ( n46901 , n46320 , n46900 );
or ( n46902 , n46319 , n46901 );
and ( n46903 , n46316 , n46902 );
or ( n46904 , n46315 , n46903 );
and ( n46905 , n46312 , n46904 );
or ( n46906 , n46311 , n46905 );
and ( n46907 , n46308 , n46906 );
or ( n46908 , n46307 , n46907 );
xor ( n46909 , n46304 , n46908 );
buf ( n46910 , n18054 );
and ( n46911 , n29909 , n46910 );
xor ( n46912 , n46909 , n46911 );
xor ( n46913 , n46308 , n46906 );
and ( n46914 , n29914 , n46910 );
and ( n46915 , n46913 , n46914 );
xor ( n46916 , n46913 , n46914 );
xor ( n46917 , n46312 , n46904 );
and ( n46918 , n29919 , n46910 );
and ( n46919 , n46917 , n46918 );
xor ( n46920 , n46917 , n46918 );
xor ( n46921 , n46316 , n46902 );
and ( n46922 , n29924 , n46910 );
and ( n46923 , n46921 , n46922 );
xor ( n46924 , n46921 , n46922 );
xor ( n46925 , n46320 , n46900 );
and ( n46926 , n29929 , n46910 );
and ( n46927 , n46925 , n46926 );
xor ( n46928 , n46925 , n46926 );
xor ( n46929 , n46324 , n46898 );
and ( n46930 , n29934 , n46910 );
and ( n46931 , n46929 , n46930 );
xor ( n46932 , n46929 , n46930 );
xor ( n46933 , n46328 , n46896 );
and ( n46934 , n29939 , n46910 );
and ( n46935 , n46933 , n46934 );
xor ( n46936 , n46933 , n46934 );
xor ( n46937 , n46332 , n46894 );
and ( n46938 , n29944 , n46910 );
and ( n46939 , n46937 , n46938 );
xor ( n46940 , n46937 , n46938 );
xor ( n46941 , n46336 , n46892 );
and ( n46942 , n29949 , n46910 );
and ( n46943 , n46941 , n46942 );
xor ( n46944 , n46941 , n46942 );
xor ( n46945 , n46340 , n46890 );
and ( n46946 , n29954 , n46910 );
and ( n46947 , n46945 , n46946 );
xor ( n46948 , n46945 , n46946 );
xor ( n46949 , n46344 , n46888 );
and ( n46950 , n29959 , n46910 );
and ( n46951 , n46949 , n46950 );
xor ( n46952 , n46949 , n46950 );
xor ( n46953 , n46348 , n46886 );
and ( n46954 , n29964 , n46910 );
and ( n46955 , n46953 , n46954 );
xor ( n46956 , n46953 , n46954 );
xor ( n46957 , n46352 , n46884 );
and ( n46958 , n29969 , n46910 );
and ( n46959 , n46957 , n46958 );
xor ( n46960 , n46957 , n46958 );
xor ( n46961 , n46356 , n46882 );
and ( n46962 , n29974 , n46910 );
and ( n46963 , n46961 , n46962 );
xor ( n46964 , n46961 , n46962 );
xor ( n46965 , n46360 , n46880 );
and ( n46966 , n29979 , n46910 );
and ( n46967 , n46965 , n46966 );
xor ( n46968 , n46965 , n46966 );
xor ( n46969 , n46364 , n46878 );
and ( n46970 , n29984 , n46910 );
and ( n46971 , n46969 , n46970 );
xor ( n46972 , n46969 , n46970 );
xor ( n46973 , n46368 , n46876 );
and ( n46974 , n29989 , n46910 );
and ( n46975 , n46973 , n46974 );
xor ( n46976 , n46973 , n46974 );
xor ( n46977 , n46372 , n46874 );
and ( n46978 , n29994 , n46910 );
and ( n46979 , n46977 , n46978 );
xor ( n46980 , n46977 , n46978 );
xor ( n46981 , n46376 , n46872 );
and ( n46982 , n29999 , n46910 );
and ( n46983 , n46981 , n46982 );
xor ( n46984 , n46981 , n46982 );
xor ( n46985 , n46380 , n46870 );
and ( n46986 , n30004 , n46910 );
and ( n46987 , n46985 , n46986 );
xor ( n46988 , n46985 , n46986 );
xor ( n46989 , n46384 , n46868 );
and ( n46990 , n30009 , n46910 );
and ( n46991 , n46989 , n46990 );
xor ( n46992 , n46989 , n46990 );
xor ( n46993 , n46388 , n46866 );
and ( n46994 , n30014 , n46910 );
and ( n46995 , n46993 , n46994 );
xor ( n46996 , n46993 , n46994 );
xor ( n46997 , n46392 , n46864 );
and ( n46998 , n30019 , n46910 );
and ( n46999 , n46997 , n46998 );
xor ( n47000 , n46997 , n46998 );
xor ( n47001 , n46396 , n46862 );
and ( n47002 , n30024 , n46910 );
and ( n47003 , n47001 , n47002 );
xor ( n47004 , n47001 , n47002 );
xor ( n47005 , n46400 , n46860 );
and ( n47006 , n30029 , n46910 );
and ( n47007 , n47005 , n47006 );
xor ( n47008 , n47005 , n47006 );
xor ( n47009 , n46404 , n46858 );
and ( n47010 , n30034 , n46910 );
and ( n47011 , n47009 , n47010 );
xor ( n47012 , n47009 , n47010 );
xor ( n47013 , n46408 , n46856 );
and ( n47014 , n30039 , n46910 );
and ( n47015 , n47013 , n47014 );
xor ( n47016 , n47013 , n47014 );
xor ( n47017 , n46412 , n46854 );
and ( n47018 , n30044 , n46910 );
and ( n47019 , n47017 , n47018 );
xor ( n47020 , n47017 , n47018 );
xor ( n47021 , n46416 , n46852 );
and ( n47022 , n30049 , n46910 );
and ( n47023 , n47021 , n47022 );
xor ( n47024 , n47021 , n47022 );
xor ( n47025 , n46420 , n46850 );
and ( n47026 , n30054 , n46910 );
and ( n47027 , n47025 , n47026 );
xor ( n47028 , n47025 , n47026 );
xor ( n47029 , n46424 , n46848 );
and ( n47030 , n30059 , n46910 );
and ( n47031 , n47029 , n47030 );
xor ( n47032 , n47029 , n47030 );
xor ( n47033 , n46428 , n46846 );
and ( n47034 , n30064 , n46910 );
and ( n47035 , n47033 , n47034 );
xor ( n47036 , n47033 , n47034 );
xor ( n47037 , n46432 , n46844 );
and ( n47038 , n30069 , n46910 );
and ( n47039 , n47037 , n47038 );
xor ( n47040 , n47037 , n47038 );
xor ( n47041 , n46436 , n46842 );
and ( n47042 , n30074 , n46910 );
and ( n47043 , n47041 , n47042 );
xor ( n47044 , n47041 , n47042 );
xor ( n47045 , n46440 , n46840 );
and ( n47046 , n30079 , n46910 );
and ( n47047 , n47045 , n47046 );
xor ( n47048 , n47045 , n47046 );
xor ( n47049 , n46444 , n46838 );
and ( n47050 , n30084 , n46910 );
and ( n47051 , n47049 , n47050 );
xor ( n47052 , n47049 , n47050 );
xor ( n47053 , n46448 , n46836 );
and ( n47054 , n30089 , n46910 );
and ( n47055 , n47053 , n47054 );
xor ( n47056 , n47053 , n47054 );
xor ( n47057 , n46452 , n46834 );
and ( n47058 , n30094 , n46910 );
and ( n47059 , n47057 , n47058 );
xor ( n47060 , n47057 , n47058 );
xor ( n47061 , n46456 , n46832 );
and ( n47062 , n30099 , n46910 );
and ( n47063 , n47061 , n47062 );
xor ( n47064 , n47061 , n47062 );
xor ( n47065 , n46460 , n46830 );
and ( n47066 , n30104 , n46910 );
and ( n47067 , n47065 , n47066 );
xor ( n47068 , n47065 , n47066 );
xor ( n47069 , n46464 , n46828 );
and ( n47070 , n30109 , n46910 );
and ( n47071 , n47069 , n47070 );
xor ( n47072 , n47069 , n47070 );
xor ( n47073 , n46468 , n46826 );
and ( n47074 , n30114 , n46910 );
and ( n47075 , n47073 , n47074 );
xor ( n47076 , n47073 , n47074 );
xor ( n47077 , n46472 , n46824 );
and ( n47078 , n30119 , n46910 );
and ( n47079 , n47077 , n47078 );
xor ( n47080 , n47077 , n47078 );
xor ( n47081 , n46476 , n46822 );
and ( n47082 , n30124 , n46910 );
and ( n47083 , n47081 , n47082 );
xor ( n47084 , n47081 , n47082 );
xor ( n47085 , n46480 , n46820 );
and ( n47086 , n30129 , n46910 );
and ( n47087 , n47085 , n47086 );
xor ( n47088 , n47085 , n47086 );
xor ( n47089 , n46484 , n46818 );
and ( n47090 , n30134 , n46910 );
and ( n47091 , n47089 , n47090 );
xor ( n47092 , n47089 , n47090 );
xor ( n47093 , n46488 , n46816 );
and ( n47094 , n30139 , n46910 );
and ( n47095 , n47093 , n47094 );
xor ( n47096 , n47093 , n47094 );
xor ( n47097 , n46492 , n46814 );
and ( n47098 , n30144 , n46910 );
and ( n47099 , n47097 , n47098 );
xor ( n47100 , n47097 , n47098 );
xor ( n47101 , n46496 , n46812 );
and ( n47102 , n30149 , n46910 );
and ( n47103 , n47101 , n47102 );
xor ( n47104 , n47101 , n47102 );
xor ( n47105 , n46500 , n46810 );
and ( n47106 , n30154 , n46910 );
and ( n47107 , n47105 , n47106 );
xor ( n47108 , n47105 , n47106 );
xor ( n47109 , n46504 , n46808 );
and ( n47110 , n30159 , n46910 );
and ( n47111 , n47109 , n47110 );
xor ( n47112 , n47109 , n47110 );
xor ( n47113 , n46508 , n46806 );
and ( n47114 , n30164 , n46910 );
and ( n47115 , n47113 , n47114 );
xor ( n47116 , n47113 , n47114 );
xor ( n47117 , n46512 , n46804 );
and ( n47118 , n30169 , n46910 );
and ( n47119 , n47117 , n47118 );
xor ( n47120 , n47117 , n47118 );
xor ( n47121 , n46516 , n46802 );
and ( n47122 , n30174 , n46910 );
and ( n47123 , n47121 , n47122 );
xor ( n47124 , n47121 , n47122 );
xor ( n47125 , n46520 , n46800 );
and ( n47126 , n30179 , n46910 );
and ( n47127 , n47125 , n47126 );
xor ( n47128 , n47125 , n47126 );
xor ( n47129 , n46524 , n46798 );
and ( n47130 , n30184 , n46910 );
and ( n47131 , n47129 , n47130 );
xor ( n47132 , n47129 , n47130 );
xor ( n47133 , n46528 , n46796 );
and ( n47134 , n30189 , n46910 );
and ( n47135 , n47133 , n47134 );
xor ( n47136 , n47133 , n47134 );
xor ( n47137 , n46532 , n46794 );
and ( n47138 , n30194 , n46910 );
and ( n47139 , n47137 , n47138 );
xor ( n47140 , n47137 , n47138 );
xor ( n47141 , n46536 , n46792 );
and ( n47142 , n30199 , n46910 );
and ( n47143 , n47141 , n47142 );
xor ( n47144 , n47141 , n47142 );
xor ( n47145 , n46540 , n46790 );
and ( n47146 , n30204 , n46910 );
and ( n47147 , n47145 , n47146 );
xor ( n47148 , n47145 , n47146 );
xor ( n47149 , n46544 , n46788 );
and ( n47150 , n30209 , n46910 );
and ( n47151 , n47149 , n47150 );
xor ( n47152 , n47149 , n47150 );
xor ( n47153 , n46548 , n46786 );
and ( n47154 , n30214 , n46910 );
and ( n47155 , n47153 , n47154 );
xor ( n47156 , n47153 , n47154 );
xor ( n47157 , n46552 , n46784 );
and ( n47158 , n30219 , n46910 );
and ( n47159 , n47157 , n47158 );
xor ( n47160 , n47157 , n47158 );
xor ( n47161 , n46556 , n46782 );
and ( n47162 , n30224 , n46910 );
and ( n47163 , n47161 , n47162 );
xor ( n47164 , n47161 , n47162 );
xor ( n47165 , n46560 , n46780 );
and ( n47166 , n30229 , n46910 );
and ( n47167 , n47165 , n47166 );
xor ( n47168 , n47165 , n47166 );
xor ( n47169 , n46564 , n46778 );
and ( n47170 , n30234 , n46910 );
and ( n47171 , n47169 , n47170 );
xor ( n47172 , n47169 , n47170 );
xor ( n47173 , n46568 , n46776 );
and ( n47174 , n30239 , n46910 );
and ( n47175 , n47173 , n47174 );
xor ( n47176 , n47173 , n47174 );
xor ( n47177 , n46572 , n46774 );
and ( n47178 , n30244 , n46910 );
and ( n47179 , n47177 , n47178 );
xor ( n47180 , n47177 , n47178 );
xor ( n47181 , n46576 , n46772 );
and ( n47182 , n30249 , n46910 );
and ( n47183 , n47181 , n47182 );
xor ( n47184 , n47181 , n47182 );
xor ( n47185 , n46580 , n46770 );
and ( n47186 , n30254 , n46910 );
and ( n47187 , n47185 , n47186 );
xor ( n47188 , n47185 , n47186 );
xor ( n47189 , n46584 , n46768 );
and ( n47190 , n30259 , n46910 );
and ( n47191 , n47189 , n47190 );
xor ( n47192 , n47189 , n47190 );
xor ( n47193 , n46588 , n46766 );
and ( n47194 , n30264 , n46910 );
and ( n47195 , n47193 , n47194 );
xor ( n47196 , n47193 , n47194 );
xor ( n47197 , n46592 , n46764 );
and ( n47198 , n30269 , n46910 );
and ( n47199 , n47197 , n47198 );
xor ( n47200 , n47197 , n47198 );
xor ( n47201 , n46596 , n46762 );
and ( n47202 , n30274 , n46910 );
and ( n47203 , n47201 , n47202 );
xor ( n47204 , n47201 , n47202 );
xor ( n47205 , n46600 , n46760 );
and ( n47206 , n30279 , n46910 );
and ( n47207 , n47205 , n47206 );
xor ( n47208 , n47205 , n47206 );
xor ( n47209 , n46604 , n46758 );
and ( n47210 , n30284 , n46910 );
and ( n47211 , n47209 , n47210 );
xor ( n47212 , n47209 , n47210 );
xor ( n47213 , n46608 , n46756 );
and ( n47214 , n30289 , n46910 );
and ( n47215 , n47213 , n47214 );
xor ( n47216 , n47213 , n47214 );
xor ( n47217 , n46612 , n46754 );
and ( n47218 , n30294 , n46910 );
and ( n47219 , n47217 , n47218 );
xor ( n47220 , n47217 , n47218 );
xor ( n47221 , n46616 , n46752 );
and ( n47222 , n30299 , n46910 );
and ( n47223 , n47221 , n47222 );
xor ( n47224 , n47221 , n47222 );
xor ( n47225 , n46620 , n46750 );
and ( n47226 , n30304 , n46910 );
and ( n47227 , n47225 , n47226 );
xor ( n47228 , n47225 , n47226 );
xor ( n47229 , n46624 , n46748 );
and ( n47230 , n30309 , n46910 );
and ( n47231 , n47229 , n47230 );
xor ( n47232 , n47229 , n47230 );
xor ( n47233 , n46628 , n46746 );
and ( n47234 , n30314 , n46910 );
and ( n47235 , n47233 , n47234 );
xor ( n47236 , n47233 , n47234 );
xor ( n47237 , n46632 , n46744 );
and ( n47238 , n30319 , n46910 );
and ( n47239 , n47237 , n47238 );
xor ( n47240 , n47237 , n47238 );
xor ( n47241 , n46636 , n46742 );
and ( n47242 , n30324 , n46910 );
and ( n47243 , n47241 , n47242 );
xor ( n47244 , n47241 , n47242 );
xor ( n47245 , n46640 , n46740 );
and ( n47246 , n30329 , n46910 );
and ( n47247 , n47245 , n47246 );
xor ( n47248 , n47245 , n47246 );
xor ( n47249 , n46644 , n46738 );
and ( n47250 , n30334 , n46910 );
and ( n47251 , n47249 , n47250 );
xor ( n47252 , n47249 , n47250 );
xor ( n47253 , n46648 , n46736 );
and ( n47254 , n30339 , n46910 );
and ( n47255 , n47253 , n47254 );
xor ( n47256 , n47253 , n47254 );
xor ( n47257 , n46652 , n46734 );
and ( n47258 , n30344 , n46910 );
and ( n47259 , n47257 , n47258 );
xor ( n47260 , n47257 , n47258 );
xor ( n47261 , n46656 , n46732 );
and ( n47262 , n30349 , n46910 );
and ( n47263 , n47261 , n47262 );
xor ( n47264 , n47261 , n47262 );
xor ( n47265 , n46660 , n46730 );
and ( n47266 , n30354 , n46910 );
and ( n47267 , n47265 , n47266 );
xor ( n47268 , n47265 , n47266 );
xor ( n47269 , n46664 , n46728 );
and ( n47270 , n30359 , n46910 );
and ( n47271 , n47269 , n47270 );
xor ( n47272 , n47269 , n47270 );
xor ( n47273 , n46668 , n46726 );
and ( n47274 , n30364 , n46910 );
and ( n47275 , n47273 , n47274 );
xor ( n47276 , n47273 , n47274 );
xor ( n47277 , n46672 , n46724 );
and ( n47278 , n30369 , n46910 );
and ( n47279 , n47277 , n47278 );
xor ( n47280 , n47277 , n47278 );
xor ( n47281 , n46676 , n46722 );
and ( n47282 , n30374 , n46910 );
and ( n47283 , n47281 , n47282 );
xor ( n47284 , n47281 , n47282 );
xor ( n47285 , n46680 , n46720 );
and ( n47286 , n30379 , n46910 );
and ( n47287 , n47285 , n47286 );
xor ( n47288 , n47285 , n47286 );
xor ( n47289 , n46684 , n46718 );
and ( n47290 , n30384 , n46910 );
and ( n47291 , n47289 , n47290 );
xor ( n47292 , n47289 , n47290 );
xor ( n47293 , n46688 , n46716 );
and ( n47294 , n30389 , n46910 );
and ( n47295 , n47293 , n47294 );
xor ( n47296 , n47293 , n47294 );
xor ( n47297 , n46692 , n46714 );
and ( n47298 , n30394 , n46910 );
and ( n47299 , n47297 , n47298 );
xor ( n47300 , n47297 , n47298 );
xor ( n47301 , n46696 , n46712 );
and ( n47302 , n30399 , n46910 );
and ( n47303 , n47301 , n47302 );
xor ( n47304 , n47301 , n47302 );
xor ( n47305 , n46700 , n46710 );
and ( n47306 , n30404 , n46910 );
and ( n47307 , n47305 , n47306 );
xor ( n47308 , n47305 , n47306 );
xor ( n47309 , n46704 , n46708 );
and ( n47310 , n30409 , n46910 );
and ( n47311 , n47309 , n47310 );
buf ( n47312 , n47311 );
and ( n47313 , n47308 , n47312 );
or ( n47314 , n47307 , n47313 );
and ( n47315 , n47304 , n47314 );
or ( n47316 , n47303 , n47315 );
and ( n47317 , n47300 , n47316 );
or ( n47318 , n47299 , n47317 );
and ( n47319 , n47296 , n47318 );
or ( n47320 , n47295 , n47319 );
and ( n47321 , n47292 , n47320 );
or ( n47322 , n47291 , n47321 );
and ( n47323 , n47288 , n47322 );
or ( n47324 , n47287 , n47323 );
and ( n47325 , n47284 , n47324 );
or ( n47326 , n47283 , n47325 );
and ( n47327 , n47280 , n47326 );
or ( n47328 , n47279 , n47327 );
and ( n47329 , n47276 , n47328 );
or ( n47330 , n47275 , n47329 );
and ( n47331 , n47272 , n47330 );
or ( n47332 , n47271 , n47331 );
and ( n47333 , n47268 , n47332 );
or ( n47334 , n47267 , n47333 );
and ( n47335 , n47264 , n47334 );
or ( n47336 , n47263 , n47335 );
and ( n47337 , n47260 , n47336 );
or ( n47338 , n47259 , n47337 );
and ( n47339 , n47256 , n47338 );
or ( n47340 , n47255 , n47339 );
and ( n47341 , n47252 , n47340 );
or ( n47342 , n47251 , n47341 );
and ( n47343 , n47248 , n47342 );
or ( n47344 , n47247 , n47343 );
and ( n47345 , n47244 , n47344 );
or ( n47346 , n47243 , n47345 );
and ( n47347 , n47240 , n47346 );
or ( n47348 , n47239 , n47347 );
and ( n47349 , n47236 , n47348 );
or ( n47350 , n47235 , n47349 );
and ( n47351 , n47232 , n47350 );
or ( n47352 , n47231 , n47351 );
and ( n47353 , n47228 , n47352 );
or ( n47354 , n47227 , n47353 );
and ( n47355 , n47224 , n47354 );
or ( n47356 , n47223 , n47355 );
and ( n47357 , n47220 , n47356 );
or ( n47358 , n47219 , n47357 );
and ( n47359 , n47216 , n47358 );
or ( n47360 , n47215 , n47359 );
and ( n47361 , n47212 , n47360 );
or ( n47362 , n47211 , n47361 );
and ( n47363 , n47208 , n47362 );
or ( n47364 , n47207 , n47363 );
and ( n47365 , n47204 , n47364 );
or ( n47366 , n47203 , n47365 );
and ( n47367 , n47200 , n47366 );
or ( n47368 , n47199 , n47367 );
and ( n47369 , n47196 , n47368 );
or ( n47370 , n47195 , n47369 );
and ( n47371 , n47192 , n47370 );
or ( n47372 , n47191 , n47371 );
and ( n47373 , n47188 , n47372 );
or ( n47374 , n47187 , n47373 );
and ( n47375 , n47184 , n47374 );
or ( n47376 , n47183 , n47375 );
and ( n47377 , n47180 , n47376 );
or ( n47378 , n47179 , n47377 );
and ( n47379 , n47176 , n47378 );
or ( n47380 , n47175 , n47379 );
and ( n47381 , n47172 , n47380 );
or ( n47382 , n47171 , n47381 );
and ( n47383 , n47168 , n47382 );
or ( n47384 , n47167 , n47383 );
and ( n47385 , n47164 , n47384 );
or ( n47386 , n47163 , n47385 );
and ( n47387 , n47160 , n47386 );
or ( n47388 , n47159 , n47387 );
and ( n47389 , n47156 , n47388 );
or ( n47390 , n47155 , n47389 );
and ( n47391 , n47152 , n47390 );
or ( n47392 , n47151 , n47391 );
and ( n47393 , n47148 , n47392 );
or ( n47394 , n47147 , n47393 );
and ( n47395 , n47144 , n47394 );
or ( n47396 , n47143 , n47395 );
and ( n47397 , n47140 , n47396 );
or ( n47398 , n47139 , n47397 );
and ( n47399 , n47136 , n47398 );
or ( n47400 , n47135 , n47399 );
and ( n47401 , n47132 , n47400 );
or ( n47402 , n47131 , n47401 );
and ( n47403 , n47128 , n47402 );
or ( n47404 , n47127 , n47403 );
and ( n47405 , n47124 , n47404 );
or ( n47406 , n47123 , n47405 );
and ( n47407 , n47120 , n47406 );
or ( n47408 , n47119 , n47407 );
and ( n47409 , n47116 , n47408 );
or ( n47410 , n47115 , n47409 );
and ( n47411 , n47112 , n47410 );
or ( n47412 , n47111 , n47411 );
and ( n47413 , n47108 , n47412 );
or ( n47414 , n47107 , n47413 );
and ( n47415 , n47104 , n47414 );
or ( n47416 , n47103 , n47415 );
and ( n47417 , n47100 , n47416 );
or ( n47418 , n47099 , n47417 );
and ( n47419 , n47096 , n47418 );
or ( n47420 , n47095 , n47419 );
and ( n47421 , n47092 , n47420 );
or ( n47422 , n47091 , n47421 );
and ( n47423 , n47088 , n47422 );
or ( n47424 , n47087 , n47423 );
and ( n47425 , n47084 , n47424 );
or ( n47426 , n47083 , n47425 );
and ( n47427 , n47080 , n47426 );
or ( n47428 , n47079 , n47427 );
and ( n47429 , n47076 , n47428 );
or ( n47430 , n47075 , n47429 );
and ( n47431 , n47072 , n47430 );
or ( n47432 , n47071 , n47431 );
and ( n47433 , n47068 , n47432 );
or ( n47434 , n47067 , n47433 );
and ( n47435 , n47064 , n47434 );
or ( n47436 , n47063 , n47435 );
and ( n47437 , n47060 , n47436 );
or ( n47438 , n47059 , n47437 );
and ( n47439 , n47056 , n47438 );
or ( n47440 , n47055 , n47439 );
and ( n47441 , n47052 , n47440 );
or ( n47442 , n47051 , n47441 );
and ( n47443 , n47048 , n47442 );
or ( n47444 , n47047 , n47443 );
and ( n47445 , n47044 , n47444 );
or ( n47446 , n47043 , n47445 );
and ( n47447 , n47040 , n47446 );
or ( n47448 , n47039 , n47447 );
and ( n47449 , n47036 , n47448 );
or ( n47450 , n47035 , n47449 );
and ( n47451 , n47032 , n47450 );
or ( n47452 , n47031 , n47451 );
and ( n47453 , n47028 , n47452 );
or ( n47454 , n47027 , n47453 );
and ( n47455 , n47024 , n47454 );
or ( n47456 , n47023 , n47455 );
and ( n47457 , n47020 , n47456 );
or ( n47458 , n47019 , n47457 );
and ( n47459 , n47016 , n47458 );
or ( n47460 , n47015 , n47459 );
and ( n47461 , n47012 , n47460 );
or ( n47462 , n47011 , n47461 );
and ( n47463 , n47008 , n47462 );
or ( n47464 , n47007 , n47463 );
and ( n47465 , n47004 , n47464 );
or ( n47466 , n47003 , n47465 );
and ( n47467 , n47000 , n47466 );
or ( n47468 , n46999 , n47467 );
and ( n47469 , n46996 , n47468 );
or ( n47470 , n46995 , n47469 );
and ( n47471 , n46992 , n47470 );
or ( n47472 , n46991 , n47471 );
and ( n47473 , n46988 , n47472 );
or ( n47474 , n46987 , n47473 );
and ( n47475 , n46984 , n47474 );
or ( n47476 , n46983 , n47475 );
and ( n47477 , n46980 , n47476 );
or ( n47478 , n46979 , n47477 );
and ( n47479 , n46976 , n47478 );
or ( n47480 , n46975 , n47479 );
and ( n47481 , n46972 , n47480 );
or ( n47482 , n46971 , n47481 );
and ( n47483 , n46968 , n47482 );
or ( n47484 , n46967 , n47483 );
and ( n47485 , n46964 , n47484 );
or ( n47486 , n46963 , n47485 );
and ( n47487 , n46960 , n47486 );
or ( n47488 , n46959 , n47487 );
and ( n47489 , n46956 , n47488 );
or ( n47490 , n46955 , n47489 );
and ( n47491 , n46952 , n47490 );
or ( n47492 , n46951 , n47491 );
and ( n47493 , n46948 , n47492 );
or ( n47494 , n46947 , n47493 );
and ( n47495 , n46944 , n47494 );
or ( n47496 , n46943 , n47495 );
and ( n47497 , n46940 , n47496 );
or ( n47498 , n46939 , n47497 );
and ( n47499 , n46936 , n47498 );
or ( n47500 , n46935 , n47499 );
and ( n47501 , n46932 , n47500 );
or ( n47502 , n46931 , n47501 );
and ( n47503 , n46928 , n47502 );
or ( n47504 , n46927 , n47503 );
and ( n47505 , n46924 , n47504 );
or ( n47506 , n46923 , n47505 );
and ( n47507 , n46920 , n47506 );
or ( n47508 , n46919 , n47507 );
and ( n47509 , n46916 , n47508 );
or ( n47510 , n46915 , n47509 );
xor ( n47511 , n46912 , n47510 );
buf ( n47512 , n18052 );
and ( n47513 , n29914 , n47512 );
xor ( n47514 , n47511 , n47513 );
xor ( n47515 , n46916 , n47508 );
and ( n47516 , n29919 , n47512 );
and ( n47517 , n47515 , n47516 );
xor ( n47518 , n47515 , n47516 );
xor ( n47519 , n46920 , n47506 );
and ( n47520 , n29924 , n47512 );
and ( n47521 , n47519 , n47520 );
xor ( n47522 , n47519 , n47520 );
xor ( n47523 , n46924 , n47504 );
and ( n47524 , n29929 , n47512 );
and ( n47525 , n47523 , n47524 );
xor ( n47526 , n47523 , n47524 );
xor ( n47527 , n46928 , n47502 );
and ( n47528 , n29934 , n47512 );
and ( n47529 , n47527 , n47528 );
xor ( n47530 , n47527 , n47528 );
xor ( n47531 , n46932 , n47500 );
and ( n47532 , n29939 , n47512 );
and ( n47533 , n47531 , n47532 );
xor ( n47534 , n47531 , n47532 );
xor ( n47535 , n46936 , n47498 );
and ( n47536 , n29944 , n47512 );
and ( n47537 , n47535 , n47536 );
xor ( n47538 , n47535 , n47536 );
xor ( n47539 , n46940 , n47496 );
and ( n47540 , n29949 , n47512 );
and ( n47541 , n47539 , n47540 );
xor ( n47542 , n47539 , n47540 );
xor ( n47543 , n46944 , n47494 );
and ( n47544 , n29954 , n47512 );
and ( n47545 , n47543 , n47544 );
xor ( n47546 , n47543 , n47544 );
xor ( n47547 , n46948 , n47492 );
and ( n47548 , n29959 , n47512 );
and ( n47549 , n47547 , n47548 );
xor ( n47550 , n47547 , n47548 );
xor ( n47551 , n46952 , n47490 );
and ( n47552 , n29964 , n47512 );
and ( n47553 , n47551 , n47552 );
xor ( n47554 , n47551 , n47552 );
xor ( n47555 , n46956 , n47488 );
and ( n47556 , n29969 , n47512 );
and ( n47557 , n47555 , n47556 );
xor ( n47558 , n47555 , n47556 );
xor ( n47559 , n46960 , n47486 );
and ( n47560 , n29974 , n47512 );
and ( n47561 , n47559 , n47560 );
xor ( n47562 , n47559 , n47560 );
xor ( n47563 , n46964 , n47484 );
and ( n47564 , n29979 , n47512 );
and ( n47565 , n47563 , n47564 );
xor ( n47566 , n47563 , n47564 );
xor ( n47567 , n46968 , n47482 );
and ( n47568 , n29984 , n47512 );
and ( n47569 , n47567 , n47568 );
xor ( n47570 , n47567 , n47568 );
xor ( n47571 , n46972 , n47480 );
and ( n47572 , n29989 , n47512 );
and ( n47573 , n47571 , n47572 );
xor ( n47574 , n47571 , n47572 );
xor ( n47575 , n46976 , n47478 );
and ( n47576 , n29994 , n47512 );
and ( n47577 , n47575 , n47576 );
xor ( n47578 , n47575 , n47576 );
xor ( n47579 , n46980 , n47476 );
and ( n47580 , n29999 , n47512 );
and ( n47581 , n47579 , n47580 );
xor ( n47582 , n47579 , n47580 );
xor ( n47583 , n46984 , n47474 );
and ( n47584 , n30004 , n47512 );
and ( n47585 , n47583 , n47584 );
xor ( n47586 , n47583 , n47584 );
xor ( n47587 , n46988 , n47472 );
and ( n47588 , n30009 , n47512 );
and ( n47589 , n47587 , n47588 );
xor ( n47590 , n47587 , n47588 );
xor ( n47591 , n46992 , n47470 );
and ( n47592 , n30014 , n47512 );
and ( n47593 , n47591 , n47592 );
xor ( n47594 , n47591 , n47592 );
xor ( n47595 , n46996 , n47468 );
and ( n47596 , n30019 , n47512 );
and ( n47597 , n47595 , n47596 );
xor ( n47598 , n47595 , n47596 );
xor ( n47599 , n47000 , n47466 );
and ( n47600 , n30024 , n47512 );
and ( n47601 , n47599 , n47600 );
xor ( n47602 , n47599 , n47600 );
xor ( n47603 , n47004 , n47464 );
and ( n47604 , n30029 , n47512 );
and ( n47605 , n47603 , n47604 );
xor ( n47606 , n47603 , n47604 );
xor ( n47607 , n47008 , n47462 );
and ( n47608 , n30034 , n47512 );
and ( n47609 , n47607 , n47608 );
xor ( n47610 , n47607 , n47608 );
xor ( n47611 , n47012 , n47460 );
and ( n47612 , n30039 , n47512 );
and ( n47613 , n47611 , n47612 );
xor ( n47614 , n47611 , n47612 );
xor ( n47615 , n47016 , n47458 );
and ( n47616 , n30044 , n47512 );
and ( n47617 , n47615 , n47616 );
xor ( n47618 , n47615 , n47616 );
xor ( n47619 , n47020 , n47456 );
and ( n47620 , n30049 , n47512 );
and ( n47621 , n47619 , n47620 );
xor ( n47622 , n47619 , n47620 );
xor ( n47623 , n47024 , n47454 );
and ( n47624 , n30054 , n47512 );
and ( n47625 , n47623 , n47624 );
xor ( n47626 , n47623 , n47624 );
xor ( n47627 , n47028 , n47452 );
and ( n47628 , n30059 , n47512 );
and ( n47629 , n47627 , n47628 );
xor ( n47630 , n47627 , n47628 );
xor ( n47631 , n47032 , n47450 );
and ( n47632 , n30064 , n47512 );
and ( n47633 , n47631 , n47632 );
xor ( n47634 , n47631 , n47632 );
xor ( n47635 , n47036 , n47448 );
and ( n47636 , n30069 , n47512 );
and ( n47637 , n47635 , n47636 );
xor ( n47638 , n47635 , n47636 );
xor ( n47639 , n47040 , n47446 );
and ( n47640 , n30074 , n47512 );
and ( n47641 , n47639 , n47640 );
xor ( n47642 , n47639 , n47640 );
xor ( n47643 , n47044 , n47444 );
and ( n47644 , n30079 , n47512 );
and ( n47645 , n47643 , n47644 );
xor ( n47646 , n47643 , n47644 );
xor ( n47647 , n47048 , n47442 );
and ( n47648 , n30084 , n47512 );
and ( n47649 , n47647 , n47648 );
xor ( n47650 , n47647 , n47648 );
xor ( n47651 , n47052 , n47440 );
and ( n47652 , n30089 , n47512 );
and ( n47653 , n47651 , n47652 );
xor ( n47654 , n47651 , n47652 );
xor ( n47655 , n47056 , n47438 );
and ( n47656 , n30094 , n47512 );
and ( n47657 , n47655 , n47656 );
xor ( n47658 , n47655 , n47656 );
xor ( n47659 , n47060 , n47436 );
and ( n47660 , n30099 , n47512 );
and ( n47661 , n47659 , n47660 );
xor ( n47662 , n47659 , n47660 );
xor ( n47663 , n47064 , n47434 );
and ( n47664 , n30104 , n47512 );
and ( n47665 , n47663 , n47664 );
xor ( n47666 , n47663 , n47664 );
xor ( n47667 , n47068 , n47432 );
and ( n47668 , n30109 , n47512 );
and ( n47669 , n47667 , n47668 );
xor ( n47670 , n47667 , n47668 );
xor ( n47671 , n47072 , n47430 );
and ( n47672 , n30114 , n47512 );
and ( n47673 , n47671 , n47672 );
xor ( n47674 , n47671 , n47672 );
xor ( n47675 , n47076 , n47428 );
and ( n47676 , n30119 , n47512 );
and ( n47677 , n47675 , n47676 );
xor ( n47678 , n47675 , n47676 );
xor ( n47679 , n47080 , n47426 );
and ( n47680 , n30124 , n47512 );
and ( n47681 , n47679 , n47680 );
xor ( n47682 , n47679 , n47680 );
xor ( n47683 , n47084 , n47424 );
and ( n47684 , n30129 , n47512 );
and ( n47685 , n47683 , n47684 );
xor ( n47686 , n47683 , n47684 );
xor ( n47687 , n47088 , n47422 );
and ( n47688 , n30134 , n47512 );
and ( n47689 , n47687 , n47688 );
xor ( n47690 , n47687 , n47688 );
xor ( n47691 , n47092 , n47420 );
and ( n47692 , n30139 , n47512 );
and ( n47693 , n47691 , n47692 );
xor ( n47694 , n47691 , n47692 );
xor ( n47695 , n47096 , n47418 );
and ( n47696 , n30144 , n47512 );
and ( n47697 , n47695 , n47696 );
xor ( n47698 , n47695 , n47696 );
xor ( n47699 , n47100 , n47416 );
and ( n47700 , n30149 , n47512 );
and ( n47701 , n47699 , n47700 );
xor ( n47702 , n47699 , n47700 );
xor ( n47703 , n47104 , n47414 );
and ( n47704 , n30154 , n47512 );
and ( n47705 , n47703 , n47704 );
xor ( n47706 , n47703 , n47704 );
xor ( n47707 , n47108 , n47412 );
and ( n47708 , n30159 , n47512 );
and ( n47709 , n47707 , n47708 );
xor ( n47710 , n47707 , n47708 );
xor ( n47711 , n47112 , n47410 );
and ( n47712 , n30164 , n47512 );
and ( n47713 , n47711 , n47712 );
xor ( n47714 , n47711 , n47712 );
xor ( n47715 , n47116 , n47408 );
and ( n47716 , n30169 , n47512 );
and ( n47717 , n47715 , n47716 );
xor ( n47718 , n47715 , n47716 );
xor ( n47719 , n47120 , n47406 );
and ( n47720 , n30174 , n47512 );
and ( n47721 , n47719 , n47720 );
xor ( n47722 , n47719 , n47720 );
xor ( n47723 , n47124 , n47404 );
and ( n47724 , n30179 , n47512 );
and ( n47725 , n47723 , n47724 );
xor ( n47726 , n47723 , n47724 );
xor ( n47727 , n47128 , n47402 );
and ( n47728 , n30184 , n47512 );
and ( n47729 , n47727 , n47728 );
xor ( n47730 , n47727 , n47728 );
xor ( n47731 , n47132 , n47400 );
and ( n47732 , n30189 , n47512 );
and ( n47733 , n47731 , n47732 );
xor ( n47734 , n47731 , n47732 );
xor ( n47735 , n47136 , n47398 );
and ( n47736 , n30194 , n47512 );
and ( n47737 , n47735 , n47736 );
xor ( n47738 , n47735 , n47736 );
xor ( n47739 , n47140 , n47396 );
and ( n47740 , n30199 , n47512 );
and ( n47741 , n47739 , n47740 );
xor ( n47742 , n47739 , n47740 );
xor ( n47743 , n47144 , n47394 );
and ( n47744 , n30204 , n47512 );
and ( n47745 , n47743 , n47744 );
xor ( n47746 , n47743 , n47744 );
xor ( n47747 , n47148 , n47392 );
and ( n47748 , n30209 , n47512 );
and ( n47749 , n47747 , n47748 );
xor ( n47750 , n47747 , n47748 );
xor ( n47751 , n47152 , n47390 );
and ( n47752 , n30214 , n47512 );
and ( n47753 , n47751 , n47752 );
xor ( n47754 , n47751 , n47752 );
xor ( n47755 , n47156 , n47388 );
and ( n47756 , n30219 , n47512 );
and ( n47757 , n47755 , n47756 );
xor ( n47758 , n47755 , n47756 );
xor ( n47759 , n47160 , n47386 );
and ( n47760 , n30224 , n47512 );
and ( n47761 , n47759 , n47760 );
xor ( n47762 , n47759 , n47760 );
xor ( n47763 , n47164 , n47384 );
and ( n47764 , n30229 , n47512 );
and ( n47765 , n47763 , n47764 );
xor ( n47766 , n47763 , n47764 );
xor ( n47767 , n47168 , n47382 );
and ( n47768 , n30234 , n47512 );
and ( n47769 , n47767 , n47768 );
xor ( n47770 , n47767 , n47768 );
xor ( n47771 , n47172 , n47380 );
and ( n47772 , n30239 , n47512 );
and ( n47773 , n47771 , n47772 );
xor ( n47774 , n47771 , n47772 );
xor ( n47775 , n47176 , n47378 );
and ( n47776 , n30244 , n47512 );
and ( n47777 , n47775 , n47776 );
xor ( n47778 , n47775 , n47776 );
xor ( n47779 , n47180 , n47376 );
and ( n47780 , n30249 , n47512 );
and ( n47781 , n47779 , n47780 );
xor ( n47782 , n47779 , n47780 );
xor ( n47783 , n47184 , n47374 );
and ( n47784 , n30254 , n47512 );
and ( n47785 , n47783 , n47784 );
xor ( n47786 , n47783 , n47784 );
xor ( n47787 , n47188 , n47372 );
and ( n47788 , n30259 , n47512 );
and ( n47789 , n47787 , n47788 );
xor ( n47790 , n47787 , n47788 );
xor ( n47791 , n47192 , n47370 );
and ( n47792 , n30264 , n47512 );
and ( n47793 , n47791 , n47792 );
xor ( n47794 , n47791 , n47792 );
xor ( n47795 , n47196 , n47368 );
and ( n47796 , n30269 , n47512 );
and ( n47797 , n47795 , n47796 );
xor ( n47798 , n47795 , n47796 );
xor ( n47799 , n47200 , n47366 );
and ( n47800 , n30274 , n47512 );
and ( n47801 , n47799 , n47800 );
xor ( n47802 , n47799 , n47800 );
xor ( n47803 , n47204 , n47364 );
and ( n47804 , n30279 , n47512 );
and ( n47805 , n47803 , n47804 );
xor ( n47806 , n47803 , n47804 );
xor ( n47807 , n47208 , n47362 );
and ( n47808 , n30284 , n47512 );
and ( n47809 , n47807 , n47808 );
xor ( n47810 , n47807 , n47808 );
xor ( n47811 , n47212 , n47360 );
and ( n47812 , n30289 , n47512 );
and ( n47813 , n47811 , n47812 );
xor ( n47814 , n47811 , n47812 );
xor ( n47815 , n47216 , n47358 );
and ( n47816 , n30294 , n47512 );
and ( n47817 , n47815 , n47816 );
xor ( n47818 , n47815 , n47816 );
xor ( n47819 , n47220 , n47356 );
and ( n47820 , n30299 , n47512 );
and ( n47821 , n47819 , n47820 );
xor ( n47822 , n47819 , n47820 );
xor ( n47823 , n47224 , n47354 );
and ( n47824 , n30304 , n47512 );
and ( n47825 , n47823 , n47824 );
xor ( n47826 , n47823 , n47824 );
xor ( n47827 , n47228 , n47352 );
and ( n47828 , n30309 , n47512 );
and ( n47829 , n47827 , n47828 );
xor ( n47830 , n47827 , n47828 );
xor ( n47831 , n47232 , n47350 );
and ( n47832 , n30314 , n47512 );
and ( n47833 , n47831 , n47832 );
xor ( n47834 , n47831 , n47832 );
xor ( n47835 , n47236 , n47348 );
and ( n47836 , n30319 , n47512 );
and ( n47837 , n47835 , n47836 );
xor ( n47838 , n47835 , n47836 );
xor ( n47839 , n47240 , n47346 );
and ( n47840 , n30324 , n47512 );
and ( n47841 , n47839 , n47840 );
xor ( n47842 , n47839 , n47840 );
xor ( n47843 , n47244 , n47344 );
and ( n47844 , n30329 , n47512 );
and ( n47845 , n47843 , n47844 );
xor ( n47846 , n47843 , n47844 );
xor ( n47847 , n47248 , n47342 );
and ( n47848 , n30334 , n47512 );
and ( n47849 , n47847 , n47848 );
xor ( n47850 , n47847 , n47848 );
xor ( n47851 , n47252 , n47340 );
and ( n47852 , n30339 , n47512 );
and ( n47853 , n47851 , n47852 );
xor ( n47854 , n47851 , n47852 );
xor ( n47855 , n47256 , n47338 );
and ( n47856 , n30344 , n47512 );
and ( n47857 , n47855 , n47856 );
xor ( n47858 , n47855 , n47856 );
xor ( n47859 , n47260 , n47336 );
and ( n47860 , n30349 , n47512 );
and ( n47861 , n47859 , n47860 );
xor ( n47862 , n47859 , n47860 );
xor ( n47863 , n47264 , n47334 );
and ( n47864 , n30354 , n47512 );
and ( n47865 , n47863 , n47864 );
xor ( n47866 , n47863 , n47864 );
xor ( n47867 , n47268 , n47332 );
and ( n47868 , n30359 , n47512 );
and ( n47869 , n47867 , n47868 );
xor ( n47870 , n47867 , n47868 );
xor ( n47871 , n47272 , n47330 );
and ( n47872 , n30364 , n47512 );
and ( n47873 , n47871 , n47872 );
xor ( n47874 , n47871 , n47872 );
xor ( n47875 , n47276 , n47328 );
and ( n47876 , n30369 , n47512 );
and ( n47877 , n47875 , n47876 );
xor ( n47878 , n47875 , n47876 );
xor ( n47879 , n47280 , n47326 );
and ( n47880 , n30374 , n47512 );
and ( n47881 , n47879 , n47880 );
xor ( n47882 , n47879 , n47880 );
xor ( n47883 , n47284 , n47324 );
and ( n47884 , n30379 , n47512 );
and ( n47885 , n47883 , n47884 );
xor ( n47886 , n47883 , n47884 );
xor ( n47887 , n47288 , n47322 );
and ( n47888 , n30384 , n47512 );
and ( n47889 , n47887 , n47888 );
xor ( n47890 , n47887 , n47888 );
xor ( n47891 , n47292 , n47320 );
and ( n47892 , n30389 , n47512 );
and ( n47893 , n47891 , n47892 );
xor ( n47894 , n47891 , n47892 );
xor ( n47895 , n47296 , n47318 );
and ( n47896 , n30394 , n47512 );
and ( n47897 , n47895 , n47896 );
xor ( n47898 , n47895 , n47896 );
xor ( n47899 , n47300 , n47316 );
and ( n47900 , n30399 , n47512 );
and ( n47901 , n47899 , n47900 );
xor ( n47902 , n47899 , n47900 );
xor ( n47903 , n47304 , n47314 );
and ( n47904 , n30404 , n47512 );
and ( n47905 , n47903 , n47904 );
xor ( n47906 , n47903 , n47904 );
xor ( n47907 , n47308 , n47312 );
and ( n47908 , n30409 , n47512 );
and ( n47909 , n47907 , n47908 );
buf ( n47910 , n47909 );
and ( n47911 , n47906 , n47910 );
or ( n47912 , n47905 , n47911 );
and ( n47913 , n47902 , n47912 );
or ( n47914 , n47901 , n47913 );
and ( n47915 , n47898 , n47914 );
or ( n47916 , n47897 , n47915 );
and ( n47917 , n47894 , n47916 );
or ( n47918 , n47893 , n47917 );
and ( n47919 , n47890 , n47918 );
or ( n47920 , n47889 , n47919 );
and ( n47921 , n47886 , n47920 );
or ( n47922 , n47885 , n47921 );
and ( n47923 , n47882 , n47922 );
or ( n47924 , n47881 , n47923 );
and ( n47925 , n47878 , n47924 );
or ( n47926 , n47877 , n47925 );
and ( n47927 , n47874 , n47926 );
or ( n47928 , n47873 , n47927 );
and ( n47929 , n47870 , n47928 );
or ( n47930 , n47869 , n47929 );
and ( n47931 , n47866 , n47930 );
or ( n47932 , n47865 , n47931 );
and ( n47933 , n47862 , n47932 );
or ( n47934 , n47861 , n47933 );
and ( n47935 , n47858 , n47934 );
or ( n47936 , n47857 , n47935 );
and ( n47937 , n47854 , n47936 );
or ( n47938 , n47853 , n47937 );
and ( n47939 , n47850 , n47938 );
or ( n47940 , n47849 , n47939 );
and ( n47941 , n47846 , n47940 );
or ( n47942 , n47845 , n47941 );
and ( n47943 , n47842 , n47942 );
or ( n47944 , n47841 , n47943 );
and ( n47945 , n47838 , n47944 );
or ( n47946 , n47837 , n47945 );
and ( n47947 , n47834 , n47946 );
or ( n47948 , n47833 , n47947 );
and ( n47949 , n47830 , n47948 );
or ( n47950 , n47829 , n47949 );
and ( n47951 , n47826 , n47950 );
or ( n47952 , n47825 , n47951 );
and ( n47953 , n47822 , n47952 );
or ( n47954 , n47821 , n47953 );
and ( n47955 , n47818 , n47954 );
or ( n47956 , n47817 , n47955 );
and ( n47957 , n47814 , n47956 );
or ( n47958 , n47813 , n47957 );
and ( n47959 , n47810 , n47958 );
or ( n47960 , n47809 , n47959 );
and ( n47961 , n47806 , n47960 );
or ( n47962 , n47805 , n47961 );
and ( n47963 , n47802 , n47962 );
or ( n47964 , n47801 , n47963 );
and ( n47965 , n47798 , n47964 );
or ( n47966 , n47797 , n47965 );
and ( n47967 , n47794 , n47966 );
or ( n47968 , n47793 , n47967 );
and ( n47969 , n47790 , n47968 );
or ( n47970 , n47789 , n47969 );
and ( n47971 , n47786 , n47970 );
or ( n47972 , n47785 , n47971 );
and ( n47973 , n47782 , n47972 );
or ( n47974 , n47781 , n47973 );
and ( n47975 , n47778 , n47974 );
or ( n47976 , n47777 , n47975 );
and ( n47977 , n47774 , n47976 );
or ( n47978 , n47773 , n47977 );
and ( n47979 , n47770 , n47978 );
or ( n47980 , n47769 , n47979 );
and ( n47981 , n47766 , n47980 );
or ( n47982 , n47765 , n47981 );
and ( n47983 , n47762 , n47982 );
or ( n47984 , n47761 , n47983 );
and ( n47985 , n47758 , n47984 );
or ( n47986 , n47757 , n47985 );
and ( n47987 , n47754 , n47986 );
or ( n47988 , n47753 , n47987 );
and ( n47989 , n47750 , n47988 );
or ( n47990 , n47749 , n47989 );
and ( n47991 , n47746 , n47990 );
or ( n47992 , n47745 , n47991 );
and ( n47993 , n47742 , n47992 );
or ( n47994 , n47741 , n47993 );
and ( n47995 , n47738 , n47994 );
or ( n47996 , n47737 , n47995 );
and ( n47997 , n47734 , n47996 );
or ( n47998 , n47733 , n47997 );
and ( n47999 , n47730 , n47998 );
or ( n48000 , n47729 , n47999 );
and ( n48001 , n47726 , n48000 );
or ( n48002 , n47725 , n48001 );
and ( n48003 , n47722 , n48002 );
or ( n48004 , n47721 , n48003 );
and ( n48005 , n47718 , n48004 );
or ( n48006 , n47717 , n48005 );
and ( n48007 , n47714 , n48006 );
or ( n48008 , n47713 , n48007 );
and ( n48009 , n47710 , n48008 );
or ( n48010 , n47709 , n48009 );
and ( n48011 , n47706 , n48010 );
or ( n48012 , n47705 , n48011 );
and ( n48013 , n47702 , n48012 );
or ( n48014 , n47701 , n48013 );
and ( n48015 , n47698 , n48014 );
or ( n48016 , n47697 , n48015 );
and ( n48017 , n47694 , n48016 );
or ( n48018 , n47693 , n48017 );
and ( n48019 , n47690 , n48018 );
or ( n48020 , n47689 , n48019 );
and ( n48021 , n47686 , n48020 );
or ( n48022 , n47685 , n48021 );
and ( n48023 , n47682 , n48022 );
or ( n48024 , n47681 , n48023 );
and ( n48025 , n47678 , n48024 );
or ( n48026 , n47677 , n48025 );
and ( n48027 , n47674 , n48026 );
or ( n48028 , n47673 , n48027 );
and ( n48029 , n47670 , n48028 );
or ( n48030 , n47669 , n48029 );
and ( n48031 , n47666 , n48030 );
or ( n48032 , n47665 , n48031 );
and ( n48033 , n47662 , n48032 );
or ( n48034 , n47661 , n48033 );
and ( n48035 , n47658 , n48034 );
or ( n48036 , n47657 , n48035 );
and ( n48037 , n47654 , n48036 );
or ( n48038 , n47653 , n48037 );
and ( n48039 , n47650 , n48038 );
or ( n48040 , n47649 , n48039 );
and ( n48041 , n47646 , n48040 );
or ( n48042 , n47645 , n48041 );
and ( n48043 , n47642 , n48042 );
or ( n48044 , n47641 , n48043 );
and ( n48045 , n47638 , n48044 );
or ( n48046 , n47637 , n48045 );
and ( n48047 , n47634 , n48046 );
or ( n48048 , n47633 , n48047 );
and ( n48049 , n47630 , n48048 );
or ( n48050 , n47629 , n48049 );
and ( n48051 , n47626 , n48050 );
or ( n48052 , n47625 , n48051 );
and ( n48053 , n47622 , n48052 );
or ( n48054 , n47621 , n48053 );
and ( n48055 , n47618 , n48054 );
or ( n48056 , n47617 , n48055 );
and ( n48057 , n47614 , n48056 );
or ( n48058 , n47613 , n48057 );
and ( n48059 , n47610 , n48058 );
or ( n48060 , n47609 , n48059 );
and ( n48061 , n47606 , n48060 );
or ( n48062 , n47605 , n48061 );
and ( n48063 , n47602 , n48062 );
or ( n48064 , n47601 , n48063 );
and ( n48065 , n47598 , n48064 );
or ( n48066 , n47597 , n48065 );
and ( n48067 , n47594 , n48066 );
or ( n48068 , n47593 , n48067 );
and ( n48069 , n47590 , n48068 );
or ( n48070 , n47589 , n48069 );
and ( n48071 , n47586 , n48070 );
or ( n48072 , n47585 , n48071 );
and ( n48073 , n47582 , n48072 );
or ( n48074 , n47581 , n48073 );
and ( n48075 , n47578 , n48074 );
or ( n48076 , n47577 , n48075 );
and ( n48077 , n47574 , n48076 );
or ( n48078 , n47573 , n48077 );
and ( n48079 , n47570 , n48078 );
or ( n48080 , n47569 , n48079 );
and ( n48081 , n47566 , n48080 );
or ( n48082 , n47565 , n48081 );
and ( n48083 , n47562 , n48082 );
or ( n48084 , n47561 , n48083 );
and ( n48085 , n47558 , n48084 );
or ( n48086 , n47557 , n48085 );
and ( n48087 , n47554 , n48086 );
or ( n48088 , n47553 , n48087 );
and ( n48089 , n47550 , n48088 );
or ( n48090 , n47549 , n48089 );
and ( n48091 , n47546 , n48090 );
or ( n48092 , n47545 , n48091 );
and ( n48093 , n47542 , n48092 );
or ( n48094 , n47541 , n48093 );
and ( n48095 , n47538 , n48094 );
or ( n48096 , n47537 , n48095 );
and ( n48097 , n47534 , n48096 );
or ( n48098 , n47533 , n48097 );
and ( n48099 , n47530 , n48098 );
or ( n48100 , n47529 , n48099 );
and ( n48101 , n47526 , n48100 );
or ( n48102 , n47525 , n48101 );
and ( n48103 , n47522 , n48102 );
or ( n48104 , n47521 , n48103 );
and ( n48105 , n47518 , n48104 );
or ( n48106 , n47517 , n48105 );
xor ( n48107 , n47514 , n48106 );
buf ( n48108 , n18050 );
and ( n48109 , n29919 , n48108 );
xor ( n48110 , n48107 , n48109 );
xor ( n48111 , n47518 , n48104 );
and ( n48112 , n29924 , n48108 );
and ( n48113 , n48111 , n48112 );
xor ( n48114 , n48111 , n48112 );
xor ( n48115 , n47522 , n48102 );
and ( n48116 , n29929 , n48108 );
and ( n48117 , n48115 , n48116 );
xor ( n48118 , n48115 , n48116 );
xor ( n48119 , n47526 , n48100 );
and ( n48120 , n29934 , n48108 );
and ( n48121 , n48119 , n48120 );
xor ( n48122 , n48119 , n48120 );
xor ( n48123 , n47530 , n48098 );
and ( n48124 , n29939 , n48108 );
and ( n48125 , n48123 , n48124 );
xor ( n48126 , n48123 , n48124 );
xor ( n48127 , n47534 , n48096 );
and ( n48128 , n29944 , n48108 );
and ( n48129 , n48127 , n48128 );
xor ( n48130 , n48127 , n48128 );
xor ( n48131 , n47538 , n48094 );
and ( n48132 , n29949 , n48108 );
and ( n48133 , n48131 , n48132 );
xor ( n48134 , n48131 , n48132 );
xor ( n48135 , n47542 , n48092 );
and ( n48136 , n29954 , n48108 );
and ( n48137 , n48135 , n48136 );
xor ( n48138 , n48135 , n48136 );
xor ( n48139 , n47546 , n48090 );
and ( n48140 , n29959 , n48108 );
and ( n48141 , n48139 , n48140 );
xor ( n48142 , n48139 , n48140 );
xor ( n48143 , n47550 , n48088 );
and ( n48144 , n29964 , n48108 );
and ( n48145 , n48143 , n48144 );
xor ( n48146 , n48143 , n48144 );
xor ( n48147 , n47554 , n48086 );
and ( n48148 , n29969 , n48108 );
and ( n48149 , n48147 , n48148 );
xor ( n48150 , n48147 , n48148 );
xor ( n48151 , n47558 , n48084 );
and ( n48152 , n29974 , n48108 );
and ( n48153 , n48151 , n48152 );
xor ( n48154 , n48151 , n48152 );
xor ( n48155 , n47562 , n48082 );
and ( n48156 , n29979 , n48108 );
and ( n48157 , n48155 , n48156 );
xor ( n48158 , n48155 , n48156 );
xor ( n48159 , n47566 , n48080 );
and ( n48160 , n29984 , n48108 );
and ( n48161 , n48159 , n48160 );
xor ( n48162 , n48159 , n48160 );
xor ( n48163 , n47570 , n48078 );
and ( n48164 , n29989 , n48108 );
and ( n48165 , n48163 , n48164 );
xor ( n48166 , n48163 , n48164 );
xor ( n48167 , n47574 , n48076 );
and ( n48168 , n29994 , n48108 );
and ( n48169 , n48167 , n48168 );
xor ( n48170 , n48167 , n48168 );
xor ( n48171 , n47578 , n48074 );
and ( n48172 , n29999 , n48108 );
and ( n48173 , n48171 , n48172 );
xor ( n48174 , n48171 , n48172 );
xor ( n48175 , n47582 , n48072 );
and ( n48176 , n30004 , n48108 );
and ( n48177 , n48175 , n48176 );
xor ( n48178 , n48175 , n48176 );
xor ( n48179 , n47586 , n48070 );
and ( n48180 , n30009 , n48108 );
and ( n48181 , n48179 , n48180 );
xor ( n48182 , n48179 , n48180 );
xor ( n48183 , n47590 , n48068 );
and ( n48184 , n30014 , n48108 );
and ( n48185 , n48183 , n48184 );
xor ( n48186 , n48183 , n48184 );
xor ( n48187 , n47594 , n48066 );
and ( n48188 , n30019 , n48108 );
and ( n48189 , n48187 , n48188 );
xor ( n48190 , n48187 , n48188 );
xor ( n48191 , n47598 , n48064 );
and ( n48192 , n30024 , n48108 );
and ( n48193 , n48191 , n48192 );
xor ( n48194 , n48191 , n48192 );
xor ( n48195 , n47602 , n48062 );
and ( n48196 , n30029 , n48108 );
and ( n48197 , n48195 , n48196 );
xor ( n48198 , n48195 , n48196 );
xor ( n48199 , n47606 , n48060 );
and ( n48200 , n30034 , n48108 );
and ( n48201 , n48199 , n48200 );
xor ( n48202 , n48199 , n48200 );
xor ( n48203 , n47610 , n48058 );
and ( n48204 , n30039 , n48108 );
and ( n48205 , n48203 , n48204 );
xor ( n48206 , n48203 , n48204 );
xor ( n48207 , n47614 , n48056 );
and ( n48208 , n30044 , n48108 );
and ( n48209 , n48207 , n48208 );
xor ( n48210 , n48207 , n48208 );
xor ( n48211 , n47618 , n48054 );
and ( n48212 , n30049 , n48108 );
and ( n48213 , n48211 , n48212 );
xor ( n48214 , n48211 , n48212 );
xor ( n48215 , n47622 , n48052 );
and ( n48216 , n30054 , n48108 );
and ( n48217 , n48215 , n48216 );
xor ( n48218 , n48215 , n48216 );
xor ( n48219 , n47626 , n48050 );
and ( n48220 , n30059 , n48108 );
and ( n48221 , n48219 , n48220 );
xor ( n48222 , n48219 , n48220 );
xor ( n48223 , n47630 , n48048 );
and ( n48224 , n30064 , n48108 );
and ( n48225 , n48223 , n48224 );
xor ( n48226 , n48223 , n48224 );
xor ( n48227 , n47634 , n48046 );
and ( n48228 , n30069 , n48108 );
and ( n48229 , n48227 , n48228 );
xor ( n48230 , n48227 , n48228 );
xor ( n48231 , n47638 , n48044 );
and ( n48232 , n30074 , n48108 );
and ( n48233 , n48231 , n48232 );
xor ( n48234 , n48231 , n48232 );
xor ( n48235 , n47642 , n48042 );
and ( n48236 , n30079 , n48108 );
and ( n48237 , n48235 , n48236 );
xor ( n48238 , n48235 , n48236 );
xor ( n48239 , n47646 , n48040 );
and ( n48240 , n30084 , n48108 );
and ( n48241 , n48239 , n48240 );
xor ( n48242 , n48239 , n48240 );
xor ( n48243 , n47650 , n48038 );
and ( n48244 , n30089 , n48108 );
and ( n48245 , n48243 , n48244 );
xor ( n48246 , n48243 , n48244 );
xor ( n48247 , n47654 , n48036 );
and ( n48248 , n30094 , n48108 );
and ( n48249 , n48247 , n48248 );
xor ( n48250 , n48247 , n48248 );
xor ( n48251 , n47658 , n48034 );
and ( n48252 , n30099 , n48108 );
and ( n48253 , n48251 , n48252 );
xor ( n48254 , n48251 , n48252 );
xor ( n48255 , n47662 , n48032 );
and ( n48256 , n30104 , n48108 );
and ( n48257 , n48255 , n48256 );
xor ( n48258 , n48255 , n48256 );
xor ( n48259 , n47666 , n48030 );
and ( n48260 , n30109 , n48108 );
and ( n48261 , n48259 , n48260 );
xor ( n48262 , n48259 , n48260 );
xor ( n48263 , n47670 , n48028 );
and ( n48264 , n30114 , n48108 );
and ( n48265 , n48263 , n48264 );
xor ( n48266 , n48263 , n48264 );
xor ( n48267 , n47674 , n48026 );
and ( n48268 , n30119 , n48108 );
and ( n48269 , n48267 , n48268 );
xor ( n48270 , n48267 , n48268 );
xor ( n48271 , n47678 , n48024 );
and ( n48272 , n30124 , n48108 );
and ( n48273 , n48271 , n48272 );
xor ( n48274 , n48271 , n48272 );
xor ( n48275 , n47682 , n48022 );
and ( n48276 , n30129 , n48108 );
and ( n48277 , n48275 , n48276 );
xor ( n48278 , n48275 , n48276 );
xor ( n48279 , n47686 , n48020 );
and ( n48280 , n30134 , n48108 );
and ( n48281 , n48279 , n48280 );
xor ( n48282 , n48279 , n48280 );
xor ( n48283 , n47690 , n48018 );
and ( n48284 , n30139 , n48108 );
and ( n48285 , n48283 , n48284 );
xor ( n48286 , n48283 , n48284 );
xor ( n48287 , n47694 , n48016 );
and ( n48288 , n30144 , n48108 );
and ( n48289 , n48287 , n48288 );
xor ( n48290 , n48287 , n48288 );
xor ( n48291 , n47698 , n48014 );
and ( n48292 , n30149 , n48108 );
and ( n48293 , n48291 , n48292 );
xor ( n48294 , n48291 , n48292 );
xor ( n48295 , n47702 , n48012 );
and ( n48296 , n30154 , n48108 );
and ( n48297 , n48295 , n48296 );
xor ( n48298 , n48295 , n48296 );
xor ( n48299 , n47706 , n48010 );
and ( n48300 , n30159 , n48108 );
and ( n48301 , n48299 , n48300 );
xor ( n48302 , n48299 , n48300 );
xor ( n48303 , n47710 , n48008 );
and ( n48304 , n30164 , n48108 );
and ( n48305 , n48303 , n48304 );
xor ( n48306 , n48303 , n48304 );
xor ( n48307 , n47714 , n48006 );
and ( n48308 , n30169 , n48108 );
and ( n48309 , n48307 , n48308 );
xor ( n48310 , n48307 , n48308 );
xor ( n48311 , n47718 , n48004 );
and ( n48312 , n30174 , n48108 );
and ( n48313 , n48311 , n48312 );
xor ( n48314 , n48311 , n48312 );
xor ( n48315 , n47722 , n48002 );
and ( n48316 , n30179 , n48108 );
and ( n48317 , n48315 , n48316 );
xor ( n48318 , n48315 , n48316 );
xor ( n48319 , n47726 , n48000 );
and ( n48320 , n30184 , n48108 );
and ( n48321 , n48319 , n48320 );
xor ( n48322 , n48319 , n48320 );
xor ( n48323 , n47730 , n47998 );
and ( n48324 , n30189 , n48108 );
and ( n48325 , n48323 , n48324 );
xor ( n48326 , n48323 , n48324 );
xor ( n48327 , n47734 , n47996 );
and ( n48328 , n30194 , n48108 );
and ( n48329 , n48327 , n48328 );
xor ( n48330 , n48327 , n48328 );
xor ( n48331 , n47738 , n47994 );
and ( n48332 , n30199 , n48108 );
and ( n48333 , n48331 , n48332 );
xor ( n48334 , n48331 , n48332 );
xor ( n48335 , n47742 , n47992 );
and ( n48336 , n30204 , n48108 );
and ( n48337 , n48335 , n48336 );
xor ( n48338 , n48335 , n48336 );
xor ( n48339 , n47746 , n47990 );
and ( n48340 , n30209 , n48108 );
and ( n48341 , n48339 , n48340 );
xor ( n48342 , n48339 , n48340 );
xor ( n48343 , n47750 , n47988 );
and ( n48344 , n30214 , n48108 );
and ( n48345 , n48343 , n48344 );
xor ( n48346 , n48343 , n48344 );
xor ( n48347 , n47754 , n47986 );
and ( n48348 , n30219 , n48108 );
and ( n48349 , n48347 , n48348 );
xor ( n48350 , n48347 , n48348 );
xor ( n48351 , n47758 , n47984 );
and ( n48352 , n30224 , n48108 );
and ( n48353 , n48351 , n48352 );
xor ( n48354 , n48351 , n48352 );
xor ( n48355 , n47762 , n47982 );
and ( n48356 , n30229 , n48108 );
and ( n48357 , n48355 , n48356 );
xor ( n48358 , n48355 , n48356 );
xor ( n48359 , n47766 , n47980 );
and ( n48360 , n30234 , n48108 );
and ( n48361 , n48359 , n48360 );
xor ( n48362 , n48359 , n48360 );
xor ( n48363 , n47770 , n47978 );
and ( n48364 , n30239 , n48108 );
and ( n48365 , n48363 , n48364 );
xor ( n48366 , n48363 , n48364 );
xor ( n48367 , n47774 , n47976 );
and ( n48368 , n30244 , n48108 );
and ( n48369 , n48367 , n48368 );
xor ( n48370 , n48367 , n48368 );
xor ( n48371 , n47778 , n47974 );
and ( n48372 , n30249 , n48108 );
and ( n48373 , n48371 , n48372 );
xor ( n48374 , n48371 , n48372 );
xor ( n48375 , n47782 , n47972 );
and ( n48376 , n30254 , n48108 );
and ( n48377 , n48375 , n48376 );
xor ( n48378 , n48375 , n48376 );
xor ( n48379 , n47786 , n47970 );
and ( n48380 , n30259 , n48108 );
and ( n48381 , n48379 , n48380 );
xor ( n48382 , n48379 , n48380 );
xor ( n48383 , n47790 , n47968 );
and ( n48384 , n30264 , n48108 );
and ( n48385 , n48383 , n48384 );
xor ( n48386 , n48383 , n48384 );
xor ( n48387 , n47794 , n47966 );
and ( n48388 , n30269 , n48108 );
and ( n48389 , n48387 , n48388 );
xor ( n48390 , n48387 , n48388 );
xor ( n48391 , n47798 , n47964 );
and ( n48392 , n30274 , n48108 );
and ( n48393 , n48391 , n48392 );
xor ( n48394 , n48391 , n48392 );
xor ( n48395 , n47802 , n47962 );
and ( n48396 , n30279 , n48108 );
and ( n48397 , n48395 , n48396 );
xor ( n48398 , n48395 , n48396 );
xor ( n48399 , n47806 , n47960 );
and ( n48400 , n30284 , n48108 );
and ( n48401 , n48399 , n48400 );
xor ( n48402 , n48399 , n48400 );
xor ( n48403 , n47810 , n47958 );
and ( n48404 , n30289 , n48108 );
and ( n48405 , n48403 , n48404 );
xor ( n48406 , n48403 , n48404 );
xor ( n48407 , n47814 , n47956 );
and ( n48408 , n30294 , n48108 );
and ( n48409 , n48407 , n48408 );
xor ( n48410 , n48407 , n48408 );
xor ( n48411 , n47818 , n47954 );
and ( n48412 , n30299 , n48108 );
and ( n48413 , n48411 , n48412 );
xor ( n48414 , n48411 , n48412 );
xor ( n48415 , n47822 , n47952 );
and ( n48416 , n30304 , n48108 );
and ( n48417 , n48415 , n48416 );
xor ( n48418 , n48415 , n48416 );
xor ( n48419 , n47826 , n47950 );
and ( n48420 , n30309 , n48108 );
and ( n48421 , n48419 , n48420 );
xor ( n48422 , n48419 , n48420 );
xor ( n48423 , n47830 , n47948 );
and ( n48424 , n30314 , n48108 );
and ( n48425 , n48423 , n48424 );
xor ( n48426 , n48423 , n48424 );
xor ( n48427 , n47834 , n47946 );
and ( n48428 , n30319 , n48108 );
and ( n48429 , n48427 , n48428 );
xor ( n48430 , n48427 , n48428 );
xor ( n48431 , n47838 , n47944 );
and ( n48432 , n30324 , n48108 );
and ( n48433 , n48431 , n48432 );
xor ( n48434 , n48431 , n48432 );
xor ( n48435 , n47842 , n47942 );
and ( n48436 , n30329 , n48108 );
and ( n48437 , n48435 , n48436 );
xor ( n48438 , n48435 , n48436 );
xor ( n48439 , n47846 , n47940 );
and ( n48440 , n30334 , n48108 );
and ( n48441 , n48439 , n48440 );
xor ( n48442 , n48439 , n48440 );
xor ( n48443 , n47850 , n47938 );
and ( n48444 , n30339 , n48108 );
and ( n48445 , n48443 , n48444 );
xor ( n48446 , n48443 , n48444 );
xor ( n48447 , n47854 , n47936 );
and ( n48448 , n30344 , n48108 );
and ( n48449 , n48447 , n48448 );
xor ( n48450 , n48447 , n48448 );
xor ( n48451 , n47858 , n47934 );
and ( n48452 , n30349 , n48108 );
and ( n48453 , n48451 , n48452 );
xor ( n48454 , n48451 , n48452 );
xor ( n48455 , n47862 , n47932 );
and ( n48456 , n30354 , n48108 );
and ( n48457 , n48455 , n48456 );
xor ( n48458 , n48455 , n48456 );
xor ( n48459 , n47866 , n47930 );
and ( n48460 , n30359 , n48108 );
and ( n48461 , n48459 , n48460 );
xor ( n48462 , n48459 , n48460 );
xor ( n48463 , n47870 , n47928 );
and ( n48464 , n30364 , n48108 );
and ( n48465 , n48463 , n48464 );
xor ( n48466 , n48463 , n48464 );
xor ( n48467 , n47874 , n47926 );
and ( n48468 , n30369 , n48108 );
and ( n48469 , n48467 , n48468 );
xor ( n48470 , n48467 , n48468 );
xor ( n48471 , n47878 , n47924 );
and ( n48472 , n30374 , n48108 );
and ( n48473 , n48471 , n48472 );
xor ( n48474 , n48471 , n48472 );
xor ( n48475 , n47882 , n47922 );
and ( n48476 , n30379 , n48108 );
and ( n48477 , n48475 , n48476 );
xor ( n48478 , n48475 , n48476 );
xor ( n48479 , n47886 , n47920 );
and ( n48480 , n30384 , n48108 );
and ( n48481 , n48479 , n48480 );
xor ( n48482 , n48479 , n48480 );
xor ( n48483 , n47890 , n47918 );
and ( n48484 , n30389 , n48108 );
and ( n48485 , n48483 , n48484 );
xor ( n48486 , n48483 , n48484 );
xor ( n48487 , n47894 , n47916 );
and ( n48488 , n30394 , n48108 );
and ( n48489 , n48487 , n48488 );
xor ( n48490 , n48487 , n48488 );
xor ( n48491 , n47898 , n47914 );
and ( n48492 , n30399 , n48108 );
and ( n48493 , n48491 , n48492 );
xor ( n48494 , n48491 , n48492 );
xor ( n48495 , n47902 , n47912 );
and ( n48496 , n30404 , n48108 );
and ( n48497 , n48495 , n48496 );
xor ( n48498 , n48495 , n48496 );
xor ( n48499 , n47906 , n47910 );
and ( n48500 , n30409 , n48108 );
and ( n48501 , n48499 , n48500 );
buf ( n48502 , n48501 );
and ( n48503 , n48498 , n48502 );
or ( n48504 , n48497 , n48503 );
and ( n48505 , n48494 , n48504 );
or ( n48506 , n48493 , n48505 );
and ( n48507 , n48490 , n48506 );
or ( n48508 , n48489 , n48507 );
and ( n48509 , n48486 , n48508 );
or ( n48510 , n48485 , n48509 );
and ( n48511 , n48482 , n48510 );
or ( n48512 , n48481 , n48511 );
and ( n48513 , n48478 , n48512 );
or ( n48514 , n48477 , n48513 );
and ( n48515 , n48474 , n48514 );
or ( n48516 , n48473 , n48515 );
and ( n48517 , n48470 , n48516 );
or ( n48518 , n48469 , n48517 );
and ( n48519 , n48466 , n48518 );
or ( n48520 , n48465 , n48519 );
and ( n48521 , n48462 , n48520 );
or ( n48522 , n48461 , n48521 );
and ( n48523 , n48458 , n48522 );
or ( n48524 , n48457 , n48523 );
and ( n48525 , n48454 , n48524 );
or ( n48526 , n48453 , n48525 );
and ( n48527 , n48450 , n48526 );
or ( n48528 , n48449 , n48527 );
and ( n48529 , n48446 , n48528 );
or ( n48530 , n48445 , n48529 );
and ( n48531 , n48442 , n48530 );
or ( n48532 , n48441 , n48531 );
and ( n48533 , n48438 , n48532 );
or ( n48534 , n48437 , n48533 );
and ( n48535 , n48434 , n48534 );
or ( n48536 , n48433 , n48535 );
and ( n48537 , n48430 , n48536 );
or ( n48538 , n48429 , n48537 );
and ( n48539 , n48426 , n48538 );
or ( n48540 , n48425 , n48539 );
and ( n48541 , n48422 , n48540 );
or ( n48542 , n48421 , n48541 );
and ( n48543 , n48418 , n48542 );
or ( n48544 , n48417 , n48543 );
and ( n48545 , n48414 , n48544 );
or ( n48546 , n48413 , n48545 );
and ( n48547 , n48410 , n48546 );
or ( n48548 , n48409 , n48547 );
and ( n48549 , n48406 , n48548 );
or ( n48550 , n48405 , n48549 );
and ( n48551 , n48402 , n48550 );
or ( n48552 , n48401 , n48551 );
and ( n48553 , n48398 , n48552 );
or ( n48554 , n48397 , n48553 );
and ( n48555 , n48394 , n48554 );
or ( n48556 , n48393 , n48555 );
and ( n48557 , n48390 , n48556 );
or ( n48558 , n48389 , n48557 );
and ( n48559 , n48386 , n48558 );
or ( n48560 , n48385 , n48559 );
and ( n48561 , n48382 , n48560 );
or ( n48562 , n48381 , n48561 );
and ( n48563 , n48378 , n48562 );
or ( n48564 , n48377 , n48563 );
and ( n48565 , n48374 , n48564 );
or ( n48566 , n48373 , n48565 );
and ( n48567 , n48370 , n48566 );
or ( n48568 , n48369 , n48567 );
and ( n48569 , n48366 , n48568 );
or ( n48570 , n48365 , n48569 );
and ( n48571 , n48362 , n48570 );
or ( n48572 , n48361 , n48571 );
and ( n48573 , n48358 , n48572 );
or ( n48574 , n48357 , n48573 );
and ( n48575 , n48354 , n48574 );
or ( n48576 , n48353 , n48575 );
and ( n48577 , n48350 , n48576 );
or ( n48578 , n48349 , n48577 );
and ( n48579 , n48346 , n48578 );
or ( n48580 , n48345 , n48579 );
and ( n48581 , n48342 , n48580 );
or ( n48582 , n48341 , n48581 );
and ( n48583 , n48338 , n48582 );
or ( n48584 , n48337 , n48583 );
and ( n48585 , n48334 , n48584 );
or ( n48586 , n48333 , n48585 );
and ( n48587 , n48330 , n48586 );
or ( n48588 , n48329 , n48587 );
and ( n48589 , n48326 , n48588 );
or ( n48590 , n48325 , n48589 );
and ( n48591 , n48322 , n48590 );
or ( n48592 , n48321 , n48591 );
and ( n48593 , n48318 , n48592 );
or ( n48594 , n48317 , n48593 );
and ( n48595 , n48314 , n48594 );
or ( n48596 , n48313 , n48595 );
and ( n48597 , n48310 , n48596 );
or ( n48598 , n48309 , n48597 );
and ( n48599 , n48306 , n48598 );
or ( n48600 , n48305 , n48599 );
and ( n48601 , n48302 , n48600 );
or ( n48602 , n48301 , n48601 );
and ( n48603 , n48298 , n48602 );
or ( n48604 , n48297 , n48603 );
and ( n48605 , n48294 , n48604 );
or ( n48606 , n48293 , n48605 );
and ( n48607 , n48290 , n48606 );
or ( n48608 , n48289 , n48607 );
and ( n48609 , n48286 , n48608 );
or ( n48610 , n48285 , n48609 );
and ( n48611 , n48282 , n48610 );
or ( n48612 , n48281 , n48611 );
and ( n48613 , n48278 , n48612 );
or ( n48614 , n48277 , n48613 );
and ( n48615 , n48274 , n48614 );
or ( n48616 , n48273 , n48615 );
and ( n48617 , n48270 , n48616 );
or ( n48618 , n48269 , n48617 );
and ( n48619 , n48266 , n48618 );
or ( n48620 , n48265 , n48619 );
and ( n48621 , n48262 , n48620 );
or ( n48622 , n48261 , n48621 );
and ( n48623 , n48258 , n48622 );
or ( n48624 , n48257 , n48623 );
and ( n48625 , n48254 , n48624 );
or ( n48626 , n48253 , n48625 );
and ( n48627 , n48250 , n48626 );
or ( n48628 , n48249 , n48627 );
and ( n48629 , n48246 , n48628 );
or ( n48630 , n48245 , n48629 );
and ( n48631 , n48242 , n48630 );
or ( n48632 , n48241 , n48631 );
and ( n48633 , n48238 , n48632 );
or ( n48634 , n48237 , n48633 );
and ( n48635 , n48234 , n48634 );
or ( n48636 , n48233 , n48635 );
and ( n48637 , n48230 , n48636 );
or ( n48638 , n48229 , n48637 );
and ( n48639 , n48226 , n48638 );
or ( n48640 , n48225 , n48639 );
and ( n48641 , n48222 , n48640 );
or ( n48642 , n48221 , n48641 );
and ( n48643 , n48218 , n48642 );
or ( n48644 , n48217 , n48643 );
and ( n48645 , n48214 , n48644 );
or ( n48646 , n48213 , n48645 );
and ( n48647 , n48210 , n48646 );
or ( n48648 , n48209 , n48647 );
and ( n48649 , n48206 , n48648 );
or ( n48650 , n48205 , n48649 );
and ( n48651 , n48202 , n48650 );
or ( n48652 , n48201 , n48651 );
and ( n48653 , n48198 , n48652 );
or ( n48654 , n48197 , n48653 );
and ( n48655 , n48194 , n48654 );
or ( n48656 , n48193 , n48655 );
and ( n48657 , n48190 , n48656 );
or ( n48658 , n48189 , n48657 );
and ( n48659 , n48186 , n48658 );
or ( n48660 , n48185 , n48659 );
and ( n48661 , n48182 , n48660 );
or ( n48662 , n48181 , n48661 );
and ( n48663 , n48178 , n48662 );
or ( n48664 , n48177 , n48663 );
and ( n48665 , n48174 , n48664 );
or ( n48666 , n48173 , n48665 );
and ( n48667 , n48170 , n48666 );
or ( n48668 , n48169 , n48667 );
and ( n48669 , n48166 , n48668 );
or ( n48670 , n48165 , n48669 );
and ( n48671 , n48162 , n48670 );
or ( n48672 , n48161 , n48671 );
and ( n48673 , n48158 , n48672 );
or ( n48674 , n48157 , n48673 );
and ( n48675 , n48154 , n48674 );
or ( n48676 , n48153 , n48675 );
and ( n48677 , n48150 , n48676 );
or ( n48678 , n48149 , n48677 );
and ( n48679 , n48146 , n48678 );
or ( n48680 , n48145 , n48679 );
and ( n48681 , n48142 , n48680 );
or ( n48682 , n48141 , n48681 );
and ( n48683 , n48138 , n48682 );
or ( n48684 , n48137 , n48683 );
and ( n48685 , n48134 , n48684 );
or ( n48686 , n48133 , n48685 );
and ( n48687 , n48130 , n48686 );
or ( n48688 , n48129 , n48687 );
and ( n48689 , n48126 , n48688 );
or ( n48690 , n48125 , n48689 );
and ( n48691 , n48122 , n48690 );
or ( n48692 , n48121 , n48691 );
and ( n48693 , n48118 , n48692 );
or ( n48694 , n48117 , n48693 );
and ( n48695 , n48114 , n48694 );
or ( n48696 , n48113 , n48695 );
xor ( n48697 , n48110 , n48696 );
buf ( n48698 , n18048 );
and ( n48699 , n29924 , n48698 );
xor ( n48700 , n48697 , n48699 );
xor ( n48701 , n48114 , n48694 );
and ( n48702 , n29929 , n48698 );
and ( n48703 , n48701 , n48702 );
xor ( n48704 , n48701 , n48702 );
xor ( n48705 , n48118 , n48692 );
and ( n48706 , n29934 , n48698 );
and ( n48707 , n48705 , n48706 );
xor ( n48708 , n48705 , n48706 );
xor ( n48709 , n48122 , n48690 );
and ( n48710 , n29939 , n48698 );
and ( n48711 , n48709 , n48710 );
xor ( n48712 , n48709 , n48710 );
xor ( n48713 , n48126 , n48688 );
and ( n48714 , n29944 , n48698 );
and ( n48715 , n48713 , n48714 );
xor ( n48716 , n48713 , n48714 );
xor ( n48717 , n48130 , n48686 );
and ( n48718 , n29949 , n48698 );
and ( n48719 , n48717 , n48718 );
xor ( n48720 , n48717 , n48718 );
xor ( n48721 , n48134 , n48684 );
and ( n48722 , n29954 , n48698 );
and ( n48723 , n48721 , n48722 );
xor ( n48724 , n48721 , n48722 );
xor ( n48725 , n48138 , n48682 );
and ( n48726 , n29959 , n48698 );
and ( n48727 , n48725 , n48726 );
xor ( n48728 , n48725 , n48726 );
xor ( n48729 , n48142 , n48680 );
and ( n48730 , n29964 , n48698 );
and ( n48731 , n48729 , n48730 );
xor ( n48732 , n48729 , n48730 );
xor ( n48733 , n48146 , n48678 );
and ( n48734 , n29969 , n48698 );
and ( n48735 , n48733 , n48734 );
xor ( n48736 , n48733 , n48734 );
xor ( n48737 , n48150 , n48676 );
and ( n48738 , n29974 , n48698 );
and ( n48739 , n48737 , n48738 );
xor ( n48740 , n48737 , n48738 );
xor ( n48741 , n48154 , n48674 );
and ( n48742 , n29979 , n48698 );
and ( n48743 , n48741 , n48742 );
xor ( n48744 , n48741 , n48742 );
xor ( n48745 , n48158 , n48672 );
and ( n48746 , n29984 , n48698 );
and ( n48747 , n48745 , n48746 );
xor ( n48748 , n48745 , n48746 );
xor ( n48749 , n48162 , n48670 );
and ( n48750 , n29989 , n48698 );
and ( n48751 , n48749 , n48750 );
xor ( n48752 , n48749 , n48750 );
xor ( n48753 , n48166 , n48668 );
and ( n48754 , n29994 , n48698 );
and ( n48755 , n48753 , n48754 );
xor ( n48756 , n48753 , n48754 );
xor ( n48757 , n48170 , n48666 );
and ( n48758 , n29999 , n48698 );
and ( n48759 , n48757 , n48758 );
xor ( n48760 , n48757 , n48758 );
xor ( n48761 , n48174 , n48664 );
and ( n48762 , n30004 , n48698 );
and ( n48763 , n48761 , n48762 );
xor ( n48764 , n48761 , n48762 );
xor ( n48765 , n48178 , n48662 );
and ( n48766 , n30009 , n48698 );
and ( n48767 , n48765 , n48766 );
xor ( n48768 , n48765 , n48766 );
xor ( n48769 , n48182 , n48660 );
and ( n48770 , n30014 , n48698 );
and ( n48771 , n48769 , n48770 );
xor ( n48772 , n48769 , n48770 );
xor ( n48773 , n48186 , n48658 );
and ( n48774 , n30019 , n48698 );
and ( n48775 , n48773 , n48774 );
xor ( n48776 , n48773 , n48774 );
xor ( n48777 , n48190 , n48656 );
and ( n48778 , n30024 , n48698 );
and ( n48779 , n48777 , n48778 );
xor ( n48780 , n48777 , n48778 );
xor ( n48781 , n48194 , n48654 );
and ( n48782 , n30029 , n48698 );
and ( n48783 , n48781 , n48782 );
xor ( n48784 , n48781 , n48782 );
xor ( n48785 , n48198 , n48652 );
and ( n48786 , n30034 , n48698 );
and ( n48787 , n48785 , n48786 );
xor ( n48788 , n48785 , n48786 );
xor ( n48789 , n48202 , n48650 );
and ( n48790 , n30039 , n48698 );
and ( n48791 , n48789 , n48790 );
xor ( n48792 , n48789 , n48790 );
xor ( n48793 , n48206 , n48648 );
and ( n48794 , n30044 , n48698 );
and ( n48795 , n48793 , n48794 );
xor ( n48796 , n48793 , n48794 );
xor ( n48797 , n48210 , n48646 );
and ( n48798 , n30049 , n48698 );
and ( n48799 , n48797 , n48798 );
xor ( n48800 , n48797 , n48798 );
xor ( n48801 , n48214 , n48644 );
and ( n48802 , n30054 , n48698 );
and ( n48803 , n48801 , n48802 );
xor ( n48804 , n48801 , n48802 );
xor ( n48805 , n48218 , n48642 );
and ( n48806 , n30059 , n48698 );
and ( n48807 , n48805 , n48806 );
xor ( n48808 , n48805 , n48806 );
xor ( n48809 , n48222 , n48640 );
and ( n48810 , n30064 , n48698 );
and ( n48811 , n48809 , n48810 );
xor ( n48812 , n48809 , n48810 );
xor ( n48813 , n48226 , n48638 );
and ( n48814 , n30069 , n48698 );
and ( n48815 , n48813 , n48814 );
xor ( n48816 , n48813 , n48814 );
xor ( n48817 , n48230 , n48636 );
and ( n48818 , n30074 , n48698 );
and ( n48819 , n48817 , n48818 );
xor ( n48820 , n48817 , n48818 );
xor ( n48821 , n48234 , n48634 );
and ( n48822 , n30079 , n48698 );
and ( n48823 , n48821 , n48822 );
xor ( n48824 , n48821 , n48822 );
xor ( n48825 , n48238 , n48632 );
and ( n48826 , n30084 , n48698 );
and ( n48827 , n48825 , n48826 );
xor ( n48828 , n48825 , n48826 );
xor ( n48829 , n48242 , n48630 );
and ( n48830 , n30089 , n48698 );
and ( n48831 , n48829 , n48830 );
xor ( n48832 , n48829 , n48830 );
xor ( n48833 , n48246 , n48628 );
and ( n48834 , n30094 , n48698 );
and ( n48835 , n48833 , n48834 );
xor ( n48836 , n48833 , n48834 );
xor ( n48837 , n48250 , n48626 );
and ( n48838 , n30099 , n48698 );
and ( n48839 , n48837 , n48838 );
xor ( n48840 , n48837 , n48838 );
xor ( n48841 , n48254 , n48624 );
and ( n48842 , n30104 , n48698 );
and ( n48843 , n48841 , n48842 );
xor ( n48844 , n48841 , n48842 );
xor ( n48845 , n48258 , n48622 );
and ( n48846 , n30109 , n48698 );
and ( n48847 , n48845 , n48846 );
xor ( n48848 , n48845 , n48846 );
xor ( n48849 , n48262 , n48620 );
and ( n48850 , n30114 , n48698 );
and ( n48851 , n48849 , n48850 );
xor ( n48852 , n48849 , n48850 );
xor ( n48853 , n48266 , n48618 );
and ( n48854 , n30119 , n48698 );
and ( n48855 , n48853 , n48854 );
xor ( n48856 , n48853 , n48854 );
xor ( n48857 , n48270 , n48616 );
and ( n48858 , n30124 , n48698 );
and ( n48859 , n48857 , n48858 );
xor ( n48860 , n48857 , n48858 );
xor ( n48861 , n48274 , n48614 );
and ( n48862 , n30129 , n48698 );
and ( n48863 , n48861 , n48862 );
xor ( n48864 , n48861 , n48862 );
xor ( n48865 , n48278 , n48612 );
and ( n48866 , n30134 , n48698 );
and ( n48867 , n48865 , n48866 );
xor ( n48868 , n48865 , n48866 );
xor ( n48869 , n48282 , n48610 );
and ( n48870 , n30139 , n48698 );
and ( n48871 , n48869 , n48870 );
xor ( n48872 , n48869 , n48870 );
xor ( n48873 , n48286 , n48608 );
and ( n48874 , n30144 , n48698 );
and ( n48875 , n48873 , n48874 );
xor ( n48876 , n48873 , n48874 );
xor ( n48877 , n48290 , n48606 );
and ( n48878 , n30149 , n48698 );
and ( n48879 , n48877 , n48878 );
xor ( n48880 , n48877 , n48878 );
xor ( n48881 , n48294 , n48604 );
and ( n48882 , n30154 , n48698 );
and ( n48883 , n48881 , n48882 );
xor ( n48884 , n48881 , n48882 );
xor ( n48885 , n48298 , n48602 );
and ( n48886 , n30159 , n48698 );
and ( n48887 , n48885 , n48886 );
xor ( n48888 , n48885 , n48886 );
xor ( n48889 , n48302 , n48600 );
and ( n48890 , n30164 , n48698 );
and ( n48891 , n48889 , n48890 );
xor ( n48892 , n48889 , n48890 );
xor ( n48893 , n48306 , n48598 );
and ( n48894 , n30169 , n48698 );
and ( n48895 , n48893 , n48894 );
xor ( n48896 , n48893 , n48894 );
xor ( n48897 , n48310 , n48596 );
and ( n48898 , n30174 , n48698 );
and ( n48899 , n48897 , n48898 );
xor ( n48900 , n48897 , n48898 );
xor ( n48901 , n48314 , n48594 );
and ( n48902 , n30179 , n48698 );
and ( n48903 , n48901 , n48902 );
xor ( n48904 , n48901 , n48902 );
xor ( n48905 , n48318 , n48592 );
and ( n48906 , n30184 , n48698 );
and ( n48907 , n48905 , n48906 );
xor ( n48908 , n48905 , n48906 );
xor ( n48909 , n48322 , n48590 );
and ( n48910 , n30189 , n48698 );
and ( n48911 , n48909 , n48910 );
xor ( n48912 , n48909 , n48910 );
xor ( n48913 , n48326 , n48588 );
and ( n48914 , n30194 , n48698 );
and ( n48915 , n48913 , n48914 );
xor ( n48916 , n48913 , n48914 );
xor ( n48917 , n48330 , n48586 );
and ( n48918 , n30199 , n48698 );
and ( n48919 , n48917 , n48918 );
xor ( n48920 , n48917 , n48918 );
xor ( n48921 , n48334 , n48584 );
and ( n48922 , n30204 , n48698 );
and ( n48923 , n48921 , n48922 );
xor ( n48924 , n48921 , n48922 );
xor ( n48925 , n48338 , n48582 );
and ( n48926 , n30209 , n48698 );
and ( n48927 , n48925 , n48926 );
xor ( n48928 , n48925 , n48926 );
xor ( n48929 , n48342 , n48580 );
and ( n48930 , n30214 , n48698 );
and ( n48931 , n48929 , n48930 );
xor ( n48932 , n48929 , n48930 );
xor ( n48933 , n48346 , n48578 );
and ( n48934 , n30219 , n48698 );
and ( n48935 , n48933 , n48934 );
xor ( n48936 , n48933 , n48934 );
xor ( n48937 , n48350 , n48576 );
and ( n48938 , n30224 , n48698 );
and ( n48939 , n48937 , n48938 );
xor ( n48940 , n48937 , n48938 );
xor ( n48941 , n48354 , n48574 );
and ( n48942 , n30229 , n48698 );
and ( n48943 , n48941 , n48942 );
xor ( n48944 , n48941 , n48942 );
xor ( n48945 , n48358 , n48572 );
and ( n48946 , n30234 , n48698 );
and ( n48947 , n48945 , n48946 );
xor ( n48948 , n48945 , n48946 );
xor ( n48949 , n48362 , n48570 );
and ( n48950 , n30239 , n48698 );
and ( n48951 , n48949 , n48950 );
xor ( n48952 , n48949 , n48950 );
xor ( n48953 , n48366 , n48568 );
and ( n48954 , n30244 , n48698 );
and ( n48955 , n48953 , n48954 );
xor ( n48956 , n48953 , n48954 );
xor ( n48957 , n48370 , n48566 );
and ( n48958 , n30249 , n48698 );
and ( n48959 , n48957 , n48958 );
xor ( n48960 , n48957 , n48958 );
xor ( n48961 , n48374 , n48564 );
and ( n48962 , n30254 , n48698 );
and ( n48963 , n48961 , n48962 );
xor ( n48964 , n48961 , n48962 );
xor ( n48965 , n48378 , n48562 );
and ( n48966 , n30259 , n48698 );
and ( n48967 , n48965 , n48966 );
xor ( n48968 , n48965 , n48966 );
xor ( n48969 , n48382 , n48560 );
and ( n48970 , n30264 , n48698 );
and ( n48971 , n48969 , n48970 );
xor ( n48972 , n48969 , n48970 );
xor ( n48973 , n48386 , n48558 );
and ( n48974 , n30269 , n48698 );
and ( n48975 , n48973 , n48974 );
xor ( n48976 , n48973 , n48974 );
xor ( n48977 , n48390 , n48556 );
and ( n48978 , n30274 , n48698 );
and ( n48979 , n48977 , n48978 );
xor ( n48980 , n48977 , n48978 );
xor ( n48981 , n48394 , n48554 );
and ( n48982 , n30279 , n48698 );
and ( n48983 , n48981 , n48982 );
xor ( n48984 , n48981 , n48982 );
xor ( n48985 , n48398 , n48552 );
and ( n48986 , n30284 , n48698 );
and ( n48987 , n48985 , n48986 );
xor ( n48988 , n48985 , n48986 );
xor ( n48989 , n48402 , n48550 );
and ( n48990 , n30289 , n48698 );
and ( n48991 , n48989 , n48990 );
xor ( n48992 , n48989 , n48990 );
xor ( n48993 , n48406 , n48548 );
and ( n48994 , n30294 , n48698 );
and ( n48995 , n48993 , n48994 );
xor ( n48996 , n48993 , n48994 );
xor ( n48997 , n48410 , n48546 );
and ( n48998 , n30299 , n48698 );
and ( n48999 , n48997 , n48998 );
xor ( n49000 , n48997 , n48998 );
xor ( n49001 , n48414 , n48544 );
and ( n49002 , n30304 , n48698 );
and ( n49003 , n49001 , n49002 );
xor ( n49004 , n49001 , n49002 );
xor ( n49005 , n48418 , n48542 );
and ( n49006 , n30309 , n48698 );
and ( n49007 , n49005 , n49006 );
xor ( n49008 , n49005 , n49006 );
xor ( n49009 , n48422 , n48540 );
and ( n49010 , n30314 , n48698 );
and ( n49011 , n49009 , n49010 );
xor ( n49012 , n49009 , n49010 );
xor ( n49013 , n48426 , n48538 );
and ( n49014 , n30319 , n48698 );
and ( n49015 , n49013 , n49014 );
xor ( n49016 , n49013 , n49014 );
xor ( n49017 , n48430 , n48536 );
and ( n49018 , n30324 , n48698 );
and ( n49019 , n49017 , n49018 );
xor ( n49020 , n49017 , n49018 );
xor ( n49021 , n48434 , n48534 );
and ( n49022 , n30329 , n48698 );
and ( n49023 , n49021 , n49022 );
xor ( n49024 , n49021 , n49022 );
xor ( n49025 , n48438 , n48532 );
and ( n49026 , n30334 , n48698 );
and ( n49027 , n49025 , n49026 );
xor ( n49028 , n49025 , n49026 );
xor ( n49029 , n48442 , n48530 );
and ( n49030 , n30339 , n48698 );
and ( n49031 , n49029 , n49030 );
xor ( n49032 , n49029 , n49030 );
xor ( n49033 , n48446 , n48528 );
and ( n49034 , n30344 , n48698 );
and ( n49035 , n49033 , n49034 );
xor ( n49036 , n49033 , n49034 );
xor ( n49037 , n48450 , n48526 );
and ( n49038 , n30349 , n48698 );
and ( n49039 , n49037 , n49038 );
xor ( n49040 , n49037 , n49038 );
xor ( n49041 , n48454 , n48524 );
and ( n49042 , n30354 , n48698 );
and ( n49043 , n49041 , n49042 );
xor ( n49044 , n49041 , n49042 );
xor ( n49045 , n48458 , n48522 );
and ( n49046 , n30359 , n48698 );
and ( n49047 , n49045 , n49046 );
xor ( n49048 , n49045 , n49046 );
xor ( n49049 , n48462 , n48520 );
and ( n49050 , n30364 , n48698 );
and ( n49051 , n49049 , n49050 );
xor ( n49052 , n49049 , n49050 );
xor ( n49053 , n48466 , n48518 );
and ( n49054 , n30369 , n48698 );
and ( n49055 , n49053 , n49054 );
xor ( n49056 , n49053 , n49054 );
xor ( n49057 , n48470 , n48516 );
and ( n49058 , n30374 , n48698 );
and ( n49059 , n49057 , n49058 );
xor ( n49060 , n49057 , n49058 );
xor ( n49061 , n48474 , n48514 );
and ( n49062 , n30379 , n48698 );
and ( n49063 , n49061 , n49062 );
xor ( n49064 , n49061 , n49062 );
xor ( n49065 , n48478 , n48512 );
and ( n49066 , n30384 , n48698 );
and ( n49067 , n49065 , n49066 );
xor ( n49068 , n49065 , n49066 );
xor ( n49069 , n48482 , n48510 );
and ( n49070 , n30389 , n48698 );
and ( n49071 , n49069 , n49070 );
xor ( n49072 , n49069 , n49070 );
xor ( n49073 , n48486 , n48508 );
and ( n49074 , n30394 , n48698 );
and ( n49075 , n49073 , n49074 );
xor ( n49076 , n49073 , n49074 );
xor ( n49077 , n48490 , n48506 );
and ( n49078 , n30399 , n48698 );
and ( n49079 , n49077 , n49078 );
xor ( n49080 , n49077 , n49078 );
xor ( n49081 , n48494 , n48504 );
and ( n49082 , n30404 , n48698 );
and ( n49083 , n49081 , n49082 );
xor ( n49084 , n49081 , n49082 );
xor ( n49085 , n48498 , n48502 );
and ( n49086 , n30409 , n48698 );
and ( n49087 , n49085 , n49086 );
buf ( n49088 , n49087 );
and ( n49089 , n49084 , n49088 );
or ( n49090 , n49083 , n49089 );
and ( n49091 , n49080 , n49090 );
or ( n49092 , n49079 , n49091 );
and ( n49093 , n49076 , n49092 );
or ( n49094 , n49075 , n49093 );
and ( n49095 , n49072 , n49094 );
or ( n49096 , n49071 , n49095 );
and ( n49097 , n49068 , n49096 );
or ( n49098 , n49067 , n49097 );
and ( n49099 , n49064 , n49098 );
or ( n49100 , n49063 , n49099 );
and ( n49101 , n49060 , n49100 );
or ( n49102 , n49059 , n49101 );
and ( n49103 , n49056 , n49102 );
or ( n49104 , n49055 , n49103 );
and ( n49105 , n49052 , n49104 );
or ( n49106 , n49051 , n49105 );
and ( n49107 , n49048 , n49106 );
or ( n49108 , n49047 , n49107 );
and ( n49109 , n49044 , n49108 );
or ( n49110 , n49043 , n49109 );
and ( n49111 , n49040 , n49110 );
or ( n49112 , n49039 , n49111 );
and ( n49113 , n49036 , n49112 );
or ( n49114 , n49035 , n49113 );
and ( n49115 , n49032 , n49114 );
or ( n49116 , n49031 , n49115 );
and ( n49117 , n49028 , n49116 );
or ( n49118 , n49027 , n49117 );
and ( n49119 , n49024 , n49118 );
or ( n49120 , n49023 , n49119 );
and ( n49121 , n49020 , n49120 );
or ( n49122 , n49019 , n49121 );
and ( n49123 , n49016 , n49122 );
or ( n49124 , n49015 , n49123 );
and ( n49125 , n49012 , n49124 );
or ( n49126 , n49011 , n49125 );
and ( n49127 , n49008 , n49126 );
or ( n49128 , n49007 , n49127 );
and ( n49129 , n49004 , n49128 );
or ( n49130 , n49003 , n49129 );
and ( n49131 , n49000 , n49130 );
or ( n49132 , n48999 , n49131 );
and ( n49133 , n48996 , n49132 );
or ( n49134 , n48995 , n49133 );
and ( n49135 , n48992 , n49134 );
or ( n49136 , n48991 , n49135 );
and ( n49137 , n48988 , n49136 );
or ( n49138 , n48987 , n49137 );
and ( n49139 , n48984 , n49138 );
or ( n49140 , n48983 , n49139 );
and ( n49141 , n48980 , n49140 );
or ( n49142 , n48979 , n49141 );
and ( n49143 , n48976 , n49142 );
or ( n49144 , n48975 , n49143 );
and ( n49145 , n48972 , n49144 );
or ( n49146 , n48971 , n49145 );
and ( n49147 , n48968 , n49146 );
or ( n49148 , n48967 , n49147 );
and ( n49149 , n48964 , n49148 );
or ( n49150 , n48963 , n49149 );
and ( n49151 , n48960 , n49150 );
or ( n49152 , n48959 , n49151 );
and ( n49153 , n48956 , n49152 );
or ( n49154 , n48955 , n49153 );
and ( n49155 , n48952 , n49154 );
or ( n49156 , n48951 , n49155 );
and ( n49157 , n48948 , n49156 );
or ( n49158 , n48947 , n49157 );
and ( n49159 , n48944 , n49158 );
or ( n49160 , n48943 , n49159 );
and ( n49161 , n48940 , n49160 );
or ( n49162 , n48939 , n49161 );
and ( n49163 , n48936 , n49162 );
or ( n49164 , n48935 , n49163 );
and ( n49165 , n48932 , n49164 );
or ( n49166 , n48931 , n49165 );
and ( n49167 , n48928 , n49166 );
or ( n49168 , n48927 , n49167 );
and ( n49169 , n48924 , n49168 );
or ( n49170 , n48923 , n49169 );
and ( n49171 , n48920 , n49170 );
or ( n49172 , n48919 , n49171 );
and ( n49173 , n48916 , n49172 );
or ( n49174 , n48915 , n49173 );
and ( n49175 , n48912 , n49174 );
or ( n49176 , n48911 , n49175 );
and ( n49177 , n48908 , n49176 );
or ( n49178 , n48907 , n49177 );
and ( n49179 , n48904 , n49178 );
or ( n49180 , n48903 , n49179 );
and ( n49181 , n48900 , n49180 );
or ( n49182 , n48899 , n49181 );
and ( n49183 , n48896 , n49182 );
or ( n49184 , n48895 , n49183 );
and ( n49185 , n48892 , n49184 );
or ( n49186 , n48891 , n49185 );
and ( n49187 , n48888 , n49186 );
or ( n49188 , n48887 , n49187 );
and ( n49189 , n48884 , n49188 );
or ( n49190 , n48883 , n49189 );
and ( n49191 , n48880 , n49190 );
or ( n49192 , n48879 , n49191 );
and ( n49193 , n48876 , n49192 );
or ( n49194 , n48875 , n49193 );
and ( n49195 , n48872 , n49194 );
or ( n49196 , n48871 , n49195 );
and ( n49197 , n48868 , n49196 );
or ( n49198 , n48867 , n49197 );
and ( n49199 , n48864 , n49198 );
or ( n49200 , n48863 , n49199 );
and ( n49201 , n48860 , n49200 );
or ( n49202 , n48859 , n49201 );
and ( n49203 , n48856 , n49202 );
or ( n49204 , n48855 , n49203 );
and ( n49205 , n48852 , n49204 );
or ( n49206 , n48851 , n49205 );
and ( n49207 , n48848 , n49206 );
or ( n49208 , n48847 , n49207 );
and ( n49209 , n48844 , n49208 );
or ( n49210 , n48843 , n49209 );
and ( n49211 , n48840 , n49210 );
or ( n49212 , n48839 , n49211 );
and ( n49213 , n48836 , n49212 );
or ( n49214 , n48835 , n49213 );
and ( n49215 , n48832 , n49214 );
or ( n49216 , n48831 , n49215 );
and ( n49217 , n48828 , n49216 );
or ( n49218 , n48827 , n49217 );
and ( n49219 , n48824 , n49218 );
or ( n49220 , n48823 , n49219 );
and ( n49221 , n48820 , n49220 );
or ( n49222 , n48819 , n49221 );
and ( n49223 , n48816 , n49222 );
or ( n49224 , n48815 , n49223 );
and ( n49225 , n48812 , n49224 );
or ( n49226 , n48811 , n49225 );
and ( n49227 , n48808 , n49226 );
or ( n49228 , n48807 , n49227 );
and ( n49229 , n48804 , n49228 );
or ( n49230 , n48803 , n49229 );
and ( n49231 , n48800 , n49230 );
or ( n49232 , n48799 , n49231 );
and ( n49233 , n48796 , n49232 );
or ( n49234 , n48795 , n49233 );
and ( n49235 , n48792 , n49234 );
or ( n49236 , n48791 , n49235 );
and ( n49237 , n48788 , n49236 );
or ( n49238 , n48787 , n49237 );
and ( n49239 , n48784 , n49238 );
or ( n49240 , n48783 , n49239 );
and ( n49241 , n48780 , n49240 );
or ( n49242 , n48779 , n49241 );
and ( n49243 , n48776 , n49242 );
or ( n49244 , n48775 , n49243 );
and ( n49245 , n48772 , n49244 );
or ( n49246 , n48771 , n49245 );
and ( n49247 , n48768 , n49246 );
or ( n49248 , n48767 , n49247 );
and ( n49249 , n48764 , n49248 );
or ( n49250 , n48763 , n49249 );
and ( n49251 , n48760 , n49250 );
or ( n49252 , n48759 , n49251 );
and ( n49253 , n48756 , n49252 );
or ( n49254 , n48755 , n49253 );
and ( n49255 , n48752 , n49254 );
or ( n49256 , n48751 , n49255 );
and ( n49257 , n48748 , n49256 );
or ( n49258 , n48747 , n49257 );
and ( n49259 , n48744 , n49258 );
or ( n49260 , n48743 , n49259 );
and ( n49261 , n48740 , n49260 );
or ( n49262 , n48739 , n49261 );
and ( n49263 , n48736 , n49262 );
or ( n49264 , n48735 , n49263 );
and ( n49265 , n48732 , n49264 );
or ( n49266 , n48731 , n49265 );
and ( n49267 , n48728 , n49266 );
or ( n49268 , n48727 , n49267 );
and ( n49269 , n48724 , n49268 );
or ( n49270 , n48723 , n49269 );
and ( n49271 , n48720 , n49270 );
or ( n49272 , n48719 , n49271 );
and ( n49273 , n48716 , n49272 );
or ( n49274 , n48715 , n49273 );
and ( n49275 , n48712 , n49274 );
or ( n49276 , n48711 , n49275 );
and ( n49277 , n48708 , n49276 );
or ( n49278 , n48707 , n49277 );
and ( n49279 , n48704 , n49278 );
or ( n49280 , n48703 , n49279 );
xor ( n49281 , n48700 , n49280 );
buf ( n49282 , n18046 );
and ( n49283 , n29929 , n49282 );
xor ( n49284 , n49281 , n49283 );
xor ( n49285 , n48704 , n49278 );
and ( n49286 , n29934 , n49282 );
and ( n49287 , n49285 , n49286 );
xor ( n49288 , n49285 , n49286 );
xor ( n49289 , n48708 , n49276 );
and ( n49290 , n29939 , n49282 );
and ( n49291 , n49289 , n49290 );
xor ( n49292 , n49289 , n49290 );
xor ( n49293 , n48712 , n49274 );
and ( n49294 , n29944 , n49282 );
and ( n49295 , n49293 , n49294 );
xor ( n49296 , n49293 , n49294 );
xor ( n49297 , n48716 , n49272 );
and ( n49298 , n29949 , n49282 );
and ( n49299 , n49297 , n49298 );
xor ( n49300 , n49297 , n49298 );
xor ( n49301 , n48720 , n49270 );
and ( n49302 , n29954 , n49282 );
and ( n49303 , n49301 , n49302 );
xor ( n49304 , n49301 , n49302 );
xor ( n49305 , n48724 , n49268 );
and ( n49306 , n29959 , n49282 );
and ( n49307 , n49305 , n49306 );
xor ( n49308 , n49305 , n49306 );
xor ( n49309 , n48728 , n49266 );
and ( n49310 , n29964 , n49282 );
and ( n49311 , n49309 , n49310 );
xor ( n49312 , n49309 , n49310 );
xor ( n49313 , n48732 , n49264 );
and ( n49314 , n29969 , n49282 );
and ( n49315 , n49313 , n49314 );
xor ( n49316 , n49313 , n49314 );
xor ( n49317 , n48736 , n49262 );
and ( n49318 , n29974 , n49282 );
and ( n49319 , n49317 , n49318 );
xor ( n49320 , n49317 , n49318 );
xor ( n49321 , n48740 , n49260 );
and ( n49322 , n29979 , n49282 );
and ( n49323 , n49321 , n49322 );
xor ( n49324 , n49321 , n49322 );
xor ( n49325 , n48744 , n49258 );
and ( n49326 , n29984 , n49282 );
and ( n49327 , n49325 , n49326 );
xor ( n49328 , n49325 , n49326 );
xor ( n49329 , n48748 , n49256 );
and ( n49330 , n29989 , n49282 );
and ( n49331 , n49329 , n49330 );
xor ( n49332 , n49329 , n49330 );
xor ( n49333 , n48752 , n49254 );
and ( n49334 , n29994 , n49282 );
and ( n49335 , n49333 , n49334 );
xor ( n49336 , n49333 , n49334 );
xor ( n49337 , n48756 , n49252 );
and ( n49338 , n29999 , n49282 );
and ( n49339 , n49337 , n49338 );
xor ( n49340 , n49337 , n49338 );
xor ( n49341 , n48760 , n49250 );
and ( n49342 , n30004 , n49282 );
and ( n49343 , n49341 , n49342 );
xor ( n49344 , n49341 , n49342 );
xor ( n49345 , n48764 , n49248 );
and ( n49346 , n30009 , n49282 );
and ( n49347 , n49345 , n49346 );
xor ( n49348 , n49345 , n49346 );
xor ( n49349 , n48768 , n49246 );
and ( n49350 , n30014 , n49282 );
and ( n49351 , n49349 , n49350 );
xor ( n49352 , n49349 , n49350 );
xor ( n49353 , n48772 , n49244 );
and ( n49354 , n30019 , n49282 );
and ( n49355 , n49353 , n49354 );
xor ( n49356 , n49353 , n49354 );
xor ( n49357 , n48776 , n49242 );
and ( n49358 , n30024 , n49282 );
and ( n49359 , n49357 , n49358 );
xor ( n49360 , n49357 , n49358 );
xor ( n49361 , n48780 , n49240 );
and ( n49362 , n30029 , n49282 );
and ( n49363 , n49361 , n49362 );
xor ( n49364 , n49361 , n49362 );
xor ( n49365 , n48784 , n49238 );
and ( n49366 , n30034 , n49282 );
and ( n49367 , n49365 , n49366 );
xor ( n49368 , n49365 , n49366 );
xor ( n49369 , n48788 , n49236 );
and ( n49370 , n30039 , n49282 );
and ( n49371 , n49369 , n49370 );
xor ( n49372 , n49369 , n49370 );
xor ( n49373 , n48792 , n49234 );
and ( n49374 , n30044 , n49282 );
and ( n49375 , n49373 , n49374 );
xor ( n49376 , n49373 , n49374 );
xor ( n49377 , n48796 , n49232 );
and ( n49378 , n30049 , n49282 );
and ( n49379 , n49377 , n49378 );
xor ( n49380 , n49377 , n49378 );
xor ( n49381 , n48800 , n49230 );
and ( n49382 , n30054 , n49282 );
and ( n49383 , n49381 , n49382 );
xor ( n49384 , n49381 , n49382 );
xor ( n49385 , n48804 , n49228 );
and ( n49386 , n30059 , n49282 );
and ( n49387 , n49385 , n49386 );
xor ( n49388 , n49385 , n49386 );
xor ( n49389 , n48808 , n49226 );
and ( n49390 , n30064 , n49282 );
and ( n49391 , n49389 , n49390 );
xor ( n49392 , n49389 , n49390 );
xor ( n49393 , n48812 , n49224 );
and ( n49394 , n30069 , n49282 );
and ( n49395 , n49393 , n49394 );
xor ( n49396 , n49393 , n49394 );
xor ( n49397 , n48816 , n49222 );
and ( n49398 , n30074 , n49282 );
and ( n49399 , n49397 , n49398 );
xor ( n49400 , n49397 , n49398 );
xor ( n49401 , n48820 , n49220 );
and ( n49402 , n30079 , n49282 );
and ( n49403 , n49401 , n49402 );
xor ( n49404 , n49401 , n49402 );
xor ( n49405 , n48824 , n49218 );
and ( n49406 , n30084 , n49282 );
and ( n49407 , n49405 , n49406 );
xor ( n49408 , n49405 , n49406 );
xor ( n49409 , n48828 , n49216 );
and ( n49410 , n30089 , n49282 );
and ( n49411 , n49409 , n49410 );
xor ( n49412 , n49409 , n49410 );
xor ( n49413 , n48832 , n49214 );
and ( n49414 , n30094 , n49282 );
and ( n49415 , n49413 , n49414 );
xor ( n49416 , n49413 , n49414 );
xor ( n49417 , n48836 , n49212 );
and ( n49418 , n30099 , n49282 );
and ( n49419 , n49417 , n49418 );
xor ( n49420 , n49417 , n49418 );
xor ( n49421 , n48840 , n49210 );
and ( n49422 , n30104 , n49282 );
and ( n49423 , n49421 , n49422 );
xor ( n49424 , n49421 , n49422 );
xor ( n49425 , n48844 , n49208 );
and ( n49426 , n30109 , n49282 );
and ( n49427 , n49425 , n49426 );
xor ( n49428 , n49425 , n49426 );
xor ( n49429 , n48848 , n49206 );
and ( n49430 , n30114 , n49282 );
and ( n49431 , n49429 , n49430 );
xor ( n49432 , n49429 , n49430 );
xor ( n49433 , n48852 , n49204 );
and ( n49434 , n30119 , n49282 );
and ( n49435 , n49433 , n49434 );
xor ( n49436 , n49433 , n49434 );
xor ( n49437 , n48856 , n49202 );
and ( n49438 , n30124 , n49282 );
and ( n49439 , n49437 , n49438 );
xor ( n49440 , n49437 , n49438 );
xor ( n49441 , n48860 , n49200 );
and ( n49442 , n30129 , n49282 );
and ( n49443 , n49441 , n49442 );
xor ( n49444 , n49441 , n49442 );
xor ( n49445 , n48864 , n49198 );
and ( n49446 , n30134 , n49282 );
and ( n49447 , n49445 , n49446 );
xor ( n49448 , n49445 , n49446 );
xor ( n49449 , n48868 , n49196 );
and ( n49450 , n30139 , n49282 );
and ( n49451 , n49449 , n49450 );
xor ( n49452 , n49449 , n49450 );
xor ( n49453 , n48872 , n49194 );
and ( n49454 , n30144 , n49282 );
and ( n49455 , n49453 , n49454 );
xor ( n49456 , n49453 , n49454 );
xor ( n49457 , n48876 , n49192 );
and ( n49458 , n30149 , n49282 );
and ( n49459 , n49457 , n49458 );
xor ( n49460 , n49457 , n49458 );
xor ( n49461 , n48880 , n49190 );
and ( n49462 , n30154 , n49282 );
and ( n49463 , n49461 , n49462 );
xor ( n49464 , n49461 , n49462 );
xor ( n49465 , n48884 , n49188 );
and ( n49466 , n30159 , n49282 );
and ( n49467 , n49465 , n49466 );
xor ( n49468 , n49465 , n49466 );
xor ( n49469 , n48888 , n49186 );
and ( n49470 , n30164 , n49282 );
and ( n49471 , n49469 , n49470 );
xor ( n49472 , n49469 , n49470 );
xor ( n49473 , n48892 , n49184 );
and ( n49474 , n30169 , n49282 );
and ( n49475 , n49473 , n49474 );
xor ( n49476 , n49473 , n49474 );
xor ( n49477 , n48896 , n49182 );
and ( n49478 , n30174 , n49282 );
and ( n49479 , n49477 , n49478 );
xor ( n49480 , n49477 , n49478 );
xor ( n49481 , n48900 , n49180 );
and ( n49482 , n30179 , n49282 );
and ( n49483 , n49481 , n49482 );
xor ( n49484 , n49481 , n49482 );
xor ( n49485 , n48904 , n49178 );
and ( n49486 , n30184 , n49282 );
and ( n49487 , n49485 , n49486 );
xor ( n49488 , n49485 , n49486 );
xor ( n49489 , n48908 , n49176 );
and ( n49490 , n30189 , n49282 );
and ( n49491 , n49489 , n49490 );
xor ( n49492 , n49489 , n49490 );
xor ( n49493 , n48912 , n49174 );
and ( n49494 , n30194 , n49282 );
and ( n49495 , n49493 , n49494 );
xor ( n49496 , n49493 , n49494 );
xor ( n49497 , n48916 , n49172 );
and ( n49498 , n30199 , n49282 );
and ( n49499 , n49497 , n49498 );
xor ( n49500 , n49497 , n49498 );
xor ( n49501 , n48920 , n49170 );
and ( n49502 , n30204 , n49282 );
and ( n49503 , n49501 , n49502 );
xor ( n49504 , n49501 , n49502 );
xor ( n49505 , n48924 , n49168 );
and ( n49506 , n30209 , n49282 );
and ( n49507 , n49505 , n49506 );
xor ( n49508 , n49505 , n49506 );
xor ( n49509 , n48928 , n49166 );
and ( n49510 , n30214 , n49282 );
and ( n49511 , n49509 , n49510 );
xor ( n49512 , n49509 , n49510 );
xor ( n49513 , n48932 , n49164 );
and ( n49514 , n30219 , n49282 );
and ( n49515 , n49513 , n49514 );
xor ( n49516 , n49513 , n49514 );
xor ( n49517 , n48936 , n49162 );
and ( n49518 , n30224 , n49282 );
and ( n49519 , n49517 , n49518 );
xor ( n49520 , n49517 , n49518 );
xor ( n49521 , n48940 , n49160 );
and ( n49522 , n30229 , n49282 );
and ( n49523 , n49521 , n49522 );
xor ( n49524 , n49521 , n49522 );
xor ( n49525 , n48944 , n49158 );
and ( n49526 , n30234 , n49282 );
and ( n49527 , n49525 , n49526 );
xor ( n49528 , n49525 , n49526 );
xor ( n49529 , n48948 , n49156 );
and ( n49530 , n30239 , n49282 );
and ( n49531 , n49529 , n49530 );
xor ( n49532 , n49529 , n49530 );
xor ( n49533 , n48952 , n49154 );
and ( n49534 , n30244 , n49282 );
and ( n49535 , n49533 , n49534 );
xor ( n49536 , n49533 , n49534 );
xor ( n49537 , n48956 , n49152 );
and ( n49538 , n30249 , n49282 );
and ( n49539 , n49537 , n49538 );
xor ( n49540 , n49537 , n49538 );
xor ( n49541 , n48960 , n49150 );
and ( n49542 , n30254 , n49282 );
and ( n49543 , n49541 , n49542 );
xor ( n49544 , n49541 , n49542 );
xor ( n49545 , n48964 , n49148 );
and ( n49546 , n30259 , n49282 );
and ( n49547 , n49545 , n49546 );
xor ( n49548 , n49545 , n49546 );
xor ( n49549 , n48968 , n49146 );
and ( n49550 , n30264 , n49282 );
and ( n49551 , n49549 , n49550 );
xor ( n49552 , n49549 , n49550 );
xor ( n49553 , n48972 , n49144 );
and ( n49554 , n30269 , n49282 );
and ( n49555 , n49553 , n49554 );
xor ( n49556 , n49553 , n49554 );
xor ( n49557 , n48976 , n49142 );
and ( n49558 , n30274 , n49282 );
and ( n49559 , n49557 , n49558 );
xor ( n49560 , n49557 , n49558 );
xor ( n49561 , n48980 , n49140 );
and ( n49562 , n30279 , n49282 );
and ( n49563 , n49561 , n49562 );
xor ( n49564 , n49561 , n49562 );
xor ( n49565 , n48984 , n49138 );
and ( n49566 , n30284 , n49282 );
and ( n49567 , n49565 , n49566 );
xor ( n49568 , n49565 , n49566 );
xor ( n49569 , n48988 , n49136 );
and ( n49570 , n30289 , n49282 );
and ( n49571 , n49569 , n49570 );
xor ( n49572 , n49569 , n49570 );
xor ( n49573 , n48992 , n49134 );
and ( n49574 , n30294 , n49282 );
and ( n49575 , n49573 , n49574 );
xor ( n49576 , n49573 , n49574 );
xor ( n49577 , n48996 , n49132 );
and ( n49578 , n30299 , n49282 );
and ( n49579 , n49577 , n49578 );
xor ( n49580 , n49577 , n49578 );
xor ( n49581 , n49000 , n49130 );
and ( n49582 , n30304 , n49282 );
and ( n49583 , n49581 , n49582 );
xor ( n49584 , n49581 , n49582 );
xor ( n49585 , n49004 , n49128 );
and ( n49586 , n30309 , n49282 );
and ( n49587 , n49585 , n49586 );
xor ( n49588 , n49585 , n49586 );
xor ( n49589 , n49008 , n49126 );
and ( n49590 , n30314 , n49282 );
and ( n49591 , n49589 , n49590 );
xor ( n49592 , n49589 , n49590 );
xor ( n49593 , n49012 , n49124 );
and ( n49594 , n30319 , n49282 );
and ( n49595 , n49593 , n49594 );
xor ( n49596 , n49593 , n49594 );
xor ( n49597 , n49016 , n49122 );
and ( n49598 , n30324 , n49282 );
and ( n49599 , n49597 , n49598 );
xor ( n49600 , n49597 , n49598 );
xor ( n49601 , n49020 , n49120 );
and ( n49602 , n30329 , n49282 );
and ( n49603 , n49601 , n49602 );
xor ( n49604 , n49601 , n49602 );
xor ( n49605 , n49024 , n49118 );
and ( n49606 , n30334 , n49282 );
and ( n49607 , n49605 , n49606 );
xor ( n49608 , n49605 , n49606 );
xor ( n49609 , n49028 , n49116 );
and ( n49610 , n30339 , n49282 );
and ( n49611 , n49609 , n49610 );
xor ( n49612 , n49609 , n49610 );
xor ( n49613 , n49032 , n49114 );
and ( n49614 , n30344 , n49282 );
and ( n49615 , n49613 , n49614 );
xor ( n49616 , n49613 , n49614 );
xor ( n49617 , n49036 , n49112 );
and ( n49618 , n30349 , n49282 );
and ( n49619 , n49617 , n49618 );
xor ( n49620 , n49617 , n49618 );
xor ( n49621 , n49040 , n49110 );
and ( n49622 , n30354 , n49282 );
and ( n49623 , n49621 , n49622 );
xor ( n49624 , n49621 , n49622 );
xor ( n49625 , n49044 , n49108 );
and ( n49626 , n30359 , n49282 );
and ( n49627 , n49625 , n49626 );
xor ( n49628 , n49625 , n49626 );
xor ( n49629 , n49048 , n49106 );
and ( n49630 , n30364 , n49282 );
and ( n49631 , n49629 , n49630 );
xor ( n49632 , n49629 , n49630 );
xor ( n49633 , n49052 , n49104 );
and ( n49634 , n30369 , n49282 );
and ( n49635 , n49633 , n49634 );
xor ( n49636 , n49633 , n49634 );
xor ( n49637 , n49056 , n49102 );
and ( n49638 , n30374 , n49282 );
and ( n49639 , n49637 , n49638 );
xor ( n49640 , n49637 , n49638 );
xor ( n49641 , n49060 , n49100 );
and ( n49642 , n30379 , n49282 );
and ( n49643 , n49641 , n49642 );
xor ( n49644 , n49641 , n49642 );
xor ( n49645 , n49064 , n49098 );
and ( n49646 , n30384 , n49282 );
and ( n49647 , n49645 , n49646 );
xor ( n49648 , n49645 , n49646 );
xor ( n49649 , n49068 , n49096 );
and ( n49650 , n30389 , n49282 );
and ( n49651 , n49649 , n49650 );
xor ( n49652 , n49649 , n49650 );
xor ( n49653 , n49072 , n49094 );
and ( n49654 , n30394 , n49282 );
and ( n49655 , n49653 , n49654 );
xor ( n49656 , n49653 , n49654 );
xor ( n49657 , n49076 , n49092 );
and ( n49658 , n30399 , n49282 );
and ( n49659 , n49657 , n49658 );
xor ( n49660 , n49657 , n49658 );
xor ( n49661 , n49080 , n49090 );
and ( n49662 , n30404 , n49282 );
and ( n49663 , n49661 , n49662 );
xor ( n49664 , n49661 , n49662 );
xor ( n49665 , n49084 , n49088 );
and ( n49666 , n30409 , n49282 );
and ( n49667 , n49665 , n49666 );
buf ( n49668 , n49667 );
and ( n49669 , n49664 , n49668 );
or ( n49670 , n49663 , n49669 );
and ( n49671 , n49660 , n49670 );
or ( n49672 , n49659 , n49671 );
and ( n49673 , n49656 , n49672 );
or ( n49674 , n49655 , n49673 );
and ( n49675 , n49652 , n49674 );
or ( n49676 , n49651 , n49675 );
and ( n49677 , n49648 , n49676 );
or ( n49678 , n49647 , n49677 );
and ( n49679 , n49644 , n49678 );
or ( n49680 , n49643 , n49679 );
and ( n49681 , n49640 , n49680 );
or ( n49682 , n49639 , n49681 );
and ( n49683 , n49636 , n49682 );
or ( n49684 , n49635 , n49683 );
and ( n49685 , n49632 , n49684 );
or ( n49686 , n49631 , n49685 );
and ( n49687 , n49628 , n49686 );
or ( n49688 , n49627 , n49687 );
and ( n49689 , n49624 , n49688 );
or ( n49690 , n49623 , n49689 );
and ( n49691 , n49620 , n49690 );
or ( n49692 , n49619 , n49691 );
and ( n49693 , n49616 , n49692 );
or ( n49694 , n49615 , n49693 );
and ( n49695 , n49612 , n49694 );
or ( n49696 , n49611 , n49695 );
and ( n49697 , n49608 , n49696 );
or ( n49698 , n49607 , n49697 );
and ( n49699 , n49604 , n49698 );
or ( n49700 , n49603 , n49699 );
and ( n49701 , n49600 , n49700 );
or ( n49702 , n49599 , n49701 );
and ( n49703 , n49596 , n49702 );
or ( n49704 , n49595 , n49703 );
and ( n49705 , n49592 , n49704 );
or ( n49706 , n49591 , n49705 );
and ( n49707 , n49588 , n49706 );
or ( n49708 , n49587 , n49707 );
and ( n49709 , n49584 , n49708 );
or ( n49710 , n49583 , n49709 );
and ( n49711 , n49580 , n49710 );
or ( n49712 , n49579 , n49711 );
and ( n49713 , n49576 , n49712 );
or ( n49714 , n49575 , n49713 );
and ( n49715 , n49572 , n49714 );
or ( n49716 , n49571 , n49715 );
and ( n49717 , n49568 , n49716 );
or ( n49718 , n49567 , n49717 );
and ( n49719 , n49564 , n49718 );
or ( n49720 , n49563 , n49719 );
and ( n49721 , n49560 , n49720 );
or ( n49722 , n49559 , n49721 );
and ( n49723 , n49556 , n49722 );
or ( n49724 , n49555 , n49723 );
and ( n49725 , n49552 , n49724 );
or ( n49726 , n49551 , n49725 );
and ( n49727 , n49548 , n49726 );
or ( n49728 , n49547 , n49727 );
and ( n49729 , n49544 , n49728 );
or ( n49730 , n49543 , n49729 );
and ( n49731 , n49540 , n49730 );
or ( n49732 , n49539 , n49731 );
and ( n49733 , n49536 , n49732 );
or ( n49734 , n49535 , n49733 );
and ( n49735 , n49532 , n49734 );
or ( n49736 , n49531 , n49735 );
and ( n49737 , n49528 , n49736 );
or ( n49738 , n49527 , n49737 );
and ( n49739 , n49524 , n49738 );
or ( n49740 , n49523 , n49739 );
and ( n49741 , n49520 , n49740 );
or ( n49742 , n49519 , n49741 );
and ( n49743 , n49516 , n49742 );
or ( n49744 , n49515 , n49743 );
and ( n49745 , n49512 , n49744 );
or ( n49746 , n49511 , n49745 );
and ( n49747 , n49508 , n49746 );
or ( n49748 , n49507 , n49747 );
and ( n49749 , n49504 , n49748 );
or ( n49750 , n49503 , n49749 );
and ( n49751 , n49500 , n49750 );
or ( n49752 , n49499 , n49751 );
and ( n49753 , n49496 , n49752 );
or ( n49754 , n49495 , n49753 );
and ( n49755 , n49492 , n49754 );
or ( n49756 , n49491 , n49755 );
and ( n49757 , n49488 , n49756 );
or ( n49758 , n49487 , n49757 );
and ( n49759 , n49484 , n49758 );
or ( n49760 , n49483 , n49759 );
and ( n49761 , n49480 , n49760 );
or ( n49762 , n49479 , n49761 );
and ( n49763 , n49476 , n49762 );
or ( n49764 , n49475 , n49763 );
and ( n49765 , n49472 , n49764 );
or ( n49766 , n49471 , n49765 );
and ( n49767 , n49468 , n49766 );
or ( n49768 , n49467 , n49767 );
and ( n49769 , n49464 , n49768 );
or ( n49770 , n49463 , n49769 );
and ( n49771 , n49460 , n49770 );
or ( n49772 , n49459 , n49771 );
and ( n49773 , n49456 , n49772 );
or ( n49774 , n49455 , n49773 );
and ( n49775 , n49452 , n49774 );
or ( n49776 , n49451 , n49775 );
and ( n49777 , n49448 , n49776 );
or ( n49778 , n49447 , n49777 );
and ( n49779 , n49444 , n49778 );
or ( n49780 , n49443 , n49779 );
and ( n49781 , n49440 , n49780 );
or ( n49782 , n49439 , n49781 );
and ( n49783 , n49436 , n49782 );
or ( n49784 , n49435 , n49783 );
and ( n49785 , n49432 , n49784 );
or ( n49786 , n49431 , n49785 );
and ( n49787 , n49428 , n49786 );
or ( n49788 , n49427 , n49787 );
and ( n49789 , n49424 , n49788 );
or ( n49790 , n49423 , n49789 );
and ( n49791 , n49420 , n49790 );
or ( n49792 , n49419 , n49791 );
and ( n49793 , n49416 , n49792 );
or ( n49794 , n49415 , n49793 );
and ( n49795 , n49412 , n49794 );
or ( n49796 , n49411 , n49795 );
and ( n49797 , n49408 , n49796 );
or ( n49798 , n49407 , n49797 );
and ( n49799 , n49404 , n49798 );
or ( n49800 , n49403 , n49799 );
and ( n49801 , n49400 , n49800 );
or ( n49802 , n49399 , n49801 );
and ( n49803 , n49396 , n49802 );
or ( n49804 , n49395 , n49803 );
and ( n49805 , n49392 , n49804 );
or ( n49806 , n49391 , n49805 );
and ( n49807 , n49388 , n49806 );
or ( n49808 , n49387 , n49807 );
and ( n49809 , n49384 , n49808 );
or ( n49810 , n49383 , n49809 );
and ( n49811 , n49380 , n49810 );
or ( n49812 , n49379 , n49811 );
and ( n49813 , n49376 , n49812 );
or ( n49814 , n49375 , n49813 );
and ( n49815 , n49372 , n49814 );
or ( n49816 , n49371 , n49815 );
and ( n49817 , n49368 , n49816 );
or ( n49818 , n49367 , n49817 );
and ( n49819 , n49364 , n49818 );
or ( n49820 , n49363 , n49819 );
and ( n49821 , n49360 , n49820 );
or ( n49822 , n49359 , n49821 );
and ( n49823 , n49356 , n49822 );
or ( n49824 , n49355 , n49823 );
and ( n49825 , n49352 , n49824 );
or ( n49826 , n49351 , n49825 );
and ( n49827 , n49348 , n49826 );
or ( n49828 , n49347 , n49827 );
and ( n49829 , n49344 , n49828 );
or ( n49830 , n49343 , n49829 );
and ( n49831 , n49340 , n49830 );
or ( n49832 , n49339 , n49831 );
and ( n49833 , n49336 , n49832 );
or ( n49834 , n49335 , n49833 );
and ( n49835 , n49332 , n49834 );
or ( n49836 , n49331 , n49835 );
and ( n49837 , n49328 , n49836 );
or ( n49838 , n49327 , n49837 );
and ( n49839 , n49324 , n49838 );
or ( n49840 , n49323 , n49839 );
and ( n49841 , n49320 , n49840 );
or ( n49842 , n49319 , n49841 );
and ( n49843 , n49316 , n49842 );
or ( n49844 , n49315 , n49843 );
and ( n49845 , n49312 , n49844 );
or ( n49846 , n49311 , n49845 );
and ( n49847 , n49308 , n49846 );
or ( n49848 , n49307 , n49847 );
and ( n49849 , n49304 , n49848 );
or ( n49850 , n49303 , n49849 );
and ( n49851 , n49300 , n49850 );
or ( n49852 , n49299 , n49851 );
and ( n49853 , n49296 , n49852 );
or ( n49854 , n49295 , n49853 );
and ( n49855 , n49292 , n49854 );
or ( n49856 , n49291 , n49855 );
and ( n49857 , n49288 , n49856 );
or ( n49858 , n49287 , n49857 );
xor ( n49859 , n49284 , n49858 );
buf ( n49860 , n18044 );
and ( n49861 , n29934 , n49860 );
xor ( n49862 , n49859 , n49861 );
xor ( n49863 , n49288 , n49856 );
and ( n49864 , n29939 , n49860 );
and ( n49865 , n49863 , n49864 );
xor ( n49866 , n49863 , n49864 );
xor ( n49867 , n49292 , n49854 );
and ( n49868 , n29944 , n49860 );
and ( n49869 , n49867 , n49868 );
xor ( n49870 , n49867 , n49868 );
xor ( n49871 , n49296 , n49852 );
and ( n49872 , n29949 , n49860 );
and ( n49873 , n49871 , n49872 );
xor ( n49874 , n49871 , n49872 );
xor ( n49875 , n49300 , n49850 );
and ( n49876 , n29954 , n49860 );
and ( n49877 , n49875 , n49876 );
xor ( n49878 , n49875 , n49876 );
xor ( n49879 , n49304 , n49848 );
and ( n49880 , n29959 , n49860 );
and ( n49881 , n49879 , n49880 );
xor ( n49882 , n49879 , n49880 );
xor ( n49883 , n49308 , n49846 );
and ( n49884 , n29964 , n49860 );
and ( n49885 , n49883 , n49884 );
xor ( n49886 , n49883 , n49884 );
xor ( n49887 , n49312 , n49844 );
and ( n49888 , n29969 , n49860 );
and ( n49889 , n49887 , n49888 );
xor ( n49890 , n49887 , n49888 );
xor ( n49891 , n49316 , n49842 );
and ( n49892 , n29974 , n49860 );
and ( n49893 , n49891 , n49892 );
xor ( n49894 , n49891 , n49892 );
xor ( n49895 , n49320 , n49840 );
and ( n49896 , n29979 , n49860 );
and ( n49897 , n49895 , n49896 );
xor ( n49898 , n49895 , n49896 );
xor ( n49899 , n49324 , n49838 );
and ( n49900 , n29984 , n49860 );
and ( n49901 , n49899 , n49900 );
xor ( n49902 , n49899 , n49900 );
xor ( n49903 , n49328 , n49836 );
and ( n49904 , n29989 , n49860 );
and ( n49905 , n49903 , n49904 );
xor ( n49906 , n49903 , n49904 );
xor ( n49907 , n49332 , n49834 );
and ( n49908 , n29994 , n49860 );
and ( n49909 , n49907 , n49908 );
xor ( n49910 , n49907 , n49908 );
xor ( n49911 , n49336 , n49832 );
and ( n49912 , n29999 , n49860 );
and ( n49913 , n49911 , n49912 );
xor ( n49914 , n49911 , n49912 );
xor ( n49915 , n49340 , n49830 );
and ( n49916 , n30004 , n49860 );
and ( n49917 , n49915 , n49916 );
xor ( n49918 , n49915 , n49916 );
xor ( n49919 , n49344 , n49828 );
and ( n49920 , n30009 , n49860 );
and ( n49921 , n49919 , n49920 );
xor ( n49922 , n49919 , n49920 );
xor ( n49923 , n49348 , n49826 );
and ( n49924 , n30014 , n49860 );
and ( n49925 , n49923 , n49924 );
xor ( n49926 , n49923 , n49924 );
xor ( n49927 , n49352 , n49824 );
and ( n49928 , n30019 , n49860 );
and ( n49929 , n49927 , n49928 );
xor ( n49930 , n49927 , n49928 );
xor ( n49931 , n49356 , n49822 );
and ( n49932 , n30024 , n49860 );
and ( n49933 , n49931 , n49932 );
xor ( n49934 , n49931 , n49932 );
xor ( n49935 , n49360 , n49820 );
and ( n49936 , n30029 , n49860 );
and ( n49937 , n49935 , n49936 );
xor ( n49938 , n49935 , n49936 );
xor ( n49939 , n49364 , n49818 );
and ( n49940 , n30034 , n49860 );
and ( n49941 , n49939 , n49940 );
xor ( n49942 , n49939 , n49940 );
xor ( n49943 , n49368 , n49816 );
and ( n49944 , n30039 , n49860 );
and ( n49945 , n49943 , n49944 );
xor ( n49946 , n49943 , n49944 );
xor ( n49947 , n49372 , n49814 );
and ( n49948 , n30044 , n49860 );
and ( n49949 , n49947 , n49948 );
xor ( n49950 , n49947 , n49948 );
xor ( n49951 , n49376 , n49812 );
and ( n49952 , n30049 , n49860 );
and ( n49953 , n49951 , n49952 );
xor ( n49954 , n49951 , n49952 );
xor ( n49955 , n49380 , n49810 );
and ( n49956 , n30054 , n49860 );
and ( n49957 , n49955 , n49956 );
xor ( n49958 , n49955 , n49956 );
xor ( n49959 , n49384 , n49808 );
and ( n49960 , n30059 , n49860 );
and ( n49961 , n49959 , n49960 );
xor ( n49962 , n49959 , n49960 );
xor ( n49963 , n49388 , n49806 );
and ( n49964 , n30064 , n49860 );
and ( n49965 , n49963 , n49964 );
xor ( n49966 , n49963 , n49964 );
xor ( n49967 , n49392 , n49804 );
and ( n49968 , n30069 , n49860 );
and ( n49969 , n49967 , n49968 );
xor ( n49970 , n49967 , n49968 );
xor ( n49971 , n49396 , n49802 );
and ( n49972 , n30074 , n49860 );
and ( n49973 , n49971 , n49972 );
xor ( n49974 , n49971 , n49972 );
xor ( n49975 , n49400 , n49800 );
and ( n49976 , n30079 , n49860 );
and ( n49977 , n49975 , n49976 );
xor ( n49978 , n49975 , n49976 );
xor ( n49979 , n49404 , n49798 );
and ( n49980 , n30084 , n49860 );
and ( n49981 , n49979 , n49980 );
xor ( n49982 , n49979 , n49980 );
xor ( n49983 , n49408 , n49796 );
and ( n49984 , n30089 , n49860 );
and ( n49985 , n49983 , n49984 );
xor ( n49986 , n49983 , n49984 );
xor ( n49987 , n49412 , n49794 );
and ( n49988 , n30094 , n49860 );
and ( n49989 , n49987 , n49988 );
xor ( n49990 , n49987 , n49988 );
xor ( n49991 , n49416 , n49792 );
and ( n49992 , n30099 , n49860 );
and ( n49993 , n49991 , n49992 );
xor ( n49994 , n49991 , n49992 );
xor ( n49995 , n49420 , n49790 );
and ( n49996 , n30104 , n49860 );
and ( n49997 , n49995 , n49996 );
xor ( n49998 , n49995 , n49996 );
xor ( n49999 , n49424 , n49788 );
and ( n50000 , n30109 , n49860 );
and ( n50001 , n49999 , n50000 );
xor ( n50002 , n49999 , n50000 );
xor ( n50003 , n49428 , n49786 );
and ( n50004 , n30114 , n49860 );
and ( n50005 , n50003 , n50004 );
xor ( n50006 , n50003 , n50004 );
xor ( n50007 , n49432 , n49784 );
and ( n50008 , n30119 , n49860 );
and ( n50009 , n50007 , n50008 );
xor ( n50010 , n50007 , n50008 );
xor ( n50011 , n49436 , n49782 );
and ( n50012 , n30124 , n49860 );
and ( n50013 , n50011 , n50012 );
xor ( n50014 , n50011 , n50012 );
xor ( n50015 , n49440 , n49780 );
and ( n50016 , n30129 , n49860 );
and ( n50017 , n50015 , n50016 );
xor ( n50018 , n50015 , n50016 );
xor ( n50019 , n49444 , n49778 );
and ( n50020 , n30134 , n49860 );
and ( n50021 , n50019 , n50020 );
xor ( n50022 , n50019 , n50020 );
xor ( n50023 , n49448 , n49776 );
and ( n50024 , n30139 , n49860 );
and ( n50025 , n50023 , n50024 );
xor ( n50026 , n50023 , n50024 );
xor ( n50027 , n49452 , n49774 );
and ( n50028 , n30144 , n49860 );
and ( n50029 , n50027 , n50028 );
xor ( n50030 , n50027 , n50028 );
xor ( n50031 , n49456 , n49772 );
and ( n50032 , n30149 , n49860 );
and ( n50033 , n50031 , n50032 );
xor ( n50034 , n50031 , n50032 );
xor ( n50035 , n49460 , n49770 );
and ( n50036 , n30154 , n49860 );
and ( n50037 , n50035 , n50036 );
xor ( n50038 , n50035 , n50036 );
xor ( n50039 , n49464 , n49768 );
and ( n50040 , n30159 , n49860 );
and ( n50041 , n50039 , n50040 );
xor ( n50042 , n50039 , n50040 );
xor ( n50043 , n49468 , n49766 );
and ( n50044 , n30164 , n49860 );
and ( n50045 , n50043 , n50044 );
xor ( n50046 , n50043 , n50044 );
xor ( n50047 , n49472 , n49764 );
and ( n50048 , n30169 , n49860 );
and ( n50049 , n50047 , n50048 );
xor ( n50050 , n50047 , n50048 );
xor ( n50051 , n49476 , n49762 );
and ( n50052 , n30174 , n49860 );
and ( n50053 , n50051 , n50052 );
xor ( n50054 , n50051 , n50052 );
xor ( n50055 , n49480 , n49760 );
and ( n50056 , n30179 , n49860 );
and ( n50057 , n50055 , n50056 );
xor ( n50058 , n50055 , n50056 );
xor ( n50059 , n49484 , n49758 );
and ( n50060 , n30184 , n49860 );
and ( n50061 , n50059 , n50060 );
xor ( n50062 , n50059 , n50060 );
xor ( n50063 , n49488 , n49756 );
and ( n50064 , n30189 , n49860 );
and ( n50065 , n50063 , n50064 );
xor ( n50066 , n50063 , n50064 );
xor ( n50067 , n49492 , n49754 );
and ( n50068 , n30194 , n49860 );
and ( n50069 , n50067 , n50068 );
xor ( n50070 , n50067 , n50068 );
xor ( n50071 , n49496 , n49752 );
and ( n50072 , n30199 , n49860 );
and ( n50073 , n50071 , n50072 );
xor ( n50074 , n50071 , n50072 );
xor ( n50075 , n49500 , n49750 );
and ( n50076 , n30204 , n49860 );
and ( n50077 , n50075 , n50076 );
xor ( n50078 , n50075 , n50076 );
xor ( n50079 , n49504 , n49748 );
and ( n50080 , n30209 , n49860 );
and ( n50081 , n50079 , n50080 );
xor ( n50082 , n50079 , n50080 );
xor ( n50083 , n49508 , n49746 );
and ( n50084 , n30214 , n49860 );
and ( n50085 , n50083 , n50084 );
xor ( n50086 , n50083 , n50084 );
xor ( n50087 , n49512 , n49744 );
and ( n50088 , n30219 , n49860 );
and ( n50089 , n50087 , n50088 );
xor ( n50090 , n50087 , n50088 );
xor ( n50091 , n49516 , n49742 );
and ( n50092 , n30224 , n49860 );
and ( n50093 , n50091 , n50092 );
xor ( n50094 , n50091 , n50092 );
xor ( n50095 , n49520 , n49740 );
and ( n50096 , n30229 , n49860 );
and ( n50097 , n50095 , n50096 );
xor ( n50098 , n50095 , n50096 );
xor ( n50099 , n49524 , n49738 );
and ( n50100 , n30234 , n49860 );
and ( n50101 , n50099 , n50100 );
xor ( n50102 , n50099 , n50100 );
xor ( n50103 , n49528 , n49736 );
and ( n50104 , n30239 , n49860 );
and ( n50105 , n50103 , n50104 );
xor ( n50106 , n50103 , n50104 );
xor ( n50107 , n49532 , n49734 );
and ( n50108 , n30244 , n49860 );
and ( n50109 , n50107 , n50108 );
xor ( n50110 , n50107 , n50108 );
xor ( n50111 , n49536 , n49732 );
and ( n50112 , n30249 , n49860 );
and ( n50113 , n50111 , n50112 );
xor ( n50114 , n50111 , n50112 );
xor ( n50115 , n49540 , n49730 );
and ( n50116 , n30254 , n49860 );
and ( n50117 , n50115 , n50116 );
xor ( n50118 , n50115 , n50116 );
xor ( n50119 , n49544 , n49728 );
and ( n50120 , n30259 , n49860 );
and ( n50121 , n50119 , n50120 );
xor ( n50122 , n50119 , n50120 );
xor ( n50123 , n49548 , n49726 );
and ( n50124 , n30264 , n49860 );
and ( n50125 , n50123 , n50124 );
xor ( n50126 , n50123 , n50124 );
xor ( n50127 , n49552 , n49724 );
and ( n50128 , n30269 , n49860 );
and ( n50129 , n50127 , n50128 );
xor ( n50130 , n50127 , n50128 );
xor ( n50131 , n49556 , n49722 );
and ( n50132 , n30274 , n49860 );
and ( n50133 , n50131 , n50132 );
xor ( n50134 , n50131 , n50132 );
xor ( n50135 , n49560 , n49720 );
and ( n50136 , n30279 , n49860 );
and ( n50137 , n50135 , n50136 );
xor ( n50138 , n50135 , n50136 );
xor ( n50139 , n49564 , n49718 );
and ( n50140 , n30284 , n49860 );
and ( n50141 , n50139 , n50140 );
xor ( n50142 , n50139 , n50140 );
xor ( n50143 , n49568 , n49716 );
and ( n50144 , n30289 , n49860 );
and ( n50145 , n50143 , n50144 );
xor ( n50146 , n50143 , n50144 );
xor ( n50147 , n49572 , n49714 );
and ( n50148 , n30294 , n49860 );
and ( n50149 , n50147 , n50148 );
xor ( n50150 , n50147 , n50148 );
xor ( n50151 , n49576 , n49712 );
and ( n50152 , n30299 , n49860 );
and ( n50153 , n50151 , n50152 );
xor ( n50154 , n50151 , n50152 );
xor ( n50155 , n49580 , n49710 );
and ( n50156 , n30304 , n49860 );
and ( n50157 , n50155 , n50156 );
xor ( n50158 , n50155 , n50156 );
xor ( n50159 , n49584 , n49708 );
and ( n50160 , n30309 , n49860 );
and ( n50161 , n50159 , n50160 );
xor ( n50162 , n50159 , n50160 );
xor ( n50163 , n49588 , n49706 );
and ( n50164 , n30314 , n49860 );
and ( n50165 , n50163 , n50164 );
xor ( n50166 , n50163 , n50164 );
xor ( n50167 , n49592 , n49704 );
and ( n50168 , n30319 , n49860 );
and ( n50169 , n50167 , n50168 );
xor ( n50170 , n50167 , n50168 );
xor ( n50171 , n49596 , n49702 );
and ( n50172 , n30324 , n49860 );
and ( n50173 , n50171 , n50172 );
xor ( n50174 , n50171 , n50172 );
xor ( n50175 , n49600 , n49700 );
and ( n50176 , n30329 , n49860 );
and ( n50177 , n50175 , n50176 );
xor ( n50178 , n50175 , n50176 );
xor ( n50179 , n49604 , n49698 );
and ( n50180 , n30334 , n49860 );
and ( n50181 , n50179 , n50180 );
xor ( n50182 , n50179 , n50180 );
xor ( n50183 , n49608 , n49696 );
and ( n50184 , n30339 , n49860 );
and ( n50185 , n50183 , n50184 );
xor ( n50186 , n50183 , n50184 );
xor ( n50187 , n49612 , n49694 );
and ( n50188 , n30344 , n49860 );
and ( n50189 , n50187 , n50188 );
xor ( n50190 , n50187 , n50188 );
xor ( n50191 , n49616 , n49692 );
and ( n50192 , n30349 , n49860 );
and ( n50193 , n50191 , n50192 );
xor ( n50194 , n50191 , n50192 );
xor ( n50195 , n49620 , n49690 );
and ( n50196 , n30354 , n49860 );
and ( n50197 , n50195 , n50196 );
xor ( n50198 , n50195 , n50196 );
xor ( n50199 , n49624 , n49688 );
and ( n50200 , n30359 , n49860 );
and ( n50201 , n50199 , n50200 );
xor ( n50202 , n50199 , n50200 );
xor ( n50203 , n49628 , n49686 );
and ( n50204 , n30364 , n49860 );
and ( n50205 , n50203 , n50204 );
xor ( n50206 , n50203 , n50204 );
xor ( n50207 , n49632 , n49684 );
and ( n50208 , n30369 , n49860 );
and ( n50209 , n50207 , n50208 );
xor ( n50210 , n50207 , n50208 );
xor ( n50211 , n49636 , n49682 );
and ( n50212 , n30374 , n49860 );
and ( n50213 , n50211 , n50212 );
xor ( n50214 , n50211 , n50212 );
xor ( n50215 , n49640 , n49680 );
and ( n50216 , n30379 , n49860 );
and ( n50217 , n50215 , n50216 );
xor ( n50218 , n50215 , n50216 );
xor ( n50219 , n49644 , n49678 );
and ( n50220 , n30384 , n49860 );
and ( n50221 , n50219 , n50220 );
xor ( n50222 , n50219 , n50220 );
xor ( n50223 , n49648 , n49676 );
and ( n50224 , n30389 , n49860 );
and ( n50225 , n50223 , n50224 );
xor ( n50226 , n50223 , n50224 );
xor ( n50227 , n49652 , n49674 );
and ( n50228 , n30394 , n49860 );
and ( n50229 , n50227 , n50228 );
xor ( n50230 , n50227 , n50228 );
xor ( n50231 , n49656 , n49672 );
and ( n50232 , n30399 , n49860 );
and ( n50233 , n50231 , n50232 );
xor ( n50234 , n50231 , n50232 );
xor ( n50235 , n49660 , n49670 );
and ( n50236 , n30404 , n49860 );
and ( n50237 , n50235 , n50236 );
xor ( n50238 , n50235 , n50236 );
xor ( n50239 , n49664 , n49668 );
and ( n50240 , n30409 , n49860 );
and ( n50241 , n50239 , n50240 );
buf ( n50242 , n50241 );
and ( n50243 , n50238 , n50242 );
or ( n50244 , n50237 , n50243 );
and ( n50245 , n50234 , n50244 );
or ( n50246 , n50233 , n50245 );
and ( n50247 , n50230 , n50246 );
or ( n50248 , n50229 , n50247 );
and ( n50249 , n50226 , n50248 );
or ( n50250 , n50225 , n50249 );
and ( n50251 , n50222 , n50250 );
or ( n50252 , n50221 , n50251 );
and ( n50253 , n50218 , n50252 );
or ( n50254 , n50217 , n50253 );
and ( n50255 , n50214 , n50254 );
or ( n50256 , n50213 , n50255 );
and ( n50257 , n50210 , n50256 );
or ( n50258 , n50209 , n50257 );
and ( n50259 , n50206 , n50258 );
or ( n50260 , n50205 , n50259 );
and ( n50261 , n50202 , n50260 );
or ( n50262 , n50201 , n50261 );
and ( n50263 , n50198 , n50262 );
or ( n50264 , n50197 , n50263 );
and ( n50265 , n50194 , n50264 );
or ( n50266 , n50193 , n50265 );
and ( n50267 , n50190 , n50266 );
or ( n50268 , n50189 , n50267 );
and ( n50269 , n50186 , n50268 );
or ( n50270 , n50185 , n50269 );
and ( n50271 , n50182 , n50270 );
or ( n50272 , n50181 , n50271 );
and ( n50273 , n50178 , n50272 );
or ( n50274 , n50177 , n50273 );
and ( n50275 , n50174 , n50274 );
or ( n50276 , n50173 , n50275 );
and ( n50277 , n50170 , n50276 );
or ( n50278 , n50169 , n50277 );
and ( n50279 , n50166 , n50278 );
or ( n50280 , n50165 , n50279 );
and ( n50281 , n50162 , n50280 );
or ( n50282 , n50161 , n50281 );
and ( n50283 , n50158 , n50282 );
or ( n50284 , n50157 , n50283 );
and ( n50285 , n50154 , n50284 );
or ( n50286 , n50153 , n50285 );
and ( n50287 , n50150 , n50286 );
or ( n50288 , n50149 , n50287 );
and ( n50289 , n50146 , n50288 );
or ( n50290 , n50145 , n50289 );
and ( n50291 , n50142 , n50290 );
or ( n50292 , n50141 , n50291 );
and ( n50293 , n50138 , n50292 );
or ( n50294 , n50137 , n50293 );
and ( n50295 , n50134 , n50294 );
or ( n50296 , n50133 , n50295 );
and ( n50297 , n50130 , n50296 );
or ( n50298 , n50129 , n50297 );
and ( n50299 , n50126 , n50298 );
or ( n50300 , n50125 , n50299 );
and ( n50301 , n50122 , n50300 );
or ( n50302 , n50121 , n50301 );
and ( n50303 , n50118 , n50302 );
or ( n50304 , n50117 , n50303 );
and ( n50305 , n50114 , n50304 );
or ( n50306 , n50113 , n50305 );
and ( n50307 , n50110 , n50306 );
or ( n50308 , n50109 , n50307 );
and ( n50309 , n50106 , n50308 );
or ( n50310 , n50105 , n50309 );
and ( n50311 , n50102 , n50310 );
or ( n50312 , n50101 , n50311 );
and ( n50313 , n50098 , n50312 );
or ( n50314 , n50097 , n50313 );
and ( n50315 , n50094 , n50314 );
or ( n50316 , n50093 , n50315 );
and ( n50317 , n50090 , n50316 );
or ( n50318 , n50089 , n50317 );
and ( n50319 , n50086 , n50318 );
or ( n50320 , n50085 , n50319 );
and ( n50321 , n50082 , n50320 );
or ( n50322 , n50081 , n50321 );
and ( n50323 , n50078 , n50322 );
or ( n50324 , n50077 , n50323 );
and ( n50325 , n50074 , n50324 );
or ( n50326 , n50073 , n50325 );
and ( n50327 , n50070 , n50326 );
or ( n50328 , n50069 , n50327 );
and ( n50329 , n50066 , n50328 );
or ( n50330 , n50065 , n50329 );
and ( n50331 , n50062 , n50330 );
or ( n50332 , n50061 , n50331 );
and ( n50333 , n50058 , n50332 );
or ( n50334 , n50057 , n50333 );
and ( n50335 , n50054 , n50334 );
or ( n50336 , n50053 , n50335 );
and ( n50337 , n50050 , n50336 );
or ( n50338 , n50049 , n50337 );
and ( n50339 , n50046 , n50338 );
or ( n50340 , n50045 , n50339 );
and ( n50341 , n50042 , n50340 );
or ( n50342 , n50041 , n50341 );
and ( n50343 , n50038 , n50342 );
or ( n50344 , n50037 , n50343 );
and ( n50345 , n50034 , n50344 );
or ( n50346 , n50033 , n50345 );
and ( n50347 , n50030 , n50346 );
or ( n50348 , n50029 , n50347 );
and ( n50349 , n50026 , n50348 );
or ( n50350 , n50025 , n50349 );
and ( n50351 , n50022 , n50350 );
or ( n50352 , n50021 , n50351 );
and ( n50353 , n50018 , n50352 );
or ( n50354 , n50017 , n50353 );
and ( n50355 , n50014 , n50354 );
or ( n50356 , n50013 , n50355 );
and ( n50357 , n50010 , n50356 );
or ( n50358 , n50009 , n50357 );
and ( n50359 , n50006 , n50358 );
or ( n50360 , n50005 , n50359 );
and ( n50361 , n50002 , n50360 );
or ( n50362 , n50001 , n50361 );
and ( n50363 , n49998 , n50362 );
or ( n50364 , n49997 , n50363 );
and ( n50365 , n49994 , n50364 );
or ( n50366 , n49993 , n50365 );
and ( n50367 , n49990 , n50366 );
or ( n50368 , n49989 , n50367 );
and ( n50369 , n49986 , n50368 );
or ( n50370 , n49985 , n50369 );
and ( n50371 , n49982 , n50370 );
or ( n50372 , n49981 , n50371 );
and ( n50373 , n49978 , n50372 );
or ( n50374 , n49977 , n50373 );
and ( n50375 , n49974 , n50374 );
or ( n50376 , n49973 , n50375 );
and ( n50377 , n49970 , n50376 );
or ( n50378 , n49969 , n50377 );
and ( n50379 , n49966 , n50378 );
or ( n50380 , n49965 , n50379 );
and ( n50381 , n49962 , n50380 );
or ( n50382 , n49961 , n50381 );
and ( n50383 , n49958 , n50382 );
or ( n50384 , n49957 , n50383 );
and ( n50385 , n49954 , n50384 );
or ( n50386 , n49953 , n50385 );
and ( n50387 , n49950 , n50386 );
or ( n50388 , n49949 , n50387 );
and ( n50389 , n49946 , n50388 );
or ( n50390 , n49945 , n50389 );
and ( n50391 , n49942 , n50390 );
or ( n50392 , n49941 , n50391 );
and ( n50393 , n49938 , n50392 );
or ( n50394 , n49937 , n50393 );
and ( n50395 , n49934 , n50394 );
or ( n50396 , n49933 , n50395 );
and ( n50397 , n49930 , n50396 );
or ( n50398 , n49929 , n50397 );
and ( n50399 , n49926 , n50398 );
or ( n50400 , n49925 , n50399 );
and ( n50401 , n49922 , n50400 );
or ( n50402 , n49921 , n50401 );
and ( n50403 , n49918 , n50402 );
or ( n50404 , n49917 , n50403 );
and ( n50405 , n49914 , n50404 );
or ( n50406 , n49913 , n50405 );
and ( n50407 , n49910 , n50406 );
or ( n50408 , n49909 , n50407 );
and ( n50409 , n49906 , n50408 );
or ( n50410 , n49905 , n50409 );
and ( n50411 , n49902 , n50410 );
or ( n50412 , n49901 , n50411 );
and ( n50413 , n49898 , n50412 );
or ( n50414 , n49897 , n50413 );
and ( n50415 , n49894 , n50414 );
or ( n50416 , n49893 , n50415 );
and ( n50417 , n49890 , n50416 );
or ( n50418 , n49889 , n50417 );
and ( n50419 , n49886 , n50418 );
or ( n50420 , n49885 , n50419 );
and ( n50421 , n49882 , n50420 );
or ( n50422 , n49881 , n50421 );
and ( n50423 , n49878 , n50422 );
or ( n50424 , n49877 , n50423 );
and ( n50425 , n49874 , n50424 );
or ( n50426 , n49873 , n50425 );
and ( n50427 , n49870 , n50426 );
or ( n50428 , n49869 , n50427 );
and ( n50429 , n49866 , n50428 );
or ( n50430 , n49865 , n50429 );
xor ( n50431 , n49862 , n50430 );
buf ( n50432 , n18042 );
and ( n50433 , n29939 , n50432 );
xor ( n50434 , n50431 , n50433 );
xor ( n50435 , n49866 , n50428 );
and ( n50436 , n29944 , n50432 );
and ( n50437 , n50435 , n50436 );
xor ( n50438 , n50435 , n50436 );
xor ( n50439 , n49870 , n50426 );
and ( n50440 , n29949 , n50432 );
and ( n50441 , n50439 , n50440 );
xor ( n50442 , n50439 , n50440 );
xor ( n50443 , n49874 , n50424 );
and ( n50444 , n29954 , n50432 );
and ( n50445 , n50443 , n50444 );
xor ( n50446 , n50443 , n50444 );
xor ( n50447 , n49878 , n50422 );
and ( n50448 , n29959 , n50432 );
and ( n50449 , n50447 , n50448 );
xor ( n50450 , n50447 , n50448 );
xor ( n50451 , n49882 , n50420 );
and ( n50452 , n29964 , n50432 );
and ( n50453 , n50451 , n50452 );
xor ( n50454 , n50451 , n50452 );
xor ( n50455 , n49886 , n50418 );
and ( n50456 , n29969 , n50432 );
and ( n50457 , n50455 , n50456 );
xor ( n50458 , n50455 , n50456 );
xor ( n50459 , n49890 , n50416 );
and ( n50460 , n29974 , n50432 );
and ( n50461 , n50459 , n50460 );
xor ( n50462 , n50459 , n50460 );
xor ( n50463 , n49894 , n50414 );
and ( n50464 , n29979 , n50432 );
and ( n50465 , n50463 , n50464 );
xor ( n50466 , n50463 , n50464 );
xor ( n50467 , n49898 , n50412 );
and ( n50468 , n29984 , n50432 );
and ( n50469 , n50467 , n50468 );
xor ( n50470 , n50467 , n50468 );
xor ( n50471 , n49902 , n50410 );
and ( n50472 , n29989 , n50432 );
and ( n50473 , n50471 , n50472 );
xor ( n50474 , n50471 , n50472 );
xor ( n50475 , n49906 , n50408 );
and ( n50476 , n29994 , n50432 );
and ( n50477 , n50475 , n50476 );
xor ( n50478 , n50475 , n50476 );
xor ( n50479 , n49910 , n50406 );
and ( n50480 , n29999 , n50432 );
and ( n50481 , n50479 , n50480 );
xor ( n50482 , n50479 , n50480 );
xor ( n50483 , n49914 , n50404 );
and ( n50484 , n30004 , n50432 );
and ( n50485 , n50483 , n50484 );
xor ( n50486 , n50483 , n50484 );
xor ( n50487 , n49918 , n50402 );
and ( n50488 , n30009 , n50432 );
and ( n50489 , n50487 , n50488 );
xor ( n50490 , n50487 , n50488 );
xor ( n50491 , n49922 , n50400 );
and ( n50492 , n30014 , n50432 );
and ( n50493 , n50491 , n50492 );
xor ( n50494 , n50491 , n50492 );
xor ( n50495 , n49926 , n50398 );
and ( n50496 , n30019 , n50432 );
and ( n50497 , n50495 , n50496 );
xor ( n50498 , n50495 , n50496 );
xor ( n50499 , n49930 , n50396 );
and ( n50500 , n30024 , n50432 );
and ( n50501 , n50499 , n50500 );
xor ( n50502 , n50499 , n50500 );
xor ( n50503 , n49934 , n50394 );
and ( n50504 , n30029 , n50432 );
and ( n50505 , n50503 , n50504 );
xor ( n50506 , n50503 , n50504 );
xor ( n50507 , n49938 , n50392 );
and ( n50508 , n30034 , n50432 );
and ( n50509 , n50507 , n50508 );
xor ( n50510 , n50507 , n50508 );
xor ( n50511 , n49942 , n50390 );
and ( n50512 , n30039 , n50432 );
and ( n50513 , n50511 , n50512 );
xor ( n50514 , n50511 , n50512 );
xor ( n50515 , n49946 , n50388 );
and ( n50516 , n30044 , n50432 );
and ( n50517 , n50515 , n50516 );
xor ( n50518 , n50515 , n50516 );
xor ( n50519 , n49950 , n50386 );
and ( n50520 , n30049 , n50432 );
and ( n50521 , n50519 , n50520 );
xor ( n50522 , n50519 , n50520 );
xor ( n50523 , n49954 , n50384 );
and ( n50524 , n30054 , n50432 );
and ( n50525 , n50523 , n50524 );
xor ( n50526 , n50523 , n50524 );
xor ( n50527 , n49958 , n50382 );
and ( n50528 , n30059 , n50432 );
and ( n50529 , n50527 , n50528 );
xor ( n50530 , n50527 , n50528 );
xor ( n50531 , n49962 , n50380 );
and ( n50532 , n30064 , n50432 );
and ( n50533 , n50531 , n50532 );
xor ( n50534 , n50531 , n50532 );
xor ( n50535 , n49966 , n50378 );
and ( n50536 , n30069 , n50432 );
and ( n50537 , n50535 , n50536 );
xor ( n50538 , n50535 , n50536 );
xor ( n50539 , n49970 , n50376 );
and ( n50540 , n30074 , n50432 );
and ( n50541 , n50539 , n50540 );
xor ( n50542 , n50539 , n50540 );
xor ( n50543 , n49974 , n50374 );
and ( n50544 , n30079 , n50432 );
and ( n50545 , n50543 , n50544 );
xor ( n50546 , n50543 , n50544 );
xor ( n50547 , n49978 , n50372 );
and ( n50548 , n30084 , n50432 );
and ( n50549 , n50547 , n50548 );
xor ( n50550 , n50547 , n50548 );
xor ( n50551 , n49982 , n50370 );
and ( n50552 , n30089 , n50432 );
and ( n50553 , n50551 , n50552 );
xor ( n50554 , n50551 , n50552 );
xor ( n50555 , n49986 , n50368 );
and ( n50556 , n30094 , n50432 );
and ( n50557 , n50555 , n50556 );
xor ( n50558 , n50555 , n50556 );
xor ( n50559 , n49990 , n50366 );
and ( n50560 , n30099 , n50432 );
and ( n50561 , n50559 , n50560 );
xor ( n50562 , n50559 , n50560 );
xor ( n50563 , n49994 , n50364 );
and ( n50564 , n30104 , n50432 );
and ( n50565 , n50563 , n50564 );
xor ( n50566 , n50563 , n50564 );
xor ( n50567 , n49998 , n50362 );
and ( n50568 , n30109 , n50432 );
and ( n50569 , n50567 , n50568 );
xor ( n50570 , n50567 , n50568 );
xor ( n50571 , n50002 , n50360 );
and ( n50572 , n30114 , n50432 );
and ( n50573 , n50571 , n50572 );
xor ( n50574 , n50571 , n50572 );
xor ( n50575 , n50006 , n50358 );
and ( n50576 , n30119 , n50432 );
and ( n50577 , n50575 , n50576 );
xor ( n50578 , n50575 , n50576 );
xor ( n50579 , n50010 , n50356 );
and ( n50580 , n30124 , n50432 );
and ( n50581 , n50579 , n50580 );
xor ( n50582 , n50579 , n50580 );
xor ( n50583 , n50014 , n50354 );
and ( n50584 , n30129 , n50432 );
and ( n50585 , n50583 , n50584 );
xor ( n50586 , n50583 , n50584 );
xor ( n50587 , n50018 , n50352 );
and ( n50588 , n30134 , n50432 );
and ( n50589 , n50587 , n50588 );
xor ( n50590 , n50587 , n50588 );
xor ( n50591 , n50022 , n50350 );
and ( n50592 , n30139 , n50432 );
and ( n50593 , n50591 , n50592 );
xor ( n50594 , n50591 , n50592 );
xor ( n50595 , n50026 , n50348 );
and ( n50596 , n30144 , n50432 );
and ( n50597 , n50595 , n50596 );
xor ( n50598 , n50595 , n50596 );
xor ( n50599 , n50030 , n50346 );
and ( n50600 , n30149 , n50432 );
and ( n50601 , n50599 , n50600 );
xor ( n50602 , n50599 , n50600 );
xor ( n50603 , n50034 , n50344 );
and ( n50604 , n30154 , n50432 );
and ( n50605 , n50603 , n50604 );
xor ( n50606 , n50603 , n50604 );
xor ( n50607 , n50038 , n50342 );
and ( n50608 , n30159 , n50432 );
and ( n50609 , n50607 , n50608 );
xor ( n50610 , n50607 , n50608 );
xor ( n50611 , n50042 , n50340 );
and ( n50612 , n30164 , n50432 );
and ( n50613 , n50611 , n50612 );
xor ( n50614 , n50611 , n50612 );
xor ( n50615 , n50046 , n50338 );
and ( n50616 , n30169 , n50432 );
and ( n50617 , n50615 , n50616 );
xor ( n50618 , n50615 , n50616 );
xor ( n50619 , n50050 , n50336 );
and ( n50620 , n30174 , n50432 );
and ( n50621 , n50619 , n50620 );
xor ( n50622 , n50619 , n50620 );
xor ( n50623 , n50054 , n50334 );
and ( n50624 , n30179 , n50432 );
and ( n50625 , n50623 , n50624 );
xor ( n50626 , n50623 , n50624 );
xor ( n50627 , n50058 , n50332 );
and ( n50628 , n30184 , n50432 );
and ( n50629 , n50627 , n50628 );
xor ( n50630 , n50627 , n50628 );
xor ( n50631 , n50062 , n50330 );
and ( n50632 , n30189 , n50432 );
and ( n50633 , n50631 , n50632 );
xor ( n50634 , n50631 , n50632 );
xor ( n50635 , n50066 , n50328 );
and ( n50636 , n30194 , n50432 );
and ( n50637 , n50635 , n50636 );
xor ( n50638 , n50635 , n50636 );
xor ( n50639 , n50070 , n50326 );
and ( n50640 , n30199 , n50432 );
and ( n50641 , n50639 , n50640 );
xor ( n50642 , n50639 , n50640 );
xor ( n50643 , n50074 , n50324 );
and ( n50644 , n30204 , n50432 );
and ( n50645 , n50643 , n50644 );
xor ( n50646 , n50643 , n50644 );
xor ( n50647 , n50078 , n50322 );
and ( n50648 , n30209 , n50432 );
and ( n50649 , n50647 , n50648 );
xor ( n50650 , n50647 , n50648 );
xor ( n50651 , n50082 , n50320 );
and ( n50652 , n30214 , n50432 );
and ( n50653 , n50651 , n50652 );
xor ( n50654 , n50651 , n50652 );
xor ( n50655 , n50086 , n50318 );
and ( n50656 , n30219 , n50432 );
and ( n50657 , n50655 , n50656 );
xor ( n50658 , n50655 , n50656 );
xor ( n50659 , n50090 , n50316 );
and ( n50660 , n30224 , n50432 );
and ( n50661 , n50659 , n50660 );
xor ( n50662 , n50659 , n50660 );
xor ( n50663 , n50094 , n50314 );
and ( n50664 , n30229 , n50432 );
and ( n50665 , n50663 , n50664 );
xor ( n50666 , n50663 , n50664 );
xor ( n50667 , n50098 , n50312 );
and ( n50668 , n30234 , n50432 );
and ( n50669 , n50667 , n50668 );
xor ( n50670 , n50667 , n50668 );
xor ( n50671 , n50102 , n50310 );
and ( n50672 , n30239 , n50432 );
and ( n50673 , n50671 , n50672 );
xor ( n50674 , n50671 , n50672 );
xor ( n50675 , n50106 , n50308 );
and ( n50676 , n30244 , n50432 );
and ( n50677 , n50675 , n50676 );
xor ( n50678 , n50675 , n50676 );
xor ( n50679 , n50110 , n50306 );
and ( n50680 , n30249 , n50432 );
and ( n50681 , n50679 , n50680 );
xor ( n50682 , n50679 , n50680 );
xor ( n50683 , n50114 , n50304 );
and ( n50684 , n30254 , n50432 );
and ( n50685 , n50683 , n50684 );
xor ( n50686 , n50683 , n50684 );
xor ( n50687 , n50118 , n50302 );
and ( n50688 , n30259 , n50432 );
and ( n50689 , n50687 , n50688 );
xor ( n50690 , n50687 , n50688 );
xor ( n50691 , n50122 , n50300 );
and ( n50692 , n30264 , n50432 );
and ( n50693 , n50691 , n50692 );
xor ( n50694 , n50691 , n50692 );
xor ( n50695 , n50126 , n50298 );
and ( n50696 , n30269 , n50432 );
and ( n50697 , n50695 , n50696 );
xor ( n50698 , n50695 , n50696 );
xor ( n50699 , n50130 , n50296 );
and ( n50700 , n30274 , n50432 );
and ( n50701 , n50699 , n50700 );
xor ( n50702 , n50699 , n50700 );
xor ( n50703 , n50134 , n50294 );
and ( n50704 , n30279 , n50432 );
and ( n50705 , n50703 , n50704 );
xor ( n50706 , n50703 , n50704 );
xor ( n50707 , n50138 , n50292 );
and ( n50708 , n30284 , n50432 );
and ( n50709 , n50707 , n50708 );
xor ( n50710 , n50707 , n50708 );
xor ( n50711 , n50142 , n50290 );
and ( n50712 , n30289 , n50432 );
and ( n50713 , n50711 , n50712 );
xor ( n50714 , n50711 , n50712 );
xor ( n50715 , n50146 , n50288 );
and ( n50716 , n30294 , n50432 );
and ( n50717 , n50715 , n50716 );
xor ( n50718 , n50715 , n50716 );
xor ( n50719 , n50150 , n50286 );
and ( n50720 , n30299 , n50432 );
and ( n50721 , n50719 , n50720 );
xor ( n50722 , n50719 , n50720 );
xor ( n50723 , n50154 , n50284 );
and ( n50724 , n30304 , n50432 );
and ( n50725 , n50723 , n50724 );
xor ( n50726 , n50723 , n50724 );
xor ( n50727 , n50158 , n50282 );
and ( n50728 , n30309 , n50432 );
and ( n50729 , n50727 , n50728 );
xor ( n50730 , n50727 , n50728 );
xor ( n50731 , n50162 , n50280 );
and ( n50732 , n30314 , n50432 );
and ( n50733 , n50731 , n50732 );
xor ( n50734 , n50731 , n50732 );
xor ( n50735 , n50166 , n50278 );
and ( n50736 , n30319 , n50432 );
and ( n50737 , n50735 , n50736 );
xor ( n50738 , n50735 , n50736 );
xor ( n50739 , n50170 , n50276 );
and ( n50740 , n30324 , n50432 );
and ( n50741 , n50739 , n50740 );
xor ( n50742 , n50739 , n50740 );
xor ( n50743 , n50174 , n50274 );
and ( n50744 , n30329 , n50432 );
and ( n50745 , n50743 , n50744 );
xor ( n50746 , n50743 , n50744 );
xor ( n50747 , n50178 , n50272 );
and ( n50748 , n30334 , n50432 );
and ( n50749 , n50747 , n50748 );
xor ( n50750 , n50747 , n50748 );
xor ( n50751 , n50182 , n50270 );
and ( n50752 , n30339 , n50432 );
and ( n50753 , n50751 , n50752 );
xor ( n50754 , n50751 , n50752 );
xor ( n50755 , n50186 , n50268 );
and ( n50756 , n30344 , n50432 );
and ( n50757 , n50755 , n50756 );
xor ( n50758 , n50755 , n50756 );
xor ( n50759 , n50190 , n50266 );
and ( n50760 , n30349 , n50432 );
and ( n50761 , n50759 , n50760 );
xor ( n50762 , n50759 , n50760 );
xor ( n50763 , n50194 , n50264 );
and ( n50764 , n30354 , n50432 );
and ( n50765 , n50763 , n50764 );
xor ( n50766 , n50763 , n50764 );
xor ( n50767 , n50198 , n50262 );
and ( n50768 , n30359 , n50432 );
and ( n50769 , n50767 , n50768 );
xor ( n50770 , n50767 , n50768 );
xor ( n50771 , n50202 , n50260 );
and ( n50772 , n30364 , n50432 );
and ( n50773 , n50771 , n50772 );
xor ( n50774 , n50771 , n50772 );
xor ( n50775 , n50206 , n50258 );
and ( n50776 , n30369 , n50432 );
and ( n50777 , n50775 , n50776 );
xor ( n50778 , n50775 , n50776 );
xor ( n50779 , n50210 , n50256 );
and ( n50780 , n30374 , n50432 );
and ( n50781 , n50779 , n50780 );
xor ( n50782 , n50779 , n50780 );
xor ( n50783 , n50214 , n50254 );
and ( n50784 , n30379 , n50432 );
and ( n50785 , n50783 , n50784 );
xor ( n50786 , n50783 , n50784 );
xor ( n50787 , n50218 , n50252 );
and ( n50788 , n30384 , n50432 );
and ( n50789 , n50787 , n50788 );
xor ( n50790 , n50787 , n50788 );
xor ( n50791 , n50222 , n50250 );
and ( n50792 , n30389 , n50432 );
and ( n50793 , n50791 , n50792 );
xor ( n50794 , n50791 , n50792 );
xor ( n50795 , n50226 , n50248 );
and ( n50796 , n30394 , n50432 );
and ( n50797 , n50795 , n50796 );
xor ( n50798 , n50795 , n50796 );
xor ( n50799 , n50230 , n50246 );
and ( n50800 , n30399 , n50432 );
and ( n50801 , n50799 , n50800 );
xor ( n50802 , n50799 , n50800 );
xor ( n50803 , n50234 , n50244 );
and ( n50804 , n30404 , n50432 );
and ( n50805 , n50803 , n50804 );
xor ( n50806 , n50803 , n50804 );
xor ( n50807 , n50238 , n50242 );
and ( n50808 , n30409 , n50432 );
and ( n50809 , n50807 , n50808 );
buf ( n50810 , n50809 );
and ( n50811 , n50806 , n50810 );
or ( n50812 , n50805 , n50811 );
and ( n50813 , n50802 , n50812 );
or ( n50814 , n50801 , n50813 );
and ( n50815 , n50798 , n50814 );
or ( n50816 , n50797 , n50815 );
and ( n50817 , n50794 , n50816 );
or ( n50818 , n50793 , n50817 );
and ( n50819 , n50790 , n50818 );
or ( n50820 , n50789 , n50819 );
and ( n50821 , n50786 , n50820 );
or ( n50822 , n50785 , n50821 );
and ( n50823 , n50782 , n50822 );
or ( n50824 , n50781 , n50823 );
and ( n50825 , n50778 , n50824 );
or ( n50826 , n50777 , n50825 );
and ( n50827 , n50774 , n50826 );
or ( n50828 , n50773 , n50827 );
and ( n50829 , n50770 , n50828 );
or ( n50830 , n50769 , n50829 );
and ( n50831 , n50766 , n50830 );
or ( n50832 , n50765 , n50831 );
and ( n50833 , n50762 , n50832 );
or ( n50834 , n50761 , n50833 );
and ( n50835 , n50758 , n50834 );
or ( n50836 , n50757 , n50835 );
and ( n50837 , n50754 , n50836 );
or ( n50838 , n50753 , n50837 );
and ( n50839 , n50750 , n50838 );
or ( n50840 , n50749 , n50839 );
and ( n50841 , n50746 , n50840 );
or ( n50842 , n50745 , n50841 );
and ( n50843 , n50742 , n50842 );
or ( n50844 , n50741 , n50843 );
and ( n50845 , n50738 , n50844 );
or ( n50846 , n50737 , n50845 );
and ( n50847 , n50734 , n50846 );
or ( n50848 , n50733 , n50847 );
and ( n50849 , n50730 , n50848 );
or ( n50850 , n50729 , n50849 );
and ( n50851 , n50726 , n50850 );
or ( n50852 , n50725 , n50851 );
and ( n50853 , n50722 , n50852 );
or ( n50854 , n50721 , n50853 );
and ( n50855 , n50718 , n50854 );
or ( n50856 , n50717 , n50855 );
and ( n50857 , n50714 , n50856 );
or ( n50858 , n50713 , n50857 );
and ( n50859 , n50710 , n50858 );
or ( n50860 , n50709 , n50859 );
and ( n50861 , n50706 , n50860 );
or ( n50862 , n50705 , n50861 );
and ( n50863 , n50702 , n50862 );
or ( n50864 , n50701 , n50863 );
and ( n50865 , n50698 , n50864 );
or ( n50866 , n50697 , n50865 );
and ( n50867 , n50694 , n50866 );
or ( n50868 , n50693 , n50867 );
and ( n50869 , n50690 , n50868 );
or ( n50870 , n50689 , n50869 );
and ( n50871 , n50686 , n50870 );
or ( n50872 , n50685 , n50871 );
and ( n50873 , n50682 , n50872 );
or ( n50874 , n50681 , n50873 );
and ( n50875 , n50678 , n50874 );
or ( n50876 , n50677 , n50875 );
and ( n50877 , n50674 , n50876 );
or ( n50878 , n50673 , n50877 );
and ( n50879 , n50670 , n50878 );
or ( n50880 , n50669 , n50879 );
and ( n50881 , n50666 , n50880 );
or ( n50882 , n50665 , n50881 );
and ( n50883 , n50662 , n50882 );
or ( n50884 , n50661 , n50883 );
and ( n50885 , n50658 , n50884 );
or ( n50886 , n50657 , n50885 );
and ( n50887 , n50654 , n50886 );
or ( n50888 , n50653 , n50887 );
and ( n50889 , n50650 , n50888 );
or ( n50890 , n50649 , n50889 );
and ( n50891 , n50646 , n50890 );
or ( n50892 , n50645 , n50891 );
and ( n50893 , n50642 , n50892 );
or ( n50894 , n50641 , n50893 );
and ( n50895 , n50638 , n50894 );
or ( n50896 , n50637 , n50895 );
and ( n50897 , n50634 , n50896 );
or ( n50898 , n50633 , n50897 );
and ( n50899 , n50630 , n50898 );
or ( n50900 , n50629 , n50899 );
and ( n50901 , n50626 , n50900 );
or ( n50902 , n50625 , n50901 );
and ( n50903 , n50622 , n50902 );
or ( n50904 , n50621 , n50903 );
and ( n50905 , n50618 , n50904 );
or ( n50906 , n50617 , n50905 );
and ( n50907 , n50614 , n50906 );
or ( n50908 , n50613 , n50907 );
and ( n50909 , n50610 , n50908 );
or ( n50910 , n50609 , n50909 );
and ( n50911 , n50606 , n50910 );
or ( n50912 , n50605 , n50911 );
and ( n50913 , n50602 , n50912 );
or ( n50914 , n50601 , n50913 );
and ( n50915 , n50598 , n50914 );
or ( n50916 , n50597 , n50915 );
and ( n50917 , n50594 , n50916 );
or ( n50918 , n50593 , n50917 );
and ( n50919 , n50590 , n50918 );
or ( n50920 , n50589 , n50919 );
and ( n50921 , n50586 , n50920 );
or ( n50922 , n50585 , n50921 );
and ( n50923 , n50582 , n50922 );
or ( n50924 , n50581 , n50923 );
and ( n50925 , n50578 , n50924 );
or ( n50926 , n50577 , n50925 );
and ( n50927 , n50574 , n50926 );
or ( n50928 , n50573 , n50927 );
and ( n50929 , n50570 , n50928 );
or ( n50930 , n50569 , n50929 );
and ( n50931 , n50566 , n50930 );
or ( n50932 , n50565 , n50931 );
and ( n50933 , n50562 , n50932 );
or ( n50934 , n50561 , n50933 );
and ( n50935 , n50558 , n50934 );
or ( n50936 , n50557 , n50935 );
and ( n50937 , n50554 , n50936 );
or ( n50938 , n50553 , n50937 );
and ( n50939 , n50550 , n50938 );
or ( n50940 , n50549 , n50939 );
and ( n50941 , n50546 , n50940 );
or ( n50942 , n50545 , n50941 );
and ( n50943 , n50542 , n50942 );
or ( n50944 , n50541 , n50943 );
and ( n50945 , n50538 , n50944 );
or ( n50946 , n50537 , n50945 );
and ( n50947 , n50534 , n50946 );
or ( n50948 , n50533 , n50947 );
and ( n50949 , n50530 , n50948 );
or ( n50950 , n50529 , n50949 );
and ( n50951 , n50526 , n50950 );
or ( n50952 , n50525 , n50951 );
and ( n50953 , n50522 , n50952 );
or ( n50954 , n50521 , n50953 );
and ( n50955 , n50518 , n50954 );
or ( n50956 , n50517 , n50955 );
and ( n50957 , n50514 , n50956 );
or ( n50958 , n50513 , n50957 );
and ( n50959 , n50510 , n50958 );
or ( n50960 , n50509 , n50959 );
and ( n50961 , n50506 , n50960 );
or ( n50962 , n50505 , n50961 );
and ( n50963 , n50502 , n50962 );
or ( n50964 , n50501 , n50963 );
and ( n50965 , n50498 , n50964 );
or ( n50966 , n50497 , n50965 );
and ( n50967 , n50494 , n50966 );
or ( n50968 , n50493 , n50967 );
and ( n50969 , n50490 , n50968 );
or ( n50970 , n50489 , n50969 );
and ( n50971 , n50486 , n50970 );
or ( n50972 , n50485 , n50971 );
and ( n50973 , n50482 , n50972 );
or ( n50974 , n50481 , n50973 );
and ( n50975 , n50478 , n50974 );
or ( n50976 , n50477 , n50975 );
and ( n50977 , n50474 , n50976 );
or ( n50978 , n50473 , n50977 );
and ( n50979 , n50470 , n50978 );
or ( n50980 , n50469 , n50979 );
and ( n50981 , n50466 , n50980 );
or ( n50982 , n50465 , n50981 );
and ( n50983 , n50462 , n50982 );
or ( n50984 , n50461 , n50983 );
and ( n50985 , n50458 , n50984 );
or ( n50986 , n50457 , n50985 );
and ( n50987 , n50454 , n50986 );
or ( n50988 , n50453 , n50987 );
and ( n50989 , n50450 , n50988 );
or ( n50990 , n50449 , n50989 );
and ( n50991 , n50446 , n50990 );
or ( n50992 , n50445 , n50991 );
and ( n50993 , n50442 , n50992 );
or ( n50994 , n50441 , n50993 );
and ( n50995 , n50438 , n50994 );
or ( n50996 , n50437 , n50995 );
xor ( n50997 , n50434 , n50996 );
buf ( n50998 , n18040 );
and ( n50999 , n29944 , n50998 );
xor ( n51000 , n50997 , n50999 );
xor ( n51001 , n50438 , n50994 );
and ( n51002 , n29949 , n50998 );
and ( n51003 , n51001 , n51002 );
xor ( n51004 , n51001 , n51002 );
xor ( n51005 , n50442 , n50992 );
and ( n51006 , n29954 , n50998 );
and ( n51007 , n51005 , n51006 );
xor ( n51008 , n51005 , n51006 );
xor ( n51009 , n50446 , n50990 );
and ( n51010 , n29959 , n50998 );
and ( n51011 , n51009 , n51010 );
xor ( n51012 , n51009 , n51010 );
xor ( n51013 , n50450 , n50988 );
and ( n51014 , n29964 , n50998 );
and ( n51015 , n51013 , n51014 );
xor ( n51016 , n51013 , n51014 );
xor ( n51017 , n50454 , n50986 );
and ( n51018 , n29969 , n50998 );
and ( n51019 , n51017 , n51018 );
xor ( n51020 , n51017 , n51018 );
xor ( n51021 , n50458 , n50984 );
and ( n51022 , n29974 , n50998 );
and ( n51023 , n51021 , n51022 );
xor ( n51024 , n51021 , n51022 );
xor ( n51025 , n50462 , n50982 );
and ( n51026 , n29979 , n50998 );
and ( n51027 , n51025 , n51026 );
xor ( n51028 , n51025 , n51026 );
xor ( n51029 , n50466 , n50980 );
and ( n51030 , n29984 , n50998 );
and ( n51031 , n51029 , n51030 );
xor ( n51032 , n51029 , n51030 );
xor ( n51033 , n50470 , n50978 );
and ( n51034 , n29989 , n50998 );
and ( n51035 , n51033 , n51034 );
xor ( n51036 , n51033 , n51034 );
xor ( n51037 , n50474 , n50976 );
and ( n51038 , n29994 , n50998 );
and ( n51039 , n51037 , n51038 );
xor ( n51040 , n51037 , n51038 );
xor ( n51041 , n50478 , n50974 );
and ( n51042 , n29999 , n50998 );
and ( n51043 , n51041 , n51042 );
xor ( n51044 , n51041 , n51042 );
xor ( n51045 , n50482 , n50972 );
and ( n51046 , n30004 , n50998 );
and ( n51047 , n51045 , n51046 );
xor ( n51048 , n51045 , n51046 );
xor ( n51049 , n50486 , n50970 );
and ( n51050 , n30009 , n50998 );
and ( n51051 , n51049 , n51050 );
xor ( n51052 , n51049 , n51050 );
xor ( n51053 , n50490 , n50968 );
and ( n51054 , n30014 , n50998 );
and ( n51055 , n51053 , n51054 );
xor ( n51056 , n51053 , n51054 );
xor ( n51057 , n50494 , n50966 );
and ( n51058 , n30019 , n50998 );
and ( n51059 , n51057 , n51058 );
xor ( n51060 , n51057 , n51058 );
xor ( n51061 , n50498 , n50964 );
and ( n51062 , n30024 , n50998 );
and ( n51063 , n51061 , n51062 );
xor ( n51064 , n51061 , n51062 );
xor ( n51065 , n50502 , n50962 );
and ( n51066 , n30029 , n50998 );
and ( n51067 , n51065 , n51066 );
xor ( n51068 , n51065 , n51066 );
xor ( n51069 , n50506 , n50960 );
and ( n51070 , n30034 , n50998 );
and ( n51071 , n51069 , n51070 );
xor ( n51072 , n51069 , n51070 );
xor ( n51073 , n50510 , n50958 );
and ( n51074 , n30039 , n50998 );
and ( n51075 , n51073 , n51074 );
xor ( n51076 , n51073 , n51074 );
xor ( n51077 , n50514 , n50956 );
and ( n51078 , n30044 , n50998 );
and ( n51079 , n51077 , n51078 );
xor ( n51080 , n51077 , n51078 );
xor ( n51081 , n50518 , n50954 );
and ( n51082 , n30049 , n50998 );
and ( n51083 , n51081 , n51082 );
xor ( n51084 , n51081 , n51082 );
xor ( n51085 , n50522 , n50952 );
and ( n51086 , n30054 , n50998 );
and ( n51087 , n51085 , n51086 );
xor ( n51088 , n51085 , n51086 );
xor ( n51089 , n50526 , n50950 );
and ( n51090 , n30059 , n50998 );
and ( n51091 , n51089 , n51090 );
xor ( n51092 , n51089 , n51090 );
xor ( n51093 , n50530 , n50948 );
and ( n51094 , n30064 , n50998 );
and ( n51095 , n51093 , n51094 );
xor ( n51096 , n51093 , n51094 );
xor ( n51097 , n50534 , n50946 );
and ( n51098 , n30069 , n50998 );
and ( n51099 , n51097 , n51098 );
xor ( n51100 , n51097 , n51098 );
xor ( n51101 , n50538 , n50944 );
and ( n51102 , n30074 , n50998 );
and ( n51103 , n51101 , n51102 );
xor ( n51104 , n51101 , n51102 );
xor ( n51105 , n50542 , n50942 );
and ( n51106 , n30079 , n50998 );
and ( n51107 , n51105 , n51106 );
xor ( n51108 , n51105 , n51106 );
xor ( n51109 , n50546 , n50940 );
and ( n51110 , n30084 , n50998 );
and ( n51111 , n51109 , n51110 );
xor ( n51112 , n51109 , n51110 );
xor ( n51113 , n50550 , n50938 );
and ( n51114 , n30089 , n50998 );
and ( n51115 , n51113 , n51114 );
xor ( n51116 , n51113 , n51114 );
xor ( n51117 , n50554 , n50936 );
and ( n51118 , n30094 , n50998 );
and ( n51119 , n51117 , n51118 );
xor ( n51120 , n51117 , n51118 );
xor ( n51121 , n50558 , n50934 );
and ( n51122 , n30099 , n50998 );
and ( n51123 , n51121 , n51122 );
xor ( n51124 , n51121 , n51122 );
xor ( n51125 , n50562 , n50932 );
and ( n51126 , n30104 , n50998 );
and ( n51127 , n51125 , n51126 );
xor ( n51128 , n51125 , n51126 );
xor ( n51129 , n50566 , n50930 );
and ( n51130 , n30109 , n50998 );
and ( n51131 , n51129 , n51130 );
xor ( n51132 , n51129 , n51130 );
xor ( n51133 , n50570 , n50928 );
and ( n51134 , n30114 , n50998 );
and ( n51135 , n51133 , n51134 );
xor ( n51136 , n51133 , n51134 );
xor ( n51137 , n50574 , n50926 );
and ( n51138 , n30119 , n50998 );
and ( n51139 , n51137 , n51138 );
xor ( n51140 , n51137 , n51138 );
xor ( n51141 , n50578 , n50924 );
and ( n51142 , n30124 , n50998 );
and ( n51143 , n51141 , n51142 );
xor ( n51144 , n51141 , n51142 );
xor ( n51145 , n50582 , n50922 );
and ( n51146 , n30129 , n50998 );
and ( n51147 , n51145 , n51146 );
xor ( n51148 , n51145 , n51146 );
xor ( n51149 , n50586 , n50920 );
and ( n51150 , n30134 , n50998 );
and ( n51151 , n51149 , n51150 );
xor ( n51152 , n51149 , n51150 );
xor ( n51153 , n50590 , n50918 );
and ( n51154 , n30139 , n50998 );
and ( n51155 , n51153 , n51154 );
xor ( n51156 , n51153 , n51154 );
xor ( n51157 , n50594 , n50916 );
and ( n51158 , n30144 , n50998 );
and ( n51159 , n51157 , n51158 );
xor ( n51160 , n51157 , n51158 );
xor ( n51161 , n50598 , n50914 );
and ( n51162 , n30149 , n50998 );
and ( n51163 , n51161 , n51162 );
xor ( n51164 , n51161 , n51162 );
xor ( n51165 , n50602 , n50912 );
and ( n51166 , n30154 , n50998 );
and ( n51167 , n51165 , n51166 );
xor ( n51168 , n51165 , n51166 );
xor ( n51169 , n50606 , n50910 );
and ( n51170 , n30159 , n50998 );
and ( n51171 , n51169 , n51170 );
xor ( n51172 , n51169 , n51170 );
xor ( n51173 , n50610 , n50908 );
and ( n51174 , n30164 , n50998 );
and ( n51175 , n51173 , n51174 );
xor ( n51176 , n51173 , n51174 );
xor ( n51177 , n50614 , n50906 );
and ( n51178 , n30169 , n50998 );
and ( n51179 , n51177 , n51178 );
xor ( n51180 , n51177 , n51178 );
xor ( n51181 , n50618 , n50904 );
and ( n51182 , n30174 , n50998 );
and ( n51183 , n51181 , n51182 );
xor ( n51184 , n51181 , n51182 );
xor ( n51185 , n50622 , n50902 );
and ( n51186 , n30179 , n50998 );
and ( n51187 , n51185 , n51186 );
xor ( n51188 , n51185 , n51186 );
xor ( n51189 , n50626 , n50900 );
and ( n51190 , n30184 , n50998 );
and ( n51191 , n51189 , n51190 );
xor ( n51192 , n51189 , n51190 );
xor ( n51193 , n50630 , n50898 );
and ( n51194 , n30189 , n50998 );
and ( n51195 , n51193 , n51194 );
xor ( n51196 , n51193 , n51194 );
xor ( n51197 , n50634 , n50896 );
and ( n51198 , n30194 , n50998 );
and ( n51199 , n51197 , n51198 );
xor ( n51200 , n51197 , n51198 );
xor ( n51201 , n50638 , n50894 );
and ( n51202 , n30199 , n50998 );
and ( n51203 , n51201 , n51202 );
xor ( n51204 , n51201 , n51202 );
xor ( n51205 , n50642 , n50892 );
and ( n51206 , n30204 , n50998 );
and ( n51207 , n51205 , n51206 );
xor ( n51208 , n51205 , n51206 );
xor ( n51209 , n50646 , n50890 );
and ( n51210 , n30209 , n50998 );
and ( n51211 , n51209 , n51210 );
xor ( n51212 , n51209 , n51210 );
xor ( n51213 , n50650 , n50888 );
and ( n51214 , n30214 , n50998 );
and ( n51215 , n51213 , n51214 );
xor ( n51216 , n51213 , n51214 );
xor ( n51217 , n50654 , n50886 );
and ( n51218 , n30219 , n50998 );
and ( n51219 , n51217 , n51218 );
xor ( n51220 , n51217 , n51218 );
xor ( n51221 , n50658 , n50884 );
and ( n51222 , n30224 , n50998 );
and ( n51223 , n51221 , n51222 );
xor ( n51224 , n51221 , n51222 );
xor ( n51225 , n50662 , n50882 );
and ( n51226 , n30229 , n50998 );
and ( n51227 , n51225 , n51226 );
xor ( n51228 , n51225 , n51226 );
xor ( n51229 , n50666 , n50880 );
and ( n51230 , n30234 , n50998 );
and ( n51231 , n51229 , n51230 );
xor ( n51232 , n51229 , n51230 );
xor ( n51233 , n50670 , n50878 );
and ( n51234 , n30239 , n50998 );
and ( n51235 , n51233 , n51234 );
xor ( n51236 , n51233 , n51234 );
xor ( n51237 , n50674 , n50876 );
and ( n51238 , n30244 , n50998 );
and ( n51239 , n51237 , n51238 );
xor ( n51240 , n51237 , n51238 );
xor ( n51241 , n50678 , n50874 );
and ( n51242 , n30249 , n50998 );
and ( n51243 , n51241 , n51242 );
xor ( n51244 , n51241 , n51242 );
xor ( n51245 , n50682 , n50872 );
and ( n51246 , n30254 , n50998 );
and ( n51247 , n51245 , n51246 );
xor ( n51248 , n51245 , n51246 );
xor ( n51249 , n50686 , n50870 );
and ( n51250 , n30259 , n50998 );
and ( n51251 , n51249 , n51250 );
xor ( n51252 , n51249 , n51250 );
xor ( n51253 , n50690 , n50868 );
and ( n51254 , n30264 , n50998 );
and ( n51255 , n51253 , n51254 );
xor ( n51256 , n51253 , n51254 );
xor ( n51257 , n50694 , n50866 );
and ( n51258 , n30269 , n50998 );
and ( n51259 , n51257 , n51258 );
xor ( n51260 , n51257 , n51258 );
xor ( n51261 , n50698 , n50864 );
and ( n51262 , n30274 , n50998 );
and ( n51263 , n51261 , n51262 );
xor ( n51264 , n51261 , n51262 );
xor ( n51265 , n50702 , n50862 );
and ( n51266 , n30279 , n50998 );
and ( n51267 , n51265 , n51266 );
xor ( n51268 , n51265 , n51266 );
xor ( n51269 , n50706 , n50860 );
and ( n51270 , n30284 , n50998 );
and ( n51271 , n51269 , n51270 );
xor ( n51272 , n51269 , n51270 );
xor ( n51273 , n50710 , n50858 );
and ( n51274 , n30289 , n50998 );
and ( n51275 , n51273 , n51274 );
xor ( n51276 , n51273 , n51274 );
xor ( n51277 , n50714 , n50856 );
and ( n51278 , n30294 , n50998 );
and ( n51279 , n51277 , n51278 );
xor ( n51280 , n51277 , n51278 );
xor ( n51281 , n50718 , n50854 );
and ( n51282 , n30299 , n50998 );
and ( n51283 , n51281 , n51282 );
xor ( n51284 , n51281 , n51282 );
xor ( n51285 , n50722 , n50852 );
and ( n51286 , n30304 , n50998 );
and ( n51287 , n51285 , n51286 );
xor ( n51288 , n51285 , n51286 );
xor ( n51289 , n50726 , n50850 );
and ( n51290 , n30309 , n50998 );
and ( n51291 , n51289 , n51290 );
xor ( n51292 , n51289 , n51290 );
xor ( n51293 , n50730 , n50848 );
and ( n51294 , n30314 , n50998 );
and ( n51295 , n51293 , n51294 );
xor ( n51296 , n51293 , n51294 );
xor ( n51297 , n50734 , n50846 );
and ( n51298 , n30319 , n50998 );
and ( n51299 , n51297 , n51298 );
xor ( n51300 , n51297 , n51298 );
xor ( n51301 , n50738 , n50844 );
and ( n51302 , n30324 , n50998 );
and ( n51303 , n51301 , n51302 );
xor ( n51304 , n51301 , n51302 );
xor ( n51305 , n50742 , n50842 );
and ( n51306 , n30329 , n50998 );
and ( n51307 , n51305 , n51306 );
xor ( n51308 , n51305 , n51306 );
xor ( n51309 , n50746 , n50840 );
and ( n51310 , n30334 , n50998 );
and ( n51311 , n51309 , n51310 );
xor ( n51312 , n51309 , n51310 );
xor ( n51313 , n50750 , n50838 );
and ( n51314 , n30339 , n50998 );
and ( n51315 , n51313 , n51314 );
xor ( n51316 , n51313 , n51314 );
xor ( n51317 , n50754 , n50836 );
and ( n51318 , n30344 , n50998 );
and ( n51319 , n51317 , n51318 );
xor ( n51320 , n51317 , n51318 );
xor ( n51321 , n50758 , n50834 );
and ( n51322 , n30349 , n50998 );
and ( n51323 , n51321 , n51322 );
xor ( n51324 , n51321 , n51322 );
xor ( n51325 , n50762 , n50832 );
and ( n51326 , n30354 , n50998 );
and ( n51327 , n51325 , n51326 );
xor ( n51328 , n51325 , n51326 );
xor ( n51329 , n50766 , n50830 );
and ( n51330 , n30359 , n50998 );
and ( n51331 , n51329 , n51330 );
xor ( n51332 , n51329 , n51330 );
xor ( n51333 , n50770 , n50828 );
and ( n51334 , n30364 , n50998 );
and ( n51335 , n51333 , n51334 );
xor ( n51336 , n51333 , n51334 );
xor ( n51337 , n50774 , n50826 );
and ( n51338 , n30369 , n50998 );
and ( n51339 , n51337 , n51338 );
xor ( n51340 , n51337 , n51338 );
xor ( n51341 , n50778 , n50824 );
and ( n51342 , n30374 , n50998 );
and ( n51343 , n51341 , n51342 );
xor ( n51344 , n51341 , n51342 );
xor ( n51345 , n50782 , n50822 );
and ( n51346 , n30379 , n50998 );
and ( n51347 , n51345 , n51346 );
xor ( n51348 , n51345 , n51346 );
xor ( n51349 , n50786 , n50820 );
and ( n51350 , n30384 , n50998 );
and ( n51351 , n51349 , n51350 );
xor ( n51352 , n51349 , n51350 );
xor ( n51353 , n50790 , n50818 );
and ( n51354 , n30389 , n50998 );
and ( n51355 , n51353 , n51354 );
xor ( n51356 , n51353 , n51354 );
xor ( n51357 , n50794 , n50816 );
and ( n51358 , n30394 , n50998 );
and ( n51359 , n51357 , n51358 );
xor ( n51360 , n51357 , n51358 );
xor ( n51361 , n50798 , n50814 );
and ( n51362 , n30399 , n50998 );
and ( n51363 , n51361 , n51362 );
xor ( n51364 , n51361 , n51362 );
xor ( n51365 , n50802 , n50812 );
and ( n51366 , n30404 , n50998 );
and ( n51367 , n51365 , n51366 );
xor ( n51368 , n51365 , n51366 );
xor ( n51369 , n50806 , n50810 );
and ( n51370 , n30409 , n50998 );
and ( n51371 , n51369 , n51370 );
buf ( n51372 , n51371 );
and ( n51373 , n51368 , n51372 );
or ( n51374 , n51367 , n51373 );
and ( n51375 , n51364 , n51374 );
or ( n51376 , n51363 , n51375 );
and ( n51377 , n51360 , n51376 );
or ( n51378 , n51359 , n51377 );
and ( n51379 , n51356 , n51378 );
or ( n51380 , n51355 , n51379 );
and ( n51381 , n51352 , n51380 );
or ( n51382 , n51351 , n51381 );
and ( n51383 , n51348 , n51382 );
or ( n51384 , n51347 , n51383 );
and ( n51385 , n51344 , n51384 );
or ( n51386 , n51343 , n51385 );
and ( n51387 , n51340 , n51386 );
or ( n51388 , n51339 , n51387 );
and ( n51389 , n51336 , n51388 );
or ( n51390 , n51335 , n51389 );
and ( n51391 , n51332 , n51390 );
or ( n51392 , n51331 , n51391 );
and ( n51393 , n51328 , n51392 );
or ( n51394 , n51327 , n51393 );
and ( n51395 , n51324 , n51394 );
or ( n51396 , n51323 , n51395 );
and ( n51397 , n51320 , n51396 );
or ( n51398 , n51319 , n51397 );
and ( n51399 , n51316 , n51398 );
or ( n51400 , n51315 , n51399 );
and ( n51401 , n51312 , n51400 );
or ( n51402 , n51311 , n51401 );
and ( n51403 , n51308 , n51402 );
or ( n51404 , n51307 , n51403 );
and ( n51405 , n51304 , n51404 );
or ( n51406 , n51303 , n51405 );
and ( n51407 , n51300 , n51406 );
or ( n51408 , n51299 , n51407 );
and ( n51409 , n51296 , n51408 );
or ( n51410 , n51295 , n51409 );
and ( n51411 , n51292 , n51410 );
or ( n51412 , n51291 , n51411 );
and ( n51413 , n51288 , n51412 );
or ( n51414 , n51287 , n51413 );
and ( n51415 , n51284 , n51414 );
or ( n51416 , n51283 , n51415 );
and ( n51417 , n51280 , n51416 );
or ( n51418 , n51279 , n51417 );
and ( n51419 , n51276 , n51418 );
or ( n51420 , n51275 , n51419 );
and ( n51421 , n51272 , n51420 );
or ( n51422 , n51271 , n51421 );
and ( n51423 , n51268 , n51422 );
or ( n51424 , n51267 , n51423 );
and ( n51425 , n51264 , n51424 );
or ( n51426 , n51263 , n51425 );
and ( n51427 , n51260 , n51426 );
or ( n51428 , n51259 , n51427 );
and ( n51429 , n51256 , n51428 );
or ( n51430 , n51255 , n51429 );
and ( n51431 , n51252 , n51430 );
or ( n51432 , n51251 , n51431 );
and ( n51433 , n51248 , n51432 );
or ( n51434 , n51247 , n51433 );
and ( n51435 , n51244 , n51434 );
or ( n51436 , n51243 , n51435 );
and ( n51437 , n51240 , n51436 );
or ( n51438 , n51239 , n51437 );
and ( n51439 , n51236 , n51438 );
or ( n51440 , n51235 , n51439 );
and ( n51441 , n51232 , n51440 );
or ( n51442 , n51231 , n51441 );
and ( n51443 , n51228 , n51442 );
or ( n51444 , n51227 , n51443 );
and ( n51445 , n51224 , n51444 );
or ( n51446 , n51223 , n51445 );
and ( n51447 , n51220 , n51446 );
or ( n51448 , n51219 , n51447 );
and ( n51449 , n51216 , n51448 );
or ( n51450 , n51215 , n51449 );
and ( n51451 , n51212 , n51450 );
or ( n51452 , n51211 , n51451 );
and ( n51453 , n51208 , n51452 );
or ( n51454 , n51207 , n51453 );
and ( n51455 , n51204 , n51454 );
or ( n51456 , n51203 , n51455 );
and ( n51457 , n51200 , n51456 );
or ( n51458 , n51199 , n51457 );
and ( n51459 , n51196 , n51458 );
or ( n51460 , n51195 , n51459 );
and ( n51461 , n51192 , n51460 );
or ( n51462 , n51191 , n51461 );
and ( n51463 , n51188 , n51462 );
or ( n51464 , n51187 , n51463 );
and ( n51465 , n51184 , n51464 );
or ( n51466 , n51183 , n51465 );
and ( n51467 , n51180 , n51466 );
or ( n51468 , n51179 , n51467 );
and ( n51469 , n51176 , n51468 );
or ( n51470 , n51175 , n51469 );
and ( n51471 , n51172 , n51470 );
or ( n51472 , n51171 , n51471 );
and ( n51473 , n51168 , n51472 );
or ( n51474 , n51167 , n51473 );
and ( n51475 , n51164 , n51474 );
or ( n51476 , n51163 , n51475 );
and ( n51477 , n51160 , n51476 );
or ( n51478 , n51159 , n51477 );
and ( n51479 , n51156 , n51478 );
or ( n51480 , n51155 , n51479 );
and ( n51481 , n51152 , n51480 );
or ( n51482 , n51151 , n51481 );
and ( n51483 , n51148 , n51482 );
or ( n51484 , n51147 , n51483 );
and ( n51485 , n51144 , n51484 );
or ( n51486 , n51143 , n51485 );
and ( n51487 , n51140 , n51486 );
or ( n51488 , n51139 , n51487 );
and ( n51489 , n51136 , n51488 );
or ( n51490 , n51135 , n51489 );
and ( n51491 , n51132 , n51490 );
or ( n51492 , n51131 , n51491 );
and ( n51493 , n51128 , n51492 );
or ( n51494 , n51127 , n51493 );
and ( n51495 , n51124 , n51494 );
or ( n51496 , n51123 , n51495 );
and ( n51497 , n51120 , n51496 );
or ( n51498 , n51119 , n51497 );
and ( n51499 , n51116 , n51498 );
or ( n51500 , n51115 , n51499 );
and ( n51501 , n51112 , n51500 );
or ( n51502 , n51111 , n51501 );
and ( n51503 , n51108 , n51502 );
or ( n51504 , n51107 , n51503 );
and ( n51505 , n51104 , n51504 );
or ( n51506 , n51103 , n51505 );
and ( n51507 , n51100 , n51506 );
or ( n51508 , n51099 , n51507 );
and ( n51509 , n51096 , n51508 );
or ( n51510 , n51095 , n51509 );
and ( n51511 , n51092 , n51510 );
or ( n51512 , n51091 , n51511 );
and ( n51513 , n51088 , n51512 );
or ( n51514 , n51087 , n51513 );
and ( n51515 , n51084 , n51514 );
or ( n51516 , n51083 , n51515 );
and ( n51517 , n51080 , n51516 );
or ( n51518 , n51079 , n51517 );
and ( n51519 , n51076 , n51518 );
or ( n51520 , n51075 , n51519 );
and ( n51521 , n51072 , n51520 );
or ( n51522 , n51071 , n51521 );
and ( n51523 , n51068 , n51522 );
or ( n51524 , n51067 , n51523 );
and ( n51525 , n51064 , n51524 );
or ( n51526 , n51063 , n51525 );
and ( n51527 , n51060 , n51526 );
or ( n51528 , n51059 , n51527 );
and ( n51529 , n51056 , n51528 );
or ( n51530 , n51055 , n51529 );
and ( n51531 , n51052 , n51530 );
or ( n51532 , n51051 , n51531 );
and ( n51533 , n51048 , n51532 );
or ( n51534 , n51047 , n51533 );
and ( n51535 , n51044 , n51534 );
or ( n51536 , n51043 , n51535 );
and ( n51537 , n51040 , n51536 );
or ( n51538 , n51039 , n51537 );
and ( n51539 , n51036 , n51538 );
or ( n51540 , n51035 , n51539 );
and ( n51541 , n51032 , n51540 );
or ( n51542 , n51031 , n51541 );
and ( n51543 , n51028 , n51542 );
or ( n51544 , n51027 , n51543 );
and ( n51545 , n51024 , n51544 );
or ( n51546 , n51023 , n51545 );
and ( n51547 , n51020 , n51546 );
or ( n51548 , n51019 , n51547 );
and ( n51549 , n51016 , n51548 );
or ( n51550 , n51015 , n51549 );
and ( n51551 , n51012 , n51550 );
or ( n51552 , n51011 , n51551 );
and ( n51553 , n51008 , n51552 );
or ( n51554 , n51007 , n51553 );
and ( n51555 , n51004 , n51554 );
or ( n51556 , n51003 , n51555 );
xor ( n51557 , n51000 , n51556 );
buf ( n51558 , n18038 );
and ( n51559 , n29949 , n51558 );
xor ( n51560 , n51557 , n51559 );
xor ( n51561 , n51004 , n51554 );
and ( n51562 , n29954 , n51558 );
and ( n51563 , n51561 , n51562 );
xor ( n51564 , n51561 , n51562 );
xor ( n51565 , n51008 , n51552 );
and ( n51566 , n29959 , n51558 );
and ( n51567 , n51565 , n51566 );
xor ( n51568 , n51565 , n51566 );
xor ( n51569 , n51012 , n51550 );
and ( n51570 , n29964 , n51558 );
and ( n51571 , n51569 , n51570 );
xor ( n51572 , n51569 , n51570 );
xor ( n51573 , n51016 , n51548 );
and ( n51574 , n29969 , n51558 );
and ( n51575 , n51573 , n51574 );
xor ( n51576 , n51573 , n51574 );
xor ( n51577 , n51020 , n51546 );
and ( n51578 , n29974 , n51558 );
and ( n51579 , n51577 , n51578 );
xor ( n51580 , n51577 , n51578 );
xor ( n51581 , n51024 , n51544 );
and ( n51582 , n29979 , n51558 );
and ( n51583 , n51581 , n51582 );
xor ( n51584 , n51581 , n51582 );
xor ( n51585 , n51028 , n51542 );
and ( n51586 , n29984 , n51558 );
and ( n51587 , n51585 , n51586 );
xor ( n51588 , n51585 , n51586 );
xor ( n51589 , n51032 , n51540 );
and ( n51590 , n29989 , n51558 );
and ( n51591 , n51589 , n51590 );
xor ( n51592 , n51589 , n51590 );
xor ( n51593 , n51036 , n51538 );
and ( n51594 , n29994 , n51558 );
and ( n51595 , n51593 , n51594 );
xor ( n51596 , n51593 , n51594 );
xor ( n51597 , n51040 , n51536 );
and ( n51598 , n29999 , n51558 );
and ( n51599 , n51597 , n51598 );
xor ( n51600 , n51597 , n51598 );
xor ( n51601 , n51044 , n51534 );
and ( n51602 , n30004 , n51558 );
and ( n51603 , n51601 , n51602 );
xor ( n51604 , n51601 , n51602 );
xor ( n51605 , n51048 , n51532 );
and ( n51606 , n30009 , n51558 );
and ( n51607 , n51605 , n51606 );
xor ( n51608 , n51605 , n51606 );
xor ( n51609 , n51052 , n51530 );
and ( n51610 , n30014 , n51558 );
and ( n51611 , n51609 , n51610 );
xor ( n51612 , n51609 , n51610 );
xor ( n51613 , n51056 , n51528 );
and ( n51614 , n30019 , n51558 );
and ( n51615 , n51613 , n51614 );
xor ( n51616 , n51613 , n51614 );
xor ( n51617 , n51060 , n51526 );
and ( n51618 , n30024 , n51558 );
and ( n51619 , n51617 , n51618 );
xor ( n51620 , n51617 , n51618 );
xor ( n51621 , n51064 , n51524 );
and ( n51622 , n30029 , n51558 );
and ( n51623 , n51621 , n51622 );
xor ( n51624 , n51621 , n51622 );
xor ( n51625 , n51068 , n51522 );
and ( n51626 , n30034 , n51558 );
and ( n51627 , n51625 , n51626 );
xor ( n51628 , n51625 , n51626 );
xor ( n51629 , n51072 , n51520 );
and ( n51630 , n30039 , n51558 );
and ( n51631 , n51629 , n51630 );
xor ( n51632 , n51629 , n51630 );
xor ( n51633 , n51076 , n51518 );
and ( n51634 , n30044 , n51558 );
and ( n51635 , n51633 , n51634 );
xor ( n51636 , n51633 , n51634 );
xor ( n51637 , n51080 , n51516 );
and ( n51638 , n30049 , n51558 );
and ( n51639 , n51637 , n51638 );
xor ( n51640 , n51637 , n51638 );
xor ( n51641 , n51084 , n51514 );
and ( n51642 , n30054 , n51558 );
and ( n51643 , n51641 , n51642 );
xor ( n51644 , n51641 , n51642 );
xor ( n51645 , n51088 , n51512 );
and ( n51646 , n30059 , n51558 );
and ( n51647 , n51645 , n51646 );
xor ( n51648 , n51645 , n51646 );
xor ( n51649 , n51092 , n51510 );
and ( n51650 , n30064 , n51558 );
and ( n51651 , n51649 , n51650 );
xor ( n51652 , n51649 , n51650 );
xor ( n51653 , n51096 , n51508 );
and ( n51654 , n30069 , n51558 );
and ( n51655 , n51653 , n51654 );
xor ( n51656 , n51653 , n51654 );
xor ( n51657 , n51100 , n51506 );
and ( n51658 , n30074 , n51558 );
and ( n51659 , n51657 , n51658 );
xor ( n51660 , n51657 , n51658 );
xor ( n51661 , n51104 , n51504 );
and ( n51662 , n30079 , n51558 );
and ( n51663 , n51661 , n51662 );
xor ( n51664 , n51661 , n51662 );
xor ( n51665 , n51108 , n51502 );
and ( n51666 , n30084 , n51558 );
and ( n51667 , n51665 , n51666 );
xor ( n51668 , n51665 , n51666 );
xor ( n51669 , n51112 , n51500 );
and ( n51670 , n30089 , n51558 );
and ( n51671 , n51669 , n51670 );
xor ( n51672 , n51669 , n51670 );
xor ( n51673 , n51116 , n51498 );
and ( n51674 , n30094 , n51558 );
and ( n51675 , n51673 , n51674 );
xor ( n51676 , n51673 , n51674 );
xor ( n51677 , n51120 , n51496 );
and ( n51678 , n30099 , n51558 );
and ( n51679 , n51677 , n51678 );
xor ( n51680 , n51677 , n51678 );
xor ( n51681 , n51124 , n51494 );
and ( n51682 , n30104 , n51558 );
and ( n51683 , n51681 , n51682 );
xor ( n51684 , n51681 , n51682 );
xor ( n51685 , n51128 , n51492 );
and ( n51686 , n30109 , n51558 );
and ( n51687 , n51685 , n51686 );
xor ( n51688 , n51685 , n51686 );
xor ( n51689 , n51132 , n51490 );
and ( n51690 , n30114 , n51558 );
and ( n51691 , n51689 , n51690 );
xor ( n51692 , n51689 , n51690 );
xor ( n51693 , n51136 , n51488 );
and ( n51694 , n30119 , n51558 );
and ( n51695 , n51693 , n51694 );
xor ( n51696 , n51693 , n51694 );
xor ( n51697 , n51140 , n51486 );
and ( n51698 , n30124 , n51558 );
and ( n51699 , n51697 , n51698 );
xor ( n51700 , n51697 , n51698 );
xor ( n51701 , n51144 , n51484 );
and ( n51702 , n30129 , n51558 );
and ( n51703 , n51701 , n51702 );
xor ( n51704 , n51701 , n51702 );
xor ( n51705 , n51148 , n51482 );
and ( n51706 , n30134 , n51558 );
and ( n51707 , n51705 , n51706 );
xor ( n51708 , n51705 , n51706 );
xor ( n51709 , n51152 , n51480 );
and ( n51710 , n30139 , n51558 );
and ( n51711 , n51709 , n51710 );
xor ( n51712 , n51709 , n51710 );
xor ( n51713 , n51156 , n51478 );
and ( n51714 , n30144 , n51558 );
and ( n51715 , n51713 , n51714 );
xor ( n51716 , n51713 , n51714 );
xor ( n51717 , n51160 , n51476 );
and ( n51718 , n30149 , n51558 );
and ( n51719 , n51717 , n51718 );
xor ( n51720 , n51717 , n51718 );
xor ( n51721 , n51164 , n51474 );
and ( n51722 , n30154 , n51558 );
and ( n51723 , n51721 , n51722 );
xor ( n51724 , n51721 , n51722 );
xor ( n51725 , n51168 , n51472 );
and ( n51726 , n30159 , n51558 );
and ( n51727 , n51725 , n51726 );
xor ( n51728 , n51725 , n51726 );
xor ( n51729 , n51172 , n51470 );
and ( n51730 , n30164 , n51558 );
and ( n51731 , n51729 , n51730 );
xor ( n51732 , n51729 , n51730 );
xor ( n51733 , n51176 , n51468 );
and ( n51734 , n30169 , n51558 );
and ( n51735 , n51733 , n51734 );
xor ( n51736 , n51733 , n51734 );
xor ( n51737 , n51180 , n51466 );
and ( n51738 , n30174 , n51558 );
and ( n51739 , n51737 , n51738 );
xor ( n51740 , n51737 , n51738 );
xor ( n51741 , n51184 , n51464 );
and ( n51742 , n30179 , n51558 );
and ( n51743 , n51741 , n51742 );
xor ( n51744 , n51741 , n51742 );
xor ( n51745 , n51188 , n51462 );
and ( n51746 , n30184 , n51558 );
and ( n51747 , n51745 , n51746 );
xor ( n51748 , n51745 , n51746 );
xor ( n51749 , n51192 , n51460 );
and ( n51750 , n30189 , n51558 );
and ( n51751 , n51749 , n51750 );
xor ( n51752 , n51749 , n51750 );
xor ( n51753 , n51196 , n51458 );
and ( n51754 , n30194 , n51558 );
and ( n51755 , n51753 , n51754 );
xor ( n51756 , n51753 , n51754 );
xor ( n51757 , n51200 , n51456 );
and ( n51758 , n30199 , n51558 );
and ( n51759 , n51757 , n51758 );
xor ( n51760 , n51757 , n51758 );
xor ( n51761 , n51204 , n51454 );
and ( n51762 , n30204 , n51558 );
and ( n51763 , n51761 , n51762 );
xor ( n51764 , n51761 , n51762 );
xor ( n51765 , n51208 , n51452 );
and ( n51766 , n30209 , n51558 );
and ( n51767 , n51765 , n51766 );
xor ( n51768 , n51765 , n51766 );
xor ( n51769 , n51212 , n51450 );
and ( n51770 , n30214 , n51558 );
and ( n51771 , n51769 , n51770 );
xor ( n51772 , n51769 , n51770 );
xor ( n51773 , n51216 , n51448 );
and ( n51774 , n30219 , n51558 );
and ( n51775 , n51773 , n51774 );
xor ( n51776 , n51773 , n51774 );
xor ( n51777 , n51220 , n51446 );
and ( n51778 , n30224 , n51558 );
and ( n51779 , n51777 , n51778 );
xor ( n51780 , n51777 , n51778 );
xor ( n51781 , n51224 , n51444 );
and ( n51782 , n30229 , n51558 );
and ( n51783 , n51781 , n51782 );
xor ( n51784 , n51781 , n51782 );
xor ( n51785 , n51228 , n51442 );
and ( n51786 , n30234 , n51558 );
and ( n51787 , n51785 , n51786 );
xor ( n51788 , n51785 , n51786 );
xor ( n51789 , n51232 , n51440 );
and ( n51790 , n30239 , n51558 );
and ( n51791 , n51789 , n51790 );
xor ( n51792 , n51789 , n51790 );
xor ( n51793 , n51236 , n51438 );
and ( n51794 , n30244 , n51558 );
and ( n51795 , n51793 , n51794 );
xor ( n51796 , n51793 , n51794 );
xor ( n51797 , n51240 , n51436 );
and ( n51798 , n30249 , n51558 );
and ( n51799 , n51797 , n51798 );
xor ( n51800 , n51797 , n51798 );
xor ( n51801 , n51244 , n51434 );
and ( n51802 , n30254 , n51558 );
and ( n51803 , n51801 , n51802 );
xor ( n51804 , n51801 , n51802 );
xor ( n51805 , n51248 , n51432 );
and ( n51806 , n30259 , n51558 );
and ( n51807 , n51805 , n51806 );
xor ( n51808 , n51805 , n51806 );
xor ( n51809 , n51252 , n51430 );
and ( n51810 , n30264 , n51558 );
and ( n51811 , n51809 , n51810 );
xor ( n51812 , n51809 , n51810 );
xor ( n51813 , n51256 , n51428 );
and ( n51814 , n30269 , n51558 );
and ( n51815 , n51813 , n51814 );
xor ( n51816 , n51813 , n51814 );
xor ( n51817 , n51260 , n51426 );
and ( n51818 , n30274 , n51558 );
and ( n51819 , n51817 , n51818 );
xor ( n51820 , n51817 , n51818 );
xor ( n51821 , n51264 , n51424 );
and ( n51822 , n30279 , n51558 );
and ( n51823 , n51821 , n51822 );
xor ( n51824 , n51821 , n51822 );
xor ( n51825 , n51268 , n51422 );
and ( n51826 , n30284 , n51558 );
and ( n51827 , n51825 , n51826 );
xor ( n51828 , n51825 , n51826 );
xor ( n51829 , n51272 , n51420 );
and ( n51830 , n30289 , n51558 );
and ( n51831 , n51829 , n51830 );
xor ( n51832 , n51829 , n51830 );
xor ( n51833 , n51276 , n51418 );
and ( n51834 , n30294 , n51558 );
and ( n51835 , n51833 , n51834 );
xor ( n51836 , n51833 , n51834 );
xor ( n51837 , n51280 , n51416 );
and ( n51838 , n30299 , n51558 );
and ( n51839 , n51837 , n51838 );
xor ( n51840 , n51837 , n51838 );
xor ( n51841 , n51284 , n51414 );
and ( n51842 , n30304 , n51558 );
and ( n51843 , n51841 , n51842 );
xor ( n51844 , n51841 , n51842 );
xor ( n51845 , n51288 , n51412 );
and ( n51846 , n30309 , n51558 );
and ( n51847 , n51845 , n51846 );
xor ( n51848 , n51845 , n51846 );
xor ( n51849 , n51292 , n51410 );
and ( n51850 , n30314 , n51558 );
and ( n51851 , n51849 , n51850 );
xor ( n51852 , n51849 , n51850 );
xor ( n51853 , n51296 , n51408 );
and ( n51854 , n30319 , n51558 );
and ( n51855 , n51853 , n51854 );
xor ( n51856 , n51853 , n51854 );
xor ( n51857 , n51300 , n51406 );
and ( n51858 , n30324 , n51558 );
and ( n51859 , n51857 , n51858 );
xor ( n51860 , n51857 , n51858 );
xor ( n51861 , n51304 , n51404 );
and ( n51862 , n30329 , n51558 );
and ( n51863 , n51861 , n51862 );
xor ( n51864 , n51861 , n51862 );
xor ( n51865 , n51308 , n51402 );
and ( n51866 , n30334 , n51558 );
and ( n51867 , n51865 , n51866 );
xor ( n51868 , n51865 , n51866 );
xor ( n51869 , n51312 , n51400 );
and ( n51870 , n30339 , n51558 );
and ( n51871 , n51869 , n51870 );
xor ( n51872 , n51869 , n51870 );
xor ( n51873 , n51316 , n51398 );
and ( n51874 , n30344 , n51558 );
and ( n51875 , n51873 , n51874 );
xor ( n51876 , n51873 , n51874 );
xor ( n51877 , n51320 , n51396 );
and ( n51878 , n30349 , n51558 );
and ( n51879 , n51877 , n51878 );
xor ( n51880 , n51877 , n51878 );
xor ( n51881 , n51324 , n51394 );
and ( n51882 , n30354 , n51558 );
and ( n51883 , n51881 , n51882 );
xor ( n51884 , n51881 , n51882 );
xor ( n51885 , n51328 , n51392 );
and ( n51886 , n30359 , n51558 );
and ( n51887 , n51885 , n51886 );
xor ( n51888 , n51885 , n51886 );
xor ( n51889 , n51332 , n51390 );
and ( n51890 , n30364 , n51558 );
and ( n51891 , n51889 , n51890 );
xor ( n51892 , n51889 , n51890 );
xor ( n51893 , n51336 , n51388 );
and ( n51894 , n30369 , n51558 );
and ( n51895 , n51893 , n51894 );
xor ( n51896 , n51893 , n51894 );
xor ( n51897 , n51340 , n51386 );
and ( n51898 , n30374 , n51558 );
and ( n51899 , n51897 , n51898 );
xor ( n51900 , n51897 , n51898 );
xor ( n51901 , n51344 , n51384 );
and ( n51902 , n30379 , n51558 );
and ( n51903 , n51901 , n51902 );
xor ( n51904 , n51901 , n51902 );
xor ( n51905 , n51348 , n51382 );
and ( n51906 , n30384 , n51558 );
and ( n51907 , n51905 , n51906 );
xor ( n51908 , n51905 , n51906 );
xor ( n51909 , n51352 , n51380 );
and ( n51910 , n30389 , n51558 );
and ( n51911 , n51909 , n51910 );
xor ( n51912 , n51909 , n51910 );
xor ( n51913 , n51356 , n51378 );
and ( n51914 , n30394 , n51558 );
and ( n51915 , n51913 , n51914 );
xor ( n51916 , n51913 , n51914 );
xor ( n51917 , n51360 , n51376 );
and ( n51918 , n30399 , n51558 );
and ( n51919 , n51917 , n51918 );
xor ( n51920 , n51917 , n51918 );
xor ( n51921 , n51364 , n51374 );
and ( n51922 , n30404 , n51558 );
and ( n51923 , n51921 , n51922 );
xor ( n51924 , n51921 , n51922 );
xor ( n51925 , n51368 , n51372 );
and ( n51926 , n30409 , n51558 );
and ( n51927 , n51925 , n51926 );
buf ( n51928 , n51927 );
and ( n51929 , n51924 , n51928 );
or ( n51930 , n51923 , n51929 );
and ( n51931 , n51920 , n51930 );
or ( n51932 , n51919 , n51931 );
and ( n51933 , n51916 , n51932 );
or ( n51934 , n51915 , n51933 );
and ( n51935 , n51912 , n51934 );
or ( n51936 , n51911 , n51935 );
and ( n51937 , n51908 , n51936 );
or ( n51938 , n51907 , n51937 );
and ( n51939 , n51904 , n51938 );
or ( n51940 , n51903 , n51939 );
and ( n51941 , n51900 , n51940 );
or ( n51942 , n51899 , n51941 );
and ( n51943 , n51896 , n51942 );
or ( n51944 , n51895 , n51943 );
and ( n51945 , n51892 , n51944 );
or ( n51946 , n51891 , n51945 );
and ( n51947 , n51888 , n51946 );
or ( n51948 , n51887 , n51947 );
and ( n51949 , n51884 , n51948 );
or ( n51950 , n51883 , n51949 );
and ( n51951 , n51880 , n51950 );
or ( n51952 , n51879 , n51951 );
and ( n51953 , n51876 , n51952 );
or ( n51954 , n51875 , n51953 );
and ( n51955 , n51872 , n51954 );
or ( n51956 , n51871 , n51955 );
and ( n51957 , n51868 , n51956 );
or ( n51958 , n51867 , n51957 );
and ( n51959 , n51864 , n51958 );
or ( n51960 , n51863 , n51959 );
and ( n51961 , n51860 , n51960 );
or ( n51962 , n51859 , n51961 );
and ( n51963 , n51856 , n51962 );
or ( n51964 , n51855 , n51963 );
and ( n51965 , n51852 , n51964 );
or ( n51966 , n51851 , n51965 );
and ( n51967 , n51848 , n51966 );
or ( n51968 , n51847 , n51967 );
and ( n51969 , n51844 , n51968 );
or ( n51970 , n51843 , n51969 );
and ( n51971 , n51840 , n51970 );
or ( n51972 , n51839 , n51971 );
and ( n51973 , n51836 , n51972 );
or ( n51974 , n51835 , n51973 );
and ( n51975 , n51832 , n51974 );
or ( n51976 , n51831 , n51975 );
and ( n51977 , n51828 , n51976 );
or ( n51978 , n51827 , n51977 );
and ( n51979 , n51824 , n51978 );
or ( n51980 , n51823 , n51979 );
and ( n51981 , n51820 , n51980 );
or ( n51982 , n51819 , n51981 );
and ( n51983 , n51816 , n51982 );
or ( n51984 , n51815 , n51983 );
and ( n51985 , n51812 , n51984 );
or ( n51986 , n51811 , n51985 );
and ( n51987 , n51808 , n51986 );
or ( n51988 , n51807 , n51987 );
and ( n51989 , n51804 , n51988 );
or ( n51990 , n51803 , n51989 );
and ( n51991 , n51800 , n51990 );
or ( n51992 , n51799 , n51991 );
and ( n51993 , n51796 , n51992 );
or ( n51994 , n51795 , n51993 );
and ( n51995 , n51792 , n51994 );
or ( n51996 , n51791 , n51995 );
and ( n51997 , n51788 , n51996 );
or ( n51998 , n51787 , n51997 );
and ( n51999 , n51784 , n51998 );
or ( n52000 , n51783 , n51999 );
and ( n52001 , n51780 , n52000 );
or ( n52002 , n51779 , n52001 );
and ( n52003 , n51776 , n52002 );
or ( n52004 , n51775 , n52003 );
and ( n52005 , n51772 , n52004 );
or ( n52006 , n51771 , n52005 );
and ( n52007 , n51768 , n52006 );
or ( n52008 , n51767 , n52007 );
and ( n52009 , n51764 , n52008 );
or ( n52010 , n51763 , n52009 );
and ( n52011 , n51760 , n52010 );
or ( n52012 , n51759 , n52011 );
and ( n52013 , n51756 , n52012 );
or ( n52014 , n51755 , n52013 );
and ( n52015 , n51752 , n52014 );
or ( n52016 , n51751 , n52015 );
and ( n52017 , n51748 , n52016 );
or ( n52018 , n51747 , n52017 );
and ( n52019 , n51744 , n52018 );
or ( n52020 , n51743 , n52019 );
and ( n52021 , n51740 , n52020 );
or ( n52022 , n51739 , n52021 );
and ( n52023 , n51736 , n52022 );
or ( n52024 , n51735 , n52023 );
and ( n52025 , n51732 , n52024 );
or ( n52026 , n51731 , n52025 );
and ( n52027 , n51728 , n52026 );
or ( n52028 , n51727 , n52027 );
and ( n52029 , n51724 , n52028 );
or ( n52030 , n51723 , n52029 );
and ( n52031 , n51720 , n52030 );
or ( n52032 , n51719 , n52031 );
and ( n52033 , n51716 , n52032 );
or ( n52034 , n51715 , n52033 );
and ( n52035 , n51712 , n52034 );
or ( n52036 , n51711 , n52035 );
and ( n52037 , n51708 , n52036 );
or ( n52038 , n51707 , n52037 );
and ( n52039 , n51704 , n52038 );
or ( n52040 , n51703 , n52039 );
and ( n52041 , n51700 , n52040 );
or ( n52042 , n51699 , n52041 );
and ( n52043 , n51696 , n52042 );
or ( n52044 , n51695 , n52043 );
and ( n52045 , n51692 , n52044 );
or ( n52046 , n51691 , n52045 );
and ( n52047 , n51688 , n52046 );
or ( n52048 , n51687 , n52047 );
and ( n52049 , n51684 , n52048 );
or ( n52050 , n51683 , n52049 );
and ( n52051 , n51680 , n52050 );
or ( n52052 , n51679 , n52051 );
and ( n52053 , n51676 , n52052 );
or ( n52054 , n51675 , n52053 );
and ( n52055 , n51672 , n52054 );
or ( n52056 , n51671 , n52055 );
and ( n52057 , n51668 , n52056 );
or ( n52058 , n51667 , n52057 );
and ( n52059 , n51664 , n52058 );
or ( n52060 , n51663 , n52059 );
and ( n52061 , n51660 , n52060 );
or ( n52062 , n51659 , n52061 );
and ( n52063 , n51656 , n52062 );
or ( n52064 , n51655 , n52063 );
and ( n52065 , n51652 , n52064 );
or ( n52066 , n51651 , n52065 );
and ( n52067 , n51648 , n52066 );
or ( n52068 , n51647 , n52067 );
and ( n52069 , n51644 , n52068 );
or ( n52070 , n51643 , n52069 );
and ( n52071 , n51640 , n52070 );
or ( n52072 , n51639 , n52071 );
and ( n52073 , n51636 , n52072 );
or ( n52074 , n51635 , n52073 );
and ( n52075 , n51632 , n52074 );
or ( n52076 , n51631 , n52075 );
and ( n52077 , n51628 , n52076 );
or ( n52078 , n51627 , n52077 );
and ( n52079 , n51624 , n52078 );
or ( n52080 , n51623 , n52079 );
and ( n52081 , n51620 , n52080 );
or ( n52082 , n51619 , n52081 );
and ( n52083 , n51616 , n52082 );
or ( n52084 , n51615 , n52083 );
and ( n52085 , n51612 , n52084 );
or ( n52086 , n51611 , n52085 );
and ( n52087 , n51608 , n52086 );
or ( n52088 , n51607 , n52087 );
and ( n52089 , n51604 , n52088 );
or ( n52090 , n51603 , n52089 );
and ( n52091 , n51600 , n52090 );
or ( n52092 , n51599 , n52091 );
and ( n52093 , n51596 , n52092 );
or ( n52094 , n51595 , n52093 );
and ( n52095 , n51592 , n52094 );
or ( n52096 , n51591 , n52095 );
and ( n52097 , n51588 , n52096 );
or ( n52098 , n51587 , n52097 );
and ( n52099 , n51584 , n52098 );
or ( n52100 , n51583 , n52099 );
and ( n52101 , n51580 , n52100 );
or ( n52102 , n51579 , n52101 );
and ( n52103 , n51576 , n52102 );
or ( n52104 , n51575 , n52103 );
and ( n52105 , n51572 , n52104 );
or ( n52106 , n51571 , n52105 );
and ( n52107 , n51568 , n52106 );
or ( n52108 , n51567 , n52107 );
and ( n52109 , n51564 , n52108 );
or ( n52110 , n51563 , n52109 );
xor ( n52111 , n51560 , n52110 );
buf ( n52112 , n18036 );
and ( n52113 , n29954 , n52112 );
xor ( n52114 , n52111 , n52113 );
xor ( n52115 , n51564 , n52108 );
and ( n52116 , n29959 , n52112 );
and ( n52117 , n52115 , n52116 );
xor ( n52118 , n52115 , n52116 );
xor ( n52119 , n51568 , n52106 );
and ( n52120 , n29964 , n52112 );
and ( n52121 , n52119 , n52120 );
xor ( n52122 , n52119 , n52120 );
xor ( n52123 , n51572 , n52104 );
and ( n52124 , n29969 , n52112 );
and ( n52125 , n52123 , n52124 );
xor ( n52126 , n52123 , n52124 );
xor ( n52127 , n51576 , n52102 );
and ( n52128 , n29974 , n52112 );
and ( n52129 , n52127 , n52128 );
xor ( n52130 , n52127 , n52128 );
xor ( n52131 , n51580 , n52100 );
and ( n52132 , n29979 , n52112 );
and ( n52133 , n52131 , n52132 );
xor ( n52134 , n52131 , n52132 );
xor ( n52135 , n51584 , n52098 );
and ( n52136 , n29984 , n52112 );
and ( n52137 , n52135 , n52136 );
xor ( n52138 , n52135 , n52136 );
xor ( n52139 , n51588 , n52096 );
and ( n52140 , n29989 , n52112 );
and ( n52141 , n52139 , n52140 );
xor ( n52142 , n52139 , n52140 );
xor ( n52143 , n51592 , n52094 );
and ( n52144 , n29994 , n52112 );
and ( n52145 , n52143 , n52144 );
xor ( n52146 , n52143 , n52144 );
xor ( n52147 , n51596 , n52092 );
and ( n52148 , n29999 , n52112 );
and ( n52149 , n52147 , n52148 );
xor ( n52150 , n52147 , n52148 );
xor ( n52151 , n51600 , n52090 );
and ( n52152 , n30004 , n52112 );
and ( n52153 , n52151 , n52152 );
xor ( n52154 , n52151 , n52152 );
xor ( n52155 , n51604 , n52088 );
and ( n52156 , n30009 , n52112 );
and ( n52157 , n52155 , n52156 );
xor ( n52158 , n52155 , n52156 );
xor ( n52159 , n51608 , n52086 );
and ( n52160 , n30014 , n52112 );
and ( n52161 , n52159 , n52160 );
xor ( n52162 , n52159 , n52160 );
xor ( n52163 , n51612 , n52084 );
and ( n52164 , n30019 , n52112 );
and ( n52165 , n52163 , n52164 );
xor ( n52166 , n52163 , n52164 );
xor ( n52167 , n51616 , n52082 );
and ( n52168 , n30024 , n52112 );
and ( n52169 , n52167 , n52168 );
xor ( n52170 , n52167 , n52168 );
xor ( n52171 , n51620 , n52080 );
and ( n52172 , n30029 , n52112 );
and ( n52173 , n52171 , n52172 );
xor ( n52174 , n52171 , n52172 );
xor ( n52175 , n51624 , n52078 );
and ( n52176 , n30034 , n52112 );
and ( n52177 , n52175 , n52176 );
xor ( n52178 , n52175 , n52176 );
xor ( n52179 , n51628 , n52076 );
and ( n52180 , n30039 , n52112 );
and ( n52181 , n52179 , n52180 );
xor ( n52182 , n52179 , n52180 );
xor ( n52183 , n51632 , n52074 );
and ( n52184 , n30044 , n52112 );
and ( n52185 , n52183 , n52184 );
xor ( n52186 , n52183 , n52184 );
xor ( n52187 , n51636 , n52072 );
and ( n52188 , n30049 , n52112 );
and ( n52189 , n52187 , n52188 );
xor ( n52190 , n52187 , n52188 );
xor ( n52191 , n51640 , n52070 );
and ( n52192 , n30054 , n52112 );
and ( n52193 , n52191 , n52192 );
xor ( n52194 , n52191 , n52192 );
xor ( n52195 , n51644 , n52068 );
and ( n52196 , n30059 , n52112 );
and ( n52197 , n52195 , n52196 );
xor ( n52198 , n52195 , n52196 );
xor ( n52199 , n51648 , n52066 );
and ( n52200 , n30064 , n52112 );
and ( n52201 , n52199 , n52200 );
xor ( n52202 , n52199 , n52200 );
xor ( n52203 , n51652 , n52064 );
and ( n52204 , n30069 , n52112 );
and ( n52205 , n52203 , n52204 );
xor ( n52206 , n52203 , n52204 );
xor ( n52207 , n51656 , n52062 );
and ( n52208 , n30074 , n52112 );
and ( n52209 , n52207 , n52208 );
xor ( n52210 , n52207 , n52208 );
xor ( n52211 , n51660 , n52060 );
and ( n52212 , n30079 , n52112 );
and ( n52213 , n52211 , n52212 );
xor ( n52214 , n52211 , n52212 );
xor ( n52215 , n51664 , n52058 );
and ( n52216 , n30084 , n52112 );
and ( n52217 , n52215 , n52216 );
xor ( n52218 , n52215 , n52216 );
xor ( n52219 , n51668 , n52056 );
and ( n52220 , n30089 , n52112 );
and ( n52221 , n52219 , n52220 );
xor ( n52222 , n52219 , n52220 );
xor ( n52223 , n51672 , n52054 );
and ( n52224 , n30094 , n52112 );
and ( n52225 , n52223 , n52224 );
xor ( n52226 , n52223 , n52224 );
xor ( n52227 , n51676 , n52052 );
and ( n52228 , n30099 , n52112 );
and ( n52229 , n52227 , n52228 );
xor ( n52230 , n52227 , n52228 );
xor ( n52231 , n51680 , n52050 );
and ( n52232 , n30104 , n52112 );
and ( n52233 , n52231 , n52232 );
xor ( n52234 , n52231 , n52232 );
xor ( n52235 , n51684 , n52048 );
and ( n52236 , n30109 , n52112 );
and ( n52237 , n52235 , n52236 );
xor ( n52238 , n52235 , n52236 );
xor ( n52239 , n51688 , n52046 );
and ( n52240 , n30114 , n52112 );
and ( n52241 , n52239 , n52240 );
xor ( n52242 , n52239 , n52240 );
xor ( n52243 , n51692 , n52044 );
and ( n52244 , n30119 , n52112 );
and ( n52245 , n52243 , n52244 );
xor ( n52246 , n52243 , n52244 );
xor ( n52247 , n51696 , n52042 );
and ( n52248 , n30124 , n52112 );
and ( n52249 , n52247 , n52248 );
xor ( n52250 , n52247 , n52248 );
xor ( n52251 , n51700 , n52040 );
and ( n52252 , n30129 , n52112 );
and ( n52253 , n52251 , n52252 );
xor ( n52254 , n52251 , n52252 );
xor ( n52255 , n51704 , n52038 );
and ( n52256 , n30134 , n52112 );
and ( n52257 , n52255 , n52256 );
xor ( n52258 , n52255 , n52256 );
xor ( n52259 , n51708 , n52036 );
and ( n52260 , n30139 , n52112 );
and ( n52261 , n52259 , n52260 );
xor ( n52262 , n52259 , n52260 );
xor ( n52263 , n51712 , n52034 );
and ( n52264 , n30144 , n52112 );
and ( n52265 , n52263 , n52264 );
xor ( n52266 , n52263 , n52264 );
xor ( n52267 , n51716 , n52032 );
and ( n52268 , n30149 , n52112 );
and ( n52269 , n52267 , n52268 );
xor ( n52270 , n52267 , n52268 );
xor ( n52271 , n51720 , n52030 );
and ( n52272 , n30154 , n52112 );
and ( n52273 , n52271 , n52272 );
xor ( n52274 , n52271 , n52272 );
xor ( n52275 , n51724 , n52028 );
and ( n52276 , n30159 , n52112 );
and ( n52277 , n52275 , n52276 );
xor ( n52278 , n52275 , n52276 );
xor ( n52279 , n51728 , n52026 );
and ( n52280 , n30164 , n52112 );
and ( n52281 , n52279 , n52280 );
xor ( n52282 , n52279 , n52280 );
xor ( n52283 , n51732 , n52024 );
and ( n52284 , n30169 , n52112 );
and ( n52285 , n52283 , n52284 );
xor ( n52286 , n52283 , n52284 );
xor ( n52287 , n51736 , n52022 );
and ( n52288 , n30174 , n52112 );
and ( n52289 , n52287 , n52288 );
xor ( n52290 , n52287 , n52288 );
xor ( n52291 , n51740 , n52020 );
and ( n52292 , n30179 , n52112 );
and ( n52293 , n52291 , n52292 );
xor ( n52294 , n52291 , n52292 );
xor ( n52295 , n51744 , n52018 );
and ( n52296 , n30184 , n52112 );
and ( n52297 , n52295 , n52296 );
xor ( n52298 , n52295 , n52296 );
xor ( n52299 , n51748 , n52016 );
and ( n52300 , n30189 , n52112 );
and ( n52301 , n52299 , n52300 );
xor ( n52302 , n52299 , n52300 );
xor ( n52303 , n51752 , n52014 );
and ( n52304 , n30194 , n52112 );
and ( n52305 , n52303 , n52304 );
xor ( n52306 , n52303 , n52304 );
xor ( n52307 , n51756 , n52012 );
and ( n52308 , n30199 , n52112 );
and ( n52309 , n52307 , n52308 );
xor ( n52310 , n52307 , n52308 );
xor ( n52311 , n51760 , n52010 );
and ( n52312 , n30204 , n52112 );
and ( n52313 , n52311 , n52312 );
xor ( n52314 , n52311 , n52312 );
xor ( n52315 , n51764 , n52008 );
and ( n52316 , n30209 , n52112 );
and ( n52317 , n52315 , n52316 );
xor ( n52318 , n52315 , n52316 );
xor ( n52319 , n51768 , n52006 );
and ( n52320 , n30214 , n52112 );
and ( n52321 , n52319 , n52320 );
xor ( n52322 , n52319 , n52320 );
xor ( n52323 , n51772 , n52004 );
and ( n52324 , n30219 , n52112 );
and ( n52325 , n52323 , n52324 );
xor ( n52326 , n52323 , n52324 );
xor ( n52327 , n51776 , n52002 );
and ( n52328 , n30224 , n52112 );
and ( n52329 , n52327 , n52328 );
xor ( n52330 , n52327 , n52328 );
xor ( n52331 , n51780 , n52000 );
and ( n52332 , n30229 , n52112 );
and ( n52333 , n52331 , n52332 );
xor ( n52334 , n52331 , n52332 );
xor ( n52335 , n51784 , n51998 );
and ( n52336 , n30234 , n52112 );
and ( n52337 , n52335 , n52336 );
xor ( n52338 , n52335 , n52336 );
xor ( n52339 , n51788 , n51996 );
and ( n52340 , n30239 , n52112 );
and ( n52341 , n52339 , n52340 );
xor ( n52342 , n52339 , n52340 );
xor ( n52343 , n51792 , n51994 );
and ( n52344 , n30244 , n52112 );
and ( n52345 , n52343 , n52344 );
xor ( n52346 , n52343 , n52344 );
xor ( n52347 , n51796 , n51992 );
and ( n52348 , n30249 , n52112 );
and ( n52349 , n52347 , n52348 );
xor ( n52350 , n52347 , n52348 );
xor ( n52351 , n51800 , n51990 );
and ( n52352 , n30254 , n52112 );
and ( n52353 , n52351 , n52352 );
xor ( n52354 , n52351 , n52352 );
xor ( n52355 , n51804 , n51988 );
and ( n52356 , n30259 , n52112 );
and ( n52357 , n52355 , n52356 );
xor ( n52358 , n52355 , n52356 );
xor ( n52359 , n51808 , n51986 );
and ( n52360 , n30264 , n52112 );
and ( n52361 , n52359 , n52360 );
xor ( n52362 , n52359 , n52360 );
xor ( n52363 , n51812 , n51984 );
and ( n52364 , n30269 , n52112 );
and ( n52365 , n52363 , n52364 );
xor ( n52366 , n52363 , n52364 );
xor ( n52367 , n51816 , n51982 );
and ( n52368 , n30274 , n52112 );
and ( n52369 , n52367 , n52368 );
xor ( n52370 , n52367 , n52368 );
xor ( n52371 , n51820 , n51980 );
and ( n52372 , n30279 , n52112 );
and ( n52373 , n52371 , n52372 );
xor ( n52374 , n52371 , n52372 );
xor ( n52375 , n51824 , n51978 );
and ( n52376 , n30284 , n52112 );
and ( n52377 , n52375 , n52376 );
xor ( n52378 , n52375 , n52376 );
xor ( n52379 , n51828 , n51976 );
and ( n52380 , n30289 , n52112 );
and ( n52381 , n52379 , n52380 );
xor ( n52382 , n52379 , n52380 );
xor ( n52383 , n51832 , n51974 );
and ( n52384 , n30294 , n52112 );
and ( n52385 , n52383 , n52384 );
xor ( n52386 , n52383 , n52384 );
xor ( n52387 , n51836 , n51972 );
and ( n52388 , n30299 , n52112 );
and ( n52389 , n52387 , n52388 );
xor ( n52390 , n52387 , n52388 );
xor ( n52391 , n51840 , n51970 );
and ( n52392 , n30304 , n52112 );
and ( n52393 , n52391 , n52392 );
xor ( n52394 , n52391 , n52392 );
xor ( n52395 , n51844 , n51968 );
and ( n52396 , n30309 , n52112 );
and ( n52397 , n52395 , n52396 );
xor ( n52398 , n52395 , n52396 );
xor ( n52399 , n51848 , n51966 );
and ( n52400 , n30314 , n52112 );
and ( n52401 , n52399 , n52400 );
xor ( n52402 , n52399 , n52400 );
xor ( n52403 , n51852 , n51964 );
and ( n52404 , n30319 , n52112 );
and ( n52405 , n52403 , n52404 );
xor ( n52406 , n52403 , n52404 );
xor ( n52407 , n51856 , n51962 );
and ( n52408 , n30324 , n52112 );
and ( n52409 , n52407 , n52408 );
xor ( n52410 , n52407 , n52408 );
xor ( n52411 , n51860 , n51960 );
and ( n52412 , n30329 , n52112 );
and ( n52413 , n52411 , n52412 );
xor ( n52414 , n52411 , n52412 );
xor ( n52415 , n51864 , n51958 );
and ( n52416 , n30334 , n52112 );
and ( n52417 , n52415 , n52416 );
xor ( n52418 , n52415 , n52416 );
xor ( n52419 , n51868 , n51956 );
and ( n52420 , n30339 , n52112 );
and ( n52421 , n52419 , n52420 );
xor ( n52422 , n52419 , n52420 );
xor ( n52423 , n51872 , n51954 );
and ( n52424 , n30344 , n52112 );
and ( n52425 , n52423 , n52424 );
xor ( n52426 , n52423 , n52424 );
xor ( n52427 , n51876 , n51952 );
and ( n52428 , n30349 , n52112 );
and ( n52429 , n52427 , n52428 );
xor ( n52430 , n52427 , n52428 );
xor ( n52431 , n51880 , n51950 );
and ( n52432 , n30354 , n52112 );
and ( n52433 , n52431 , n52432 );
xor ( n52434 , n52431 , n52432 );
xor ( n52435 , n51884 , n51948 );
and ( n52436 , n30359 , n52112 );
and ( n52437 , n52435 , n52436 );
xor ( n52438 , n52435 , n52436 );
xor ( n52439 , n51888 , n51946 );
and ( n52440 , n30364 , n52112 );
and ( n52441 , n52439 , n52440 );
xor ( n52442 , n52439 , n52440 );
xor ( n52443 , n51892 , n51944 );
and ( n52444 , n30369 , n52112 );
and ( n52445 , n52443 , n52444 );
xor ( n52446 , n52443 , n52444 );
xor ( n52447 , n51896 , n51942 );
and ( n52448 , n30374 , n52112 );
and ( n52449 , n52447 , n52448 );
xor ( n52450 , n52447 , n52448 );
xor ( n52451 , n51900 , n51940 );
and ( n52452 , n30379 , n52112 );
and ( n52453 , n52451 , n52452 );
xor ( n52454 , n52451 , n52452 );
xor ( n52455 , n51904 , n51938 );
and ( n52456 , n30384 , n52112 );
and ( n52457 , n52455 , n52456 );
xor ( n52458 , n52455 , n52456 );
xor ( n52459 , n51908 , n51936 );
and ( n52460 , n30389 , n52112 );
and ( n52461 , n52459 , n52460 );
xor ( n52462 , n52459 , n52460 );
xor ( n52463 , n51912 , n51934 );
and ( n52464 , n30394 , n52112 );
and ( n52465 , n52463 , n52464 );
xor ( n52466 , n52463 , n52464 );
xor ( n52467 , n51916 , n51932 );
and ( n52468 , n30399 , n52112 );
and ( n52469 , n52467 , n52468 );
xor ( n52470 , n52467 , n52468 );
xor ( n52471 , n51920 , n51930 );
and ( n52472 , n30404 , n52112 );
and ( n52473 , n52471 , n52472 );
xor ( n52474 , n52471 , n52472 );
xor ( n52475 , n51924 , n51928 );
and ( n52476 , n30409 , n52112 );
and ( n52477 , n52475 , n52476 );
buf ( n52478 , n52477 );
and ( n52479 , n52474 , n52478 );
or ( n52480 , n52473 , n52479 );
and ( n52481 , n52470 , n52480 );
or ( n52482 , n52469 , n52481 );
and ( n52483 , n52466 , n52482 );
or ( n52484 , n52465 , n52483 );
and ( n52485 , n52462 , n52484 );
or ( n52486 , n52461 , n52485 );
and ( n52487 , n52458 , n52486 );
or ( n52488 , n52457 , n52487 );
and ( n52489 , n52454 , n52488 );
or ( n52490 , n52453 , n52489 );
and ( n52491 , n52450 , n52490 );
or ( n52492 , n52449 , n52491 );
and ( n52493 , n52446 , n52492 );
or ( n52494 , n52445 , n52493 );
and ( n52495 , n52442 , n52494 );
or ( n52496 , n52441 , n52495 );
and ( n52497 , n52438 , n52496 );
or ( n52498 , n52437 , n52497 );
and ( n52499 , n52434 , n52498 );
or ( n52500 , n52433 , n52499 );
and ( n52501 , n52430 , n52500 );
or ( n52502 , n52429 , n52501 );
and ( n52503 , n52426 , n52502 );
or ( n52504 , n52425 , n52503 );
and ( n52505 , n52422 , n52504 );
or ( n52506 , n52421 , n52505 );
and ( n52507 , n52418 , n52506 );
or ( n52508 , n52417 , n52507 );
and ( n52509 , n52414 , n52508 );
or ( n52510 , n52413 , n52509 );
and ( n52511 , n52410 , n52510 );
or ( n52512 , n52409 , n52511 );
and ( n52513 , n52406 , n52512 );
or ( n52514 , n52405 , n52513 );
and ( n52515 , n52402 , n52514 );
or ( n52516 , n52401 , n52515 );
and ( n52517 , n52398 , n52516 );
or ( n52518 , n52397 , n52517 );
and ( n52519 , n52394 , n52518 );
or ( n52520 , n52393 , n52519 );
and ( n52521 , n52390 , n52520 );
or ( n52522 , n52389 , n52521 );
and ( n52523 , n52386 , n52522 );
or ( n52524 , n52385 , n52523 );
and ( n52525 , n52382 , n52524 );
or ( n52526 , n52381 , n52525 );
and ( n52527 , n52378 , n52526 );
or ( n52528 , n52377 , n52527 );
and ( n52529 , n52374 , n52528 );
or ( n52530 , n52373 , n52529 );
and ( n52531 , n52370 , n52530 );
or ( n52532 , n52369 , n52531 );
and ( n52533 , n52366 , n52532 );
or ( n52534 , n52365 , n52533 );
and ( n52535 , n52362 , n52534 );
or ( n52536 , n52361 , n52535 );
and ( n52537 , n52358 , n52536 );
or ( n52538 , n52357 , n52537 );
and ( n52539 , n52354 , n52538 );
or ( n52540 , n52353 , n52539 );
and ( n52541 , n52350 , n52540 );
or ( n52542 , n52349 , n52541 );
and ( n52543 , n52346 , n52542 );
or ( n52544 , n52345 , n52543 );
and ( n52545 , n52342 , n52544 );
or ( n52546 , n52341 , n52545 );
and ( n52547 , n52338 , n52546 );
or ( n52548 , n52337 , n52547 );
and ( n52549 , n52334 , n52548 );
or ( n52550 , n52333 , n52549 );
and ( n52551 , n52330 , n52550 );
or ( n52552 , n52329 , n52551 );
and ( n52553 , n52326 , n52552 );
or ( n52554 , n52325 , n52553 );
and ( n52555 , n52322 , n52554 );
or ( n52556 , n52321 , n52555 );
and ( n52557 , n52318 , n52556 );
or ( n52558 , n52317 , n52557 );
and ( n52559 , n52314 , n52558 );
or ( n52560 , n52313 , n52559 );
and ( n52561 , n52310 , n52560 );
or ( n52562 , n52309 , n52561 );
and ( n52563 , n52306 , n52562 );
or ( n52564 , n52305 , n52563 );
and ( n52565 , n52302 , n52564 );
or ( n52566 , n52301 , n52565 );
and ( n52567 , n52298 , n52566 );
or ( n52568 , n52297 , n52567 );
and ( n52569 , n52294 , n52568 );
or ( n52570 , n52293 , n52569 );
and ( n52571 , n52290 , n52570 );
or ( n52572 , n52289 , n52571 );
and ( n52573 , n52286 , n52572 );
or ( n52574 , n52285 , n52573 );
and ( n52575 , n52282 , n52574 );
or ( n52576 , n52281 , n52575 );
and ( n52577 , n52278 , n52576 );
or ( n52578 , n52277 , n52577 );
and ( n52579 , n52274 , n52578 );
or ( n52580 , n52273 , n52579 );
and ( n52581 , n52270 , n52580 );
or ( n52582 , n52269 , n52581 );
and ( n52583 , n52266 , n52582 );
or ( n52584 , n52265 , n52583 );
and ( n52585 , n52262 , n52584 );
or ( n52586 , n52261 , n52585 );
and ( n52587 , n52258 , n52586 );
or ( n52588 , n52257 , n52587 );
and ( n52589 , n52254 , n52588 );
or ( n52590 , n52253 , n52589 );
and ( n52591 , n52250 , n52590 );
or ( n52592 , n52249 , n52591 );
and ( n52593 , n52246 , n52592 );
or ( n52594 , n52245 , n52593 );
and ( n52595 , n52242 , n52594 );
or ( n52596 , n52241 , n52595 );
and ( n52597 , n52238 , n52596 );
or ( n52598 , n52237 , n52597 );
and ( n52599 , n52234 , n52598 );
or ( n52600 , n52233 , n52599 );
and ( n52601 , n52230 , n52600 );
or ( n52602 , n52229 , n52601 );
and ( n52603 , n52226 , n52602 );
or ( n52604 , n52225 , n52603 );
and ( n52605 , n52222 , n52604 );
or ( n52606 , n52221 , n52605 );
and ( n52607 , n52218 , n52606 );
or ( n52608 , n52217 , n52607 );
and ( n52609 , n52214 , n52608 );
or ( n52610 , n52213 , n52609 );
and ( n52611 , n52210 , n52610 );
or ( n52612 , n52209 , n52611 );
and ( n52613 , n52206 , n52612 );
or ( n52614 , n52205 , n52613 );
and ( n52615 , n52202 , n52614 );
or ( n52616 , n52201 , n52615 );
and ( n52617 , n52198 , n52616 );
or ( n52618 , n52197 , n52617 );
and ( n52619 , n52194 , n52618 );
or ( n52620 , n52193 , n52619 );
and ( n52621 , n52190 , n52620 );
or ( n52622 , n52189 , n52621 );
and ( n52623 , n52186 , n52622 );
or ( n52624 , n52185 , n52623 );
and ( n52625 , n52182 , n52624 );
or ( n52626 , n52181 , n52625 );
and ( n52627 , n52178 , n52626 );
or ( n52628 , n52177 , n52627 );
and ( n52629 , n52174 , n52628 );
or ( n52630 , n52173 , n52629 );
and ( n52631 , n52170 , n52630 );
or ( n52632 , n52169 , n52631 );
and ( n52633 , n52166 , n52632 );
or ( n52634 , n52165 , n52633 );
and ( n52635 , n52162 , n52634 );
or ( n52636 , n52161 , n52635 );
and ( n52637 , n52158 , n52636 );
or ( n52638 , n52157 , n52637 );
and ( n52639 , n52154 , n52638 );
or ( n52640 , n52153 , n52639 );
and ( n52641 , n52150 , n52640 );
or ( n52642 , n52149 , n52641 );
and ( n52643 , n52146 , n52642 );
or ( n52644 , n52145 , n52643 );
and ( n52645 , n52142 , n52644 );
or ( n52646 , n52141 , n52645 );
and ( n52647 , n52138 , n52646 );
or ( n52648 , n52137 , n52647 );
and ( n52649 , n52134 , n52648 );
or ( n52650 , n52133 , n52649 );
and ( n52651 , n52130 , n52650 );
or ( n52652 , n52129 , n52651 );
and ( n52653 , n52126 , n52652 );
or ( n52654 , n52125 , n52653 );
and ( n52655 , n52122 , n52654 );
or ( n52656 , n52121 , n52655 );
and ( n52657 , n52118 , n52656 );
or ( n52658 , n52117 , n52657 );
xor ( n52659 , n52114 , n52658 );
buf ( n52660 , n18034 );
and ( n52661 , n29959 , n52660 );
xor ( n52662 , n52659 , n52661 );
xor ( n52663 , n52118 , n52656 );
and ( n52664 , n29964 , n52660 );
and ( n52665 , n52663 , n52664 );
xor ( n52666 , n52663 , n52664 );
xor ( n52667 , n52122 , n52654 );
and ( n52668 , n29969 , n52660 );
and ( n52669 , n52667 , n52668 );
xor ( n52670 , n52667 , n52668 );
xor ( n52671 , n52126 , n52652 );
and ( n52672 , n29974 , n52660 );
and ( n52673 , n52671 , n52672 );
xor ( n52674 , n52671 , n52672 );
xor ( n52675 , n52130 , n52650 );
and ( n52676 , n29979 , n52660 );
and ( n52677 , n52675 , n52676 );
xor ( n52678 , n52675 , n52676 );
xor ( n52679 , n52134 , n52648 );
and ( n52680 , n29984 , n52660 );
and ( n52681 , n52679 , n52680 );
xor ( n52682 , n52679 , n52680 );
xor ( n52683 , n52138 , n52646 );
and ( n52684 , n29989 , n52660 );
and ( n52685 , n52683 , n52684 );
xor ( n52686 , n52683 , n52684 );
xor ( n52687 , n52142 , n52644 );
and ( n52688 , n29994 , n52660 );
and ( n52689 , n52687 , n52688 );
xor ( n52690 , n52687 , n52688 );
xor ( n52691 , n52146 , n52642 );
and ( n52692 , n29999 , n52660 );
and ( n52693 , n52691 , n52692 );
xor ( n52694 , n52691 , n52692 );
xor ( n52695 , n52150 , n52640 );
and ( n52696 , n30004 , n52660 );
and ( n52697 , n52695 , n52696 );
xor ( n52698 , n52695 , n52696 );
xor ( n52699 , n52154 , n52638 );
and ( n52700 , n30009 , n52660 );
and ( n52701 , n52699 , n52700 );
xor ( n52702 , n52699 , n52700 );
xor ( n52703 , n52158 , n52636 );
and ( n52704 , n30014 , n52660 );
and ( n52705 , n52703 , n52704 );
xor ( n52706 , n52703 , n52704 );
xor ( n52707 , n52162 , n52634 );
and ( n52708 , n30019 , n52660 );
and ( n52709 , n52707 , n52708 );
xor ( n52710 , n52707 , n52708 );
xor ( n52711 , n52166 , n52632 );
and ( n52712 , n30024 , n52660 );
and ( n52713 , n52711 , n52712 );
xor ( n52714 , n52711 , n52712 );
xor ( n52715 , n52170 , n52630 );
and ( n52716 , n30029 , n52660 );
and ( n52717 , n52715 , n52716 );
xor ( n52718 , n52715 , n52716 );
xor ( n52719 , n52174 , n52628 );
and ( n52720 , n30034 , n52660 );
and ( n52721 , n52719 , n52720 );
xor ( n52722 , n52719 , n52720 );
xor ( n52723 , n52178 , n52626 );
and ( n52724 , n30039 , n52660 );
and ( n52725 , n52723 , n52724 );
xor ( n52726 , n52723 , n52724 );
xor ( n52727 , n52182 , n52624 );
and ( n52728 , n30044 , n52660 );
and ( n52729 , n52727 , n52728 );
xor ( n52730 , n52727 , n52728 );
xor ( n52731 , n52186 , n52622 );
and ( n52732 , n30049 , n52660 );
and ( n52733 , n52731 , n52732 );
xor ( n52734 , n52731 , n52732 );
xor ( n52735 , n52190 , n52620 );
and ( n52736 , n30054 , n52660 );
and ( n52737 , n52735 , n52736 );
xor ( n52738 , n52735 , n52736 );
xor ( n52739 , n52194 , n52618 );
and ( n52740 , n30059 , n52660 );
and ( n52741 , n52739 , n52740 );
xor ( n52742 , n52739 , n52740 );
xor ( n52743 , n52198 , n52616 );
and ( n52744 , n30064 , n52660 );
and ( n52745 , n52743 , n52744 );
xor ( n52746 , n52743 , n52744 );
xor ( n52747 , n52202 , n52614 );
and ( n52748 , n30069 , n52660 );
and ( n52749 , n52747 , n52748 );
xor ( n52750 , n52747 , n52748 );
xor ( n52751 , n52206 , n52612 );
and ( n52752 , n30074 , n52660 );
and ( n52753 , n52751 , n52752 );
xor ( n52754 , n52751 , n52752 );
xor ( n52755 , n52210 , n52610 );
and ( n52756 , n30079 , n52660 );
and ( n52757 , n52755 , n52756 );
xor ( n52758 , n52755 , n52756 );
xor ( n52759 , n52214 , n52608 );
and ( n52760 , n30084 , n52660 );
and ( n52761 , n52759 , n52760 );
xor ( n52762 , n52759 , n52760 );
xor ( n52763 , n52218 , n52606 );
and ( n52764 , n30089 , n52660 );
and ( n52765 , n52763 , n52764 );
xor ( n52766 , n52763 , n52764 );
xor ( n52767 , n52222 , n52604 );
and ( n52768 , n30094 , n52660 );
and ( n52769 , n52767 , n52768 );
xor ( n52770 , n52767 , n52768 );
xor ( n52771 , n52226 , n52602 );
and ( n52772 , n30099 , n52660 );
and ( n52773 , n52771 , n52772 );
xor ( n52774 , n52771 , n52772 );
xor ( n52775 , n52230 , n52600 );
and ( n52776 , n30104 , n52660 );
and ( n52777 , n52775 , n52776 );
xor ( n52778 , n52775 , n52776 );
xor ( n52779 , n52234 , n52598 );
and ( n52780 , n30109 , n52660 );
and ( n52781 , n52779 , n52780 );
xor ( n52782 , n52779 , n52780 );
xor ( n52783 , n52238 , n52596 );
and ( n52784 , n30114 , n52660 );
and ( n52785 , n52783 , n52784 );
xor ( n52786 , n52783 , n52784 );
xor ( n52787 , n52242 , n52594 );
and ( n52788 , n30119 , n52660 );
and ( n52789 , n52787 , n52788 );
xor ( n52790 , n52787 , n52788 );
xor ( n52791 , n52246 , n52592 );
and ( n52792 , n30124 , n52660 );
and ( n52793 , n52791 , n52792 );
xor ( n52794 , n52791 , n52792 );
xor ( n52795 , n52250 , n52590 );
and ( n52796 , n30129 , n52660 );
and ( n52797 , n52795 , n52796 );
xor ( n52798 , n52795 , n52796 );
xor ( n52799 , n52254 , n52588 );
and ( n52800 , n30134 , n52660 );
and ( n52801 , n52799 , n52800 );
xor ( n52802 , n52799 , n52800 );
xor ( n52803 , n52258 , n52586 );
and ( n52804 , n30139 , n52660 );
and ( n52805 , n52803 , n52804 );
xor ( n52806 , n52803 , n52804 );
xor ( n52807 , n52262 , n52584 );
and ( n52808 , n30144 , n52660 );
and ( n52809 , n52807 , n52808 );
xor ( n52810 , n52807 , n52808 );
xor ( n52811 , n52266 , n52582 );
and ( n52812 , n30149 , n52660 );
and ( n52813 , n52811 , n52812 );
xor ( n52814 , n52811 , n52812 );
xor ( n52815 , n52270 , n52580 );
and ( n52816 , n30154 , n52660 );
and ( n52817 , n52815 , n52816 );
xor ( n52818 , n52815 , n52816 );
xor ( n52819 , n52274 , n52578 );
and ( n52820 , n30159 , n52660 );
and ( n52821 , n52819 , n52820 );
xor ( n52822 , n52819 , n52820 );
xor ( n52823 , n52278 , n52576 );
and ( n52824 , n30164 , n52660 );
and ( n52825 , n52823 , n52824 );
xor ( n52826 , n52823 , n52824 );
xor ( n52827 , n52282 , n52574 );
and ( n52828 , n30169 , n52660 );
and ( n52829 , n52827 , n52828 );
xor ( n52830 , n52827 , n52828 );
xor ( n52831 , n52286 , n52572 );
and ( n52832 , n30174 , n52660 );
and ( n52833 , n52831 , n52832 );
xor ( n52834 , n52831 , n52832 );
xor ( n52835 , n52290 , n52570 );
and ( n52836 , n30179 , n52660 );
and ( n52837 , n52835 , n52836 );
xor ( n52838 , n52835 , n52836 );
xor ( n52839 , n52294 , n52568 );
and ( n52840 , n30184 , n52660 );
and ( n52841 , n52839 , n52840 );
xor ( n52842 , n52839 , n52840 );
xor ( n52843 , n52298 , n52566 );
and ( n52844 , n30189 , n52660 );
and ( n52845 , n52843 , n52844 );
xor ( n52846 , n52843 , n52844 );
xor ( n52847 , n52302 , n52564 );
and ( n52848 , n30194 , n52660 );
and ( n52849 , n52847 , n52848 );
xor ( n52850 , n52847 , n52848 );
xor ( n52851 , n52306 , n52562 );
and ( n52852 , n30199 , n52660 );
and ( n52853 , n52851 , n52852 );
xor ( n52854 , n52851 , n52852 );
xor ( n52855 , n52310 , n52560 );
and ( n52856 , n30204 , n52660 );
and ( n52857 , n52855 , n52856 );
xor ( n52858 , n52855 , n52856 );
xor ( n52859 , n52314 , n52558 );
and ( n52860 , n30209 , n52660 );
and ( n52861 , n52859 , n52860 );
xor ( n52862 , n52859 , n52860 );
xor ( n52863 , n52318 , n52556 );
and ( n52864 , n30214 , n52660 );
and ( n52865 , n52863 , n52864 );
xor ( n52866 , n52863 , n52864 );
xor ( n52867 , n52322 , n52554 );
and ( n52868 , n30219 , n52660 );
and ( n52869 , n52867 , n52868 );
xor ( n52870 , n52867 , n52868 );
xor ( n52871 , n52326 , n52552 );
and ( n52872 , n30224 , n52660 );
and ( n52873 , n52871 , n52872 );
xor ( n52874 , n52871 , n52872 );
xor ( n52875 , n52330 , n52550 );
and ( n52876 , n30229 , n52660 );
and ( n52877 , n52875 , n52876 );
xor ( n52878 , n52875 , n52876 );
xor ( n52879 , n52334 , n52548 );
and ( n52880 , n30234 , n52660 );
and ( n52881 , n52879 , n52880 );
xor ( n52882 , n52879 , n52880 );
xor ( n52883 , n52338 , n52546 );
and ( n52884 , n30239 , n52660 );
and ( n52885 , n52883 , n52884 );
xor ( n52886 , n52883 , n52884 );
xor ( n52887 , n52342 , n52544 );
and ( n52888 , n30244 , n52660 );
and ( n52889 , n52887 , n52888 );
xor ( n52890 , n52887 , n52888 );
xor ( n52891 , n52346 , n52542 );
and ( n52892 , n30249 , n52660 );
and ( n52893 , n52891 , n52892 );
xor ( n52894 , n52891 , n52892 );
xor ( n52895 , n52350 , n52540 );
and ( n52896 , n30254 , n52660 );
and ( n52897 , n52895 , n52896 );
xor ( n52898 , n52895 , n52896 );
xor ( n52899 , n52354 , n52538 );
and ( n52900 , n30259 , n52660 );
and ( n52901 , n52899 , n52900 );
xor ( n52902 , n52899 , n52900 );
xor ( n52903 , n52358 , n52536 );
and ( n52904 , n30264 , n52660 );
and ( n52905 , n52903 , n52904 );
xor ( n52906 , n52903 , n52904 );
xor ( n52907 , n52362 , n52534 );
and ( n52908 , n30269 , n52660 );
and ( n52909 , n52907 , n52908 );
xor ( n52910 , n52907 , n52908 );
xor ( n52911 , n52366 , n52532 );
and ( n52912 , n30274 , n52660 );
and ( n52913 , n52911 , n52912 );
xor ( n52914 , n52911 , n52912 );
xor ( n52915 , n52370 , n52530 );
and ( n52916 , n30279 , n52660 );
and ( n52917 , n52915 , n52916 );
xor ( n52918 , n52915 , n52916 );
xor ( n52919 , n52374 , n52528 );
and ( n52920 , n30284 , n52660 );
and ( n52921 , n52919 , n52920 );
xor ( n52922 , n52919 , n52920 );
xor ( n52923 , n52378 , n52526 );
and ( n52924 , n30289 , n52660 );
and ( n52925 , n52923 , n52924 );
xor ( n52926 , n52923 , n52924 );
xor ( n52927 , n52382 , n52524 );
and ( n52928 , n30294 , n52660 );
and ( n52929 , n52927 , n52928 );
xor ( n52930 , n52927 , n52928 );
xor ( n52931 , n52386 , n52522 );
and ( n52932 , n30299 , n52660 );
and ( n52933 , n52931 , n52932 );
xor ( n52934 , n52931 , n52932 );
xor ( n52935 , n52390 , n52520 );
and ( n52936 , n30304 , n52660 );
and ( n52937 , n52935 , n52936 );
xor ( n52938 , n52935 , n52936 );
xor ( n52939 , n52394 , n52518 );
and ( n52940 , n30309 , n52660 );
and ( n52941 , n52939 , n52940 );
xor ( n52942 , n52939 , n52940 );
xor ( n52943 , n52398 , n52516 );
and ( n52944 , n30314 , n52660 );
and ( n52945 , n52943 , n52944 );
xor ( n52946 , n52943 , n52944 );
xor ( n52947 , n52402 , n52514 );
and ( n52948 , n30319 , n52660 );
and ( n52949 , n52947 , n52948 );
xor ( n52950 , n52947 , n52948 );
xor ( n52951 , n52406 , n52512 );
and ( n52952 , n30324 , n52660 );
and ( n52953 , n52951 , n52952 );
xor ( n52954 , n52951 , n52952 );
xor ( n52955 , n52410 , n52510 );
and ( n52956 , n30329 , n52660 );
and ( n52957 , n52955 , n52956 );
xor ( n52958 , n52955 , n52956 );
xor ( n52959 , n52414 , n52508 );
and ( n52960 , n30334 , n52660 );
and ( n52961 , n52959 , n52960 );
xor ( n52962 , n52959 , n52960 );
xor ( n52963 , n52418 , n52506 );
and ( n52964 , n30339 , n52660 );
and ( n52965 , n52963 , n52964 );
xor ( n52966 , n52963 , n52964 );
xor ( n52967 , n52422 , n52504 );
and ( n52968 , n30344 , n52660 );
and ( n52969 , n52967 , n52968 );
xor ( n52970 , n52967 , n52968 );
xor ( n52971 , n52426 , n52502 );
and ( n52972 , n30349 , n52660 );
and ( n52973 , n52971 , n52972 );
xor ( n52974 , n52971 , n52972 );
xor ( n52975 , n52430 , n52500 );
and ( n52976 , n30354 , n52660 );
and ( n52977 , n52975 , n52976 );
xor ( n52978 , n52975 , n52976 );
xor ( n52979 , n52434 , n52498 );
and ( n52980 , n30359 , n52660 );
and ( n52981 , n52979 , n52980 );
xor ( n52982 , n52979 , n52980 );
xor ( n52983 , n52438 , n52496 );
and ( n52984 , n30364 , n52660 );
and ( n52985 , n52983 , n52984 );
xor ( n52986 , n52983 , n52984 );
xor ( n52987 , n52442 , n52494 );
and ( n52988 , n30369 , n52660 );
and ( n52989 , n52987 , n52988 );
xor ( n52990 , n52987 , n52988 );
xor ( n52991 , n52446 , n52492 );
and ( n52992 , n30374 , n52660 );
and ( n52993 , n52991 , n52992 );
xor ( n52994 , n52991 , n52992 );
xor ( n52995 , n52450 , n52490 );
and ( n52996 , n30379 , n52660 );
and ( n52997 , n52995 , n52996 );
xor ( n52998 , n52995 , n52996 );
xor ( n52999 , n52454 , n52488 );
and ( n53000 , n30384 , n52660 );
and ( n53001 , n52999 , n53000 );
xor ( n53002 , n52999 , n53000 );
xor ( n53003 , n52458 , n52486 );
and ( n53004 , n30389 , n52660 );
and ( n53005 , n53003 , n53004 );
xor ( n53006 , n53003 , n53004 );
xor ( n53007 , n52462 , n52484 );
and ( n53008 , n30394 , n52660 );
and ( n53009 , n53007 , n53008 );
xor ( n53010 , n53007 , n53008 );
xor ( n53011 , n52466 , n52482 );
and ( n53012 , n30399 , n52660 );
and ( n53013 , n53011 , n53012 );
xor ( n53014 , n53011 , n53012 );
xor ( n53015 , n52470 , n52480 );
and ( n53016 , n30404 , n52660 );
and ( n53017 , n53015 , n53016 );
xor ( n53018 , n53015 , n53016 );
xor ( n53019 , n52474 , n52478 );
and ( n53020 , n30409 , n52660 );
and ( n53021 , n53019 , n53020 );
buf ( n53022 , n53021 );
and ( n53023 , n53018 , n53022 );
or ( n53024 , n53017 , n53023 );
and ( n53025 , n53014 , n53024 );
or ( n53026 , n53013 , n53025 );
and ( n53027 , n53010 , n53026 );
or ( n53028 , n53009 , n53027 );
and ( n53029 , n53006 , n53028 );
or ( n53030 , n53005 , n53029 );
and ( n53031 , n53002 , n53030 );
or ( n53032 , n53001 , n53031 );
and ( n53033 , n52998 , n53032 );
or ( n53034 , n52997 , n53033 );
and ( n53035 , n52994 , n53034 );
or ( n53036 , n52993 , n53035 );
and ( n53037 , n52990 , n53036 );
or ( n53038 , n52989 , n53037 );
and ( n53039 , n52986 , n53038 );
or ( n53040 , n52985 , n53039 );
and ( n53041 , n52982 , n53040 );
or ( n53042 , n52981 , n53041 );
and ( n53043 , n52978 , n53042 );
or ( n53044 , n52977 , n53043 );
and ( n53045 , n52974 , n53044 );
or ( n53046 , n52973 , n53045 );
and ( n53047 , n52970 , n53046 );
or ( n53048 , n52969 , n53047 );
and ( n53049 , n52966 , n53048 );
or ( n53050 , n52965 , n53049 );
and ( n53051 , n52962 , n53050 );
or ( n53052 , n52961 , n53051 );
and ( n53053 , n52958 , n53052 );
or ( n53054 , n52957 , n53053 );
and ( n53055 , n52954 , n53054 );
or ( n53056 , n52953 , n53055 );
and ( n53057 , n52950 , n53056 );
or ( n53058 , n52949 , n53057 );
and ( n53059 , n52946 , n53058 );
or ( n53060 , n52945 , n53059 );
and ( n53061 , n52942 , n53060 );
or ( n53062 , n52941 , n53061 );
and ( n53063 , n52938 , n53062 );
or ( n53064 , n52937 , n53063 );
and ( n53065 , n52934 , n53064 );
or ( n53066 , n52933 , n53065 );
and ( n53067 , n52930 , n53066 );
or ( n53068 , n52929 , n53067 );
and ( n53069 , n52926 , n53068 );
or ( n53070 , n52925 , n53069 );
and ( n53071 , n52922 , n53070 );
or ( n53072 , n52921 , n53071 );
and ( n53073 , n52918 , n53072 );
or ( n53074 , n52917 , n53073 );
and ( n53075 , n52914 , n53074 );
or ( n53076 , n52913 , n53075 );
and ( n53077 , n52910 , n53076 );
or ( n53078 , n52909 , n53077 );
and ( n53079 , n52906 , n53078 );
or ( n53080 , n52905 , n53079 );
and ( n53081 , n52902 , n53080 );
or ( n53082 , n52901 , n53081 );
and ( n53083 , n52898 , n53082 );
or ( n53084 , n52897 , n53083 );
and ( n53085 , n52894 , n53084 );
or ( n53086 , n52893 , n53085 );
and ( n53087 , n52890 , n53086 );
or ( n53088 , n52889 , n53087 );
and ( n53089 , n52886 , n53088 );
or ( n53090 , n52885 , n53089 );
and ( n53091 , n52882 , n53090 );
or ( n53092 , n52881 , n53091 );
and ( n53093 , n52878 , n53092 );
or ( n53094 , n52877 , n53093 );
and ( n53095 , n52874 , n53094 );
or ( n53096 , n52873 , n53095 );
and ( n53097 , n52870 , n53096 );
or ( n53098 , n52869 , n53097 );
and ( n53099 , n52866 , n53098 );
or ( n53100 , n52865 , n53099 );
and ( n53101 , n52862 , n53100 );
or ( n53102 , n52861 , n53101 );
and ( n53103 , n52858 , n53102 );
or ( n53104 , n52857 , n53103 );
and ( n53105 , n52854 , n53104 );
or ( n53106 , n52853 , n53105 );
and ( n53107 , n52850 , n53106 );
or ( n53108 , n52849 , n53107 );
and ( n53109 , n52846 , n53108 );
or ( n53110 , n52845 , n53109 );
and ( n53111 , n52842 , n53110 );
or ( n53112 , n52841 , n53111 );
and ( n53113 , n52838 , n53112 );
or ( n53114 , n52837 , n53113 );
and ( n53115 , n52834 , n53114 );
or ( n53116 , n52833 , n53115 );
and ( n53117 , n52830 , n53116 );
or ( n53118 , n52829 , n53117 );
and ( n53119 , n52826 , n53118 );
or ( n53120 , n52825 , n53119 );
and ( n53121 , n52822 , n53120 );
or ( n53122 , n52821 , n53121 );
and ( n53123 , n52818 , n53122 );
or ( n53124 , n52817 , n53123 );
and ( n53125 , n52814 , n53124 );
or ( n53126 , n52813 , n53125 );
and ( n53127 , n52810 , n53126 );
or ( n53128 , n52809 , n53127 );
and ( n53129 , n52806 , n53128 );
or ( n53130 , n52805 , n53129 );
and ( n53131 , n52802 , n53130 );
or ( n53132 , n52801 , n53131 );
and ( n53133 , n52798 , n53132 );
or ( n53134 , n52797 , n53133 );
and ( n53135 , n52794 , n53134 );
or ( n53136 , n52793 , n53135 );
and ( n53137 , n52790 , n53136 );
or ( n53138 , n52789 , n53137 );
and ( n53139 , n52786 , n53138 );
or ( n53140 , n52785 , n53139 );
and ( n53141 , n52782 , n53140 );
or ( n53142 , n52781 , n53141 );
and ( n53143 , n52778 , n53142 );
or ( n53144 , n52777 , n53143 );
and ( n53145 , n52774 , n53144 );
or ( n53146 , n52773 , n53145 );
and ( n53147 , n52770 , n53146 );
or ( n53148 , n52769 , n53147 );
and ( n53149 , n52766 , n53148 );
or ( n53150 , n52765 , n53149 );
and ( n53151 , n52762 , n53150 );
or ( n53152 , n52761 , n53151 );
and ( n53153 , n52758 , n53152 );
or ( n53154 , n52757 , n53153 );
and ( n53155 , n52754 , n53154 );
or ( n53156 , n52753 , n53155 );
and ( n53157 , n52750 , n53156 );
or ( n53158 , n52749 , n53157 );
and ( n53159 , n52746 , n53158 );
or ( n53160 , n52745 , n53159 );
and ( n53161 , n52742 , n53160 );
or ( n53162 , n52741 , n53161 );
and ( n53163 , n52738 , n53162 );
or ( n53164 , n52737 , n53163 );
and ( n53165 , n52734 , n53164 );
or ( n53166 , n52733 , n53165 );
and ( n53167 , n52730 , n53166 );
or ( n53168 , n52729 , n53167 );
and ( n53169 , n52726 , n53168 );
or ( n53170 , n52725 , n53169 );
and ( n53171 , n52722 , n53170 );
or ( n53172 , n52721 , n53171 );
and ( n53173 , n52718 , n53172 );
or ( n53174 , n52717 , n53173 );
and ( n53175 , n52714 , n53174 );
or ( n53176 , n52713 , n53175 );
and ( n53177 , n52710 , n53176 );
or ( n53178 , n52709 , n53177 );
and ( n53179 , n52706 , n53178 );
or ( n53180 , n52705 , n53179 );
and ( n53181 , n52702 , n53180 );
or ( n53182 , n52701 , n53181 );
and ( n53183 , n52698 , n53182 );
or ( n53184 , n52697 , n53183 );
and ( n53185 , n52694 , n53184 );
or ( n53186 , n52693 , n53185 );
and ( n53187 , n52690 , n53186 );
or ( n53188 , n52689 , n53187 );
and ( n53189 , n52686 , n53188 );
or ( n53190 , n52685 , n53189 );
and ( n53191 , n52682 , n53190 );
or ( n53192 , n52681 , n53191 );
and ( n53193 , n52678 , n53192 );
or ( n53194 , n52677 , n53193 );
and ( n53195 , n52674 , n53194 );
or ( n53196 , n52673 , n53195 );
and ( n53197 , n52670 , n53196 );
or ( n53198 , n52669 , n53197 );
and ( n53199 , n52666 , n53198 );
or ( n53200 , n52665 , n53199 );
xor ( n53201 , n52662 , n53200 );
buf ( n53202 , n18032 );
and ( n53203 , n29964 , n53202 );
xor ( n53204 , n53201 , n53203 );
xor ( n53205 , n52666 , n53198 );
and ( n53206 , n29969 , n53202 );
and ( n53207 , n53205 , n53206 );
xor ( n53208 , n53205 , n53206 );
xor ( n53209 , n52670 , n53196 );
and ( n53210 , n29974 , n53202 );
and ( n53211 , n53209 , n53210 );
xor ( n53212 , n53209 , n53210 );
xor ( n53213 , n52674 , n53194 );
and ( n53214 , n29979 , n53202 );
and ( n53215 , n53213 , n53214 );
xor ( n53216 , n53213 , n53214 );
xor ( n53217 , n52678 , n53192 );
and ( n53218 , n29984 , n53202 );
and ( n53219 , n53217 , n53218 );
xor ( n53220 , n53217 , n53218 );
xor ( n53221 , n52682 , n53190 );
and ( n53222 , n29989 , n53202 );
and ( n53223 , n53221 , n53222 );
xor ( n53224 , n53221 , n53222 );
xor ( n53225 , n52686 , n53188 );
and ( n53226 , n29994 , n53202 );
and ( n53227 , n53225 , n53226 );
xor ( n53228 , n53225 , n53226 );
xor ( n53229 , n52690 , n53186 );
and ( n53230 , n29999 , n53202 );
and ( n53231 , n53229 , n53230 );
xor ( n53232 , n53229 , n53230 );
xor ( n53233 , n52694 , n53184 );
and ( n53234 , n30004 , n53202 );
and ( n53235 , n53233 , n53234 );
xor ( n53236 , n53233 , n53234 );
xor ( n53237 , n52698 , n53182 );
and ( n53238 , n30009 , n53202 );
and ( n53239 , n53237 , n53238 );
xor ( n53240 , n53237 , n53238 );
xor ( n53241 , n52702 , n53180 );
and ( n53242 , n30014 , n53202 );
and ( n53243 , n53241 , n53242 );
xor ( n53244 , n53241 , n53242 );
xor ( n53245 , n52706 , n53178 );
and ( n53246 , n30019 , n53202 );
and ( n53247 , n53245 , n53246 );
xor ( n53248 , n53245 , n53246 );
xor ( n53249 , n52710 , n53176 );
and ( n53250 , n30024 , n53202 );
and ( n53251 , n53249 , n53250 );
xor ( n53252 , n53249 , n53250 );
xor ( n53253 , n52714 , n53174 );
and ( n53254 , n30029 , n53202 );
and ( n53255 , n53253 , n53254 );
xor ( n53256 , n53253 , n53254 );
xor ( n53257 , n52718 , n53172 );
and ( n53258 , n30034 , n53202 );
and ( n53259 , n53257 , n53258 );
xor ( n53260 , n53257 , n53258 );
xor ( n53261 , n52722 , n53170 );
and ( n53262 , n30039 , n53202 );
and ( n53263 , n53261 , n53262 );
xor ( n53264 , n53261 , n53262 );
xor ( n53265 , n52726 , n53168 );
and ( n53266 , n30044 , n53202 );
and ( n53267 , n53265 , n53266 );
xor ( n53268 , n53265 , n53266 );
xor ( n53269 , n52730 , n53166 );
and ( n53270 , n30049 , n53202 );
and ( n53271 , n53269 , n53270 );
xor ( n53272 , n53269 , n53270 );
xor ( n53273 , n52734 , n53164 );
and ( n53274 , n30054 , n53202 );
and ( n53275 , n53273 , n53274 );
xor ( n53276 , n53273 , n53274 );
xor ( n53277 , n52738 , n53162 );
and ( n53278 , n30059 , n53202 );
and ( n53279 , n53277 , n53278 );
xor ( n53280 , n53277 , n53278 );
xor ( n53281 , n52742 , n53160 );
and ( n53282 , n30064 , n53202 );
and ( n53283 , n53281 , n53282 );
xor ( n53284 , n53281 , n53282 );
xor ( n53285 , n52746 , n53158 );
and ( n53286 , n30069 , n53202 );
and ( n53287 , n53285 , n53286 );
xor ( n53288 , n53285 , n53286 );
xor ( n53289 , n52750 , n53156 );
and ( n53290 , n30074 , n53202 );
and ( n53291 , n53289 , n53290 );
xor ( n53292 , n53289 , n53290 );
xor ( n53293 , n52754 , n53154 );
and ( n53294 , n30079 , n53202 );
and ( n53295 , n53293 , n53294 );
xor ( n53296 , n53293 , n53294 );
xor ( n53297 , n52758 , n53152 );
and ( n53298 , n30084 , n53202 );
and ( n53299 , n53297 , n53298 );
xor ( n53300 , n53297 , n53298 );
xor ( n53301 , n52762 , n53150 );
and ( n53302 , n30089 , n53202 );
and ( n53303 , n53301 , n53302 );
xor ( n53304 , n53301 , n53302 );
xor ( n53305 , n52766 , n53148 );
and ( n53306 , n30094 , n53202 );
and ( n53307 , n53305 , n53306 );
xor ( n53308 , n53305 , n53306 );
xor ( n53309 , n52770 , n53146 );
and ( n53310 , n30099 , n53202 );
and ( n53311 , n53309 , n53310 );
xor ( n53312 , n53309 , n53310 );
xor ( n53313 , n52774 , n53144 );
and ( n53314 , n30104 , n53202 );
and ( n53315 , n53313 , n53314 );
xor ( n53316 , n53313 , n53314 );
xor ( n53317 , n52778 , n53142 );
and ( n53318 , n30109 , n53202 );
and ( n53319 , n53317 , n53318 );
xor ( n53320 , n53317 , n53318 );
xor ( n53321 , n52782 , n53140 );
and ( n53322 , n30114 , n53202 );
and ( n53323 , n53321 , n53322 );
xor ( n53324 , n53321 , n53322 );
xor ( n53325 , n52786 , n53138 );
and ( n53326 , n30119 , n53202 );
and ( n53327 , n53325 , n53326 );
xor ( n53328 , n53325 , n53326 );
xor ( n53329 , n52790 , n53136 );
and ( n53330 , n30124 , n53202 );
and ( n53331 , n53329 , n53330 );
xor ( n53332 , n53329 , n53330 );
xor ( n53333 , n52794 , n53134 );
and ( n53334 , n30129 , n53202 );
and ( n53335 , n53333 , n53334 );
xor ( n53336 , n53333 , n53334 );
xor ( n53337 , n52798 , n53132 );
and ( n53338 , n30134 , n53202 );
and ( n53339 , n53337 , n53338 );
xor ( n53340 , n53337 , n53338 );
xor ( n53341 , n52802 , n53130 );
and ( n53342 , n30139 , n53202 );
and ( n53343 , n53341 , n53342 );
xor ( n53344 , n53341 , n53342 );
xor ( n53345 , n52806 , n53128 );
and ( n53346 , n30144 , n53202 );
and ( n53347 , n53345 , n53346 );
xor ( n53348 , n53345 , n53346 );
xor ( n53349 , n52810 , n53126 );
and ( n53350 , n30149 , n53202 );
and ( n53351 , n53349 , n53350 );
xor ( n53352 , n53349 , n53350 );
xor ( n53353 , n52814 , n53124 );
and ( n53354 , n30154 , n53202 );
and ( n53355 , n53353 , n53354 );
xor ( n53356 , n53353 , n53354 );
xor ( n53357 , n52818 , n53122 );
and ( n53358 , n30159 , n53202 );
and ( n53359 , n53357 , n53358 );
xor ( n53360 , n53357 , n53358 );
xor ( n53361 , n52822 , n53120 );
and ( n53362 , n30164 , n53202 );
and ( n53363 , n53361 , n53362 );
xor ( n53364 , n53361 , n53362 );
xor ( n53365 , n52826 , n53118 );
and ( n53366 , n30169 , n53202 );
and ( n53367 , n53365 , n53366 );
xor ( n53368 , n53365 , n53366 );
xor ( n53369 , n52830 , n53116 );
and ( n53370 , n30174 , n53202 );
and ( n53371 , n53369 , n53370 );
xor ( n53372 , n53369 , n53370 );
xor ( n53373 , n52834 , n53114 );
and ( n53374 , n30179 , n53202 );
and ( n53375 , n53373 , n53374 );
xor ( n53376 , n53373 , n53374 );
xor ( n53377 , n52838 , n53112 );
and ( n53378 , n30184 , n53202 );
and ( n53379 , n53377 , n53378 );
xor ( n53380 , n53377 , n53378 );
xor ( n53381 , n52842 , n53110 );
and ( n53382 , n30189 , n53202 );
and ( n53383 , n53381 , n53382 );
xor ( n53384 , n53381 , n53382 );
xor ( n53385 , n52846 , n53108 );
and ( n53386 , n30194 , n53202 );
and ( n53387 , n53385 , n53386 );
xor ( n53388 , n53385 , n53386 );
xor ( n53389 , n52850 , n53106 );
and ( n53390 , n30199 , n53202 );
and ( n53391 , n53389 , n53390 );
xor ( n53392 , n53389 , n53390 );
xor ( n53393 , n52854 , n53104 );
and ( n53394 , n30204 , n53202 );
and ( n53395 , n53393 , n53394 );
xor ( n53396 , n53393 , n53394 );
xor ( n53397 , n52858 , n53102 );
and ( n53398 , n30209 , n53202 );
and ( n53399 , n53397 , n53398 );
xor ( n53400 , n53397 , n53398 );
xor ( n53401 , n52862 , n53100 );
and ( n53402 , n30214 , n53202 );
and ( n53403 , n53401 , n53402 );
xor ( n53404 , n53401 , n53402 );
xor ( n53405 , n52866 , n53098 );
and ( n53406 , n30219 , n53202 );
and ( n53407 , n53405 , n53406 );
xor ( n53408 , n53405 , n53406 );
xor ( n53409 , n52870 , n53096 );
and ( n53410 , n30224 , n53202 );
and ( n53411 , n53409 , n53410 );
xor ( n53412 , n53409 , n53410 );
xor ( n53413 , n52874 , n53094 );
and ( n53414 , n30229 , n53202 );
and ( n53415 , n53413 , n53414 );
xor ( n53416 , n53413 , n53414 );
xor ( n53417 , n52878 , n53092 );
and ( n53418 , n30234 , n53202 );
and ( n53419 , n53417 , n53418 );
xor ( n53420 , n53417 , n53418 );
xor ( n53421 , n52882 , n53090 );
and ( n53422 , n30239 , n53202 );
and ( n53423 , n53421 , n53422 );
xor ( n53424 , n53421 , n53422 );
xor ( n53425 , n52886 , n53088 );
and ( n53426 , n30244 , n53202 );
and ( n53427 , n53425 , n53426 );
xor ( n53428 , n53425 , n53426 );
xor ( n53429 , n52890 , n53086 );
and ( n53430 , n30249 , n53202 );
and ( n53431 , n53429 , n53430 );
xor ( n53432 , n53429 , n53430 );
xor ( n53433 , n52894 , n53084 );
and ( n53434 , n30254 , n53202 );
and ( n53435 , n53433 , n53434 );
xor ( n53436 , n53433 , n53434 );
xor ( n53437 , n52898 , n53082 );
and ( n53438 , n30259 , n53202 );
and ( n53439 , n53437 , n53438 );
xor ( n53440 , n53437 , n53438 );
xor ( n53441 , n52902 , n53080 );
and ( n53442 , n30264 , n53202 );
and ( n53443 , n53441 , n53442 );
xor ( n53444 , n53441 , n53442 );
xor ( n53445 , n52906 , n53078 );
and ( n53446 , n30269 , n53202 );
and ( n53447 , n53445 , n53446 );
xor ( n53448 , n53445 , n53446 );
xor ( n53449 , n52910 , n53076 );
and ( n53450 , n30274 , n53202 );
and ( n53451 , n53449 , n53450 );
xor ( n53452 , n53449 , n53450 );
xor ( n53453 , n52914 , n53074 );
and ( n53454 , n30279 , n53202 );
and ( n53455 , n53453 , n53454 );
xor ( n53456 , n53453 , n53454 );
xor ( n53457 , n52918 , n53072 );
and ( n53458 , n30284 , n53202 );
and ( n53459 , n53457 , n53458 );
xor ( n53460 , n53457 , n53458 );
xor ( n53461 , n52922 , n53070 );
and ( n53462 , n30289 , n53202 );
and ( n53463 , n53461 , n53462 );
xor ( n53464 , n53461 , n53462 );
xor ( n53465 , n52926 , n53068 );
and ( n53466 , n30294 , n53202 );
and ( n53467 , n53465 , n53466 );
xor ( n53468 , n53465 , n53466 );
xor ( n53469 , n52930 , n53066 );
and ( n53470 , n30299 , n53202 );
and ( n53471 , n53469 , n53470 );
xor ( n53472 , n53469 , n53470 );
xor ( n53473 , n52934 , n53064 );
and ( n53474 , n30304 , n53202 );
and ( n53475 , n53473 , n53474 );
xor ( n53476 , n53473 , n53474 );
xor ( n53477 , n52938 , n53062 );
and ( n53478 , n30309 , n53202 );
and ( n53479 , n53477 , n53478 );
xor ( n53480 , n53477 , n53478 );
xor ( n53481 , n52942 , n53060 );
and ( n53482 , n30314 , n53202 );
and ( n53483 , n53481 , n53482 );
xor ( n53484 , n53481 , n53482 );
xor ( n53485 , n52946 , n53058 );
and ( n53486 , n30319 , n53202 );
and ( n53487 , n53485 , n53486 );
xor ( n53488 , n53485 , n53486 );
xor ( n53489 , n52950 , n53056 );
and ( n53490 , n30324 , n53202 );
and ( n53491 , n53489 , n53490 );
xor ( n53492 , n53489 , n53490 );
xor ( n53493 , n52954 , n53054 );
and ( n53494 , n30329 , n53202 );
and ( n53495 , n53493 , n53494 );
xor ( n53496 , n53493 , n53494 );
xor ( n53497 , n52958 , n53052 );
and ( n53498 , n30334 , n53202 );
and ( n53499 , n53497 , n53498 );
xor ( n53500 , n53497 , n53498 );
xor ( n53501 , n52962 , n53050 );
and ( n53502 , n30339 , n53202 );
and ( n53503 , n53501 , n53502 );
xor ( n53504 , n53501 , n53502 );
xor ( n53505 , n52966 , n53048 );
and ( n53506 , n30344 , n53202 );
and ( n53507 , n53505 , n53506 );
xor ( n53508 , n53505 , n53506 );
xor ( n53509 , n52970 , n53046 );
and ( n53510 , n30349 , n53202 );
and ( n53511 , n53509 , n53510 );
xor ( n53512 , n53509 , n53510 );
xor ( n53513 , n52974 , n53044 );
and ( n53514 , n30354 , n53202 );
and ( n53515 , n53513 , n53514 );
xor ( n53516 , n53513 , n53514 );
xor ( n53517 , n52978 , n53042 );
and ( n53518 , n30359 , n53202 );
and ( n53519 , n53517 , n53518 );
xor ( n53520 , n53517 , n53518 );
xor ( n53521 , n52982 , n53040 );
and ( n53522 , n30364 , n53202 );
and ( n53523 , n53521 , n53522 );
xor ( n53524 , n53521 , n53522 );
xor ( n53525 , n52986 , n53038 );
and ( n53526 , n30369 , n53202 );
and ( n53527 , n53525 , n53526 );
xor ( n53528 , n53525 , n53526 );
xor ( n53529 , n52990 , n53036 );
and ( n53530 , n30374 , n53202 );
and ( n53531 , n53529 , n53530 );
xor ( n53532 , n53529 , n53530 );
xor ( n53533 , n52994 , n53034 );
and ( n53534 , n30379 , n53202 );
and ( n53535 , n53533 , n53534 );
xor ( n53536 , n53533 , n53534 );
xor ( n53537 , n52998 , n53032 );
and ( n53538 , n30384 , n53202 );
and ( n53539 , n53537 , n53538 );
xor ( n53540 , n53537 , n53538 );
xor ( n53541 , n53002 , n53030 );
and ( n53542 , n30389 , n53202 );
and ( n53543 , n53541 , n53542 );
xor ( n53544 , n53541 , n53542 );
xor ( n53545 , n53006 , n53028 );
and ( n53546 , n30394 , n53202 );
and ( n53547 , n53545 , n53546 );
xor ( n53548 , n53545 , n53546 );
xor ( n53549 , n53010 , n53026 );
and ( n53550 , n30399 , n53202 );
and ( n53551 , n53549 , n53550 );
xor ( n53552 , n53549 , n53550 );
xor ( n53553 , n53014 , n53024 );
and ( n53554 , n30404 , n53202 );
and ( n53555 , n53553 , n53554 );
xor ( n53556 , n53553 , n53554 );
xor ( n53557 , n53018 , n53022 );
and ( n53558 , n30409 , n53202 );
and ( n53559 , n53557 , n53558 );
buf ( n53560 , n53559 );
and ( n53561 , n53556 , n53560 );
or ( n53562 , n53555 , n53561 );
and ( n53563 , n53552 , n53562 );
or ( n53564 , n53551 , n53563 );
and ( n53565 , n53548 , n53564 );
or ( n53566 , n53547 , n53565 );
and ( n53567 , n53544 , n53566 );
or ( n53568 , n53543 , n53567 );
and ( n53569 , n53540 , n53568 );
or ( n53570 , n53539 , n53569 );
and ( n53571 , n53536 , n53570 );
or ( n53572 , n53535 , n53571 );
and ( n53573 , n53532 , n53572 );
or ( n53574 , n53531 , n53573 );
and ( n53575 , n53528 , n53574 );
or ( n53576 , n53527 , n53575 );
and ( n53577 , n53524 , n53576 );
or ( n53578 , n53523 , n53577 );
and ( n53579 , n53520 , n53578 );
or ( n53580 , n53519 , n53579 );
and ( n53581 , n53516 , n53580 );
or ( n53582 , n53515 , n53581 );
and ( n53583 , n53512 , n53582 );
or ( n53584 , n53511 , n53583 );
and ( n53585 , n53508 , n53584 );
or ( n53586 , n53507 , n53585 );
and ( n53587 , n53504 , n53586 );
or ( n53588 , n53503 , n53587 );
and ( n53589 , n53500 , n53588 );
or ( n53590 , n53499 , n53589 );
and ( n53591 , n53496 , n53590 );
or ( n53592 , n53495 , n53591 );
and ( n53593 , n53492 , n53592 );
or ( n53594 , n53491 , n53593 );
and ( n53595 , n53488 , n53594 );
or ( n53596 , n53487 , n53595 );
and ( n53597 , n53484 , n53596 );
or ( n53598 , n53483 , n53597 );
and ( n53599 , n53480 , n53598 );
or ( n53600 , n53479 , n53599 );
and ( n53601 , n53476 , n53600 );
or ( n53602 , n53475 , n53601 );
and ( n53603 , n53472 , n53602 );
or ( n53604 , n53471 , n53603 );
and ( n53605 , n53468 , n53604 );
or ( n53606 , n53467 , n53605 );
and ( n53607 , n53464 , n53606 );
or ( n53608 , n53463 , n53607 );
and ( n53609 , n53460 , n53608 );
or ( n53610 , n53459 , n53609 );
and ( n53611 , n53456 , n53610 );
or ( n53612 , n53455 , n53611 );
and ( n53613 , n53452 , n53612 );
or ( n53614 , n53451 , n53613 );
and ( n53615 , n53448 , n53614 );
or ( n53616 , n53447 , n53615 );
and ( n53617 , n53444 , n53616 );
or ( n53618 , n53443 , n53617 );
and ( n53619 , n53440 , n53618 );
or ( n53620 , n53439 , n53619 );
and ( n53621 , n53436 , n53620 );
or ( n53622 , n53435 , n53621 );
and ( n53623 , n53432 , n53622 );
or ( n53624 , n53431 , n53623 );
and ( n53625 , n53428 , n53624 );
or ( n53626 , n53427 , n53625 );
and ( n53627 , n53424 , n53626 );
or ( n53628 , n53423 , n53627 );
and ( n53629 , n53420 , n53628 );
or ( n53630 , n53419 , n53629 );
and ( n53631 , n53416 , n53630 );
or ( n53632 , n53415 , n53631 );
and ( n53633 , n53412 , n53632 );
or ( n53634 , n53411 , n53633 );
and ( n53635 , n53408 , n53634 );
or ( n53636 , n53407 , n53635 );
and ( n53637 , n53404 , n53636 );
or ( n53638 , n53403 , n53637 );
and ( n53639 , n53400 , n53638 );
or ( n53640 , n53399 , n53639 );
and ( n53641 , n53396 , n53640 );
or ( n53642 , n53395 , n53641 );
and ( n53643 , n53392 , n53642 );
or ( n53644 , n53391 , n53643 );
and ( n53645 , n53388 , n53644 );
or ( n53646 , n53387 , n53645 );
and ( n53647 , n53384 , n53646 );
or ( n53648 , n53383 , n53647 );
and ( n53649 , n53380 , n53648 );
or ( n53650 , n53379 , n53649 );
and ( n53651 , n53376 , n53650 );
or ( n53652 , n53375 , n53651 );
and ( n53653 , n53372 , n53652 );
or ( n53654 , n53371 , n53653 );
and ( n53655 , n53368 , n53654 );
or ( n53656 , n53367 , n53655 );
and ( n53657 , n53364 , n53656 );
or ( n53658 , n53363 , n53657 );
and ( n53659 , n53360 , n53658 );
or ( n53660 , n53359 , n53659 );
and ( n53661 , n53356 , n53660 );
or ( n53662 , n53355 , n53661 );
and ( n53663 , n53352 , n53662 );
or ( n53664 , n53351 , n53663 );
and ( n53665 , n53348 , n53664 );
or ( n53666 , n53347 , n53665 );
and ( n53667 , n53344 , n53666 );
or ( n53668 , n53343 , n53667 );
and ( n53669 , n53340 , n53668 );
or ( n53670 , n53339 , n53669 );
and ( n53671 , n53336 , n53670 );
or ( n53672 , n53335 , n53671 );
and ( n53673 , n53332 , n53672 );
or ( n53674 , n53331 , n53673 );
and ( n53675 , n53328 , n53674 );
or ( n53676 , n53327 , n53675 );
and ( n53677 , n53324 , n53676 );
or ( n53678 , n53323 , n53677 );
and ( n53679 , n53320 , n53678 );
or ( n53680 , n53319 , n53679 );
and ( n53681 , n53316 , n53680 );
or ( n53682 , n53315 , n53681 );
and ( n53683 , n53312 , n53682 );
or ( n53684 , n53311 , n53683 );
and ( n53685 , n53308 , n53684 );
or ( n53686 , n53307 , n53685 );
and ( n53687 , n53304 , n53686 );
or ( n53688 , n53303 , n53687 );
and ( n53689 , n53300 , n53688 );
or ( n53690 , n53299 , n53689 );
and ( n53691 , n53296 , n53690 );
or ( n53692 , n53295 , n53691 );
and ( n53693 , n53292 , n53692 );
or ( n53694 , n53291 , n53693 );
and ( n53695 , n53288 , n53694 );
or ( n53696 , n53287 , n53695 );
and ( n53697 , n53284 , n53696 );
or ( n53698 , n53283 , n53697 );
and ( n53699 , n53280 , n53698 );
or ( n53700 , n53279 , n53699 );
and ( n53701 , n53276 , n53700 );
or ( n53702 , n53275 , n53701 );
and ( n53703 , n53272 , n53702 );
or ( n53704 , n53271 , n53703 );
and ( n53705 , n53268 , n53704 );
or ( n53706 , n53267 , n53705 );
and ( n53707 , n53264 , n53706 );
or ( n53708 , n53263 , n53707 );
and ( n53709 , n53260 , n53708 );
or ( n53710 , n53259 , n53709 );
and ( n53711 , n53256 , n53710 );
or ( n53712 , n53255 , n53711 );
and ( n53713 , n53252 , n53712 );
or ( n53714 , n53251 , n53713 );
and ( n53715 , n53248 , n53714 );
or ( n53716 , n53247 , n53715 );
and ( n53717 , n53244 , n53716 );
or ( n53718 , n53243 , n53717 );
and ( n53719 , n53240 , n53718 );
or ( n53720 , n53239 , n53719 );
and ( n53721 , n53236 , n53720 );
or ( n53722 , n53235 , n53721 );
and ( n53723 , n53232 , n53722 );
or ( n53724 , n53231 , n53723 );
and ( n53725 , n53228 , n53724 );
or ( n53726 , n53227 , n53725 );
and ( n53727 , n53224 , n53726 );
or ( n53728 , n53223 , n53727 );
and ( n53729 , n53220 , n53728 );
or ( n53730 , n53219 , n53729 );
and ( n53731 , n53216 , n53730 );
or ( n53732 , n53215 , n53731 );
and ( n53733 , n53212 , n53732 );
or ( n53734 , n53211 , n53733 );
and ( n53735 , n53208 , n53734 );
or ( n53736 , n53207 , n53735 );
xor ( n53737 , n53204 , n53736 );
buf ( n53738 , n18030 );
and ( n53739 , n29969 , n53738 );
xor ( n53740 , n53737 , n53739 );
xor ( n53741 , n53208 , n53734 );
and ( n53742 , n29974 , n53738 );
and ( n53743 , n53741 , n53742 );
xor ( n53744 , n53741 , n53742 );
xor ( n53745 , n53212 , n53732 );
and ( n53746 , n29979 , n53738 );
and ( n53747 , n53745 , n53746 );
xor ( n53748 , n53745 , n53746 );
xor ( n53749 , n53216 , n53730 );
and ( n53750 , n29984 , n53738 );
and ( n53751 , n53749 , n53750 );
xor ( n53752 , n53749 , n53750 );
xor ( n53753 , n53220 , n53728 );
and ( n53754 , n29989 , n53738 );
and ( n53755 , n53753 , n53754 );
xor ( n53756 , n53753 , n53754 );
xor ( n53757 , n53224 , n53726 );
and ( n53758 , n29994 , n53738 );
and ( n53759 , n53757 , n53758 );
xor ( n53760 , n53757 , n53758 );
xor ( n53761 , n53228 , n53724 );
and ( n53762 , n29999 , n53738 );
and ( n53763 , n53761 , n53762 );
xor ( n53764 , n53761 , n53762 );
xor ( n53765 , n53232 , n53722 );
and ( n53766 , n30004 , n53738 );
and ( n53767 , n53765 , n53766 );
xor ( n53768 , n53765 , n53766 );
xor ( n53769 , n53236 , n53720 );
and ( n53770 , n30009 , n53738 );
and ( n53771 , n53769 , n53770 );
xor ( n53772 , n53769 , n53770 );
xor ( n53773 , n53240 , n53718 );
and ( n53774 , n30014 , n53738 );
and ( n53775 , n53773 , n53774 );
xor ( n53776 , n53773 , n53774 );
xor ( n53777 , n53244 , n53716 );
and ( n53778 , n30019 , n53738 );
and ( n53779 , n53777 , n53778 );
xor ( n53780 , n53777 , n53778 );
xor ( n53781 , n53248 , n53714 );
and ( n53782 , n30024 , n53738 );
and ( n53783 , n53781 , n53782 );
xor ( n53784 , n53781 , n53782 );
xor ( n53785 , n53252 , n53712 );
and ( n53786 , n30029 , n53738 );
and ( n53787 , n53785 , n53786 );
xor ( n53788 , n53785 , n53786 );
xor ( n53789 , n53256 , n53710 );
and ( n53790 , n30034 , n53738 );
and ( n53791 , n53789 , n53790 );
xor ( n53792 , n53789 , n53790 );
xor ( n53793 , n53260 , n53708 );
and ( n53794 , n30039 , n53738 );
and ( n53795 , n53793 , n53794 );
xor ( n53796 , n53793 , n53794 );
xor ( n53797 , n53264 , n53706 );
and ( n53798 , n30044 , n53738 );
and ( n53799 , n53797 , n53798 );
xor ( n53800 , n53797 , n53798 );
xor ( n53801 , n53268 , n53704 );
and ( n53802 , n30049 , n53738 );
and ( n53803 , n53801 , n53802 );
xor ( n53804 , n53801 , n53802 );
xor ( n53805 , n53272 , n53702 );
and ( n53806 , n30054 , n53738 );
and ( n53807 , n53805 , n53806 );
xor ( n53808 , n53805 , n53806 );
xor ( n53809 , n53276 , n53700 );
and ( n53810 , n30059 , n53738 );
and ( n53811 , n53809 , n53810 );
xor ( n53812 , n53809 , n53810 );
xor ( n53813 , n53280 , n53698 );
and ( n53814 , n30064 , n53738 );
and ( n53815 , n53813 , n53814 );
xor ( n53816 , n53813 , n53814 );
xor ( n53817 , n53284 , n53696 );
and ( n53818 , n30069 , n53738 );
and ( n53819 , n53817 , n53818 );
xor ( n53820 , n53817 , n53818 );
xor ( n53821 , n53288 , n53694 );
and ( n53822 , n30074 , n53738 );
and ( n53823 , n53821 , n53822 );
xor ( n53824 , n53821 , n53822 );
xor ( n53825 , n53292 , n53692 );
and ( n53826 , n30079 , n53738 );
and ( n53827 , n53825 , n53826 );
xor ( n53828 , n53825 , n53826 );
xor ( n53829 , n53296 , n53690 );
and ( n53830 , n30084 , n53738 );
and ( n53831 , n53829 , n53830 );
xor ( n53832 , n53829 , n53830 );
xor ( n53833 , n53300 , n53688 );
and ( n53834 , n30089 , n53738 );
and ( n53835 , n53833 , n53834 );
xor ( n53836 , n53833 , n53834 );
xor ( n53837 , n53304 , n53686 );
and ( n53838 , n30094 , n53738 );
and ( n53839 , n53837 , n53838 );
xor ( n53840 , n53837 , n53838 );
xor ( n53841 , n53308 , n53684 );
and ( n53842 , n30099 , n53738 );
and ( n53843 , n53841 , n53842 );
xor ( n53844 , n53841 , n53842 );
xor ( n53845 , n53312 , n53682 );
and ( n53846 , n30104 , n53738 );
and ( n53847 , n53845 , n53846 );
xor ( n53848 , n53845 , n53846 );
xor ( n53849 , n53316 , n53680 );
and ( n53850 , n30109 , n53738 );
and ( n53851 , n53849 , n53850 );
xor ( n53852 , n53849 , n53850 );
xor ( n53853 , n53320 , n53678 );
and ( n53854 , n30114 , n53738 );
and ( n53855 , n53853 , n53854 );
xor ( n53856 , n53853 , n53854 );
xor ( n53857 , n53324 , n53676 );
and ( n53858 , n30119 , n53738 );
and ( n53859 , n53857 , n53858 );
xor ( n53860 , n53857 , n53858 );
xor ( n53861 , n53328 , n53674 );
and ( n53862 , n30124 , n53738 );
and ( n53863 , n53861 , n53862 );
xor ( n53864 , n53861 , n53862 );
xor ( n53865 , n53332 , n53672 );
and ( n53866 , n30129 , n53738 );
and ( n53867 , n53865 , n53866 );
xor ( n53868 , n53865 , n53866 );
xor ( n53869 , n53336 , n53670 );
and ( n53870 , n30134 , n53738 );
and ( n53871 , n53869 , n53870 );
xor ( n53872 , n53869 , n53870 );
xor ( n53873 , n53340 , n53668 );
and ( n53874 , n30139 , n53738 );
and ( n53875 , n53873 , n53874 );
xor ( n53876 , n53873 , n53874 );
xor ( n53877 , n53344 , n53666 );
and ( n53878 , n30144 , n53738 );
and ( n53879 , n53877 , n53878 );
xor ( n53880 , n53877 , n53878 );
xor ( n53881 , n53348 , n53664 );
and ( n53882 , n30149 , n53738 );
and ( n53883 , n53881 , n53882 );
xor ( n53884 , n53881 , n53882 );
xor ( n53885 , n53352 , n53662 );
and ( n53886 , n30154 , n53738 );
and ( n53887 , n53885 , n53886 );
xor ( n53888 , n53885 , n53886 );
xor ( n53889 , n53356 , n53660 );
and ( n53890 , n30159 , n53738 );
and ( n53891 , n53889 , n53890 );
xor ( n53892 , n53889 , n53890 );
xor ( n53893 , n53360 , n53658 );
and ( n53894 , n30164 , n53738 );
and ( n53895 , n53893 , n53894 );
xor ( n53896 , n53893 , n53894 );
xor ( n53897 , n53364 , n53656 );
and ( n53898 , n30169 , n53738 );
and ( n53899 , n53897 , n53898 );
xor ( n53900 , n53897 , n53898 );
xor ( n53901 , n53368 , n53654 );
and ( n53902 , n30174 , n53738 );
and ( n53903 , n53901 , n53902 );
xor ( n53904 , n53901 , n53902 );
xor ( n53905 , n53372 , n53652 );
and ( n53906 , n30179 , n53738 );
and ( n53907 , n53905 , n53906 );
xor ( n53908 , n53905 , n53906 );
xor ( n53909 , n53376 , n53650 );
and ( n53910 , n30184 , n53738 );
and ( n53911 , n53909 , n53910 );
xor ( n53912 , n53909 , n53910 );
xor ( n53913 , n53380 , n53648 );
and ( n53914 , n30189 , n53738 );
and ( n53915 , n53913 , n53914 );
xor ( n53916 , n53913 , n53914 );
xor ( n53917 , n53384 , n53646 );
and ( n53918 , n30194 , n53738 );
and ( n53919 , n53917 , n53918 );
xor ( n53920 , n53917 , n53918 );
xor ( n53921 , n53388 , n53644 );
and ( n53922 , n30199 , n53738 );
and ( n53923 , n53921 , n53922 );
xor ( n53924 , n53921 , n53922 );
xor ( n53925 , n53392 , n53642 );
and ( n53926 , n30204 , n53738 );
and ( n53927 , n53925 , n53926 );
xor ( n53928 , n53925 , n53926 );
xor ( n53929 , n53396 , n53640 );
and ( n53930 , n30209 , n53738 );
and ( n53931 , n53929 , n53930 );
xor ( n53932 , n53929 , n53930 );
xor ( n53933 , n53400 , n53638 );
and ( n53934 , n30214 , n53738 );
and ( n53935 , n53933 , n53934 );
xor ( n53936 , n53933 , n53934 );
xor ( n53937 , n53404 , n53636 );
and ( n53938 , n30219 , n53738 );
and ( n53939 , n53937 , n53938 );
xor ( n53940 , n53937 , n53938 );
xor ( n53941 , n53408 , n53634 );
and ( n53942 , n30224 , n53738 );
and ( n53943 , n53941 , n53942 );
xor ( n53944 , n53941 , n53942 );
xor ( n53945 , n53412 , n53632 );
and ( n53946 , n30229 , n53738 );
and ( n53947 , n53945 , n53946 );
xor ( n53948 , n53945 , n53946 );
xor ( n53949 , n53416 , n53630 );
and ( n53950 , n30234 , n53738 );
and ( n53951 , n53949 , n53950 );
xor ( n53952 , n53949 , n53950 );
xor ( n53953 , n53420 , n53628 );
and ( n53954 , n30239 , n53738 );
and ( n53955 , n53953 , n53954 );
xor ( n53956 , n53953 , n53954 );
xor ( n53957 , n53424 , n53626 );
and ( n53958 , n30244 , n53738 );
and ( n53959 , n53957 , n53958 );
xor ( n53960 , n53957 , n53958 );
xor ( n53961 , n53428 , n53624 );
and ( n53962 , n30249 , n53738 );
and ( n53963 , n53961 , n53962 );
xor ( n53964 , n53961 , n53962 );
xor ( n53965 , n53432 , n53622 );
and ( n53966 , n30254 , n53738 );
and ( n53967 , n53965 , n53966 );
xor ( n53968 , n53965 , n53966 );
xor ( n53969 , n53436 , n53620 );
and ( n53970 , n30259 , n53738 );
and ( n53971 , n53969 , n53970 );
xor ( n53972 , n53969 , n53970 );
xor ( n53973 , n53440 , n53618 );
and ( n53974 , n30264 , n53738 );
and ( n53975 , n53973 , n53974 );
xor ( n53976 , n53973 , n53974 );
xor ( n53977 , n53444 , n53616 );
and ( n53978 , n30269 , n53738 );
and ( n53979 , n53977 , n53978 );
xor ( n53980 , n53977 , n53978 );
xor ( n53981 , n53448 , n53614 );
and ( n53982 , n30274 , n53738 );
and ( n53983 , n53981 , n53982 );
xor ( n53984 , n53981 , n53982 );
xor ( n53985 , n53452 , n53612 );
and ( n53986 , n30279 , n53738 );
and ( n53987 , n53985 , n53986 );
xor ( n53988 , n53985 , n53986 );
xor ( n53989 , n53456 , n53610 );
and ( n53990 , n30284 , n53738 );
and ( n53991 , n53989 , n53990 );
xor ( n53992 , n53989 , n53990 );
xor ( n53993 , n53460 , n53608 );
and ( n53994 , n30289 , n53738 );
and ( n53995 , n53993 , n53994 );
xor ( n53996 , n53993 , n53994 );
xor ( n53997 , n53464 , n53606 );
and ( n53998 , n30294 , n53738 );
and ( n53999 , n53997 , n53998 );
xor ( n54000 , n53997 , n53998 );
xor ( n54001 , n53468 , n53604 );
and ( n54002 , n30299 , n53738 );
and ( n54003 , n54001 , n54002 );
xor ( n54004 , n54001 , n54002 );
xor ( n54005 , n53472 , n53602 );
and ( n54006 , n30304 , n53738 );
and ( n54007 , n54005 , n54006 );
xor ( n54008 , n54005 , n54006 );
xor ( n54009 , n53476 , n53600 );
and ( n54010 , n30309 , n53738 );
and ( n54011 , n54009 , n54010 );
xor ( n54012 , n54009 , n54010 );
xor ( n54013 , n53480 , n53598 );
and ( n54014 , n30314 , n53738 );
and ( n54015 , n54013 , n54014 );
xor ( n54016 , n54013 , n54014 );
xor ( n54017 , n53484 , n53596 );
and ( n54018 , n30319 , n53738 );
and ( n54019 , n54017 , n54018 );
xor ( n54020 , n54017 , n54018 );
xor ( n54021 , n53488 , n53594 );
and ( n54022 , n30324 , n53738 );
and ( n54023 , n54021 , n54022 );
xor ( n54024 , n54021 , n54022 );
xor ( n54025 , n53492 , n53592 );
and ( n54026 , n30329 , n53738 );
and ( n54027 , n54025 , n54026 );
xor ( n54028 , n54025 , n54026 );
xor ( n54029 , n53496 , n53590 );
and ( n54030 , n30334 , n53738 );
and ( n54031 , n54029 , n54030 );
xor ( n54032 , n54029 , n54030 );
xor ( n54033 , n53500 , n53588 );
and ( n54034 , n30339 , n53738 );
and ( n54035 , n54033 , n54034 );
xor ( n54036 , n54033 , n54034 );
xor ( n54037 , n53504 , n53586 );
and ( n54038 , n30344 , n53738 );
and ( n54039 , n54037 , n54038 );
xor ( n54040 , n54037 , n54038 );
xor ( n54041 , n53508 , n53584 );
and ( n54042 , n30349 , n53738 );
and ( n54043 , n54041 , n54042 );
xor ( n54044 , n54041 , n54042 );
xor ( n54045 , n53512 , n53582 );
and ( n54046 , n30354 , n53738 );
and ( n54047 , n54045 , n54046 );
xor ( n54048 , n54045 , n54046 );
xor ( n54049 , n53516 , n53580 );
and ( n54050 , n30359 , n53738 );
and ( n54051 , n54049 , n54050 );
xor ( n54052 , n54049 , n54050 );
xor ( n54053 , n53520 , n53578 );
and ( n54054 , n30364 , n53738 );
and ( n54055 , n54053 , n54054 );
xor ( n54056 , n54053 , n54054 );
xor ( n54057 , n53524 , n53576 );
and ( n54058 , n30369 , n53738 );
and ( n54059 , n54057 , n54058 );
xor ( n54060 , n54057 , n54058 );
xor ( n54061 , n53528 , n53574 );
and ( n54062 , n30374 , n53738 );
and ( n54063 , n54061 , n54062 );
xor ( n54064 , n54061 , n54062 );
xor ( n54065 , n53532 , n53572 );
and ( n54066 , n30379 , n53738 );
and ( n54067 , n54065 , n54066 );
xor ( n54068 , n54065 , n54066 );
xor ( n54069 , n53536 , n53570 );
and ( n54070 , n30384 , n53738 );
and ( n54071 , n54069 , n54070 );
xor ( n54072 , n54069 , n54070 );
xor ( n54073 , n53540 , n53568 );
and ( n54074 , n30389 , n53738 );
and ( n54075 , n54073 , n54074 );
xor ( n54076 , n54073 , n54074 );
xor ( n54077 , n53544 , n53566 );
and ( n54078 , n30394 , n53738 );
and ( n54079 , n54077 , n54078 );
xor ( n54080 , n54077 , n54078 );
xor ( n54081 , n53548 , n53564 );
and ( n54082 , n30399 , n53738 );
and ( n54083 , n54081 , n54082 );
xor ( n54084 , n54081 , n54082 );
xor ( n54085 , n53552 , n53562 );
and ( n54086 , n30404 , n53738 );
and ( n54087 , n54085 , n54086 );
xor ( n54088 , n54085 , n54086 );
xor ( n54089 , n53556 , n53560 );
and ( n54090 , n30409 , n53738 );
and ( n54091 , n54089 , n54090 );
buf ( n54092 , n54091 );
and ( n54093 , n54088 , n54092 );
or ( n54094 , n54087 , n54093 );
and ( n54095 , n54084 , n54094 );
or ( n54096 , n54083 , n54095 );
and ( n54097 , n54080 , n54096 );
or ( n54098 , n54079 , n54097 );
and ( n54099 , n54076 , n54098 );
or ( n54100 , n54075 , n54099 );
and ( n54101 , n54072 , n54100 );
or ( n54102 , n54071 , n54101 );
and ( n54103 , n54068 , n54102 );
or ( n54104 , n54067 , n54103 );
and ( n54105 , n54064 , n54104 );
or ( n54106 , n54063 , n54105 );
and ( n54107 , n54060 , n54106 );
or ( n54108 , n54059 , n54107 );
and ( n54109 , n54056 , n54108 );
or ( n54110 , n54055 , n54109 );
and ( n54111 , n54052 , n54110 );
or ( n54112 , n54051 , n54111 );
and ( n54113 , n54048 , n54112 );
or ( n54114 , n54047 , n54113 );
and ( n54115 , n54044 , n54114 );
or ( n54116 , n54043 , n54115 );
and ( n54117 , n54040 , n54116 );
or ( n54118 , n54039 , n54117 );
and ( n54119 , n54036 , n54118 );
or ( n54120 , n54035 , n54119 );
and ( n54121 , n54032 , n54120 );
or ( n54122 , n54031 , n54121 );
and ( n54123 , n54028 , n54122 );
or ( n54124 , n54027 , n54123 );
and ( n54125 , n54024 , n54124 );
or ( n54126 , n54023 , n54125 );
and ( n54127 , n54020 , n54126 );
or ( n54128 , n54019 , n54127 );
and ( n54129 , n54016 , n54128 );
or ( n54130 , n54015 , n54129 );
and ( n54131 , n54012 , n54130 );
or ( n54132 , n54011 , n54131 );
and ( n54133 , n54008 , n54132 );
or ( n54134 , n54007 , n54133 );
and ( n54135 , n54004 , n54134 );
or ( n54136 , n54003 , n54135 );
and ( n54137 , n54000 , n54136 );
or ( n54138 , n53999 , n54137 );
and ( n54139 , n53996 , n54138 );
or ( n54140 , n53995 , n54139 );
and ( n54141 , n53992 , n54140 );
or ( n54142 , n53991 , n54141 );
and ( n54143 , n53988 , n54142 );
or ( n54144 , n53987 , n54143 );
and ( n54145 , n53984 , n54144 );
or ( n54146 , n53983 , n54145 );
and ( n54147 , n53980 , n54146 );
or ( n54148 , n53979 , n54147 );
and ( n54149 , n53976 , n54148 );
or ( n54150 , n53975 , n54149 );
and ( n54151 , n53972 , n54150 );
or ( n54152 , n53971 , n54151 );
and ( n54153 , n53968 , n54152 );
or ( n54154 , n53967 , n54153 );
and ( n54155 , n53964 , n54154 );
or ( n54156 , n53963 , n54155 );
and ( n54157 , n53960 , n54156 );
or ( n54158 , n53959 , n54157 );
and ( n54159 , n53956 , n54158 );
or ( n54160 , n53955 , n54159 );
and ( n54161 , n53952 , n54160 );
or ( n54162 , n53951 , n54161 );
and ( n54163 , n53948 , n54162 );
or ( n54164 , n53947 , n54163 );
and ( n54165 , n53944 , n54164 );
or ( n54166 , n53943 , n54165 );
and ( n54167 , n53940 , n54166 );
or ( n54168 , n53939 , n54167 );
and ( n54169 , n53936 , n54168 );
or ( n54170 , n53935 , n54169 );
and ( n54171 , n53932 , n54170 );
or ( n54172 , n53931 , n54171 );
and ( n54173 , n53928 , n54172 );
or ( n54174 , n53927 , n54173 );
and ( n54175 , n53924 , n54174 );
or ( n54176 , n53923 , n54175 );
and ( n54177 , n53920 , n54176 );
or ( n54178 , n53919 , n54177 );
and ( n54179 , n53916 , n54178 );
or ( n54180 , n53915 , n54179 );
and ( n54181 , n53912 , n54180 );
or ( n54182 , n53911 , n54181 );
and ( n54183 , n53908 , n54182 );
or ( n54184 , n53907 , n54183 );
and ( n54185 , n53904 , n54184 );
or ( n54186 , n53903 , n54185 );
and ( n54187 , n53900 , n54186 );
or ( n54188 , n53899 , n54187 );
and ( n54189 , n53896 , n54188 );
or ( n54190 , n53895 , n54189 );
and ( n54191 , n53892 , n54190 );
or ( n54192 , n53891 , n54191 );
and ( n54193 , n53888 , n54192 );
or ( n54194 , n53887 , n54193 );
and ( n54195 , n53884 , n54194 );
or ( n54196 , n53883 , n54195 );
and ( n54197 , n53880 , n54196 );
or ( n54198 , n53879 , n54197 );
and ( n54199 , n53876 , n54198 );
or ( n54200 , n53875 , n54199 );
and ( n54201 , n53872 , n54200 );
or ( n54202 , n53871 , n54201 );
and ( n54203 , n53868 , n54202 );
or ( n54204 , n53867 , n54203 );
and ( n54205 , n53864 , n54204 );
or ( n54206 , n53863 , n54205 );
and ( n54207 , n53860 , n54206 );
or ( n54208 , n53859 , n54207 );
and ( n54209 , n53856 , n54208 );
or ( n54210 , n53855 , n54209 );
and ( n54211 , n53852 , n54210 );
or ( n54212 , n53851 , n54211 );
and ( n54213 , n53848 , n54212 );
or ( n54214 , n53847 , n54213 );
and ( n54215 , n53844 , n54214 );
or ( n54216 , n53843 , n54215 );
and ( n54217 , n53840 , n54216 );
or ( n54218 , n53839 , n54217 );
and ( n54219 , n53836 , n54218 );
or ( n54220 , n53835 , n54219 );
and ( n54221 , n53832 , n54220 );
or ( n54222 , n53831 , n54221 );
and ( n54223 , n53828 , n54222 );
or ( n54224 , n53827 , n54223 );
and ( n54225 , n53824 , n54224 );
or ( n54226 , n53823 , n54225 );
and ( n54227 , n53820 , n54226 );
or ( n54228 , n53819 , n54227 );
and ( n54229 , n53816 , n54228 );
or ( n54230 , n53815 , n54229 );
and ( n54231 , n53812 , n54230 );
or ( n54232 , n53811 , n54231 );
and ( n54233 , n53808 , n54232 );
or ( n54234 , n53807 , n54233 );
and ( n54235 , n53804 , n54234 );
or ( n54236 , n53803 , n54235 );
and ( n54237 , n53800 , n54236 );
or ( n54238 , n53799 , n54237 );
and ( n54239 , n53796 , n54238 );
or ( n54240 , n53795 , n54239 );
and ( n54241 , n53792 , n54240 );
or ( n54242 , n53791 , n54241 );
and ( n54243 , n53788 , n54242 );
or ( n54244 , n53787 , n54243 );
and ( n54245 , n53784 , n54244 );
or ( n54246 , n53783 , n54245 );
and ( n54247 , n53780 , n54246 );
or ( n54248 , n53779 , n54247 );
and ( n54249 , n53776 , n54248 );
or ( n54250 , n53775 , n54249 );
and ( n54251 , n53772 , n54250 );
or ( n54252 , n53771 , n54251 );
and ( n54253 , n53768 , n54252 );
or ( n54254 , n53767 , n54253 );
and ( n54255 , n53764 , n54254 );
or ( n54256 , n53763 , n54255 );
and ( n54257 , n53760 , n54256 );
or ( n54258 , n53759 , n54257 );
and ( n54259 , n53756 , n54258 );
or ( n54260 , n53755 , n54259 );
and ( n54261 , n53752 , n54260 );
or ( n54262 , n53751 , n54261 );
and ( n54263 , n53748 , n54262 );
or ( n54264 , n53747 , n54263 );
and ( n54265 , n53744 , n54264 );
or ( n54266 , n53743 , n54265 );
xor ( n54267 , n53740 , n54266 );
buf ( n54268 , n18028 );
and ( n54269 , n29974 , n54268 );
xor ( n54270 , n54267 , n54269 );
xor ( n54271 , n53744 , n54264 );
and ( n54272 , n29979 , n54268 );
and ( n54273 , n54271 , n54272 );
xor ( n54274 , n54271 , n54272 );
xor ( n54275 , n53748 , n54262 );
and ( n54276 , n29984 , n54268 );
and ( n54277 , n54275 , n54276 );
xor ( n54278 , n54275 , n54276 );
xor ( n54279 , n53752 , n54260 );
and ( n54280 , n29989 , n54268 );
and ( n54281 , n54279 , n54280 );
xor ( n54282 , n54279 , n54280 );
xor ( n54283 , n53756 , n54258 );
and ( n54284 , n29994 , n54268 );
and ( n54285 , n54283 , n54284 );
xor ( n54286 , n54283 , n54284 );
xor ( n54287 , n53760 , n54256 );
and ( n54288 , n29999 , n54268 );
and ( n54289 , n54287 , n54288 );
xor ( n54290 , n54287 , n54288 );
xor ( n54291 , n53764 , n54254 );
and ( n54292 , n30004 , n54268 );
and ( n54293 , n54291 , n54292 );
xor ( n54294 , n54291 , n54292 );
xor ( n54295 , n53768 , n54252 );
and ( n54296 , n30009 , n54268 );
and ( n54297 , n54295 , n54296 );
xor ( n54298 , n54295 , n54296 );
xor ( n54299 , n53772 , n54250 );
and ( n54300 , n30014 , n54268 );
and ( n54301 , n54299 , n54300 );
xor ( n54302 , n54299 , n54300 );
xor ( n54303 , n53776 , n54248 );
and ( n54304 , n30019 , n54268 );
and ( n54305 , n54303 , n54304 );
xor ( n54306 , n54303 , n54304 );
xor ( n54307 , n53780 , n54246 );
and ( n54308 , n30024 , n54268 );
and ( n54309 , n54307 , n54308 );
xor ( n54310 , n54307 , n54308 );
xor ( n54311 , n53784 , n54244 );
and ( n54312 , n30029 , n54268 );
and ( n54313 , n54311 , n54312 );
xor ( n54314 , n54311 , n54312 );
xor ( n54315 , n53788 , n54242 );
and ( n54316 , n30034 , n54268 );
and ( n54317 , n54315 , n54316 );
xor ( n54318 , n54315 , n54316 );
xor ( n54319 , n53792 , n54240 );
and ( n54320 , n30039 , n54268 );
and ( n54321 , n54319 , n54320 );
xor ( n54322 , n54319 , n54320 );
xor ( n54323 , n53796 , n54238 );
and ( n54324 , n30044 , n54268 );
and ( n54325 , n54323 , n54324 );
xor ( n54326 , n54323 , n54324 );
xor ( n54327 , n53800 , n54236 );
and ( n54328 , n30049 , n54268 );
and ( n54329 , n54327 , n54328 );
xor ( n54330 , n54327 , n54328 );
xor ( n54331 , n53804 , n54234 );
and ( n54332 , n30054 , n54268 );
and ( n54333 , n54331 , n54332 );
xor ( n54334 , n54331 , n54332 );
xor ( n54335 , n53808 , n54232 );
and ( n54336 , n30059 , n54268 );
and ( n54337 , n54335 , n54336 );
xor ( n54338 , n54335 , n54336 );
xor ( n54339 , n53812 , n54230 );
and ( n54340 , n30064 , n54268 );
and ( n54341 , n54339 , n54340 );
xor ( n54342 , n54339 , n54340 );
xor ( n54343 , n53816 , n54228 );
and ( n54344 , n30069 , n54268 );
and ( n54345 , n54343 , n54344 );
xor ( n54346 , n54343 , n54344 );
xor ( n54347 , n53820 , n54226 );
and ( n54348 , n30074 , n54268 );
and ( n54349 , n54347 , n54348 );
xor ( n54350 , n54347 , n54348 );
xor ( n54351 , n53824 , n54224 );
and ( n54352 , n30079 , n54268 );
and ( n54353 , n54351 , n54352 );
xor ( n54354 , n54351 , n54352 );
xor ( n54355 , n53828 , n54222 );
and ( n54356 , n30084 , n54268 );
and ( n54357 , n54355 , n54356 );
xor ( n54358 , n54355 , n54356 );
xor ( n54359 , n53832 , n54220 );
and ( n54360 , n30089 , n54268 );
and ( n54361 , n54359 , n54360 );
xor ( n54362 , n54359 , n54360 );
xor ( n54363 , n53836 , n54218 );
and ( n54364 , n30094 , n54268 );
and ( n54365 , n54363 , n54364 );
xor ( n54366 , n54363 , n54364 );
xor ( n54367 , n53840 , n54216 );
and ( n54368 , n30099 , n54268 );
and ( n54369 , n54367 , n54368 );
xor ( n54370 , n54367 , n54368 );
xor ( n54371 , n53844 , n54214 );
and ( n54372 , n30104 , n54268 );
and ( n54373 , n54371 , n54372 );
xor ( n54374 , n54371 , n54372 );
xor ( n54375 , n53848 , n54212 );
and ( n54376 , n30109 , n54268 );
and ( n54377 , n54375 , n54376 );
xor ( n54378 , n54375 , n54376 );
xor ( n54379 , n53852 , n54210 );
and ( n54380 , n30114 , n54268 );
and ( n54381 , n54379 , n54380 );
xor ( n54382 , n54379 , n54380 );
xor ( n54383 , n53856 , n54208 );
and ( n54384 , n30119 , n54268 );
and ( n54385 , n54383 , n54384 );
xor ( n54386 , n54383 , n54384 );
xor ( n54387 , n53860 , n54206 );
and ( n54388 , n30124 , n54268 );
and ( n54389 , n54387 , n54388 );
xor ( n54390 , n54387 , n54388 );
xor ( n54391 , n53864 , n54204 );
and ( n54392 , n30129 , n54268 );
and ( n54393 , n54391 , n54392 );
xor ( n54394 , n54391 , n54392 );
xor ( n54395 , n53868 , n54202 );
and ( n54396 , n30134 , n54268 );
and ( n54397 , n54395 , n54396 );
xor ( n54398 , n54395 , n54396 );
xor ( n54399 , n53872 , n54200 );
and ( n54400 , n30139 , n54268 );
and ( n54401 , n54399 , n54400 );
xor ( n54402 , n54399 , n54400 );
xor ( n54403 , n53876 , n54198 );
and ( n54404 , n30144 , n54268 );
and ( n54405 , n54403 , n54404 );
xor ( n54406 , n54403 , n54404 );
xor ( n54407 , n53880 , n54196 );
and ( n54408 , n30149 , n54268 );
and ( n54409 , n54407 , n54408 );
xor ( n54410 , n54407 , n54408 );
xor ( n54411 , n53884 , n54194 );
and ( n54412 , n30154 , n54268 );
and ( n54413 , n54411 , n54412 );
xor ( n54414 , n54411 , n54412 );
xor ( n54415 , n53888 , n54192 );
and ( n54416 , n30159 , n54268 );
and ( n54417 , n54415 , n54416 );
xor ( n54418 , n54415 , n54416 );
xor ( n54419 , n53892 , n54190 );
and ( n54420 , n30164 , n54268 );
and ( n54421 , n54419 , n54420 );
xor ( n54422 , n54419 , n54420 );
xor ( n54423 , n53896 , n54188 );
and ( n54424 , n30169 , n54268 );
and ( n54425 , n54423 , n54424 );
xor ( n54426 , n54423 , n54424 );
xor ( n54427 , n53900 , n54186 );
and ( n54428 , n30174 , n54268 );
and ( n54429 , n54427 , n54428 );
xor ( n54430 , n54427 , n54428 );
xor ( n54431 , n53904 , n54184 );
and ( n54432 , n30179 , n54268 );
and ( n54433 , n54431 , n54432 );
xor ( n54434 , n54431 , n54432 );
xor ( n54435 , n53908 , n54182 );
and ( n54436 , n30184 , n54268 );
and ( n54437 , n54435 , n54436 );
xor ( n54438 , n54435 , n54436 );
xor ( n54439 , n53912 , n54180 );
and ( n54440 , n30189 , n54268 );
and ( n54441 , n54439 , n54440 );
xor ( n54442 , n54439 , n54440 );
xor ( n54443 , n53916 , n54178 );
and ( n54444 , n30194 , n54268 );
and ( n54445 , n54443 , n54444 );
xor ( n54446 , n54443 , n54444 );
xor ( n54447 , n53920 , n54176 );
and ( n54448 , n30199 , n54268 );
and ( n54449 , n54447 , n54448 );
xor ( n54450 , n54447 , n54448 );
xor ( n54451 , n53924 , n54174 );
and ( n54452 , n30204 , n54268 );
and ( n54453 , n54451 , n54452 );
xor ( n54454 , n54451 , n54452 );
xor ( n54455 , n53928 , n54172 );
and ( n54456 , n30209 , n54268 );
and ( n54457 , n54455 , n54456 );
xor ( n54458 , n54455 , n54456 );
xor ( n54459 , n53932 , n54170 );
and ( n54460 , n30214 , n54268 );
and ( n54461 , n54459 , n54460 );
xor ( n54462 , n54459 , n54460 );
xor ( n54463 , n53936 , n54168 );
and ( n54464 , n30219 , n54268 );
and ( n54465 , n54463 , n54464 );
xor ( n54466 , n54463 , n54464 );
xor ( n54467 , n53940 , n54166 );
and ( n54468 , n30224 , n54268 );
and ( n54469 , n54467 , n54468 );
xor ( n54470 , n54467 , n54468 );
xor ( n54471 , n53944 , n54164 );
and ( n54472 , n30229 , n54268 );
and ( n54473 , n54471 , n54472 );
xor ( n54474 , n54471 , n54472 );
xor ( n54475 , n53948 , n54162 );
and ( n54476 , n30234 , n54268 );
and ( n54477 , n54475 , n54476 );
xor ( n54478 , n54475 , n54476 );
xor ( n54479 , n53952 , n54160 );
and ( n54480 , n30239 , n54268 );
and ( n54481 , n54479 , n54480 );
xor ( n54482 , n54479 , n54480 );
xor ( n54483 , n53956 , n54158 );
and ( n54484 , n30244 , n54268 );
and ( n54485 , n54483 , n54484 );
xor ( n54486 , n54483 , n54484 );
xor ( n54487 , n53960 , n54156 );
and ( n54488 , n30249 , n54268 );
and ( n54489 , n54487 , n54488 );
xor ( n54490 , n54487 , n54488 );
xor ( n54491 , n53964 , n54154 );
and ( n54492 , n30254 , n54268 );
and ( n54493 , n54491 , n54492 );
xor ( n54494 , n54491 , n54492 );
xor ( n54495 , n53968 , n54152 );
and ( n54496 , n30259 , n54268 );
and ( n54497 , n54495 , n54496 );
xor ( n54498 , n54495 , n54496 );
xor ( n54499 , n53972 , n54150 );
and ( n54500 , n30264 , n54268 );
and ( n54501 , n54499 , n54500 );
xor ( n54502 , n54499 , n54500 );
xor ( n54503 , n53976 , n54148 );
and ( n54504 , n30269 , n54268 );
and ( n54505 , n54503 , n54504 );
xor ( n54506 , n54503 , n54504 );
xor ( n54507 , n53980 , n54146 );
and ( n54508 , n30274 , n54268 );
and ( n54509 , n54507 , n54508 );
xor ( n54510 , n54507 , n54508 );
xor ( n54511 , n53984 , n54144 );
and ( n54512 , n30279 , n54268 );
and ( n54513 , n54511 , n54512 );
xor ( n54514 , n54511 , n54512 );
xor ( n54515 , n53988 , n54142 );
and ( n54516 , n30284 , n54268 );
and ( n54517 , n54515 , n54516 );
xor ( n54518 , n54515 , n54516 );
xor ( n54519 , n53992 , n54140 );
and ( n54520 , n30289 , n54268 );
and ( n54521 , n54519 , n54520 );
xor ( n54522 , n54519 , n54520 );
xor ( n54523 , n53996 , n54138 );
and ( n54524 , n30294 , n54268 );
and ( n54525 , n54523 , n54524 );
xor ( n54526 , n54523 , n54524 );
xor ( n54527 , n54000 , n54136 );
and ( n54528 , n30299 , n54268 );
and ( n54529 , n54527 , n54528 );
xor ( n54530 , n54527 , n54528 );
xor ( n54531 , n54004 , n54134 );
and ( n54532 , n30304 , n54268 );
and ( n54533 , n54531 , n54532 );
xor ( n54534 , n54531 , n54532 );
xor ( n54535 , n54008 , n54132 );
and ( n54536 , n30309 , n54268 );
and ( n54537 , n54535 , n54536 );
xor ( n54538 , n54535 , n54536 );
xor ( n54539 , n54012 , n54130 );
and ( n54540 , n30314 , n54268 );
and ( n54541 , n54539 , n54540 );
xor ( n54542 , n54539 , n54540 );
xor ( n54543 , n54016 , n54128 );
and ( n54544 , n30319 , n54268 );
and ( n54545 , n54543 , n54544 );
xor ( n54546 , n54543 , n54544 );
xor ( n54547 , n54020 , n54126 );
and ( n54548 , n30324 , n54268 );
and ( n54549 , n54547 , n54548 );
xor ( n54550 , n54547 , n54548 );
xor ( n54551 , n54024 , n54124 );
and ( n54552 , n30329 , n54268 );
and ( n54553 , n54551 , n54552 );
xor ( n54554 , n54551 , n54552 );
xor ( n54555 , n54028 , n54122 );
and ( n54556 , n30334 , n54268 );
and ( n54557 , n54555 , n54556 );
xor ( n54558 , n54555 , n54556 );
xor ( n54559 , n54032 , n54120 );
and ( n54560 , n30339 , n54268 );
and ( n54561 , n54559 , n54560 );
xor ( n54562 , n54559 , n54560 );
xor ( n54563 , n54036 , n54118 );
and ( n54564 , n30344 , n54268 );
and ( n54565 , n54563 , n54564 );
xor ( n54566 , n54563 , n54564 );
xor ( n54567 , n54040 , n54116 );
and ( n54568 , n30349 , n54268 );
and ( n54569 , n54567 , n54568 );
xor ( n54570 , n54567 , n54568 );
xor ( n54571 , n54044 , n54114 );
and ( n54572 , n30354 , n54268 );
and ( n54573 , n54571 , n54572 );
xor ( n54574 , n54571 , n54572 );
xor ( n54575 , n54048 , n54112 );
and ( n54576 , n30359 , n54268 );
and ( n54577 , n54575 , n54576 );
xor ( n54578 , n54575 , n54576 );
xor ( n54579 , n54052 , n54110 );
and ( n54580 , n30364 , n54268 );
and ( n54581 , n54579 , n54580 );
xor ( n54582 , n54579 , n54580 );
xor ( n54583 , n54056 , n54108 );
and ( n54584 , n30369 , n54268 );
and ( n54585 , n54583 , n54584 );
xor ( n54586 , n54583 , n54584 );
xor ( n54587 , n54060 , n54106 );
and ( n54588 , n30374 , n54268 );
and ( n54589 , n54587 , n54588 );
xor ( n54590 , n54587 , n54588 );
xor ( n54591 , n54064 , n54104 );
and ( n54592 , n30379 , n54268 );
and ( n54593 , n54591 , n54592 );
xor ( n54594 , n54591 , n54592 );
xor ( n54595 , n54068 , n54102 );
and ( n54596 , n30384 , n54268 );
and ( n54597 , n54595 , n54596 );
xor ( n54598 , n54595 , n54596 );
xor ( n54599 , n54072 , n54100 );
and ( n54600 , n30389 , n54268 );
and ( n54601 , n54599 , n54600 );
xor ( n54602 , n54599 , n54600 );
xor ( n54603 , n54076 , n54098 );
and ( n54604 , n30394 , n54268 );
and ( n54605 , n54603 , n54604 );
xor ( n54606 , n54603 , n54604 );
xor ( n54607 , n54080 , n54096 );
and ( n54608 , n30399 , n54268 );
and ( n54609 , n54607 , n54608 );
xor ( n54610 , n54607 , n54608 );
xor ( n54611 , n54084 , n54094 );
and ( n54612 , n30404 , n54268 );
and ( n54613 , n54611 , n54612 );
xor ( n54614 , n54611 , n54612 );
xor ( n54615 , n54088 , n54092 );
and ( n54616 , n30409 , n54268 );
and ( n54617 , n54615 , n54616 );
buf ( n54618 , n54617 );
and ( n54619 , n54614 , n54618 );
or ( n54620 , n54613 , n54619 );
and ( n54621 , n54610 , n54620 );
or ( n54622 , n54609 , n54621 );
and ( n54623 , n54606 , n54622 );
or ( n54624 , n54605 , n54623 );
and ( n54625 , n54602 , n54624 );
or ( n54626 , n54601 , n54625 );
and ( n54627 , n54598 , n54626 );
or ( n54628 , n54597 , n54627 );
and ( n54629 , n54594 , n54628 );
or ( n54630 , n54593 , n54629 );
and ( n54631 , n54590 , n54630 );
or ( n54632 , n54589 , n54631 );
and ( n54633 , n54586 , n54632 );
or ( n54634 , n54585 , n54633 );
and ( n54635 , n54582 , n54634 );
or ( n54636 , n54581 , n54635 );
and ( n54637 , n54578 , n54636 );
or ( n54638 , n54577 , n54637 );
and ( n54639 , n54574 , n54638 );
or ( n54640 , n54573 , n54639 );
and ( n54641 , n54570 , n54640 );
or ( n54642 , n54569 , n54641 );
and ( n54643 , n54566 , n54642 );
or ( n54644 , n54565 , n54643 );
and ( n54645 , n54562 , n54644 );
or ( n54646 , n54561 , n54645 );
and ( n54647 , n54558 , n54646 );
or ( n54648 , n54557 , n54647 );
and ( n54649 , n54554 , n54648 );
or ( n54650 , n54553 , n54649 );
and ( n54651 , n54550 , n54650 );
or ( n54652 , n54549 , n54651 );
and ( n54653 , n54546 , n54652 );
or ( n54654 , n54545 , n54653 );
and ( n54655 , n54542 , n54654 );
or ( n54656 , n54541 , n54655 );
and ( n54657 , n54538 , n54656 );
or ( n54658 , n54537 , n54657 );
and ( n54659 , n54534 , n54658 );
or ( n54660 , n54533 , n54659 );
and ( n54661 , n54530 , n54660 );
or ( n54662 , n54529 , n54661 );
and ( n54663 , n54526 , n54662 );
or ( n54664 , n54525 , n54663 );
and ( n54665 , n54522 , n54664 );
or ( n54666 , n54521 , n54665 );
and ( n54667 , n54518 , n54666 );
or ( n54668 , n54517 , n54667 );
and ( n54669 , n54514 , n54668 );
or ( n54670 , n54513 , n54669 );
and ( n54671 , n54510 , n54670 );
or ( n54672 , n54509 , n54671 );
and ( n54673 , n54506 , n54672 );
or ( n54674 , n54505 , n54673 );
and ( n54675 , n54502 , n54674 );
or ( n54676 , n54501 , n54675 );
and ( n54677 , n54498 , n54676 );
or ( n54678 , n54497 , n54677 );
and ( n54679 , n54494 , n54678 );
or ( n54680 , n54493 , n54679 );
and ( n54681 , n54490 , n54680 );
or ( n54682 , n54489 , n54681 );
and ( n54683 , n54486 , n54682 );
or ( n54684 , n54485 , n54683 );
and ( n54685 , n54482 , n54684 );
or ( n54686 , n54481 , n54685 );
and ( n54687 , n54478 , n54686 );
or ( n54688 , n54477 , n54687 );
and ( n54689 , n54474 , n54688 );
or ( n54690 , n54473 , n54689 );
and ( n54691 , n54470 , n54690 );
or ( n54692 , n54469 , n54691 );
and ( n54693 , n54466 , n54692 );
or ( n54694 , n54465 , n54693 );
and ( n54695 , n54462 , n54694 );
or ( n54696 , n54461 , n54695 );
and ( n54697 , n54458 , n54696 );
or ( n54698 , n54457 , n54697 );
and ( n54699 , n54454 , n54698 );
or ( n54700 , n54453 , n54699 );
and ( n54701 , n54450 , n54700 );
or ( n54702 , n54449 , n54701 );
and ( n54703 , n54446 , n54702 );
or ( n54704 , n54445 , n54703 );
and ( n54705 , n54442 , n54704 );
or ( n54706 , n54441 , n54705 );
and ( n54707 , n54438 , n54706 );
or ( n54708 , n54437 , n54707 );
and ( n54709 , n54434 , n54708 );
or ( n54710 , n54433 , n54709 );
and ( n54711 , n54430 , n54710 );
or ( n54712 , n54429 , n54711 );
and ( n54713 , n54426 , n54712 );
or ( n54714 , n54425 , n54713 );
and ( n54715 , n54422 , n54714 );
or ( n54716 , n54421 , n54715 );
and ( n54717 , n54418 , n54716 );
or ( n54718 , n54417 , n54717 );
and ( n54719 , n54414 , n54718 );
or ( n54720 , n54413 , n54719 );
and ( n54721 , n54410 , n54720 );
or ( n54722 , n54409 , n54721 );
and ( n54723 , n54406 , n54722 );
or ( n54724 , n54405 , n54723 );
and ( n54725 , n54402 , n54724 );
or ( n54726 , n54401 , n54725 );
and ( n54727 , n54398 , n54726 );
or ( n54728 , n54397 , n54727 );
and ( n54729 , n54394 , n54728 );
or ( n54730 , n54393 , n54729 );
and ( n54731 , n54390 , n54730 );
or ( n54732 , n54389 , n54731 );
and ( n54733 , n54386 , n54732 );
or ( n54734 , n54385 , n54733 );
and ( n54735 , n54382 , n54734 );
or ( n54736 , n54381 , n54735 );
and ( n54737 , n54378 , n54736 );
or ( n54738 , n54377 , n54737 );
and ( n54739 , n54374 , n54738 );
or ( n54740 , n54373 , n54739 );
and ( n54741 , n54370 , n54740 );
or ( n54742 , n54369 , n54741 );
and ( n54743 , n54366 , n54742 );
or ( n54744 , n54365 , n54743 );
and ( n54745 , n54362 , n54744 );
or ( n54746 , n54361 , n54745 );
and ( n54747 , n54358 , n54746 );
or ( n54748 , n54357 , n54747 );
and ( n54749 , n54354 , n54748 );
or ( n54750 , n54353 , n54749 );
and ( n54751 , n54350 , n54750 );
or ( n54752 , n54349 , n54751 );
and ( n54753 , n54346 , n54752 );
or ( n54754 , n54345 , n54753 );
and ( n54755 , n54342 , n54754 );
or ( n54756 , n54341 , n54755 );
and ( n54757 , n54338 , n54756 );
or ( n54758 , n54337 , n54757 );
and ( n54759 , n54334 , n54758 );
or ( n54760 , n54333 , n54759 );
and ( n54761 , n54330 , n54760 );
or ( n54762 , n54329 , n54761 );
and ( n54763 , n54326 , n54762 );
or ( n54764 , n54325 , n54763 );
and ( n54765 , n54322 , n54764 );
or ( n54766 , n54321 , n54765 );
and ( n54767 , n54318 , n54766 );
or ( n54768 , n54317 , n54767 );
and ( n54769 , n54314 , n54768 );
or ( n54770 , n54313 , n54769 );
and ( n54771 , n54310 , n54770 );
or ( n54772 , n54309 , n54771 );
and ( n54773 , n54306 , n54772 );
or ( n54774 , n54305 , n54773 );
and ( n54775 , n54302 , n54774 );
or ( n54776 , n54301 , n54775 );
and ( n54777 , n54298 , n54776 );
or ( n54778 , n54297 , n54777 );
and ( n54779 , n54294 , n54778 );
or ( n54780 , n54293 , n54779 );
and ( n54781 , n54290 , n54780 );
or ( n54782 , n54289 , n54781 );
and ( n54783 , n54286 , n54782 );
or ( n54784 , n54285 , n54783 );
and ( n54785 , n54282 , n54784 );
or ( n54786 , n54281 , n54785 );
and ( n54787 , n54278 , n54786 );
or ( n54788 , n54277 , n54787 );
and ( n54789 , n54274 , n54788 );
or ( n54790 , n54273 , n54789 );
xor ( n54791 , n54270 , n54790 );
buf ( n54792 , n18026 );
and ( n54793 , n29979 , n54792 );
xor ( n54794 , n54791 , n54793 );
xor ( n54795 , n54274 , n54788 );
and ( n54796 , n29984 , n54792 );
and ( n54797 , n54795 , n54796 );
xor ( n54798 , n54795 , n54796 );
xor ( n54799 , n54278 , n54786 );
and ( n54800 , n29989 , n54792 );
and ( n54801 , n54799 , n54800 );
xor ( n54802 , n54799 , n54800 );
xor ( n54803 , n54282 , n54784 );
and ( n54804 , n29994 , n54792 );
and ( n54805 , n54803 , n54804 );
xor ( n54806 , n54803 , n54804 );
xor ( n54807 , n54286 , n54782 );
and ( n54808 , n29999 , n54792 );
and ( n54809 , n54807 , n54808 );
xor ( n54810 , n54807 , n54808 );
xor ( n54811 , n54290 , n54780 );
and ( n54812 , n30004 , n54792 );
and ( n54813 , n54811 , n54812 );
xor ( n54814 , n54811 , n54812 );
xor ( n54815 , n54294 , n54778 );
and ( n54816 , n30009 , n54792 );
and ( n54817 , n54815 , n54816 );
xor ( n54818 , n54815 , n54816 );
xor ( n54819 , n54298 , n54776 );
and ( n54820 , n30014 , n54792 );
and ( n54821 , n54819 , n54820 );
xor ( n54822 , n54819 , n54820 );
xor ( n54823 , n54302 , n54774 );
and ( n54824 , n30019 , n54792 );
and ( n54825 , n54823 , n54824 );
xor ( n54826 , n54823 , n54824 );
xor ( n54827 , n54306 , n54772 );
and ( n54828 , n30024 , n54792 );
and ( n54829 , n54827 , n54828 );
xor ( n54830 , n54827 , n54828 );
xor ( n54831 , n54310 , n54770 );
and ( n54832 , n30029 , n54792 );
and ( n54833 , n54831 , n54832 );
xor ( n54834 , n54831 , n54832 );
xor ( n54835 , n54314 , n54768 );
and ( n54836 , n30034 , n54792 );
and ( n54837 , n54835 , n54836 );
xor ( n54838 , n54835 , n54836 );
xor ( n54839 , n54318 , n54766 );
and ( n54840 , n30039 , n54792 );
and ( n54841 , n54839 , n54840 );
xor ( n54842 , n54839 , n54840 );
xor ( n54843 , n54322 , n54764 );
and ( n54844 , n30044 , n54792 );
and ( n54845 , n54843 , n54844 );
xor ( n54846 , n54843 , n54844 );
xor ( n54847 , n54326 , n54762 );
and ( n54848 , n30049 , n54792 );
and ( n54849 , n54847 , n54848 );
xor ( n54850 , n54847 , n54848 );
xor ( n54851 , n54330 , n54760 );
and ( n54852 , n30054 , n54792 );
and ( n54853 , n54851 , n54852 );
xor ( n54854 , n54851 , n54852 );
xor ( n54855 , n54334 , n54758 );
and ( n54856 , n30059 , n54792 );
and ( n54857 , n54855 , n54856 );
xor ( n54858 , n54855 , n54856 );
xor ( n54859 , n54338 , n54756 );
and ( n54860 , n30064 , n54792 );
and ( n54861 , n54859 , n54860 );
xor ( n54862 , n54859 , n54860 );
xor ( n54863 , n54342 , n54754 );
and ( n54864 , n30069 , n54792 );
and ( n54865 , n54863 , n54864 );
xor ( n54866 , n54863 , n54864 );
xor ( n54867 , n54346 , n54752 );
and ( n54868 , n30074 , n54792 );
and ( n54869 , n54867 , n54868 );
xor ( n54870 , n54867 , n54868 );
xor ( n54871 , n54350 , n54750 );
and ( n54872 , n30079 , n54792 );
and ( n54873 , n54871 , n54872 );
xor ( n54874 , n54871 , n54872 );
xor ( n54875 , n54354 , n54748 );
and ( n54876 , n30084 , n54792 );
and ( n54877 , n54875 , n54876 );
xor ( n54878 , n54875 , n54876 );
xor ( n54879 , n54358 , n54746 );
and ( n54880 , n30089 , n54792 );
and ( n54881 , n54879 , n54880 );
xor ( n54882 , n54879 , n54880 );
xor ( n54883 , n54362 , n54744 );
and ( n54884 , n30094 , n54792 );
and ( n54885 , n54883 , n54884 );
xor ( n54886 , n54883 , n54884 );
xor ( n54887 , n54366 , n54742 );
and ( n54888 , n30099 , n54792 );
and ( n54889 , n54887 , n54888 );
xor ( n54890 , n54887 , n54888 );
xor ( n54891 , n54370 , n54740 );
and ( n54892 , n30104 , n54792 );
and ( n54893 , n54891 , n54892 );
xor ( n54894 , n54891 , n54892 );
xor ( n54895 , n54374 , n54738 );
and ( n54896 , n30109 , n54792 );
and ( n54897 , n54895 , n54896 );
xor ( n54898 , n54895 , n54896 );
xor ( n54899 , n54378 , n54736 );
and ( n54900 , n30114 , n54792 );
and ( n54901 , n54899 , n54900 );
xor ( n54902 , n54899 , n54900 );
xor ( n54903 , n54382 , n54734 );
and ( n54904 , n30119 , n54792 );
and ( n54905 , n54903 , n54904 );
xor ( n54906 , n54903 , n54904 );
xor ( n54907 , n54386 , n54732 );
and ( n54908 , n30124 , n54792 );
and ( n54909 , n54907 , n54908 );
xor ( n54910 , n54907 , n54908 );
xor ( n54911 , n54390 , n54730 );
and ( n54912 , n30129 , n54792 );
and ( n54913 , n54911 , n54912 );
xor ( n54914 , n54911 , n54912 );
xor ( n54915 , n54394 , n54728 );
and ( n54916 , n30134 , n54792 );
and ( n54917 , n54915 , n54916 );
xor ( n54918 , n54915 , n54916 );
xor ( n54919 , n54398 , n54726 );
and ( n54920 , n30139 , n54792 );
and ( n54921 , n54919 , n54920 );
xor ( n54922 , n54919 , n54920 );
xor ( n54923 , n54402 , n54724 );
and ( n54924 , n30144 , n54792 );
and ( n54925 , n54923 , n54924 );
xor ( n54926 , n54923 , n54924 );
xor ( n54927 , n54406 , n54722 );
and ( n54928 , n30149 , n54792 );
and ( n54929 , n54927 , n54928 );
xor ( n54930 , n54927 , n54928 );
xor ( n54931 , n54410 , n54720 );
and ( n54932 , n30154 , n54792 );
and ( n54933 , n54931 , n54932 );
xor ( n54934 , n54931 , n54932 );
xor ( n54935 , n54414 , n54718 );
and ( n54936 , n30159 , n54792 );
and ( n54937 , n54935 , n54936 );
xor ( n54938 , n54935 , n54936 );
xor ( n54939 , n54418 , n54716 );
and ( n54940 , n30164 , n54792 );
and ( n54941 , n54939 , n54940 );
xor ( n54942 , n54939 , n54940 );
xor ( n54943 , n54422 , n54714 );
and ( n54944 , n30169 , n54792 );
and ( n54945 , n54943 , n54944 );
xor ( n54946 , n54943 , n54944 );
xor ( n54947 , n54426 , n54712 );
and ( n54948 , n30174 , n54792 );
and ( n54949 , n54947 , n54948 );
xor ( n54950 , n54947 , n54948 );
xor ( n54951 , n54430 , n54710 );
and ( n54952 , n30179 , n54792 );
and ( n54953 , n54951 , n54952 );
xor ( n54954 , n54951 , n54952 );
xor ( n54955 , n54434 , n54708 );
and ( n54956 , n30184 , n54792 );
and ( n54957 , n54955 , n54956 );
xor ( n54958 , n54955 , n54956 );
xor ( n54959 , n54438 , n54706 );
and ( n54960 , n30189 , n54792 );
and ( n54961 , n54959 , n54960 );
xor ( n54962 , n54959 , n54960 );
xor ( n54963 , n54442 , n54704 );
and ( n54964 , n30194 , n54792 );
and ( n54965 , n54963 , n54964 );
xor ( n54966 , n54963 , n54964 );
xor ( n54967 , n54446 , n54702 );
and ( n54968 , n30199 , n54792 );
and ( n54969 , n54967 , n54968 );
xor ( n54970 , n54967 , n54968 );
xor ( n54971 , n54450 , n54700 );
and ( n54972 , n30204 , n54792 );
and ( n54973 , n54971 , n54972 );
xor ( n54974 , n54971 , n54972 );
xor ( n54975 , n54454 , n54698 );
and ( n54976 , n30209 , n54792 );
and ( n54977 , n54975 , n54976 );
xor ( n54978 , n54975 , n54976 );
xor ( n54979 , n54458 , n54696 );
and ( n54980 , n30214 , n54792 );
and ( n54981 , n54979 , n54980 );
xor ( n54982 , n54979 , n54980 );
xor ( n54983 , n54462 , n54694 );
and ( n54984 , n30219 , n54792 );
and ( n54985 , n54983 , n54984 );
xor ( n54986 , n54983 , n54984 );
xor ( n54987 , n54466 , n54692 );
and ( n54988 , n30224 , n54792 );
and ( n54989 , n54987 , n54988 );
xor ( n54990 , n54987 , n54988 );
xor ( n54991 , n54470 , n54690 );
and ( n54992 , n30229 , n54792 );
and ( n54993 , n54991 , n54992 );
xor ( n54994 , n54991 , n54992 );
xor ( n54995 , n54474 , n54688 );
and ( n54996 , n30234 , n54792 );
and ( n54997 , n54995 , n54996 );
xor ( n54998 , n54995 , n54996 );
xor ( n54999 , n54478 , n54686 );
and ( n55000 , n30239 , n54792 );
and ( n55001 , n54999 , n55000 );
xor ( n55002 , n54999 , n55000 );
xor ( n55003 , n54482 , n54684 );
and ( n55004 , n30244 , n54792 );
and ( n55005 , n55003 , n55004 );
xor ( n55006 , n55003 , n55004 );
xor ( n55007 , n54486 , n54682 );
and ( n55008 , n30249 , n54792 );
and ( n55009 , n55007 , n55008 );
xor ( n55010 , n55007 , n55008 );
xor ( n55011 , n54490 , n54680 );
and ( n55012 , n30254 , n54792 );
and ( n55013 , n55011 , n55012 );
xor ( n55014 , n55011 , n55012 );
xor ( n55015 , n54494 , n54678 );
and ( n55016 , n30259 , n54792 );
and ( n55017 , n55015 , n55016 );
xor ( n55018 , n55015 , n55016 );
xor ( n55019 , n54498 , n54676 );
and ( n55020 , n30264 , n54792 );
and ( n55021 , n55019 , n55020 );
xor ( n55022 , n55019 , n55020 );
xor ( n55023 , n54502 , n54674 );
and ( n55024 , n30269 , n54792 );
and ( n55025 , n55023 , n55024 );
xor ( n55026 , n55023 , n55024 );
xor ( n55027 , n54506 , n54672 );
and ( n55028 , n30274 , n54792 );
and ( n55029 , n55027 , n55028 );
xor ( n55030 , n55027 , n55028 );
xor ( n55031 , n54510 , n54670 );
and ( n55032 , n30279 , n54792 );
and ( n55033 , n55031 , n55032 );
xor ( n55034 , n55031 , n55032 );
xor ( n55035 , n54514 , n54668 );
and ( n55036 , n30284 , n54792 );
and ( n55037 , n55035 , n55036 );
xor ( n55038 , n55035 , n55036 );
xor ( n55039 , n54518 , n54666 );
and ( n55040 , n30289 , n54792 );
and ( n55041 , n55039 , n55040 );
xor ( n55042 , n55039 , n55040 );
xor ( n55043 , n54522 , n54664 );
and ( n55044 , n30294 , n54792 );
and ( n55045 , n55043 , n55044 );
xor ( n55046 , n55043 , n55044 );
xor ( n55047 , n54526 , n54662 );
and ( n55048 , n30299 , n54792 );
and ( n55049 , n55047 , n55048 );
xor ( n55050 , n55047 , n55048 );
xor ( n55051 , n54530 , n54660 );
and ( n55052 , n30304 , n54792 );
and ( n55053 , n55051 , n55052 );
xor ( n55054 , n55051 , n55052 );
xor ( n55055 , n54534 , n54658 );
and ( n55056 , n30309 , n54792 );
and ( n55057 , n55055 , n55056 );
xor ( n55058 , n55055 , n55056 );
xor ( n55059 , n54538 , n54656 );
and ( n55060 , n30314 , n54792 );
and ( n55061 , n55059 , n55060 );
xor ( n55062 , n55059 , n55060 );
xor ( n55063 , n54542 , n54654 );
and ( n55064 , n30319 , n54792 );
and ( n55065 , n55063 , n55064 );
xor ( n55066 , n55063 , n55064 );
xor ( n55067 , n54546 , n54652 );
and ( n55068 , n30324 , n54792 );
and ( n55069 , n55067 , n55068 );
xor ( n55070 , n55067 , n55068 );
xor ( n55071 , n54550 , n54650 );
and ( n55072 , n30329 , n54792 );
and ( n55073 , n55071 , n55072 );
xor ( n55074 , n55071 , n55072 );
xor ( n55075 , n54554 , n54648 );
and ( n55076 , n30334 , n54792 );
and ( n55077 , n55075 , n55076 );
xor ( n55078 , n55075 , n55076 );
xor ( n55079 , n54558 , n54646 );
and ( n55080 , n30339 , n54792 );
and ( n55081 , n55079 , n55080 );
xor ( n55082 , n55079 , n55080 );
xor ( n55083 , n54562 , n54644 );
and ( n55084 , n30344 , n54792 );
and ( n55085 , n55083 , n55084 );
xor ( n55086 , n55083 , n55084 );
xor ( n55087 , n54566 , n54642 );
and ( n55088 , n30349 , n54792 );
and ( n55089 , n55087 , n55088 );
xor ( n55090 , n55087 , n55088 );
xor ( n55091 , n54570 , n54640 );
and ( n55092 , n30354 , n54792 );
and ( n55093 , n55091 , n55092 );
xor ( n55094 , n55091 , n55092 );
xor ( n55095 , n54574 , n54638 );
and ( n55096 , n30359 , n54792 );
and ( n55097 , n55095 , n55096 );
xor ( n55098 , n55095 , n55096 );
xor ( n55099 , n54578 , n54636 );
and ( n55100 , n30364 , n54792 );
and ( n55101 , n55099 , n55100 );
xor ( n55102 , n55099 , n55100 );
xor ( n55103 , n54582 , n54634 );
and ( n55104 , n30369 , n54792 );
and ( n55105 , n55103 , n55104 );
xor ( n55106 , n55103 , n55104 );
xor ( n55107 , n54586 , n54632 );
and ( n55108 , n30374 , n54792 );
and ( n55109 , n55107 , n55108 );
xor ( n55110 , n55107 , n55108 );
xor ( n55111 , n54590 , n54630 );
and ( n55112 , n30379 , n54792 );
and ( n55113 , n55111 , n55112 );
xor ( n55114 , n55111 , n55112 );
xor ( n55115 , n54594 , n54628 );
and ( n55116 , n30384 , n54792 );
and ( n55117 , n55115 , n55116 );
xor ( n55118 , n55115 , n55116 );
xor ( n55119 , n54598 , n54626 );
and ( n55120 , n30389 , n54792 );
and ( n55121 , n55119 , n55120 );
xor ( n55122 , n55119 , n55120 );
xor ( n55123 , n54602 , n54624 );
and ( n55124 , n30394 , n54792 );
and ( n55125 , n55123 , n55124 );
xor ( n55126 , n55123 , n55124 );
xor ( n55127 , n54606 , n54622 );
and ( n55128 , n30399 , n54792 );
and ( n55129 , n55127 , n55128 );
xor ( n55130 , n55127 , n55128 );
xor ( n55131 , n54610 , n54620 );
and ( n55132 , n30404 , n54792 );
and ( n55133 , n55131 , n55132 );
xor ( n55134 , n55131 , n55132 );
xor ( n55135 , n54614 , n54618 );
and ( n55136 , n30409 , n54792 );
and ( n55137 , n55135 , n55136 );
buf ( n55138 , n55137 );
and ( n55139 , n55134 , n55138 );
or ( n55140 , n55133 , n55139 );
and ( n55141 , n55130 , n55140 );
or ( n55142 , n55129 , n55141 );
and ( n55143 , n55126 , n55142 );
or ( n55144 , n55125 , n55143 );
and ( n55145 , n55122 , n55144 );
or ( n55146 , n55121 , n55145 );
and ( n55147 , n55118 , n55146 );
or ( n55148 , n55117 , n55147 );
and ( n55149 , n55114 , n55148 );
or ( n55150 , n55113 , n55149 );
and ( n55151 , n55110 , n55150 );
or ( n55152 , n55109 , n55151 );
and ( n55153 , n55106 , n55152 );
or ( n55154 , n55105 , n55153 );
and ( n55155 , n55102 , n55154 );
or ( n55156 , n55101 , n55155 );
and ( n55157 , n55098 , n55156 );
or ( n55158 , n55097 , n55157 );
and ( n55159 , n55094 , n55158 );
or ( n55160 , n55093 , n55159 );
and ( n55161 , n55090 , n55160 );
or ( n55162 , n55089 , n55161 );
and ( n55163 , n55086 , n55162 );
or ( n55164 , n55085 , n55163 );
and ( n55165 , n55082 , n55164 );
or ( n55166 , n55081 , n55165 );
and ( n55167 , n55078 , n55166 );
or ( n55168 , n55077 , n55167 );
and ( n55169 , n55074 , n55168 );
or ( n55170 , n55073 , n55169 );
and ( n55171 , n55070 , n55170 );
or ( n55172 , n55069 , n55171 );
and ( n55173 , n55066 , n55172 );
or ( n55174 , n55065 , n55173 );
and ( n55175 , n55062 , n55174 );
or ( n55176 , n55061 , n55175 );
and ( n55177 , n55058 , n55176 );
or ( n55178 , n55057 , n55177 );
and ( n55179 , n55054 , n55178 );
or ( n55180 , n55053 , n55179 );
and ( n55181 , n55050 , n55180 );
or ( n55182 , n55049 , n55181 );
and ( n55183 , n55046 , n55182 );
or ( n55184 , n55045 , n55183 );
and ( n55185 , n55042 , n55184 );
or ( n55186 , n55041 , n55185 );
and ( n55187 , n55038 , n55186 );
or ( n55188 , n55037 , n55187 );
and ( n55189 , n55034 , n55188 );
or ( n55190 , n55033 , n55189 );
and ( n55191 , n55030 , n55190 );
or ( n55192 , n55029 , n55191 );
and ( n55193 , n55026 , n55192 );
or ( n55194 , n55025 , n55193 );
and ( n55195 , n55022 , n55194 );
or ( n55196 , n55021 , n55195 );
and ( n55197 , n55018 , n55196 );
or ( n55198 , n55017 , n55197 );
and ( n55199 , n55014 , n55198 );
or ( n55200 , n55013 , n55199 );
and ( n55201 , n55010 , n55200 );
or ( n55202 , n55009 , n55201 );
and ( n55203 , n55006 , n55202 );
or ( n55204 , n55005 , n55203 );
and ( n55205 , n55002 , n55204 );
or ( n55206 , n55001 , n55205 );
and ( n55207 , n54998 , n55206 );
or ( n55208 , n54997 , n55207 );
and ( n55209 , n54994 , n55208 );
or ( n55210 , n54993 , n55209 );
and ( n55211 , n54990 , n55210 );
or ( n55212 , n54989 , n55211 );
and ( n55213 , n54986 , n55212 );
or ( n55214 , n54985 , n55213 );
and ( n55215 , n54982 , n55214 );
or ( n55216 , n54981 , n55215 );
and ( n55217 , n54978 , n55216 );
or ( n55218 , n54977 , n55217 );
and ( n55219 , n54974 , n55218 );
or ( n55220 , n54973 , n55219 );
and ( n55221 , n54970 , n55220 );
or ( n55222 , n54969 , n55221 );
and ( n55223 , n54966 , n55222 );
or ( n55224 , n54965 , n55223 );
and ( n55225 , n54962 , n55224 );
or ( n55226 , n54961 , n55225 );
and ( n55227 , n54958 , n55226 );
or ( n55228 , n54957 , n55227 );
and ( n55229 , n54954 , n55228 );
or ( n55230 , n54953 , n55229 );
and ( n55231 , n54950 , n55230 );
or ( n55232 , n54949 , n55231 );
and ( n55233 , n54946 , n55232 );
or ( n55234 , n54945 , n55233 );
and ( n55235 , n54942 , n55234 );
or ( n55236 , n54941 , n55235 );
and ( n55237 , n54938 , n55236 );
or ( n55238 , n54937 , n55237 );
and ( n55239 , n54934 , n55238 );
or ( n55240 , n54933 , n55239 );
and ( n55241 , n54930 , n55240 );
or ( n55242 , n54929 , n55241 );
and ( n55243 , n54926 , n55242 );
or ( n55244 , n54925 , n55243 );
and ( n55245 , n54922 , n55244 );
or ( n55246 , n54921 , n55245 );
and ( n55247 , n54918 , n55246 );
or ( n55248 , n54917 , n55247 );
and ( n55249 , n54914 , n55248 );
or ( n55250 , n54913 , n55249 );
and ( n55251 , n54910 , n55250 );
or ( n55252 , n54909 , n55251 );
and ( n55253 , n54906 , n55252 );
or ( n55254 , n54905 , n55253 );
and ( n55255 , n54902 , n55254 );
or ( n55256 , n54901 , n55255 );
and ( n55257 , n54898 , n55256 );
or ( n55258 , n54897 , n55257 );
and ( n55259 , n54894 , n55258 );
or ( n55260 , n54893 , n55259 );
and ( n55261 , n54890 , n55260 );
or ( n55262 , n54889 , n55261 );
and ( n55263 , n54886 , n55262 );
or ( n55264 , n54885 , n55263 );
and ( n55265 , n54882 , n55264 );
or ( n55266 , n54881 , n55265 );
and ( n55267 , n54878 , n55266 );
or ( n55268 , n54877 , n55267 );
and ( n55269 , n54874 , n55268 );
or ( n55270 , n54873 , n55269 );
and ( n55271 , n54870 , n55270 );
or ( n55272 , n54869 , n55271 );
and ( n55273 , n54866 , n55272 );
or ( n55274 , n54865 , n55273 );
and ( n55275 , n54862 , n55274 );
or ( n55276 , n54861 , n55275 );
and ( n55277 , n54858 , n55276 );
or ( n55278 , n54857 , n55277 );
and ( n55279 , n54854 , n55278 );
or ( n55280 , n54853 , n55279 );
and ( n55281 , n54850 , n55280 );
or ( n55282 , n54849 , n55281 );
and ( n55283 , n54846 , n55282 );
or ( n55284 , n54845 , n55283 );
and ( n55285 , n54842 , n55284 );
or ( n55286 , n54841 , n55285 );
and ( n55287 , n54838 , n55286 );
or ( n55288 , n54837 , n55287 );
and ( n55289 , n54834 , n55288 );
or ( n55290 , n54833 , n55289 );
and ( n55291 , n54830 , n55290 );
or ( n55292 , n54829 , n55291 );
and ( n55293 , n54826 , n55292 );
or ( n55294 , n54825 , n55293 );
and ( n55295 , n54822 , n55294 );
or ( n55296 , n54821 , n55295 );
and ( n55297 , n54818 , n55296 );
or ( n55298 , n54817 , n55297 );
and ( n55299 , n54814 , n55298 );
or ( n55300 , n54813 , n55299 );
and ( n55301 , n54810 , n55300 );
or ( n55302 , n54809 , n55301 );
and ( n55303 , n54806 , n55302 );
or ( n55304 , n54805 , n55303 );
and ( n55305 , n54802 , n55304 );
or ( n55306 , n54801 , n55305 );
and ( n55307 , n54798 , n55306 );
or ( n55308 , n54797 , n55307 );
xor ( n55309 , n54794 , n55308 );
buf ( n55310 , n18024 );
and ( n55311 , n29984 , n55310 );
xor ( n55312 , n55309 , n55311 );
xor ( n55313 , n54798 , n55306 );
and ( n55314 , n29989 , n55310 );
and ( n55315 , n55313 , n55314 );
xor ( n55316 , n55313 , n55314 );
xor ( n55317 , n54802 , n55304 );
and ( n55318 , n29994 , n55310 );
and ( n55319 , n55317 , n55318 );
xor ( n55320 , n55317 , n55318 );
xor ( n55321 , n54806 , n55302 );
and ( n55322 , n29999 , n55310 );
and ( n55323 , n55321 , n55322 );
xor ( n55324 , n55321 , n55322 );
xor ( n55325 , n54810 , n55300 );
and ( n55326 , n30004 , n55310 );
and ( n55327 , n55325 , n55326 );
xor ( n55328 , n55325 , n55326 );
xor ( n55329 , n54814 , n55298 );
and ( n55330 , n30009 , n55310 );
and ( n55331 , n55329 , n55330 );
xor ( n55332 , n55329 , n55330 );
xor ( n55333 , n54818 , n55296 );
and ( n55334 , n30014 , n55310 );
and ( n55335 , n55333 , n55334 );
xor ( n55336 , n55333 , n55334 );
xor ( n55337 , n54822 , n55294 );
and ( n55338 , n30019 , n55310 );
and ( n55339 , n55337 , n55338 );
xor ( n55340 , n55337 , n55338 );
xor ( n55341 , n54826 , n55292 );
and ( n55342 , n30024 , n55310 );
and ( n55343 , n55341 , n55342 );
xor ( n55344 , n55341 , n55342 );
xor ( n55345 , n54830 , n55290 );
and ( n55346 , n30029 , n55310 );
and ( n55347 , n55345 , n55346 );
xor ( n55348 , n55345 , n55346 );
xor ( n55349 , n54834 , n55288 );
and ( n55350 , n30034 , n55310 );
and ( n55351 , n55349 , n55350 );
xor ( n55352 , n55349 , n55350 );
xor ( n55353 , n54838 , n55286 );
and ( n55354 , n30039 , n55310 );
and ( n55355 , n55353 , n55354 );
xor ( n55356 , n55353 , n55354 );
xor ( n55357 , n54842 , n55284 );
and ( n55358 , n30044 , n55310 );
and ( n55359 , n55357 , n55358 );
xor ( n55360 , n55357 , n55358 );
xor ( n55361 , n54846 , n55282 );
and ( n55362 , n30049 , n55310 );
and ( n55363 , n55361 , n55362 );
xor ( n55364 , n55361 , n55362 );
xor ( n55365 , n54850 , n55280 );
and ( n55366 , n30054 , n55310 );
and ( n55367 , n55365 , n55366 );
xor ( n55368 , n55365 , n55366 );
xor ( n55369 , n54854 , n55278 );
and ( n55370 , n30059 , n55310 );
and ( n55371 , n55369 , n55370 );
xor ( n55372 , n55369 , n55370 );
xor ( n55373 , n54858 , n55276 );
and ( n55374 , n30064 , n55310 );
and ( n55375 , n55373 , n55374 );
xor ( n55376 , n55373 , n55374 );
xor ( n55377 , n54862 , n55274 );
and ( n55378 , n30069 , n55310 );
and ( n55379 , n55377 , n55378 );
xor ( n55380 , n55377 , n55378 );
xor ( n55381 , n54866 , n55272 );
and ( n55382 , n30074 , n55310 );
and ( n55383 , n55381 , n55382 );
xor ( n55384 , n55381 , n55382 );
xor ( n55385 , n54870 , n55270 );
and ( n55386 , n30079 , n55310 );
and ( n55387 , n55385 , n55386 );
xor ( n55388 , n55385 , n55386 );
xor ( n55389 , n54874 , n55268 );
and ( n55390 , n30084 , n55310 );
and ( n55391 , n55389 , n55390 );
xor ( n55392 , n55389 , n55390 );
xor ( n55393 , n54878 , n55266 );
and ( n55394 , n30089 , n55310 );
and ( n55395 , n55393 , n55394 );
xor ( n55396 , n55393 , n55394 );
xor ( n55397 , n54882 , n55264 );
and ( n55398 , n30094 , n55310 );
and ( n55399 , n55397 , n55398 );
xor ( n55400 , n55397 , n55398 );
xor ( n55401 , n54886 , n55262 );
and ( n55402 , n30099 , n55310 );
and ( n55403 , n55401 , n55402 );
xor ( n55404 , n55401 , n55402 );
xor ( n55405 , n54890 , n55260 );
and ( n55406 , n30104 , n55310 );
and ( n55407 , n55405 , n55406 );
xor ( n55408 , n55405 , n55406 );
xor ( n55409 , n54894 , n55258 );
and ( n55410 , n30109 , n55310 );
and ( n55411 , n55409 , n55410 );
xor ( n55412 , n55409 , n55410 );
xor ( n55413 , n54898 , n55256 );
and ( n55414 , n30114 , n55310 );
and ( n55415 , n55413 , n55414 );
xor ( n55416 , n55413 , n55414 );
xor ( n55417 , n54902 , n55254 );
and ( n55418 , n30119 , n55310 );
and ( n55419 , n55417 , n55418 );
xor ( n55420 , n55417 , n55418 );
xor ( n55421 , n54906 , n55252 );
and ( n55422 , n30124 , n55310 );
and ( n55423 , n55421 , n55422 );
xor ( n55424 , n55421 , n55422 );
xor ( n55425 , n54910 , n55250 );
and ( n55426 , n30129 , n55310 );
and ( n55427 , n55425 , n55426 );
xor ( n55428 , n55425 , n55426 );
xor ( n55429 , n54914 , n55248 );
and ( n55430 , n30134 , n55310 );
and ( n55431 , n55429 , n55430 );
xor ( n55432 , n55429 , n55430 );
xor ( n55433 , n54918 , n55246 );
and ( n55434 , n30139 , n55310 );
and ( n55435 , n55433 , n55434 );
xor ( n55436 , n55433 , n55434 );
xor ( n55437 , n54922 , n55244 );
and ( n55438 , n30144 , n55310 );
and ( n55439 , n55437 , n55438 );
xor ( n55440 , n55437 , n55438 );
xor ( n55441 , n54926 , n55242 );
and ( n55442 , n30149 , n55310 );
and ( n55443 , n55441 , n55442 );
xor ( n55444 , n55441 , n55442 );
xor ( n55445 , n54930 , n55240 );
and ( n55446 , n30154 , n55310 );
and ( n55447 , n55445 , n55446 );
xor ( n55448 , n55445 , n55446 );
xor ( n55449 , n54934 , n55238 );
and ( n55450 , n30159 , n55310 );
and ( n55451 , n55449 , n55450 );
xor ( n55452 , n55449 , n55450 );
xor ( n55453 , n54938 , n55236 );
and ( n55454 , n30164 , n55310 );
and ( n55455 , n55453 , n55454 );
xor ( n55456 , n55453 , n55454 );
xor ( n55457 , n54942 , n55234 );
and ( n55458 , n30169 , n55310 );
and ( n55459 , n55457 , n55458 );
xor ( n55460 , n55457 , n55458 );
xor ( n55461 , n54946 , n55232 );
and ( n55462 , n30174 , n55310 );
and ( n55463 , n55461 , n55462 );
xor ( n55464 , n55461 , n55462 );
xor ( n55465 , n54950 , n55230 );
and ( n55466 , n30179 , n55310 );
and ( n55467 , n55465 , n55466 );
xor ( n55468 , n55465 , n55466 );
xor ( n55469 , n54954 , n55228 );
and ( n55470 , n30184 , n55310 );
and ( n55471 , n55469 , n55470 );
xor ( n55472 , n55469 , n55470 );
xor ( n55473 , n54958 , n55226 );
and ( n55474 , n30189 , n55310 );
and ( n55475 , n55473 , n55474 );
xor ( n55476 , n55473 , n55474 );
xor ( n55477 , n54962 , n55224 );
and ( n55478 , n30194 , n55310 );
and ( n55479 , n55477 , n55478 );
xor ( n55480 , n55477 , n55478 );
xor ( n55481 , n54966 , n55222 );
and ( n55482 , n30199 , n55310 );
and ( n55483 , n55481 , n55482 );
xor ( n55484 , n55481 , n55482 );
xor ( n55485 , n54970 , n55220 );
and ( n55486 , n30204 , n55310 );
and ( n55487 , n55485 , n55486 );
xor ( n55488 , n55485 , n55486 );
xor ( n55489 , n54974 , n55218 );
and ( n55490 , n30209 , n55310 );
and ( n55491 , n55489 , n55490 );
xor ( n55492 , n55489 , n55490 );
xor ( n55493 , n54978 , n55216 );
and ( n55494 , n30214 , n55310 );
and ( n55495 , n55493 , n55494 );
xor ( n55496 , n55493 , n55494 );
xor ( n55497 , n54982 , n55214 );
and ( n55498 , n30219 , n55310 );
and ( n55499 , n55497 , n55498 );
xor ( n55500 , n55497 , n55498 );
xor ( n55501 , n54986 , n55212 );
and ( n55502 , n30224 , n55310 );
and ( n55503 , n55501 , n55502 );
xor ( n55504 , n55501 , n55502 );
xor ( n55505 , n54990 , n55210 );
and ( n55506 , n30229 , n55310 );
and ( n55507 , n55505 , n55506 );
xor ( n55508 , n55505 , n55506 );
xor ( n55509 , n54994 , n55208 );
and ( n55510 , n30234 , n55310 );
and ( n55511 , n55509 , n55510 );
xor ( n55512 , n55509 , n55510 );
xor ( n55513 , n54998 , n55206 );
and ( n55514 , n30239 , n55310 );
and ( n55515 , n55513 , n55514 );
xor ( n55516 , n55513 , n55514 );
xor ( n55517 , n55002 , n55204 );
and ( n55518 , n30244 , n55310 );
and ( n55519 , n55517 , n55518 );
xor ( n55520 , n55517 , n55518 );
xor ( n55521 , n55006 , n55202 );
and ( n55522 , n30249 , n55310 );
and ( n55523 , n55521 , n55522 );
xor ( n55524 , n55521 , n55522 );
xor ( n55525 , n55010 , n55200 );
and ( n55526 , n30254 , n55310 );
and ( n55527 , n55525 , n55526 );
xor ( n55528 , n55525 , n55526 );
xor ( n55529 , n55014 , n55198 );
and ( n55530 , n30259 , n55310 );
and ( n55531 , n55529 , n55530 );
xor ( n55532 , n55529 , n55530 );
xor ( n55533 , n55018 , n55196 );
and ( n55534 , n30264 , n55310 );
and ( n55535 , n55533 , n55534 );
xor ( n55536 , n55533 , n55534 );
xor ( n55537 , n55022 , n55194 );
and ( n55538 , n30269 , n55310 );
and ( n55539 , n55537 , n55538 );
xor ( n55540 , n55537 , n55538 );
xor ( n55541 , n55026 , n55192 );
and ( n55542 , n30274 , n55310 );
and ( n55543 , n55541 , n55542 );
xor ( n55544 , n55541 , n55542 );
xor ( n55545 , n55030 , n55190 );
and ( n55546 , n30279 , n55310 );
and ( n55547 , n55545 , n55546 );
xor ( n55548 , n55545 , n55546 );
xor ( n55549 , n55034 , n55188 );
and ( n55550 , n30284 , n55310 );
and ( n55551 , n55549 , n55550 );
xor ( n55552 , n55549 , n55550 );
xor ( n55553 , n55038 , n55186 );
and ( n55554 , n30289 , n55310 );
and ( n55555 , n55553 , n55554 );
xor ( n55556 , n55553 , n55554 );
xor ( n55557 , n55042 , n55184 );
and ( n55558 , n30294 , n55310 );
and ( n55559 , n55557 , n55558 );
xor ( n55560 , n55557 , n55558 );
xor ( n55561 , n55046 , n55182 );
and ( n55562 , n30299 , n55310 );
and ( n55563 , n55561 , n55562 );
xor ( n55564 , n55561 , n55562 );
xor ( n55565 , n55050 , n55180 );
and ( n55566 , n30304 , n55310 );
and ( n55567 , n55565 , n55566 );
xor ( n55568 , n55565 , n55566 );
xor ( n55569 , n55054 , n55178 );
and ( n55570 , n30309 , n55310 );
and ( n55571 , n55569 , n55570 );
xor ( n55572 , n55569 , n55570 );
xor ( n55573 , n55058 , n55176 );
and ( n55574 , n30314 , n55310 );
and ( n55575 , n55573 , n55574 );
xor ( n55576 , n55573 , n55574 );
xor ( n55577 , n55062 , n55174 );
and ( n55578 , n30319 , n55310 );
and ( n55579 , n55577 , n55578 );
xor ( n55580 , n55577 , n55578 );
xor ( n55581 , n55066 , n55172 );
and ( n55582 , n30324 , n55310 );
and ( n55583 , n55581 , n55582 );
xor ( n55584 , n55581 , n55582 );
xor ( n55585 , n55070 , n55170 );
and ( n55586 , n30329 , n55310 );
and ( n55587 , n55585 , n55586 );
xor ( n55588 , n55585 , n55586 );
xor ( n55589 , n55074 , n55168 );
and ( n55590 , n30334 , n55310 );
and ( n55591 , n55589 , n55590 );
xor ( n55592 , n55589 , n55590 );
xor ( n55593 , n55078 , n55166 );
and ( n55594 , n30339 , n55310 );
and ( n55595 , n55593 , n55594 );
xor ( n55596 , n55593 , n55594 );
xor ( n55597 , n55082 , n55164 );
and ( n55598 , n30344 , n55310 );
and ( n55599 , n55597 , n55598 );
xor ( n55600 , n55597 , n55598 );
xor ( n55601 , n55086 , n55162 );
and ( n55602 , n30349 , n55310 );
and ( n55603 , n55601 , n55602 );
xor ( n55604 , n55601 , n55602 );
xor ( n55605 , n55090 , n55160 );
and ( n55606 , n30354 , n55310 );
and ( n55607 , n55605 , n55606 );
xor ( n55608 , n55605 , n55606 );
xor ( n55609 , n55094 , n55158 );
and ( n55610 , n30359 , n55310 );
and ( n55611 , n55609 , n55610 );
xor ( n55612 , n55609 , n55610 );
xor ( n55613 , n55098 , n55156 );
and ( n55614 , n30364 , n55310 );
and ( n55615 , n55613 , n55614 );
xor ( n55616 , n55613 , n55614 );
xor ( n55617 , n55102 , n55154 );
and ( n55618 , n30369 , n55310 );
and ( n55619 , n55617 , n55618 );
xor ( n55620 , n55617 , n55618 );
xor ( n55621 , n55106 , n55152 );
and ( n55622 , n30374 , n55310 );
and ( n55623 , n55621 , n55622 );
xor ( n55624 , n55621 , n55622 );
xor ( n55625 , n55110 , n55150 );
and ( n55626 , n30379 , n55310 );
and ( n55627 , n55625 , n55626 );
xor ( n55628 , n55625 , n55626 );
xor ( n55629 , n55114 , n55148 );
and ( n55630 , n30384 , n55310 );
and ( n55631 , n55629 , n55630 );
xor ( n55632 , n55629 , n55630 );
xor ( n55633 , n55118 , n55146 );
and ( n55634 , n30389 , n55310 );
and ( n55635 , n55633 , n55634 );
xor ( n55636 , n55633 , n55634 );
xor ( n55637 , n55122 , n55144 );
and ( n55638 , n30394 , n55310 );
and ( n55639 , n55637 , n55638 );
xor ( n55640 , n55637 , n55638 );
xor ( n55641 , n55126 , n55142 );
and ( n55642 , n30399 , n55310 );
and ( n55643 , n55641 , n55642 );
xor ( n55644 , n55641 , n55642 );
xor ( n55645 , n55130 , n55140 );
and ( n55646 , n30404 , n55310 );
and ( n55647 , n55645 , n55646 );
xor ( n55648 , n55645 , n55646 );
xor ( n55649 , n55134 , n55138 );
and ( n55650 , n30409 , n55310 );
and ( n55651 , n55649 , n55650 );
buf ( n55652 , n55651 );
and ( n55653 , n55648 , n55652 );
or ( n55654 , n55647 , n55653 );
and ( n55655 , n55644 , n55654 );
or ( n55656 , n55643 , n55655 );
and ( n55657 , n55640 , n55656 );
or ( n55658 , n55639 , n55657 );
and ( n55659 , n55636 , n55658 );
or ( n55660 , n55635 , n55659 );
and ( n55661 , n55632 , n55660 );
or ( n55662 , n55631 , n55661 );
and ( n55663 , n55628 , n55662 );
or ( n55664 , n55627 , n55663 );
and ( n55665 , n55624 , n55664 );
or ( n55666 , n55623 , n55665 );
and ( n55667 , n55620 , n55666 );
or ( n55668 , n55619 , n55667 );
and ( n55669 , n55616 , n55668 );
or ( n55670 , n55615 , n55669 );
and ( n55671 , n55612 , n55670 );
or ( n55672 , n55611 , n55671 );
and ( n55673 , n55608 , n55672 );
or ( n55674 , n55607 , n55673 );
and ( n55675 , n55604 , n55674 );
or ( n55676 , n55603 , n55675 );
and ( n55677 , n55600 , n55676 );
or ( n55678 , n55599 , n55677 );
and ( n55679 , n55596 , n55678 );
or ( n55680 , n55595 , n55679 );
and ( n55681 , n55592 , n55680 );
or ( n55682 , n55591 , n55681 );
and ( n55683 , n55588 , n55682 );
or ( n55684 , n55587 , n55683 );
and ( n55685 , n55584 , n55684 );
or ( n55686 , n55583 , n55685 );
and ( n55687 , n55580 , n55686 );
or ( n55688 , n55579 , n55687 );
and ( n55689 , n55576 , n55688 );
or ( n55690 , n55575 , n55689 );
and ( n55691 , n55572 , n55690 );
or ( n55692 , n55571 , n55691 );
and ( n55693 , n55568 , n55692 );
or ( n55694 , n55567 , n55693 );
and ( n55695 , n55564 , n55694 );
or ( n55696 , n55563 , n55695 );
and ( n55697 , n55560 , n55696 );
or ( n55698 , n55559 , n55697 );
and ( n55699 , n55556 , n55698 );
or ( n55700 , n55555 , n55699 );
and ( n55701 , n55552 , n55700 );
or ( n55702 , n55551 , n55701 );
and ( n55703 , n55548 , n55702 );
or ( n55704 , n55547 , n55703 );
and ( n55705 , n55544 , n55704 );
or ( n55706 , n55543 , n55705 );
and ( n55707 , n55540 , n55706 );
or ( n55708 , n55539 , n55707 );
and ( n55709 , n55536 , n55708 );
or ( n55710 , n55535 , n55709 );
and ( n55711 , n55532 , n55710 );
or ( n55712 , n55531 , n55711 );
and ( n55713 , n55528 , n55712 );
or ( n55714 , n55527 , n55713 );
and ( n55715 , n55524 , n55714 );
or ( n55716 , n55523 , n55715 );
and ( n55717 , n55520 , n55716 );
or ( n55718 , n55519 , n55717 );
and ( n55719 , n55516 , n55718 );
or ( n55720 , n55515 , n55719 );
and ( n55721 , n55512 , n55720 );
or ( n55722 , n55511 , n55721 );
and ( n55723 , n55508 , n55722 );
or ( n55724 , n55507 , n55723 );
and ( n55725 , n55504 , n55724 );
or ( n55726 , n55503 , n55725 );
and ( n55727 , n55500 , n55726 );
or ( n55728 , n55499 , n55727 );
and ( n55729 , n55496 , n55728 );
or ( n55730 , n55495 , n55729 );
and ( n55731 , n55492 , n55730 );
or ( n55732 , n55491 , n55731 );
and ( n55733 , n55488 , n55732 );
or ( n55734 , n55487 , n55733 );
and ( n55735 , n55484 , n55734 );
or ( n55736 , n55483 , n55735 );
and ( n55737 , n55480 , n55736 );
or ( n55738 , n55479 , n55737 );
and ( n55739 , n55476 , n55738 );
or ( n55740 , n55475 , n55739 );
and ( n55741 , n55472 , n55740 );
or ( n55742 , n55471 , n55741 );
and ( n55743 , n55468 , n55742 );
or ( n55744 , n55467 , n55743 );
and ( n55745 , n55464 , n55744 );
or ( n55746 , n55463 , n55745 );
and ( n55747 , n55460 , n55746 );
or ( n55748 , n55459 , n55747 );
and ( n55749 , n55456 , n55748 );
or ( n55750 , n55455 , n55749 );
and ( n55751 , n55452 , n55750 );
or ( n55752 , n55451 , n55751 );
and ( n55753 , n55448 , n55752 );
or ( n55754 , n55447 , n55753 );
and ( n55755 , n55444 , n55754 );
or ( n55756 , n55443 , n55755 );
and ( n55757 , n55440 , n55756 );
or ( n55758 , n55439 , n55757 );
and ( n55759 , n55436 , n55758 );
or ( n55760 , n55435 , n55759 );
and ( n55761 , n55432 , n55760 );
or ( n55762 , n55431 , n55761 );
and ( n55763 , n55428 , n55762 );
or ( n55764 , n55427 , n55763 );
and ( n55765 , n55424 , n55764 );
or ( n55766 , n55423 , n55765 );
and ( n55767 , n55420 , n55766 );
or ( n55768 , n55419 , n55767 );
and ( n55769 , n55416 , n55768 );
or ( n55770 , n55415 , n55769 );
and ( n55771 , n55412 , n55770 );
or ( n55772 , n55411 , n55771 );
and ( n55773 , n55408 , n55772 );
or ( n55774 , n55407 , n55773 );
and ( n55775 , n55404 , n55774 );
or ( n55776 , n55403 , n55775 );
and ( n55777 , n55400 , n55776 );
or ( n55778 , n55399 , n55777 );
and ( n55779 , n55396 , n55778 );
or ( n55780 , n55395 , n55779 );
and ( n55781 , n55392 , n55780 );
or ( n55782 , n55391 , n55781 );
and ( n55783 , n55388 , n55782 );
or ( n55784 , n55387 , n55783 );
and ( n55785 , n55384 , n55784 );
or ( n55786 , n55383 , n55785 );
and ( n55787 , n55380 , n55786 );
or ( n55788 , n55379 , n55787 );
and ( n55789 , n55376 , n55788 );
or ( n55790 , n55375 , n55789 );
and ( n55791 , n55372 , n55790 );
or ( n55792 , n55371 , n55791 );
and ( n55793 , n55368 , n55792 );
or ( n55794 , n55367 , n55793 );
and ( n55795 , n55364 , n55794 );
or ( n55796 , n55363 , n55795 );
and ( n55797 , n55360 , n55796 );
or ( n55798 , n55359 , n55797 );
and ( n55799 , n55356 , n55798 );
or ( n55800 , n55355 , n55799 );
and ( n55801 , n55352 , n55800 );
or ( n55802 , n55351 , n55801 );
and ( n55803 , n55348 , n55802 );
or ( n55804 , n55347 , n55803 );
and ( n55805 , n55344 , n55804 );
or ( n55806 , n55343 , n55805 );
and ( n55807 , n55340 , n55806 );
or ( n55808 , n55339 , n55807 );
and ( n55809 , n55336 , n55808 );
or ( n55810 , n55335 , n55809 );
and ( n55811 , n55332 , n55810 );
or ( n55812 , n55331 , n55811 );
and ( n55813 , n55328 , n55812 );
or ( n55814 , n55327 , n55813 );
and ( n55815 , n55324 , n55814 );
or ( n55816 , n55323 , n55815 );
and ( n55817 , n55320 , n55816 );
or ( n55818 , n55319 , n55817 );
and ( n55819 , n55316 , n55818 );
or ( n55820 , n55315 , n55819 );
xor ( n55821 , n55312 , n55820 );
buf ( n55822 , n18022 );
and ( n55823 , n29989 , n55822 );
xor ( n55824 , n55821 , n55823 );
xor ( n55825 , n55316 , n55818 );
and ( n55826 , n29994 , n55822 );
and ( n55827 , n55825 , n55826 );
xor ( n55828 , n55825 , n55826 );
xor ( n55829 , n55320 , n55816 );
and ( n55830 , n29999 , n55822 );
and ( n55831 , n55829 , n55830 );
xor ( n55832 , n55829 , n55830 );
xor ( n55833 , n55324 , n55814 );
and ( n55834 , n30004 , n55822 );
and ( n55835 , n55833 , n55834 );
xor ( n55836 , n55833 , n55834 );
xor ( n55837 , n55328 , n55812 );
and ( n55838 , n30009 , n55822 );
and ( n55839 , n55837 , n55838 );
xor ( n55840 , n55837 , n55838 );
xor ( n55841 , n55332 , n55810 );
and ( n55842 , n30014 , n55822 );
and ( n55843 , n55841 , n55842 );
xor ( n55844 , n55841 , n55842 );
xor ( n55845 , n55336 , n55808 );
and ( n55846 , n30019 , n55822 );
and ( n55847 , n55845 , n55846 );
xor ( n55848 , n55845 , n55846 );
xor ( n55849 , n55340 , n55806 );
and ( n55850 , n30024 , n55822 );
and ( n55851 , n55849 , n55850 );
xor ( n55852 , n55849 , n55850 );
xor ( n55853 , n55344 , n55804 );
and ( n55854 , n30029 , n55822 );
and ( n55855 , n55853 , n55854 );
xor ( n55856 , n55853 , n55854 );
xor ( n55857 , n55348 , n55802 );
and ( n55858 , n30034 , n55822 );
and ( n55859 , n55857 , n55858 );
xor ( n55860 , n55857 , n55858 );
xor ( n55861 , n55352 , n55800 );
and ( n55862 , n30039 , n55822 );
and ( n55863 , n55861 , n55862 );
xor ( n55864 , n55861 , n55862 );
xor ( n55865 , n55356 , n55798 );
and ( n55866 , n30044 , n55822 );
and ( n55867 , n55865 , n55866 );
xor ( n55868 , n55865 , n55866 );
xor ( n55869 , n55360 , n55796 );
and ( n55870 , n30049 , n55822 );
and ( n55871 , n55869 , n55870 );
xor ( n55872 , n55869 , n55870 );
xor ( n55873 , n55364 , n55794 );
and ( n55874 , n30054 , n55822 );
and ( n55875 , n55873 , n55874 );
xor ( n55876 , n55873 , n55874 );
xor ( n55877 , n55368 , n55792 );
and ( n55878 , n30059 , n55822 );
and ( n55879 , n55877 , n55878 );
xor ( n55880 , n55877 , n55878 );
xor ( n55881 , n55372 , n55790 );
and ( n55882 , n30064 , n55822 );
and ( n55883 , n55881 , n55882 );
xor ( n55884 , n55881 , n55882 );
xor ( n55885 , n55376 , n55788 );
and ( n55886 , n30069 , n55822 );
and ( n55887 , n55885 , n55886 );
xor ( n55888 , n55885 , n55886 );
xor ( n55889 , n55380 , n55786 );
and ( n55890 , n30074 , n55822 );
and ( n55891 , n55889 , n55890 );
xor ( n55892 , n55889 , n55890 );
xor ( n55893 , n55384 , n55784 );
and ( n55894 , n30079 , n55822 );
and ( n55895 , n55893 , n55894 );
xor ( n55896 , n55893 , n55894 );
xor ( n55897 , n55388 , n55782 );
and ( n55898 , n30084 , n55822 );
and ( n55899 , n55897 , n55898 );
xor ( n55900 , n55897 , n55898 );
xor ( n55901 , n55392 , n55780 );
and ( n55902 , n30089 , n55822 );
and ( n55903 , n55901 , n55902 );
xor ( n55904 , n55901 , n55902 );
xor ( n55905 , n55396 , n55778 );
and ( n55906 , n30094 , n55822 );
and ( n55907 , n55905 , n55906 );
xor ( n55908 , n55905 , n55906 );
xor ( n55909 , n55400 , n55776 );
and ( n55910 , n30099 , n55822 );
and ( n55911 , n55909 , n55910 );
xor ( n55912 , n55909 , n55910 );
xor ( n55913 , n55404 , n55774 );
and ( n55914 , n30104 , n55822 );
and ( n55915 , n55913 , n55914 );
xor ( n55916 , n55913 , n55914 );
xor ( n55917 , n55408 , n55772 );
and ( n55918 , n30109 , n55822 );
and ( n55919 , n55917 , n55918 );
xor ( n55920 , n55917 , n55918 );
xor ( n55921 , n55412 , n55770 );
and ( n55922 , n30114 , n55822 );
and ( n55923 , n55921 , n55922 );
xor ( n55924 , n55921 , n55922 );
xor ( n55925 , n55416 , n55768 );
and ( n55926 , n30119 , n55822 );
and ( n55927 , n55925 , n55926 );
xor ( n55928 , n55925 , n55926 );
xor ( n55929 , n55420 , n55766 );
and ( n55930 , n30124 , n55822 );
and ( n55931 , n55929 , n55930 );
xor ( n55932 , n55929 , n55930 );
xor ( n55933 , n55424 , n55764 );
and ( n55934 , n30129 , n55822 );
and ( n55935 , n55933 , n55934 );
xor ( n55936 , n55933 , n55934 );
xor ( n55937 , n55428 , n55762 );
and ( n55938 , n30134 , n55822 );
and ( n55939 , n55937 , n55938 );
xor ( n55940 , n55937 , n55938 );
xor ( n55941 , n55432 , n55760 );
and ( n55942 , n30139 , n55822 );
and ( n55943 , n55941 , n55942 );
xor ( n55944 , n55941 , n55942 );
xor ( n55945 , n55436 , n55758 );
and ( n55946 , n30144 , n55822 );
and ( n55947 , n55945 , n55946 );
xor ( n55948 , n55945 , n55946 );
xor ( n55949 , n55440 , n55756 );
and ( n55950 , n30149 , n55822 );
and ( n55951 , n55949 , n55950 );
xor ( n55952 , n55949 , n55950 );
xor ( n55953 , n55444 , n55754 );
and ( n55954 , n30154 , n55822 );
and ( n55955 , n55953 , n55954 );
xor ( n55956 , n55953 , n55954 );
xor ( n55957 , n55448 , n55752 );
and ( n55958 , n30159 , n55822 );
and ( n55959 , n55957 , n55958 );
xor ( n55960 , n55957 , n55958 );
xor ( n55961 , n55452 , n55750 );
and ( n55962 , n30164 , n55822 );
and ( n55963 , n55961 , n55962 );
xor ( n55964 , n55961 , n55962 );
xor ( n55965 , n55456 , n55748 );
and ( n55966 , n30169 , n55822 );
and ( n55967 , n55965 , n55966 );
xor ( n55968 , n55965 , n55966 );
xor ( n55969 , n55460 , n55746 );
and ( n55970 , n30174 , n55822 );
and ( n55971 , n55969 , n55970 );
xor ( n55972 , n55969 , n55970 );
xor ( n55973 , n55464 , n55744 );
and ( n55974 , n30179 , n55822 );
and ( n55975 , n55973 , n55974 );
xor ( n55976 , n55973 , n55974 );
xor ( n55977 , n55468 , n55742 );
and ( n55978 , n30184 , n55822 );
and ( n55979 , n55977 , n55978 );
xor ( n55980 , n55977 , n55978 );
xor ( n55981 , n55472 , n55740 );
and ( n55982 , n30189 , n55822 );
and ( n55983 , n55981 , n55982 );
xor ( n55984 , n55981 , n55982 );
xor ( n55985 , n55476 , n55738 );
and ( n55986 , n30194 , n55822 );
and ( n55987 , n55985 , n55986 );
xor ( n55988 , n55985 , n55986 );
xor ( n55989 , n55480 , n55736 );
and ( n55990 , n30199 , n55822 );
and ( n55991 , n55989 , n55990 );
xor ( n55992 , n55989 , n55990 );
xor ( n55993 , n55484 , n55734 );
and ( n55994 , n30204 , n55822 );
and ( n55995 , n55993 , n55994 );
xor ( n55996 , n55993 , n55994 );
xor ( n55997 , n55488 , n55732 );
and ( n55998 , n30209 , n55822 );
and ( n55999 , n55997 , n55998 );
xor ( n56000 , n55997 , n55998 );
xor ( n56001 , n55492 , n55730 );
and ( n56002 , n30214 , n55822 );
and ( n56003 , n56001 , n56002 );
xor ( n56004 , n56001 , n56002 );
xor ( n56005 , n55496 , n55728 );
and ( n56006 , n30219 , n55822 );
and ( n56007 , n56005 , n56006 );
xor ( n56008 , n56005 , n56006 );
xor ( n56009 , n55500 , n55726 );
and ( n56010 , n30224 , n55822 );
and ( n56011 , n56009 , n56010 );
xor ( n56012 , n56009 , n56010 );
xor ( n56013 , n55504 , n55724 );
and ( n56014 , n30229 , n55822 );
and ( n56015 , n56013 , n56014 );
xor ( n56016 , n56013 , n56014 );
xor ( n56017 , n55508 , n55722 );
and ( n56018 , n30234 , n55822 );
and ( n56019 , n56017 , n56018 );
xor ( n56020 , n56017 , n56018 );
xor ( n56021 , n55512 , n55720 );
and ( n56022 , n30239 , n55822 );
and ( n56023 , n56021 , n56022 );
xor ( n56024 , n56021 , n56022 );
xor ( n56025 , n55516 , n55718 );
and ( n56026 , n30244 , n55822 );
and ( n56027 , n56025 , n56026 );
xor ( n56028 , n56025 , n56026 );
xor ( n56029 , n55520 , n55716 );
and ( n56030 , n30249 , n55822 );
and ( n56031 , n56029 , n56030 );
xor ( n56032 , n56029 , n56030 );
xor ( n56033 , n55524 , n55714 );
and ( n56034 , n30254 , n55822 );
and ( n56035 , n56033 , n56034 );
xor ( n56036 , n56033 , n56034 );
xor ( n56037 , n55528 , n55712 );
and ( n56038 , n30259 , n55822 );
and ( n56039 , n56037 , n56038 );
xor ( n56040 , n56037 , n56038 );
xor ( n56041 , n55532 , n55710 );
and ( n56042 , n30264 , n55822 );
and ( n56043 , n56041 , n56042 );
xor ( n56044 , n56041 , n56042 );
xor ( n56045 , n55536 , n55708 );
and ( n56046 , n30269 , n55822 );
and ( n56047 , n56045 , n56046 );
xor ( n56048 , n56045 , n56046 );
xor ( n56049 , n55540 , n55706 );
and ( n56050 , n30274 , n55822 );
and ( n56051 , n56049 , n56050 );
xor ( n56052 , n56049 , n56050 );
xor ( n56053 , n55544 , n55704 );
and ( n56054 , n30279 , n55822 );
and ( n56055 , n56053 , n56054 );
xor ( n56056 , n56053 , n56054 );
xor ( n56057 , n55548 , n55702 );
and ( n56058 , n30284 , n55822 );
and ( n56059 , n56057 , n56058 );
xor ( n56060 , n56057 , n56058 );
xor ( n56061 , n55552 , n55700 );
and ( n56062 , n30289 , n55822 );
and ( n56063 , n56061 , n56062 );
xor ( n56064 , n56061 , n56062 );
xor ( n56065 , n55556 , n55698 );
and ( n56066 , n30294 , n55822 );
and ( n56067 , n56065 , n56066 );
xor ( n56068 , n56065 , n56066 );
xor ( n56069 , n55560 , n55696 );
and ( n56070 , n30299 , n55822 );
and ( n56071 , n56069 , n56070 );
xor ( n56072 , n56069 , n56070 );
xor ( n56073 , n55564 , n55694 );
and ( n56074 , n30304 , n55822 );
and ( n56075 , n56073 , n56074 );
xor ( n56076 , n56073 , n56074 );
xor ( n56077 , n55568 , n55692 );
and ( n56078 , n30309 , n55822 );
and ( n56079 , n56077 , n56078 );
xor ( n56080 , n56077 , n56078 );
xor ( n56081 , n55572 , n55690 );
and ( n56082 , n30314 , n55822 );
and ( n56083 , n56081 , n56082 );
xor ( n56084 , n56081 , n56082 );
xor ( n56085 , n55576 , n55688 );
and ( n56086 , n30319 , n55822 );
and ( n56087 , n56085 , n56086 );
xor ( n56088 , n56085 , n56086 );
xor ( n56089 , n55580 , n55686 );
and ( n56090 , n30324 , n55822 );
and ( n56091 , n56089 , n56090 );
xor ( n56092 , n56089 , n56090 );
xor ( n56093 , n55584 , n55684 );
and ( n56094 , n30329 , n55822 );
and ( n56095 , n56093 , n56094 );
xor ( n56096 , n56093 , n56094 );
xor ( n56097 , n55588 , n55682 );
and ( n56098 , n30334 , n55822 );
and ( n56099 , n56097 , n56098 );
xor ( n56100 , n56097 , n56098 );
xor ( n56101 , n55592 , n55680 );
and ( n56102 , n30339 , n55822 );
and ( n56103 , n56101 , n56102 );
xor ( n56104 , n56101 , n56102 );
xor ( n56105 , n55596 , n55678 );
and ( n56106 , n30344 , n55822 );
and ( n56107 , n56105 , n56106 );
xor ( n56108 , n56105 , n56106 );
xor ( n56109 , n55600 , n55676 );
and ( n56110 , n30349 , n55822 );
and ( n56111 , n56109 , n56110 );
xor ( n56112 , n56109 , n56110 );
xor ( n56113 , n55604 , n55674 );
and ( n56114 , n30354 , n55822 );
and ( n56115 , n56113 , n56114 );
xor ( n56116 , n56113 , n56114 );
xor ( n56117 , n55608 , n55672 );
and ( n56118 , n30359 , n55822 );
and ( n56119 , n56117 , n56118 );
xor ( n56120 , n56117 , n56118 );
xor ( n56121 , n55612 , n55670 );
and ( n56122 , n30364 , n55822 );
and ( n56123 , n56121 , n56122 );
xor ( n56124 , n56121 , n56122 );
xor ( n56125 , n55616 , n55668 );
and ( n56126 , n30369 , n55822 );
and ( n56127 , n56125 , n56126 );
xor ( n56128 , n56125 , n56126 );
xor ( n56129 , n55620 , n55666 );
and ( n56130 , n30374 , n55822 );
and ( n56131 , n56129 , n56130 );
xor ( n56132 , n56129 , n56130 );
xor ( n56133 , n55624 , n55664 );
and ( n56134 , n30379 , n55822 );
and ( n56135 , n56133 , n56134 );
xor ( n56136 , n56133 , n56134 );
xor ( n56137 , n55628 , n55662 );
and ( n56138 , n30384 , n55822 );
and ( n56139 , n56137 , n56138 );
xor ( n56140 , n56137 , n56138 );
xor ( n56141 , n55632 , n55660 );
and ( n56142 , n30389 , n55822 );
and ( n56143 , n56141 , n56142 );
xor ( n56144 , n56141 , n56142 );
xor ( n56145 , n55636 , n55658 );
and ( n56146 , n30394 , n55822 );
and ( n56147 , n56145 , n56146 );
xor ( n56148 , n56145 , n56146 );
xor ( n56149 , n55640 , n55656 );
and ( n56150 , n30399 , n55822 );
and ( n56151 , n56149 , n56150 );
xor ( n56152 , n56149 , n56150 );
xor ( n56153 , n55644 , n55654 );
and ( n56154 , n30404 , n55822 );
and ( n56155 , n56153 , n56154 );
xor ( n56156 , n56153 , n56154 );
xor ( n56157 , n55648 , n55652 );
and ( n56158 , n30409 , n55822 );
and ( n56159 , n56157 , n56158 );
buf ( n56160 , n56159 );
and ( n56161 , n56156 , n56160 );
or ( n56162 , n56155 , n56161 );
and ( n56163 , n56152 , n56162 );
or ( n56164 , n56151 , n56163 );
and ( n56165 , n56148 , n56164 );
or ( n56166 , n56147 , n56165 );
and ( n56167 , n56144 , n56166 );
or ( n56168 , n56143 , n56167 );
and ( n56169 , n56140 , n56168 );
or ( n56170 , n56139 , n56169 );
and ( n56171 , n56136 , n56170 );
or ( n56172 , n56135 , n56171 );
and ( n56173 , n56132 , n56172 );
or ( n56174 , n56131 , n56173 );
and ( n56175 , n56128 , n56174 );
or ( n56176 , n56127 , n56175 );
and ( n56177 , n56124 , n56176 );
or ( n56178 , n56123 , n56177 );
and ( n56179 , n56120 , n56178 );
or ( n56180 , n56119 , n56179 );
and ( n56181 , n56116 , n56180 );
or ( n56182 , n56115 , n56181 );
and ( n56183 , n56112 , n56182 );
or ( n56184 , n56111 , n56183 );
and ( n56185 , n56108 , n56184 );
or ( n56186 , n56107 , n56185 );
and ( n56187 , n56104 , n56186 );
or ( n56188 , n56103 , n56187 );
and ( n56189 , n56100 , n56188 );
or ( n56190 , n56099 , n56189 );
and ( n56191 , n56096 , n56190 );
or ( n56192 , n56095 , n56191 );
and ( n56193 , n56092 , n56192 );
or ( n56194 , n56091 , n56193 );
and ( n56195 , n56088 , n56194 );
or ( n56196 , n56087 , n56195 );
and ( n56197 , n56084 , n56196 );
or ( n56198 , n56083 , n56197 );
and ( n56199 , n56080 , n56198 );
or ( n56200 , n56079 , n56199 );
and ( n56201 , n56076 , n56200 );
or ( n56202 , n56075 , n56201 );
and ( n56203 , n56072 , n56202 );
or ( n56204 , n56071 , n56203 );
and ( n56205 , n56068 , n56204 );
or ( n56206 , n56067 , n56205 );
and ( n56207 , n56064 , n56206 );
or ( n56208 , n56063 , n56207 );
and ( n56209 , n56060 , n56208 );
or ( n56210 , n56059 , n56209 );
and ( n56211 , n56056 , n56210 );
or ( n56212 , n56055 , n56211 );
and ( n56213 , n56052 , n56212 );
or ( n56214 , n56051 , n56213 );
and ( n56215 , n56048 , n56214 );
or ( n56216 , n56047 , n56215 );
and ( n56217 , n56044 , n56216 );
or ( n56218 , n56043 , n56217 );
and ( n56219 , n56040 , n56218 );
or ( n56220 , n56039 , n56219 );
and ( n56221 , n56036 , n56220 );
or ( n56222 , n56035 , n56221 );
and ( n56223 , n56032 , n56222 );
or ( n56224 , n56031 , n56223 );
and ( n56225 , n56028 , n56224 );
or ( n56226 , n56027 , n56225 );
and ( n56227 , n56024 , n56226 );
or ( n56228 , n56023 , n56227 );
and ( n56229 , n56020 , n56228 );
or ( n56230 , n56019 , n56229 );
and ( n56231 , n56016 , n56230 );
or ( n56232 , n56015 , n56231 );
and ( n56233 , n56012 , n56232 );
or ( n56234 , n56011 , n56233 );
and ( n56235 , n56008 , n56234 );
or ( n56236 , n56007 , n56235 );
and ( n56237 , n56004 , n56236 );
or ( n56238 , n56003 , n56237 );
and ( n56239 , n56000 , n56238 );
or ( n56240 , n55999 , n56239 );
and ( n56241 , n55996 , n56240 );
or ( n56242 , n55995 , n56241 );
and ( n56243 , n55992 , n56242 );
or ( n56244 , n55991 , n56243 );
and ( n56245 , n55988 , n56244 );
or ( n56246 , n55987 , n56245 );
and ( n56247 , n55984 , n56246 );
or ( n56248 , n55983 , n56247 );
and ( n56249 , n55980 , n56248 );
or ( n56250 , n55979 , n56249 );
and ( n56251 , n55976 , n56250 );
or ( n56252 , n55975 , n56251 );
and ( n56253 , n55972 , n56252 );
or ( n56254 , n55971 , n56253 );
and ( n56255 , n55968 , n56254 );
or ( n56256 , n55967 , n56255 );
and ( n56257 , n55964 , n56256 );
or ( n56258 , n55963 , n56257 );
and ( n56259 , n55960 , n56258 );
or ( n56260 , n55959 , n56259 );
and ( n56261 , n55956 , n56260 );
or ( n56262 , n55955 , n56261 );
and ( n56263 , n55952 , n56262 );
or ( n56264 , n55951 , n56263 );
and ( n56265 , n55948 , n56264 );
or ( n56266 , n55947 , n56265 );
and ( n56267 , n55944 , n56266 );
or ( n56268 , n55943 , n56267 );
and ( n56269 , n55940 , n56268 );
or ( n56270 , n55939 , n56269 );
and ( n56271 , n55936 , n56270 );
or ( n56272 , n55935 , n56271 );
and ( n56273 , n55932 , n56272 );
or ( n56274 , n55931 , n56273 );
and ( n56275 , n55928 , n56274 );
or ( n56276 , n55927 , n56275 );
and ( n56277 , n55924 , n56276 );
or ( n56278 , n55923 , n56277 );
and ( n56279 , n55920 , n56278 );
or ( n56280 , n55919 , n56279 );
and ( n56281 , n55916 , n56280 );
or ( n56282 , n55915 , n56281 );
and ( n56283 , n55912 , n56282 );
or ( n56284 , n55911 , n56283 );
and ( n56285 , n55908 , n56284 );
or ( n56286 , n55907 , n56285 );
and ( n56287 , n55904 , n56286 );
or ( n56288 , n55903 , n56287 );
and ( n56289 , n55900 , n56288 );
or ( n56290 , n55899 , n56289 );
and ( n56291 , n55896 , n56290 );
or ( n56292 , n55895 , n56291 );
and ( n56293 , n55892 , n56292 );
or ( n56294 , n55891 , n56293 );
and ( n56295 , n55888 , n56294 );
or ( n56296 , n55887 , n56295 );
and ( n56297 , n55884 , n56296 );
or ( n56298 , n55883 , n56297 );
and ( n56299 , n55880 , n56298 );
or ( n56300 , n55879 , n56299 );
and ( n56301 , n55876 , n56300 );
or ( n56302 , n55875 , n56301 );
and ( n56303 , n55872 , n56302 );
or ( n56304 , n55871 , n56303 );
and ( n56305 , n55868 , n56304 );
or ( n56306 , n55867 , n56305 );
and ( n56307 , n55864 , n56306 );
or ( n56308 , n55863 , n56307 );
and ( n56309 , n55860 , n56308 );
or ( n56310 , n55859 , n56309 );
and ( n56311 , n55856 , n56310 );
or ( n56312 , n55855 , n56311 );
and ( n56313 , n55852 , n56312 );
or ( n56314 , n55851 , n56313 );
and ( n56315 , n55848 , n56314 );
or ( n56316 , n55847 , n56315 );
and ( n56317 , n55844 , n56316 );
or ( n56318 , n55843 , n56317 );
and ( n56319 , n55840 , n56318 );
or ( n56320 , n55839 , n56319 );
and ( n56321 , n55836 , n56320 );
or ( n56322 , n55835 , n56321 );
and ( n56323 , n55832 , n56322 );
or ( n56324 , n55831 , n56323 );
and ( n56325 , n55828 , n56324 );
or ( n56326 , n55827 , n56325 );
xor ( n56327 , n55824 , n56326 );
buf ( n56328 , n18020 );
and ( n56329 , n29994 , n56328 );
xor ( n56330 , n56327 , n56329 );
xor ( n56331 , n55828 , n56324 );
and ( n56332 , n29999 , n56328 );
and ( n56333 , n56331 , n56332 );
xor ( n56334 , n56331 , n56332 );
xor ( n56335 , n55832 , n56322 );
and ( n56336 , n30004 , n56328 );
and ( n56337 , n56335 , n56336 );
xor ( n56338 , n56335 , n56336 );
xor ( n56339 , n55836 , n56320 );
and ( n56340 , n30009 , n56328 );
and ( n56341 , n56339 , n56340 );
xor ( n56342 , n56339 , n56340 );
xor ( n56343 , n55840 , n56318 );
and ( n56344 , n30014 , n56328 );
and ( n56345 , n56343 , n56344 );
xor ( n56346 , n56343 , n56344 );
xor ( n56347 , n55844 , n56316 );
and ( n56348 , n30019 , n56328 );
and ( n56349 , n56347 , n56348 );
xor ( n56350 , n56347 , n56348 );
xor ( n56351 , n55848 , n56314 );
and ( n56352 , n30024 , n56328 );
and ( n56353 , n56351 , n56352 );
xor ( n56354 , n56351 , n56352 );
xor ( n56355 , n55852 , n56312 );
and ( n56356 , n30029 , n56328 );
and ( n56357 , n56355 , n56356 );
xor ( n56358 , n56355 , n56356 );
xor ( n56359 , n55856 , n56310 );
and ( n56360 , n30034 , n56328 );
and ( n56361 , n56359 , n56360 );
xor ( n56362 , n56359 , n56360 );
xor ( n56363 , n55860 , n56308 );
and ( n56364 , n30039 , n56328 );
and ( n56365 , n56363 , n56364 );
xor ( n56366 , n56363 , n56364 );
xor ( n56367 , n55864 , n56306 );
and ( n56368 , n30044 , n56328 );
and ( n56369 , n56367 , n56368 );
xor ( n56370 , n56367 , n56368 );
xor ( n56371 , n55868 , n56304 );
and ( n56372 , n30049 , n56328 );
and ( n56373 , n56371 , n56372 );
xor ( n56374 , n56371 , n56372 );
xor ( n56375 , n55872 , n56302 );
and ( n56376 , n30054 , n56328 );
and ( n56377 , n56375 , n56376 );
xor ( n56378 , n56375 , n56376 );
xor ( n56379 , n55876 , n56300 );
and ( n56380 , n30059 , n56328 );
and ( n56381 , n56379 , n56380 );
xor ( n56382 , n56379 , n56380 );
xor ( n56383 , n55880 , n56298 );
and ( n56384 , n30064 , n56328 );
and ( n56385 , n56383 , n56384 );
xor ( n56386 , n56383 , n56384 );
xor ( n56387 , n55884 , n56296 );
and ( n56388 , n30069 , n56328 );
and ( n56389 , n56387 , n56388 );
xor ( n56390 , n56387 , n56388 );
xor ( n56391 , n55888 , n56294 );
and ( n56392 , n30074 , n56328 );
and ( n56393 , n56391 , n56392 );
xor ( n56394 , n56391 , n56392 );
xor ( n56395 , n55892 , n56292 );
and ( n56396 , n30079 , n56328 );
and ( n56397 , n56395 , n56396 );
xor ( n56398 , n56395 , n56396 );
xor ( n56399 , n55896 , n56290 );
and ( n56400 , n30084 , n56328 );
and ( n56401 , n56399 , n56400 );
xor ( n56402 , n56399 , n56400 );
xor ( n56403 , n55900 , n56288 );
and ( n56404 , n30089 , n56328 );
and ( n56405 , n56403 , n56404 );
xor ( n56406 , n56403 , n56404 );
xor ( n56407 , n55904 , n56286 );
and ( n56408 , n30094 , n56328 );
and ( n56409 , n56407 , n56408 );
xor ( n56410 , n56407 , n56408 );
xor ( n56411 , n55908 , n56284 );
and ( n56412 , n30099 , n56328 );
and ( n56413 , n56411 , n56412 );
xor ( n56414 , n56411 , n56412 );
xor ( n56415 , n55912 , n56282 );
and ( n56416 , n30104 , n56328 );
and ( n56417 , n56415 , n56416 );
xor ( n56418 , n56415 , n56416 );
xor ( n56419 , n55916 , n56280 );
and ( n56420 , n30109 , n56328 );
and ( n56421 , n56419 , n56420 );
xor ( n56422 , n56419 , n56420 );
xor ( n56423 , n55920 , n56278 );
and ( n56424 , n30114 , n56328 );
and ( n56425 , n56423 , n56424 );
xor ( n56426 , n56423 , n56424 );
xor ( n56427 , n55924 , n56276 );
and ( n56428 , n30119 , n56328 );
and ( n56429 , n56427 , n56428 );
xor ( n56430 , n56427 , n56428 );
xor ( n56431 , n55928 , n56274 );
and ( n56432 , n30124 , n56328 );
and ( n56433 , n56431 , n56432 );
xor ( n56434 , n56431 , n56432 );
xor ( n56435 , n55932 , n56272 );
and ( n56436 , n30129 , n56328 );
and ( n56437 , n56435 , n56436 );
xor ( n56438 , n56435 , n56436 );
xor ( n56439 , n55936 , n56270 );
and ( n56440 , n30134 , n56328 );
and ( n56441 , n56439 , n56440 );
xor ( n56442 , n56439 , n56440 );
xor ( n56443 , n55940 , n56268 );
and ( n56444 , n30139 , n56328 );
and ( n56445 , n56443 , n56444 );
xor ( n56446 , n56443 , n56444 );
xor ( n56447 , n55944 , n56266 );
and ( n56448 , n30144 , n56328 );
and ( n56449 , n56447 , n56448 );
xor ( n56450 , n56447 , n56448 );
xor ( n56451 , n55948 , n56264 );
and ( n56452 , n30149 , n56328 );
and ( n56453 , n56451 , n56452 );
xor ( n56454 , n56451 , n56452 );
xor ( n56455 , n55952 , n56262 );
and ( n56456 , n30154 , n56328 );
and ( n56457 , n56455 , n56456 );
xor ( n56458 , n56455 , n56456 );
xor ( n56459 , n55956 , n56260 );
and ( n56460 , n30159 , n56328 );
and ( n56461 , n56459 , n56460 );
xor ( n56462 , n56459 , n56460 );
xor ( n56463 , n55960 , n56258 );
and ( n56464 , n30164 , n56328 );
and ( n56465 , n56463 , n56464 );
xor ( n56466 , n56463 , n56464 );
xor ( n56467 , n55964 , n56256 );
and ( n56468 , n30169 , n56328 );
and ( n56469 , n56467 , n56468 );
xor ( n56470 , n56467 , n56468 );
xor ( n56471 , n55968 , n56254 );
and ( n56472 , n30174 , n56328 );
and ( n56473 , n56471 , n56472 );
xor ( n56474 , n56471 , n56472 );
xor ( n56475 , n55972 , n56252 );
and ( n56476 , n30179 , n56328 );
and ( n56477 , n56475 , n56476 );
xor ( n56478 , n56475 , n56476 );
xor ( n56479 , n55976 , n56250 );
and ( n56480 , n30184 , n56328 );
and ( n56481 , n56479 , n56480 );
xor ( n56482 , n56479 , n56480 );
xor ( n56483 , n55980 , n56248 );
and ( n56484 , n30189 , n56328 );
and ( n56485 , n56483 , n56484 );
xor ( n56486 , n56483 , n56484 );
xor ( n56487 , n55984 , n56246 );
and ( n56488 , n30194 , n56328 );
and ( n56489 , n56487 , n56488 );
xor ( n56490 , n56487 , n56488 );
xor ( n56491 , n55988 , n56244 );
and ( n56492 , n30199 , n56328 );
and ( n56493 , n56491 , n56492 );
xor ( n56494 , n56491 , n56492 );
xor ( n56495 , n55992 , n56242 );
and ( n56496 , n30204 , n56328 );
and ( n56497 , n56495 , n56496 );
xor ( n56498 , n56495 , n56496 );
xor ( n56499 , n55996 , n56240 );
and ( n56500 , n30209 , n56328 );
and ( n56501 , n56499 , n56500 );
xor ( n56502 , n56499 , n56500 );
xor ( n56503 , n56000 , n56238 );
and ( n56504 , n30214 , n56328 );
and ( n56505 , n56503 , n56504 );
xor ( n56506 , n56503 , n56504 );
xor ( n56507 , n56004 , n56236 );
and ( n56508 , n30219 , n56328 );
and ( n56509 , n56507 , n56508 );
xor ( n56510 , n56507 , n56508 );
xor ( n56511 , n56008 , n56234 );
and ( n56512 , n30224 , n56328 );
and ( n56513 , n56511 , n56512 );
xor ( n56514 , n56511 , n56512 );
xor ( n56515 , n56012 , n56232 );
and ( n56516 , n30229 , n56328 );
and ( n56517 , n56515 , n56516 );
xor ( n56518 , n56515 , n56516 );
xor ( n56519 , n56016 , n56230 );
and ( n56520 , n30234 , n56328 );
and ( n56521 , n56519 , n56520 );
xor ( n56522 , n56519 , n56520 );
xor ( n56523 , n56020 , n56228 );
and ( n56524 , n30239 , n56328 );
and ( n56525 , n56523 , n56524 );
xor ( n56526 , n56523 , n56524 );
xor ( n56527 , n56024 , n56226 );
and ( n56528 , n30244 , n56328 );
and ( n56529 , n56527 , n56528 );
xor ( n56530 , n56527 , n56528 );
xor ( n56531 , n56028 , n56224 );
and ( n56532 , n30249 , n56328 );
and ( n56533 , n56531 , n56532 );
xor ( n56534 , n56531 , n56532 );
xor ( n56535 , n56032 , n56222 );
and ( n56536 , n30254 , n56328 );
and ( n56537 , n56535 , n56536 );
xor ( n56538 , n56535 , n56536 );
xor ( n56539 , n56036 , n56220 );
and ( n56540 , n30259 , n56328 );
and ( n56541 , n56539 , n56540 );
xor ( n56542 , n56539 , n56540 );
xor ( n56543 , n56040 , n56218 );
and ( n56544 , n30264 , n56328 );
and ( n56545 , n56543 , n56544 );
xor ( n56546 , n56543 , n56544 );
xor ( n56547 , n56044 , n56216 );
and ( n56548 , n30269 , n56328 );
and ( n56549 , n56547 , n56548 );
xor ( n56550 , n56547 , n56548 );
xor ( n56551 , n56048 , n56214 );
and ( n56552 , n30274 , n56328 );
and ( n56553 , n56551 , n56552 );
xor ( n56554 , n56551 , n56552 );
xor ( n56555 , n56052 , n56212 );
and ( n56556 , n30279 , n56328 );
and ( n56557 , n56555 , n56556 );
xor ( n56558 , n56555 , n56556 );
xor ( n56559 , n56056 , n56210 );
and ( n56560 , n30284 , n56328 );
and ( n56561 , n56559 , n56560 );
xor ( n56562 , n56559 , n56560 );
xor ( n56563 , n56060 , n56208 );
and ( n56564 , n30289 , n56328 );
and ( n56565 , n56563 , n56564 );
xor ( n56566 , n56563 , n56564 );
xor ( n56567 , n56064 , n56206 );
and ( n56568 , n30294 , n56328 );
and ( n56569 , n56567 , n56568 );
xor ( n56570 , n56567 , n56568 );
xor ( n56571 , n56068 , n56204 );
and ( n56572 , n30299 , n56328 );
and ( n56573 , n56571 , n56572 );
xor ( n56574 , n56571 , n56572 );
xor ( n56575 , n56072 , n56202 );
and ( n56576 , n30304 , n56328 );
and ( n56577 , n56575 , n56576 );
xor ( n56578 , n56575 , n56576 );
xor ( n56579 , n56076 , n56200 );
and ( n56580 , n30309 , n56328 );
and ( n56581 , n56579 , n56580 );
xor ( n56582 , n56579 , n56580 );
xor ( n56583 , n56080 , n56198 );
and ( n56584 , n30314 , n56328 );
and ( n56585 , n56583 , n56584 );
xor ( n56586 , n56583 , n56584 );
xor ( n56587 , n56084 , n56196 );
and ( n56588 , n30319 , n56328 );
and ( n56589 , n56587 , n56588 );
xor ( n56590 , n56587 , n56588 );
xor ( n56591 , n56088 , n56194 );
and ( n56592 , n30324 , n56328 );
and ( n56593 , n56591 , n56592 );
xor ( n56594 , n56591 , n56592 );
xor ( n56595 , n56092 , n56192 );
and ( n56596 , n30329 , n56328 );
and ( n56597 , n56595 , n56596 );
xor ( n56598 , n56595 , n56596 );
xor ( n56599 , n56096 , n56190 );
and ( n56600 , n30334 , n56328 );
and ( n56601 , n56599 , n56600 );
xor ( n56602 , n56599 , n56600 );
xor ( n56603 , n56100 , n56188 );
and ( n56604 , n30339 , n56328 );
and ( n56605 , n56603 , n56604 );
xor ( n56606 , n56603 , n56604 );
xor ( n56607 , n56104 , n56186 );
and ( n56608 , n30344 , n56328 );
and ( n56609 , n56607 , n56608 );
xor ( n56610 , n56607 , n56608 );
xor ( n56611 , n56108 , n56184 );
and ( n56612 , n30349 , n56328 );
and ( n56613 , n56611 , n56612 );
xor ( n56614 , n56611 , n56612 );
xor ( n56615 , n56112 , n56182 );
and ( n56616 , n30354 , n56328 );
and ( n56617 , n56615 , n56616 );
xor ( n56618 , n56615 , n56616 );
xor ( n56619 , n56116 , n56180 );
and ( n56620 , n30359 , n56328 );
and ( n56621 , n56619 , n56620 );
xor ( n56622 , n56619 , n56620 );
xor ( n56623 , n56120 , n56178 );
and ( n56624 , n30364 , n56328 );
and ( n56625 , n56623 , n56624 );
xor ( n56626 , n56623 , n56624 );
xor ( n56627 , n56124 , n56176 );
and ( n56628 , n30369 , n56328 );
and ( n56629 , n56627 , n56628 );
xor ( n56630 , n56627 , n56628 );
xor ( n56631 , n56128 , n56174 );
and ( n56632 , n30374 , n56328 );
and ( n56633 , n56631 , n56632 );
xor ( n56634 , n56631 , n56632 );
xor ( n56635 , n56132 , n56172 );
and ( n56636 , n30379 , n56328 );
and ( n56637 , n56635 , n56636 );
xor ( n56638 , n56635 , n56636 );
xor ( n56639 , n56136 , n56170 );
and ( n56640 , n30384 , n56328 );
and ( n56641 , n56639 , n56640 );
xor ( n56642 , n56639 , n56640 );
xor ( n56643 , n56140 , n56168 );
and ( n56644 , n30389 , n56328 );
and ( n56645 , n56643 , n56644 );
xor ( n56646 , n56643 , n56644 );
xor ( n56647 , n56144 , n56166 );
and ( n56648 , n30394 , n56328 );
and ( n56649 , n56647 , n56648 );
xor ( n56650 , n56647 , n56648 );
xor ( n56651 , n56148 , n56164 );
and ( n56652 , n30399 , n56328 );
and ( n56653 , n56651 , n56652 );
xor ( n56654 , n56651 , n56652 );
xor ( n56655 , n56152 , n56162 );
and ( n56656 , n30404 , n56328 );
and ( n56657 , n56655 , n56656 );
xor ( n56658 , n56655 , n56656 );
xor ( n56659 , n56156 , n56160 );
and ( n56660 , n30409 , n56328 );
and ( n56661 , n56659 , n56660 );
buf ( n56662 , n56661 );
and ( n56663 , n56658 , n56662 );
or ( n56664 , n56657 , n56663 );
and ( n56665 , n56654 , n56664 );
or ( n56666 , n56653 , n56665 );
and ( n56667 , n56650 , n56666 );
or ( n56668 , n56649 , n56667 );
and ( n56669 , n56646 , n56668 );
or ( n56670 , n56645 , n56669 );
and ( n56671 , n56642 , n56670 );
or ( n56672 , n56641 , n56671 );
and ( n56673 , n56638 , n56672 );
or ( n56674 , n56637 , n56673 );
and ( n56675 , n56634 , n56674 );
or ( n56676 , n56633 , n56675 );
and ( n56677 , n56630 , n56676 );
or ( n56678 , n56629 , n56677 );
and ( n56679 , n56626 , n56678 );
or ( n56680 , n56625 , n56679 );
and ( n56681 , n56622 , n56680 );
or ( n56682 , n56621 , n56681 );
and ( n56683 , n56618 , n56682 );
or ( n56684 , n56617 , n56683 );
and ( n56685 , n56614 , n56684 );
or ( n56686 , n56613 , n56685 );
and ( n56687 , n56610 , n56686 );
or ( n56688 , n56609 , n56687 );
and ( n56689 , n56606 , n56688 );
or ( n56690 , n56605 , n56689 );
and ( n56691 , n56602 , n56690 );
or ( n56692 , n56601 , n56691 );
and ( n56693 , n56598 , n56692 );
or ( n56694 , n56597 , n56693 );
and ( n56695 , n56594 , n56694 );
or ( n56696 , n56593 , n56695 );
and ( n56697 , n56590 , n56696 );
or ( n56698 , n56589 , n56697 );
and ( n56699 , n56586 , n56698 );
or ( n56700 , n56585 , n56699 );
and ( n56701 , n56582 , n56700 );
or ( n56702 , n56581 , n56701 );
and ( n56703 , n56578 , n56702 );
or ( n56704 , n56577 , n56703 );
and ( n56705 , n56574 , n56704 );
or ( n56706 , n56573 , n56705 );
and ( n56707 , n56570 , n56706 );
or ( n56708 , n56569 , n56707 );
and ( n56709 , n56566 , n56708 );
or ( n56710 , n56565 , n56709 );
and ( n56711 , n56562 , n56710 );
or ( n56712 , n56561 , n56711 );
and ( n56713 , n56558 , n56712 );
or ( n56714 , n56557 , n56713 );
and ( n56715 , n56554 , n56714 );
or ( n56716 , n56553 , n56715 );
and ( n56717 , n56550 , n56716 );
or ( n56718 , n56549 , n56717 );
and ( n56719 , n56546 , n56718 );
or ( n56720 , n56545 , n56719 );
and ( n56721 , n56542 , n56720 );
or ( n56722 , n56541 , n56721 );
and ( n56723 , n56538 , n56722 );
or ( n56724 , n56537 , n56723 );
and ( n56725 , n56534 , n56724 );
or ( n56726 , n56533 , n56725 );
and ( n56727 , n56530 , n56726 );
or ( n56728 , n56529 , n56727 );
and ( n56729 , n56526 , n56728 );
or ( n56730 , n56525 , n56729 );
and ( n56731 , n56522 , n56730 );
or ( n56732 , n56521 , n56731 );
and ( n56733 , n56518 , n56732 );
or ( n56734 , n56517 , n56733 );
and ( n56735 , n56514 , n56734 );
or ( n56736 , n56513 , n56735 );
and ( n56737 , n56510 , n56736 );
or ( n56738 , n56509 , n56737 );
and ( n56739 , n56506 , n56738 );
or ( n56740 , n56505 , n56739 );
and ( n56741 , n56502 , n56740 );
or ( n56742 , n56501 , n56741 );
and ( n56743 , n56498 , n56742 );
or ( n56744 , n56497 , n56743 );
and ( n56745 , n56494 , n56744 );
or ( n56746 , n56493 , n56745 );
and ( n56747 , n56490 , n56746 );
or ( n56748 , n56489 , n56747 );
and ( n56749 , n56486 , n56748 );
or ( n56750 , n56485 , n56749 );
and ( n56751 , n56482 , n56750 );
or ( n56752 , n56481 , n56751 );
and ( n56753 , n56478 , n56752 );
or ( n56754 , n56477 , n56753 );
and ( n56755 , n56474 , n56754 );
or ( n56756 , n56473 , n56755 );
and ( n56757 , n56470 , n56756 );
or ( n56758 , n56469 , n56757 );
and ( n56759 , n56466 , n56758 );
or ( n56760 , n56465 , n56759 );
and ( n56761 , n56462 , n56760 );
or ( n56762 , n56461 , n56761 );
and ( n56763 , n56458 , n56762 );
or ( n56764 , n56457 , n56763 );
and ( n56765 , n56454 , n56764 );
or ( n56766 , n56453 , n56765 );
and ( n56767 , n56450 , n56766 );
or ( n56768 , n56449 , n56767 );
and ( n56769 , n56446 , n56768 );
or ( n56770 , n56445 , n56769 );
and ( n56771 , n56442 , n56770 );
or ( n56772 , n56441 , n56771 );
and ( n56773 , n56438 , n56772 );
or ( n56774 , n56437 , n56773 );
and ( n56775 , n56434 , n56774 );
or ( n56776 , n56433 , n56775 );
and ( n56777 , n56430 , n56776 );
or ( n56778 , n56429 , n56777 );
and ( n56779 , n56426 , n56778 );
or ( n56780 , n56425 , n56779 );
and ( n56781 , n56422 , n56780 );
or ( n56782 , n56421 , n56781 );
and ( n56783 , n56418 , n56782 );
or ( n56784 , n56417 , n56783 );
and ( n56785 , n56414 , n56784 );
or ( n56786 , n56413 , n56785 );
and ( n56787 , n56410 , n56786 );
or ( n56788 , n56409 , n56787 );
and ( n56789 , n56406 , n56788 );
or ( n56790 , n56405 , n56789 );
and ( n56791 , n56402 , n56790 );
or ( n56792 , n56401 , n56791 );
and ( n56793 , n56398 , n56792 );
or ( n56794 , n56397 , n56793 );
and ( n56795 , n56394 , n56794 );
or ( n56796 , n56393 , n56795 );
and ( n56797 , n56390 , n56796 );
or ( n56798 , n56389 , n56797 );
and ( n56799 , n56386 , n56798 );
or ( n56800 , n56385 , n56799 );
and ( n56801 , n56382 , n56800 );
or ( n56802 , n56381 , n56801 );
and ( n56803 , n56378 , n56802 );
or ( n56804 , n56377 , n56803 );
and ( n56805 , n56374 , n56804 );
or ( n56806 , n56373 , n56805 );
and ( n56807 , n56370 , n56806 );
or ( n56808 , n56369 , n56807 );
and ( n56809 , n56366 , n56808 );
or ( n56810 , n56365 , n56809 );
and ( n56811 , n56362 , n56810 );
or ( n56812 , n56361 , n56811 );
and ( n56813 , n56358 , n56812 );
or ( n56814 , n56357 , n56813 );
and ( n56815 , n56354 , n56814 );
or ( n56816 , n56353 , n56815 );
and ( n56817 , n56350 , n56816 );
or ( n56818 , n56349 , n56817 );
and ( n56819 , n56346 , n56818 );
or ( n56820 , n56345 , n56819 );
and ( n56821 , n56342 , n56820 );
or ( n56822 , n56341 , n56821 );
and ( n56823 , n56338 , n56822 );
or ( n56824 , n56337 , n56823 );
and ( n56825 , n56334 , n56824 );
or ( n56826 , n56333 , n56825 );
xor ( n56827 , n56330 , n56826 );
buf ( n56828 , n18018 );
and ( n56829 , n29999 , n56828 );
xor ( n56830 , n56827 , n56829 );
xor ( n56831 , n56334 , n56824 );
and ( n56832 , n30004 , n56828 );
and ( n56833 , n56831 , n56832 );
xor ( n56834 , n56831 , n56832 );
xor ( n56835 , n56338 , n56822 );
and ( n56836 , n30009 , n56828 );
and ( n56837 , n56835 , n56836 );
xor ( n56838 , n56835 , n56836 );
xor ( n56839 , n56342 , n56820 );
and ( n56840 , n30014 , n56828 );
and ( n56841 , n56839 , n56840 );
xor ( n56842 , n56839 , n56840 );
xor ( n56843 , n56346 , n56818 );
and ( n56844 , n30019 , n56828 );
and ( n56845 , n56843 , n56844 );
xor ( n56846 , n56843 , n56844 );
xor ( n56847 , n56350 , n56816 );
and ( n56848 , n30024 , n56828 );
and ( n56849 , n56847 , n56848 );
xor ( n56850 , n56847 , n56848 );
xor ( n56851 , n56354 , n56814 );
and ( n56852 , n30029 , n56828 );
and ( n56853 , n56851 , n56852 );
xor ( n56854 , n56851 , n56852 );
xor ( n56855 , n56358 , n56812 );
and ( n56856 , n30034 , n56828 );
and ( n56857 , n56855 , n56856 );
xor ( n56858 , n56855 , n56856 );
xor ( n56859 , n56362 , n56810 );
and ( n56860 , n30039 , n56828 );
and ( n56861 , n56859 , n56860 );
xor ( n56862 , n56859 , n56860 );
xor ( n56863 , n56366 , n56808 );
and ( n56864 , n30044 , n56828 );
and ( n56865 , n56863 , n56864 );
xor ( n56866 , n56863 , n56864 );
xor ( n56867 , n56370 , n56806 );
and ( n56868 , n30049 , n56828 );
and ( n56869 , n56867 , n56868 );
xor ( n56870 , n56867 , n56868 );
xor ( n56871 , n56374 , n56804 );
and ( n56872 , n30054 , n56828 );
and ( n56873 , n56871 , n56872 );
xor ( n56874 , n56871 , n56872 );
xor ( n56875 , n56378 , n56802 );
and ( n56876 , n30059 , n56828 );
and ( n56877 , n56875 , n56876 );
xor ( n56878 , n56875 , n56876 );
xor ( n56879 , n56382 , n56800 );
and ( n56880 , n30064 , n56828 );
and ( n56881 , n56879 , n56880 );
xor ( n56882 , n56879 , n56880 );
xor ( n56883 , n56386 , n56798 );
and ( n56884 , n30069 , n56828 );
and ( n56885 , n56883 , n56884 );
xor ( n56886 , n56883 , n56884 );
xor ( n56887 , n56390 , n56796 );
and ( n56888 , n30074 , n56828 );
and ( n56889 , n56887 , n56888 );
xor ( n56890 , n56887 , n56888 );
xor ( n56891 , n56394 , n56794 );
and ( n56892 , n30079 , n56828 );
and ( n56893 , n56891 , n56892 );
xor ( n56894 , n56891 , n56892 );
xor ( n56895 , n56398 , n56792 );
and ( n56896 , n30084 , n56828 );
and ( n56897 , n56895 , n56896 );
xor ( n56898 , n56895 , n56896 );
xor ( n56899 , n56402 , n56790 );
and ( n56900 , n30089 , n56828 );
and ( n56901 , n56899 , n56900 );
xor ( n56902 , n56899 , n56900 );
xor ( n56903 , n56406 , n56788 );
and ( n56904 , n30094 , n56828 );
and ( n56905 , n56903 , n56904 );
xor ( n56906 , n56903 , n56904 );
xor ( n56907 , n56410 , n56786 );
and ( n56908 , n30099 , n56828 );
and ( n56909 , n56907 , n56908 );
xor ( n56910 , n56907 , n56908 );
xor ( n56911 , n56414 , n56784 );
and ( n56912 , n30104 , n56828 );
and ( n56913 , n56911 , n56912 );
xor ( n56914 , n56911 , n56912 );
xor ( n56915 , n56418 , n56782 );
and ( n56916 , n30109 , n56828 );
and ( n56917 , n56915 , n56916 );
xor ( n56918 , n56915 , n56916 );
xor ( n56919 , n56422 , n56780 );
and ( n56920 , n30114 , n56828 );
and ( n56921 , n56919 , n56920 );
xor ( n56922 , n56919 , n56920 );
xor ( n56923 , n56426 , n56778 );
and ( n56924 , n30119 , n56828 );
and ( n56925 , n56923 , n56924 );
xor ( n56926 , n56923 , n56924 );
xor ( n56927 , n56430 , n56776 );
and ( n56928 , n30124 , n56828 );
and ( n56929 , n56927 , n56928 );
xor ( n56930 , n56927 , n56928 );
xor ( n56931 , n56434 , n56774 );
and ( n56932 , n30129 , n56828 );
and ( n56933 , n56931 , n56932 );
xor ( n56934 , n56931 , n56932 );
xor ( n56935 , n56438 , n56772 );
and ( n56936 , n30134 , n56828 );
and ( n56937 , n56935 , n56936 );
xor ( n56938 , n56935 , n56936 );
xor ( n56939 , n56442 , n56770 );
and ( n56940 , n30139 , n56828 );
and ( n56941 , n56939 , n56940 );
xor ( n56942 , n56939 , n56940 );
xor ( n56943 , n56446 , n56768 );
and ( n56944 , n30144 , n56828 );
and ( n56945 , n56943 , n56944 );
xor ( n56946 , n56943 , n56944 );
xor ( n56947 , n56450 , n56766 );
and ( n56948 , n30149 , n56828 );
and ( n56949 , n56947 , n56948 );
xor ( n56950 , n56947 , n56948 );
xor ( n56951 , n56454 , n56764 );
and ( n56952 , n30154 , n56828 );
and ( n56953 , n56951 , n56952 );
xor ( n56954 , n56951 , n56952 );
xor ( n56955 , n56458 , n56762 );
and ( n56956 , n30159 , n56828 );
and ( n56957 , n56955 , n56956 );
xor ( n56958 , n56955 , n56956 );
xor ( n56959 , n56462 , n56760 );
and ( n56960 , n30164 , n56828 );
and ( n56961 , n56959 , n56960 );
xor ( n56962 , n56959 , n56960 );
xor ( n56963 , n56466 , n56758 );
and ( n56964 , n30169 , n56828 );
and ( n56965 , n56963 , n56964 );
xor ( n56966 , n56963 , n56964 );
xor ( n56967 , n56470 , n56756 );
and ( n56968 , n30174 , n56828 );
and ( n56969 , n56967 , n56968 );
xor ( n56970 , n56967 , n56968 );
xor ( n56971 , n56474 , n56754 );
and ( n56972 , n30179 , n56828 );
and ( n56973 , n56971 , n56972 );
xor ( n56974 , n56971 , n56972 );
xor ( n56975 , n56478 , n56752 );
and ( n56976 , n30184 , n56828 );
and ( n56977 , n56975 , n56976 );
xor ( n56978 , n56975 , n56976 );
xor ( n56979 , n56482 , n56750 );
and ( n56980 , n30189 , n56828 );
and ( n56981 , n56979 , n56980 );
xor ( n56982 , n56979 , n56980 );
xor ( n56983 , n56486 , n56748 );
and ( n56984 , n30194 , n56828 );
and ( n56985 , n56983 , n56984 );
xor ( n56986 , n56983 , n56984 );
xor ( n56987 , n56490 , n56746 );
and ( n56988 , n30199 , n56828 );
and ( n56989 , n56987 , n56988 );
xor ( n56990 , n56987 , n56988 );
xor ( n56991 , n56494 , n56744 );
and ( n56992 , n30204 , n56828 );
and ( n56993 , n56991 , n56992 );
xor ( n56994 , n56991 , n56992 );
xor ( n56995 , n56498 , n56742 );
and ( n56996 , n30209 , n56828 );
and ( n56997 , n56995 , n56996 );
xor ( n56998 , n56995 , n56996 );
xor ( n56999 , n56502 , n56740 );
and ( n57000 , n30214 , n56828 );
and ( n57001 , n56999 , n57000 );
xor ( n57002 , n56999 , n57000 );
xor ( n57003 , n56506 , n56738 );
and ( n57004 , n30219 , n56828 );
and ( n57005 , n57003 , n57004 );
xor ( n57006 , n57003 , n57004 );
xor ( n57007 , n56510 , n56736 );
and ( n57008 , n30224 , n56828 );
and ( n57009 , n57007 , n57008 );
xor ( n57010 , n57007 , n57008 );
xor ( n57011 , n56514 , n56734 );
and ( n57012 , n30229 , n56828 );
and ( n57013 , n57011 , n57012 );
xor ( n57014 , n57011 , n57012 );
xor ( n57015 , n56518 , n56732 );
and ( n57016 , n30234 , n56828 );
and ( n57017 , n57015 , n57016 );
xor ( n57018 , n57015 , n57016 );
xor ( n57019 , n56522 , n56730 );
and ( n57020 , n30239 , n56828 );
and ( n57021 , n57019 , n57020 );
xor ( n57022 , n57019 , n57020 );
xor ( n57023 , n56526 , n56728 );
and ( n57024 , n30244 , n56828 );
and ( n57025 , n57023 , n57024 );
xor ( n57026 , n57023 , n57024 );
xor ( n57027 , n56530 , n56726 );
and ( n57028 , n30249 , n56828 );
and ( n57029 , n57027 , n57028 );
xor ( n57030 , n57027 , n57028 );
xor ( n57031 , n56534 , n56724 );
and ( n57032 , n30254 , n56828 );
and ( n57033 , n57031 , n57032 );
xor ( n57034 , n57031 , n57032 );
xor ( n57035 , n56538 , n56722 );
and ( n57036 , n30259 , n56828 );
and ( n57037 , n57035 , n57036 );
xor ( n57038 , n57035 , n57036 );
xor ( n57039 , n56542 , n56720 );
and ( n57040 , n30264 , n56828 );
and ( n57041 , n57039 , n57040 );
xor ( n57042 , n57039 , n57040 );
xor ( n57043 , n56546 , n56718 );
and ( n57044 , n30269 , n56828 );
and ( n57045 , n57043 , n57044 );
xor ( n57046 , n57043 , n57044 );
xor ( n57047 , n56550 , n56716 );
and ( n57048 , n30274 , n56828 );
and ( n57049 , n57047 , n57048 );
xor ( n57050 , n57047 , n57048 );
xor ( n57051 , n56554 , n56714 );
and ( n57052 , n30279 , n56828 );
and ( n57053 , n57051 , n57052 );
xor ( n57054 , n57051 , n57052 );
xor ( n57055 , n56558 , n56712 );
and ( n57056 , n30284 , n56828 );
and ( n57057 , n57055 , n57056 );
xor ( n57058 , n57055 , n57056 );
xor ( n57059 , n56562 , n56710 );
and ( n57060 , n30289 , n56828 );
and ( n57061 , n57059 , n57060 );
xor ( n57062 , n57059 , n57060 );
xor ( n57063 , n56566 , n56708 );
and ( n57064 , n30294 , n56828 );
and ( n57065 , n57063 , n57064 );
xor ( n57066 , n57063 , n57064 );
xor ( n57067 , n56570 , n56706 );
and ( n57068 , n30299 , n56828 );
and ( n57069 , n57067 , n57068 );
xor ( n57070 , n57067 , n57068 );
xor ( n57071 , n56574 , n56704 );
and ( n57072 , n30304 , n56828 );
and ( n57073 , n57071 , n57072 );
xor ( n57074 , n57071 , n57072 );
xor ( n57075 , n56578 , n56702 );
and ( n57076 , n30309 , n56828 );
and ( n57077 , n57075 , n57076 );
xor ( n57078 , n57075 , n57076 );
xor ( n57079 , n56582 , n56700 );
and ( n57080 , n30314 , n56828 );
and ( n57081 , n57079 , n57080 );
xor ( n57082 , n57079 , n57080 );
xor ( n57083 , n56586 , n56698 );
and ( n57084 , n30319 , n56828 );
and ( n57085 , n57083 , n57084 );
xor ( n57086 , n57083 , n57084 );
xor ( n57087 , n56590 , n56696 );
and ( n57088 , n30324 , n56828 );
and ( n57089 , n57087 , n57088 );
xor ( n57090 , n57087 , n57088 );
xor ( n57091 , n56594 , n56694 );
and ( n57092 , n30329 , n56828 );
and ( n57093 , n57091 , n57092 );
xor ( n57094 , n57091 , n57092 );
xor ( n57095 , n56598 , n56692 );
and ( n57096 , n30334 , n56828 );
and ( n57097 , n57095 , n57096 );
xor ( n57098 , n57095 , n57096 );
xor ( n57099 , n56602 , n56690 );
and ( n57100 , n30339 , n56828 );
and ( n57101 , n57099 , n57100 );
xor ( n57102 , n57099 , n57100 );
xor ( n57103 , n56606 , n56688 );
and ( n57104 , n30344 , n56828 );
and ( n57105 , n57103 , n57104 );
xor ( n57106 , n57103 , n57104 );
xor ( n57107 , n56610 , n56686 );
and ( n57108 , n30349 , n56828 );
and ( n57109 , n57107 , n57108 );
xor ( n57110 , n57107 , n57108 );
xor ( n57111 , n56614 , n56684 );
and ( n57112 , n30354 , n56828 );
and ( n57113 , n57111 , n57112 );
xor ( n57114 , n57111 , n57112 );
xor ( n57115 , n56618 , n56682 );
and ( n57116 , n30359 , n56828 );
and ( n57117 , n57115 , n57116 );
xor ( n57118 , n57115 , n57116 );
xor ( n57119 , n56622 , n56680 );
and ( n57120 , n30364 , n56828 );
and ( n57121 , n57119 , n57120 );
xor ( n57122 , n57119 , n57120 );
xor ( n57123 , n56626 , n56678 );
and ( n57124 , n30369 , n56828 );
and ( n57125 , n57123 , n57124 );
xor ( n57126 , n57123 , n57124 );
xor ( n57127 , n56630 , n56676 );
and ( n57128 , n30374 , n56828 );
and ( n57129 , n57127 , n57128 );
xor ( n57130 , n57127 , n57128 );
xor ( n57131 , n56634 , n56674 );
and ( n57132 , n30379 , n56828 );
and ( n57133 , n57131 , n57132 );
xor ( n57134 , n57131 , n57132 );
xor ( n57135 , n56638 , n56672 );
and ( n57136 , n30384 , n56828 );
and ( n57137 , n57135 , n57136 );
xor ( n57138 , n57135 , n57136 );
xor ( n57139 , n56642 , n56670 );
and ( n57140 , n30389 , n56828 );
and ( n57141 , n57139 , n57140 );
xor ( n57142 , n57139 , n57140 );
xor ( n57143 , n56646 , n56668 );
and ( n57144 , n30394 , n56828 );
and ( n57145 , n57143 , n57144 );
xor ( n57146 , n57143 , n57144 );
xor ( n57147 , n56650 , n56666 );
and ( n57148 , n30399 , n56828 );
and ( n57149 , n57147 , n57148 );
xor ( n57150 , n57147 , n57148 );
xor ( n57151 , n56654 , n56664 );
and ( n57152 , n30404 , n56828 );
and ( n57153 , n57151 , n57152 );
xor ( n57154 , n57151 , n57152 );
xor ( n57155 , n56658 , n56662 );
and ( n57156 , n30409 , n56828 );
and ( n57157 , n57155 , n57156 );
buf ( n57158 , n57157 );
and ( n57159 , n57154 , n57158 );
or ( n57160 , n57153 , n57159 );
and ( n57161 , n57150 , n57160 );
or ( n57162 , n57149 , n57161 );
and ( n57163 , n57146 , n57162 );
or ( n57164 , n57145 , n57163 );
and ( n57165 , n57142 , n57164 );
or ( n57166 , n57141 , n57165 );
and ( n57167 , n57138 , n57166 );
or ( n57168 , n57137 , n57167 );
and ( n57169 , n57134 , n57168 );
or ( n57170 , n57133 , n57169 );
and ( n57171 , n57130 , n57170 );
or ( n57172 , n57129 , n57171 );
and ( n57173 , n57126 , n57172 );
or ( n57174 , n57125 , n57173 );
and ( n57175 , n57122 , n57174 );
or ( n57176 , n57121 , n57175 );
and ( n57177 , n57118 , n57176 );
or ( n57178 , n57117 , n57177 );
and ( n57179 , n57114 , n57178 );
or ( n57180 , n57113 , n57179 );
and ( n57181 , n57110 , n57180 );
or ( n57182 , n57109 , n57181 );
and ( n57183 , n57106 , n57182 );
or ( n57184 , n57105 , n57183 );
and ( n57185 , n57102 , n57184 );
or ( n57186 , n57101 , n57185 );
and ( n57187 , n57098 , n57186 );
or ( n57188 , n57097 , n57187 );
and ( n57189 , n57094 , n57188 );
or ( n57190 , n57093 , n57189 );
and ( n57191 , n57090 , n57190 );
or ( n57192 , n57089 , n57191 );
and ( n57193 , n57086 , n57192 );
or ( n57194 , n57085 , n57193 );
and ( n57195 , n57082 , n57194 );
or ( n57196 , n57081 , n57195 );
and ( n57197 , n57078 , n57196 );
or ( n57198 , n57077 , n57197 );
and ( n57199 , n57074 , n57198 );
or ( n57200 , n57073 , n57199 );
and ( n57201 , n57070 , n57200 );
or ( n57202 , n57069 , n57201 );
and ( n57203 , n57066 , n57202 );
or ( n57204 , n57065 , n57203 );
and ( n57205 , n57062 , n57204 );
or ( n57206 , n57061 , n57205 );
and ( n57207 , n57058 , n57206 );
or ( n57208 , n57057 , n57207 );
and ( n57209 , n57054 , n57208 );
or ( n57210 , n57053 , n57209 );
and ( n57211 , n57050 , n57210 );
or ( n57212 , n57049 , n57211 );
and ( n57213 , n57046 , n57212 );
or ( n57214 , n57045 , n57213 );
and ( n57215 , n57042 , n57214 );
or ( n57216 , n57041 , n57215 );
and ( n57217 , n57038 , n57216 );
or ( n57218 , n57037 , n57217 );
and ( n57219 , n57034 , n57218 );
or ( n57220 , n57033 , n57219 );
and ( n57221 , n57030 , n57220 );
or ( n57222 , n57029 , n57221 );
and ( n57223 , n57026 , n57222 );
or ( n57224 , n57025 , n57223 );
and ( n57225 , n57022 , n57224 );
or ( n57226 , n57021 , n57225 );
and ( n57227 , n57018 , n57226 );
or ( n57228 , n57017 , n57227 );
and ( n57229 , n57014 , n57228 );
or ( n57230 , n57013 , n57229 );
and ( n57231 , n57010 , n57230 );
or ( n57232 , n57009 , n57231 );
and ( n57233 , n57006 , n57232 );
or ( n57234 , n57005 , n57233 );
and ( n57235 , n57002 , n57234 );
or ( n57236 , n57001 , n57235 );
and ( n57237 , n56998 , n57236 );
or ( n57238 , n56997 , n57237 );
and ( n57239 , n56994 , n57238 );
or ( n57240 , n56993 , n57239 );
and ( n57241 , n56990 , n57240 );
or ( n57242 , n56989 , n57241 );
and ( n57243 , n56986 , n57242 );
or ( n57244 , n56985 , n57243 );
and ( n57245 , n56982 , n57244 );
or ( n57246 , n56981 , n57245 );
and ( n57247 , n56978 , n57246 );
or ( n57248 , n56977 , n57247 );
and ( n57249 , n56974 , n57248 );
or ( n57250 , n56973 , n57249 );
and ( n57251 , n56970 , n57250 );
or ( n57252 , n56969 , n57251 );
and ( n57253 , n56966 , n57252 );
or ( n57254 , n56965 , n57253 );
and ( n57255 , n56962 , n57254 );
or ( n57256 , n56961 , n57255 );
and ( n57257 , n56958 , n57256 );
or ( n57258 , n56957 , n57257 );
and ( n57259 , n56954 , n57258 );
or ( n57260 , n56953 , n57259 );
and ( n57261 , n56950 , n57260 );
or ( n57262 , n56949 , n57261 );
and ( n57263 , n56946 , n57262 );
or ( n57264 , n56945 , n57263 );
and ( n57265 , n56942 , n57264 );
or ( n57266 , n56941 , n57265 );
and ( n57267 , n56938 , n57266 );
or ( n57268 , n56937 , n57267 );
and ( n57269 , n56934 , n57268 );
or ( n57270 , n56933 , n57269 );
and ( n57271 , n56930 , n57270 );
or ( n57272 , n56929 , n57271 );
and ( n57273 , n56926 , n57272 );
or ( n57274 , n56925 , n57273 );
and ( n57275 , n56922 , n57274 );
or ( n57276 , n56921 , n57275 );
and ( n57277 , n56918 , n57276 );
or ( n57278 , n56917 , n57277 );
and ( n57279 , n56914 , n57278 );
or ( n57280 , n56913 , n57279 );
and ( n57281 , n56910 , n57280 );
or ( n57282 , n56909 , n57281 );
and ( n57283 , n56906 , n57282 );
or ( n57284 , n56905 , n57283 );
and ( n57285 , n56902 , n57284 );
or ( n57286 , n56901 , n57285 );
and ( n57287 , n56898 , n57286 );
or ( n57288 , n56897 , n57287 );
and ( n57289 , n56894 , n57288 );
or ( n57290 , n56893 , n57289 );
and ( n57291 , n56890 , n57290 );
or ( n57292 , n56889 , n57291 );
and ( n57293 , n56886 , n57292 );
or ( n57294 , n56885 , n57293 );
and ( n57295 , n56882 , n57294 );
or ( n57296 , n56881 , n57295 );
and ( n57297 , n56878 , n57296 );
or ( n57298 , n56877 , n57297 );
and ( n57299 , n56874 , n57298 );
or ( n57300 , n56873 , n57299 );
and ( n57301 , n56870 , n57300 );
or ( n57302 , n56869 , n57301 );
and ( n57303 , n56866 , n57302 );
or ( n57304 , n56865 , n57303 );
and ( n57305 , n56862 , n57304 );
or ( n57306 , n56861 , n57305 );
and ( n57307 , n56858 , n57306 );
or ( n57308 , n56857 , n57307 );
and ( n57309 , n56854 , n57308 );
or ( n57310 , n56853 , n57309 );
and ( n57311 , n56850 , n57310 );
or ( n57312 , n56849 , n57311 );
and ( n57313 , n56846 , n57312 );
or ( n57314 , n56845 , n57313 );
and ( n57315 , n56842 , n57314 );
or ( n57316 , n56841 , n57315 );
and ( n57317 , n56838 , n57316 );
or ( n57318 , n56837 , n57317 );
and ( n57319 , n56834 , n57318 );
or ( n57320 , n56833 , n57319 );
xor ( n57321 , n56830 , n57320 );
buf ( n57322 , n18016 );
and ( n57323 , n30004 , n57322 );
xor ( n57324 , n57321 , n57323 );
xor ( n57325 , n56834 , n57318 );
and ( n57326 , n30009 , n57322 );
and ( n57327 , n57325 , n57326 );
xor ( n57328 , n57325 , n57326 );
xor ( n57329 , n56838 , n57316 );
and ( n57330 , n30014 , n57322 );
and ( n57331 , n57329 , n57330 );
xor ( n57332 , n57329 , n57330 );
xor ( n57333 , n56842 , n57314 );
and ( n57334 , n30019 , n57322 );
and ( n57335 , n57333 , n57334 );
xor ( n57336 , n57333 , n57334 );
xor ( n57337 , n56846 , n57312 );
and ( n57338 , n30024 , n57322 );
and ( n57339 , n57337 , n57338 );
xor ( n57340 , n57337 , n57338 );
xor ( n57341 , n56850 , n57310 );
and ( n57342 , n30029 , n57322 );
and ( n57343 , n57341 , n57342 );
xor ( n57344 , n57341 , n57342 );
xor ( n57345 , n56854 , n57308 );
and ( n57346 , n30034 , n57322 );
and ( n57347 , n57345 , n57346 );
xor ( n57348 , n57345 , n57346 );
xor ( n57349 , n56858 , n57306 );
and ( n57350 , n30039 , n57322 );
and ( n57351 , n57349 , n57350 );
xor ( n57352 , n57349 , n57350 );
xor ( n57353 , n56862 , n57304 );
and ( n57354 , n30044 , n57322 );
and ( n57355 , n57353 , n57354 );
xor ( n57356 , n57353 , n57354 );
xor ( n57357 , n56866 , n57302 );
and ( n57358 , n30049 , n57322 );
and ( n57359 , n57357 , n57358 );
xor ( n57360 , n57357 , n57358 );
xor ( n57361 , n56870 , n57300 );
and ( n57362 , n30054 , n57322 );
and ( n57363 , n57361 , n57362 );
xor ( n57364 , n57361 , n57362 );
xor ( n57365 , n56874 , n57298 );
and ( n57366 , n30059 , n57322 );
and ( n57367 , n57365 , n57366 );
xor ( n57368 , n57365 , n57366 );
xor ( n57369 , n56878 , n57296 );
and ( n57370 , n30064 , n57322 );
and ( n57371 , n57369 , n57370 );
xor ( n57372 , n57369 , n57370 );
xor ( n57373 , n56882 , n57294 );
and ( n57374 , n30069 , n57322 );
and ( n57375 , n57373 , n57374 );
xor ( n57376 , n57373 , n57374 );
xor ( n57377 , n56886 , n57292 );
and ( n57378 , n30074 , n57322 );
and ( n57379 , n57377 , n57378 );
xor ( n57380 , n57377 , n57378 );
xor ( n57381 , n56890 , n57290 );
and ( n57382 , n30079 , n57322 );
and ( n57383 , n57381 , n57382 );
xor ( n57384 , n57381 , n57382 );
xor ( n57385 , n56894 , n57288 );
and ( n57386 , n30084 , n57322 );
and ( n57387 , n57385 , n57386 );
xor ( n57388 , n57385 , n57386 );
xor ( n57389 , n56898 , n57286 );
and ( n57390 , n30089 , n57322 );
and ( n57391 , n57389 , n57390 );
xor ( n57392 , n57389 , n57390 );
xor ( n57393 , n56902 , n57284 );
and ( n57394 , n30094 , n57322 );
and ( n57395 , n57393 , n57394 );
xor ( n57396 , n57393 , n57394 );
xor ( n57397 , n56906 , n57282 );
and ( n57398 , n30099 , n57322 );
and ( n57399 , n57397 , n57398 );
xor ( n57400 , n57397 , n57398 );
xor ( n57401 , n56910 , n57280 );
and ( n57402 , n30104 , n57322 );
and ( n57403 , n57401 , n57402 );
xor ( n57404 , n57401 , n57402 );
xor ( n57405 , n56914 , n57278 );
and ( n57406 , n30109 , n57322 );
and ( n57407 , n57405 , n57406 );
xor ( n57408 , n57405 , n57406 );
xor ( n57409 , n56918 , n57276 );
and ( n57410 , n30114 , n57322 );
and ( n57411 , n57409 , n57410 );
xor ( n57412 , n57409 , n57410 );
xor ( n57413 , n56922 , n57274 );
and ( n57414 , n30119 , n57322 );
and ( n57415 , n57413 , n57414 );
xor ( n57416 , n57413 , n57414 );
xor ( n57417 , n56926 , n57272 );
and ( n57418 , n30124 , n57322 );
and ( n57419 , n57417 , n57418 );
xor ( n57420 , n57417 , n57418 );
xor ( n57421 , n56930 , n57270 );
and ( n57422 , n30129 , n57322 );
and ( n57423 , n57421 , n57422 );
xor ( n57424 , n57421 , n57422 );
xor ( n57425 , n56934 , n57268 );
and ( n57426 , n30134 , n57322 );
and ( n57427 , n57425 , n57426 );
xor ( n57428 , n57425 , n57426 );
xor ( n57429 , n56938 , n57266 );
and ( n57430 , n30139 , n57322 );
and ( n57431 , n57429 , n57430 );
xor ( n57432 , n57429 , n57430 );
xor ( n57433 , n56942 , n57264 );
and ( n57434 , n30144 , n57322 );
and ( n57435 , n57433 , n57434 );
xor ( n57436 , n57433 , n57434 );
xor ( n57437 , n56946 , n57262 );
and ( n57438 , n30149 , n57322 );
and ( n57439 , n57437 , n57438 );
xor ( n57440 , n57437 , n57438 );
xor ( n57441 , n56950 , n57260 );
and ( n57442 , n30154 , n57322 );
and ( n57443 , n57441 , n57442 );
xor ( n57444 , n57441 , n57442 );
xor ( n57445 , n56954 , n57258 );
and ( n57446 , n30159 , n57322 );
and ( n57447 , n57445 , n57446 );
xor ( n57448 , n57445 , n57446 );
xor ( n57449 , n56958 , n57256 );
and ( n57450 , n30164 , n57322 );
and ( n57451 , n57449 , n57450 );
xor ( n57452 , n57449 , n57450 );
xor ( n57453 , n56962 , n57254 );
and ( n57454 , n30169 , n57322 );
and ( n57455 , n57453 , n57454 );
xor ( n57456 , n57453 , n57454 );
xor ( n57457 , n56966 , n57252 );
and ( n57458 , n30174 , n57322 );
and ( n57459 , n57457 , n57458 );
xor ( n57460 , n57457 , n57458 );
xor ( n57461 , n56970 , n57250 );
and ( n57462 , n30179 , n57322 );
and ( n57463 , n57461 , n57462 );
xor ( n57464 , n57461 , n57462 );
xor ( n57465 , n56974 , n57248 );
and ( n57466 , n30184 , n57322 );
and ( n57467 , n57465 , n57466 );
xor ( n57468 , n57465 , n57466 );
xor ( n57469 , n56978 , n57246 );
and ( n57470 , n30189 , n57322 );
and ( n57471 , n57469 , n57470 );
xor ( n57472 , n57469 , n57470 );
xor ( n57473 , n56982 , n57244 );
and ( n57474 , n30194 , n57322 );
and ( n57475 , n57473 , n57474 );
xor ( n57476 , n57473 , n57474 );
xor ( n57477 , n56986 , n57242 );
and ( n57478 , n30199 , n57322 );
and ( n57479 , n57477 , n57478 );
xor ( n57480 , n57477 , n57478 );
xor ( n57481 , n56990 , n57240 );
and ( n57482 , n30204 , n57322 );
and ( n57483 , n57481 , n57482 );
xor ( n57484 , n57481 , n57482 );
xor ( n57485 , n56994 , n57238 );
and ( n57486 , n30209 , n57322 );
and ( n57487 , n57485 , n57486 );
xor ( n57488 , n57485 , n57486 );
xor ( n57489 , n56998 , n57236 );
and ( n57490 , n30214 , n57322 );
and ( n57491 , n57489 , n57490 );
xor ( n57492 , n57489 , n57490 );
xor ( n57493 , n57002 , n57234 );
and ( n57494 , n30219 , n57322 );
and ( n57495 , n57493 , n57494 );
xor ( n57496 , n57493 , n57494 );
xor ( n57497 , n57006 , n57232 );
and ( n57498 , n30224 , n57322 );
and ( n57499 , n57497 , n57498 );
xor ( n57500 , n57497 , n57498 );
xor ( n57501 , n57010 , n57230 );
and ( n57502 , n30229 , n57322 );
and ( n57503 , n57501 , n57502 );
xor ( n57504 , n57501 , n57502 );
xor ( n57505 , n57014 , n57228 );
and ( n57506 , n30234 , n57322 );
and ( n57507 , n57505 , n57506 );
xor ( n57508 , n57505 , n57506 );
xor ( n57509 , n57018 , n57226 );
and ( n57510 , n30239 , n57322 );
and ( n57511 , n57509 , n57510 );
xor ( n57512 , n57509 , n57510 );
xor ( n57513 , n57022 , n57224 );
and ( n57514 , n30244 , n57322 );
and ( n57515 , n57513 , n57514 );
xor ( n57516 , n57513 , n57514 );
xor ( n57517 , n57026 , n57222 );
and ( n57518 , n30249 , n57322 );
and ( n57519 , n57517 , n57518 );
xor ( n57520 , n57517 , n57518 );
xor ( n57521 , n57030 , n57220 );
and ( n57522 , n30254 , n57322 );
and ( n57523 , n57521 , n57522 );
xor ( n57524 , n57521 , n57522 );
xor ( n57525 , n57034 , n57218 );
and ( n57526 , n30259 , n57322 );
and ( n57527 , n57525 , n57526 );
xor ( n57528 , n57525 , n57526 );
xor ( n57529 , n57038 , n57216 );
and ( n57530 , n30264 , n57322 );
and ( n57531 , n57529 , n57530 );
xor ( n57532 , n57529 , n57530 );
xor ( n57533 , n57042 , n57214 );
and ( n57534 , n30269 , n57322 );
and ( n57535 , n57533 , n57534 );
xor ( n57536 , n57533 , n57534 );
xor ( n57537 , n57046 , n57212 );
and ( n57538 , n30274 , n57322 );
and ( n57539 , n57537 , n57538 );
xor ( n57540 , n57537 , n57538 );
xor ( n57541 , n57050 , n57210 );
and ( n57542 , n30279 , n57322 );
and ( n57543 , n57541 , n57542 );
xor ( n57544 , n57541 , n57542 );
xor ( n57545 , n57054 , n57208 );
and ( n57546 , n30284 , n57322 );
and ( n57547 , n57545 , n57546 );
xor ( n57548 , n57545 , n57546 );
xor ( n57549 , n57058 , n57206 );
and ( n57550 , n30289 , n57322 );
and ( n57551 , n57549 , n57550 );
xor ( n57552 , n57549 , n57550 );
xor ( n57553 , n57062 , n57204 );
and ( n57554 , n30294 , n57322 );
and ( n57555 , n57553 , n57554 );
xor ( n57556 , n57553 , n57554 );
xor ( n57557 , n57066 , n57202 );
and ( n57558 , n30299 , n57322 );
and ( n57559 , n57557 , n57558 );
xor ( n57560 , n57557 , n57558 );
xor ( n57561 , n57070 , n57200 );
and ( n57562 , n30304 , n57322 );
and ( n57563 , n57561 , n57562 );
xor ( n57564 , n57561 , n57562 );
xor ( n57565 , n57074 , n57198 );
and ( n57566 , n30309 , n57322 );
and ( n57567 , n57565 , n57566 );
xor ( n57568 , n57565 , n57566 );
xor ( n57569 , n57078 , n57196 );
and ( n57570 , n30314 , n57322 );
and ( n57571 , n57569 , n57570 );
xor ( n57572 , n57569 , n57570 );
xor ( n57573 , n57082 , n57194 );
and ( n57574 , n30319 , n57322 );
and ( n57575 , n57573 , n57574 );
xor ( n57576 , n57573 , n57574 );
xor ( n57577 , n57086 , n57192 );
and ( n57578 , n30324 , n57322 );
and ( n57579 , n57577 , n57578 );
xor ( n57580 , n57577 , n57578 );
xor ( n57581 , n57090 , n57190 );
and ( n57582 , n30329 , n57322 );
and ( n57583 , n57581 , n57582 );
xor ( n57584 , n57581 , n57582 );
xor ( n57585 , n57094 , n57188 );
and ( n57586 , n30334 , n57322 );
and ( n57587 , n57585 , n57586 );
xor ( n57588 , n57585 , n57586 );
xor ( n57589 , n57098 , n57186 );
and ( n57590 , n30339 , n57322 );
and ( n57591 , n57589 , n57590 );
xor ( n57592 , n57589 , n57590 );
xor ( n57593 , n57102 , n57184 );
and ( n57594 , n30344 , n57322 );
and ( n57595 , n57593 , n57594 );
xor ( n57596 , n57593 , n57594 );
xor ( n57597 , n57106 , n57182 );
and ( n57598 , n30349 , n57322 );
and ( n57599 , n57597 , n57598 );
xor ( n57600 , n57597 , n57598 );
xor ( n57601 , n57110 , n57180 );
and ( n57602 , n30354 , n57322 );
and ( n57603 , n57601 , n57602 );
xor ( n57604 , n57601 , n57602 );
xor ( n57605 , n57114 , n57178 );
and ( n57606 , n30359 , n57322 );
and ( n57607 , n57605 , n57606 );
xor ( n57608 , n57605 , n57606 );
xor ( n57609 , n57118 , n57176 );
and ( n57610 , n30364 , n57322 );
and ( n57611 , n57609 , n57610 );
xor ( n57612 , n57609 , n57610 );
xor ( n57613 , n57122 , n57174 );
and ( n57614 , n30369 , n57322 );
and ( n57615 , n57613 , n57614 );
xor ( n57616 , n57613 , n57614 );
xor ( n57617 , n57126 , n57172 );
and ( n57618 , n30374 , n57322 );
and ( n57619 , n57617 , n57618 );
xor ( n57620 , n57617 , n57618 );
xor ( n57621 , n57130 , n57170 );
and ( n57622 , n30379 , n57322 );
and ( n57623 , n57621 , n57622 );
xor ( n57624 , n57621 , n57622 );
xor ( n57625 , n57134 , n57168 );
and ( n57626 , n30384 , n57322 );
and ( n57627 , n57625 , n57626 );
xor ( n57628 , n57625 , n57626 );
xor ( n57629 , n57138 , n57166 );
and ( n57630 , n30389 , n57322 );
and ( n57631 , n57629 , n57630 );
xor ( n57632 , n57629 , n57630 );
xor ( n57633 , n57142 , n57164 );
and ( n57634 , n30394 , n57322 );
and ( n57635 , n57633 , n57634 );
xor ( n57636 , n57633 , n57634 );
xor ( n57637 , n57146 , n57162 );
and ( n57638 , n30399 , n57322 );
and ( n57639 , n57637 , n57638 );
xor ( n57640 , n57637 , n57638 );
xor ( n57641 , n57150 , n57160 );
and ( n57642 , n30404 , n57322 );
and ( n57643 , n57641 , n57642 );
xor ( n57644 , n57641 , n57642 );
xor ( n57645 , n57154 , n57158 );
and ( n57646 , n30409 , n57322 );
and ( n57647 , n57645 , n57646 );
buf ( n57648 , n57647 );
and ( n57649 , n57644 , n57648 );
or ( n57650 , n57643 , n57649 );
and ( n57651 , n57640 , n57650 );
or ( n57652 , n57639 , n57651 );
and ( n57653 , n57636 , n57652 );
or ( n57654 , n57635 , n57653 );
and ( n57655 , n57632 , n57654 );
or ( n57656 , n57631 , n57655 );
and ( n57657 , n57628 , n57656 );
or ( n57658 , n57627 , n57657 );
and ( n57659 , n57624 , n57658 );
or ( n57660 , n57623 , n57659 );
and ( n57661 , n57620 , n57660 );
or ( n57662 , n57619 , n57661 );
and ( n57663 , n57616 , n57662 );
or ( n57664 , n57615 , n57663 );
and ( n57665 , n57612 , n57664 );
or ( n57666 , n57611 , n57665 );
and ( n57667 , n57608 , n57666 );
or ( n57668 , n57607 , n57667 );
and ( n57669 , n57604 , n57668 );
or ( n57670 , n57603 , n57669 );
and ( n57671 , n57600 , n57670 );
or ( n57672 , n57599 , n57671 );
and ( n57673 , n57596 , n57672 );
or ( n57674 , n57595 , n57673 );
and ( n57675 , n57592 , n57674 );
or ( n57676 , n57591 , n57675 );
and ( n57677 , n57588 , n57676 );
or ( n57678 , n57587 , n57677 );
and ( n57679 , n57584 , n57678 );
or ( n57680 , n57583 , n57679 );
and ( n57681 , n57580 , n57680 );
or ( n57682 , n57579 , n57681 );
and ( n57683 , n57576 , n57682 );
or ( n57684 , n57575 , n57683 );
and ( n57685 , n57572 , n57684 );
or ( n57686 , n57571 , n57685 );
and ( n57687 , n57568 , n57686 );
or ( n57688 , n57567 , n57687 );
and ( n57689 , n57564 , n57688 );
or ( n57690 , n57563 , n57689 );
and ( n57691 , n57560 , n57690 );
or ( n57692 , n57559 , n57691 );
and ( n57693 , n57556 , n57692 );
or ( n57694 , n57555 , n57693 );
and ( n57695 , n57552 , n57694 );
or ( n57696 , n57551 , n57695 );
and ( n57697 , n57548 , n57696 );
or ( n57698 , n57547 , n57697 );
and ( n57699 , n57544 , n57698 );
or ( n57700 , n57543 , n57699 );
and ( n57701 , n57540 , n57700 );
or ( n57702 , n57539 , n57701 );
and ( n57703 , n57536 , n57702 );
or ( n57704 , n57535 , n57703 );
and ( n57705 , n57532 , n57704 );
or ( n57706 , n57531 , n57705 );
and ( n57707 , n57528 , n57706 );
or ( n57708 , n57527 , n57707 );
and ( n57709 , n57524 , n57708 );
or ( n57710 , n57523 , n57709 );
and ( n57711 , n57520 , n57710 );
or ( n57712 , n57519 , n57711 );
and ( n57713 , n57516 , n57712 );
or ( n57714 , n57515 , n57713 );
and ( n57715 , n57512 , n57714 );
or ( n57716 , n57511 , n57715 );
and ( n57717 , n57508 , n57716 );
or ( n57718 , n57507 , n57717 );
and ( n57719 , n57504 , n57718 );
or ( n57720 , n57503 , n57719 );
and ( n57721 , n57500 , n57720 );
or ( n57722 , n57499 , n57721 );
and ( n57723 , n57496 , n57722 );
or ( n57724 , n57495 , n57723 );
and ( n57725 , n57492 , n57724 );
or ( n57726 , n57491 , n57725 );
and ( n57727 , n57488 , n57726 );
or ( n57728 , n57487 , n57727 );
and ( n57729 , n57484 , n57728 );
or ( n57730 , n57483 , n57729 );
and ( n57731 , n57480 , n57730 );
or ( n57732 , n57479 , n57731 );
and ( n57733 , n57476 , n57732 );
or ( n57734 , n57475 , n57733 );
and ( n57735 , n57472 , n57734 );
or ( n57736 , n57471 , n57735 );
and ( n57737 , n57468 , n57736 );
or ( n57738 , n57467 , n57737 );
and ( n57739 , n57464 , n57738 );
or ( n57740 , n57463 , n57739 );
and ( n57741 , n57460 , n57740 );
or ( n57742 , n57459 , n57741 );
and ( n57743 , n57456 , n57742 );
or ( n57744 , n57455 , n57743 );
and ( n57745 , n57452 , n57744 );
or ( n57746 , n57451 , n57745 );
and ( n57747 , n57448 , n57746 );
or ( n57748 , n57447 , n57747 );
and ( n57749 , n57444 , n57748 );
or ( n57750 , n57443 , n57749 );
and ( n57751 , n57440 , n57750 );
or ( n57752 , n57439 , n57751 );
and ( n57753 , n57436 , n57752 );
or ( n57754 , n57435 , n57753 );
and ( n57755 , n57432 , n57754 );
or ( n57756 , n57431 , n57755 );
and ( n57757 , n57428 , n57756 );
or ( n57758 , n57427 , n57757 );
and ( n57759 , n57424 , n57758 );
or ( n57760 , n57423 , n57759 );
and ( n57761 , n57420 , n57760 );
or ( n57762 , n57419 , n57761 );
and ( n57763 , n57416 , n57762 );
or ( n57764 , n57415 , n57763 );
and ( n57765 , n57412 , n57764 );
or ( n57766 , n57411 , n57765 );
and ( n57767 , n57408 , n57766 );
or ( n57768 , n57407 , n57767 );
and ( n57769 , n57404 , n57768 );
or ( n57770 , n57403 , n57769 );
and ( n57771 , n57400 , n57770 );
or ( n57772 , n57399 , n57771 );
and ( n57773 , n57396 , n57772 );
or ( n57774 , n57395 , n57773 );
and ( n57775 , n57392 , n57774 );
or ( n57776 , n57391 , n57775 );
and ( n57777 , n57388 , n57776 );
or ( n57778 , n57387 , n57777 );
and ( n57779 , n57384 , n57778 );
or ( n57780 , n57383 , n57779 );
and ( n57781 , n57380 , n57780 );
or ( n57782 , n57379 , n57781 );
and ( n57783 , n57376 , n57782 );
or ( n57784 , n57375 , n57783 );
and ( n57785 , n57372 , n57784 );
or ( n57786 , n57371 , n57785 );
and ( n57787 , n57368 , n57786 );
or ( n57788 , n57367 , n57787 );
and ( n57789 , n57364 , n57788 );
or ( n57790 , n57363 , n57789 );
and ( n57791 , n57360 , n57790 );
or ( n57792 , n57359 , n57791 );
and ( n57793 , n57356 , n57792 );
or ( n57794 , n57355 , n57793 );
and ( n57795 , n57352 , n57794 );
or ( n57796 , n57351 , n57795 );
and ( n57797 , n57348 , n57796 );
or ( n57798 , n57347 , n57797 );
and ( n57799 , n57344 , n57798 );
or ( n57800 , n57343 , n57799 );
and ( n57801 , n57340 , n57800 );
or ( n57802 , n57339 , n57801 );
and ( n57803 , n57336 , n57802 );
or ( n57804 , n57335 , n57803 );
and ( n57805 , n57332 , n57804 );
or ( n57806 , n57331 , n57805 );
and ( n57807 , n57328 , n57806 );
or ( n57808 , n57327 , n57807 );
xor ( n57809 , n57324 , n57808 );
buf ( n57810 , n18014 );
and ( n57811 , n30009 , n57810 );
xor ( n57812 , n57809 , n57811 );
xor ( n57813 , n57328 , n57806 );
and ( n57814 , n30014 , n57810 );
and ( n57815 , n57813 , n57814 );
xor ( n57816 , n57813 , n57814 );
xor ( n57817 , n57332 , n57804 );
and ( n57818 , n30019 , n57810 );
and ( n57819 , n57817 , n57818 );
xor ( n57820 , n57817 , n57818 );
xor ( n57821 , n57336 , n57802 );
and ( n57822 , n30024 , n57810 );
and ( n57823 , n57821 , n57822 );
xor ( n57824 , n57821 , n57822 );
xor ( n57825 , n57340 , n57800 );
and ( n57826 , n30029 , n57810 );
and ( n57827 , n57825 , n57826 );
xor ( n57828 , n57825 , n57826 );
xor ( n57829 , n57344 , n57798 );
and ( n57830 , n30034 , n57810 );
and ( n57831 , n57829 , n57830 );
xor ( n57832 , n57829 , n57830 );
xor ( n57833 , n57348 , n57796 );
and ( n57834 , n30039 , n57810 );
and ( n57835 , n57833 , n57834 );
xor ( n57836 , n57833 , n57834 );
xor ( n57837 , n57352 , n57794 );
and ( n57838 , n30044 , n57810 );
and ( n57839 , n57837 , n57838 );
xor ( n57840 , n57837 , n57838 );
xor ( n57841 , n57356 , n57792 );
and ( n57842 , n30049 , n57810 );
and ( n57843 , n57841 , n57842 );
xor ( n57844 , n57841 , n57842 );
xor ( n57845 , n57360 , n57790 );
and ( n57846 , n30054 , n57810 );
and ( n57847 , n57845 , n57846 );
xor ( n57848 , n57845 , n57846 );
xor ( n57849 , n57364 , n57788 );
and ( n57850 , n30059 , n57810 );
and ( n57851 , n57849 , n57850 );
xor ( n57852 , n57849 , n57850 );
xor ( n57853 , n57368 , n57786 );
and ( n57854 , n30064 , n57810 );
and ( n57855 , n57853 , n57854 );
xor ( n57856 , n57853 , n57854 );
xor ( n57857 , n57372 , n57784 );
and ( n57858 , n30069 , n57810 );
and ( n57859 , n57857 , n57858 );
xor ( n57860 , n57857 , n57858 );
xor ( n57861 , n57376 , n57782 );
and ( n57862 , n30074 , n57810 );
and ( n57863 , n57861 , n57862 );
xor ( n57864 , n57861 , n57862 );
xor ( n57865 , n57380 , n57780 );
and ( n57866 , n30079 , n57810 );
and ( n57867 , n57865 , n57866 );
xor ( n57868 , n57865 , n57866 );
xor ( n57869 , n57384 , n57778 );
and ( n57870 , n30084 , n57810 );
and ( n57871 , n57869 , n57870 );
xor ( n57872 , n57869 , n57870 );
xor ( n57873 , n57388 , n57776 );
and ( n57874 , n30089 , n57810 );
and ( n57875 , n57873 , n57874 );
xor ( n57876 , n57873 , n57874 );
xor ( n57877 , n57392 , n57774 );
and ( n57878 , n30094 , n57810 );
and ( n57879 , n57877 , n57878 );
xor ( n57880 , n57877 , n57878 );
xor ( n57881 , n57396 , n57772 );
and ( n57882 , n30099 , n57810 );
and ( n57883 , n57881 , n57882 );
xor ( n57884 , n57881 , n57882 );
xor ( n57885 , n57400 , n57770 );
and ( n57886 , n30104 , n57810 );
and ( n57887 , n57885 , n57886 );
xor ( n57888 , n57885 , n57886 );
xor ( n57889 , n57404 , n57768 );
and ( n57890 , n30109 , n57810 );
and ( n57891 , n57889 , n57890 );
xor ( n57892 , n57889 , n57890 );
xor ( n57893 , n57408 , n57766 );
and ( n57894 , n30114 , n57810 );
and ( n57895 , n57893 , n57894 );
xor ( n57896 , n57893 , n57894 );
xor ( n57897 , n57412 , n57764 );
and ( n57898 , n30119 , n57810 );
and ( n57899 , n57897 , n57898 );
xor ( n57900 , n57897 , n57898 );
xor ( n57901 , n57416 , n57762 );
and ( n57902 , n30124 , n57810 );
and ( n57903 , n57901 , n57902 );
xor ( n57904 , n57901 , n57902 );
xor ( n57905 , n57420 , n57760 );
and ( n57906 , n30129 , n57810 );
and ( n57907 , n57905 , n57906 );
xor ( n57908 , n57905 , n57906 );
xor ( n57909 , n57424 , n57758 );
and ( n57910 , n30134 , n57810 );
and ( n57911 , n57909 , n57910 );
xor ( n57912 , n57909 , n57910 );
xor ( n57913 , n57428 , n57756 );
and ( n57914 , n30139 , n57810 );
and ( n57915 , n57913 , n57914 );
xor ( n57916 , n57913 , n57914 );
xor ( n57917 , n57432 , n57754 );
and ( n57918 , n30144 , n57810 );
and ( n57919 , n57917 , n57918 );
xor ( n57920 , n57917 , n57918 );
xor ( n57921 , n57436 , n57752 );
and ( n57922 , n30149 , n57810 );
and ( n57923 , n57921 , n57922 );
xor ( n57924 , n57921 , n57922 );
xor ( n57925 , n57440 , n57750 );
and ( n57926 , n30154 , n57810 );
and ( n57927 , n57925 , n57926 );
xor ( n57928 , n57925 , n57926 );
xor ( n57929 , n57444 , n57748 );
and ( n57930 , n30159 , n57810 );
and ( n57931 , n57929 , n57930 );
xor ( n57932 , n57929 , n57930 );
xor ( n57933 , n57448 , n57746 );
and ( n57934 , n30164 , n57810 );
and ( n57935 , n57933 , n57934 );
xor ( n57936 , n57933 , n57934 );
xor ( n57937 , n57452 , n57744 );
and ( n57938 , n30169 , n57810 );
and ( n57939 , n57937 , n57938 );
xor ( n57940 , n57937 , n57938 );
xor ( n57941 , n57456 , n57742 );
and ( n57942 , n30174 , n57810 );
and ( n57943 , n57941 , n57942 );
xor ( n57944 , n57941 , n57942 );
xor ( n57945 , n57460 , n57740 );
and ( n57946 , n30179 , n57810 );
and ( n57947 , n57945 , n57946 );
xor ( n57948 , n57945 , n57946 );
xor ( n57949 , n57464 , n57738 );
and ( n57950 , n30184 , n57810 );
and ( n57951 , n57949 , n57950 );
xor ( n57952 , n57949 , n57950 );
xor ( n57953 , n57468 , n57736 );
and ( n57954 , n30189 , n57810 );
and ( n57955 , n57953 , n57954 );
xor ( n57956 , n57953 , n57954 );
xor ( n57957 , n57472 , n57734 );
and ( n57958 , n30194 , n57810 );
and ( n57959 , n57957 , n57958 );
xor ( n57960 , n57957 , n57958 );
xor ( n57961 , n57476 , n57732 );
and ( n57962 , n30199 , n57810 );
and ( n57963 , n57961 , n57962 );
xor ( n57964 , n57961 , n57962 );
xor ( n57965 , n57480 , n57730 );
and ( n57966 , n30204 , n57810 );
and ( n57967 , n57965 , n57966 );
xor ( n57968 , n57965 , n57966 );
xor ( n57969 , n57484 , n57728 );
and ( n57970 , n30209 , n57810 );
and ( n57971 , n57969 , n57970 );
xor ( n57972 , n57969 , n57970 );
xor ( n57973 , n57488 , n57726 );
and ( n57974 , n30214 , n57810 );
and ( n57975 , n57973 , n57974 );
xor ( n57976 , n57973 , n57974 );
xor ( n57977 , n57492 , n57724 );
and ( n57978 , n30219 , n57810 );
and ( n57979 , n57977 , n57978 );
xor ( n57980 , n57977 , n57978 );
xor ( n57981 , n57496 , n57722 );
and ( n57982 , n30224 , n57810 );
and ( n57983 , n57981 , n57982 );
xor ( n57984 , n57981 , n57982 );
xor ( n57985 , n57500 , n57720 );
and ( n57986 , n30229 , n57810 );
and ( n57987 , n57985 , n57986 );
xor ( n57988 , n57985 , n57986 );
xor ( n57989 , n57504 , n57718 );
and ( n57990 , n30234 , n57810 );
and ( n57991 , n57989 , n57990 );
xor ( n57992 , n57989 , n57990 );
xor ( n57993 , n57508 , n57716 );
and ( n57994 , n30239 , n57810 );
and ( n57995 , n57993 , n57994 );
xor ( n57996 , n57993 , n57994 );
xor ( n57997 , n57512 , n57714 );
and ( n57998 , n30244 , n57810 );
and ( n57999 , n57997 , n57998 );
xor ( n58000 , n57997 , n57998 );
xor ( n58001 , n57516 , n57712 );
and ( n58002 , n30249 , n57810 );
and ( n58003 , n58001 , n58002 );
xor ( n58004 , n58001 , n58002 );
xor ( n58005 , n57520 , n57710 );
and ( n58006 , n30254 , n57810 );
and ( n58007 , n58005 , n58006 );
xor ( n58008 , n58005 , n58006 );
xor ( n58009 , n57524 , n57708 );
and ( n58010 , n30259 , n57810 );
and ( n58011 , n58009 , n58010 );
xor ( n58012 , n58009 , n58010 );
xor ( n58013 , n57528 , n57706 );
and ( n58014 , n30264 , n57810 );
and ( n58015 , n58013 , n58014 );
xor ( n58016 , n58013 , n58014 );
xor ( n58017 , n57532 , n57704 );
and ( n58018 , n30269 , n57810 );
and ( n58019 , n58017 , n58018 );
xor ( n58020 , n58017 , n58018 );
xor ( n58021 , n57536 , n57702 );
and ( n58022 , n30274 , n57810 );
and ( n58023 , n58021 , n58022 );
xor ( n58024 , n58021 , n58022 );
xor ( n58025 , n57540 , n57700 );
and ( n58026 , n30279 , n57810 );
and ( n58027 , n58025 , n58026 );
xor ( n58028 , n58025 , n58026 );
xor ( n58029 , n57544 , n57698 );
and ( n58030 , n30284 , n57810 );
and ( n58031 , n58029 , n58030 );
xor ( n58032 , n58029 , n58030 );
xor ( n58033 , n57548 , n57696 );
and ( n58034 , n30289 , n57810 );
and ( n58035 , n58033 , n58034 );
xor ( n58036 , n58033 , n58034 );
xor ( n58037 , n57552 , n57694 );
and ( n58038 , n30294 , n57810 );
and ( n58039 , n58037 , n58038 );
xor ( n58040 , n58037 , n58038 );
xor ( n58041 , n57556 , n57692 );
and ( n58042 , n30299 , n57810 );
and ( n58043 , n58041 , n58042 );
xor ( n58044 , n58041 , n58042 );
xor ( n58045 , n57560 , n57690 );
and ( n58046 , n30304 , n57810 );
and ( n58047 , n58045 , n58046 );
xor ( n58048 , n58045 , n58046 );
xor ( n58049 , n57564 , n57688 );
and ( n58050 , n30309 , n57810 );
and ( n58051 , n58049 , n58050 );
xor ( n58052 , n58049 , n58050 );
xor ( n58053 , n57568 , n57686 );
and ( n58054 , n30314 , n57810 );
and ( n58055 , n58053 , n58054 );
xor ( n58056 , n58053 , n58054 );
xor ( n58057 , n57572 , n57684 );
and ( n58058 , n30319 , n57810 );
and ( n58059 , n58057 , n58058 );
xor ( n58060 , n58057 , n58058 );
xor ( n58061 , n57576 , n57682 );
and ( n58062 , n30324 , n57810 );
and ( n58063 , n58061 , n58062 );
xor ( n58064 , n58061 , n58062 );
xor ( n58065 , n57580 , n57680 );
and ( n58066 , n30329 , n57810 );
and ( n58067 , n58065 , n58066 );
xor ( n58068 , n58065 , n58066 );
xor ( n58069 , n57584 , n57678 );
and ( n58070 , n30334 , n57810 );
and ( n58071 , n58069 , n58070 );
xor ( n58072 , n58069 , n58070 );
xor ( n58073 , n57588 , n57676 );
and ( n58074 , n30339 , n57810 );
and ( n58075 , n58073 , n58074 );
xor ( n58076 , n58073 , n58074 );
xor ( n58077 , n57592 , n57674 );
and ( n58078 , n30344 , n57810 );
and ( n58079 , n58077 , n58078 );
xor ( n58080 , n58077 , n58078 );
xor ( n58081 , n57596 , n57672 );
and ( n58082 , n30349 , n57810 );
and ( n58083 , n58081 , n58082 );
xor ( n58084 , n58081 , n58082 );
xor ( n58085 , n57600 , n57670 );
and ( n58086 , n30354 , n57810 );
and ( n58087 , n58085 , n58086 );
xor ( n58088 , n58085 , n58086 );
xor ( n58089 , n57604 , n57668 );
and ( n58090 , n30359 , n57810 );
and ( n58091 , n58089 , n58090 );
xor ( n58092 , n58089 , n58090 );
xor ( n58093 , n57608 , n57666 );
and ( n58094 , n30364 , n57810 );
and ( n58095 , n58093 , n58094 );
xor ( n58096 , n58093 , n58094 );
xor ( n58097 , n57612 , n57664 );
and ( n58098 , n30369 , n57810 );
and ( n58099 , n58097 , n58098 );
xor ( n58100 , n58097 , n58098 );
xor ( n58101 , n57616 , n57662 );
and ( n58102 , n30374 , n57810 );
and ( n58103 , n58101 , n58102 );
xor ( n58104 , n58101 , n58102 );
xor ( n58105 , n57620 , n57660 );
and ( n58106 , n30379 , n57810 );
and ( n58107 , n58105 , n58106 );
xor ( n58108 , n58105 , n58106 );
xor ( n58109 , n57624 , n57658 );
and ( n58110 , n30384 , n57810 );
and ( n58111 , n58109 , n58110 );
xor ( n58112 , n58109 , n58110 );
xor ( n58113 , n57628 , n57656 );
and ( n58114 , n30389 , n57810 );
and ( n58115 , n58113 , n58114 );
xor ( n58116 , n58113 , n58114 );
xor ( n58117 , n57632 , n57654 );
and ( n58118 , n30394 , n57810 );
and ( n58119 , n58117 , n58118 );
xor ( n58120 , n58117 , n58118 );
xor ( n58121 , n57636 , n57652 );
and ( n58122 , n30399 , n57810 );
and ( n58123 , n58121 , n58122 );
xor ( n58124 , n58121 , n58122 );
xor ( n58125 , n57640 , n57650 );
and ( n58126 , n30404 , n57810 );
and ( n58127 , n58125 , n58126 );
xor ( n58128 , n58125 , n58126 );
xor ( n58129 , n57644 , n57648 );
and ( n58130 , n30409 , n57810 );
and ( n58131 , n58129 , n58130 );
buf ( n58132 , n58131 );
and ( n58133 , n58128 , n58132 );
or ( n58134 , n58127 , n58133 );
and ( n58135 , n58124 , n58134 );
or ( n58136 , n58123 , n58135 );
and ( n58137 , n58120 , n58136 );
or ( n58138 , n58119 , n58137 );
and ( n58139 , n58116 , n58138 );
or ( n58140 , n58115 , n58139 );
and ( n58141 , n58112 , n58140 );
or ( n58142 , n58111 , n58141 );
and ( n58143 , n58108 , n58142 );
or ( n58144 , n58107 , n58143 );
and ( n58145 , n58104 , n58144 );
or ( n58146 , n58103 , n58145 );
and ( n58147 , n58100 , n58146 );
or ( n58148 , n58099 , n58147 );
and ( n58149 , n58096 , n58148 );
or ( n58150 , n58095 , n58149 );
and ( n58151 , n58092 , n58150 );
or ( n58152 , n58091 , n58151 );
and ( n58153 , n58088 , n58152 );
or ( n58154 , n58087 , n58153 );
and ( n58155 , n58084 , n58154 );
or ( n58156 , n58083 , n58155 );
and ( n58157 , n58080 , n58156 );
or ( n58158 , n58079 , n58157 );
and ( n58159 , n58076 , n58158 );
or ( n58160 , n58075 , n58159 );
and ( n58161 , n58072 , n58160 );
or ( n58162 , n58071 , n58161 );
and ( n58163 , n58068 , n58162 );
or ( n58164 , n58067 , n58163 );
and ( n58165 , n58064 , n58164 );
or ( n58166 , n58063 , n58165 );
and ( n58167 , n58060 , n58166 );
or ( n58168 , n58059 , n58167 );
and ( n58169 , n58056 , n58168 );
or ( n58170 , n58055 , n58169 );
and ( n58171 , n58052 , n58170 );
or ( n58172 , n58051 , n58171 );
and ( n58173 , n58048 , n58172 );
or ( n58174 , n58047 , n58173 );
and ( n58175 , n58044 , n58174 );
or ( n58176 , n58043 , n58175 );
and ( n58177 , n58040 , n58176 );
or ( n58178 , n58039 , n58177 );
and ( n58179 , n58036 , n58178 );
or ( n58180 , n58035 , n58179 );
and ( n58181 , n58032 , n58180 );
or ( n58182 , n58031 , n58181 );
and ( n58183 , n58028 , n58182 );
or ( n58184 , n58027 , n58183 );
and ( n58185 , n58024 , n58184 );
or ( n58186 , n58023 , n58185 );
and ( n58187 , n58020 , n58186 );
or ( n58188 , n58019 , n58187 );
and ( n58189 , n58016 , n58188 );
or ( n58190 , n58015 , n58189 );
and ( n58191 , n58012 , n58190 );
or ( n58192 , n58011 , n58191 );
and ( n58193 , n58008 , n58192 );
or ( n58194 , n58007 , n58193 );
and ( n58195 , n58004 , n58194 );
or ( n58196 , n58003 , n58195 );
and ( n58197 , n58000 , n58196 );
or ( n58198 , n57999 , n58197 );
and ( n58199 , n57996 , n58198 );
or ( n58200 , n57995 , n58199 );
and ( n58201 , n57992 , n58200 );
or ( n58202 , n57991 , n58201 );
and ( n58203 , n57988 , n58202 );
or ( n58204 , n57987 , n58203 );
and ( n58205 , n57984 , n58204 );
or ( n58206 , n57983 , n58205 );
and ( n58207 , n57980 , n58206 );
or ( n58208 , n57979 , n58207 );
and ( n58209 , n57976 , n58208 );
or ( n58210 , n57975 , n58209 );
and ( n58211 , n57972 , n58210 );
or ( n58212 , n57971 , n58211 );
and ( n58213 , n57968 , n58212 );
or ( n58214 , n57967 , n58213 );
and ( n58215 , n57964 , n58214 );
or ( n58216 , n57963 , n58215 );
and ( n58217 , n57960 , n58216 );
or ( n58218 , n57959 , n58217 );
and ( n58219 , n57956 , n58218 );
or ( n58220 , n57955 , n58219 );
and ( n58221 , n57952 , n58220 );
or ( n58222 , n57951 , n58221 );
and ( n58223 , n57948 , n58222 );
or ( n58224 , n57947 , n58223 );
and ( n58225 , n57944 , n58224 );
or ( n58226 , n57943 , n58225 );
and ( n58227 , n57940 , n58226 );
or ( n58228 , n57939 , n58227 );
and ( n58229 , n57936 , n58228 );
or ( n58230 , n57935 , n58229 );
and ( n58231 , n57932 , n58230 );
or ( n58232 , n57931 , n58231 );
and ( n58233 , n57928 , n58232 );
or ( n58234 , n57927 , n58233 );
and ( n58235 , n57924 , n58234 );
or ( n58236 , n57923 , n58235 );
and ( n58237 , n57920 , n58236 );
or ( n58238 , n57919 , n58237 );
and ( n58239 , n57916 , n58238 );
or ( n58240 , n57915 , n58239 );
and ( n58241 , n57912 , n58240 );
or ( n58242 , n57911 , n58241 );
and ( n58243 , n57908 , n58242 );
or ( n58244 , n57907 , n58243 );
and ( n58245 , n57904 , n58244 );
or ( n58246 , n57903 , n58245 );
and ( n58247 , n57900 , n58246 );
or ( n58248 , n57899 , n58247 );
and ( n58249 , n57896 , n58248 );
or ( n58250 , n57895 , n58249 );
and ( n58251 , n57892 , n58250 );
or ( n58252 , n57891 , n58251 );
and ( n58253 , n57888 , n58252 );
or ( n58254 , n57887 , n58253 );
and ( n58255 , n57884 , n58254 );
or ( n58256 , n57883 , n58255 );
and ( n58257 , n57880 , n58256 );
or ( n58258 , n57879 , n58257 );
and ( n58259 , n57876 , n58258 );
or ( n58260 , n57875 , n58259 );
and ( n58261 , n57872 , n58260 );
or ( n58262 , n57871 , n58261 );
and ( n58263 , n57868 , n58262 );
or ( n58264 , n57867 , n58263 );
and ( n58265 , n57864 , n58264 );
or ( n58266 , n57863 , n58265 );
and ( n58267 , n57860 , n58266 );
or ( n58268 , n57859 , n58267 );
and ( n58269 , n57856 , n58268 );
or ( n58270 , n57855 , n58269 );
and ( n58271 , n57852 , n58270 );
or ( n58272 , n57851 , n58271 );
and ( n58273 , n57848 , n58272 );
or ( n58274 , n57847 , n58273 );
and ( n58275 , n57844 , n58274 );
or ( n58276 , n57843 , n58275 );
and ( n58277 , n57840 , n58276 );
or ( n58278 , n57839 , n58277 );
and ( n58279 , n57836 , n58278 );
or ( n58280 , n57835 , n58279 );
and ( n58281 , n57832 , n58280 );
or ( n58282 , n57831 , n58281 );
and ( n58283 , n57828 , n58282 );
or ( n58284 , n57827 , n58283 );
and ( n58285 , n57824 , n58284 );
or ( n58286 , n57823 , n58285 );
and ( n58287 , n57820 , n58286 );
or ( n58288 , n57819 , n58287 );
and ( n58289 , n57816 , n58288 );
or ( n58290 , n57815 , n58289 );
xor ( n58291 , n57812 , n58290 );
buf ( n58292 , n18012 );
and ( n58293 , n30014 , n58292 );
xor ( n58294 , n58291 , n58293 );
xor ( n58295 , n57816 , n58288 );
and ( n58296 , n30019 , n58292 );
and ( n58297 , n58295 , n58296 );
xor ( n58298 , n58295 , n58296 );
xor ( n58299 , n57820 , n58286 );
and ( n58300 , n30024 , n58292 );
and ( n58301 , n58299 , n58300 );
xor ( n58302 , n58299 , n58300 );
xor ( n58303 , n57824 , n58284 );
and ( n58304 , n30029 , n58292 );
and ( n58305 , n58303 , n58304 );
xor ( n58306 , n58303 , n58304 );
xor ( n58307 , n57828 , n58282 );
and ( n58308 , n30034 , n58292 );
and ( n58309 , n58307 , n58308 );
xor ( n58310 , n58307 , n58308 );
xor ( n58311 , n57832 , n58280 );
and ( n58312 , n30039 , n58292 );
and ( n58313 , n58311 , n58312 );
xor ( n58314 , n58311 , n58312 );
xor ( n58315 , n57836 , n58278 );
and ( n58316 , n30044 , n58292 );
and ( n58317 , n58315 , n58316 );
xor ( n58318 , n58315 , n58316 );
xor ( n58319 , n57840 , n58276 );
and ( n58320 , n30049 , n58292 );
and ( n58321 , n58319 , n58320 );
xor ( n58322 , n58319 , n58320 );
xor ( n58323 , n57844 , n58274 );
and ( n58324 , n30054 , n58292 );
and ( n58325 , n58323 , n58324 );
xor ( n58326 , n58323 , n58324 );
xor ( n58327 , n57848 , n58272 );
and ( n58328 , n30059 , n58292 );
and ( n58329 , n58327 , n58328 );
xor ( n58330 , n58327 , n58328 );
xor ( n58331 , n57852 , n58270 );
and ( n58332 , n30064 , n58292 );
and ( n58333 , n58331 , n58332 );
xor ( n58334 , n58331 , n58332 );
xor ( n58335 , n57856 , n58268 );
and ( n58336 , n30069 , n58292 );
and ( n58337 , n58335 , n58336 );
xor ( n58338 , n58335 , n58336 );
xor ( n58339 , n57860 , n58266 );
and ( n58340 , n30074 , n58292 );
and ( n58341 , n58339 , n58340 );
xor ( n58342 , n58339 , n58340 );
xor ( n58343 , n57864 , n58264 );
and ( n58344 , n30079 , n58292 );
and ( n58345 , n58343 , n58344 );
xor ( n58346 , n58343 , n58344 );
xor ( n58347 , n57868 , n58262 );
and ( n58348 , n30084 , n58292 );
and ( n58349 , n58347 , n58348 );
xor ( n58350 , n58347 , n58348 );
xor ( n58351 , n57872 , n58260 );
and ( n58352 , n30089 , n58292 );
and ( n58353 , n58351 , n58352 );
xor ( n58354 , n58351 , n58352 );
xor ( n58355 , n57876 , n58258 );
and ( n58356 , n30094 , n58292 );
and ( n58357 , n58355 , n58356 );
xor ( n58358 , n58355 , n58356 );
xor ( n58359 , n57880 , n58256 );
and ( n58360 , n30099 , n58292 );
and ( n58361 , n58359 , n58360 );
xor ( n58362 , n58359 , n58360 );
xor ( n58363 , n57884 , n58254 );
and ( n58364 , n30104 , n58292 );
and ( n58365 , n58363 , n58364 );
xor ( n58366 , n58363 , n58364 );
xor ( n58367 , n57888 , n58252 );
and ( n58368 , n30109 , n58292 );
and ( n58369 , n58367 , n58368 );
xor ( n58370 , n58367 , n58368 );
xor ( n58371 , n57892 , n58250 );
and ( n58372 , n30114 , n58292 );
and ( n58373 , n58371 , n58372 );
xor ( n58374 , n58371 , n58372 );
xor ( n58375 , n57896 , n58248 );
and ( n58376 , n30119 , n58292 );
and ( n58377 , n58375 , n58376 );
xor ( n58378 , n58375 , n58376 );
xor ( n58379 , n57900 , n58246 );
and ( n58380 , n30124 , n58292 );
and ( n58381 , n58379 , n58380 );
xor ( n58382 , n58379 , n58380 );
xor ( n58383 , n57904 , n58244 );
and ( n58384 , n30129 , n58292 );
and ( n58385 , n58383 , n58384 );
xor ( n58386 , n58383 , n58384 );
xor ( n58387 , n57908 , n58242 );
and ( n58388 , n30134 , n58292 );
and ( n58389 , n58387 , n58388 );
xor ( n58390 , n58387 , n58388 );
xor ( n58391 , n57912 , n58240 );
and ( n58392 , n30139 , n58292 );
and ( n58393 , n58391 , n58392 );
xor ( n58394 , n58391 , n58392 );
xor ( n58395 , n57916 , n58238 );
and ( n58396 , n30144 , n58292 );
and ( n58397 , n58395 , n58396 );
xor ( n58398 , n58395 , n58396 );
xor ( n58399 , n57920 , n58236 );
and ( n58400 , n30149 , n58292 );
and ( n58401 , n58399 , n58400 );
xor ( n58402 , n58399 , n58400 );
xor ( n58403 , n57924 , n58234 );
and ( n58404 , n30154 , n58292 );
and ( n58405 , n58403 , n58404 );
xor ( n58406 , n58403 , n58404 );
xor ( n58407 , n57928 , n58232 );
and ( n58408 , n30159 , n58292 );
and ( n58409 , n58407 , n58408 );
xor ( n58410 , n58407 , n58408 );
xor ( n58411 , n57932 , n58230 );
and ( n58412 , n30164 , n58292 );
and ( n58413 , n58411 , n58412 );
xor ( n58414 , n58411 , n58412 );
xor ( n58415 , n57936 , n58228 );
and ( n58416 , n30169 , n58292 );
and ( n58417 , n58415 , n58416 );
xor ( n58418 , n58415 , n58416 );
xor ( n58419 , n57940 , n58226 );
and ( n58420 , n30174 , n58292 );
and ( n58421 , n58419 , n58420 );
xor ( n58422 , n58419 , n58420 );
xor ( n58423 , n57944 , n58224 );
and ( n58424 , n30179 , n58292 );
and ( n58425 , n58423 , n58424 );
xor ( n58426 , n58423 , n58424 );
xor ( n58427 , n57948 , n58222 );
and ( n58428 , n30184 , n58292 );
and ( n58429 , n58427 , n58428 );
xor ( n58430 , n58427 , n58428 );
xor ( n58431 , n57952 , n58220 );
and ( n58432 , n30189 , n58292 );
and ( n58433 , n58431 , n58432 );
xor ( n58434 , n58431 , n58432 );
xor ( n58435 , n57956 , n58218 );
and ( n58436 , n30194 , n58292 );
and ( n58437 , n58435 , n58436 );
xor ( n58438 , n58435 , n58436 );
xor ( n58439 , n57960 , n58216 );
and ( n58440 , n30199 , n58292 );
and ( n58441 , n58439 , n58440 );
xor ( n58442 , n58439 , n58440 );
xor ( n58443 , n57964 , n58214 );
and ( n58444 , n30204 , n58292 );
and ( n58445 , n58443 , n58444 );
xor ( n58446 , n58443 , n58444 );
xor ( n58447 , n57968 , n58212 );
and ( n58448 , n30209 , n58292 );
and ( n58449 , n58447 , n58448 );
xor ( n58450 , n58447 , n58448 );
xor ( n58451 , n57972 , n58210 );
and ( n58452 , n30214 , n58292 );
and ( n58453 , n58451 , n58452 );
xor ( n58454 , n58451 , n58452 );
xor ( n58455 , n57976 , n58208 );
and ( n58456 , n30219 , n58292 );
and ( n58457 , n58455 , n58456 );
xor ( n58458 , n58455 , n58456 );
xor ( n58459 , n57980 , n58206 );
and ( n58460 , n30224 , n58292 );
and ( n58461 , n58459 , n58460 );
xor ( n58462 , n58459 , n58460 );
xor ( n58463 , n57984 , n58204 );
and ( n58464 , n30229 , n58292 );
and ( n58465 , n58463 , n58464 );
xor ( n58466 , n58463 , n58464 );
xor ( n58467 , n57988 , n58202 );
and ( n58468 , n30234 , n58292 );
and ( n58469 , n58467 , n58468 );
xor ( n58470 , n58467 , n58468 );
xor ( n58471 , n57992 , n58200 );
and ( n58472 , n30239 , n58292 );
and ( n58473 , n58471 , n58472 );
xor ( n58474 , n58471 , n58472 );
xor ( n58475 , n57996 , n58198 );
and ( n58476 , n30244 , n58292 );
and ( n58477 , n58475 , n58476 );
xor ( n58478 , n58475 , n58476 );
xor ( n58479 , n58000 , n58196 );
and ( n58480 , n30249 , n58292 );
and ( n58481 , n58479 , n58480 );
xor ( n58482 , n58479 , n58480 );
xor ( n58483 , n58004 , n58194 );
and ( n58484 , n30254 , n58292 );
and ( n58485 , n58483 , n58484 );
xor ( n58486 , n58483 , n58484 );
xor ( n58487 , n58008 , n58192 );
and ( n58488 , n30259 , n58292 );
and ( n58489 , n58487 , n58488 );
xor ( n58490 , n58487 , n58488 );
xor ( n58491 , n58012 , n58190 );
and ( n58492 , n30264 , n58292 );
and ( n58493 , n58491 , n58492 );
xor ( n58494 , n58491 , n58492 );
xor ( n58495 , n58016 , n58188 );
and ( n58496 , n30269 , n58292 );
and ( n58497 , n58495 , n58496 );
xor ( n58498 , n58495 , n58496 );
xor ( n58499 , n58020 , n58186 );
and ( n58500 , n30274 , n58292 );
and ( n58501 , n58499 , n58500 );
xor ( n58502 , n58499 , n58500 );
xor ( n58503 , n58024 , n58184 );
and ( n58504 , n30279 , n58292 );
and ( n58505 , n58503 , n58504 );
xor ( n58506 , n58503 , n58504 );
xor ( n58507 , n58028 , n58182 );
and ( n58508 , n30284 , n58292 );
and ( n58509 , n58507 , n58508 );
xor ( n58510 , n58507 , n58508 );
xor ( n58511 , n58032 , n58180 );
and ( n58512 , n30289 , n58292 );
and ( n58513 , n58511 , n58512 );
xor ( n58514 , n58511 , n58512 );
xor ( n58515 , n58036 , n58178 );
and ( n58516 , n30294 , n58292 );
and ( n58517 , n58515 , n58516 );
xor ( n58518 , n58515 , n58516 );
xor ( n58519 , n58040 , n58176 );
and ( n58520 , n30299 , n58292 );
and ( n58521 , n58519 , n58520 );
xor ( n58522 , n58519 , n58520 );
xor ( n58523 , n58044 , n58174 );
and ( n58524 , n30304 , n58292 );
and ( n58525 , n58523 , n58524 );
xor ( n58526 , n58523 , n58524 );
xor ( n58527 , n58048 , n58172 );
and ( n58528 , n30309 , n58292 );
and ( n58529 , n58527 , n58528 );
xor ( n58530 , n58527 , n58528 );
xor ( n58531 , n58052 , n58170 );
and ( n58532 , n30314 , n58292 );
and ( n58533 , n58531 , n58532 );
xor ( n58534 , n58531 , n58532 );
xor ( n58535 , n58056 , n58168 );
and ( n58536 , n30319 , n58292 );
and ( n58537 , n58535 , n58536 );
xor ( n58538 , n58535 , n58536 );
xor ( n58539 , n58060 , n58166 );
and ( n58540 , n30324 , n58292 );
and ( n58541 , n58539 , n58540 );
xor ( n58542 , n58539 , n58540 );
xor ( n58543 , n58064 , n58164 );
and ( n58544 , n30329 , n58292 );
and ( n58545 , n58543 , n58544 );
xor ( n58546 , n58543 , n58544 );
xor ( n58547 , n58068 , n58162 );
and ( n58548 , n30334 , n58292 );
and ( n58549 , n58547 , n58548 );
xor ( n58550 , n58547 , n58548 );
xor ( n58551 , n58072 , n58160 );
and ( n58552 , n30339 , n58292 );
and ( n58553 , n58551 , n58552 );
xor ( n58554 , n58551 , n58552 );
xor ( n58555 , n58076 , n58158 );
and ( n58556 , n30344 , n58292 );
and ( n58557 , n58555 , n58556 );
xor ( n58558 , n58555 , n58556 );
xor ( n58559 , n58080 , n58156 );
and ( n58560 , n30349 , n58292 );
and ( n58561 , n58559 , n58560 );
xor ( n58562 , n58559 , n58560 );
xor ( n58563 , n58084 , n58154 );
and ( n58564 , n30354 , n58292 );
and ( n58565 , n58563 , n58564 );
xor ( n58566 , n58563 , n58564 );
xor ( n58567 , n58088 , n58152 );
and ( n58568 , n30359 , n58292 );
and ( n58569 , n58567 , n58568 );
xor ( n58570 , n58567 , n58568 );
xor ( n58571 , n58092 , n58150 );
and ( n58572 , n30364 , n58292 );
and ( n58573 , n58571 , n58572 );
xor ( n58574 , n58571 , n58572 );
xor ( n58575 , n58096 , n58148 );
and ( n58576 , n30369 , n58292 );
and ( n58577 , n58575 , n58576 );
xor ( n58578 , n58575 , n58576 );
xor ( n58579 , n58100 , n58146 );
and ( n58580 , n30374 , n58292 );
and ( n58581 , n58579 , n58580 );
xor ( n58582 , n58579 , n58580 );
xor ( n58583 , n58104 , n58144 );
and ( n58584 , n30379 , n58292 );
and ( n58585 , n58583 , n58584 );
xor ( n58586 , n58583 , n58584 );
xor ( n58587 , n58108 , n58142 );
and ( n58588 , n30384 , n58292 );
and ( n58589 , n58587 , n58588 );
xor ( n58590 , n58587 , n58588 );
xor ( n58591 , n58112 , n58140 );
and ( n58592 , n30389 , n58292 );
and ( n58593 , n58591 , n58592 );
xor ( n58594 , n58591 , n58592 );
xor ( n58595 , n58116 , n58138 );
and ( n58596 , n30394 , n58292 );
and ( n58597 , n58595 , n58596 );
xor ( n58598 , n58595 , n58596 );
xor ( n58599 , n58120 , n58136 );
and ( n58600 , n30399 , n58292 );
and ( n58601 , n58599 , n58600 );
xor ( n58602 , n58599 , n58600 );
xor ( n58603 , n58124 , n58134 );
and ( n58604 , n30404 , n58292 );
and ( n58605 , n58603 , n58604 );
xor ( n58606 , n58603 , n58604 );
xor ( n58607 , n58128 , n58132 );
and ( n58608 , n30409 , n58292 );
and ( n58609 , n58607 , n58608 );
buf ( n58610 , n58609 );
and ( n58611 , n58606 , n58610 );
or ( n58612 , n58605 , n58611 );
and ( n58613 , n58602 , n58612 );
or ( n58614 , n58601 , n58613 );
and ( n58615 , n58598 , n58614 );
or ( n58616 , n58597 , n58615 );
and ( n58617 , n58594 , n58616 );
or ( n58618 , n58593 , n58617 );
and ( n58619 , n58590 , n58618 );
or ( n58620 , n58589 , n58619 );
and ( n58621 , n58586 , n58620 );
or ( n58622 , n58585 , n58621 );
and ( n58623 , n58582 , n58622 );
or ( n58624 , n58581 , n58623 );
and ( n58625 , n58578 , n58624 );
or ( n58626 , n58577 , n58625 );
and ( n58627 , n58574 , n58626 );
or ( n58628 , n58573 , n58627 );
and ( n58629 , n58570 , n58628 );
or ( n58630 , n58569 , n58629 );
and ( n58631 , n58566 , n58630 );
or ( n58632 , n58565 , n58631 );
and ( n58633 , n58562 , n58632 );
or ( n58634 , n58561 , n58633 );
and ( n58635 , n58558 , n58634 );
or ( n58636 , n58557 , n58635 );
and ( n58637 , n58554 , n58636 );
or ( n58638 , n58553 , n58637 );
and ( n58639 , n58550 , n58638 );
or ( n58640 , n58549 , n58639 );
and ( n58641 , n58546 , n58640 );
or ( n58642 , n58545 , n58641 );
and ( n58643 , n58542 , n58642 );
or ( n58644 , n58541 , n58643 );
and ( n58645 , n58538 , n58644 );
or ( n58646 , n58537 , n58645 );
and ( n58647 , n58534 , n58646 );
or ( n58648 , n58533 , n58647 );
and ( n58649 , n58530 , n58648 );
or ( n58650 , n58529 , n58649 );
and ( n58651 , n58526 , n58650 );
or ( n58652 , n58525 , n58651 );
and ( n58653 , n58522 , n58652 );
or ( n58654 , n58521 , n58653 );
and ( n58655 , n58518 , n58654 );
or ( n58656 , n58517 , n58655 );
and ( n58657 , n58514 , n58656 );
or ( n58658 , n58513 , n58657 );
and ( n58659 , n58510 , n58658 );
or ( n58660 , n58509 , n58659 );
and ( n58661 , n58506 , n58660 );
or ( n58662 , n58505 , n58661 );
and ( n58663 , n58502 , n58662 );
or ( n58664 , n58501 , n58663 );
and ( n58665 , n58498 , n58664 );
or ( n58666 , n58497 , n58665 );
and ( n58667 , n58494 , n58666 );
or ( n58668 , n58493 , n58667 );
and ( n58669 , n58490 , n58668 );
or ( n58670 , n58489 , n58669 );
and ( n58671 , n58486 , n58670 );
or ( n58672 , n58485 , n58671 );
and ( n58673 , n58482 , n58672 );
or ( n58674 , n58481 , n58673 );
and ( n58675 , n58478 , n58674 );
or ( n58676 , n58477 , n58675 );
and ( n58677 , n58474 , n58676 );
or ( n58678 , n58473 , n58677 );
and ( n58679 , n58470 , n58678 );
or ( n58680 , n58469 , n58679 );
and ( n58681 , n58466 , n58680 );
or ( n58682 , n58465 , n58681 );
and ( n58683 , n58462 , n58682 );
or ( n58684 , n58461 , n58683 );
and ( n58685 , n58458 , n58684 );
or ( n58686 , n58457 , n58685 );
and ( n58687 , n58454 , n58686 );
or ( n58688 , n58453 , n58687 );
and ( n58689 , n58450 , n58688 );
or ( n58690 , n58449 , n58689 );
and ( n58691 , n58446 , n58690 );
or ( n58692 , n58445 , n58691 );
and ( n58693 , n58442 , n58692 );
or ( n58694 , n58441 , n58693 );
and ( n58695 , n58438 , n58694 );
or ( n58696 , n58437 , n58695 );
and ( n58697 , n58434 , n58696 );
or ( n58698 , n58433 , n58697 );
and ( n58699 , n58430 , n58698 );
or ( n58700 , n58429 , n58699 );
and ( n58701 , n58426 , n58700 );
or ( n58702 , n58425 , n58701 );
and ( n58703 , n58422 , n58702 );
or ( n58704 , n58421 , n58703 );
and ( n58705 , n58418 , n58704 );
or ( n58706 , n58417 , n58705 );
and ( n58707 , n58414 , n58706 );
or ( n58708 , n58413 , n58707 );
and ( n58709 , n58410 , n58708 );
or ( n58710 , n58409 , n58709 );
and ( n58711 , n58406 , n58710 );
or ( n58712 , n58405 , n58711 );
and ( n58713 , n58402 , n58712 );
or ( n58714 , n58401 , n58713 );
and ( n58715 , n58398 , n58714 );
or ( n58716 , n58397 , n58715 );
and ( n58717 , n58394 , n58716 );
or ( n58718 , n58393 , n58717 );
and ( n58719 , n58390 , n58718 );
or ( n58720 , n58389 , n58719 );
and ( n58721 , n58386 , n58720 );
or ( n58722 , n58385 , n58721 );
and ( n58723 , n58382 , n58722 );
or ( n58724 , n58381 , n58723 );
and ( n58725 , n58378 , n58724 );
or ( n58726 , n58377 , n58725 );
and ( n58727 , n58374 , n58726 );
or ( n58728 , n58373 , n58727 );
and ( n58729 , n58370 , n58728 );
or ( n58730 , n58369 , n58729 );
and ( n58731 , n58366 , n58730 );
or ( n58732 , n58365 , n58731 );
and ( n58733 , n58362 , n58732 );
or ( n58734 , n58361 , n58733 );
and ( n58735 , n58358 , n58734 );
or ( n58736 , n58357 , n58735 );
and ( n58737 , n58354 , n58736 );
or ( n58738 , n58353 , n58737 );
and ( n58739 , n58350 , n58738 );
or ( n58740 , n58349 , n58739 );
and ( n58741 , n58346 , n58740 );
or ( n58742 , n58345 , n58741 );
and ( n58743 , n58342 , n58742 );
or ( n58744 , n58341 , n58743 );
and ( n58745 , n58338 , n58744 );
or ( n58746 , n58337 , n58745 );
and ( n58747 , n58334 , n58746 );
or ( n58748 , n58333 , n58747 );
and ( n58749 , n58330 , n58748 );
or ( n58750 , n58329 , n58749 );
and ( n58751 , n58326 , n58750 );
or ( n58752 , n58325 , n58751 );
and ( n58753 , n58322 , n58752 );
or ( n58754 , n58321 , n58753 );
and ( n58755 , n58318 , n58754 );
or ( n58756 , n58317 , n58755 );
and ( n58757 , n58314 , n58756 );
or ( n58758 , n58313 , n58757 );
and ( n58759 , n58310 , n58758 );
or ( n58760 , n58309 , n58759 );
and ( n58761 , n58306 , n58760 );
or ( n58762 , n58305 , n58761 );
and ( n58763 , n58302 , n58762 );
or ( n58764 , n58301 , n58763 );
and ( n58765 , n58298 , n58764 );
or ( n58766 , n58297 , n58765 );
xor ( n58767 , n58294 , n58766 );
buf ( n58768 , n18010 );
and ( n58769 , n30019 , n58768 );
xor ( n58770 , n58767 , n58769 );
xor ( n58771 , n58298 , n58764 );
and ( n58772 , n30024 , n58768 );
and ( n58773 , n58771 , n58772 );
xor ( n58774 , n58771 , n58772 );
xor ( n58775 , n58302 , n58762 );
and ( n58776 , n30029 , n58768 );
and ( n58777 , n58775 , n58776 );
xor ( n58778 , n58775 , n58776 );
xor ( n58779 , n58306 , n58760 );
and ( n58780 , n30034 , n58768 );
and ( n58781 , n58779 , n58780 );
xor ( n58782 , n58779 , n58780 );
xor ( n58783 , n58310 , n58758 );
and ( n58784 , n30039 , n58768 );
and ( n58785 , n58783 , n58784 );
xor ( n58786 , n58783 , n58784 );
xor ( n58787 , n58314 , n58756 );
and ( n58788 , n30044 , n58768 );
and ( n58789 , n58787 , n58788 );
xor ( n58790 , n58787 , n58788 );
xor ( n58791 , n58318 , n58754 );
and ( n58792 , n30049 , n58768 );
and ( n58793 , n58791 , n58792 );
xor ( n58794 , n58791 , n58792 );
xor ( n58795 , n58322 , n58752 );
and ( n58796 , n30054 , n58768 );
and ( n58797 , n58795 , n58796 );
xor ( n58798 , n58795 , n58796 );
xor ( n58799 , n58326 , n58750 );
and ( n58800 , n30059 , n58768 );
and ( n58801 , n58799 , n58800 );
xor ( n58802 , n58799 , n58800 );
xor ( n58803 , n58330 , n58748 );
and ( n58804 , n30064 , n58768 );
and ( n58805 , n58803 , n58804 );
xor ( n58806 , n58803 , n58804 );
xor ( n58807 , n58334 , n58746 );
and ( n58808 , n30069 , n58768 );
and ( n58809 , n58807 , n58808 );
xor ( n58810 , n58807 , n58808 );
xor ( n58811 , n58338 , n58744 );
and ( n58812 , n30074 , n58768 );
and ( n58813 , n58811 , n58812 );
xor ( n58814 , n58811 , n58812 );
xor ( n58815 , n58342 , n58742 );
and ( n58816 , n30079 , n58768 );
and ( n58817 , n58815 , n58816 );
xor ( n58818 , n58815 , n58816 );
xor ( n58819 , n58346 , n58740 );
and ( n58820 , n30084 , n58768 );
and ( n58821 , n58819 , n58820 );
xor ( n58822 , n58819 , n58820 );
xor ( n58823 , n58350 , n58738 );
and ( n58824 , n30089 , n58768 );
and ( n58825 , n58823 , n58824 );
xor ( n58826 , n58823 , n58824 );
xor ( n58827 , n58354 , n58736 );
and ( n58828 , n30094 , n58768 );
and ( n58829 , n58827 , n58828 );
xor ( n58830 , n58827 , n58828 );
xor ( n58831 , n58358 , n58734 );
and ( n58832 , n30099 , n58768 );
and ( n58833 , n58831 , n58832 );
xor ( n58834 , n58831 , n58832 );
xor ( n58835 , n58362 , n58732 );
and ( n58836 , n30104 , n58768 );
and ( n58837 , n58835 , n58836 );
xor ( n58838 , n58835 , n58836 );
xor ( n58839 , n58366 , n58730 );
and ( n58840 , n30109 , n58768 );
and ( n58841 , n58839 , n58840 );
xor ( n58842 , n58839 , n58840 );
xor ( n58843 , n58370 , n58728 );
and ( n58844 , n30114 , n58768 );
and ( n58845 , n58843 , n58844 );
xor ( n58846 , n58843 , n58844 );
xor ( n58847 , n58374 , n58726 );
and ( n58848 , n30119 , n58768 );
and ( n58849 , n58847 , n58848 );
xor ( n58850 , n58847 , n58848 );
xor ( n58851 , n58378 , n58724 );
and ( n58852 , n30124 , n58768 );
and ( n58853 , n58851 , n58852 );
xor ( n58854 , n58851 , n58852 );
xor ( n58855 , n58382 , n58722 );
and ( n58856 , n30129 , n58768 );
and ( n58857 , n58855 , n58856 );
xor ( n58858 , n58855 , n58856 );
xor ( n58859 , n58386 , n58720 );
and ( n58860 , n30134 , n58768 );
and ( n58861 , n58859 , n58860 );
xor ( n58862 , n58859 , n58860 );
xor ( n58863 , n58390 , n58718 );
and ( n58864 , n30139 , n58768 );
and ( n58865 , n58863 , n58864 );
xor ( n58866 , n58863 , n58864 );
xor ( n58867 , n58394 , n58716 );
and ( n58868 , n30144 , n58768 );
and ( n58869 , n58867 , n58868 );
xor ( n58870 , n58867 , n58868 );
xor ( n58871 , n58398 , n58714 );
and ( n58872 , n30149 , n58768 );
and ( n58873 , n58871 , n58872 );
xor ( n58874 , n58871 , n58872 );
xor ( n58875 , n58402 , n58712 );
and ( n58876 , n30154 , n58768 );
and ( n58877 , n58875 , n58876 );
xor ( n58878 , n58875 , n58876 );
xor ( n58879 , n58406 , n58710 );
and ( n58880 , n30159 , n58768 );
and ( n58881 , n58879 , n58880 );
xor ( n58882 , n58879 , n58880 );
xor ( n58883 , n58410 , n58708 );
and ( n58884 , n30164 , n58768 );
and ( n58885 , n58883 , n58884 );
xor ( n58886 , n58883 , n58884 );
xor ( n58887 , n58414 , n58706 );
and ( n58888 , n30169 , n58768 );
and ( n58889 , n58887 , n58888 );
xor ( n58890 , n58887 , n58888 );
xor ( n58891 , n58418 , n58704 );
and ( n58892 , n30174 , n58768 );
and ( n58893 , n58891 , n58892 );
xor ( n58894 , n58891 , n58892 );
xor ( n58895 , n58422 , n58702 );
and ( n58896 , n30179 , n58768 );
and ( n58897 , n58895 , n58896 );
xor ( n58898 , n58895 , n58896 );
xor ( n58899 , n58426 , n58700 );
and ( n58900 , n30184 , n58768 );
and ( n58901 , n58899 , n58900 );
xor ( n58902 , n58899 , n58900 );
xor ( n58903 , n58430 , n58698 );
and ( n58904 , n30189 , n58768 );
and ( n58905 , n58903 , n58904 );
xor ( n58906 , n58903 , n58904 );
xor ( n58907 , n58434 , n58696 );
and ( n58908 , n30194 , n58768 );
and ( n58909 , n58907 , n58908 );
xor ( n58910 , n58907 , n58908 );
xor ( n58911 , n58438 , n58694 );
and ( n58912 , n30199 , n58768 );
and ( n58913 , n58911 , n58912 );
xor ( n58914 , n58911 , n58912 );
xor ( n58915 , n58442 , n58692 );
and ( n58916 , n30204 , n58768 );
and ( n58917 , n58915 , n58916 );
xor ( n58918 , n58915 , n58916 );
xor ( n58919 , n58446 , n58690 );
and ( n58920 , n30209 , n58768 );
and ( n58921 , n58919 , n58920 );
xor ( n58922 , n58919 , n58920 );
xor ( n58923 , n58450 , n58688 );
and ( n58924 , n30214 , n58768 );
and ( n58925 , n58923 , n58924 );
xor ( n58926 , n58923 , n58924 );
xor ( n58927 , n58454 , n58686 );
and ( n58928 , n30219 , n58768 );
and ( n58929 , n58927 , n58928 );
xor ( n58930 , n58927 , n58928 );
xor ( n58931 , n58458 , n58684 );
and ( n58932 , n30224 , n58768 );
and ( n58933 , n58931 , n58932 );
xor ( n58934 , n58931 , n58932 );
xor ( n58935 , n58462 , n58682 );
and ( n58936 , n30229 , n58768 );
and ( n58937 , n58935 , n58936 );
xor ( n58938 , n58935 , n58936 );
xor ( n58939 , n58466 , n58680 );
and ( n58940 , n30234 , n58768 );
and ( n58941 , n58939 , n58940 );
xor ( n58942 , n58939 , n58940 );
xor ( n58943 , n58470 , n58678 );
and ( n58944 , n30239 , n58768 );
and ( n58945 , n58943 , n58944 );
xor ( n58946 , n58943 , n58944 );
xor ( n58947 , n58474 , n58676 );
and ( n58948 , n30244 , n58768 );
and ( n58949 , n58947 , n58948 );
xor ( n58950 , n58947 , n58948 );
xor ( n58951 , n58478 , n58674 );
and ( n58952 , n30249 , n58768 );
and ( n58953 , n58951 , n58952 );
xor ( n58954 , n58951 , n58952 );
xor ( n58955 , n58482 , n58672 );
and ( n58956 , n30254 , n58768 );
and ( n58957 , n58955 , n58956 );
xor ( n58958 , n58955 , n58956 );
xor ( n58959 , n58486 , n58670 );
and ( n58960 , n30259 , n58768 );
and ( n58961 , n58959 , n58960 );
xor ( n58962 , n58959 , n58960 );
xor ( n58963 , n58490 , n58668 );
and ( n58964 , n30264 , n58768 );
and ( n58965 , n58963 , n58964 );
xor ( n58966 , n58963 , n58964 );
xor ( n58967 , n58494 , n58666 );
and ( n58968 , n30269 , n58768 );
and ( n58969 , n58967 , n58968 );
xor ( n58970 , n58967 , n58968 );
xor ( n58971 , n58498 , n58664 );
and ( n58972 , n30274 , n58768 );
and ( n58973 , n58971 , n58972 );
xor ( n58974 , n58971 , n58972 );
xor ( n58975 , n58502 , n58662 );
and ( n58976 , n30279 , n58768 );
and ( n58977 , n58975 , n58976 );
xor ( n58978 , n58975 , n58976 );
xor ( n58979 , n58506 , n58660 );
and ( n58980 , n30284 , n58768 );
and ( n58981 , n58979 , n58980 );
xor ( n58982 , n58979 , n58980 );
xor ( n58983 , n58510 , n58658 );
and ( n58984 , n30289 , n58768 );
and ( n58985 , n58983 , n58984 );
xor ( n58986 , n58983 , n58984 );
xor ( n58987 , n58514 , n58656 );
and ( n58988 , n30294 , n58768 );
and ( n58989 , n58987 , n58988 );
xor ( n58990 , n58987 , n58988 );
xor ( n58991 , n58518 , n58654 );
and ( n58992 , n30299 , n58768 );
and ( n58993 , n58991 , n58992 );
xor ( n58994 , n58991 , n58992 );
xor ( n58995 , n58522 , n58652 );
and ( n58996 , n30304 , n58768 );
and ( n58997 , n58995 , n58996 );
xor ( n58998 , n58995 , n58996 );
xor ( n58999 , n58526 , n58650 );
and ( n59000 , n30309 , n58768 );
and ( n59001 , n58999 , n59000 );
xor ( n59002 , n58999 , n59000 );
xor ( n59003 , n58530 , n58648 );
and ( n59004 , n30314 , n58768 );
and ( n59005 , n59003 , n59004 );
xor ( n59006 , n59003 , n59004 );
xor ( n59007 , n58534 , n58646 );
and ( n59008 , n30319 , n58768 );
and ( n59009 , n59007 , n59008 );
xor ( n59010 , n59007 , n59008 );
xor ( n59011 , n58538 , n58644 );
and ( n59012 , n30324 , n58768 );
and ( n59013 , n59011 , n59012 );
xor ( n59014 , n59011 , n59012 );
xor ( n59015 , n58542 , n58642 );
and ( n59016 , n30329 , n58768 );
and ( n59017 , n59015 , n59016 );
xor ( n59018 , n59015 , n59016 );
xor ( n59019 , n58546 , n58640 );
and ( n59020 , n30334 , n58768 );
and ( n59021 , n59019 , n59020 );
xor ( n59022 , n59019 , n59020 );
xor ( n59023 , n58550 , n58638 );
and ( n59024 , n30339 , n58768 );
and ( n59025 , n59023 , n59024 );
xor ( n59026 , n59023 , n59024 );
xor ( n59027 , n58554 , n58636 );
and ( n59028 , n30344 , n58768 );
and ( n59029 , n59027 , n59028 );
xor ( n59030 , n59027 , n59028 );
xor ( n59031 , n58558 , n58634 );
and ( n59032 , n30349 , n58768 );
and ( n59033 , n59031 , n59032 );
xor ( n59034 , n59031 , n59032 );
xor ( n59035 , n58562 , n58632 );
and ( n59036 , n30354 , n58768 );
and ( n59037 , n59035 , n59036 );
xor ( n59038 , n59035 , n59036 );
xor ( n59039 , n58566 , n58630 );
and ( n59040 , n30359 , n58768 );
and ( n59041 , n59039 , n59040 );
xor ( n59042 , n59039 , n59040 );
xor ( n59043 , n58570 , n58628 );
and ( n59044 , n30364 , n58768 );
and ( n59045 , n59043 , n59044 );
xor ( n59046 , n59043 , n59044 );
xor ( n59047 , n58574 , n58626 );
and ( n59048 , n30369 , n58768 );
and ( n59049 , n59047 , n59048 );
xor ( n59050 , n59047 , n59048 );
xor ( n59051 , n58578 , n58624 );
and ( n59052 , n30374 , n58768 );
and ( n59053 , n59051 , n59052 );
xor ( n59054 , n59051 , n59052 );
xor ( n59055 , n58582 , n58622 );
and ( n59056 , n30379 , n58768 );
and ( n59057 , n59055 , n59056 );
xor ( n59058 , n59055 , n59056 );
xor ( n59059 , n58586 , n58620 );
and ( n59060 , n30384 , n58768 );
and ( n59061 , n59059 , n59060 );
xor ( n59062 , n59059 , n59060 );
xor ( n59063 , n58590 , n58618 );
and ( n59064 , n30389 , n58768 );
and ( n59065 , n59063 , n59064 );
xor ( n59066 , n59063 , n59064 );
xor ( n59067 , n58594 , n58616 );
and ( n59068 , n30394 , n58768 );
and ( n59069 , n59067 , n59068 );
xor ( n59070 , n59067 , n59068 );
xor ( n59071 , n58598 , n58614 );
and ( n59072 , n30399 , n58768 );
and ( n59073 , n59071 , n59072 );
xor ( n59074 , n59071 , n59072 );
xor ( n59075 , n58602 , n58612 );
and ( n59076 , n30404 , n58768 );
and ( n59077 , n59075 , n59076 );
xor ( n59078 , n59075 , n59076 );
xor ( n59079 , n58606 , n58610 );
and ( n59080 , n30409 , n58768 );
and ( n59081 , n59079 , n59080 );
buf ( n59082 , n59081 );
and ( n59083 , n59078 , n59082 );
or ( n59084 , n59077 , n59083 );
and ( n59085 , n59074 , n59084 );
or ( n59086 , n59073 , n59085 );
and ( n59087 , n59070 , n59086 );
or ( n59088 , n59069 , n59087 );
and ( n59089 , n59066 , n59088 );
or ( n59090 , n59065 , n59089 );
and ( n59091 , n59062 , n59090 );
or ( n59092 , n59061 , n59091 );
and ( n59093 , n59058 , n59092 );
or ( n59094 , n59057 , n59093 );
and ( n59095 , n59054 , n59094 );
or ( n59096 , n59053 , n59095 );
and ( n59097 , n59050 , n59096 );
or ( n59098 , n59049 , n59097 );
and ( n59099 , n59046 , n59098 );
or ( n59100 , n59045 , n59099 );
and ( n59101 , n59042 , n59100 );
or ( n59102 , n59041 , n59101 );
and ( n59103 , n59038 , n59102 );
or ( n59104 , n59037 , n59103 );
and ( n59105 , n59034 , n59104 );
or ( n59106 , n59033 , n59105 );
and ( n59107 , n59030 , n59106 );
or ( n59108 , n59029 , n59107 );
and ( n59109 , n59026 , n59108 );
or ( n59110 , n59025 , n59109 );
and ( n59111 , n59022 , n59110 );
or ( n59112 , n59021 , n59111 );
and ( n59113 , n59018 , n59112 );
or ( n59114 , n59017 , n59113 );
and ( n59115 , n59014 , n59114 );
or ( n59116 , n59013 , n59115 );
and ( n59117 , n59010 , n59116 );
or ( n59118 , n59009 , n59117 );
and ( n59119 , n59006 , n59118 );
or ( n59120 , n59005 , n59119 );
and ( n59121 , n59002 , n59120 );
or ( n59122 , n59001 , n59121 );
and ( n59123 , n58998 , n59122 );
or ( n59124 , n58997 , n59123 );
and ( n59125 , n58994 , n59124 );
or ( n59126 , n58993 , n59125 );
and ( n59127 , n58990 , n59126 );
or ( n59128 , n58989 , n59127 );
and ( n59129 , n58986 , n59128 );
or ( n59130 , n58985 , n59129 );
and ( n59131 , n58982 , n59130 );
or ( n59132 , n58981 , n59131 );
and ( n59133 , n58978 , n59132 );
or ( n59134 , n58977 , n59133 );
and ( n59135 , n58974 , n59134 );
or ( n59136 , n58973 , n59135 );
and ( n59137 , n58970 , n59136 );
or ( n59138 , n58969 , n59137 );
and ( n59139 , n58966 , n59138 );
or ( n59140 , n58965 , n59139 );
and ( n59141 , n58962 , n59140 );
or ( n59142 , n58961 , n59141 );
and ( n59143 , n58958 , n59142 );
or ( n59144 , n58957 , n59143 );
and ( n59145 , n58954 , n59144 );
or ( n59146 , n58953 , n59145 );
and ( n59147 , n58950 , n59146 );
or ( n59148 , n58949 , n59147 );
and ( n59149 , n58946 , n59148 );
or ( n59150 , n58945 , n59149 );
and ( n59151 , n58942 , n59150 );
or ( n59152 , n58941 , n59151 );
and ( n59153 , n58938 , n59152 );
or ( n59154 , n58937 , n59153 );
and ( n59155 , n58934 , n59154 );
or ( n59156 , n58933 , n59155 );
and ( n59157 , n58930 , n59156 );
or ( n59158 , n58929 , n59157 );
and ( n59159 , n58926 , n59158 );
or ( n59160 , n58925 , n59159 );
and ( n59161 , n58922 , n59160 );
or ( n59162 , n58921 , n59161 );
and ( n59163 , n58918 , n59162 );
or ( n59164 , n58917 , n59163 );
and ( n59165 , n58914 , n59164 );
or ( n59166 , n58913 , n59165 );
and ( n59167 , n58910 , n59166 );
or ( n59168 , n58909 , n59167 );
and ( n59169 , n58906 , n59168 );
or ( n59170 , n58905 , n59169 );
and ( n59171 , n58902 , n59170 );
or ( n59172 , n58901 , n59171 );
and ( n59173 , n58898 , n59172 );
or ( n59174 , n58897 , n59173 );
and ( n59175 , n58894 , n59174 );
or ( n59176 , n58893 , n59175 );
and ( n59177 , n58890 , n59176 );
or ( n59178 , n58889 , n59177 );
and ( n59179 , n58886 , n59178 );
or ( n59180 , n58885 , n59179 );
and ( n59181 , n58882 , n59180 );
or ( n59182 , n58881 , n59181 );
and ( n59183 , n58878 , n59182 );
or ( n59184 , n58877 , n59183 );
and ( n59185 , n58874 , n59184 );
or ( n59186 , n58873 , n59185 );
and ( n59187 , n58870 , n59186 );
or ( n59188 , n58869 , n59187 );
and ( n59189 , n58866 , n59188 );
or ( n59190 , n58865 , n59189 );
and ( n59191 , n58862 , n59190 );
or ( n59192 , n58861 , n59191 );
and ( n59193 , n58858 , n59192 );
or ( n59194 , n58857 , n59193 );
and ( n59195 , n58854 , n59194 );
or ( n59196 , n58853 , n59195 );
and ( n59197 , n58850 , n59196 );
or ( n59198 , n58849 , n59197 );
and ( n59199 , n58846 , n59198 );
or ( n59200 , n58845 , n59199 );
and ( n59201 , n58842 , n59200 );
or ( n59202 , n58841 , n59201 );
and ( n59203 , n58838 , n59202 );
or ( n59204 , n58837 , n59203 );
and ( n59205 , n58834 , n59204 );
or ( n59206 , n58833 , n59205 );
and ( n59207 , n58830 , n59206 );
or ( n59208 , n58829 , n59207 );
and ( n59209 , n58826 , n59208 );
or ( n59210 , n58825 , n59209 );
and ( n59211 , n58822 , n59210 );
or ( n59212 , n58821 , n59211 );
and ( n59213 , n58818 , n59212 );
or ( n59214 , n58817 , n59213 );
and ( n59215 , n58814 , n59214 );
or ( n59216 , n58813 , n59215 );
and ( n59217 , n58810 , n59216 );
or ( n59218 , n58809 , n59217 );
and ( n59219 , n58806 , n59218 );
or ( n59220 , n58805 , n59219 );
and ( n59221 , n58802 , n59220 );
or ( n59222 , n58801 , n59221 );
and ( n59223 , n58798 , n59222 );
or ( n59224 , n58797 , n59223 );
and ( n59225 , n58794 , n59224 );
or ( n59226 , n58793 , n59225 );
and ( n59227 , n58790 , n59226 );
or ( n59228 , n58789 , n59227 );
and ( n59229 , n58786 , n59228 );
or ( n59230 , n58785 , n59229 );
and ( n59231 , n58782 , n59230 );
or ( n59232 , n58781 , n59231 );
and ( n59233 , n58778 , n59232 );
or ( n59234 , n58777 , n59233 );
and ( n59235 , n58774 , n59234 );
or ( n59236 , n58773 , n59235 );
xor ( n59237 , n58770 , n59236 );
buf ( n59238 , n18008 );
and ( n59239 , n30024 , n59238 );
xor ( n59240 , n59237 , n59239 );
xor ( n59241 , n58774 , n59234 );
and ( n59242 , n30029 , n59238 );
and ( n59243 , n59241 , n59242 );
xor ( n59244 , n59241 , n59242 );
xor ( n59245 , n58778 , n59232 );
and ( n59246 , n30034 , n59238 );
and ( n59247 , n59245 , n59246 );
xor ( n59248 , n59245 , n59246 );
xor ( n59249 , n58782 , n59230 );
and ( n59250 , n30039 , n59238 );
and ( n59251 , n59249 , n59250 );
xor ( n59252 , n59249 , n59250 );
xor ( n59253 , n58786 , n59228 );
and ( n59254 , n30044 , n59238 );
and ( n59255 , n59253 , n59254 );
xor ( n59256 , n59253 , n59254 );
xor ( n59257 , n58790 , n59226 );
and ( n59258 , n30049 , n59238 );
and ( n59259 , n59257 , n59258 );
xor ( n59260 , n59257 , n59258 );
xor ( n59261 , n58794 , n59224 );
and ( n59262 , n30054 , n59238 );
and ( n59263 , n59261 , n59262 );
xor ( n59264 , n59261 , n59262 );
xor ( n59265 , n58798 , n59222 );
and ( n59266 , n30059 , n59238 );
and ( n59267 , n59265 , n59266 );
xor ( n59268 , n59265 , n59266 );
xor ( n59269 , n58802 , n59220 );
and ( n59270 , n30064 , n59238 );
and ( n59271 , n59269 , n59270 );
xor ( n59272 , n59269 , n59270 );
xor ( n59273 , n58806 , n59218 );
and ( n59274 , n30069 , n59238 );
and ( n59275 , n59273 , n59274 );
xor ( n59276 , n59273 , n59274 );
xor ( n59277 , n58810 , n59216 );
and ( n59278 , n30074 , n59238 );
and ( n59279 , n59277 , n59278 );
xor ( n59280 , n59277 , n59278 );
xor ( n59281 , n58814 , n59214 );
and ( n59282 , n30079 , n59238 );
and ( n59283 , n59281 , n59282 );
xor ( n59284 , n59281 , n59282 );
xor ( n59285 , n58818 , n59212 );
and ( n59286 , n30084 , n59238 );
and ( n59287 , n59285 , n59286 );
xor ( n59288 , n59285 , n59286 );
xor ( n59289 , n58822 , n59210 );
and ( n59290 , n30089 , n59238 );
and ( n59291 , n59289 , n59290 );
xor ( n59292 , n59289 , n59290 );
xor ( n59293 , n58826 , n59208 );
and ( n59294 , n30094 , n59238 );
and ( n59295 , n59293 , n59294 );
xor ( n59296 , n59293 , n59294 );
xor ( n59297 , n58830 , n59206 );
and ( n59298 , n30099 , n59238 );
and ( n59299 , n59297 , n59298 );
xor ( n59300 , n59297 , n59298 );
xor ( n59301 , n58834 , n59204 );
and ( n59302 , n30104 , n59238 );
and ( n59303 , n59301 , n59302 );
xor ( n59304 , n59301 , n59302 );
xor ( n59305 , n58838 , n59202 );
and ( n59306 , n30109 , n59238 );
and ( n59307 , n59305 , n59306 );
xor ( n59308 , n59305 , n59306 );
xor ( n59309 , n58842 , n59200 );
and ( n59310 , n30114 , n59238 );
and ( n59311 , n59309 , n59310 );
xor ( n59312 , n59309 , n59310 );
xor ( n59313 , n58846 , n59198 );
and ( n59314 , n30119 , n59238 );
and ( n59315 , n59313 , n59314 );
xor ( n59316 , n59313 , n59314 );
xor ( n59317 , n58850 , n59196 );
and ( n59318 , n30124 , n59238 );
and ( n59319 , n59317 , n59318 );
xor ( n59320 , n59317 , n59318 );
xor ( n59321 , n58854 , n59194 );
and ( n59322 , n30129 , n59238 );
and ( n59323 , n59321 , n59322 );
xor ( n59324 , n59321 , n59322 );
xor ( n59325 , n58858 , n59192 );
and ( n59326 , n30134 , n59238 );
and ( n59327 , n59325 , n59326 );
xor ( n59328 , n59325 , n59326 );
xor ( n59329 , n58862 , n59190 );
and ( n59330 , n30139 , n59238 );
and ( n59331 , n59329 , n59330 );
xor ( n59332 , n59329 , n59330 );
xor ( n59333 , n58866 , n59188 );
and ( n59334 , n30144 , n59238 );
and ( n59335 , n59333 , n59334 );
xor ( n59336 , n59333 , n59334 );
xor ( n59337 , n58870 , n59186 );
and ( n59338 , n30149 , n59238 );
and ( n59339 , n59337 , n59338 );
xor ( n59340 , n59337 , n59338 );
xor ( n59341 , n58874 , n59184 );
and ( n59342 , n30154 , n59238 );
and ( n59343 , n59341 , n59342 );
xor ( n59344 , n59341 , n59342 );
xor ( n59345 , n58878 , n59182 );
and ( n59346 , n30159 , n59238 );
and ( n59347 , n59345 , n59346 );
xor ( n59348 , n59345 , n59346 );
xor ( n59349 , n58882 , n59180 );
and ( n59350 , n30164 , n59238 );
and ( n59351 , n59349 , n59350 );
xor ( n59352 , n59349 , n59350 );
xor ( n59353 , n58886 , n59178 );
and ( n59354 , n30169 , n59238 );
and ( n59355 , n59353 , n59354 );
xor ( n59356 , n59353 , n59354 );
xor ( n59357 , n58890 , n59176 );
and ( n59358 , n30174 , n59238 );
and ( n59359 , n59357 , n59358 );
xor ( n59360 , n59357 , n59358 );
xor ( n59361 , n58894 , n59174 );
and ( n59362 , n30179 , n59238 );
and ( n59363 , n59361 , n59362 );
xor ( n59364 , n59361 , n59362 );
xor ( n59365 , n58898 , n59172 );
and ( n59366 , n30184 , n59238 );
and ( n59367 , n59365 , n59366 );
xor ( n59368 , n59365 , n59366 );
xor ( n59369 , n58902 , n59170 );
and ( n59370 , n30189 , n59238 );
and ( n59371 , n59369 , n59370 );
xor ( n59372 , n59369 , n59370 );
xor ( n59373 , n58906 , n59168 );
and ( n59374 , n30194 , n59238 );
and ( n59375 , n59373 , n59374 );
xor ( n59376 , n59373 , n59374 );
xor ( n59377 , n58910 , n59166 );
and ( n59378 , n30199 , n59238 );
and ( n59379 , n59377 , n59378 );
xor ( n59380 , n59377 , n59378 );
xor ( n59381 , n58914 , n59164 );
and ( n59382 , n30204 , n59238 );
and ( n59383 , n59381 , n59382 );
xor ( n59384 , n59381 , n59382 );
xor ( n59385 , n58918 , n59162 );
and ( n59386 , n30209 , n59238 );
and ( n59387 , n59385 , n59386 );
xor ( n59388 , n59385 , n59386 );
xor ( n59389 , n58922 , n59160 );
and ( n59390 , n30214 , n59238 );
and ( n59391 , n59389 , n59390 );
xor ( n59392 , n59389 , n59390 );
xor ( n59393 , n58926 , n59158 );
and ( n59394 , n30219 , n59238 );
and ( n59395 , n59393 , n59394 );
xor ( n59396 , n59393 , n59394 );
xor ( n59397 , n58930 , n59156 );
and ( n59398 , n30224 , n59238 );
and ( n59399 , n59397 , n59398 );
xor ( n59400 , n59397 , n59398 );
xor ( n59401 , n58934 , n59154 );
and ( n59402 , n30229 , n59238 );
and ( n59403 , n59401 , n59402 );
xor ( n59404 , n59401 , n59402 );
xor ( n59405 , n58938 , n59152 );
and ( n59406 , n30234 , n59238 );
and ( n59407 , n59405 , n59406 );
xor ( n59408 , n59405 , n59406 );
xor ( n59409 , n58942 , n59150 );
and ( n59410 , n30239 , n59238 );
and ( n59411 , n59409 , n59410 );
xor ( n59412 , n59409 , n59410 );
xor ( n59413 , n58946 , n59148 );
and ( n59414 , n30244 , n59238 );
and ( n59415 , n59413 , n59414 );
xor ( n59416 , n59413 , n59414 );
xor ( n59417 , n58950 , n59146 );
and ( n59418 , n30249 , n59238 );
and ( n59419 , n59417 , n59418 );
xor ( n59420 , n59417 , n59418 );
xor ( n59421 , n58954 , n59144 );
and ( n59422 , n30254 , n59238 );
and ( n59423 , n59421 , n59422 );
xor ( n59424 , n59421 , n59422 );
xor ( n59425 , n58958 , n59142 );
and ( n59426 , n30259 , n59238 );
and ( n59427 , n59425 , n59426 );
xor ( n59428 , n59425 , n59426 );
xor ( n59429 , n58962 , n59140 );
and ( n59430 , n30264 , n59238 );
and ( n59431 , n59429 , n59430 );
xor ( n59432 , n59429 , n59430 );
xor ( n59433 , n58966 , n59138 );
and ( n59434 , n30269 , n59238 );
and ( n59435 , n59433 , n59434 );
xor ( n59436 , n59433 , n59434 );
xor ( n59437 , n58970 , n59136 );
and ( n59438 , n30274 , n59238 );
and ( n59439 , n59437 , n59438 );
xor ( n59440 , n59437 , n59438 );
xor ( n59441 , n58974 , n59134 );
and ( n59442 , n30279 , n59238 );
and ( n59443 , n59441 , n59442 );
xor ( n59444 , n59441 , n59442 );
xor ( n59445 , n58978 , n59132 );
and ( n59446 , n30284 , n59238 );
and ( n59447 , n59445 , n59446 );
xor ( n59448 , n59445 , n59446 );
xor ( n59449 , n58982 , n59130 );
and ( n59450 , n30289 , n59238 );
and ( n59451 , n59449 , n59450 );
xor ( n59452 , n59449 , n59450 );
xor ( n59453 , n58986 , n59128 );
and ( n59454 , n30294 , n59238 );
and ( n59455 , n59453 , n59454 );
xor ( n59456 , n59453 , n59454 );
xor ( n59457 , n58990 , n59126 );
and ( n59458 , n30299 , n59238 );
and ( n59459 , n59457 , n59458 );
xor ( n59460 , n59457 , n59458 );
xor ( n59461 , n58994 , n59124 );
and ( n59462 , n30304 , n59238 );
and ( n59463 , n59461 , n59462 );
xor ( n59464 , n59461 , n59462 );
xor ( n59465 , n58998 , n59122 );
and ( n59466 , n30309 , n59238 );
and ( n59467 , n59465 , n59466 );
xor ( n59468 , n59465 , n59466 );
xor ( n59469 , n59002 , n59120 );
and ( n59470 , n30314 , n59238 );
and ( n59471 , n59469 , n59470 );
xor ( n59472 , n59469 , n59470 );
xor ( n59473 , n59006 , n59118 );
and ( n59474 , n30319 , n59238 );
and ( n59475 , n59473 , n59474 );
xor ( n59476 , n59473 , n59474 );
xor ( n59477 , n59010 , n59116 );
and ( n59478 , n30324 , n59238 );
and ( n59479 , n59477 , n59478 );
xor ( n59480 , n59477 , n59478 );
xor ( n59481 , n59014 , n59114 );
and ( n59482 , n30329 , n59238 );
and ( n59483 , n59481 , n59482 );
xor ( n59484 , n59481 , n59482 );
xor ( n59485 , n59018 , n59112 );
and ( n59486 , n30334 , n59238 );
and ( n59487 , n59485 , n59486 );
xor ( n59488 , n59485 , n59486 );
xor ( n59489 , n59022 , n59110 );
and ( n59490 , n30339 , n59238 );
and ( n59491 , n59489 , n59490 );
xor ( n59492 , n59489 , n59490 );
xor ( n59493 , n59026 , n59108 );
and ( n59494 , n30344 , n59238 );
and ( n59495 , n59493 , n59494 );
xor ( n59496 , n59493 , n59494 );
xor ( n59497 , n59030 , n59106 );
and ( n59498 , n30349 , n59238 );
and ( n59499 , n59497 , n59498 );
xor ( n59500 , n59497 , n59498 );
xor ( n59501 , n59034 , n59104 );
and ( n59502 , n30354 , n59238 );
and ( n59503 , n59501 , n59502 );
xor ( n59504 , n59501 , n59502 );
xor ( n59505 , n59038 , n59102 );
and ( n59506 , n30359 , n59238 );
and ( n59507 , n59505 , n59506 );
xor ( n59508 , n59505 , n59506 );
xor ( n59509 , n59042 , n59100 );
and ( n59510 , n30364 , n59238 );
and ( n59511 , n59509 , n59510 );
xor ( n59512 , n59509 , n59510 );
xor ( n59513 , n59046 , n59098 );
and ( n59514 , n30369 , n59238 );
and ( n59515 , n59513 , n59514 );
xor ( n59516 , n59513 , n59514 );
xor ( n59517 , n59050 , n59096 );
and ( n59518 , n30374 , n59238 );
and ( n59519 , n59517 , n59518 );
xor ( n59520 , n59517 , n59518 );
xor ( n59521 , n59054 , n59094 );
and ( n59522 , n30379 , n59238 );
and ( n59523 , n59521 , n59522 );
xor ( n59524 , n59521 , n59522 );
xor ( n59525 , n59058 , n59092 );
and ( n59526 , n30384 , n59238 );
and ( n59527 , n59525 , n59526 );
xor ( n59528 , n59525 , n59526 );
xor ( n59529 , n59062 , n59090 );
and ( n59530 , n30389 , n59238 );
and ( n59531 , n59529 , n59530 );
xor ( n59532 , n59529 , n59530 );
xor ( n59533 , n59066 , n59088 );
and ( n59534 , n30394 , n59238 );
and ( n59535 , n59533 , n59534 );
xor ( n59536 , n59533 , n59534 );
xor ( n59537 , n59070 , n59086 );
and ( n59538 , n30399 , n59238 );
and ( n59539 , n59537 , n59538 );
xor ( n59540 , n59537 , n59538 );
xor ( n59541 , n59074 , n59084 );
and ( n59542 , n30404 , n59238 );
and ( n59543 , n59541 , n59542 );
xor ( n59544 , n59541 , n59542 );
xor ( n59545 , n59078 , n59082 );
and ( n59546 , n30409 , n59238 );
and ( n59547 , n59545 , n59546 );
buf ( n59548 , n59547 );
and ( n59549 , n59544 , n59548 );
or ( n59550 , n59543 , n59549 );
and ( n59551 , n59540 , n59550 );
or ( n59552 , n59539 , n59551 );
and ( n59553 , n59536 , n59552 );
or ( n59554 , n59535 , n59553 );
and ( n59555 , n59532 , n59554 );
or ( n59556 , n59531 , n59555 );
and ( n59557 , n59528 , n59556 );
or ( n59558 , n59527 , n59557 );
and ( n59559 , n59524 , n59558 );
or ( n59560 , n59523 , n59559 );
and ( n59561 , n59520 , n59560 );
or ( n59562 , n59519 , n59561 );
and ( n59563 , n59516 , n59562 );
or ( n59564 , n59515 , n59563 );
and ( n59565 , n59512 , n59564 );
or ( n59566 , n59511 , n59565 );
and ( n59567 , n59508 , n59566 );
or ( n59568 , n59507 , n59567 );
and ( n59569 , n59504 , n59568 );
or ( n59570 , n59503 , n59569 );
and ( n59571 , n59500 , n59570 );
or ( n59572 , n59499 , n59571 );
and ( n59573 , n59496 , n59572 );
or ( n59574 , n59495 , n59573 );
and ( n59575 , n59492 , n59574 );
or ( n59576 , n59491 , n59575 );
and ( n59577 , n59488 , n59576 );
or ( n59578 , n59487 , n59577 );
and ( n59579 , n59484 , n59578 );
or ( n59580 , n59483 , n59579 );
and ( n59581 , n59480 , n59580 );
or ( n59582 , n59479 , n59581 );
and ( n59583 , n59476 , n59582 );
or ( n59584 , n59475 , n59583 );
and ( n59585 , n59472 , n59584 );
or ( n59586 , n59471 , n59585 );
and ( n59587 , n59468 , n59586 );
or ( n59588 , n59467 , n59587 );
and ( n59589 , n59464 , n59588 );
or ( n59590 , n59463 , n59589 );
and ( n59591 , n59460 , n59590 );
or ( n59592 , n59459 , n59591 );
and ( n59593 , n59456 , n59592 );
or ( n59594 , n59455 , n59593 );
and ( n59595 , n59452 , n59594 );
or ( n59596 , n59451 , n59595 );
and ( n59597 , n59448 , n59596 );
or ( n59598 , n59447 , n59597 );
and ( n59599 , n59444 , n59598 );
or ( n59600 , n59443 , n59599 );
and ( n59601 , n59440 , n59600 );
or ( n59602 , n59439 , n59601 );
and ( n59603 , n59436 , n59602 );
or ( n59604 , n59435 , n59603 );
and ( n59605 , n59432 , n59604 );
or ( n59606 , n59431 , n59605 );
and ( n59607 , n59428 , n59606 );
or ( n59608 , n59427 , n59607 );
and ( n59609 , n59424 , n59608 );
or ( n59610 , n59423 , n59609 );
and ( n59611 , n59420 , n59610 );
or ( n59612 , n59419 , n59611 );
and ( n59613 , n59416 , n59612 );
or ( n59614 , n59415 , n59613 );
and ( n59615 , n59412 , n59614 );
or ( n59616 , n59411 , n59615 );
and ( n59617 , n59408 , n59616 );
or ( n59618 , n59407 , n59617 );
and ( n59619 , n59404 , n59618 );
or ( n59620 , n59403 , n59619 );
and ( n59621 , n59400 , n59620 );
or ( n59622 , n59399 , n59621 );
and ( n59623 , n59396 , n59622 );
or ( n59624 , n59395 , n59623 );
and ( n59625 , n59392 , n59624 );
or ( n59626 , n59391 , n59625 );
and ( n59627 , n59388 , n59626 );
or ( n59628 , n59387 , n59627 );
and ( n59629 , n59384 , n59628 );
or ( n59630 , n59383 , n59629 );
and ( n59631 , n59380 , n59630 );
or ( n59632 , n59379 , n59631 );
and ( n59633 , n59376 , n59632 );
or ( n59634 , n59375 , n59633 );
and ( n59635 , n59372 , n59634 );
or ( n59636 , n59371 , n59635 );
and ( n59637 , n59368 , n59636 );
or ( n59638 , n59367 , n59637 );
and ( n59639 , n59364 , n59638 );
or ( n59640 , n59363 , n59639 );
and ( n59641 , n59360 , n59640 );
or ( n59642 , n59359 , n59641 );
and ( n59643 , n59356 , n59642 );
or ( n59644 , n59355 , n59643 );
and ( n59645 , n59352 , n59644 );
or ( n59646 , n59351 , n59645 );
and ( n59647 , n59348 , n59646 );
or ( n59648 , n59347 , n59647 );
and ( n59649 , n59344 , n59648 );
or ( n59650 , n59343 , n59649 );
and ( n59651 , n59340 , n59650 );
or ( n59652 , n59339 , n59651 );
and ( n59653 , n59336 , n59652 );
or ( n59654 , n59335 , n59653 );
and ( n59655 , n59332 , n59654 );
or ( n59656 , n59331 , n59655 );
and ( n59657 , n59328 , n59656 );
or ( n59658 , n59327 , n59657 );
and ( n59659 , n59324 , n59658 );
or ( n59660 , n59323 , n59659 );
and ( n59661 , n59320 , n59660 );
or ( n59662 , n59319 , n59661 );
and ( n59663 , n59316 , n59662 );
or ( n59664 , n59315 , n59663 );
and ( n59665 , n59312 , n59664 );
or ( n59666 , n59311 , n59665 );
and ( n59667 , n59308 , n59666 );
or ( n59668 , n59307 , n59667 );
and ( n59669 , n59304 , n59668 );
or ( n59670 , n59303 , n59669 );
and ( n59671 , n59300 , n59670 );
or ( n59672 , n59299 , n59671 );
and ( n59673 , n59296 , n59672 );
or ( n59674 , n59295 , n59673 );
and ( n59675 , n59292 , n59674 );
or ( n59676 , n59291 , n59675 );
and ( n59677 , n59288 , n59676 );
or ( n59678 , n59287 , n59677 );
and ( n59679 , n59284 , n59678 );
or ( n59680 , n59283 , n59679 );
and ( n59681 , n59280 , n59680 );
or ( n59682 , n59279 , n59681 );
and ( n59683 , n59276 , n59682 );
or ( n59684 , n59275 , n59683 );
and ( n59685 , n59272 , n59684 );
or ( n59686 , n59271 , n59685 );
and ( n59687 , n59268 , n59686 );
or ( n59688 , n59267 , n59687 );
and ( n59689 , n59264 , n59688 );
or ( n59690 , n59263 , n59689 );
and ( n59691 , n59260 , n59690 );
or ( n59692 , n59259 , n59691 );
and ( n59693 , n59256 , n59692 );
or ( n59694 , n59255 , n59693 );
and ( n59695 , n59252 , n59694 );
or ( n59696 , n59251 , n59695 );
and ( n59697 , n59248 , n59696 );
or ( n59698 , n59247 , n59697 );
and ( n59699 , n59244 , n59698 );
or ( n59700 , n59243 , n59699 );
xor ( n59701 , n59240 , n59700 );
buf ( n59702 , n18006 );
and ( n59703 , n30029 , n59702 );
xor ( n59704 , n59701 , n59703 );
xor ( n59705 , n59244 , n59698 );
and ( n59706 , n30034 , n59702 );
and ( n59707 , n59705 , n59706 );
xor ( n59708 , n59705 , n59706 );
xor ( n59709 , n59248 , n59696 );
and ( n59710 , n30039 , n59702 );
and ( n59711 , n59709 , n59710 );
xor ( n59712 , n59709 , n59710 );
xor ( n59713 , n59252 , n59694 );
and ( n59714 , n30044 , n59702 );
and ( n59715 , n59713 , n59714 );
xor ( n59716 , n59713 , n59714 );
xor ( n59717 , n59256 , n59692 );
and ( n59718 , n30049 , n59702 );
and ( n59719 , n59717 , n59718 );
xor ( n59720 , n59717 , n59718 );
xor ( n59721 , n59260 , n59690 );
and ( n59722 , n30054 , n59702 );
and ( n59723 , n59721 , n59722 );
xor ( n59724 , n59721 , n59722 );
xor ( n59725 , n59264 , n59688 );
and ( n59726 , n30059 , n59702 );
and ( n59727 , n59725 , n59726 );
xor ( n59728 , n59725 , n59726 );
xor ( n59729 , n59268 , n59686 );
and ( n59730 , n30064 , n59702 );
and ( n59731 , n59729 , n59730 );
xor ( n59732 , n59729 , n59730 );
xor ( n59733 , n59272 , n59684 );
and ( n59734 , n30069 , n59702 );
and ( n59735 , n59733 , n59734 );
xor ( n59736 , n59733 , n59734 );
xor ( n59737 , n59276 , n59682 );
and ( n59738 , n30074 , n59702 );
and ( n59739 , n59737 , n59738 );
xor ( n59740 , n59737 , n59738 );
xor ( n59741 , n59280 , n59680 );
and ( n59742 , n30079 , n59702 );
and ( n59743 , n59741 , n59742 );
xor ( n59744 , n59741 , n59742 );
xor ( n59745 , n59284 , n59678 );
and ( n59746 , n30084 , n59702 );
and ( n59747 , n59745 , n59746 );
xor ( n59748 , n59745 , n59746 );
xor ( n59749 , n59288 , n59676 );
and ( n59750 , n30089 , n59702 );
and ( n59751 , n59749 , n59750 );
xor ( n59752 , n59749 , n59750 );
xor ( n59753 , n59292 , n59674 );
and ( n59754 , n30094 , n59702 );
and ( n59755 , n59753 , n59754 );
xor ( n59756 , n59753 , n59754 );
xor ( n59757 , n59296 , n59672 );
and ( n59758 , n30099 , n59702 );
and ( n59759 , n59757 , n59758 );
xor ( n59760 , n59757 , n59758 );
xor ( n59761 , n59300 , n59670 );
and ( n59762 , n30104 , n59702 );
and ( n59763 , n59761 , n59762 );
xor ( n59764 , n59761 , n59762 );
xor ( n59765 , n59304 , n59668 );
and ( n59766 , n30109 , n59702 );
and ( n59767 , n59765 , n59766 );
xor ( n59768 , n59765 , n59766 );
xor ( n59769 , n59308 , n59666 );
and ( n59770 , n30114 , n59702 );
and ( n59771 , n59769 , n59770 );
xor ( n59772 , n59769 , n59770 );
xor ( n59773 , n59312 , n59664 );
and ( n59774 , n30119 , n59702 );
and ( n59775 , n59773 , n59774 );
xor ( n59776 , n59773 , n59774 );
xor ( n59777 , n59316 , n59662 );
and ( n59778 , n30124 , n59702 );
and ( n59779 , n59777 , n59778 );
xor ( n59780 , n59777 , n59778 );
xor ( n59781 , n59320 , n59660 );
and ( n59782 , n30129 , n59702 );
and ( n59783 , n59781 , n59782 );
xor ( n59784 , n59781 , n59782 );
xor ( n59785 , n59324 , n59658 );
and ( n59786 , n30134 , n59702 );
and ( n59787 , n59785 , n59786 );
xor ( n59788 , n59785 , n59786 );
xor ( n59789 , n59328 , n59656 );
and ( n59790 , n30139 , n59702 );
and ( n59791 , n59789 , n59790 );
xor ( n59792 , n59789 , n59790 );
xor ( n59793 , n59332 , n59654 );
and ( n59794 , n30144 , n59702 );
and ( n59795 , n59793 , n59794 );
xor ( n59796 , n59793 , n59794 );
xor ( n59797 , n59336 , n59652 );
and ( n59798 , n30149 , n59702 );
and ( n59799 , n59797 , n59798 );
xor ( n59800 , n59797 , n59798 );
xor ( n59801 , n59340 , n59650 );
and ( n59802 , n30154 , n59702 );
and ( n59803 , n59801 , n59802 );
xor ( n59804 , n59801 , n59802 );
xor ( n59805 , n59344 , n59648 );
and ( n59806 , n30159 , n59702 );
and ( n59807 , n59805 , n59806 );
xor ( n59808 , n59805 , n59806 );
xor ( n59809 , n59348 , n59646 );
and ( n59810 , n30164 , n59702 );
and ( n59811 , n59809 , n59810 );
xor ( n59812 , n59809 , n59810 );
xor ( n59813 , n59352 , n59644 );
and ( n59814 , n30169 , n59702 );
and ( n59815 , n59813 , n59814 );
xor ( n59816 , n59813 , n59814 );
xor ( n59817 , n59356 , n59642 );
and ( n59818 , n30174 , n59702 );
and ( n59819 , n59817 , n59818 );
xor ( n59820 , n59817 , n59818 );
xor ( n59821 , n59360 , n59640 );
and ( n59822 , n30179 , n59702 );
and ( n59823 , n59821 , n59822 );
xor ( n59824 , n59821 , n59822 );
xor ( n59825 , n59364 , n59638 );
and ( n59826 , n30184 , n59702 );
and ( n59827 , n59825 , n59826 );
xor ( n59828 , n59825 , n59826 );
xor ( n59829 , n59368 , n59636 );
and ( n59830 , n30189 , n59702 );
and ( n59831 , n59829 , n59830 );
xor ( n59832 , n59829 , n59830 );
xor ( n59833 , n59372 , n59634 );
and ( n59834 , n30194 , n59702 );
and ( n59835 , n59833 , n59834 );
xor ( n59836 , n59833 , n59834 );
xor ( n59837 , n59376 , n59632 );
and ( n59838 , n30199 , n59702 );
and ( n59839 , n59837 , n59838 );
xor ( n59840 , n59837 , n59838 );
xor ( n59841 , n59380 , n59630 );
and ( n59842 , n30204 , n59702 );
and ( n59843 , n59841 , n59842 );
xor ( n59844 , n59841 , n59842 );
xor ( n59845 , n59384 , n59628 );
and ( n59846 , n30209 , n59702 );
and ( n59847 , n59845 , n59846 );
xor ( n59848 , n59845 , n59846 );
xor ( n59849 , n59388 , n59626 );
and ( n59850 , n30214 , n59702 );
and ( n59851 , n59849 , n59850 );
xor ( n59852 , n59849 , n59850 );
xor ( n59853 , n59392 , n59624 );
and ( n59854 , n30219 , n59702 );
and ( n59855 , n59853 , n59854 );
xor ( n59856 , n59853 , n59854 );
xor ( n59857 , n59396 , n59622 );
and ( n59858 , n30224 , n59702 );
and ( n59859 , n59857 , n59858 );
xor ( n59860 , n59857 , n59858 );
xor ( n59861 , n59400 , n59620 );
and ( n59862 , n30229 , n59702 );
and ( n59863 , n59861 , n59862 );
xor ( n59864 , n59861 , n59862 );
xor ( n59865 , n59404 , n59618 );
and ( n59866 , n30234 , n59702 );
and ( n59867 , n59865 , n59866 );
xor ( n59868 , n59865 , n59866 );
xor ( n59869 , n59408 , n59616 );
and ( n59870 , n30239 , n59702 );
and ( n59871 , n59869 , n59870 );
xor ( n59872 , n59869 , n59870 );
xor ( n59873 , n59412 , n59614 );
and ( n59874 , n30244 , n59702 );
and ( n59875 , n59873 , n59874 );
xor ( n59876 , n59873 , n59874 );
xor ( n59877 , n59416 , n59612 );
and ( n59878 , n30249 , n59702 );
and ( n59879 , n59877 , n59878 );
xor ( n59880 , n59877 , n59878 );
xor ( n59881 , n59420 , n59610 );
and ( n59882 , n30254 , n59702 );
and ( n59883 , n59881 , n59882 );
xor ( n59884 , n59881 , n59882 );
xor ( n59885 , n59424 , n59608 );
and ( n59886 , n30259 , n59702 );
and ( n59887 , n59885 , n59886 );
xor ( n59888 , n59885 , n59886 );
xor ( n59889 , n59428 , n59606 );
and ( n59890 , n30264 , n59702 );
and ( n59891 , n59889 , n59890 );
xor ( n59892 , n59889 , n59890 );
xor ( n59893 , n59432 , n59604 );
and ( n59894 , n30269 , n59702 );
and ( n59895 , n59893 , n59894 );
xor ( n59896 , n59893 , n59894 );
xor ( n59897 , n59436 , n59602 );
and ( n59898 , n30274 , n59702 );
and ( n59899 , n59897 , n59898 );
xor ( n59900 , n59897 , n59898 );
xor ( n59901 , n59440 , n59600 );
and ( n59902 , n30279 , n59702 );
and ( n59903 , n59901 , n59902 );
xor ( n59904 , n59901 , n59902 );
xor ( n59905 , n59444 , n59598 );
and ( n59906 , n30284 , n59702 );
and ( n59907 , n59905 , n59906 );
xor ( n59908 , n59905 , n59906 );
xor ( n59909 , n59448 , n59596 );
and ( n59910 , n30289 , n59702 );
and ( n59911 , n59909 , n59910 );
xor ( n59912 , n59909 , n59910 );
xor ( n59913 , n59452 , n59594 );
and ( n59914 , n30294 , n59702 );
and ( n59915 , n59913 , n59914 );
xor ( n59916 , n59913 , n59914 );
xor ( n59917 , n59456 , n59592 );
and ( n59918 , n30299 , n59702 );
and ( n59919 , n59917 , n59918 );
xor ( n59920 , n59917 , n59918 );
xor ( n59921 , n59460 , n59590 );
and ( n59922 , n30304 , n59702 );
and ( n59923 , n59921 , n59922 );
xor ( n59924 , n59921 , n59922 );
xor ( n59925 , n59464 , n59588 );
and ( n59926 , n30309 , n59702 );
and ( n59927 , n59925 , n59926 );
xor ( n59928 , n59925 , n59926 );
xor ( n59929 , n59468 , n59586 );
and ( n59930 , n30314 , n59702 );
and ( n59931 , n59929 , n59930 );
xor ( n59932 , n59929 , n59930 );
xor ( n59933 , n59472 , n59584 );
and ( n59934 , n30319 , n59702 );
and ( n59935 , n59933 , n59934 );
xor ( n59936 , n59933 , n59934 );
xor ( n59937 , n59476 , n59582 );
and ( n59938 , n30324 , n59702 );
and ( n59939 , n59937 , n59938 );
xor ( n59940 , n59937 , n59938 );
xor ( n59941 , n59480 , n59580 );
and ( n59942 , n30329 , n59702 );
and ( n59943 , n59941 , n59942 );
xor ( n59944 , n59941 , n59942 );
xor ( n59945 , n59484 , n59578 );
and ( n59946 , n30334 , n59702 );
and ( n59947 , n59945 , n59946 );
xor ( n59948 , n59945 , n59946 );
xor ( n59949 , n59488 , n59576 );
and ( n59950 , n30339 , n59702 );
and ( n59951 , n59949 , n59950 );
xor ( n59952 , n59949 , n59950 );
xor ( n59953 , n59492 , n59574 );
and ( n59954 , n30344 , n59702 );
and ( n59955 , n59953 , n59954 );
xor ( n59956 , n59953 , n59954 );
xor ( n59957 , n59496 , n59572 );
and ( n59958 , n30349 , n59702 );
and ( n59959 , n59957 , n59958 );
xor ( n59960 , n59957 , n59958 );
xor ( n59961 , n59500 , n59570 );
and ( n59962 , n30354 , n59702 );
and ( n59963 , n59961 , n59962 );
xor ( n59964 , n59961 , n59962 );
xor ( n59965 , n59504 , n59568 );
and ( n59966 , n30359 , n59702 );
and ( n59967 , n59965 , n59966 );
xor ( n59968 , n59965 , n59966 );
xor ( n59969 , n59508 , n59566 );
and ( n59970 , n30364 , n59702 );
and ( n59971 , n59969 , n59970 );
xor ( n59972 , n59969 , n59970 );
xor ( n59973 , n59512 , n59564 );
and ( n59974 , n30369 , n59702 );
and ( n59975 , n59973 , n59974 );
xor ( n59976 , n59973 , n59974 );
xor ( n59977 , n59516 , n59562 );
and ( n59978 , n30374 , n59702 );
and ( n59979 , n59977 , n59978 );
xor ( n59980 , n59977 , n59978 );
xor ( n59981 , n59520 , n59560 );
and ( n59982 , n30379 , n59702 );
and ( n59983 , n59981 , n59982 );
xor ( n59984 , n59981 , n59982 );
xor ( n59985 , n59524 , n59558 );
and ( n59986 , n30384 , n59702 );
and ( n59987 , n59985 , n59986 );
xor ( n59988 , n59985 , n59986 );
xor ( n59989 , n59528 , n59556 );
and ( n59990 , n30389 , n59702 );
and ( n59991 , n59989 , n59990 );
xor ( n59992 , n59989 , n59990 );
xor ( n59993 , n59532 , n59554 );
and ( n59994 , n30394 , n59702 );
and ( n59995 , n59993 , n59994 );
xor ( n59996 , n59993 , n59994 );
xor ( n59997 , n59536 , n59552 );
and ( n59998 , n30399 , n59702 );
and ( n59999 , n59997 , n59998 );
xor ( n60000 , n59997 , n59998 );
xor ( n60001 , n59540 , n59550 );
and ( n60002 , n30404 , n59702 );
and ( n60003 , n60001 , n60002 );
xor ( n60004 , n60001 , n60002 );
xor ( n60005 , n59544 , n59548 );
and ( n60006 , n30409 , n59702 );
and ( n60007 , n60005 , n60006 );
buf ( n60008 , n60007 );
and ( n60009 , n60004 , n60008 );
or ( n60010 , n60003 , n60009 );
and ( n60011 , n60000 , n60010 );
or ( n60012 , n59999 , n60011 );
and ( n60013 , n59996 , n60012 );
or ( n60014 , n59995 , n60013 );
and ( n60015 , n59992 , n60014 );
or ( n60016 , n59991 , n60015 );
and ( n60017 , n59988 , n60016 );
or ( n60018 , n59987 , n60017 );
and ( n60019 , n59984 , n60018 );
or ( n60020 , n59983 , n60019 );
and ( n60021 , n59980 , n60020 );
or ( n60022 , n59979 , n60021 );
and ( n60023 , n59976 , n60022 );
or ( n60024 , n59975 , n60023 );
and ( n60025 , n59972 , n60024 );
or ( n60026 , n59971 , n60025 );
and ( n60027 , n59968 , n60026 );
or ( n60028 , n59967 , n60027 );
and ( n60029 , n59964 , n60028 );
or ( n60030 , n59963 , n60029 );
and ( n60031 , n59960 , n60030 );
or ( n60032 , n59959 , n60031 );
and ( n60033 , n59956 , n60032 );
or ( n60034 , n59955 , n60033 );
and ( n60035 , n59952 , n60034 );
or ( n60036 , n59951 , n60035 );
and ( n60037 , n59948 , n60036 );
or ( n60038 , n59947 , n60037 );
and ( n60039 , n59944 , n60038 );
or ( n60040 , n59943 , n60039 );
and ( n60041 , n59940 , n60040 );
or ( n60042 , n59939 , n60041 );
and ( n60043 , n59936 , n60042 );
or ( n60044 , n59935 , n60043 );
and ( n60045 , n59932 , n60044 );
or ( n60046 , n59931 , n60045 );
and ( n60047 , n59928 , n60046 );
or ( n60048 , n59927 , n60047 );
and ( n60049 , n59924 , n60048 );
or ( n60050 , n59923 , n60049 );
and ( n60051 , n59920 , n60050 );
or ( n60052 , n59919 , n60051 );
and ( n60053 , n59916 , n60052 );
or ( n60054 , n59915 , n60053 );
and ( n60055 , n59912 , n60054 );
or ( n60056 , n59911 , n60055 );
and ( n60057 , n59908 , n60056 );
or ( n60058 , n59907 , n60057 );
and ( n60059 , n59904 , n60058 );
or ( n60060 , n59903 , n60059 );
and ( n60061 , n59900 , n60060 );
or ( n60062 , n59899 , n60061 );
and ( n60063 , n59896 , n60062 );
or ( n60064 , n59895 , n60063 );
and ( n60065 , n59892 , n60064 );
or ( n60066 , n59891 , n60065 );
and ( n60067 , n59888 , n60066 );
or ( n60068 , n59887 , n60067 );
and ( n60069 , n59884 , n60068 );
or ( n60070 , n59883 , n60069 );
and ( n60071 , n59880 , n60070 );
or ( n60072 , n59879 , n60071 );
and ( n60073 , n59876 , n60072 );
or ( n60074 , n59875 , n60073 );
and ( n60075 , n59872 , n60074 );
or ( n60076 , n59871 , n60075 );
and ( n60077 , n59868 , n60076 );
or ( n60078 , n59867 , n60077 );
and ( n60079 , n59864 , n60078 );
or ( n60080 , n59863 , n60079 );
and ( n60081 , n59860 , n60080 );
or ( n60082 , n59859 , n60081 );
and ( n60083 , n59856 , n60082 );
or ( n60084 , n59855 , n60083 );
and ( n60085 , n59852 , n60084 );
or ( n60086 , n59851 , n60085 );
and ( n60087 , n59848 , n60086 );
or ( n60088 , n59847 , n60087 );
and ( n60089 , n59844 , n60088 );
or ( n60090 , n59843 , n60089 );
and ( n60091 , n59840 , n60090 );
or ( n60092 , n59839 , n60091 );
and ( n60093 , n59836 , n60092 );
or ( n60094 , n59835 , n60093 );
and ( n60095 , n59832 , n60094 );
or ( n60096 , n59831 , n60095 );
and ( n60097 , n59828 , n60096 );
or ( n60098 , n59827 , n60097 );
and ( n60099 , n59824 , n60098 );
or ( n60100 , n59823 , n60099 );
and ( n60101 , n59820 , n60100 );
or ( n60102 , n59819 , n60101 );
and ( n60103 , n59816 , n60102 );
or ( n60104 , n59815 , n60103 );
and ( n60105 , n59812 , n60104 );
or ( n60106 , n59811 , n60105 );
and ( n60107 , n59808 , n60106 );
or ( n60108 , n59807 , n60107 );
and ( n60109 , n59804 , n60108 );
or ( n60110 , n59803 , n60109 );
and ( n60111 , n59800 , n60110 );
or ( n60112 , n59799 , n60111 );
and ( n60113 , n59796 , n60112 );
or ( n60114 , n59795 , n60113 );
and ( n60115 , n59792 , n60114 );
or ( n60116 , n59791 , n60115 );
and ( n60117 , n59788 , n60116 );
or ( n60118 , n59787 , n60117 );
and ( n60119 , n59784 , n60118 );
or ( n60120 , n59783 , n60119 );
and ( n60121 , n59780 , n60120 );
or ( n60122 , n59779 , n60121 );
and ( n60123 , n59776 , n60122 );
or ( n60124 , n59775 , n60123 );
and ( n60125 , n59772 , n60124 );
or ( n60126 , n59771 , n60125 );
and ( n60127 , n59768 , n60126 );
or ( n60128 , n59767 , n60127 );
and ( n60129 , n59764 , n60128 );
or ( n60130 , n59763 , n60129 );
and ( n60131 , n59760 , n60130 );
or ( n60132 , n59759 , n60131 );
and ( n60133 , n59756 , n60132 );
or ( n60134 , n59755 , n60133 );
and ( n60135 , n59752 , n60134 );
or ( n60136 , n59751 , n60135 );
and ( n60137 , n59748 , n60136 );
or ( n60138 , n59747 , n60137 );
and ( n60139 , n59744 , n60138 );
or ( n60140 , n59743 , n60139 );
and ( n60141 , n59740 , n60140 );
or ( n60142 , n59739 , n60141 );
and ( n60143 , n59736 , n60142 );
or ( n60144 , n59735 , n60143 );
and ( n60145 , n59732 , n60144 );
or ( n60146 , n59731 , n60145 );
and ( n60147 , n59728 , n60146 );
or ( n60148 , n59727 , n60147 );
and ( n60149 , n59724 , n60148 );
or ( n60150 , n59723 , n60149 );
and ( n60151 , n59720 , n60150 );
or ( n60152 , n59719 , n60151 );
and ( n60153 , n59716 , n60152 );
or ( n60154 , n59715 , n60153 );
and ( n60155 , n59712 , n60154 );
or ( n60156 , n59711 , n60155 );
and ( n60157 , n59708 , n60156 );
or ( n60158 , n59707 , n60157 );
xor ( n60159 , n59704 , n60158 );
buf ( n60160 , n18004 );
and ( n60161 , n30034 , n60160 );
xor ( n60162 , n60159 , n60161 );
xor ( n60163 , n59708 , n60156 );
and ( n60164 , n30039 , n60160 );
and ( n60165 , n60163 , n60164 );
xor ( n60166 , n60163 , n60164 );
xor ( n60167 , n59712 , n60154 );
and ( n60168 , n30044 , n60160 );
and ( n60169 , n60167 , n60168 );
xor ( n60170 , n60167 , n60168 );
xor ( n60171 , n59716 , n60152 );
and ( n60172 , n30049 , n60160 );
and ( n60173 , n60171 , n60172 );
xor ( n60174 , n60171 , n60172 );
xor ( n60175 , n59720 , n60150 );
and ( n60176 , n30054 , n60160 );
and ( n60177 , n60175 , n60176 );
xor ( n60178 , n60175 , n60176 );
xor ( n60179 , n59724 , n60148 );
and ( n60180 , n30059 , n60160 );
and ( n60181 , n60179 , n60180 );
xor ( n60182 , n60179 , n60180 );
xor ( n60183 , n59728 , n60146 );
and ( n60184 , n30064 , n60160 );
and ( n60185 , n60183 , n60184 );
xor ( n60186 , n60183 , n60184 );
xor ( n60187 , n59732 , n60144 );
and ( n60188 , n30069 , n60160 );
and ( n60189 , n60187 , n60188 );
xor ( n60190 , n60187 , n60188 );
xor ( n60191 , n59736 , n60142 );
and ( n60192 , n30074 , n60160 );
and ( n60193 , n60191 , n60192 );
xor ( n60194 , n60191 , n60192 );
xor ( n60195 , n59740 , n60140 );
and ( n60196 , n30079 , n60160 );
and ( n60197 , n60195 , n60196 );
xor ( n60198 , n60195 , n60196 );
xor ( n60199 , n59744 , n60138 );
and ( n60200 , n30084 , n60160 );
and ( n60201 , n60199 , n60200 );
xor ( n60202 , n60199 , n60200 );
xor ( n60203 , n59748 , n60136 );
and ( n60204 , n30089 , n60160 );
and ( n60205 , n60203 , n60204 );
xor ( n60206 , n60203 , n60204 );
xor ( n60207 , n59752 , n60134 );
and ( n60208 , n30094 , n60160 );
and ( n60209 , n60207 , n60208 );
xor ( n60210 , n60207 , n60208 );
xor ( n60211 , n59756 , n60132 );
and ( n60212 , n30099 , n60160 );
and ( n60213 , n60211 , n60212 );
xor ( n60214 , n60211 , n60212 );
xor ( n60215 , n59760 , n60130 );
and ( n60216 , n30104 , n60160 );
and ( n60217 , n60215 , n60216 );
xor ( n60218 , n60215 , n60216 );
xor ( n60219 , n59764 , n60128 );
and ( n60220 , n30109 , n60160 );
and ( n60221 , n60219 , n60220 );
xor ( n60222 , n60219 , n60220 );
xor ( n60223 , n59768 , n60126 );
and ( n60224 , n30114 , n60160 );
and ( n60225 , n60223 , n60224 );
xor ( n60226 , n60223 , n60224 );
xor ( n60227 , n59772 , n60124 );
and ( n60228 , n30119 , n60160 );
and ( n60229 , n60227 , n60228 );
xor ( n60230 , n60227 , n60228 );
xor ( n60231 , n59776 , n60122 );
and ( n60232 , n30124 , n60160 );
and ( n60233 , n60231 , n60232 );
xor ( n60234 , n60231 , n60232 );
xor ( n60235 , n59780 , n60120 );
and ( n60236 , n30129 , n60160 );
and ( n60237 , n60235 , n60236 );
xor ( n60238 , n60235 , n60236 );
xor ( n60239 , n59784 , n60118 );
and ( n60240 , n30134 , n60160 );
and ( n60241 , n60239 , n60240 );
xor ( n60242 , n60239 , n60240 );
xor ( n60243 , n59788 , n60116 );
and ( n60244 , n30139 , n60160 );
and ( n60245 , n60243 , n60244 );
xor ( n60246 , n60243 , n60244 );
xor ( n60247 , n59792 , n60114 );
and ( n60248 , n30144 , n60160 );
and ( n60249 , n60247 , n60248 );
xor ( n60250 , n60247 , n60248 );
xor ( n60251 , n59796 , n60112 );
and ( n60252 , n30149 , n60160 );
and ( n60253 , n60251 , n60252 );
xor ( n60254 , n60251 , n60252 );
xor ( n60255 , n59800 , n60110 );
and ( n60256 , n30154 , n60160 );
and ( n60257 , n60255 , n60256 );
xor ( n60258 , n60255 , n60256 );
xor ( n60259 , n59804 , n60108 );
and ( n60260 , n30159 , n60160 );
and ( n60261 , n60259 , n60260 );
xor ( n60262 , n60259 , n60260 );
xor ( n60263 , n59808 , n60106 );
and ( n60264 , n30164 , n60160 );
and ( n60265 , n60263 , n60264 );
xor ( n60266 , n60263 , n60264 );
xor ( n60267 , n59812 , n60104 );
and ( n60268 , n30169 , n60160 );
and ( n60269 , n60267 , n60268 );
xor ( n60270 , n60267 , n60268 );
xor ( n60271 , n59816 , n60102 );
and ( n60272 , n30174 , n60160 );
and ( n60273 , n60271 , n60272 );
xor ( n60274 , n60271 , n60272 );
xor ( n60275 , n59820 , n60100 );
and ( n60276 , n30179 , n60160 );
and ( n60277 , n60275 , n60276 );
xor ( n60278 , n60275 , n60276 );
xor ( n60279 , n59824 , n60098 );
and ( n60280 , n30184 , n60160 );
and ( n60281 , n60279 , n60280 );
xor ( n60282 , n60279 , n60280 );
xor ( n60283 , n59828 , n60096 );
and ( n60284 , n30189 , n60160 );
and ( n60285 , n60283 , n60284 );
xor ( n60286 , n60283 , n60284 );
xor ( n60287 , n59832 , n60094 );
and ( n60288 , n30194 , n60160 );
and ( n60289 , n60287 , n60288 );
xor ( n60290 , n60287 , n60288 );
xor ( n60291 , n59836 , n60092 );
and ( n60292 , n30199 , n60160 );
and ( n60293 , n60291 , n60292 );
xor ( n60294 , n60291 , n60292 );
xor ( n60295 , n59840 , n60090 );
and ( n60296 , n30204 , n60160 );
and ( n60297 , n60295 , n60296 );
xor ( n60298 , n60295 , n60296 );
xor ( n60299 , n59844 , n60088 );
and ( n60300 , n30209 , n60160 );
and ( n60301 , n60299 , n60300 );
xor ( n60302 , n60299 , n60300 );
xor ( n60303 , n59848 , n60086 );
and ( n60304 , n30214 , n60160 );
and ( n60305 , n60303 , n60304 );
xor ( n60306 , n60303 , n60304 );
xor ( n60307 , n59852 , n60084 );
and ( n60308 , n30219 , n60160 );
and ( n60309 , n60307 , n60308 );
xor ( n60310 , n60307 , n60308 );
xor ( n60311 , n59856 , n60082 );
and ( n60312 , n30224 , n60160 );
and ( n60313 , n60311 , n60312 );
xor ( n60314 , n60311 , n60312 );
xor ( n60315 , n59860 , n60080 );
and ( n60316 , n30229 , n60160 );
and ( n60317 , n60315 , n60316 );
xor ( n60318 , n60315 , n60316 );
xor ( n60319 , n59864 , n60078 );
and ( n60320 , n30234 , n60160 );
and ( n60321 , n60319 , n60320 );
xor ( n60322 , n60319 , n60320 );
xor ( n60323 , n59868 , n60076 );
and ( n60324 , n30239 , n60160 );
and ( n60325 , n60323 , n60324 );
xor ( n60326 , n60323 , n60324 );
xor ( n60327 , n59872 , n60074 );
and ( n60328 , n30244 , n60160 );
and ( n60329 , n60327 , n60328 );
xor ( n60330 , n60327 , n60328 );
xor ( n60331 , n59876 , n60072 );
and ( n60332 , n30249 , n60160 );
and ( n60333 , n60331 , n60332 );
xor ( n60334 , n60331 , n60332 );
xor ( n60335 , n59880 , n60070 );
and ( n60336 , n30254 , n60160 );
and ( n60337 , n60335 , n60336 );
xor ( n60338 , n60335 , n60336 );
xor ( n60339 , n59884 , n60068 );
and ( n60340 , n30259 , n60160 );
and ( n60341 , n60339 , n60340 );
xor ( n60342 , n60339 , n60340 );
xor ( n60343 , n59888 , n60066 );
and ( n60344 , n30264 , n60160 );
and ( n60345 , n60343 , n60344 );
xor ( n60346 , n60343 , n60344 );
xor ( n60347 , n59892 , n60064 );
and ( n60348 , n30269 , n60160 );
and ( n60349 , n60347 , n60348 );
xor ( n60350 , n60347 , n60348 );
xor ( n60351 , n59896 , n60062 );
and ( n60352 , n30274 , n60160 );
and ( n60353 , n60351 , n60352 );
xor ( n60354 , n60351 , n60352 );
xor ( n60355 , n59900 , n60060 );
and ( n60356 , n30279 , n60160 );
and ( n60357 , n60355 , n60356 );
xor ( n60358 , n60355 , n60356 );
xor ( n60359 , n59904 , n60058 );
and ( n60360 , n30284 , n60160 );
and ( n60361 , n60359 , n60360 );
xor ( n60362 , n60359 , n60360 );
xor ( n60363 , n59908 , n60056 );
and ( n60364 , n30289 , n60160 );
and ( n60365 , n60363 , n60364 );
xor ( n60366 , n60363 , n60364 );
xor ( n60367 , n59912 , n60054 );
and ( n60368 , n30294 , n60160 );
and ( n60369 , n60367 , n60368 );
xor ( n60370 , n60367 , n60368 );
xor ( n60371 , n59916 , n60052 );
and ( n60372 , n30299 , n60160 );
and ( n60373 , n60371 , n60372 );
xor ( n60374 , n60371 , n60372 );
xor ( n60375 , n59920 , n60050 );
and ( n60376 , n30304 , n60160 );
and ( n60377 , n60375 , n60376 );
xor ( n60378 , n60375 , n60376 );
xor ( n60379 , n59924 , n60048 );
and ( n60380 , n30309 , n60160 );
and ( n60381 , n60379 , n60380 );
xor ( n60382 , n60379 , n60380 );
xor ( n60383 , n59928 , n60046 );
and ( n60384 , n30314 , n60160 );
and ( n60385 , n60383 , n60384 );
xor ( n60386 , n60383 , n60384 );
xor ( n60387 , n59932 , n60044 );
and ( n60388 , n30319 , n60160 );
and ( n60389 , n60387 , n60388 );
xor ( n60390 , n60387 , n60388 );
xor ( n60391 , n59936 , n60042 );
and ( n60392 , n30324 , n60160 );
and ( n60393 , n60391 , n60392 );
xor ( n60394 , n60391 , n60392 );
xor ( n60395 , n59940 , n60040 );
and ( n60396 , n30329 , n60160 );
and ( n60397 , n60395 , n60396 );
xor ( n60398 , n60395 , n60396 );
xor ( n60399 , n59944 , n60038 );
and ( n60400 , n30334 , n60160 );
and ( n60401 , n60399 , n60400 );
xor ( n60402 , n60399 , n60400 );
xor ( n60403 , n59948 , n60036 );
and ( n60404 , n30339 , n60160 );
and ( n60405 , n60403 , n60404 );
xor ( n60406 , n60403 , n60404 );
xor ( n60407 , n59952 , n60034 );
and ( n60408 , n30344 , n60160 );
and ( n60409 , n60407 , n60408 );
xor ( n60410 , n60407 , n60408 );
xor ( n60411 , n59956 , n60032 );
and ( n60412 , n30349 , n60160 );
and ( n60413 , n60411 , n60412 );
xor ( n60414 , n60411 , n60412 );
xor ( n60415 , n59960 , n60030 );
and ( n60416 , n30354 , n60160 );
and ( n60417 , n60415 , n60416 );
xor ( n60418 , n60415 , n60416 );
xor ( n60419 , n59964 , n60028 );
and ( n60420 , n30359 , n60160 );
and ( n60421 , n60419 , n60420 );
xor ( n60422 , n60419 , n60420 );
xor ( n60423 , n59968 , n60026 );
and ( n60424 , n30364 , n60160 );
and ( n60425 , n60423 , n60424 );
xor ( n60426 , n60423 , n60424 );
xor ( n60427 , n59972 , n60024 );
and ( n60428 , n30369 , n60160 );
and ( n60429 , n60427 , n60428 );
xor ( n60430 , n60427 , n60428 );
xor ( n60431 , n59976 , n60022 );
and ( n60432 , n30374 , n60160 );
and ( n60433 , n60431 , n60432 );
xor ( n60434 , n60431 , n60432 );
xor ( n60435 , n59980 , n60020 );
and ( n60436 , n30379 , n60160 );
and ( n60437 , n60435 , n60436 );
xor ( n60438 , n60435 , n60436 );
xor ( n60439 , n59984 , n60018 );
and ( n60440 , n30384 , n60160 );
and ( n60441 , n60439 , n60440 );
xor ( n60442 , n60439 , n60440 );
xor ( n60443 , n59988 , n60016 );
and ( n60444 , n30389 , n60160 );
and ( n60445 , n60443 , n60444 );
xor ( n60446 , n60443 , n60444 );
xor ( n60447 , n59992 , n60014 );
and ( n60448 , n30394 , n60160 );
and ( n60449 , n60447 , n60448 );
xor ( n60450 , n60447 , n60448 );
xor ( n60451 , n59996 , n60012 );
and ( n60452 , n30399 , n60160 );
and ( n60453 , n60451 , n60452 );
xor ( n60454 , n60451 , n60452 );
xor ( n60455 , n60000 , n60010 );
and ( n60456 , n30404 , n60160 );
and ( n60457 , n60455 , n60456 );
xor ( n60458 , n60455 , n60456 );
xor ( n60459 , n60004 , n60008 );
and ( n60460 , n30409 , n60160 );
and ( n60461 , n60459 , n60460 );
buf ( n60462 , n60461 );
and ( n60463 , n60458 , n60462 );
or ( n60464 , n60457 , n60463 );
and ( n60465 , n60454 , n60464 );
or ( n60466 , n60453 , n60465 );
and ( n60467 , n60450 , n60466 );
or ( n60468 , n60449 , n60467 );
and ( n60469 , n60446 , n60468 );
or ( n60470 , n60445 , n60469 );
and ( n60471 , n60442 , n60470 );
or ( n60472 , n60441 , n60471 );
and ( n60473 , n60438 , n60472 );
or ( n60474 , n60437 , n60473 );
and ( n60475 , n60434 , n60474 );
or ( n60476 , n60433 , n60475 );
and ( n60477 , n60430 , n60476 );
or ( n60478 , n60429 , n60477 );
and ( n60479 , n60426 , n60478 );
or ( n60480 , n60425 , n60479 );
and ( n60481 , n60422 , n60480 );
or ( n60482 , n60421 , n60481 );
and ( n60483 , n60418 , n60482 );
or ( n60484 , n60417 , n60483 );
and ( n60485 , n60414 , n60484 );
or ( n60486 , n60413 , n60485 );
and ( n60487 , n60410 , n60486 );
or ( n60488 , n60409 , n60487 );
and ( n60489 , n60406 , n60488 );
or ( n60490 , n60405 , n60489 );
and ( n60491 , n60402 , n60490 );
or ( n60492 , n60401 , n60491 );
and ( n60493 , n60398 , n60492 );
or ( n60494 , n60397 , n60493 );
and ( n60495 , n60394 , n60494 );
or ( n60496 , n60393 , n60495 );
and ( n60497 , n60390 , n60496 );
or ( n60498 , n60389 , n60497 );
and ( n60499 , n60386 , n60498 );
or ( n60500 , n60385 , n60499 );
and ( n60501 , n60382 , n60500 );
or ( n60502 , n60381 , n60501 );
and ( n60503 , n60378 , n60502 );
or ( n60504 , n60377 , n60503 );
and ( n60505 , n60374 , n60504 );
or ( n60506 , n60373 , n60505 );
and ( n60507 , n60370 , n60506 );
or ( n60508 , n60369 , n60507 );
and ( n60509 , n60366 , n60508 );
or ( n60510 , n60365 , n60509 );
and ( n60511 , n60362 , n60510 );
or ( n60512 , n60361 , n60511 );
and ( n60513 , n60358 , n60512 );
or ( n60514 , n60357 , n60513 );
and ( n60515 , n60354 , n60514 );
or ( n60516 , n60353 , n60515 );
and ( n60517 , n60350 , n60516 );
or ( n60518 , n60349 , n60517 );
and ( n60519 , n60346 , n60518 );
or ( n60520 , n60345 , n60519 );
and ( n60521 , n60342 , n60520 );
or ( n60522 , n60341 , n60521 );
and ( n60523 , n60338 , n60522 );
or ( n60524 , n60337 , n60523 );
and ( n60525 , n60334 , n60524 );
or ( n60526 , n60333 , n60525 );
and ( n60527 , n60330 , n60526 );
or ( n60528 , n60329 , n60527 );
and ( n60529 , n60326 , n60528 );
or ( n60530 , n60325 , n60529 );
and ( n60531 , n60322 , n60530 );
or ( n60532 , n60321 , n60531 );
and ( n60533 , n60318 , n60532 );
or ( n60534 , n60317 , n60533 );
and ( n60535 , n60314 , n60534 );
or ( n60536 , n60313 , n60535 );
and ( n60537 , n60310 , n60536 );
or ( n60538 , n60309 , n60537 );
and ( n60539 , n60306 , n60538 );
or ( n60540 , n60305 , n60539 );
and ( n60541 , n60302 , n60540 );
or ( n60542 , n60301 , n60541 );
and ( n60543 , n60298 , n60542 );
or ( n60544 , n60297 , n60543 );
and ( n60545 , n60294 , n60544 );
or ( n60546 , n60293 , n60545 );
and ( n60547 , n60290 , n60546 );
or ( n60548 , n60289 , n60547 );
and ( n60549 , n60286 , n60548 );
or ( n60550 , n60285 , n60549 );
and ( n60551 , n60282 , n60550 );
or ( n60552 , n60281 , n60551 );
and ( n60553 , n60278 , n60552 );
or ( n60554 , n60277 , n60553 );
and ( n60555 , n60274 , n60554 );
or ( n60556 , n60273 , n60555 );
and ( n60557 , n60270 , n60556 );
or ( n60558 , n60269 , n60557 );
and ( n60559 , n60266 , n60558 );
or ( n60560 , n60265 , n60559 );
and ( n60561 , n60262 , n60560 );
or ( n60562 , n60261 , n60561 );
and ( n60563 , n60258 , n60562 );
or ( n60564 , n60257 , n60563 );
and ( n60565 , n60254 , n60564 );
or ( n60566 , n60253 , n60565 );
and ( n60567 , n60250 , n60566 );
or ( n60568 , n60249 , n60567 );
and ( n60569 , n60246 , n60568 );
or ( n60570 , n60245 , n60569 );
and ( n60571 , n60242 , n60570 );
or ( n60572 , n60241 , n60571 );
and ( n60573 , n60238 , n60572 );
or ( n60574 , n60237 , n60573 );
and ( n60575 , n60234 , n60574 );
or ( n60576 , n60233 , n60575 );
and ( n60577 , n60230 , n60576 );
or ( n60578 , n60229 , n60577 );
and ( n60579 , n60226 , n60578 );
or ( n60580 , n60225 , n60579 );
and ( n60581 , n60222 , n60580 );
or ( n60582 , n60221 , n60581 );
and ( n60583 , n60218 , n60582 );
or ( n60584 , n60217 , n60583 );
and ( n60585 , n60214 , n60584 );
or ( n60586 , n60213 , n60585 );
and ( n60587 , n60210 , n60586 );
or ( n60588 , n60209 , n60587 );
and ( n60589 , n60206 , n60588 );
or ( n60590 , n60205 , n60589 );
and ( n60591 , n60202 , n60590 );
or ( n60592 , n60201 , n60591 );
and ( n60593 , n60198 , n60592 );
or ( n60594 , n60197 , n60593 );
and ( n60595 , n60194 , n60594 );
or ( n60596 , n60193 , n60595 );
and ( n60597 , n60190 , n60596 );
or ( n60598 , n60189 , n60597 );
and ( n60599 , n60186 , n60598 );
or ( n60600 , n60185 , n60599 );
and ( n60601 , n60182 , n60600 );
or ( n60602 , n60181 , n60601 );
and ( n60603 , n60178 , n60602 );
or ( n60604 , n60177 , n60603 );
and ( n60605 , n60174 , n60604 );
or ( n60606 , n60173 , n60605 );
and ( n60607 , n60170 , n60606 );
or ( n60608 , n60169 , n60607 );
and ( n60609 , n60166 , n60608 );
or ( n60610 , n60165 , n60609 );
xor ( n60611 , n60162 , n60610 );
buf ( n60612 , n18002 );
and ( n60613 , n30039 , n60612 );
xor ( n60614 , n60611 , n60613 );
xor ( n60615 , n60166 , n60608 );
and ( n60616 , n30044 , n60612 );
and ( n60617 , n60615 , n60616 );
xor ( n60618 , n60615 , n60616 );
xor ( n60619 , n60170 , n60606 );
and ( n60620 , n30049 , n60612 );
and ( n60621 , n60619 , n60620 );
xor ( n60622 , n60619 , n60620 );
xor ( n60623 , n60174 , n60604 );
and ( n60624 , n30054 , n60612 );
and ( n60625 , n60623 , n60624 );
xor ( n60626 , n60623 , n60624 );
xor ( n60627 , n60178 , n60602 );
and ( n60628 , n30059 , n60612 );
and ( n60629 , n60627 , n60628 );
xor ( n60630 , n60627 , n60628 );
xor ( n60631 , n60182 , n60600 );
and ( n60632 , n30064 , n60612 );
and ( n60633 , n60631 , n60632 );
xor ( n60634 , n60631 , n60632 );
xor ( n60635 , n60186 , n60598 );
and ( n60636 , n30069 , n60612 );
and ( n60637 , n60635 , n60636 );
xor ( n60638 , n60635 , n60636 );
xor ( n60639 , n60190 , n60596 );
and ( n60640 , n30074 , n60612 );
and ( n60641 , n60639 , n60640 );
xor ( n60642 , n60639 , n60640 );
xor ( n60643 , n60194 , n60594 );
and ( n60644 , n30079 , n60612 );
and ( n60645 , n60643 , n60644 );
xor ( n60646 , n60643 , n60644 );
xor ( n60647 , n60198 , n60592 );
and ( n60648 , n30084 , n60612 );
and ( n60649 , n60647 , n60648 );
xor ( n60650 , n60647 , n60648 );
xor ( n60651 , n60202 , n60590 );
and ( n60652 , n30089 , n60612 );
and ( n60653 , n60651 , n60652 );
xor ( n60654 , n60651 , n60652 );
xor ( n60655 , n60206 , n60588 );
and ( n60656 , n30094 , n60612 );
and ( n60657 , n60655 , n60656 );
xor ( n60658 , n60655 , n60656 );
xor ( n60659 , n60210 , n60586 );
and ( n60660 , n30099 , n60612 );
and ( n60661 , n60659 , n60660 );
xor ( n60662 , n60659 , n60660 );
xor ( n60663 , n60214 , n60584 );
and ( n60664 , n30104 , n60612 );
and ( n60665 , n60663 , n60664 );
xor ( n60666 , n60663 , n60664 );
xor ( n60667 , n60218 , n60582 );
and ( n60668 , n30109 , n60612 );
and ( n60669 , n60667 , n60668 );
xor ( n60670 , n60667 , n60668 );
xor ( n60671 , n60222 , n60580 );
and ( n60672 , n30114 , n60612 );
and ( n60673 , n60671 , n60672 );
xor ( n60674 , n60671 , n60672 );
xor ( n60675 , n60226 , n60578 );
and ( n60676 , n30119 , n60612 );
and ( n60677 , n60675 , n60676 );
xor ( n60678 , n60675 , n60676 );
xor ( n60679 , n60230 , n60576 );
and ( n60680 , n30124 , n60612 );
and ( n60681 , n60679 , n60680 );
xor ( n60682 , n60679 , n60680 );
xor ( n60683 , n60234 , n60574 );
and ( n60684 , n30129 , n60612 );
and ( n60685 , n60683 , n60684 );
xor ( n60686 , n60683 , n60684 );
xor ( n60687 , n60238 , n60572 );
and ( n60688 , n30134 , n60612 );
and ( n60689 , n60687 , n60688 );
xor ( n60690 , n60687 , n60688 );
xor ( n60691 , n60242 , n60570 );
and ( n60692 , n30139 , n60612 );
and ( n60693 , n60691 , n60692 );
xor ( n60694 , n60691 , n60692 );
xor ( n60695 , n60246 , n60568 );
and ( n60696 , n30144 , n60612 );
and ( n60697 , n60695 , n60696 );
xor ( n60698 , n60695 , n60696 );
xor ( n60699 , n60250 , n60566 );
and ( n60700 , n30149 , n60612 );
and ( n60701 , n60699 , n60700 );
xor ( n60702 , n60699 , n60700 );
xor ( n60703 , n60254 , n60564 );
and ( n60704 , n30154 , n60612 );
and ( n60705 , n60703 , n60704 );
xor ( n60706 , n60703 , n60704 );
xor ( n60707 , n60258 , n60562 );
and ( n60708 , n30159 , n60612 );
and ( n60709 , n60707 , n60708 );
xor ( n60710 , n60707 , n60708 );
xor ( n60711 , n60262 , n60560 );
and ( n60712 , n30164 , n60612 );
and ( n60713 , n60711 , n60712 );
xor ( n60714 , n60711 , n60712 );
xor ( n60715 , n60266 , n60558 );
and ( n60716 , n30169 , n60612 );
and ( n60717 , n60715 , n60716 );
xor ( n60718 , n60715 , n60716 );
xor ( n60719 , n60270 , n60556 );
and ( n60720 , n30174 , n60612 );
and ( n60721 , n60719 , n60720 );
xor ( n60722 , n60719 , n60720 );
xor ( n60723 , n60274 , n60554 );
and ( n60724 , n30179 , n60612 );
and ( n60725 , n60723 , n60724 );
xor ( n60726 , n60723 , n60724 );
xor ( n60727 , n60278 , n60552 );
and ( n60728 , n30184 , n60612 );
and ( n60729 , n60727 , n60728 );
xor ( n60730 , n60727 , n60728 );
xor ( n60731 , n60282 , n60550 );
and ( n60732 , n30189 , n60612 );
and ( n60733 , n60731 , n60732 );
xor ( n60734 , n60731 , n60732 );
xor ( n60735 , n60286 , n60548 );
and ( n60736 , n30194 , n60612 );
and ( n60737 , n60735 , n60736 );
xor ( n60738 , n60735 , n60736 );
xor ( n60739 , n60290 , n60546 );
and ( n60740 , n30199 , n60612 );
and ( n60741 , n60739 , n60740 );
xor ( n60742 , n60739 , n60740 );
xor ( n60743 , n60294 , n60544 );
and ( n60744 , n30204 , n60612 );
and ( n60745 , n60743 , n60744 );
xor ( n60746 , n60743 , n60744 );
xor ( n60747 , n60298 , n60542 );
and ( n60748 , n30209 , n60612 );
and ( n60749 , n60747 , n60748 );
xor ( n60750 , n60747 , n60748 );
xor ( n60751 , n60302 , n60540 );
and ( n60752 , n30214 , n60612 );
and ( n60753 , n60751 , n60752 );
xor ( n60754 , n60751 , n60752 );
xor ( n60755 , n60306 , n60538 );
and ( n60756 , n30219 , n60612 );
and ( n60757 , n60755 , n60756 );
xor ( n60758 , n60755 , n60756 );
xor ( n60759 , n60310 , n60536 );
and ( n60760 , n30224 , n60612 );
and ( n60761 , n60759 , n60760 );
xor ( n60762 , n60759 , n60760 );
xor ( n60763 , n60314 , n60534 );
and ( n60764 , n30229 , n60612 );
and ( n60765 , n60763 , n60764 );
xor ( n60766 , n60763 , n60764 );
xor ( n60767 , n60318 , n60532 );
and ( n60768 , n30234 , n60612 );
and ( n60769 , n60767 , n60768 );
xor ( n60770 , n60767 , n60768 );
xor ( n60771 , n60322 , n60530 );
and ( n60772 , n30239 , n60612 );
and ( n60773 , n60771 , n60772 );
xor ( n60774 , n60771 , n60772 );
xor ( n60775 , n60326 , n60528 );
and ( n60776 , n30244 , n60612 );
and ( n60777 , n60775 , n60776 );
xor ( n60778 , n60775 , n60776 );
xor ( n60779 , n60330 , n60526 );
and ( n60780 , n30249 , n60612 );
and ( n60781 , n60779 , n60780 );
xor ( n60782 , n60779 , n60780 );
xor ( n60783 , n60334 , n60524 );
and ( n60784 , n30254 , n60612 );
and ( n60785 , n60783 , n60784 );
xor ( n60786 , n60783 , n60784 );
xor ( n60787 , n60338 , n60522 );
and ( n60788 , n30259 , n60612 );
and ( n60789 , n60787 , n60788 );
xor ( n60790 , n60787 , n60788 );
xor ( n60791 , n60342 , n60520 );
and ( n60792 , n30264 , n60612 );
and ( n60793 , n60791 , n60792 );
xor ( n60794 , n60791 , n60792 );
xor ( n60795 , n60346 , n60518 );
and ( n60796 , n30269 , n60612 );
and ( n60797 , n60795 , n60796 );
xor ( n60798 , n60795 , n60796 );
xor ( n60799 , n60350 , n60516 );
and ( n60800 , n30274 , n60612 );
and ( n60801 , n60799 , n60800 );
xor ( n60802 , n60799 , n60800 );
xor ( n60803 , n60354 , n60514 );
and ( n60804 , n30279 , n60612 );
and ( n60805 , n60803 , n60804 );
xor ( n60806 , n60803 , n60804 );
xor ( n60807 , n60358 , n60512 );
and ( n60808 , n30284 , n60612 );
and ( n60809 , n60807 , n60808 );
xor ( n60810 , n60807 , n60808 );
xor ( n60811 , n60362 , n60510 );
and ( n60812 , n30289 , n60612 );
and ( n60813 , n60811 , n60812 );
xor ( n60814 , n60811 , n60812 );
xor ( n60815 , n60366 , n60508 );
and ( n60816 , n30294 , n60612 );
and ( n60817 , n60815 , n60816 );
xor ( n60818 , n60815 , n60816 );
xor ( n60819 , n60370 , n60506 );
and ( n60820 , n30299 , n60612 );
and ( n60821 , n60819 , n60820 );
xor ( n60822 , n60819 , n60820 );
xor ( n60823 , n60374 , n60504 );
and ( n60824 , n30304 , n60612 );
and ( n60825 , n60823 , n60824 );
xor ( n60826 , n60823 , n60824 );
xor ( n60827 , n60378 , n60502 );
and ( n60828 , n30309 , n60612 );
and ( n60829 , n60827 , n60828 );
xor ( n60830 , n60827 , n60828 );
xor ( n60831 , n60382 , n60500 );
and ( n60832 , n30314 , n60612 );
and ( n60833 , n60831 , n60832 );
xor ( n60834 , n60831 , n60832 );
xor ( n60835 , n60386 , n60498 );
and ( n60836 , n30319 , n60612 );
and ( n60837 , n60835 , n60836 );
xor ( n60838 , n60835 , n60836 );
xor ( n60839 , n60390 , n60496 );
and ( n60840 , n30324 , n60612 );
and ( n60841 , n60839 , n60840 );
xor ( n60842 , n60839 , n60840 );
xor ( n60843 , n60394 , n60494 );
and ( n60844 , n30329 , n60612 );
and ( n60845 , n60843 , n60844 );
xor ( n60846 , n60843 , n60844 );
xor ( n60847 , n60398 , n60492 );
and ( n60848 , n30334 , n60612 );
and ( n60849 , n60847 , n60848 );
xor ( n60850 , n60847 , n60848 );
xor ( n60851 , n60402 , n60490 );
and ( n60852 , n30339 , n60612 );
and ( n60853 , n60851 , n60852 );
xor ( n60854 , n60851 , n60852 );
xor ( n60855 , n60406 , n60488 );
and ( n60856 , n30344 , n60612 );
and ( n60857 , n60855 , n60856 );
xor ( n60858 , n60855 , n60856 );
xor ( n60859 , n60410 , n60486 );
and ( n60860 , n30349 , n60612 );
and ( n60861 , n60859 , n60860 );
xor ( n60862 , n60859 , n60860 );
xor ( n60863 , n60414 , n60484 );
and ( n60864 , n30354 , n60612 );
and ( n60865 , n60863 , n60864 );
xor ( n60866 , n60863 , n60864 );
xor ( n60867 , n60418 , n60482 );
and ( n60868 , n30359 , n60612 );
and ( n60869 , n60867 , n60868 );
xor ( n60870 , n60867 , n60868 );
xor ( n60871 , n60422 , n60480 );
and ( n60872 , n30364 , n60612 );
and ( n60873 , n60871 , n60872 );
xor ( n60874 , n60871 , n60872 );
xor ( n60875 , n60426 , n60478 );
and ( n60876 , n30369 , n60612 );
and ( n60877 , n60875 , n60876 );
xor ( n60878 , n60875 , n60876 );
xor ( n60879 , n60430 , n60476 );
and ( n60880 , n30374 , n60612 );
and ( n60881 , n60879 , n60880 );
xor ( n60882 , n60879 , n60880 );
xor ( n60883 , n60434 , n60474 );
and ( n60884 , n30379 , n60612 );
and ( n60885 , n60883 , n60884 );
xor ( n60886 , n60883 , n60884 );
xor ( n60887 , n60438 , n60472 );
and ( n60888 , n30384 , n60612 );
and ( n60889 , n60887 , n60888 );
xor ( n60890 , n60887 , n60888 );
xor ( n60891 , n60442 , n60470 );
and ( n60892 , n30389 , n60612 );
and ( n60893 , n60891 , n60892 );
xor ( n60894 , n60891 , n60892 );
xor ( n60895 , n60446 , n60468 );
and ( n60896 , n30394 , n60612 );
and ( n60897 , n60895 , n60896 );
xor ( n60898 , n60895 , n60896 );
xor ( n60899 , n60450 , n60466 );
and ( n60900 , n30399 , n60612 );
and ( n60901 , n60899 , n60900 );
xor ( n60902 , n60899 , n60900 );
xor ( n60903 , n60454 , n60464 );
and ( n60904 , n30404 , n60612 );
and ( n60905 , n60903 , n60904 );
xor ( n60906 , n60903 , n60904 );
xor ( n60907 , n60458 , n60462 );
and ( n60908 , n30409 , n60612 );
and ( n60909 , n60907 , n60908 );
buf ( n60910 , n60909 );
and ( n60911 , n60906 , n60910 );
or ( n60912 , n60905 , n60911 );
and ( n60913 , n60902 , n60912 );
or ( n60914 , n60901 , n60913 );
and ( n60915 , n60898 , n60914 );
or ( n60916 , n60897 , n60915 );
and ( n60917 , n60894 , n60916 );
or ( n60918 , n60893 , n60917 );
and ( n60919 , n60890 , n60918 );
or ( n60920 , n60889 , n60919 );
and ( n60921 , n60886 , n60920 );
or ( n60922 , n60885 , n60921 );
and ( n60923 , n60882 , n60922 );
or ( n60924 , n60881 , n60923 );
and ( n60925 , n60878 , n60924 );
or ( n60926 , n60877 , n60925 );
and ( n60927 , n60874 , n60926 );
or ( n60928 , n60873 , n60927 );
and ( n60929 , n60870 , n60928 );
or ( n60930 , n60869 , n60929 );
and ( n60931 , n60866 , n60930 );
or ( n60932 , n60865 , n60931 );
and ( n60933 , n60862 , n60932 );
or ( n60934 , n60861 , n60933 );
and ( n60935 , n60858 , n60934 );
or ( n60936 , n60857 , n60935 );
and ( n60937 , n60854 , n60936 );
or ( n60938 , n60853 , n60937 );
and ( n60939 , n60850 , n60938 );
or ( n60940 , n60849 , n60939 );
and ( n60941 , n60846 , n60940 );
or ( n60942 , n60845 , n60941 );
and ( n60943 , n60842 , n60942 );
or ( n60944 , n60841 , n60943 );
and ( n60945 , n60838 , n60944 );
or ( n60946 , n60837 , n60945 );
and ( n60947 , n60834 , n60946 );
or ( n60948 , n60833 , n60947 );
and ( n60949 , n60830 , n60948 );
or ( n60950 , n60829 , n60949 );
and ( n60951 , n60826 , n60950 );
or ( n60952 , n60825 , n60951 );
and ( n60953 , n60822 , n60952 );
or ( n60954 , n60821 , n60953 );
and ( n60955 , n60818 , n60954 );
or ( n60956 , n60817 , n60955 );
and ( n60957 , n60814 , n60956 );
or ( n60958 , n60813 , n60957 );
and ( n60959 , n60810 , n60958 );
or ( n60960 , n60809 , n60959 );
and ( n60961 , n60806 , n60960 );
or ( n60962 , n60805 , n60961 );
and ( n60963 , n60802 , n60962 );
or ( n60964 , n60801 , n60963 );
and ( n60965 , n60798 , n60964 );
or ( n60966 , n60797 , n60965 );
and ( n60967 , n60794 , n60966 );
or ( n60968 , n60793 , n60967 );
and ( n60969 , n60790 , n60968 );
or ( n60970 , n60789 , n60969 );
and ( n60971 , n60786 , n60970 );
or ( n60972 , n60785 , n60971 );
and ( n60973 , n60782 , n60972 );
or ( n60974 , n60781 , n60973 );
and ( n60975 , n60778 , n60974 );
or ( n60976 , n60777 , n60975 );
and ( n60977 , n60774 , n60976 );
or ( n60978 , n60773 , n60977 );
and ( n60979 , n60770 , n60978 );
or ( n60980 , n60769 , n60979 );
and ( n60981 , n60766 , n60980 );
or ( n60982 , n60765 , n60981 );
and ( n60983 , n60762 , n60982 );
or ( n60984 , n60761 , n60983 );
and ( n60985 , n60758 , n60984 );
or ( n60986 , n60757 , n60985 );
and ( n60987 , n60754 , n60986 );
or ( n60988 , n60753 , n60987 );
and ( n60989 , n60750 , n60988 );
or ( n60990 , n60749 , n60989 );
and ( n60991 , n60746 , n60990 );
or ( n60992 , n60745 , n60991 );
and ( n60993 , n60742 , n60992 );
or ( n60994 , n60741 , n60993 );
and ( n60995 , n60738 , n60994 );
or ( n60996 , n60737 , n60995 );
and ( n60997 , n60734 , n60996 );
or ( n60998 , n60733 , n60997 );
and ( n60999 , n60730 , n60998 );
or ( n61000 , n60729 , n60999 );
and ( n61001 , n60726 , n61000 );
or ( n61002 , n60725 , n61001 );
and ( n61003 , n60722 , n61002 );
or ( n61004 , n60721 , n61003 );
and ( n61005 , n60718 , n61004 );
or ( n61006 , n60717 , n61005 );
and ( n61007 , n60714 , n61006 );
or ( n61008 , n60713 , n61007 );
and ( n61009 , n60710 , n61008 );
or ( n61010 , n60709 , n61009 );
and ( n61011 , n60706 , n61010 );
or ( n61012 , n60705 , n61011 );
and ( n61013 , n60702 , n61012 );
or ( n61014 , n60701 , n61013 );
and ( n61015 , n60698 , n61014 );
or ( n61016 , n60697 , n61015 );
and ( n61017 , n60694 , n61016 );
or ( n61018 , n60693 , n61017 );
and ( n61019 , n60690 , n61018 );
or ( n61020 , n60689 , n61019 );
and ( n61021 , n60686 , n61020 );
or ( n61022 , n60685 , n61021 );
and ( n61023 , n60682 , n61022 );
or ( n61024 , n60681 , n61023 );
and ( n61025 , n60678 , n61024 );
or ( n61026 , n60677 , n61025 );
and ( n61027 , n60674 , n61026 );
or ( n61028 , n60673 , n61027 );
and ( n61029 , n60670 , n61028 );
or ( n61030 , n60669 , n61029 );
and ( n61031 , n60666 , n61030 );
or ( n61032 , n60665 , n61031 );
and ( n61033 , n60662 , n61032 );
or ( n61034 , n60661 , n61033 );
and ( n61035 , n60658 , n61034 );
or ( n61036 , n60657 , n61035 );
and ( n61037 , n60654 , n61036 );
or ( n61038 , n60653 , n61037 );
and ( n61039 , n60650 , n61038 );
or ( n61040 , n60649 , n61039 );
and ( n61041 , n60646 , n61040 );
or ( n61042 , n60645 , n61041 );
and ( n61043 , n60642 , n61042 );
or ( n61044 , n60641 , n61043 );
and ( n61045 , n60638 , n61044 );
or ( n61046 , n60637 , n61045 );
and ( n61047 , n60634 , n61046 );
or ( n61048 , n60633 , n61047 );
and ( n61049 , n60630 , n61048 );
or ( n61050 , n60629 , n61049 );
and ( n61051 , n60626 , n61050 );
or ( n61052 , n60625 , n61051 );
and ( n61053 , n60622 , n61052 );
or ( n61054 , n60621 , n61053 );
and ( n61055 , n60618 , n61054 );
or ( n61056 , n60617 , n61055 );
xor ( n61057 , n60614 , n61056 );
buf ( n61058 , n18000 );
and ( n61059 , n30044 , n61058 );
xor ( n61060 , n61057 , n61059 );
xor ( n61061 , n60618 , n61054 );
and ( n61062 , n30049 , n61058 );
and ( n61063 , n61061 , n61062 );
xor ( n61064 , n61061 , n61062 );
xor ( n61065 , n60622 , n61052 );
and ( n61066 , n30054 , n61058 );
and ( n61067 , n61065 , n61066 );
xor ( n61068 , n61065 , n61066 );
xor ( n61069 , n60626 , n61050 );
and ( n61070 , n30059 , n61058 );
and ( n61071 , n61069 , n61070 );
xor ( n61072 , n61069 , n61070 );
xor ( n61073 , n60630 , n61048 );
and ( n61074 , n30064 , n61058 );
and ( n61075 , n61073 , n61074 );
xor ( n61076 , n61073 , n61074 );
xor ( n61077 , n60634 , n61046 );
and ( n61078 , n30069 , n61058 );
and ( n61079 , n61077 , n61078 );
xor ( n61080 , n61077 , n61078 );
xor ( n61081 , n60638 , n61044 );
and ( n61082 , n30074 , n61058 );
and ( n61083 , n61081 , n61082 );
xor ( n61084 , n61081 , n61082 );
xor ( n61085 , n60642 , n61042 );
and ( n61086 , n30079 , n61058 );
and ( n61087 , n61085 , n61086 );
xor ( n61088 , n61085 , n61086 );
xor ( n61089 , n60646 , n61040 );
and ( n61090 , n30084 , n61058 );
and ( n61091 , n61089 , n61090 );
xor ( n61092 , n61089 , n61090 );
xor ( n61093 , n60650 , n61038 );
and ( n61094 , n30089 , n61058 );
and ( n61095 , n61093 , n61094 );
xor ( n61096 , n61093 , n61094 );
xor ( n61097 , n60654 , n61036 );
and ( n61098 , n30094 , n61058 );
and ( n61099 , n61097 , n61098 );
xor ( n61100 , n61097 , n61098 );
xor ( n61101 , n60658 , n61034 );
and ( n61102 , n30099 , n61058 );
and ( n61103 , n61101 , n61102 );
xor ( n61104 , n61101 , n61102 );
xor ( n61105 , n60662 , n61032 );
and ( n61106 , n30104 , n61058 );
and ( n61107 , n61105 , n61106 );
xor ( n61108 , n61105 , n61106 );
xor ( n61109 , n60666 , n61030 );
and ( n61110 , n30109 , n61058 );
and ( n61111 , n61109 , n61110 );
xor ( n61112 , n61109 , n61110 );
xor ( n61113 , n60670 , n61028 );
and ( n61114 , n30114 , n61058 );
and ( n61115 , n61113 , n61114 );
xor ( n61116 , n61113 , n61114 );
xor ( n61117 , n60674 , n61026 );
and ( n61118 , n30119 , n61058 );
and ( n61119 , n61117 , n61118 );
xor ( n61120 , n61117 , n61118 );
xor ( n61121 , n60678 , n61024 );
and ( n61122 , n30124 , n61058 );
and ( n61123 , n61121 , n61122 );
xor ( n61124 , n61121 , n61122 );
xor ( n61125 , n60682 , n61022 );
and ( n61126 , n30129 , n61058 );
and ( n61127 , n61125 , n61126 );
xor ( n61128 , n61125 , n61126 );
xor ( n61129 , n60686 , n61020 );
and ( n61130 , n30134 , n61058 );
and ( n61131 , n61129 , n61130 );
xor ( n61132 , n61129 , n61130 );
xor ( n61133 , n60690 , n61018 );
and ( n61134 , n30139 , n61058 );
and ( n61135 , n61133 , n61134 );
xor ( n61136 , n61133 , n61134 );
xor ( n61137 , n60694 , n61016 );
and ( n61138 , n30144 , n61058 );
and ( n61139 , n61137 , n61138 );
xor ( n61140 , n61137 , n61138 );
xor ( n61141 , n60698 , n61014 );
and ( n61142 , n30149 , n61058 );
and ( n61143 , n61141 , n61142 );
xor ( n61144 , n61141 , n61142 );
xor ( n61145 , n60702 , n61012 );
and ( n61146 , n30154 , n61058 );
and ( n61147 , n61145 , n61146 );
xor ( n61148 , n61145 , n61146 );
xor ( n61149 , n60706 , n61010 );
and ( n61150 , n30159 , n61058 );
and ( n61151 , n61149 , n61150 );
xor ( n61152 , n61149 , n61150 );
xor ( n61153 , n60710 , n61008 );
and ( n61154 , n30164 , n61058 );
and ( n61155 , n61153 , n61154 );
xor ( n61156 , n61153 , n61154 );
xor ( n61157 , n60714 , n61006 );
and ( n61158 , n30169 , n61058 );
and ( n61159 , n61157 , n61158 );
xor ( n61160 , n61157 , n61158 );
xor ( n61161 , n60718 , n61004 );
and ( n61162 , n30174 , n61058 );
and ( n61163 , n61161 , n61162 );
xor ( n61164 , n61161 , n61162 );
xor ( n61165 , n60722 , n61002 );
and ( n61166 , n30179 , n61058 );
and ( n61167 , n61165 , n61166 );
xor ( n61168 , n61165 , n61166 );
xor ( n61169 , n60726 , n61000 );
and ( n61170 , n30184 , n61058 );
and ( n61171 , n61169 , n61170 );
xor ( n61172 , n61169 , n61170 );
xor ( n61173 , n60730 , n60998 );
and ( n61174 , n30189 , n61058 );
and ( n61175 , n61173 , n61174 );
xor ( n61176 , n61173 , n61174 );
xor ( n61177 , n60734 , n60996 );
and ( n61178 , n30194 , n61058 );
and ( n61179 , n61177 , n61178 );
xor ( n61180 , n61177 , n61178 );
xor ( n61181 , n60738 , n60994 );
and ( n61182 , n30199 , n61058 );
and ( n61183 , n61181 , n61182 );
xor ( n61184 , n61181 , n61182 );
xor ( n61185 , n60742 , n60992 );
and ( n61186 , n30204 , n61058 );
and ( n61187 , n61185 , n61186 );
xor ( n61188 , n61185 , n61186 );
xor ( n61189 , n60746 , n60990 );
and ( n61190 , n30209 , n61058 );
and ( n61191 , n61189 , n61190 );
xor ( n61192 , n61189 , n61190 );
xor ( n61193 , n60750 , n60988 );
and ( n61194 , n30214 , n61058 );
and ( n61195 , n61193 , n61194 );
xor ( n61196 , n61193 , n61194 );
xor ( n61197 , n60754 , n60986 );
and ( n61198 , n30219 , n61058 );
and ( n61199 , n61197 , n61198 );
xor ( n61200 , n61197 , n61198 );
xor ( n61201 , n60758 , n60984 );
and ( n61202 , n30224 , n61058 );
and ( n61203 , n61201 , n61202 );
xor ( n61204 , n61201 , n61202 );
xor ( n61205 , n60762 , n60982 );
and ( n61206 , n30229 , n61058 );
and ( n61207 , n61205 , n61206 );
xor ( n61208 , n61205 , n61206 );
xor ( n61209 , n60766 , n60980 );
and ( n61210 , n30234 , n61058 );
and ( n61211 , n61209 , n61210 );
xor ( n61212 , n61209 , n61210 );
xor ( n61213 , n60770 , n60978 );
and ( n61214 , n30239 , n61058 );
and ( n61215 , n61213 , n61214 );
xor ( n61216 , n61213 , n61214 );
xor ( n61217 , n60774 , n60976 );
and ( n61218 , n30244 , n61058 );
and ( n61219 , n61217 , n61218 );
xor ( n61220 , n61217 , n61218 );
xor ( n61221 , n60778 , n60974 );
and ( n61222 , n30249 , n61058 );
and ( n61223 , n61221 , n61222 );
xor ( n61224 , n61221 , n61222 );
xor ( n61225 , n60782 , n60972 );
and ( n61226 , n30254 , n61058 );
and ( n61227 , n61225 , n61226 );
xor ( n61228 , n61225 , n61226 );
xor ( n61229 , n60786 , n60970 );
and ( n61230 , n30259 , n61058 );
and ( n61231 , n61229 , n61230 );
xor ( n61232 , n61229 , n61230 );
xor ( n61233 , n60790 , n60968 );
and ( n61234 , n30264 , n61058 );
and ( n61235 , n61233 , n61234 );
xor ( n61236 , n61233 , n61234 );
xor ( n61237 , n60794 , n60966 );
and ( n61238 , n30269 , n61058 );
and ( n61239 , n61237 , n61238 );
xor ( n61240 , n61237 , n61238 );
xor ( n61241 , n60798 , n60964 );
and ( n61242 , n30274 , n61058 );
and ( n61243 , n61241 , n61242 );
xor ( n61244 , n61241 , n61242 );
xor ( n61245 , n60802 , n60962 );
and ( n61246 , n30279 , n61058 );
and ( n61247 , n61245 , n61246 );
xor ( n61248 , n61245 , n61246 );
xor ( n61249 , n60806 , n60960 );
and ( n61250 , n30284 , n61058 );
and ( n61251 , n61249 , n61250 );
xor ( n61252 , n61249 , n61250 );
xor ( n61253 , n60810 , n60958 );
and ( n61254 , n30289 , n61058 );
and ( n61255 , n61253 , n61254 );
xor ( n61256 , n61253 , n61254 );
xor ( n61257 , n60814 , n60956 );
and ( n61258 , n30294 , n61058 );
and ( n61259 , n61257 , n61258 );
xor ( n61260 , n61257 , n61258 );
xor ( n61261 , n60818 , n60954 );
and ( n61262 , n30299 , n61058 );
and ( n61263 , n61261 , n61262 );
xor ( n61264 , n61261 , n61262 );
xor ( n61265 , n60822 , n60952 );
and ( n61266 , n30304 , n61058 );
and ( n61267 , n61265 , n61266 );
xor ( n61268 , n61265 , n61266 );
xor ( n61269 , n60826 , n60950 );
and ( n61270 , n30309 , n61058 );
and ( n61271 , n61269 , n61270 );
xor ( n61272 , n61269 , n61270 );
xor ( n61273 , n60830 , n60948 );
and ( n61274 , n30314 , n61058 );
and ( n61275 , n61273 , n61274 );
xor ( n61276 , n61273 , n61274 );
xor ( n61277 , n60834 , n60946 );
and ( n61278 , n30319 , n61058 );
and ( n61279 , n61277 , n61278 );
xor ( n61280 , n61277 , n61278 );
xor ( n61281 , n60838 , n60944 );
and ( n61282 , n30324 , n61058 );
and ( n61283 , n61281 , n61282 );
xor ( n61284 , n61281 , n61282 );
xor ( n61285 , n60842 , n60942 );
and ( n61286 , n30329 , n61058 );
and ( n61287 , n61285 , n61286 );
xor ( n61288 , n61285 , n61286 );
xor ( n61289 , n60846 , n60940 );
and ( n61290 , n30334 , n61058 );
and ( n61291 , n61289 , n61290 );
xor ( n61292 , n61289 , n61290 );
xor ( n61293 , n60850 , n60938 );
and ( n61294 , n30339 , n61058 );
and ( n61295 , n61293 , n61294 );
xor ( n61296 , n61293 , n61294 );
xor ( n61297 , n60854 , n60936 );
and ( n61298 , n30344 , n61058 );
and ( n61299 , n61297 , n61298 );
xor ( n61300 , n61297 , n61298 );
xor ( n61301 , n60858 , n60934 );
and ( n61302 , n30349 , n61058 );
and ( n61303 , n61301 , n61302 );
xor ( n61304 , n61301 , n61302 );
xor ( n61305 , n60862 , n60932 );
and ( n61306 , n30354 , n61058 );
and ( n61307 , n61305 , n61306 );
xor ( n61308 , n61305 , n61306 );
xor ( n61309 , n60866 , n60930 );
and ( n61310 , n30359 , n61058 );
and ( n61311 , n61309 , n61310 );
xor ( n61312 , n61309 , n61310 );
xor ( n61313 , n60870 , n60928 );
and ( n61314 , n30364 , n61058 );
and ( n61315 , n61313 , n61314 );
xor ( n61316 , n61313 , n61314 );
xor ( n61317 , n60874 , n60926 );
and ( n61318 , n30369 , n61058 );
and ( n61319 , n61317 , n61318 );
xor ( n61320 , n61317 , n61318 );
xor ( n61321 , n60878 , n60924 );
and ( n61322 , n30374 , n61058 );
and ( n61323 , n61321 , n61322 );
xor ( n61324 , n61321 , n61322 );
xor ( n61325 , n60882 , n60922 );
and ( n61326 , n30379 , n61058 );
and ( n61327 , n61325 , n61326 );
xor ( n61328 , n61325 , n61326 );
xor ( n61329 , n60886 , n60920 );
and ( n61330 , n30384 , n61058 );
and ( n61331 , n61329 , n61330 );
xor ( n61332 , n61329 , n61330 );
xor ( n61333 , n60890 , n60918 );
and ( n61334 , n30389 , n61058 );
and ( n61335 , n61333 , n61334 );
xor ( n61336 , n61333 , n61334 );
xor ( n61337 , n60894 , n60916 );
and ( n61338 , n30394 , n61058 );
and ( n61339 , n61337 , n61338 );
xor ( n61340 , n61337 , n61338 );
xor ( n61341 , n60898 , n60914 );
and ( n61342 , n30399 , n61058 );
and ( n61343 , n61341 , n61342 );
xor ( n61344 , n61341 , n61342 );
xor ( n61345 , n60902 , n60912 );
and ( n61346 , n30404 , n61058 );
and ( n61347 , n61345 , n61346 );
xor ( n61348 , n61345 , n61346 );
xor ( n61349 , n60906 , n60910 );
and ( n61350 , n30409 , n61058 );
and ( n61351 , n61349 , n61350 );
buf ( n61352 , n61351 );
and ( n61353 , n61348 , n61352 );
or ( n61354 , n61347 , n61353 );
and ( n61355 , n61344 , n61354 );
or ( n61356 , n61343 , n61355 );
and ( n61357 , n61340 , n61356 );
or ( n61358 , n61339 , n61357 );
and ( n61359 , n61336 , n61358 );
or ( n61360 , n61335 , n61359 );
and ( n61361 , n61332 , n61360 );
or ( n61362 , n61331 , n61361 );
and ( n61363 , n61328 , n61362 );
or ( n61364 , n61327 , n61363 );
and ( n61365 , n61324 , n61364 );
or ( n61366 , n61323 , n61365 );
and ( n61367 , n61320 , n61366 );
or ( n61368 , n61319 , n61367 );
and ( n61369 , n61316 , n61368 );
or ( n61370 , n61315 , n61369 );
and ( n61371 , n61312 , n61370 );
or ( n61372 , n61311 , n61371 );
and ( n61373 , n61308 , n61372 );
or ( n61374 , n61307 , n61373 );
and ( n61375 , n61304 , n61374 );
or ( n61376 , n61303 , n61375 );
and ( n61377 , n61300 , n61376 );
or ( n61378 , n61299 , n61377 );
and ( n61379 , n61296 , n61378 );
or ( n61380 , n61295 , n61379 );
and ( n61381 , n61292 , n61380 );
or ( n61382 , n61291 , n61381 );
and ( n61383 , n61288 , n61382 );
or ( n61384 , n61287 , n61383 );
and ( n61385 , n61284 , n61384 );
or ( n61386 , n61283 , n61385 );
and ( n61387 , n61280 , n61386 );
or ( n61388 , n61279 , n61387 );
and ( n61389 , n61276 , n61388 );
or ( n61390 , n61275 , n61389 );
and ( n61391 , n61272 , n61390 );
or ( n61392 , n61271 , n61391 );
and ( n61393 , n61268 , n61392 );
or ( n61394 , n61267 , n61393 );
and ( n61395 , n61264 , n61394 );
or ( n61396 , n61263 , n61395 );
and ( n61397 , n61260 , n61396 );
or ( n61398 , n61259 , n61397 );
and ( n61399 , n61256 , n61398 );
or ( n61400 , n61255 , n61399 );
and ( n61401 , n61252 , n61400 );
or ( n61402 , n61251 , n61401 );
and ( n61403 , n61248 , n61402 );
or ( n61404 , n61247 , n61403 );
and ( n61405 , n61244 , n61404 );
or ( n61406 , n61243 , n61405 );
and ( n61407 , n61240 , n61406 );
or ( n61408 , n61239 , n61407 );
and ( n61409 , n61236 , n61408 );
or ( n61410 , n61235 , n61409 );
and ( n61411 , n61232 , n61410 );
or ( n61412 , n61231 , n61411 );
and ( n61413 , n61228 , n61412 );
or ( n61414 , n61227 , n61413 );
and ( n61415 , n61224 , n61414 );
or ( n61416 , n61223 , n61415 );
and ( n61417 , n61220 , n61416 );
or ( n61418 , n61219 , n61417 );
and ( n61419 , n61216 , n61418 );
or ( n61420 , n61215 , n61419 );
and ( n61421 , n61212 , n61420 );
or ( n61422 , n61211 , n61421 );
and ( n61423 , n61208 , n61422 );
or ( n61424 , n61207 , n61423 );
and ( n61425 , n61204 , n61424 );
or ( n61426 , n61203 , n61425 );
and ( n61427 , n61200 , n61426 );
or ( n61428 , n61199 , n61427 );
and ( n61429 , n61196 , n61428 );
or ( n61430 , n61195 , n61429 );
and ( n61431 , n61192 , n61430 );
or ( n61432 , n61191 , n61431 );
and ( n61433 , n61188 , n61432 );
or ( n61434 , n61187 , n61433 );
and ( n61435 , n61184 , n61434 );
or ( n61436 , n61183 , n61435 );
and ( n61437 , n61180 , n61436 );
or ( n61438 , n61179 , n61437 );
and ( n61439 , n61176 , n61438 );
or ( n61440 , n61175 , n61439 );
and ( n61441 , n61172 , n61440 );
or ( n61442 , n61171 , n61441 );
and ( n61443 , n61168 , n61442 );
or ( n61444 , n61167 , n61443 );
and ( n61445 , n61164 , n61444 );
or ( n61446 , n61163 , n61445 );
and ( n61447 , n61160 , n61446 );
or ( n61448 , n61159 , n61447 );
and ( n61449 , n61156 , n61448 );
or ( n61450 , n61155 , n61449 );
and ( n61451 , n61152 , n61450 );
or ( n61452 , n61151 , n61451 );
and ( n61453 , n61148 , n61452 );
or ( n61454 , n61147 , n61453 );
and ( n61455 , n61144 , n61454 );
or ( n61456 , n61143 , n61455 );
and ( n61457 , n61140 , n61456 );
or ( n61458 , n61139 , n61457 );
and ( n61459 , n61136 , n61458 );
or ( n61460 , n61135 , n61459 );
and ( n61461 , n61132 , n61460 );
or ( n61462 , n61131 , n61461 );
and ( n61463 , n61128 , n61462 );
or ( n61464 , n61127 , n61463 );
and ( n61465 , n61124 , n61464 );
or ( n61466 , n61123 , n61465 );
and ( n61467 , n61120 , n61466 );
or ( n61468 , n61119 , n61467 );
and ( n61469 , n61116 , n61468 );
or ( n61470 , n61115 , n61469 );
and ( n61471 , n61112 , n61470 );
or ( n61472 , n61111 , n61471 );
and ( n61473 , n61108 , n61472 );
or ( n61474 , n61107 , n61473 );
and ( n61475 , n61104 , n61474 );
or ( n61476 , n61103 , n61475 );
and ( n61477 , n61100 , n61476 );
or ( n61478 , n61099 , n61477 );
and ( n61479 , n61096 , n61478 );
or ( n61480 , n61095 , n61479 );
and ( n61481 , n61092 , n61480 );
or ( n61482 , n61091 , n61481 );
and ( n61483 , n61088 , n61482 );
or ( n61484 , n61087 , n61483 );
and ( n61485 , n61084 , n61484 );
or ( n61486 , n61083 , n61485 );
and ( n61487 , n61080 , n61486 );
or ( n61488 , n61079 , n61487 );
and ( n61489 , n61076 , n61488 );
or ( n61490 , n61075 , n61489 );
and ( n61491 , n61072 , n61490 );
or ( n61492 , n61071 , n61491 );
and ( n61493 , n61068 , n61492 );
or ( n61494 , n61067 , n61493 );
and ( n61495 , n61064 , n61494 );
or ( n61496 , n61063 , n61495 );
xor ( n61497 , n61060 , n61496 );
buf ( n61498 , n17998 );
and ( n61499 , n30049 , n61498 );
xor ( n61500 , n61497 , n61499 );
xor ( n61501 , n61064 , n61494 );
and ( n61502 , n30054 , n61498 );
and ( n61503 , n61501 , n61502 );
xor ( n61504 , n61501 , n61502 );
xor ( n61505 , n61068 , n61492 );
and ( n61506 , n30059 , n61498 );
and ( n61507 , n61505 , n61506 );
xor ( n61508 , n61505 , n61506 );
xor ( n61509 , n61072 , n61490 );
and ( n61510 , n30064 , n61498 );
and ( n61511 , n61509 , n61510 );
xor ( n61512 , n61509 , n61510 );
xor ( n61513 , n61076 , n61488 );
and ( n61514 , n30069 , n61498 );
and ( n61515 , n61513 , n61514 );
xor ( n61516 , n61513 , n61514 );
xor ( n61517 , n61080 , n61486 );
and ( n61518 , n30074 , n61498 );
and ( n61519 , n61517 , n61518 );
xor ( n61520 , n61517 , n61518 );
xor ( n61521 , n61084 , n61484 );
and ( n61522 , n30079 , n61498 );
and ( n61523 , n61521 , n61522 );
xor ( n61524 , n61521 , n61522 );
xor ( n61525 , n61088 , n61482 );
and ( n61526 , n30084 , n61498 );
and ( n61527 , n61525 , n61526 );
xor ( n61528 , n61525 , n61526 );
xor ( n61529 , n61092 , n61480 );
and ( n61530 , n30089 , n61498 );
and ( n61531 , n61529 , n61530 );
xor ( n61532 , n61529 , n61530 );
xor ( n61533 , n61096 , n61478 );
and ( n61534 , n30094 , n61498 );
and ( n61535 , n61533 , n61534 );
xor ( n61536 , n61533 , n61534 );
xor ( n61537 , n61100 , n61476 );
and ( n61538 , n30099 , n61498 );
and ( n61539 , n61537 , n61538 );
xor ( n61540 , n61537 , n61538 );
xor ( n61541 , n61104 , n61474 );
and ( n61542 , n30104 , n61498 );
and ( n61543 , n61541 , n61542 );
xor ( n61544 , n61541 , n61542 );
xor ( n61545 , n61108 , n61472 );
and ( n61546 , n30109 , n61498 );
and ( n61547 , n61545 , n61546 );
xor ( n61548 , n61545 , n61546 );
xor ( n61549 , n61112 , n61470 );
and ( n61550 , n30114 , n61498 );
and ( n61551 , n61549 , n61550 );
xor ( n61552 , n61549 , n61550 );
xor ( n61553 , n61116 , n61468 );
and ( n61554 , n30119 , n61498 );
and ( n61555 , n61553 , n61554 );
xor ( n61556 , n61553 , n61554 );
xor ( n61557 , n61120 , n61466 );
and ( n61558 , n30124 , n61498 );
and ( n61559 , n61557 , n61558 );
xor ( n61560 , n61557 , n61558 );
xor ( n61561 , n61124 , n61464 );
and ( n61562 , n30129 , n61498 );
and ( n61563 , n61561 , n61562 );
xor ( n61564 , n61561 , n61562 );
xor ( n61565 , n61128 , n61462 );
and ( n61566 , n30134 , n61498 );
and ( n61567 , n61565 , n61566 );
xor ( n61568 , n61565 , n61566 );
xor ( n61569 , n61132 , n61460 );
and ( n61570 , n30139 , n61498 );
and ( n61571 , n61569 , n61570 );
xor ( n61572 , n61569 , n61570 );
xor ( n61573 , n61136 , n61458 );
and ( n61574 , n30144 , n61498 );
and ( n61575 , n61573 , n61574 );
xor ( n61576 , n61573 , n61574 );
xor ( n61577 , n61140 , n61456 );
and ( n61578 , n30149 , n61498 );
and ( n61579 , n61577 , n61578 );
xor ( n61580 , n61577 , n61578 );
xor ( n61581 , n61144 , n61454 );
and ( n61582 , n30154 , n61498 );
and ( n61583 , n61581 , n61582 );
xor ( n61584 , n61581 , n61582 );
xor ( n61585 , n61148 , n61452 );
and ( n61586 , n30159 , n61498 );
and ( n61587 , n61585 , n61586 );
xor ( n61588 , n61585 , n61586 );
xor ( n61589 , n61152 , n61450 );
and ( n61590 , n30164 , n61498 );
and ( n61591 , n61589 , n61590 );
xor ( n61592 , n61589 , n61590 );
xor ( n61593 , n61156 , n61448 );
and ( n61594 , n30169 , n61498 );
and ( n61595 , n61593 , n61594 );
xor ( n61596 , n61593 , n61594 );
xor ( n61597 , n61160 , n61446 );
and ( n61598 , n30174 , n61498 );
and ( n61599 , n61597 , n61598 );
xor ( n61600 , n61597 , n61598 );
xor ( n61601 , n61164 , n61444 );
and ( n61602 , n30179 , n61498 );
and ( n61603 , n61601 , n61602 );
xor ( n61604 , n61601 , n61602 );
xor ( n61605 , n61168 , n61442 );
and ( n61606 , n30184 , n61498 );
and ( n61607 , n61605 , n61606 );
xor ( n61608 , n61605 , n61606 );
xor ( n61609 , n61172 , n61440 );
and ( n61610 , n30189 , n61498 );
and ( n61611 , n61609 , n61610 );
xor ( n61612 , n61609 , n61610 );
xor ( n61613 , n61176 , n61438 );
and ( n61614 , n30194 , n61498 );
and ( n61615 , n61613 , n61614 );
xor ( n61616 , n61613 , n61614 );
xor ( n61617 , n61180 , n61436 );
and ( n61618 , n30199 , n61498 );
and ( n61619 , n61617 , n61618 );
xor ( n61620 , n61617 , n61618 );
xor ( n61621 , n61184 , n61434 );
and ( n61622 , n30204 , n61498 );
and ( n61623 , n61621 , n61622 );
xor ( n61624 , n61621 , n61622 );
xor ( n61625 , n61188 , n61432 );
and ( n61626 , n30209 , n61498 );
and ( n61627 , n61625 , n61626 );
xor ( n61628 , n61625 , n61626 );
xor ( n61629 , n61192 , n61430 );
and ( n61630 , n30214 , n61498 );
and ( n61631 , n61629 , n61630 );
xor ( n61632 , n61629 , n61630 );
xor ( n61633 , n61196 , n61428 );
and ( n61634 , n30219 , n61498 );
and ( n61635 , n61633 , n61634 );
xor ( n61636 , n61633 , n61634 );
xor ( n61637 , n61200 , n61426 );
and ( n61638 , n30224 , n61498 );
and ( n61639 , n61637 , n61638 );
xor ( n61640 , n61637 , n61638 );
xor ( n61641 , n61204 , n61424 );
and ( n61642 , n30229 , n61498 );
and ( n61643 , n61641 , n61642 );
xor ( n61644 , n61641 , n61642 );
xor ( n61645 , n61208 , n61422 );
and ( n61646 , n30234 , n61498 );
and ( n61647 , n61645 , n61646 );
xor ( n61648 , n61645 , n61646 );
xor ( n61649 , n61212 , n61420 );
and ( n61650 , n30239 , n61498 );
and ( n61651 , n61649 , n61650 );
xor ( n61652 , n61649 , n61650 );
xor ( n61653 , n61216 , n61418 );
and ( n61654 , n30244 , n61498 );
and ( n61655 , n61653 , n61654 );
xor ( n61656 , n61653 , n61654 );
xor ( n61657 , n61220 , n61416 );
and ( n61658 , n30249 , n61498 );
and ( n61659 , n61657 , n61658 );
xor ( n61660 , n61657 , n61658 );
xor ( n61661 , n61224 , n61414 );
and ( n61662 , n30254 , n61498 );
and ( n61663 , n61661 , n61662 );
xor ( n61664 , n61661 , n61662 );
xor ( n61665 , n61228 , n61412 );
and ( n61666 , n30259 , n61498 );
and ( n61667 , n61665 , n61666 );
xor ( n61668 , n61665 , n61666 );
xor ( n61669 , n61232 , n61410 );
and ( n61670 , n30264 , n61498 );
and ( n61671 , n61669 , n61670 );
xor ( n61672 , n61669 , n61670 );
xor ( n61673 , n61236 , n61408 );
and ( n61674 , n30269 , n61498 );
and ( n61675 , n61673 , n61674 );
xor ( n61676 , n61673 , n61674 );
xor ( n61677 , n61240 , n61406 );
and ( n61678 , n30274 , n61498 );
and ( n61679 , n61677 , n61678 );
xor ( n61680 , n61677 , n61678 );
xor ( n61681 , n61244 , n61404 );
and ( n61682 , n30279 , n61498 );
and ( n61683 , n61681 , n61682 );
xor ( n61684 , n61681 , n61682 );
xor ( n61685 , n61248 , n61402 );
and ( n61686 , n30284 , n61498 );
and ( n61687 , n61685 , n61686 );
xor ( n61688 , n61685 , n61686 );
xor ( n61689 , n61252 , n61400 );
and ( n61690 , n30289 , n61498 );
and ( n61691 , n61689 , n61690 );
xor ( n61692 , n61689 , n61690 );
xor ( n61693 , n61256 , n61398 );
and ( n61694 , n30294 , n61498 );
and ( n61695 , n61693 , n61694 );
xor ( n61696 , n61693 , n61694 );
xor ( n61697 , n61260 , n61396 );
and ( n61698 , n30299 , n61498 );
and ( n61699 , n61697 , n61698 );
xor ( n61700 , n61697 , n61698 );
xor ( n61701 , n61264 , n61394 );
and ( n61702 , n30304 , n61498 );
and ( n61703 , n61701 , n61702 );
xor ( n61704 , n61701 , n61702 );
xor ( n61705 , n61268 , n61392 );
and ( n61706 , n30309 , n61498 );
and ( n61707 , n61705 , n61706 );
xor ( n61708 , n61705 , n61706 );
xor ( n61709 , n61272 , n61390 );
and ( n61710 , n30314 , n61498 );
and ( n61711 , n61709 , n61710 );
xor ( n61712 , n61709 , n61710 );
xor ( n61713 , n61276 , n61388 );
and ( n61714 , n30319 , n61498 );
and ( n61715 , n61713 , n61714 );
xor ( n61716 , n61713 , n61714 );
xor ( n61717 , n61280 , n61386 );
and ( n61718 , n30324 , n61498 );
and ( n61719 , n61717 , n61718 );
xor ( n61720 , n61717 , n61718 );
xor ( n61721 , n61284 , n61384 );
and ( n61722 , n30329 , n61498 );
and ( n61723 , n61721 , n61722 );
xor ( n61724 , n61721 , n61722 );
xor ( n61725 , n61288 , n61382 );
and ( n61726 , n30334 , n61498 );
and ( n61727 , n61725 , n61726 );
xor ( n61728 , n61725 , n61726 );
xor ( n61729 , n61292 , n61380 );
and ( n61730 , n30339 , n61498 );
and ( n61731 , n61729 , n61730 );
xor ( n61732 , n61729 , n61730 );
xor ( n61733 , n61296 , n61378 );
and ( n61734 , n30344 , n61498 );
and ( n61735 , n61733 , n61734 );
xor ( n61736 , n61733 , n61734 );
xor ( n61737 , n61300 , n61376 );
and ( n61738 , n30349 , n61498 );
and ( n61739 , n61737 , n61738 );
xor ( n61740 , n61737 , n61738 );
xor ( n61741 , n61304 , n61374 );
and ( n61742 , n30354 , n61498 );
and ( n61743 , n61741 , n61742 );
xor ( n61744 , n61741 , n61742 );
xor ( n61745 , n61308 , n61372 );
and ( n61746 , n30359 , n61498 );
and ( n61747 , n61745 , n61746 );
xor ( n61748 , n61745 , n61746 );
xor ( n61749 , n61312 , n61370 );
and ( n61750 , n30364 , n61498 );
and ( n61751 , n61749 , n61750 );
xor ( n61752 , n61749 , n61750 );
xor ( n61753 , n61316 , n61368 );
and ( n61754 , n30369 , n61498 );
and ( n61755 , n61753 , n61754 );
xor ( n61756 , n61753 , n61754 );
xor ( n61757 , n61320 , n61366 );
and ( n61758 , n30374 , n61498 );
and ( n61759 , n61757 , n61758 );
xor ( n61760 , n61757 , n61758 );
xor ( n61761 , n61324 , n61364 );
and ( n61762 , n30379 , n61498 );
and ( n61763 , n61761 , n61762 );
xor ( n61764 , n61761 , n61762 );
xor ( n61765 , n61328 , n61362 );
and ( n61766 , n30384 , n61498 );
and ( n61767 , n61765 , n61766 );
xor ( n61768 , n61765 , n61766 );
xor ( n61769 , n61332 , n61360 );
and ( n61770 , n30389 , n61498 );
and ( n61771 , n61769 , n61770 );
xor ( n61772 , n61769 , n61770 );
xor ( n61773 , n61336 , n61358 );
and ( n61774 , n30394 , n61498 );
and ( n61775 , n61773 , n61774 );
xor ( n61776 , n61773 , n61774 );
xor ( n61777 , n61340 , n61356 );
and ( n61778 , n30399 , n61498 );
and ( n61779 , n61777 , n61778 );
xor ( n61780 , n61777 , n61778 );
xor ( n61781 , n61344 , n61354 );
and ( n61782 , n30404 , n61498 );
and ( n61783 , n61781 , n61782 );
xor ( n61784 , n61781 , n61782 );
xor ( n61785 , n61348 , n61352 );
and ( n61786 , n30409 , n61498 );
and ( n61787 , n61785 , n61786 );
buf ( n61788 , n61787 );
and ( n61789 , n61784 , n61788 );
or ( n61790 , n61783 , n61789 );
and ( n61791 , n61780 , n61790 );
or ( n61792 , n61779 , n61791 );
and ( n61793 , n61776 , n61792 );
or ( n61794 , n61775 , n61793 );
and ( n61795 , n61772 , n61794 );
or ( n61796 , n61771 , n61795 );
and ( n61797 , n61768 , n61796 );
or ( n61798 , n61767 , n61797 );
and ( n61799 , n61764 , n61798 );
or ( n61800 , n61763 , n61799 );
and ( n61801 , n61760 , n61800 );
or ( n61802 , n61759 , n61801 );
and ( n61803 , n61756 , n61802 );
or ( n61804 , n61755 , n61803 );
and ( n61805 , n61752 , n61804 );
or ( n61806 , n61751 , n61805 );
and ( n61807 , n61748 , n61806 );
or ( n61808 , n61747 , n61807 );
and ( n61809 , n61744 , n61808 );
or ( n61810 , n61743 , n61809 );
and ( n61811 , n61740 , n61810 );
or ( n61812 , n61739 , n61811 );
and ( n61813 , n61736 , n61812 );
or ( n61814 , n61735 , n61813 );
and ( n61815 , n61732 , n61814 );
or ( n61816 , n61731 , n61815 );
and ( n61817 , n61728 , n61816 );
or ( n61818 , n61727 , n61817 );
and ( n61819 , n61724 , n61818 );
or ( n61820 , n61723 , n61819 );
and ( n61821 , n61720 , n61820 );
or ( n61822 , n61719 , n61821 );
and ( n61823 , n61716 , n61822 );
or ( n61824 , n61715 , n61823 );
and ( n61825 , n61712 , n61824 );
or ( n61826 , n61711 , n61825 );
and ( n61827 , n61708 , n61826 );
or ( n61828 , n61707 , n61827 );
and ( n61829 , n61704 , n61828 );
or ( n61830 , n61703 , n61829 );
and ( n61831 , n61700 , n61830 );
or ( n61832 , n61699 , n61831 );
and ( n61833 , n61696 , n61832 );
or ( n61834 , n61695 , n61833 );
and ( n61835 , n61692 , n61834 );
or ( n61836 , n61691 , n61835 );
and ( n61837 , n61688 , n61836 );
or ( n61838 , n61687 , n61837 );
and ( n61839 , n61684 , n61838 );
or ( n61840 , n61683 , n61839 );
and ( n61841 , n61680 , n61840 );
or ( n61842 , n61679 , n61841 );
and ( n61843 , n61676 , n61842 );
or ( n61844 , n61675 , n61843 );
and ( n61845 , n61672 , n61844 );
or ( n61846 , n61671 , n61845 );
and ( n61847 , n61668 , n61846 );
or ( n61848 , n61667 , n61847 );
and ( n61849 , n61664 , n61848 );
or ( n61850 , n61663 , n61849 );
and ( n61851 , n61660 , n61850 );
or ( n61852 , n61659 , n61851 );
and ( n61853 , n61656 , n61852 );
or ( n61854 , n61655 , n61853 );
and ( n61855 , n61652 , n61854 );
or ( n61856 , n61651 , n61855 );
and ( n61857 , n61648 , n61856 );
or ( n61858 , n61647 , n61857 );
and ( n61859 , n61644 , n61858 );
or ( n61860 , n61643 , n61859 );
and ( n61861 , n61640 , n61860 );
or ( n61862 , n61639 , n61861 );
and ( n61863 , n61636 , n61862 );
or ( n61864 , n61635 , n61863 );
and ( n61865 , n61632 , n61864 );
or ( n61866 , n61631 , n61865 );
and ( n61867 , n61628 , n61866 );
or ( n61868 , n61627 , n61867 );
and ( n61869 , n61624 , n61868 );
or ( n61870 , n61623 , n61869 );
and ( n61871 , n61620 , n61870 );
or ( n61872 , n61619 , n61871 );
and ( n61873 , n61616 , n61872 );
or ( n61874 , n61615 , n61873 );
and ( n61875 , n61612 , n61874 );
or ( n61876 , n61611 , n61875 );
and ( n61877 , n61608 , n61876 );
or ( n61878 , n61607 , n61877 );
and ( n61879 , n61604 , n61878 );
or ( n61880 , n61603 , n61879 );
and ( n61881 , n61600 , n61880 );
or ( n61882 , n61599 , n61881 );
and ( n61883 , n61596 , n61882 );
or ( n61884 , n61595 , n61883 );
and ( n61885 , n61592 , n61884 );
or ( n61886 , n61591 , n61885 );
and ( n61887 , n61588 , n61886 );
or ( n61888 , n61587 , n61887 );
and ( n61889 , n61584 , n61888 );
or ( n61890 , n61583 , n61889 );
and ( n61891 , n61580 , n61890 );
or ( n61892 , n61579 , n61891 );
and ( n61893 , n61576 , n61892 );
or ( n61894 , n61575 , n61893 );
and ( n61895 , n61572 , n61894 );
or ( n61896 , n61571 , n61895 );
and ( n61897 , n61568 , n61896 );
or ( n61898 , n61567 , n61897 );
and ( n61899 , n61564 , n61898 );
or ( n61900 , n61563 , n61899 );
and ( n61901 , n61560 , n61900 );
or ( n61902 , n61559 , n61901 );
and ( n61903 , n61556 , n61902 );
or ( n61904 , n61555 , n61903 );
and ( n61905 , n61552 , n61904 );
or ( n61906 , n61551 , n61905 );
and ( n61907 , n61548 , n61906 );
or ( n61908 , n61547 , n61907 );
and ( n61909 , n61544 , n61908 );
or ( n61910 , n61543 , n61909 );
and ( n61911 , n61540 , n61910 );
or ( n61912 , n61539 , n61911 );
and ( n61913 , n61536 , n61912 );
or ( n61914 , n61535 , n61913 );
and ( n61915 , n61532 , n61914 );
or ( n61916 , n61531 , n61915 );
and ( n61917 , n61528 , n61916 );
or ( n61918 , n61527 , n61917 );
and ( n61919 , n61524 , n61918 );
or ( n61920 , n61523 , n61919 );
and ( n61921 , n61520 , n61920 );
or ( n61922 , n61519 , n61921 );
and ( n61923 , n61516 , n61922 );
or ( n61924 , n61515 , n61923 );
and ( n61925 , n61512 , n61924 );
or ( n61926 , n61511 , n61925 );
and ( n61927 , n61508 , n61926 );
or ( n61928 , n61507 , n61927 );
and ( n61929 , n61504 , n61928 );
or ( n61930 , n61503 , n61929 );
xor ( n61931 , n61500 , n61930 );
buf ( n61932 , n17996 );
and ( n61933 , n30054 , n61932 );
xor ( n61934 , n61931 , n61933 );
xor ( n61935 , n61504 , n61928 );
and ( n61936 , n30059 , n61932 );
and ( n61937 , n61935 , n61936 );
xor ( n61938 , n61935 , n61936 );
xor ( n61939 , n61508 , n61926 );
and ( n61940 , n30064 , n61932 );
and ( n61941 , n61939 , n61940 );
xor ( n61942 , n61939 , n61940 );
xor ( n61943 , n61512 , n61924 );
and ( n61944 , n30069 , n61932 );
and ( n61945 , n61943 , n61944 );
xor ( n61946 , n61943 , n61944 );
xor ( n61947 , n61516 , n61922 );
and ( n61948 , n30074 , n61932 );
and ( n61949 , n61947 , n61948 );
xor ( n61950 , n61947 , n61948 );
xor ( n61951 , n61520 , n61920 );
and ( n61952 , n30079 , n61932 );
and ( n61953 , n61951 , n61952 );
xor ( n61954 , n61951 , n61952 );
xor ( n61955 , n61524 , n61918 );
and ( n61956 , n30084 , n61932 );
and ( n61957 , n61955 , n61956 );
xor ( n61958 , n61955 , n61956 );
xor ( n61959 , n61528 , n61916 );
and ( n61960 , n30089 , n61932 );
and ( n61961 , n61959 , n61960 );
xor ( n61962 , n61959 , n61960 );
xor ( n61963 , n61532 , n61914 );
and ( n61964 , n30094 , n61932 );
and ( n61965 , n61963 , n61964 );
xor ( n61966 , n61963 , n61964 );
xor ( n61967 , n61536 , n61912 );
and ( n61968 , n30099 , n61932 );
and ( n61969 , n61967 , n61968 );
xor ( n61970 , n61967 , n61968 );
xor ( n61971 , n61540 , n61910 );
and ( n61972 , n30104 , n61932 );
and ( n61973 , n61971 , n61972 );
xor ( n61974 , n61971 , n61972 );
xor ( n61975 , n61544 , n61908 );
and ( n61976 , n30109 , n61932 );
and ( n61977 , n61975 , n61976 );
xor ( n61978 , n61975 , n61976 );
xor ( n61979 , n61548 , n61906 );
and ( n61980 , n30114 , n61932 );
and ( n61981 , n61979 , n61980 );
xor ( n61982 , n61979 , n61980 );
xor ( n61983 , n61552 , n61904 );
and ( n61984 , n30119 , n61932 );
and ( n61985 , n61983 , n61984 );
xor ( n61986 , n61983 , n61984 );
xor ( n61987 , n61556 , n61902 );
and ( n61988 , n30124 , n61932 );
and ( n61989 , n61987 , n61988 );
xor ( n61990 , n61987 , n61988 );
xor ( n61991 , n61560 , n61900 );
and ( n61992 , n30129 , n61932 );
and ( n61993 , n61991 , n61992 );
xor ( n61994 , n61991 , n61992 );
xor ( n61995 , n61564 , n61898 );
and ( n61996 , n30134 , n61932 );
and ( n61997 , n61995 , n61996 );
xor ( n61998 , n61995 , n61996 );
xor ( n61999 , n61568 , n61896 );
and ( n62000 , n30139 , n61932 );
and ( n62001 , n61999 , n62000 );
xor ( n62002 , n61999 , n62000 );
xor ( n62003 , n61572 , n61894 );
and ( n62004 , n30144 , n61932 );
and ( n62005 , n62003 , n62004 );
xor ( n62006 , n62003 , n62004 );
xor ( n62007 , n61576 , n61892 );
and ( n62008 , n30149 , n61932 );
and ( n62009 , n62007 , n62008 );
xor ( n62010 , n62007 , n62008 );
xor ( n62011 , n61580 , n61890 );
and ( n62012 , n30154 , n61932 );
and ( n62013 , n62011 , n62012 );
xor ( n62014 , n62011 , n62012 );
xor ( n62015 , n61584 , n61888 );
and ( n62016 , n30159 , n61932 );
and ( n62017 , n62015 , n62016 );
xor ( n62018 , n62015 , n62016 );
xor ( n62019 , n61588 , n61886 );
and ( n62020 , n30164 , n61932 );
and ( n62021 , n62019 , n62020 );
xor ( n62022 , n62019 , n62020 );
xor ( n62023 , n61592 , n61884 );
and ( n62024 , n30169 , n61932 );
and ( n62025 , n62023 , n62024 );
xor ( n62026 , n62023 , n62024 );
xor ( n62027 , n61596 , n61882 );
and ( n62028 , n30174 , n61932 );
and ( n62029 , n62027 , n62028 );
xor ( n62030 , n62027 , n62028 );
xor ( n62031 , n61600 , n61880 );
and ( n62032 , n30179 , n61932 );
and ( n62033 , n62031 , n62032 );
xor ( n62034 , n62031 , n62032 );
xor ( n62035 , n61604 , n61878 );
and ( n62036 , n30184 , n61932 );
and ( n62037 , n62035 , n62036 );
xor ( n62038 , n62035 , n62036 );
xor ( n62039 , n61608 , n61876 );
and ( n62040 , n30189 , n61932 );
and ( n62041 , n62039 , n62040 );
xor ( n62042 , n62039 , n62040 );
xor ( n62043 , n61612 , n61874 );
and ( n62044 , n30194 , n61932 );
and ( n62045 , n62043 , n62044 );
xor ( n62046 , n62043 , n62044 );
xor ( n62047 , n61616 , n61872 );
and ( n62048 , n30199 , n61932 );
and ( n62049 , n62047 , n62048 );
xor ( n62050 , n62047 , n62048 );
xor ( n62051 , n61620 , n61870 );
and ( n62052 , n30204 , n61932 );
and ( n62053 , n62051 , n62052 );
xor ( n62054 , n62051 , n62052 );
xor ( n62055 , n61624 , n61868 );
and ( n62056 , n30209 , n61932 );
and ( n62057 , n62055 , n62056 );
xor ( n62058 , n62055 , n62056 );
xor ( n62059 , n61628 , n61866 );
and ( n62060 , n30214 , n61932 );
and ( n62061 , n62059 , n62060 );
xor ( n62062 , n62059 , n62060 );
xor ( n62063 , n61632 , n61864 );
and ( n62064 , n30219 , n61932 );
and ( n62065 , n62063 , n62064 );
xor ( n62066 , n62063 , n62064 );
xor ( n62067 , n61636 , n61862 );
and ( n62068 , n30224 , n61932 );
and ( n62069 , n62067 , n62068 );
xor ( n62070 , n62067 , n62068 );
xor ( n62071 , n61640 , n61860 );
and ( n62072 , n30229 , n61932 );
and ( n62073 , n62071 , n62072 );
xor ( n62074 , n62071 , n62072 );
xor ( n62075 , n61644 , n61858 );
and ( n62076 , n30234 , n61932 );
and ( n62077 , n62075 , n62076 );
xor ( n62078 , n62075 , n62076 );
xor ( n62079 , n61648 , n61856 );
and ( n62080 , n30239 , n61932 );
and ( n62081 , n62079 , n62080 );
xor ( n62082 , n62079 , n62080 );
xor ( n62083 , n61652 , n61854 );
and ( n62084 , n30244 , n61932 );
and ( n62085 , n62083 , n62084 );
xor ( n62086 , n62083 , n62084 );
xor ( n62087 , n61656 , n61852 );
and ( n62088 , n30249 , n61932 );
and ( n62089 , n62087 , n62088 );
xor ( n62090 , n62087 , n62088 );
xor ( n62091 , n61660 , n61850 );
and ( n62092 , n30254 , n61932 );
and ( n62093 , n62091 , n62092 );
xor ( n62094 , n62091 , n62092 );
xor ( n62095 , n61664 , n61848 );
and ( n62096 , n30259 , n61932 );
and ( n62097 , n62095 , n62096 );
xor ( n62098 , n62095 , n62096 );
xor ( n62099 , n61668 , n61846 );
and ( n62100 , n30264 , n61932 );
and ( n62101 , n62099 , n62100 );
xor ( n62102 , n62099 , n62100 );
xor ( n62103 , n61672 , n61844 );
and ( n62104 , n30269 , n61932 );
and ( n62105 , n62103 , n62104 );
xor ( n62106 , n62103 , n62104 );
xor ( n62107 , n61676 , n61842 );
and ( n62108 , n30274 , n61932 );
and ( n62109 , n62107 , n62108 );
xor ( n62110 , n62107 , n62108 );
xor ( n62111 , n61680 , n61840 );
and ( n62112 , n30279 , n61932 );
and ( n62113 , n62111 , n62112 );
xor ( n62114 , n62111 , n62112 );
xor ( n62115 , n61684 , n61838 );
and ( n62116 , n30284 , n61932 );
and ( n62117 , n62115 , n62116 );
xor ( n62118 , n62115 , n62116 );
xor ( n62119 , n61688 , n61836 );
and ( n62120 , n30289 , n61932 );
and ( n62121 , n62119 , n62120 );
xor ( n62122 , n62119 , n62120 );
xor ( n62123 , n61692 , n61834 );
and ( n62124 , n30294 , n61932 );
and ( n62125 , n62123 , n62124 );
xor ( n62126 , n62123 , n62124 );
xor ( n62127 , n61696 , n61832 );
and ( n62128 , n30299 , n61932 );
and ( n62129 , n62127 , n62128 );
xor ( n62130 , n62127 , n62128 );
xor ( n62131 , n61700 , n61830 );
and ( n62132 , n30304 , n61932 );
and ( n62133 , n62131 , n62132 );
xor ( n62134 , n62131 , n62132 );
xor ( n62135 , n61704 , n61828 );
and ( n62136 , n30309 , n61932 );
and ( n62137 , n62135 , n62136 );
xor ( n62138 , n62135 , n62136 );
xor ( n62139 , n61708 , n61826 );
and ( n62140 , n30314 , n61932 );
and ( n62141 , n62139 , n62140 );
xor ( n62142 , n62139 , n62140 );
xor ( n62143 , n61712 , n61824 );
and ( n62144 , n30319 , n61932 );
and ( n62145 , n62143 , n62144 );
xor ( n62146 , n62143 , n62144 );
xor ( n62147 , n61716 , n61822 );
and ( n62148 , n30324 , n61932 );
and ( n62149 , n62147 , n62148 );
xor ( n62150 , n62147 , n62148 );
xor ( n62151 , n61720 , n61820 );
and ( n62152 , n30329 , n61932 );
and ( n62153 , n62151 , n62152 );
xor ( n62154 , n62151 , n62152 );
xor ( n62155 , n61724 , n61818 );
and ( n62156 , n30334 , n61932 );
and ( n62157 , n62155 , n62156 );
xor ( n62158 , n62155 , n62156 );
xor ( n62159 , n61728 , n61816 );
and ( n62160 , n30339 , n61932 );
and ( n62161 , n62159 , n62160 );
xor ( n62162 , n62159 , n62160 );
xor ( n62163 , n61732 , n61814 );
and ( n62164 , n30344 , n61932 );
and ( n62165 , n62163 , n62164 );
xor ( n62166 , n62163 , n62164 );
xor ( n62167 , n61736 , n61812 );
and ( n62168 , n30349 , n61932 );
and ( n62169 , n62167 , n62168 );
xor ( n62170 , n62167 , n62168 );
xor ( n62171 , n61740 , n61810 );
and ( n62172 , n30354 , n61932 );
and ( n62173 , n62171 , n62172 );
xor ( n62174 , n62171 , n62172 );
xor ( n62175 , n61744 , n61808 );
and ( n62176 , n30359 , n61932 );
and ( n62177 , n62175 , n62176 );
xor ( n62178 , n62175 , n62176 );
xor ( n62179 , n61748 , n61806 );
and ( n62180 , n30364 , n61932 );
and ( n62181 , n62179 , n62180 );
xor ( n62182 , n62179 , n62180 );
xor ( n62183 , n61752 , n61804 );
and ( n62184 , n30369 , n61932 );
and ( n62185 , n62183 , n62184 );
xor ( n62186 , n62183 , n62184 );
xor ( n62187 , n61756 , n61802 );
and ( n62188 , n30374 , n61932 );
and ( n62189 , n62187 , n62188 );
xor ( n62190 , n62187 , n62188 );
xor ( n62191 , n61760 , n61800 );
and ( n62192 , n30379 , n61932 );
and ( n62193 , n62191 , n62192 );
xor ( n62194 , n62191 , n62192 );
xor ( n62195 , n61764 , n61798 );
and ( n62196 , n30384 , n61932 );
and ( n62197 , n62195 , n62196 );
xor ( n62198 , n62195 , n62196 );
xor ( n62199 , n61768 , n61796 );
and ( n62200 , n30389 , n61932 );
and ( n62201 , n62199 , n62200 );
xor ( n62202 , n62199 , n62200 );
xor ( n62203 , n61772 , n61794 );
and ( n62204 , n30394 , n61932 );
and ( n62205 , n62203 , n62204 );
xor ( n62206 , n62203 , n62204 );
xor ( n62207 , n61776 , n61792 );
and ( n62208 , n30399 , n61932 );
and ( n62209 , n62207 , n62208 );
xor ( n62210 , n62207 , n62208 );
xor ( n62211 , n61780 , n61790 );
and ( n62212 , n30404 , n61932 );
and ( n62213 , n62211 , n62212 );
xor ( n62214 , n62211 , n62212 );
xor ( n62215 , n61784 , n61788 );
and ( n62216 , n30409 , n61932 );
and ( n62217 , n62215 , n62216 );
buf ( n62218 , n62217 );
and ( n62219 , n62214 , n62218 );
or ( n62220 , n62213 , n62219 );
and ( n62221 , n62210 , n62220 );
or ( n62222 , n62209 , n62221 );
and ( n62223 , n62206 , n62222 );
or ( n62224 , n62205 , n62223 );
and ( n62225 , n62202 , n62224 );
or ( n62226 , n62201 , n62225 );
and ( n62227 , n62198 , n62226 );
or ( n62228 , n62197 , n62227 );
and ( n62229 , n62194 , n62228 );
or ( n62230 , n62193 , n62229 );
and ( n62231 , n62190 , n62230 );
or ( n62232 , n62189 , n62231 );
and ( n62233 , n62186 , n62232 );
or ( n62234 , n62185 , n62233 );
and ( n62235 , n62182 , n62234 );
or ( n62236 , n62181 , n62235 );
and ( n62237 , n62178 , n62236 );
or ( n62238 , n62177 , n62237 );
and ( n62239 , n62174 , n62238 );
or ( n62240 , n62173 , n62239 );
and ( n62241 , n62170 , n62240 );
or ( n62242 , n62169 , n62241 );
and ( n62243 , n62166 , n62242 );
or ( n62244 , n62165 , n62243 );
and ( n62245 , n62162 , n62244 );
or ( n62246 , n62161 , n62245 );
and ( n62247 , n62158 , n62246 );
or ( n62248 , n62157 , n62247 );
and ( n62249 , n62154 , n62248 );
or ( n62250 , n62153 , n62249 );
and ( n62251 , n62150 , n62250 );
or ( n62252 , n62149 , n62251 );
and ( n62253 , n62146 , n62252 );
or ( n62254 , n62145 , n62253 );
and ( n62255 , n62142 , n62254 );
or ( n62256 , n62141 , n62255 );
and ( n62257 , n62138 , n62256 );
or ( n62258 , n62137 , n62257 );
and ( n62259 , n62134 , n62258 );
or ( n62260 , n62133 , n62259 );
and ( n62261 , n62130 , n62260 );
or ( n62262 , n62129 , n62261 );
and ( n62263 , n62126 , n62262 );
or ( n62264 , n62125 , n62263 );
and ( n62265 , n62122 , n62264 );
or ( n62266 , n62121 , n62265 );
and ( n62267 , n62118 , n62266 );
or ( n62268 , n62117 , n62267 );
and ( n62269 , n62114 , n62268 );
or ( n62270 , n62113 , n62269 );
and ( n62271 , n62110 , n62270 );
or ( n62272 , n62109 , n62271 );
and ( n62273 , n62106 , n62272 );
or ( n62274 , n62105 , n62273 );
and ( n62275 , n62102 , n62274 );
or ( n62276 , n62101 , n62275 );
and ( n62277 , n62098 , n62276 );
or ( n62278 , n62097 , n62277 );
and ( n62279 , n62094 , n62278 );
or ( n62280 , n62093 , n62279 );
and ( n62281 , n62090 , n62280 );
or ( n62282 , n62089 , n62281 );
and ( n62283 , n62086 , n62282 );
or ( n62284 , n62085 , n62283 );
and ( n62285 , n62082 , n62284 );
or ( n62286 , n62081 , n62285 );
and ( n62287 , n62078 , n62286 );
or ( n62288 , n62077 , n62287 );
and ( n62289 , n62074 , n62288 );
or ( n62290 , n62073 , n62289 );
and ( n62291 , n62070 , n62290 );
or ( n62292 , n62069 , n62291 );
and ( n62293 , n62066 , n62292 );
or ( n62294 , n62065 , n62293 );
and ( n62295 , n62062 , n62294 );
or ( n62296 , n62061 , n62295 );
and ( n62297 , n62058 , n62296 );
or ( n62298 , n62057 , n62297 );
and ( n62299 , n62054 , n62298 );
or ( n62300 , n62053 , n62299 );
and ( n62301 , n62050 , n62300 );
or ( n62302 , n62049 , n62301 );
and ( n62303 , n62046 , n62302 );
or ( n62304 , n62045 , n62303 );
and ( n62305 , n62042 , n62304 );
or ( n62306 , n62041 , n62305 );
and ( n62307 , n62038 , n62306 );
or ( n62308 , n62037 , n62307 );
and ( n62309 , n62034 , n62308 );
or ( n62310 , n62033 , n62309 );
and ( n62311 , n62030 , n62310 );
or ( n62312 , n62029 , n62311 );
and ( n62313 , n62026 , n62312 );
or ( n62314 , n62025 , n62313 );
and ( n62315 , n62022 , n62314 );
or ( n62316 , n62021 , n62315 );
and ( n62317 , n62018 , n62316 );
or ( n62318 , n62017 , n62317 );
and ( n62319 , n62014 , n62318 );
or ( n62320 , n62013 , n62319 );
and ( n62321 , n62010 , n62320 );
or ( n62322 , n62009 , n62321 );
and ( n62323 , n62006 , n62322 );
or ( n62324 , n62005 , n62323 );
and ( n62325 , n62002 , n62324 );
or ( n62326 , n62001 , n62325 );
and ( n62327 , n61998 , n62326 );
or ( n62328 , n61997 , n62327 );
and ( n62329 , n61994 , n62328 );
or ( n62330 , n61993 , n62329 );
and ( n62331 , n61990 , n62330 );
or ( n62332 , n61989 , n62331 );
and ( n62333 , n61986 , n62332 );
or ( n62334 , n61985 , n62333 );
and ( n62335 , n61982 , n62334 );
or ( n62336 , n61981 , n62335 );
and ( n62337 , n61978 , n62336 );
or ( n62338 , n61977 , n62337 );
and ( n62339 , n61974 , n62338 );
or ( n62340 , n61973 , n62339 );
and ( n62341 , n61970 , n62340 );
or ( n62342 , n61969 , n62341 );
and ( n62343 , n61966 , n62342 );
or ( n62344 , n61965 , n62343 );
and ( n62345 , n61962 , n62344 );
or ( n62346 , n61961 , n62345 );
and ( n62347 , n61958 , n62346 );
or ( n62348 , n61957 , n62347 );
and ( n62349 , n61954 , n62348 );
or ( n62350 , n61953 , n62349 );
and ( n62351 , n61950 , n62350 );
or ( n62352 , n61949 , n62351 );
and ( n62353 , n61946 , n62352 );
or ( n62354 , n61945 , n62353 );
and ( n62355 , n61942 , n62354 );
or ( n62356 , n61941 , n62355 );
and ( n62357 , n61938 , n62356 );
or ( n62358 , n61937 , n62357 );
xor ( n62359 , n61934 , n62358 );
buf ( n62360 , n17994 );
and ( n62361 , n30059 , n62360 );
xor ( n62362 , n62359 , n62361 );
xor ( n62363 , n61938 , n62356 );
and ( n62364 , n30064 , n62360 );
and ( n62365 , n62363 , n62364 );
xor ( n62366 , n62363 , n62364 );
xor ( n62367 , n61942 , n62354 );
and ( n62368 , n30069 , n62360 );
and ( n62369 , n62367 , n62368 );
xor ( n62370 , n62367 , n62368 );
xor ( n62371 , n61946 , n62352 );
and ( n62372 , n30074 , n62360 );
and ( n62373 , n62371 , n62372 );
xor ( n62374 , n62371 , n62372 );
xor ( n62375 , n61950 , n62350 );
and ( n62376 , n30079 , n62360 );
and ( n62377 , n62375 , n62376 );
xor ( n62378 , n62375 , n62376 );
xor ( n62379 , n61954 , n62348 );
and ( n62380 , n30084 , n62360 );
and ( n62381 , n62379 , n62380 );
xor ( n62382 , n62379 , n62380 );
xor ( n62383 , n61958 , n62346 );
and ( n62384 , n30089 , n62360 );
and ( n62385 , n62383 , n62384 );
xor ( n62386 , n62383 , n62384 );
xor ( n62387 , n61962 , n62344 );
and ( n62388 , n30094 , n62360 );
and ( n62389 , n62387 , n62388 );
xor ( n62390 , n62387 , n62388 );
xor ( n62391 , n61966 , n62342 );
and ( n62392 , n30099 , n62360 );
and ( n62393 , n62391 , n62392 );
xor ( n62394 , n62391 , n62392 );
xor ( n62395 , n61970 , n62340 );
and ( n62396 , n30104 , n62360 );
and ( n62397 , n62395 , n62396 );
xor ( n62398 , n62395 , n62396 );
xor ( n62399 , n61974 , n62338 );
and ( n62400 , n30109 , n62360 );
and ( n62401 , n62399 , n62400 );
xor ( n62402 , n62399 , n62400 );
xor ( n62403 , n61978 , n62336 );
and ( n62404 , n30114 , n62360 );
and ( n62405 , n62403 , n62404 );
xor ( n62406 , n62403 , n62404 );
xor ( n62407 , n61982 , n62334 );
and ( n62408 , n30119 , n62360 );
and ( n62409 , n62407 , n62408 );
xor ( n62410 , n62407 , n62408 );
xor ( n62411 , n61986 , n62332 );
and ( n62412 , n30124 , n62360 );
and ( n62413 , n62411 , n62412 );
xor ( n62414 , n62411 , n62412 );
xor ( n62415 , n61990 , n62330 );
and ( n62416 , n30129 , n62360 );
and ( n62417 , n62415 , n62416 );
xor ( n62418 , n62415 , n62416 );
xor ( n62419 , n61994 , n62328 );
and ( n62420 , n30134 , n62360 );
and ( n62421 , n62419 , n62420 );
xor ( n62422 , n62419 , n62420 );
xor ( n62423 , n61998 , n62326 );
and ( n62424 , n30139 , n62360 );
and ( n62425 , n62423 , n62424 );
xor ( n62426 , n62423 , n62424 );
xor ( n62427 , n62002 , n62324 );
and ( n62428 , n30144 , n62360 );
and ( n62429 , n62427 , n62428 );
xor ( n62430 , n62427 , n62428 );
xor ( n62431 , n62006 , n62322 );
and ( n62432 , n30149 , n62360 );
and ( n62433 , n62431 , n62432 );
xor ( n62434 , n62431 , n62432 );
xor ( n62435 , n62010 , n62320 );
and ( n62436 , n30154 , n62360 );
and ( n62437 , n62435 , n62436 );
xor ( n62438 , n62435 , n62436 );
xor ( n62439 , n62014 , n62318 );
and ( n62440 , n30159 , n62360 );
and ( n62441 , n62439 , n62440 );
xor ( n62442 , n62439 , n62440 );
xor ( n62443 , n62018 , n62316 );
and ( n62444 , n30164 , n62360 );
and ( n62445 , n62443 , n62444 );
xor ( n62446 , n62443 , n62444 );
xor ( n62447 , n62022 , n62314 );
and ( n62448 , n30169 , n62360 );
and ( n62449 , n62447 , n62448 );
xor ( n62450 , n62447 , n62448 );
xor ( n62451 , n62026 , n62312 );
and ( n62452 , n30174 , n62360 );
and ( n62453 , n62451 , n62452 );
xor ( n62454 , n62451 , n62452 );
xor ( n62455 , n62030 , n62310 );
and ( n62456 , n30179 , n62360 );
and ( n62457 , n62455 , n62456 );
xor ( n62458 , n62455 , n62456 );
xor ( n62459 , n62034 , n62308 );
and ( n62460 , n30184 , n62360 );
and ( n62461 , n62459 , n62460 );
xor ( n62462 , n62459 , n62460 );
xor ( n62463 , n62038 , n62306 );
and ( n62464 , n30189 , n62360 );
and ( n62465 , n62463 , n62464 );
xor ( n62466 , n62463 , n62464 );
xor ( n62467 , n62042 , n62304 );
and ( n62468 , n30194 , n62360 );
and ( n62469 , n62467 , n62468 );
xor ( n62470 , n62467 , n62468 );
xor ( n62471 , n62046 , n62302 );
and ( n62472 , n30199 , n62360 );
and ( n62473 , n62471 , n62472 );
xor ( n62474 , n62471 , n62472 );
xor ( n62475 , n62050 , n62300 );
and ( n62476 , n30204 , n62360 );
and ( n62477 , n62475 , n62476 );
xor ( n62478 , n62475 , n62476 );
xor ( n62479 , n62054 , n62298 );
and ( n62480 , n30209 , n62360 );
and ( n62481 , n62479 , n62480 );
xor ( n62482 , n62479 , n62480 );
xor ( n62483 , n62058 , n62296 );
and ( n62484 , n30214 , n62360 );
and ( n62485 , n62483 , n62484 );
xor ( n62486 , n62483 , n62484 );
xor ( n62487 , n62062 , n62294 );
and ( n62488 , n30219 , n62360 );
and ( n62489 , n62487 , n62488 );
xor ( n62490 , n62487 , n62488 );
xor ( n62491 , n62066 , n62292 );
and ( n62492 , n30224 , n62360 );
and ( n62493 , n62491 , n62492 );
xor ( n62494 , n62491 , n62492 );
xor ( n62495 , n62070 , n62290 );
and ( n62496 , n30229 , n62360 );
and ( n62497 , n62495 , n62496 );
xor ( n62498 , n62495 , n62496 );
xor ( n62499 , n62074 , n62288 );
and ( n62500 , n30234 , n62360 );
and ( n62501 , n62499 , n62500 );
xor ( n62502 , n62499 , n62500 );
xor ( n62503 , n62078 , n62286 );
and ( n62504 , n30239 , n62360 );
and ( n62505 , n62503 , n62504 );
xor ( n62506 , n62503 , n62504 );
xor ( n62507 , n62082 , n62284 );
and ( n62508 , n30244 , n62360 );
and ( n62509 , n62507 , n62508 );
xor ( n62510 , n62507 , n62508 );
xor ( n62511 , n62086 , n62282 );
and ( n62512 , n30249 , n62360 );
and ( n62513 , n62511 , n62512 );
xor ( n62514 , n62511 , n62512 );
xor ( n62515 , n62090 , n62280 );
and ( n62516 , n30254 , n62360 );
and ( n62517 , n62515 , n62516 );
xor ( n62518 , n62515 , n62516 );
xor ( n62519 , n62094 , n62278 );
and ( n62520 , n30259 , n62360 );
and ( n62521 , n62519 , n62520 );
xor ( n62522 , n62519 , n62520 );
xor ( n62523 , n62098 , n62276 );
and ( n62524 , n30264 , n62360 );
and ( n62525 , n62523 , n62524 );
xor ( n62526 , n62523 , n62524 );
xor ( n62527 , n62102 , n62274 );
and ( n62528 , n30269 , n62360 );
and ( n62529 , n62527 , n62528 );
xor ( n62530 , n62527 , n62528 );
xor ( n62531 , n62106 , n62272 );
and ( n62532 , n30274 , n62360 );
and ( n62533 , n62531 , n62532 );
xor ( n62534 , n62531 , n62532 );
xor ( n62535 , n62110 , n62270 );
and ( n62536 , n30279 , n62360 );
and ( n62537 , n62535 , n62536 );
xor ( n62538 , n62535 , n62536 );
xor ( n62539 , n62114 , n62268 );
and ( n62540 , n30284 , n62360 );
and ( n62541 , n62539 , n62540 );
xor ( n62542 , n62539 , n62540 );
xor ( n62543 , n62118 , n62266 );
and ( n62544 , n30289 , n62360 );
and ( n62545 , n62543 , n62544 );
xor ( n62546 , n62543 , n62544 );
xor ( n62547 , n62122 , n62264 );
and ( n62548 , n30294 , n62360 );
and ( n62549 , n62547 , n62548 );
xor ( n62550 , n62547 , n62548 );
xor ( n62551 , n62126 , n62262 );
and ( n62552 , n30299 , n62360 );
and ( n62553 , n62551 , n62552 );
xor ( n62554 , n62551 , n62552 );
xor ( n62555 , n62130 , n62260 );
and ( n62556 , n30304 , n62360 );
and ( n62557 , n62555 , n62556 );
xor ( n62558 , n62555 , n62556 );
xor ( n62559 , n62134 , n62258 );
and ( n62560 , n30309 , n62360 );
and ( n62561 , n62559 , n62560 );
xor ( n62562 , n62559 , n62560 );
xor ( n62563 , n62138 , n62256 );
and ( n62564 , n30314 , n62360 );
and ( n62565 , n62563 , n62564 );
xor ( n62566 , n62563 , n62564 );
xor ( n62567 , n62142 , n62254 );
and ( n62568 , n30319 , n62360 );
and ( n62569 , n62567 , n62568 );
xor ( n62570 , n62567 , n62568 );
xor ( n62571 , n62146 , n62252 );
and ( n62572 , n30324 , n62360 );
and ( n62573 , n62571 , n62572 );
xor ( n62574 , n62571 , n62572 );
xor ( n62575 , n62150 , n62250 );
and ( n62576 , n30329 , n62360 );
and ( n62577 , n62575 , n62576 );
xor ( n62578 , n62575 , n62576 );
xor ( n62579 , n62154 , n62248 );
and ( n62580 , n30334 , n62360 );
and ( n62581 , n62579 , n62580 );
xor ( n62582 , n62579 , n62580 );
xor ( n62583 , n62158 , n62246 );
and ( n62584 , n30339 , n62360 );
and ( n62585 , n62583 , n62584 );
xor ( n62586 , n62583 , n62584 );
xor ( n62587 , n62162 , n62244 );
and ( n62588 , n30344 , n62360 );
and ( n62589 , n62587 , n62588 );
xor ( n62590 , n62587 , n62588 );
xor ( n62591 , n62166 , n62242 );
and ( n62592 , n30349 , n62360 );
and ( n62593 , n62591 , n62592 );
xor ( n62594 , n62591 , n62592 );
xor ( n62595 , n62170 , n62240 );
and ( n62596 , n30354 , n62360 );
and ( n62597 , n62595 , n62596 );
xor ( n62598 , n62595 , n62596 );
xor ( n62599 , n62174 , n62238 );
and ( n62600 , n30359 , n62360 );
and ( n62601 , n62599 , n62600 );
xor ( n62602 , n62599 , n62600 );
xor ( n62603 , n62178 , n62236 );
and ( n62604 , n30364 , n62360 );
and ( n62605 , n62603 , n62604 );
xor ( n62606 , n62603 , n62604 );
xor ( n62607 , n62182 , n62234 );
and ( n62608 , n30369 , n62360 );
and ( n62609 , n62607 , n62608 );
xor ( n62610 , n62607 , n62608 );
xor ( n62611 , n62186 , n62232 );
and ( n62612 , n30374 , n62360 );
and ( n62613 , n62611 , n62612 );
xor ( n62614 , n62611 , n62612 );
xor ( n62615 , n62190 , n62230 );
and ( n62616 , n30379 , n62360 );
and ( n62617 , n62615 , n62616 );
xor ( n62618 , n62615 , n62616 );
xor ( n62619 , n62194 , n62228 );
and ( n62620 , n30384 , n62360 );
and ( n62621 , n62619 , n62620 );
xor ( n62622 , n62619 , n62620 );
xor ( n62623 , n62198 , n62226 );
and ( n62624 , n30389 , n62360 );
and ( n62625 , n62623 , n62624 );
xor ( n62626 , n62623 , n62624 );
xor ( n62627 , n62202 , n62224 );
and ( n62628 , n30394 , n62360 );
and ( n62629 , n62627 , n62628 );
xor ( n62630 , n62627 , n62628 );
xor ( n62631 , n62206 , n62222 );
and ( n62632 , n30399 , n62360 );
and ( n62633 , n62631 , n62632 );
xor ( n62634 , n62631 , n62632 );
xor ( n62635 , n62210 , n62220 );
and ( n62636 , n30404 , n62360 );
and ( n62637 , n62635 , n62636 );
xor ( n62638 , n62635 , n62636 );
xor ( n62639 , n62214 , n62218 );
and ( n62640 , n30409 , n62360 );
and ( n62641 , n62639 , n62640 );
buf ( n62642 , n62641 );
and ( n62643 , n62638 , n62642 );
or ( n62644 , n62637 , n62643 );
and ( n62645 , n62634 , n62644 );
or ( n62646 , n62633 , n62645 );
and ( n62647 , n62630 , n62646 );
or ( n62648 , n62629 , n62647 );
and ( n62649 , n62626 , n62648 );
or ( n62650 , n62625 , n62649 );
and ( n62651 , n62622 , n62650 );
or ( n62652 , n62621 , n62651 );
and ( n62653 , n62618 , n62652 );
or ( n62654 , n62617 , n62653 );
and ( n62655 , n62614 , n62654 );
or ( n62656 , n62613 , n62655 );
and ( n62657 , n62610 , n62656 );
or ( n62658 , n62609 , n62657 );
and ( n62659 , n62606 , n62658 );
or ( n62660 , n62605 , n62659 );
and ( n62661 , n62602 , n62660 );
or ( n62662 , n62601 , n62661 );
and ( n62663 , n62598 , n62662 );
or ( n62664 , n62597 , n62663 );
and ( n62665 , n62594 , n62664 );
or ( n62666 , n62593 , n62665 );
and ( n62667 , n62590 , n62666 );
or ( n62668 , n62589 , n62667 );
and ( n62669 , n62586 , n62668 );
or ( n62670 , n62585 , n62669 );
and ( n62671 , n62582 , n62670 );
or ( n62672 , n62581 , n62671 );
and ( n62673 , n62578 , n62672 );
or ( n62674 , n62577 , n62673 );
and ( n62675 , n62574 , n62674 );
or ( n62676 , n62573 , n62675 );
and ( n62677 , n62570 , n62676 );
or ( n62678 , n62569 , n62677 );
and ( n62679 , n62566 , n62678 );
or ( n62680 , n62565 , n62679 );
and ( n62681 , n62562 , n62680 );
or ( n62682 , n62561 , n62681 );
and ( n62683 , n62558 , n62682 );
or ( n62684 , n62557 , n62683 );
and ( n62685 , n62554 , n62684 );
or ( n62686 , n62553 , n62685 );
and ( n62687 , n62550 , n62686 );
or ( n62688 , n62549 , n62687 );
and ( n62689 , n62546 , n62688 );
or ( n62690 , n62545 , n62689 );
and ( n62691 , n62542 , n62690 );
or ( n62692 , n62541 , n62691 );
and ( n62693 , n62538 , n62692 );
or ( n62694 , n62537 , n62693 );
and ( n62695 , n62534 , n62694 );
or ( n62696 , n62533 , n62695 );
and ( n62697 , n62530 , n62696 );
or ( n62698 , n62529 , n62697 );
and ( n62699 , n62526 , n62698 );
or ( n62700 , n62525 , n62699 );
and ( n62701 , n62522 , n62700 );
or ( n62702 , n62521 , n62701 );
and ( n62703 , n62518 , n62702 );
or ( n62704 , n62517 , n62703 );
and ( n62705 , n62514 , n62704 );
or ( n62706 , n62513 , n62705 );
and ( n62707 , n62510 , n62706 );
or ( n62708 , n62509 , n62707 );
and ( n62709 , n62506 , n62708 );
or ( n62710 , n62505 , n62709 );
and ( n62711 , n62502 , n62710 );
or ( n62712 , n62501 , n62711 );
and ( n62713 , n62498 , n62712 );
or ( n62714 , n62497 , n62713 );
and ( n62715 , n62494 , n62714 );
or ( n62716 , n62493 , n62715 );
and ( n62717 , n62490 , n62716 );
or ( n62718 , n62489 , n62717 );
and ( n62719 , n62486 , n62718 );
or ( n62720 , n62485 , n62719 );
and ( n62721 , n62482 , n62720 );
or ( n62722 , n62481 , n62721 );
and ( n62723 , n62478 , n62722 );
or ( n62724 , n62477 , n62723 );
and ( n62725 , n62474 , n62724 );
or ( n62726 , n62473 , n62725 );
and ( n62727 , n62470 , n62726 );
or ( n62728 , n62469 , n62727 );
and ( n62729 , n62466 , n62728 );
or ( n62730 , n62465 , n62729 );
and ( n62731 , n62462 , n62730 );
or ( n62732 , n62461 , n62731 );
and ( n62733 , n62458 , n62732 );
or ( n62734 , n62457 , n62733 );
and ( n62735 , n62454 , n62734 );
or ( n62736 , n62453 , n62735 );
and ( n62737 , n62450 , n62736 );
or ( n62738 , n62449 , n62737 );
and ( n62739 , n62446 , n62738 );
or ( n62740 , n62445 , n62739 );
and ( n62741 , n62442 , n62740 );
or ( n62742 , n62441 , n62741 );
and ( n62743 , n62438 , n62742 );
or ( n62744 , n62437 , n62743 );
and ( n62745 , n62434 , n62744 );
or ( n62746 , n62433 , n62745 );
and ( n62747 , n62430 , n62746 );
or ( n62748 , n62429 , n62747 );
and ( n62749 , n62426 , n62748 );
or ( n62750 , n62425 , n62749 );
and ( n62751 , n62422 , n62750 );
or ( n62752 , n62421 , n62751 );
and ( n62753 , n62418 , n62752 );
or ( n62754 , n62417 , n62753 );
and ( n62755 , n62414 , n62754 );
or ( n62756 , n62413 , n62755 );
and ( n62757 , n62410 , n62756 );
or ( n62758 , n62409 , n62757 );
and ( n62759 , n62406 , n62758 );
or ( n62760 , n62405 , n62759 );
and ( n62761 , n62402 , n62760 );
or ( n62762 , n62401 , n62761 );
and ( n62763 , n62398 , n62762 );
or ( n62764 , n62397 , n62763 );
and ( n62765 , n62394 , n62764 );
or ( n62766 , n62393 , n62765 );
and ( n62767 , n62390 , n62766 );
or ( n62768 , n62389 , n62767 );
and ( n62769 , n62386 , n62768 );
or ( n62770 , n62385 , n62769 );
and ( n62771 , n62382 , n62770 );
or ( n62772 , n62381 , n62771 );
and ( n62773 , n62378 , n62772 );
or ( n62774 , n62377 , n62773 );
and ( n62775 , n62374 , n62774 );
or ( n62776 , n62373 , n62775 );
and ( n62777 , n62370 , n62776 );
or ( n62778 , n62369 , n62777 );
and ( n62779 , n62366 , n62778 );
or ( n62780 , n62365 , n62779 );
xor ( n62781 , n62362 , n62780 );
buf ( n62782 , n17992 );
and ( n62783 , n30064 , n62782 );
xor ( n62784 , n62781 , n62783 );
xor ( n62785 , n62366 , n62778 );
and ( n62786 , n30069 , n62782 );
and ( n62787 , n62785 , n62786 );
xor ( n62788 , n62785 , n62786 );
xor ( n62789 , n62370 , n62776 );
and ( n62790 , n30074 , n62782 );
and ( n62791 , n62789 , n62790 );
xor ( n62792 , n62789 , n62790 );
xor ( n62793 , n62374 , n62774 );
and ( n62794 , n30079 , n62782 );
and ( n62795 , n62793 , n62794 );
xor ( n62796 , n62793 , n62794 );
xor ( n62797 , n62378 , n62772 );
and ( n62798 , n30084 , n62782 );
and ( n62799 , n62797 , n62798 );
xor ( n62800 , n62797 , n62798 );
xor ( n62801 , n62382 , n62770 );
and ( n62802 , n30089 , n62782 );
and ( n62803 , n62801 , n62802 );
xor ( n62804 , n62801 , n62802 );
xor ( n62805 , n62386 , n62768 );
and ( n62806 , n30094 , n62782 );
and ( n62807 , n62805 , n62806 );
xor ( n62808 , n62805 , n62806 );
xor ( n62809 , n62390 , n62766 );
and ( n62810 , n30099 , n62782 );
and ( n62811 , n62809 , n62810 );
xor ( n62812 , n62809 , n62810 );
xor ( n62813 , n62394 , n62764 );
and ( n62814 , n30104 , n62782 );
and ( n62815 , n62813 , n62814 );
xor ( n62816 , n62813 , n62814 );
xor ( n62817 , n62398 , n62762 );
and ( n62818 , n30109 , n62782 );
and ( n62819 , n62817 , n62818 );
xor ( n62820 , n62817 , n62818 );
xor ( n62821 , n62402 , n62760 );
and ( n62822 , n30114 , n62782 );
and ( n62823 , n62821 , n62822 );
xor ( n62824 , n62821 , n62822 );
xor ( n62825 , n62406 , n62758 );
and ( n62826 , n30119 , n62782 );
and ( n62827 , n62825 , n62826 );
xor ( n62828 , n62825 , n62826 );
xor ( n62829 , n62410 , n62756 );
and ( n62830 , n30124 , n62782 );
and ( n62831 , n62829 , n62830 );
xor ( n62832 , n62829 , n62830 );
xor ( n62833 , n62414 , n62754 );
and ( n62834 , n30129 , n62782 );
and ( n62835 , n62833 , n62834 );
xor ( n62836 , n62833 , n62834 );
xor ( n62837 , n62418 , n62752 );
and ( n62838 , n30134 , n62782 );
and ( n62839 , n62837 , n62838 );
xor ( n62840 , n62837 , n62838 );
xor ( n62841 , n62422 , n62750 );
and ( n62842 , n30139 , n62782 );
and ( n62843 , n62841 , n62842 );
xor ( n62844 , n62841 , n62842 );
xor ( n62845 , n62426 , n62748 );
and ( n62846 , n30144 , n62782 );
and ( n62847 , n62845 , n62846 );
xor ( n62848 , n62845 , n62846 );
xor ( n62849 , n62430 , n62746 );
and ( n62850 , n30149 , n62782 );
and ( n62851 , n62849 , n62850 );
xor ( n62852 , n62849 , n62850 );
xor ( n62853 , n62434 , n62744 );
and ( n62854 , n30154 , n62782 );
and ( n62855 , n62853 , n62854 );
xor ( n62856 , n62853 , n62854 );
xor ( n62857 , n62438 , n62742 );
and ( n62858 , n30159 , n62782 );
and ( n62859 , n62857 , n62858 );
xor ( n62860 , n62857 , n62858 );
xor ( n62861 , n62442 , n62740 );
and ( n62862 , n30164 , n62782 );
and ( n62863 , n62861 , n62862 );
xor ( n62864 , n62861 , n62862 );
xor ( n62865 , n62446 , n62738 );
and ( n62866 , n30169 , n62782 );
and ( n62867 , n62865 , n62866 );
xor ( n62868 , n62865 , n62866 );
xor ( n62869 , n62450 , n62736 );
and ( n62870 , n30174 , n62782 );
and ( n62871 , n62869 , n62870 );
xor ( n62872 , n62869 , n62870 );
xor ( n62873 , n62454 , n62734 );
and ( n62874 , n30179 , n62782 );
and ( n62875 , n62873 , n62874 );
xor ( n62876 , n62873 , n62874 );
xor ( n62877 , n62458 , n62732 );
and ( n62878 , n30184 , n62782 );
and ( n62879 , n62877 , n62878 );
xor ( n62880 , n62877 , n62878 );
xor ( n62881 , n62462 , n62730 );
and ( n62882 , n30189 , n62782 );
and ( n62883 , n62881 , n62882 );
xor ( n62884 , n62881 , n62882 );
xor ( n62885 , n62466 , n62728 );
and ( n62886 , n30194 , n62782 );
and ( n62887 , n62885 , n62886 );
xor ( n62888 , n62885 , n62886 );
xor ( n62889 , n62470 , n62726 );
and ( n62890 , n30199 , n62782 );
and ( n62891 , n62889 , n62890 );
xor ( n62892 , n62889 , n62890 );
xor ( n62893 , n62474 , n62724 );
and ( n62894 , n30204 , n62782 );
and ( n62895 , n62893 , n62894 );
xor ( n62896 , n62893 , n62894 );
xor ( n62897 , n62478 , n62722 );
and ( n62898 , n30209 , n62782 );
and ( n62899 , n62897 , n62898 );
xor ( n62900 , n62897 , n62898 );
xor ( n62901 , n62482 , n62720 );
and ( n62902 , n30214 , n62782 );
and ( n62903 , n62901 , n62902 );
xor ( n62904 , n62901 , n62902 );
xor ( n62905 , n62486 , n62718 );
and ( n62906 , n30219 , n62782 );
and ( n62907 , n62905 , n62906 );
xor ( n62908 , n62905 , n62906 );
xor ( n62909 , n62490 , n62716 );
and ( n62910 , n30224 , n62782 );
and ( n62911 , n62909 , n62910 );
xor ( n62912 , n62909 , n62910 );
xor ( n62913 , n62494 , n62714 );
and ( n62914 , n30229 , n62782 );
and ( n62915 , n62913 , n62914 );
xor ( n62916 , n62913 , n62914 );
xor ( n62917 , n62498 , n62712 );
and ( n62918 , n30234 , n62782 );
and ( n62919 , n62917 , n62918 );
xor ( n62920 , n62917 , n62918 );
xor ( n62921 , n62502 , n62710 );
and ( n62922 , n30239 , n62782 );
and ( n62923 , n62921 , n62922 );
xor ( n62924 , n62921 , n62922 );
xor ( n62925 , n62506 , n62708 );
and ( n62926 , n30244 , n62782 );
and ( n62927 , n62925 , n62926 );
xor ( n62928 , n62925 , n62926 );
xor ( n62929 , n62510 , n62706 );
and ( n62930 , n30249 , n62782 );
and ( n62931 , n62929 , n62930 );
xor ( n62932 , n62929 , n62930 );
xor ( n62933 , n62514 , n62704 );
and ( n62934 , n30254 , n62782 );
and ( n62935 , n62933 , n62934 );
xor ( n62936 , n62933 , n62934 );
xor ( n62937 , n62518 , n62702 );
and ( n62938 , n30259 , n62782 );
and ( n62939 , n62937 , n62938 );
xor ( n62940 , n62937 , n62938 );
xor ( n62941 , n62522 , n62700 );
and ( n62942 , n30264 , n62782 );
and ( n62943 , n62941 , n62942 );
xor ( n62944 , n62941 , n62942 );
xor ( n62945 , n62526 , n62698 );
and ( n62946 , n30269 , n62782 );
and ( n62947 , n62945 , n62946 );
xor ( n62948 , n62945 , n62946 );
xor ( n62949 , n62530 , n62696 );
and ( n62950 , n30274 , n62782 );
and ( n62951 , n62949 , n62950 );
xor ( n62952 , n62949 , n62950 );
xor ( n62953 , n62534 , n62694 );
and ( n62954 , n30279 , n62782 );
and ( n62955 , n62953 , n62954 );
xor ( n62956 , n62953 , n62954 );
xor ( n62957 , n62538 , n62692 );
and ( n62958 , n30284 , n62782 );
and ( n62959 , n62957 , n62958 );
xor ( n62960 , n62957 , n62958 );
xor ( n62961 , n62542 , n62690 );
and ( n62962 , n30289 , n62782 );
and ( n62963 , n62961 , n62962 );
xor ( n62964 , n62961 , n62962 );
xor ( n62965 , n62546 , n62688 );
and ( n62966 , n30294 , n62782 );
and ( n62967 , n62965 , n62966 );
xor ( n62968 , n62965 , n62966 );
xor ( n62969 , n62550 , n62686 );
and ( n62970 , n30299 , n62782 );
and ( n62971 , n62969 , n62970 );
xor ( n62972 , n62969 , n62970 );
xor ( n62973 , n62554 , n62684 );
and ( n62974 , n30304 , n62782 );
and ( n62975 , n62973 , n62974 );
xor ( n62976 , n62973 , n62974 );
xor ( n62977 , n62558 , n62682 );
and ( n62978 , n30309 , n62782 );
and ( n62979 , n62977 , n62978 );
xor ( n62980 , n62977 , n62978 );
xor ( n62981 , n62562 , n62680 );
and ( n62982 , n30314 , n62782 );
and ( n62983 , n62981 , n62982 );
xor ( n62984 , n62981 , n62982 );
xor ( n62985 , n62566 , n62678 );
and ( n62986 , n30319 , n62782 );
and ( n62987 , n62985 , n62986 );
xor ( n62988 , n62985 , n62986 );
xor ( n62989 , n62570 , n62676 );
and ( n62990 , n30324 , n62782 );
and ( n62991 , n62989 , n62990 );
xor ( n62992 , n62989 , n62990 );
xor ( n62993 , n62574 , n62674 );
and ( n62994 , n30329 , n62782 );
and ( n62995 , n62993 , n62994 );
xor ( n62996 , n62993 , n62994 );
xor ( n62997 , n62578 , n62672 );
and ( n62998 , n30334 , n62782 );
and ( n62999 , n62997 , n62998 );
xor ( n63000 , n62997 , n62998 );
xor ( n63001 , n62582 , n62670 );
and ( n63002 , n30339 , n62782 );
and ( n63003 , n63001 , n63002 );
xor ( n63004 , n63001 , n63002 );
xor ( n63005 , n62586 , n62668 );
and ( n63006 , n30344 , n62782 );
and ( n63007 , n63005 , n63006 );
xor ( n63008 , n63005 , n63006 );
xor ( n63009 , n62590 , n62666 );
and ( n63010 , n30349 , n62782 );
and ( n63011 , n63009 , n63010 );
xor ( n63012 , n63009 , n63010 );
xor ( n63013 , n62594 , n62664 );
and ( n63014 , n30354 , n62782 );
and ( n63015 , n63013 , n63014 );
xor ( n63016 , n63013 , n63014 );
xor ( n63017 , n62598 , n62662 );
and ( n63018 , n30359 , n62782 );
and ( n63019 , n63017 , n63018 );
xor ( n63020 , n63017 , n63018 );
xor ( n63021 , n62602 , n62660 );
and ( n63022 , n30364 , n62782 );
and ( n63023 , n63021 , n63022 );
xor ( n63024 , n63021 , n63022 );
xor ( n63025 , n62606 , n62658 );
and ( n63026 , n30369 , n62782 );
and ( n63027 , n63025 , n63026 );
xor ( n63028 , n63025 , n63026 );
xor ( n63029 , n62610 , n62656 );
and ( n63030 , n30374 , n62782 );
and ( n63031 , n63029 , n63030 );
xor ( n63032 , n63029 , n63030 );
xor ( n63033 , n62614 , n62654 );
and ( n63034 , n30379 , n62782 );
and ( n63035 , n63033 , n63034 );
xor ( n63036 , n63033 , n63034 );
xor ( n63037 , n62618 , n62652 );
and ( n63038 , n30384 , n62782 );
and ( n63039 , n63037 , n63038 );
xor ( n63040 , n63037 , n63038 );
xor ( n63041 , n62622 , n62650 );
and ( n63042 , n30389 , n62782 );
and ( n63043 , n63041 , n63042 );
xor ( n63044 , n63041 , n63042 );
xor ( n63045 , n62626 , n62648 );
and ( n63046 , n30394 , n62782 );
and ( n63047 , n63045 , n63046 );
xor ( n63048 , n63045 , n63046 );
xor ( n63049 , n62630 , n62646 );
and ( n63050 , n30399 , n62782 );
and ( n63051 , n63049 , n63050 );
xor ( n63052 , n63049 , n63050 );
xor ( n63053 , n62634 , n62644 );
and ( n63054 , n30404 , n62782 );
and ( n63055 , n63053 , n63054 );
xor ( n63056 , n63053 , n63054 );
xor ( n63057 , n62638 , n62642 );
and ( n63058 , n30409 , n62782 );
and ( n63059 , n63057 , n63058 );
buf ( n63060 , n63059 );
and ( n63061 , n63056 , n63060 );
or ( n63062 , n63055 , n63061 );
and ( n63063 , n63052 , n63062 );
or ( n63064 , n63051 , n63063 );
and ( n63065 , n63048 , n63064 );
or ( n63066 , n63047 , n63065 );
and ( n63067 , n63044 , n63066 );
or ( n63068 , n63043 , n63067 );
and ( n63069 , n63040 , n63068 );
or ( n63070 , n63039 , n63069 );
and ( n63071 , n63036 , n63070 );
or ( n63072 , n63035 , n63071 );
and ( n63073 , n63032 , n63072 );
or ( n63074 , n63031 , n63073 );
and ( n63075 , n63028 , n63074 );
or ( n63076 , n63027 , n63075 );
and ( n63077 , n63024 , n63076 );
or ( n63078 , n63023 , n63077 );
and ( n63079 , n63020 , n63078 );
or ( n63080 , n63019 , n63079 );
and ( n63081 , n63016 , n63080 );
or ( n63082 , n63015 , n63081 );
and ( n63083 , n63012 , n63082 );
or ( n63084 , n63011 , n63083 );
and ( n63085 , n63008 , n63084 );
or ( n63086 , n63007 , n63085 );
and ( n63087 , n63004 , n63086 );
or ( n63088 , n63003 , n63087 );
and ( n63089 , n63000 , n63088 );
or ( n63090 , n62999 , n63089 );
and ( n63091 , n62996 , n63090 );
or ( n63092 , n62995 , n63091 );
and ( n63093 , n62992 , n63092 );
or ( n63094 , n62991 , n63093 );
and ( n63095 , n62988 , n63094 );
or ( n63096 , n62987 , n63095 );
and ( n63097 , n62984 , n63096 );
or ( n63098 , n62983 , n63097 );
and ( n63099 , n62980 , n63098 );
or ( n63100 , n62979 , n63099 );
and ( n63101 , n62976 , n63100 );
or ( n63102 , n62975 , n63101 );
and ( n63103 , n62972 , n63102 );
or ( n63104 , n62971 , n63103 );
and ( n63105 , n62968 , n63104 );
or ( n63106 , n62967 , n63105 );
and ( n63107 , n62964 , n63106 );
or ( n63108 , n62963 , n63107 );
and ( n63109 , n62960 , n63108 );
or ( n63110 , n62959 , n63109 );
and ( n63111 , n62956 , n63110 );
or ( n63112 , n62955 , n63111 );
and ( n63113 , n62952 , n63112 );
or ( n63114 , n62951 , n63113 );
and ( n63115 , n62948 , n63114 );
or ( n63116 , n62947 , n63115 );
and ( n63117 , n62944 , n63116 );
or ( n63118 , n62943 , n63117 );
and ( n63119 , n62940 , n63118 );
or ( n63120 , n62939 , n63119 );
and ( n63121 , n62936 , n63120 );
or ( n63122 , n62935 , n63121 );
and ( n63123 , n62932 , n63122 );
or ( n63124 , n62931 , n63123 );
and ( n63125 , n62928 , n63124 );
or ( n63126 , n62927 , n63125 );
and ( n63127 , n62924 , n63126 );
or ( n63128 , n62923 , n63127 );
and ( n63129 , n62920 , n63128 );
or ( n63130 , n62919 , n63129 );
and ( n63131 , n62916 , n63130 );
or ( n63132 , n62915 , n63131 );
and ( n63133 , n62912 , n63132 );
or ( n63134 , n62911 , n63133 );
and ( n63135 , n62908 , n63134 );
or ( n63136 , n62907 , n63135 );
and ( n63137 , n62904 , n63136 );
or ( n63138 , n62903 , n63137 );
and ( n63139 , n62900 , n63138 );
or ( n63140 , n62899 , n63139 );
and ( n63141 , n62896 , n63140 );
or ( n63142 , n62895 , n63141 );
and ( n63143 , n62892 , n63142 );
or ( n63144 , n62891 , n63143 );
and ( n63145 , n62888 , n63144 );
or ( n63146 , n62887 , n63145 );
and ( n63147 , n62884 , n63146 );
or ( n63148 , n62883 , n63147 );
and ( n63149 , n62880 , n63148 );
or ( n63150 , n62879 , n63149 );
and ( n63151 , n62876 , n63150 );
or ( n63152 , n62875 , n63151 );
and ( n63153 , n62872 , n63152 );
or ( n63154 , n62871 , n63153 );
and ( n63155 , n62868 , n63154 );
or ( n63156 , n62867 , n63155 );
and ( n63157 , n62864 , n63156 );
or ( n63158 , n62863 , n63157 );
and ( n63159 , n62860 , n63158 );
or ( n63160 , n62859 , n63159 );
and ( n63161 , n62856 , n63160 );
or ( n63162 , n62855 , n63161 );
and ( n63163 , n62852 , n63162 );
or ( n63164 , n62851 , n63163 );
and ( n63165 , n62848 , n63164 );
or ( n63166 , n62847 , n63165 );
and ( n63167 , n62844 , n63166 );
or ( n63168 , n62843 , n63167 );
and ( n63169 , n62840 , n63168 );
or ( n63170 , n62839 , n63169 );
and ( n63171 , n62836 , n63170 );
or ( n63172 , n62835 , n63171 );
and ( n63173 , n62832 , n63172 );
or ( n63174 , n62831 , n63173 );
and ( n63175 , n62828 , n63174 );
or ( n63176 , n62827 , n63175 );
and ( n63177 , n62824 , n63176 );
or ( n63178 , n62823 , n63177 );
and ( n63179 , n62820 , n63178 );
or ( n63180 , n62819 , n63179 );
and ( n63181 , n62816 , n63180 );
or ( n63182 , n62815 , n63181 );
and ( n63183 , n62812 , n63182 );
or ( n63184 , n62811 , n63183 );
and ( n63185 , n62808 , n63184 );
or ( n63186 , n62807 , n63185 );
and ( n63187 , n62804 , n63186 );
or ( n63188 , n62803 , n63187 );
and ( n63189 , n62800 , n63188 );
or ( n63190 , n62799 , n63189 );
and ( n63191 , n62796 , n63190 );
or ( n63192 , n62795 , n63191 );
and ( n63193 , n62792 , n63192 );
or ( n63194 , n62791 , n63193 );
and ( n63195 , n62788 , n63194 );
or ( n63196 , n62787 , n63195 );
xor ( n63197 , n62784 , n63196 );
buf ( n63198 , n17990 );
and ( n63199 , n30069 , n63198 );
xor ( n63200 , n63197 , n63199 );
xor ( n63201 , n62788 , n63194 );
and ( n63202 , n30074 , n63198 );
and ( n63203 , n63201 , n63202 );
xor ( n63204 , n63201 , n63202 );
xor ( n63205 , n62792 , n63192 );
and ( n63206 , n30079 , n63198 );
and ( n63207 , n63205 , n63206 );
xor ( n63208 , n63205 , n63206 );
xor ( n63209 , n62796 , n63190 );
and ( n63210 , n30084 , n63198 );
and ( n63211 , n63209 , n63210 );
xor ( n63212 , n63209 , n63210 );
xor ( n63213 , n62800 , n63188 );
and ( n63214 , n30089 , n63198 );
and ( n63215 , n63213 , n63214 );
xor ( n63216 , n63213 , n63214 );
xor ( n63217 , n62804 , n63186 );
and ( n63218 , n30094 , n63198 );
and ( n63219 , n63217 , n63218 );
xor ( n63220 , n63217 , n63218 );
xor ( n63221 , n62808 , n63184 );
and ( n63222 , n30099 , n63198 );
and ( n63223 , n63221 , n63222 );
xor ( n63224 , n63221 , n63222 );
xor ( n63225 , n62812 , n63182 );
and ( n63226 , n30104 , n63198 );
and ( n63227 , n63225 , n63226 );
xor ( n63228 , n63225 , n63226 );
xor ( n63229 , n62816 , n63180 );
and ( n63230 , n30109 , n63198 );
and ( n63231 , n63229 , n63230 );
xor ( n63232 , n63229 , n63230 );
xor ( n63233 , n62820 , n63178 );
and ( n63234 , n30114 , n63198 );
and ( n63235 , n63233 , n63234 );
xor ( n63236 , n63233 , n63234 );
xor ( n63237 , n62824 , n63176 );
and ( n63238 , n30119 , n63198 );
and ( n63239 , n63237 , n63238 );
xor ( n63240 , n63237 , n63238 );
xor ( n63241 , n62828 , n63174 );
and ( n63242 , n30124 , n63198 );
and ( n63243 , n63241 , n63242 );
xor ( n63244 , n63241 , n63242 );
xor ( n63245 , n62832 , n63172 );
and ( n63246 , n30129 , n63198 );
and ( n63247 , n63245 , n63246 );
xor ( n63248 , n63245 , n63246 );
xor ( n63249 , n62836 , n63170 );
and ( n63250 , n30134 , n63198 );
and ( n63251 , n63249 , n63250 );
xor ( n63252 , n63249 , n63250 );
xor ( n63253 , n62840 , n63168 );
and ( n63254 , n30139 , n63198 );
and ( n63255 , n63253 , n63254 );
xor ( n63256 , n63253 , n63254 );
xor ( n63257 , n62844 , n63166 );
and ( n63258 , n30144 , n63198 );
and ( n63259 , n63257 , n63258 );
xor ( n63260 , n63257 , n63258 );
xor ( n63261 , n62848 , n63164 );
and ( n63262 , n30149 , n63198 );
and ( n63263 , n63261 , n63262 );
xor ( n63264 , n63261 , n63262 );
xor ( n63265 , n62852 , n63162 );
and ( n63266 , n30154 , n63198 );
and ( n63267 , n63265 , n63266 );
xor ( n63268 , n63265 , n63266 );
xor ( n63269 , n62856 , n63160 );
and ( n63270 , n30159 , n63198 );
and ( n63271 , n63269 , n63270 );
xor ( n63272 , n63269 , n63270 );
xor ( n63273 , n62860 , n63158 );
and ( n63274 , n30164 , n63198 );
and ( n63275 , n63273 , n63274 );
xor ( n63276 , n63273 , n63274 );
xor ( n63277 , n62864 , n63156 );
and ( n63278 , n30169 , n63198 );
and ( n63279 , n63277 , n63278 );
xor ( n63280 , n63277 , n63278 );
xor ( n63281 , n62868 , n63154 );
and ( n63282 , n30174 , n63198 );
and ( n63283 , n63281 , n63282 );
xor ( n63284 , n63281 , n63282 );
xor ( n63285 , n62872 , n63152 );
and ( n63286 , n30179 , n63198 );
and ( n63287 , n63285 , n63286 );
xor ( n63288 , n63285 , n63286 );
xor ( n63289 , n62876 , n63150 );
and ( n63290 , n30184 , n63198 );
and ( n63291 , n63289 , n63290 );
xor ( n63292 , n63289 , n63290 );
xor ( n63293 , n62880 , n63148 );
and ( n63294 , n30189 , n63198 );
and ( n63295 , n63293 , n63294 );
xor ( n63296 , n63293 , n63294 );
xor ( n63297 , n62884 , n63146 );
and ( n63298 , n30194 , n63198 );
and ( n63299 , n63297 , n63298 );
xor ( n63300 , n63297 , n63298 );
xor ( n63301 , n62888 , n63144 );
and ( n63302 , n30199 , n63198 );
and ( n63303 , n63301 , n63302 );
xor ( n63304 , n63301 , n63302 );
xor ( n63305 , n62892 , n63142 );
and ( n63306 , n30204 , n63198 );
and ( n63307 , n63305 , n63306 );
xor ( n63308 , n63305 , n63306 );
xor ( n63309 , n62896 , n63140 );
and ( n63310 , n30209 , n63198 );
and ( n63311 , n63309 , n63310 );
xor ( n63312 , n63309 , n63310 );
xor ( n63313 , n62900 , n63138 );
and ( n63314 , n30214 , n63198 );
and ( n63315 , n63313 , n63314 );
xor ( n63316 , n63313 , n63314 );
xor ( n63317 , n62904 , n63136 );
and ( n63318 , n30219 , n63198 );
and ( n63319 , n63317 , n63318 );
xor ( n63320 , n63317 , n63318 );
xor ( n63321 , n62908 , n63134 );
and ( n63322 , n30224 , n63198 );
and ( n63323 , n63321 , n63322 );
xor ( n63324 , n63321 , n63322 );
xor ( n63325 , n62912 , n63132 );
and ( n63326 , n30229 , n63198 );
and ( n63327 , n63325 , n63326 );
xor ( n63328 , n63325 , n63326 );
xor ( n63329 , n62916 , n63130 );
and ( n63330 , n30234 , n63198 );
and ( n63331 , n63329 , n63330 );
xor ( n63332 , n63329 , n63330 );
xor ( n63333 , n62920 , n63128 );
and ( n63334 , n30239 , n63198 );
and ( n63335 , n63333 , n63334 );
xor ( n63336 , n63333 , n63334 );
xor ( n63337 , n62924 , n63126 );
and ( n63338 , n30244 , n63198 );
and ( n63339 , n63337 , n63338 );
xor ( n63340 , n63337 , n63338 );
xor ( n63341 , n62928 , n63124 );
and ( n63342 , n30249 , n63198 );
and ( n63343 , n63341 , n63342 );
xor ( n63344 , n63341 , n63342 );
xor ( n63345 , n62932 , n63122 );
and ( n63346 , n30254 , n63198 );
and ( n63347 , n63345 , n63346 );
xor ( n63348 , n63345 , n63346 );
xor ( n63349 , n62936 , n63120 );
and ( n63350 , n30259 , n63198 );
and ( n63351 , n63349 , n63350 );
xor ( n63352 , n63349 , n63350 );
xor ( n63353 , n62940 , n63118 );
and ( n63354 , n30264 , n63198 );
and ( n63355 , n63353 , n63354 );
xor ( n63356 , n63353 , n63354 );
xor ( n63357 , n62944 , n63116 );
and ( n63358 , n30269 , n63198 );
and ( n63359 , n63357 , n63358 );
xor ( n63360 , n63357 , n63358 );
xor ( n63361 , n62948 , n63114 );
and ( n63362 , n30274 , n63198 );
and ( n63363 , n63361 , n63362 );
xor ( n63364 , n63361 , n63362 );
xor ( n63365 , n62952 , n63112 );
and ( n63366 , n30279 , n63198 );
and ( n63367 , n63365 , n63366 );
xor ( n63368 , n63365 , n63366 );
xor ( n63369 , n62956 , n63110 );
and ( n63370 , n30284 , n63198 );
and ( n63371 , n63369 , n63370 );
xor ( n63372 , n63369 , n63370 );
xor ( n63373 , n62960 , n63108 );
and ( n63374 , n30289 , n63198 );
and ( n63375 , n63373 , n63374 );
xor ( n63376 , n63373 , n63374 );
xor ( n63377 , n62964 , n63106 );
and ( n63378 , n30294 , n63198 );
and ( n63379 , n63377 , n63378 );
xor ( n63380 , n63377 , n63378 );
xor ( n63381 , n62968 , n63104 );
and ( n63382 , n30299 , n63198 );
and ( n63383 , n63381 , n63382 );
xor ( n63384 , n63381 , n63382 );
xor ( n63385 , n62972 , n63102 );
and ( n63386 , n30304 , n63198 );
and ( n63387 , n63385 , n63386 );
xor ( n63388 , n63385 , n63386 );
xor ( n63389 , n62976 , n63100 );
and ( n63390 , n30309 , n63198 );
and ( n63391 , n63389 , n63390 );
xor ( n63392 , n63389 , n63390 );
xor ( n63393 , n62980 , n63098 );
and ( n63394 , n30314 , n63198 );
and ( n63395 , n63393 , n63394 );
xor ( n63396 , n63393 , n63394 );
xor ( n63397 , n62984 , n63096 );
and ( n63398 , n30319 , n63198 );
and ( n63399 , n63397 , n63398 );
xor ( n63400 , n63397 , n63398 );
xor ( n63401 , n62988 , n63094 );
and ( n63402 , n30324 , n63198 );
and ( n63403 , n63401 , n63402 );
xor ( n63404 , n63401 , n63402 );
xor ( n63405 , n62992 , n63092 );
and ( n63406 , n30329 , n63198 );
and ( n63407 , n63405 , n63406 );
xor ( n63408 , n63405 , n63406 );
xor ( n63409 , n62996 , n63090 );
and ( n63410 , n30334 , n63198 );
and ( n63411 , n63409 , n63410 );
xor ( n63412 , n63409 , n63410 );
xor ( n63413 , n63000 , n63088 );
and ( n63414 , n30339 , n63198 );
and ( n63415 , n63413 , n63414 );
xor ( n63416 , n63413 , n63414 );
xor ( n63417 , n63004 , n63086 );
and ( n63418 , n30344 , n63198 );
and ( n63419 , n63417 , n63418 );
xor ( n63420 , n63417 , n63418 );
xor ( n63421 , n63008 , n63084 );
and ( n63422 , n30349 , n63198 );
and ( n63423 , n63421 , n63422 );
xor ( n63424 , n63421 , n63422 );
xor ( n63425 , n63012 , n63082 );
and ( n63426 , n30354 , n63198 );
and ( n63427 , n63425 , n63426 );
xor ( n63428 , n63425 , n63426 );
xor ( n63429 , n63016 , n63080 );
and ( n63430 , n30359 , n63198 );
and ( n63431 , n63429 , n63430 );
xor ( n63432 , n63429 , n63430 );
xor ( n63433 , n63020 , n63078 );
and ( n63434 , n30364 , n63198 );
and ( n63435 , n63433 , n63434 );
xor ( n63436 , n63433 , n63434 );
xor ( n63437 , n63024 , n63076 );
and ( n63438 , n30369 , n63198 );
and ( n63439 , n63437 , n63438 );
xor ( n63440 , n63437 , n63438 );
xor ( n63441 , n63028 , n63074 );
and ( n63442 , n30374 , n63198 );
and ( n63443 , n63441 , n63442 );
xor ( n63444 , n63441 , n63442 );
xor ( n63445 , n63032 , n63072 );
and ( n63446 , n30379 , n63198 );
and ( n63447 , n63445 , n63446 );
xor ( n63448 , n63445 , n63446 );
xor ( n63449 , n63036 , n63070 );
and ( n63450 , n30384 , n63198 );
and ( n63451 , n63449 , n63450 );
xor ( n63452 , n63449 , n63450 );
xor ( n63453 , n63040 , n63068 );
and ( n63454 , n30389 , n63198 );
and ( n63455 , n63453 , n63454 );
xor ( n63456 , n63453 , n63454 );
xor ( n63457 , n63044 , n63066 );
and ( n63458 , n30394 , n63198 );
and ( n63459 , n63457 , n63458 );
xor ( n63460 , n63457 , n63458 );
xor ( n63461 , n63048 , n63064 );
and ( n63462 , n30399 , n63198 );
and ( n63463 , n63461 , n63462 );
xor ( n63464 , n63461 , n63462 );
xor ( n63465 , n63052 , n63062 );
and ( n63466 , n30404 , n63198 );
and ( n63467 , n63465 , n63466 );
xor ( n63468 , n63465 , n63466 );
xor ( n63469 , n63056 , n63060 );
and ( n63470 , n30409 , n63198 );
and ( n63471 , n63469 , n63470 );
buf ( n63472 , n63471 );
and ( n63473 , n63468 , n63472 );
or ( n63474 , n63467 , n63473 );
and ( n63475 , n63464 , n63474 );
or ( n63476 , n63463 , n63475 );
and ( n63477 , n63460 , n63476 );
or ( n63478 , n63459 , n63477 );
and ( n63479 , n63456 , n63478 );
or ( n63480 , n63455 , n63479 );
and ( n63481 , n63452 , n63480 );
or ( n63482 , n63451 , n63481 );
and ( n63483 , n63448 , n63482 );
or ( n63484 , n63447 , n63483 );
and ( n63485 , n63444 , n63484 );
or ( n63486 , n63443 , n63485 );
and ( n63487 , n63440 , n63486 );
or ( n63488 , n63439 , n63487 );
and ( n63489 , n63436 , n63488 );
or ( n63490 , n63435 , n63489 );
and ( n63491 , n63432 , n63490 );
or ( n63492 , n63431 , n63491 );
and ( n63493 , n63428 , n63492 );
or ( n63494 , n63427 , n63493 );
and ( n63495 , n63424 , n63494 );
or ( n63496 , n63423 , n63495 );
and ( n63497 , n63420 , n63496 );
or ( n63498 , n63419 , n63497 );
and ( n63499 , n63416 , n63498 );
or ( n63500 , n63415 , n63499 );
and ( n63501 , n63412 , n63500 );
or ( n63502 , n63411 , n63501 );
and ( n63503 , n63408 , n63502 );
or ( n63504 , n63407 , n63503 );
and ( n63505 , n63404 , n63504 );
or ( n63506 , n63403 , n63505 );
and ( n63507 , n63400 , n63506 );
or ( n63508 , n63399 , n63507 );
and ( n63509 , n63396 , n63508 );
or ( n63510 , n63395 , n63509 );
and ( n63511 , n63392 , n63510 );
or ( n63512 , n63391 , n63511 );
and ( n63513 , n63388 , n63512 );
or ( n63514 , n63387 , n63513 );
and ( n63515 , n63384 , n63514 );
or ( n63516 , n63383 , n63515 );
and ( n63517 , n63380 , n63516 );
or ( n63518 , n63379 , n63517 );
and ( n63519 , n63376 , n63518 );
or ( n63520 , n63375 , n63519 );
and ( n63521 , n63372 , n63520 );
or ( n63522 , n63371 , n63521 );
and ( n63523 , n63368 , n63522 );
or ( n63524 , n63367 , n63523 );
and ( n63525 , n63364 , n63524 );
or ( n63526 , n63363 , n63525 );
and ( n63527 , n63360 , n63526 );
or ( n63528 , n63359 , n63527 );
and ( n63529 , n63356 , n63528 );
or ( n63530 , n63355 , n63529 );
and ( n63531 , n63352 , n63530 );
or ( n63532 , n63351 , n63531 );
and ( n63533 , n63348 , n63532 );
or ( n63534 , n63347 , n63533 );
and ( n63535 , n63344 , n63534 );
or ( n63536 , n63343 , n63535 );
and ( n63537 , n63340 , n63536 );
or ( n63538 , n63339 , n63537 );
and ( n63539 , n63336 , n63538 );
or ( n63540 , n63335 , n63539 );
and ( n63541 , n63332 , n63540 );
or ( n63542 , n63331 , n63541 );
and ( n63543 , n63328 , n63542 );
or ( n63544 , n63327 , n63543 );
and ( n63545 , n63324 , n63544 );
or ( n63546 , n63323 , n63545 );
and ( n63547 , n63320 , n63546 );
or ( n63548 , n63319 , n63547 );
and ( n63549 , n63316 , n63548 );
or ( n63550 , n63315 , n63549 );
and ( n63551 , n63312 , n63550 );
or ( n63552 , n63311 , n63551 );
and ( n63553 , n63308 , n63552 );
or ( n63554 , n63307 , n63553 );
and ( n63555 , n63304 , n63554 );
or ( n63556 , n63303 , n63555 );
and ( n63557 , n63300 , n63556 );
or ( n63558 , n63299 , n63557 );
and ( n63559 , n63296 , n63558 );
or ( n63560 , n63295 , n63559 );
and ( n63561 , n63292 , n63560 );
or ( n63562 , n63291 , n63561 );
and ( n63563 , n63288 , n63562 );
or ( n63564 , n63287 , n63563 );
and ( n63565 , n63284 , n63564 );
or ( n63566 , n63283 , n63565 );
and ( n63567 , n63280 , n63566 );
or ( n63568 , n63279 , n63567 );
and ( n63569 , n63276 , n63568 );
or ( n63570 , n63275 , n63569 );
and ( n63571 , n63272 , n63570 );
or ( n63572 , n63271 , n63571 );
and ( n63573 , n63268 , n63572 );
or ( n63574 , n63267 , n63573 );
and ( n63575 , n63264 , n63574 );
or ( n63576 , n63263 , n63575 );
and ( n63577 , n63260 , n63576 );
or ( n63578 , n63259 , n63577 );
and ( n63579 , n63256 , n63578 );
or ( n63580 , n63255 , n63579 );
and ( n63581 , n63252 , n63580 );
or ( n63582 , n63251 , n63581 );
and ( n63583 , n63248 , n63582 );
or ( n63584 , n63247 , n63583 );
and ( n63585 , n63244 , n63584 );
or ( n63586 , n63243 , n63585 );
and ( n63587 , n63240 , n63586 );
or ( n63588 , n63239 , n63587 );
and ( n63589 , n63236 , n63588 );
or ( n63590 , n63235 , n63589 );
and ( n63591 , n63232 , n63590 );
or ( n63592 , n63231 , n63591 );
and ( n63593 , n63228 , n63592 );
or ( n63594 , n63227 , n63593 );
and ( n63595 , n63224 , n63594 );
or ( n63596 , n63223 , n63595 );
and ( n63597 , n63220 , n63596 );
or ( n63598 , n63219 , n63597 );
and ( n63599 , n63216 , n63598 );
or ( n63600 , n63215 , n63599 );
and ( n63601 , n63212 , n63600 );
or ( n63602 , n63211 , n63601 );
and ( n63603 , n63208 , n63602 );
or ( n63604 , n63207 , n63603 );
and ( n63605 , n63204 , n63604 );
or ( n63606 , n63203 , n63605 );
xor ( n63607 , n63200 , n63606 );
buf ( n63608 , n17988 );
and ( n63609 , n30074 , n63608 );
xor ( n63610 , n63607 , n63609 );
xor ( n63611 , n63204 , n63604 );
and ( n63612 , n30079 , n63608 );
and ( n63613 , n63611 , n63612 );
xor ( n63614 , n63611 , n63612 );
xor ( n63615 , n63208 , n63602 );
and ( n63616 , n30084 , n63608 );
and ( n63617 , n63615 , n63616 );
xor ( n63618 , n63615 , n63616 );
xor ( n63619 , n63212 , n63600 );
and ( n63620 , n30089 , n63608 );
and ( n63621 , n63619 , n63620 );
xor ( n63622 , n63619 , n63620 );
xor ( n63623 , n63216 , n63598 );
and ( n63624 , n30094 , n63608 );
and ( n63625 , n63623 , n63624 );
xor ( n63626 , n63623 , n63624 );
xor ( n63627 , n63220 , n63596 );
and ( n63628 , n30099 , n63608 );
and ( n63629 , n63627 , n63628 );
xor ( n63630 , n63627 , n63628 );
xor ( n63631 , n63224 , n63594 );
and ( n63632 , n30104 , n63608 );
and ( n63633 , n63631 , n63632 );
xor ( n63634 , n63631 , n63632 );
xor ( n63635 , n63228 , n63592 );
and ( n63636 , n30109 , n63608 );
and ( n63637 , n63635 , n63636 );
xor ( n63638 , n63635 , n63636 );
xor ( n63639 , n63232 , n63590 );
and ( n63640 , n30114 , n63608 );
and ( n63641 , n63639 , n63640 );
xor ( n63642 , n63639 , n63640 );
xor ( n63643 , n63236 , n63588 );
and ( n63644 , n30119 , n63608 );
and ( n63645 , n63643 , n63644 );
xor ( n63646 , n63643 , n63644 );
xor ( n63647 , n63240 , n63586 );
and ( n63648 , n30124 , n63608 );
and ( n63649 , n63647 , n63648 );
xor ( n63650 , n63647 , n63648 );
xor ( n63651 , n63244 , n63584 );
and ( n63652 , n30129 , n63608 );
and ( n63653 , n63651 , n63652 );
xor ( n63654 , n63651 , n63652 );
xor ( n63655 , n63248 , n63582 );
and ( n63656 , n30134 , n63608 );
and ( n63657 , n63655 , n63656 );
xor ( n63658 , n63655 , n63656 );
xor ( n63659 , n63252 , n63580 );
and ( n63660 , n30139 , n63608 );
and ( n63661 , n63659 , n63660 );
xor ( n63662 , n63659 , n63660 );
xor ( n63663 , n63256 , n63578 );
and ( n63664 , n30144 , n63608 );
and ( n63665 , n63663 , n63664 );
xor ( n63666 , n63663 , n63664 );
xor ( n63667 , n63260 , n63576 );
and ( n63668 , n30149 , n63608 );
and ( n63669 , n63667 , n63668 );
xor ( n63670 , n63667 , n63668 );
xor ( n63671 , n63264 , n63574 );
and ( n63672 , n30154 , n63608 );
and ( n63673 , n63671 , n63672 );
xor ( n63674 , n63671 , n63672 );
xor ( n63675 , n63268 , n63572 );
and ( n63676 , n30159 , n63608 );
and ( n63677 , n63675 , n63676 );
xor ( n63678 , n63675 , n63676 );
xor ( n63679 , n63272 , n63570 );
and ( n63680 , n30164 , n63608 );
and ( n63681 , n63679 , n63680 );
xor ( n63682 , n63679 , n63680 );
xor ( n63683 , n63276 , n63568 );
and ( n63684 , n30169 , n63608 );
and ( n63685 , n63683 , n63684 );
xor ( n63686 , n63683 , n63684 );
xor ( n63687 , n63280 , n63566 );
and ( n63688 , n30174 , n63608 );
and ( n63689 , n63687 , n63688 );
xor ( n63690 , n63687 , n63688 );
xor ( n63691 , n63284 , n63564 );
and ( n63692 , n30179 , n63608 );
and ( n63693 , n63691 , n63692 );
xor ( n63694 , n63691 , n63692 );
xor ( n63695 , n63288 , n63562 );
and ( n63696 , n30184 , n63608 );
and ( n63697 , n63695 , n63696 );
xor ( n63698 , n63695 , n63696 );
xor ( n63699 , n63292 , n63560 );
and ( n63700 , n30189 , n63608 );
and ( n63701 , n63699 , n63700 );
xor ( n63702 , n63699 , n63700 );
xor ( n63703 , n63296 , n63558 );
and ( n63704 , n30194 , n63608 );
and ( n63705 , n63703 , n63704 );
xor ( n63706 , n63703 , n63704 );
xor ( n63707 , n63300 , n63556 );
and ( n63708 , n30199 , n63608 );
and ( n63709 , n63707 , n63708 );
xor ( n63710 , n63707 , n63708 );
xor ( n63711 , n63304 , n63554 );
and ( n63712 , n30204 , n63608 );
and ( n63713 , n63711 , n63712 );
xor ( n63714 , n63711 , n63712 );
xor ( n63715 , n63308 , n63552 );
and ( n63716 , n30209 , n63608 );
and ( n63717 , n63715 , n63716 );
xor ( n63718 , n63715 , n63716 );
xor ( n63719 , n63312 , n63550 );
and ( n63720 , n30214 , n63608 );
and ( n63721 , n63719 , n63720 );
xor ( n63722 , n63719 , n63720 );
xor ( n63723 , n63316 , n63548 );
and ( n63724 , n30219 , n63608 );
and ( n63725 , n63723 , n63724 );
xor ( n63726 , n63723 , n63724 );
xor ( n63727 , n63320 , n63546 );
and ( n63728 , n30224 , n63608 );
and ( n63729 , n63727 , n63728 );
xor ( n63730 , n63727 , n63728 );
xor ( n63731 , n63324 , n63544 );
and ( n63732 , n30229 , n63608 );
and ( n63733 , n63731 , n63732 );
xor ( n63734 , n63731 , n63732 );
xor ( n63735 , n63328 , n63542 );
and ( n63736 , n30234 , n63608 );
and ( n63737 , n63735 , n63736 );
xor ( n63738 , n63735 , n63736 );
xor ( n63739 , n63332 , n63540 );
and ( n63740 , n30239 , n63608 );
and ( n63741 , n63739 , n63740 );
xor ( n63742 , n63739 , n63740 );
xor ( n63743 , n63336 , n63538 );
and ( n63744 , n30244 , n63608 );
and ( n63745 , n63743 , n63744 );
xor ( n63746 , n63743 , n63744 );
xor ( n63747 , n63340 , n63536 );
and ( n63748 , n30249 , n63608 );
and ( n63749 , n63747 , n63748 );
xor ( n63750 , n63747 , n63748 );
xor ( n63751 , n63344 , n63534 );
and ( n63752 , n30254 , n63608 );
and ( n63753 , n63751 , n63752 );
xor ( n63754 , n63751 , n63752 );
xor ( n63755 , n63348 , n63532 );
and ( n63756 , n30259 , n63608 );
and ( n63757 , n63755 , n63756 );
xor ( n63758 , n63755 , n63756 );
xor ( n63759 , n63352 , n63530 );
and ( n63760 , n30264 , n63608 );
and ( n63761 , n63759 , n63760 );
xor ( n63762 , n63759 , n63760 );
xor ( n63763 , n63356 , n63528 );
and ( n63764 , n30269 , n63608 );
and ( n63765 , n63763 , n63764 );
xor ( n63766 , n63763 , n63764 );
xor ( n63767 , n63360 , n63526 );
and ( n63768 , n30274 , n63608 );
and ( n63769 , n63767 , n63768 );
xor ( n63770 , n63767 , n63768 );
xor ( n63771 , n63364 , n63524 );
and ( n63772 , n30279 , n63608 );
and ( n63773 , n63771 , n63772 );
xor ( n63774 , n63771 , n63772 );
xor ( n63775 , n63368 , n63522 );
and ( n63776 , n30284 , n63608 );
and ( n63777 , n63775 , n63776 );
xor ( n63778 , n63775 , n63776 );
xor ( n63779 , n63372 , n63520 );
and ( n63780 , n30289 , n63608 );
and ( n63781 , n63779 , n63780 );
xor ( n63782 , n63779 , n63780 );
xor ( n63783 , n63376 , n63518 );
and ( n63784 , n30294 , n63608 );
and ( n63785 , n63783 , n63784 );
xor ( n63786 , n63783 , n63784 );
xor ( n63787 , n63380 , n63516 );
and ( n63788 , n30299 , n63608 );
and ( n63789 , n63787 , n63788 );
xor ( n63790 , n63787 , n63788 );
xor ( n63791 , n63384 , n63514 );
and ( n63792 , n30304 , n63608 );
and ( n63793 , n63791 , n63792 );
xor ( n63794 , n63791 , n63792 );
xor ( n63795 , n63388 , n63512 );
and ( n63796 , n30309 , n63608 );
and ( n63797 , n63795 , n63796 );
xor ( n63798 , n63795 , n63796 );
xor ( n63799 , n63392 , n63510 );
and ( n63800 , n30314 , n63608 );
and ( n63801 , n63799 , n63800 );
xor ( n63802 , n63799 , n63800 );
xor ( n63803 , n63396 , n63508 );
and ( n63804 , n30319 , n63608 );
and ( n63805 , n63803 , n63804 );
xor ( n63806 , n63803 , n63804 );
xor ( n63807 , n63400 , n63506 );
and ( n63808 , n30324 , n63608 );
and ( n63809 , n63807 , n63808 );
xor ( n63810 , n63807 , n63808 );
xor ( n63811 , n63404 , n63504 );
and ( n63812 , n30329 , n63608 );
and ( n63813 , n63811 , n63812 );
xor ( n63814 , n63811 , n63812 );
xor ( n63815 , n63408 , n63502 );
and ( n63816 , n30334 , n63608 );
and ( n63817 , n63815 , n63816 );
xor ( n63818 , n63815 , n63816 );
xor ( n63819 , n63412 , n63500 );
and ( n63820 , n30339 , n63608 );
and ( n63821 , n63819 , n63820 );
xor ( n63822 , n63819 , n63820 );
xor ( n63823 , n63416 , n63498 );
and ( n63824 , n30344 , n63608 );
and ( n63825 , n63823 , n63824 );
xor ( n63826 , n63823 , n63824 );
xor ( n63827 , n63420 , n63496 );
and ( n63828 , n30349 , n63608 );
and ( n63829 , n63827 , n63828 );
xor ( n63830 , n63827 , n63828 );
xor ( n63831 , n63424 , n63494 );
and ( n63832 , n30354 , n63608 );
and ( n63833 , n63831 , n63832 );
xor ( n63834 , n63831 , n63832 );
xor ( n63835 , n63428 , n63492 );
and ( n63836 , n30359 , n63608 );
and ( n63837 , n63835 , n63836 );
xor ( n63838 , n63835 , n63836 );
xor ( n63839 , n63432 , n63490 );
and ( n63840 , n30364 , n63608 );
and ( n63841 , n63839 , n63840 );
xor ( n63842 , n63839 , n63840 );
xor ( n63843 , n63436 , n63488 );
and ( n63844 , n30369 , n63608 );
and ( n63845 , n63843 , n63844 );
xor ( n63846 , n63843 , n63844 );
xor ( n63847 , n63440 , n63486 );
and ( n63848 , n30374 , n63608 );
and ( n63849 , n63847 , n63848 );
xor ( n63850 , n63847 , n63848 );
xor ( n63851 , n63444 , n63484 );
and ( n63852 , n30379 , n63608 );
and ( n63853 , n63851 , n63852 );
xor ( n63854 , n63851 , n63852 );
xor ( n63855 , n63448 , n63482 );
and ( n63856 , n30384 , n63608 );
and ( n63857 , n63855 , n63856 );
xor ( n63858 , n63855 , n63856 );
xor ( n63859 , n63452 , n63480 );
and ( n63860 , n30389 , n63608 );
and ( n63861 , n63859 , n63860 );
xor ( n63862 , n63859 , n63860 );
xor ( n63863 , n63456 , n63478 );
and ( n63864 , n30394 , n63608 );
and ( n63865 , n63863 , n63864 );
xor ( n63866 , n63863 , n63864 );
xor ( n63867 , n63460 , n63476 );
and ( n63868 , n30399 , n63608 );
and ( n63869 , n63867 , n63868 );
xor ( n63870 , n63867 , n63868 );
xor ( n63871 , n63464 , n63474 );
and ( n63872 , n30404 , n63608 );
and ( n63873 , n63871 , n63872 );
xor ( n63874 , n63871 , n63872 );
xor ( n63875 , n63468 , n63472 );
and ( n63876 , n30409 , n63608 );
and ( n63877 , n63875 , n63876 );
buf ( n63878 , n63877 );
and ( n63879 , n63874 , n63878 );
or ( n63880 , n63873 , n63879 );
and ( n63881 , n63870 , n63880 );
or ( n63882 , n63869 , n63881 );
and ( n63883 , n63866 , n63882 );
or ( n63884 , n63865 , n63883 );
and ( n63885 , n63862 , n63884 );
or ( n63886 , n63861 , n63885 );
and ( n63887 , n63858 , n63886 );
or ( n63888 , n63857 , n63887 );
and ( n63889 , n63854 , n63888 );
or ( n63890 , n63853 , n63889 );
and ( n63891 , n63850 , n63890 );
or ( n63892 , n63849 , n63891 );
and ( n63893 , n63846 , n63892 );
or ( n63894 , n63845 , n63893 );
and ( n63895 , n63842 , n63894 );
or ( n63896 , n63841 , n63895 );
and ( n63897 , n63838 , n63896 );
or ( n63898 , n63837 , n63897 );
and ( n63899 , n63834 , n63898 );
or ( n63900 , n63833 , n63899 );
and ( n63901 , n63830 , n63900 );
or ( n63902 , n63829 , n63901 );
and ( n63903 , n63826 , n63902 );
or ( n63904 , n63825 , n63903 );
and ( n63905 , n63822 , n63904 );
or ( n63906 , n63821 , n63905 );
and ( n63907 , n63818 , n63906 );
or ( n63908 , n63817 , n63907 );
and ( n63909 , n63814 , n63908 );
or ( n63910 , n63813 , n63909 );
and ( n63911 , n63810 , n63910 );
or ( n63912 , n63809 , n63911 );
and ( n63913 , n63806 , n63912 );
or ( n63914 , n63805 , n63913 );
and ( n63915 , n63802 , n63914 );
or ( n63916 , n63801 , n63915 );
and ( n63917 , n63798 , n63916 );
or ( n63918 , n63797 , n63917 );
and ( n63919 , n63794 , n63918 );
or ( n63920 , n63793 , n63919 );
and ( n63921 , n63790 , n63920 );
or ( n63922 , n63789 , n63921 );
and ( n63923 , n63786 , n63922 );
or ( n63924 , n63785 , n63923 );
and ( n63925 , n63782 , n63924 );
or ( n63926 , n63781 , n63925 );
and ( n63927 , n63778 , n63926 );
or ( n63928 , n63777 , n63927 );
and ( n63929 , n63774 , n63928 );
or ( n63930 , n63773 , n63929 );
and ( n63931 , n63770 , n63930 );
or ( n63932 , n63769 , n63931 );
and ( n63933 , n63766 , n63932 );
or ( n63934 , n63765 , n63933 );
and ( n63935 , n63762 , n63934 );
or ( n63936 , n63761 , n63935 );
and ( n63937 , n63758 , n63936 );
or ( n63938 , n63757 , n63937 );
and ( n63939 , n63754 , n63938 );
or ( n63940 , n63753 , n63939 );
and ( n63941 , n63750 , n63940 );
or ( n63942 , n63749 , n63941 );
and ( n63943 , n63746 , n63942 );
or ( n63944 , n63745 , n63943 );
and ( n63945 , n63742 , n63944 );
or ( n63946 , n63741 , n63945 );
and ( n63947 , n63738 , n63946 );
or ( n63948 , n63737 , n63947 );
and ( n63949 , n63734 , n63948 );
or ( n63950 , n63733 , n63949 );
and ( n63951 , n63730 , n63950 );
or ( n63952 , n63729 , n63951 );
and ( n63953 , n63726 , n63952 );
or ( n63954 , n63725 , n63953 );
and ( n63955 , n63722 , n63954 );
or ( n63956 , n63721 , n63955 );
and ( n63957 , n63718 , n63956 );
or ( n63958 , n63717 , n63957 );
and ( n63959 , n63714 , n63958 );
or ( n63960 , n63713 , n63959 );
and ( n63961 , n63710 , n63960 );
or ( n63962 , n63709 , n63961 );
and ( n63963 , n63706 , n63962 );
or ( n63964 , n63705 , n63963 );
and ( n63965 , n63702 , n63964 );
or ( n63966 , n63701 , n63965 );
and ( n63967 , n63698 , n63966 );
or ( n63968 , n63697 , n63967 );
and ( n63969 , n63694 , n63968 );
or ( n63970 , n63693 , n63969 );
and ( n63971 , n63690 , n63970 );
or ( n63972 , n63689 , n63971 );
and ( n63973 , n63686 , n63972 );
or ( n63974 , n63685 , n63973 );
and ( n63975 , n63682 , n63974 );
or ( n63976 , n63681 , n63975 );
and ( n63977 , n63678 , n63976 );
or ( n63978 , n63677 , n63977 );
and ( n63979 , n63674 , n63978 );
or ( n63980 , n63673 , n63979 );
and ( n63981 , n63670 , n63980 );
or ( n63982 , n63669 , n63981 );
and ( n63983 , n63666 , n63982 );
or ( n63984 , n63665 , n63983 );
and ( n63985 , n63662 , n63984 );
or ( n63986 , n63661 , n63985 );
and ( n63987 , n63658 , n63986 );
or ( n63988 , n63657 , n63987 );
and ( n63989 , n63654 , n63988 );
or ( n63990 , n63653 , n63989 );
and ( n63991 , n63650 , n63990 );
or ( n63992 , n63649 , n63991 );
and ( n63993 , n63646 , n63992 );
or ( n63994 , n63645 , n63993 );
and ( n63995 , n63642 , n63994 );
or ( n63996 , n63641 , n63995 );
and ( n63997 , n63638 , n63996 );
or ( n63998 , n63637 , n63997 );
and ( n63999 , n63634 , n63998 );
or ( n64000 , n63633 , n63999 );
and ( n64001 , n63630 , n64000 );
or ( n64002 , n63629 , n64001 );
and ( n64003 , n63626 , n64002 );
or ( n64004 , n63625 , n64003 );
and ( n64005 , n63622 , n64004 );
or ( n64006 , n63621 , n64005 );
and ( n64007 , n63618 , n64006 );
or ( n64008 , n63617 , n64007 );
and ( n64009 , n63614 , n64008 );
or ( n64010 , n63613 , n64009 );
xor ( n64011 , n63610 , n64010 );
buf ( n64012 , n17986 );
and ( n64013 , n30079 , n64012 );
xor ( n64014 , n64011 , n64013 );
xor ( n64015 , n63614 , n64008 );
and ( n64016 , n30084 , n64012 );
and ( n64017 , n64015 , n64016 );
xor ( n64018 , n64015 , n64016 );
xor ( n64019 , n63618 , n64006 );
and ( n64020 , n30089 , n64012 );
and ( n64021 , n64019 , n64020 );
xor ( n64022 , n64019 , n64020 );
xor ( n64023 , n63622 , n64004 );
and ( n64024 , n30094 , n64012 );
and ( n64025 , n64023 , n64024 );
xor ( n64026 , n64023 , n64024 );
xor ( n64027 , n63626 , n64002 );
and ( n64028 , n30099 , n64012 );
and ( n64029 , n64027 , n64028 );
xor ( n64030 , n64027 , n64028 );
xor ( n64031 , n63630 , n64000 );
and ( n64032 , n30104 , n64012 );
and ( n64033 , n64031 , n64032 );
xor ( n64034 , n64031 , n64032 );
xor ( n64035 , n63634 , n63998 );
and ( n64036 , n30109 , n64012 );
and ( n64037 , n64035 , n64036 );
xor ( n64038 , n64035 , n64036 );
xor ( n64039 , n63638 , n63996 );
and ( n64040 , n30114 , n64012 );
and ( n64041 , n64039 , n64040 );
xor ( n64042 , n64039 , n64040 );
xor ( n64043 , n63642 , n63994 );
and ( n64044 , n30119 , n64012 );
and ( n64045 , n64043 , n64044 );
xor ( n64046 , n64043 , n64044 );
xor ( n64047 , n63646 , n63992 );
and ( n64048 , n30124 , n64012 );
and ( n64049 , n64047 , n64048 );
xor ( n64050 , n64047 , n64048 );
xor ( n64051 , n63650 , n63990 );
and ( n64052 , n30129 , n64012 );
and ( n64053 , n64051 , n64052 );
xor ( n64054 , n64051 , n64052 );
xor ( n64055 , n63654 , n63988 );
and ( n64056 , n30134 , n64012 );
and ( n64057 , n64055 , n64056 );
xor ( n64058 , n64055 , n64056 );
xor ( n64059 , n63658 , n63986 );
and ( n64060 , n30139 , n64012 );
and ( n64061 , n64059 , n64060 );
xor ( n64062 , n64059 , n64060 );
xor ( n64063 , n63662 , n63984 );
and ( n64064 , n30144 , n64012 );
and ( n64065 , n64063 , n64064 );
xor ( n64066 , n64063 , n64064 );
xor ( n64067 , n63666 , n63982 );
and ( n64068 , n30149 , n64012 );
and ( n64069 , n64067 , n64068 );
xor ( n64070 , n64067 , n64068 );
xor ( n64071 , n63670 , n63980 );
and ( n64072 , n30154 , n64012 );
and ( n64073 , n64071 , n64072 );
xor ( n64074 , n64071 , n64072 );
xor ( n64075 , n63674 , n63978 );
and ( n64076 , n30159 , n64012 );
and ( n64077 , n64075 , n64076 );
xor ( n64078 , n64075 , n64076 );
xor ( n64079 , n63678 , n63976 );
and ( n64080 , n30164 , n64012 );
and ( n64081 , n64079 , n64080 );
xor ( n64082 , n64079 , n64080 );
xor ( n64083 , n63682 , n63974 );
and ( n64084 , n30169 , n64012 );
and ( n64085 , n64083 , n64084 );
xor ( n64086 , n64083 , n64084 );
xor ( n64087 , n63686 , n63972 );
and ( n64088 , n30174 , n64012 );
and ( n64089 , n64087 , n64088 );
xor ( n64090 , n64087 , n64088 );
xor ( n64091 , n63690 , n63970 );
and ( n64092 , n30179 , n64012 );
and ( n64093 , n64091 , n64092 );
xor ( n64094 , n64091 , n64092 );
xor ( n64095 , n63694 , n63968 );
and ( n64096 , n30184 , n64012 );
and ( n64097 , n64095 , n64096 );
xor ( n64098 , n64095 , n64096 );
xor ( n64099 , n63698 , n63966 );
and ( n64100 , n30189 , n64012 );
and ( n64101 , n64099 , n64100 );
xor ( n64102 , n64099 , n64100 );
xor ( n64103 , n63702 , n63964 );
and ( n64104 , n30194 , n64012 );
and ( n64105 , n64103 , n64104 );
xor ( n64106 , n64103 , n64104 );
xor ( n64107 , n63706 , n63962 );
and ( n64108 , n30199 , n64012 );
and ( n64109 , n64107 , n64108 );
xor ( n64110 , n64107 , n64108 );
xor ( n64111 , n63710 , n63960 );
and ( n64112 , n30204 , n64012 );
and ( n64113 , n64111 , n64112 );
xor ( n64114 , n64111 , n64112 );
xor ( n64115 , n63714 , n63958 );
and ( n64116 , n30209 , n64012 );
and ( n64117 , n64115 , n64116 );
xor ( n64118 , n64115 , n64116 );
xor ( n64119 , n63718 , n63956 );
and ( n64120 , n30214 , n64012 );
and ( n64121 , n64119 , n64120 );
xor ( n64122 , n64119 , n64120 );
xor ( n64123 , n63722 , n63954 );
and ( n64124 , n30219 , n64012 );
and ( n64125 , n64123 , n64124 );
xor ( n64126 , n64123 , n64124 );
xor ( n64127 , n63726 , n63952 );
and ( n64128 , n30224 , n64012 );
and ( n64129 , n64127 , n64128 );
xor ( n64130 , n64127 , n64128 );
xor ( n64131 , n63730 , n63950 );
and ( n64132 , n30229 , n64012 );
and ( n64133 , n64131 , n64132 );
xor ( n64134 , n64131 , n64132 );
xor ( n64135 , n63734 , n63948 );
and ( n64136 , n30234 , n64012 );
and ( n64137 , n64135 , n64136 );
xor ( n64138 , n64135 , n64136 );
xor ( n64139 , n63738 , n63946 );
and ( n64140 , n30239 , n64012 );
and ( n64141 , n64139 , n64140 );
xor ( n64142 , n64139 , n64140 );
xor ( n64143 , n63742 , n63944 );
and ( n64144 , n30244 , n64012 );
and ( n64145 , n64143 , n64144 );
xor ( n64146 , n64143 , n64144 );
xor ( n64147 , n63746 , n63942 );
and ( n64148 , n30249 , n64012 );
and ( n64149 , n64147 , n64148 );
xor ( n64150 , n64147 , n64148 );
xor ( n64151 , n63750 , n63940 );
and ( n64152 , n30254 , n64012 );
and ( n64153 , n64151 , n64152 );
xor ( n64154 , n64151 , n64152 );
xor ( n64155 , n63754 , n63938 );
and ( n64156 , n30259 , n64012 );
and ( n64157 , n64155 , n64156 );
xor ( n64158 , n64155 , n64156 );
xor ( n64159 , n63758 , n63936 );
and ( n64160 , n30264 , n64012 );
and ( n64161 , n64159 , n64160 );
xor ( n64162 , n64159 , n64160 );
xor ( n64163 , n63762 , n63934 );
and ( n64164 , n30269 , n64012 );
and ( n64165 , n64163 , n64164 );
xor ( n64166 , n64163 , n64164 );
xor ( n64167 , n63766 , n63932 );
and ( n64168 , n30274 , n64012 );
and ( n64169 , n64167 , n64168 );
xor ( n64170 , n64167 , n64168 );
xor ( n64171 , n63770 , n63930 );
and ( n64172 , n30279 , n64012 );
and ( n64173 , n64171 , n64172 );
xor ( n64174 , n64171 , n64172 );
xor ( n64175 , n63774 , n63928 );
and ( n64176 , n30284 , n64012 );
and ( n64177 , n64175 , n64176 );
xor ( n64178 , n64175 , n64176 );
xor ( n64179 , n63778 , n63926 );
and ( n64180 , n30289 , n64012 );
and ( n64181 , n64179 , n64180 );
xor ( n64182 , n64179 , n64180 );
xor ( n64183 , n63782 , n63924 );
and ( n64184 , n30294 , n64012 );
and ( n64185 , n64183 , n64184 );
xor ( n64186 , n64183 , n64184 );
xor ( n64187 , n63786 , n63922 );
and ( n64188 , n30299 , n64012 );
and ( n64189 , n64187 , n64188 );
xor ( n64190 , n64187 , n64188 );
xor ( n64191 , n63790 , n63920 );
and ( n64192 , n30304 , n64012 );
and ( n64193 , n64191 , n64192 );
xor ( n64194 , n64191 , n64192 );
xor ( n64195 , n63794 , n63918 );
and ( n64196 , n30309 , n64012 );
and ( n64197 , n64195 , n64196 );
xor ( n64198 , n64195 , n64196 );
xor ( n64199 , n63798 , n63916 );
and ( n64200 , n30314 , n64012 );
and ( n64201 , n64199 , n64200 );
xor ( n64202 , n64199 , n64200 );
xor ( n64203 , n63802 , n63914 );
and ( n64204 , n30319 , n64012 );
and ( n64205 , n64203 , n64204 );
xor ( n64206 , n64203 , n64204 );
xor ( n64207 , n63806 , n63912 );
and ( n64208 , n30324 , n64012 );
and ( n64209 , n64207 , n64208 );
xor ( n64210 , n64207 , n64208 );
xor ( n64211 , n63810 , n63910 );
and ( n64212 , n30329 , n64012 );
and ( n64213 , n64211 , n64212 );
xor ( n64214 , n64211 , n64212 );
xor ( n64215 , n63814 , n63908 );
and ( n64216 , n30334 , n64012 );
and ( n64217 , n64215 , n64216 );
xor ( n64218 , n64215 , n64216 );
xor ( n64219 , n63818 , n63906 );
and ( n64220 , n30339 , n64012 );
and ( n64221 , n64219 , n64220 );
xor ( n64222 , n64219 , n64220 );
xor ( n64223 , n63822 , n63904 );
and ( n64224 , n30344 , n64012 );
and ( n64225 , n64223 , n64224 );
xor ( n64226 , n64223 , n64224 );
xor ( n64227 , n63826 , n63902 );
and ( n64228 , n30349 , n64012 );
and ( n64229 , n64227 , n64228 );
xor ( n64230 , n64227 , n64228 );
xor ( n64231 , n63830 , n63900 );
and ( n64232 , n30354 , n64012 );
and ( n64233 , n64231 , n64232 );
xor ( n64234 , n64231 , n64232 );
xor ( n64235 , n63834 , n63898 );
and ( n64236 , n30359 , n64012 );
and ( n64237 , n64235 , n64236 );
xor ( n64238 , n64235 , n64236 );
xor ( n64239 , n63838 , n63896 );
and ( n64240 , n30364 , n64012 );
and ( n64241 , n64239 , n64240 );
xor ( n64242 , n64239 , n64240 );
xor ( n64243 , n63842 , n63894 );
and ( n64244 , n30369 , n64012 );
and ( n64245 , n64243 , n64244 );
xor ( n64246 , n64243 , n64244 );
xor ( n64247 , n63846 , n63892 );
and ( n64248 , n30374 , n64012 );
and ( n64249 , n64247 , n64248 );
xor ( n64250 , n64247 , n64248 );
xor ( n64251 , n63850 , n63890 );
and ( n64252 , n30379 , n64012 );
and ( n64253 , n64251 , n64252 );
xor ( n64254 , n64251 , n64252 );
xor ( n64255 , n63854 , n63888 );
and ( n64256 , n30384 , n64012 );
and ( n64257 , n64255 , n64256 );
xor ( n64258 , n64255 , n64256 );
xor ( n64259 , n63858 , n63886 );
and ( n64260 , n30389 , n64012 );
and ( n64261 , n64259 , n64260 );
xor ( n64262 , n64259 , n64260 );
xor ( n64263 , n63862 , n63884 );
and ( n64264 , n30394 , n64012 );
and ( n64265 , n64263 , n64264 );
xor ( n64266 , n64263 , n64264 );
xor ( n64267 , n63866 , n63882 );
and ( n64268 , n30399 , n64012 );
and ( n64269 , n64267 , n64268 );
xor ( n64270 , n64267 , n64268 );
xor ( n64271 , n63870 , n63880 );
and ( n64272 , n30404 , n64012 );
and ( n64273 , n64271 , n64272 );
xor ( n64274 , n64271 , n64272 );
xor ( n64275 , n63874 , n63878 );
and ( n64276 , n30409 , n64012 );
and ( n64277 , n64275 , n64276 );
buf ( n64278 , n64277 );
and ( n64279 , n64274 , n64278 );
or ( n64280 , n64273 , n64279 );
and ( n64281 , n64270 , n64280 );
or ( n64282 , n64269 , n64281 );
and ( n64283 , n64266 , n64282 );
or ( n64284 , n64265 , n64283 );
and ( n64285 , n64262 , n64284 );
or ( n64286 , n64261 , n64285 );
and ( n64287 , n64258 , n64286 );
or ( n64288 , n64257 , n64287 );
and ( n64289 , n64254 , n64288 );
or ( n64290 , n64253 , n64289 );
and ( n64291 , n64250 , n64290 );
or ( n64292 , n64249 , n64291 );
and ( n64293 , n64246 , n64292 );
or ( n64294 , n64245 , n64293 );
and ( n64295 , n64242 , n64294 );
or ( n64296 , n64241 , n64295 );
and ( n64297 , n64238 , n64296 );
or ( n64298 , n64237 , n64297 );
and ( n64299 , n64234 , n64298 );
or ( n64300 , n64233 , n64299 );
and ( n64301 , n64230 , n64300 );
or ( n64302 , n64229 , n64301 );
and ( n64303 , n64226 , n64302 );
or ( n64304 , n64225 , n64303 );
and ( n64305 , n64222 , n64304 );
or ( n64306 , n64221 , n64305 );
and ( n64307 , n64218 , n64306 );
or ( n64308 , n64217 , n64307 );
and ( n64309 , n64214 , n64308 );
or ( n64310 , n64213 , n64309 );
and ( n64311 , n64210 , n64310 );
or ( n64312 , n64209 , n64311 );
and ( n64313 , n64206 , n64312 );
or ( n64314 , n64205 , n64313 );
and ( n64315 , n64202 , n64314 );
or ( n64316 , n64201 , n64315 );
and ( n64317 , n64198 , n64316 );
or ( n64318 , n64197 , n64317 );
and ( n64319 , n64194 , n64318 );
or ( n64320 , n64193 , n64319 );
and ( n64321 , n64190 , n64320 );
or ( n64322 , n64189 , n64321 );
and ( n64323 , n64186 , n64322 );
or ( n64324 , n64185 , n64323 );
and ( n64325 , n64182 , n64324 );
or ( n64326 , n64181 , n64325 );
and ( n64327 , n64178 , n64326 );
or ( n64328 , n64177 , n64327 );
and ( n64329 , n64174 , n64328 );
or ( n64330 , n64173 , n64329 );
and ( n64331 , n64170 , n64330 );
or ( n64332 , n64169 , n64331 );
and ( n64333 , n64166 , n64332 );
or ( n64334 , n64165 , n64333 );
and ( n64335 , n64162 , n64334 );
or ( n64336 , n64161 , n64335 );
and ( n64337 , n64158 , n64336 );
or ( n64338 , n64157 , n64337 );
and ( n64339 , n64154 , n64338 );
or ( n64340 , n64153 , n64339 );
and ( n64341 , n64150 , n64340 );
or ( n64342 , n64149 , n64341 );
and ( n64343 , n64146 , n64342 );
or ( n64344 , n64145 , n64343 );
and ( n64345 , n64142 , n64344 );
or ( n64346 , n64141 , n64345 );
and ( n64347 , n64138 , n64346 );
or ( n64348 , n64137 , n64347 );
and ( n64349 , n64134 , n64348 );
or ( n64350 , n64133 , n64349 );
and ( n64351 , n64130 , n64350 );
or ( n64352 , n64129 , n64351 );
and ( n64353 , n64126 , n64352 );
or ( n64354 , n64125 , n64353 );
and ( n64355 , n64122 , n64354 );
or ( n64356 , n64121 , n64355 );
and ( n64357 , n64118 , n64356 );
or ( n64358 , n64117 , n64357 );
and ( n64359 , n64114 , n64358 );
or ( n64360 , n64113 , n64359 );
and ( n64361 , n64110 , n64360 );
or ( n64362 , n64109 , n64361 );
and ( n64363 , n64106 , n64362 );
or ( n64364 , n64105 , n64363 );
and ( n64365 , n64102 , n64364 );
or ( n64366 , n64101 , n64365 );
and ( n64367 , n64098 , n64366 );
or ( n64368 , n64097 , n64367 );
and ( n64369 , n64094 , n64368 );
or ( n64370 , n64093 , n64369 );
and ( n64371 , n64090 , n64370 );
or ( n64372 , n64089 , n64371 );
and ( n64373 , n64086 , n64372 );
or ( n64374 , n64085 , n64373 );
and ( n64375 , n64082 , n64374 );
or ( n64376 , n64081 , n64375 );
and ( n64377 , n64078 , n64376 );
or ( n64378 , n64077 , n64377 );
and ( n64379 , n64074 , n64378 );
or ( n64380 , n64073 , n64379 );
and ( n64381 , n64070 , n64380 );
or ( n64382 , n64069 , n64381 );
and ( n64383 , n64066 , n64382 );
or ( n64384 , n64065 , n64383 );
and ( n64385 , n64062 , n64384 );
or ( n64386 , n64061 , n64385 );
and ( n64387 , n64058 , n64386 );
or ( n64388 , n64057 , n64387 );
and ( n64389 , n64054 , n64388 );
or ( n64390 , n64053 , n64389 );
and ( n64391 , n64050 , n64390 );
or ( n64392 , n64049 , n64391 );
and ( n64393 , n64046 , n64392 );
or ( n64394 , n64045 , n64393 );
and ( n64395 , n64042 , n64394 );
or ( n64396 , n64041 , n64395 );
and ( n64397 , n64038 , n64396 );
or ( n64398 , n64037 , n64397 );
and ( n64399 , n64034 , n64398 );
or ( n64400 , n64033 , n64399 );
and ( n64401 , n64030 , n64400 );
or ( n64402 , n64029 , n64401 );
and ( n64403 , n64026 , n64402 );
or ( n64404 , n64025 , n64403 );
and ( n64405 , n64022 , n64404 );
or ( n64406 , n64021 , n64405 );
and ( n64407 , n64018 , n64406 );
or ( n64408 , n64017 , n64407 );
xor ( n64409 , n64014 , n64408 );
buf ( n64410 , n17984 );
and ( n64411 , n30084 , n64410 );
xor ( n64412 , n64409 , n64411 );
xor ( n64413 , n64018 , n64406 );
and ( n64414 , n30089 , n64410 );
and ( n64415 , n64413 , n64414 );
xor ( n64416 , n64413 , n64414 );
xor ( n64417 , n64022 , n64404 );
and ( n64418 , n30094 , n64410 );
and ( n64419 , n64417 , n64418 );
xor ( n64420 , n64417 , n64418 );
xor ( n64421 , n64026 , n64402 );
and ( n64422 , n30099 , n64410 );
and ( n64423 , n64421 , n64422 );
xor ( n64424 , n64421 , n64422 );
xor ( n64425 , n64030 , n64400 );
and ( n64426 , n30104 , n64410 );
and ( n64427 , n64425 , n64426 );
xor ( n64428 , n64425 , n64426 );
xor ( n64429 , n64034 , n64398 );
and ( n64430 , n30109 , n64410 );
and ( n64431 , n64429 , n64430 );
xor ( n64432 , n64429 , n64430 );
xor ( n64433 , n64038 , n64396 );
and ( n64434 , n30114 , n64410 );
and ( n64435 , n64433 , n64434 );
xor ( n64436 , n64433 , n64434 );
xor ( n64437 , n64042 , n64394 );
and ( n64438 , n30119 , n64410 );
and ( n64439 , n64437 , n64438 );
xor ( n64440 , n64437 , n64438 );
xor ( n64441 , n64046 , n64392 );
and ( n64442 , n30124 , n64410 );
and ( n64443 , n64441 , n64442 );
xor ( n64444 , n64441 , n64442 );
xor ( n64445 , n64050 , n64390 );
and ( n64446 , n30129 , n64410 );
and ( n64447 , n64445 , n64446 );
xor ( n64448 , n64445 , n64446 );
xor ( n64449 , n64054 , n64388 );
and ( n64450 , n30134 , n64410 );
and ( n64451 , n64449 , n64450 );
xor ( n64452 , n64449 , n64450 );
xor ( n64453 , n64058 , n64386 );
and ( n64454 , n30139 , n64410 );
and ( n64455 , n64453 , n64454 );
xor ( n64456 , n64453 , n64454 );
xor ( n64457 , n64062 , n64384 );
and ( n64458 , n30144 , n64410 );
and ( n64459 , n64457 , n64458 );
xor ( n64460 , n64457 , n64458 );
xor ( n64461 , n64066 , n64382 );
and ( n64462 , n30149 , n64410 );
and ( n64463 , n64461 , n64462 );
xor ( n64464 , n64461 , n64462 );
xor ( n64465 , n64070 , n64380 );
and ( n64466 , n30154 , n64410 );
and ( n64467 , n64465 , n64466 );
xor ( n64468 , n64465 , n64466 );
xor ( n64469 , n64074 , n64378 );
and ( n64470 , n30159 , n64410 );
and ( n64471 , n64469 , n64470 );
xor ( n64472 , n64469 , n64470 );
xor ( n64473 , n64078 , n64376 );
and ( n64474 , n30164 , n64410 );
and ( n64475 , n64473 , n64474 );
xor ( n64476 , n64473 , n64474 );
xor ( n64477 , n64082 , n64374 );
and ( n64478 , n30169 , n64410 );
and ( n64479 , n64477 , n64478 );
xor ( n64480 , n64477 , n64478 );
xor ( n64481 , n64086 , n64372 );
and ( n64482 , n30174 , n64410 );
and ( n64483 , n64481 , n64482 );
xor ( n64484 , n64481 , n64482 );
xor ( n64485 , n64090 , n64370 );
and ( n64486 , n30179 , n64410 );
and ( n64487 , n64485 , n64486 );
xor ( n64488 , n64485 , n64486 );
xor ( n64489 , n64094 , n64368 );
and ( n64490 , n30184 , n64410 );
and ( n64491 , n64489 , n64490 );
xor ( n64492 , n64489 , n64490 );
xor ( n64493 , n64098 , n64366 );
and ( n64494 , n30189 , n64410 );
and ( n64495 , n64493 , n64494 );
xor ( n64496 , n64493 , n64494 );
xor ( n64497 , n64102 , n64364 );
and ( n64498 , n30194 , n64410 );
and ( n64499 , n64497 , n64498 );
xor ( n64500 , n64497 , n64498 );
xor ( n64501 , n64106 , n64362 );
and ( n64502 , n30199 , n64410 );
and ( n64503 , n64501 , n64502 );
xor ( n64504 , n64501 , n64502 );
xor ( n64505 , n64110 , n64360 );
and ( n64506 , n30204 , n64410 );
and ( n64507 , n64505 , n64506 );
xor ( n64508 , n64505 , n64506 );
xor ( n64509 , n64114 , n64358 );
and ( n64510 , n30209 , n64410 );
and ( n64511 , n64509 , n64510 );
xor ( n64512 , n64509 , n64510 );
xor ( n64513 , n64118 , n64356 );
and ( n64514 , n30214 , n64410 );
and ( n64515 , n64513 , n64514 );
xor ( n64516 , n64513 , n64514 );
xor ( n64517 , n64122 , n64354 );
and ( n64518 , n30219 , n64410 );
and ( n64519 , n64517 , n64518 );
xor ( n64520 , n64517 , n64518 );
xor ( n64521 , n64126 , n64352 );
and ( n64522 , n30224 , n64410 );
and ( n64523 , n64521 , n64522 );
xor ( n64524 , n64521 , n64522 );
xor ( n64525 , n64130 , n64350 );
and ( n64526 , n30229 , n64410 );
and ( n64527 , n64525 , n64526 );
xor ( n64528 , n64525 , n64526 );
xor ( n64529 , n64134 , n64348 );
and ( n64530 , n30234 , n64410 );
and ( n64531 , n64529 , n64530 );
xor ( n64532 , n64529 , n64530 );
xor ( n64533 , n64138 , n64346 );
and ( n64534 , n30239 , n64410 );
and ( n64535 , n64533 , n64534 );
xor ( n64536 , n64533 , n64534 );
xor ( n64537 , n64142 , n64344 );
and ( n64538 , n30244 , n64410 );
and ( n64539 , n64537 , n64538 );
xor ( n64540 , n64537 , n64538 );
xor ( n64541 , n64146 , n64342 );
and ( n64542 , n30249 , n64410 );
and ( n64543 , n64541 , n64542 );
xor ( n64544 , n64541 , n64542 );
xor ( n64545 , n64150 , n64340 );
and ( n64546 , n30254 , n64410 );
and ( n64547 , n64545 , n64546 );
xor ( n64548 , n64545 , n64546 );
xor ( n64549 , n64154 , n64338 );
and ( n64550 , n30259 , n64410 );
and ( n64551 , n64549 , n64550 );
xor ( n64552 , n64549 , n64550 );
xor ( n64553 , n64158 , n64336 );
and ( n64554 , n30264 , n64410 );
and ( n64555 , n64553 , n64554 );
xor ( n64556 , n64553 , n64554 );
xor ( n64557 , n64162 , n64334 );
and ( n64558 , n30269 , n64410 );
and ( n64559 , n64557 , n64558 );
xor ( n64560 , n64557 , n64558 );
xor ( n64561 , n64166 , n64332 );
and ( n64562 , n30274 , n64410 );
and ( n64563 , n64561 , n64562 );
xor ( n64564 , n64561 , n64562 );
xor ( n64565 , n64170 , n64330 );
and ( n64566 , n30279 , n64410 );
and ( n64567 , n64565 , n64566 );
xor ( n64568 , n64565 , n64566 );
xor ( n64569 , n64174 , n64328 );
and ( n64570 , n30284 , n64410 );
and ( n64571 , n64569 , n64570 );
xor ( n64572 , n64569 , n64570 );
xor ( n64573 , n64178 , n64326 );
and ( n64574 , n30289 , n64410 );
and ( n64575 , n64573 , n64574 );
xor ( n64576 , n64573 , n64574 );
xor ( n64577 , n64182 , n64324 );
and ( n64578 , n30294 , n64410 );
and ( n64579 , n64577 , n64578 );
xor ( n64580 , n64577 , n64578 );
xor ( n64581 , n64186 , n64322 );
and ( n64582 , n30299 , n64410 );
and ( n64583 , n64581 , n64582 );
xor ( n64584 , n64581 , n64582 );
xor ( n64585 , n64190 , n64320 );
and ( n64586 , n30304 , n64410 );
and ( n64587 , n64585 , n64586 );
xor ( n64588 , n64585 , n64586 );
xor ( n64589 , n64194 , n64318 );
and ( n64590 , n30309 , n64410 );
and ( n64591 , n64589 , n64590 );
xor ( n64592 , n64589 , n64590 );
xor ( n64593 , n64198 , n64316 );
and ( n64594 , n30314 , n64410 );
and ( n64595 , n64593 , n64594 );
xor ( n64596 , n64593 , n64594 );
xor ( n64597 , n64202 , n64314 );
and ( n64598 , n30319 , n64410 );
and ( n64599 , n64597 , n64598 );
xor ( n64600 , n64597 , n64598 );
xor ( n64601 , n64206 , n64312 );
and ( n64602 , n30324 , n64410 );
and ( n64603 , n64601 , n64602 );
xor ( n64604 , n64601 , n64602 );
xor ( n64605 , n64210 , n64310 );
and ( n64606 , n30329 , n64410 );
and ( n64607 , n64605 , n64606 );
xor ( n64608 , n64605 , n64606 );
xor ( n64609 , n64214 , n64308 );
and ( n64610 , n30334 , n64410 );
and ( n64611 , n64609 , n64610 );
xor ( n64612 , n64609 , n64610 );
xor ( n64613 , n64218 , n64306 );
and ( n64614 , n30339 , n64410 );
and ( n64615 , n64613 , n64614 );
xor ( n64616 , n64613 , n64614 );
xor ( n64617 , n64222 , n64304 );
and ( n64618 , n30344 , n64410 );
and ( n64619 , n64617 , n64618 );
xor ( n64620 , n64617 , n64618 );
xor ( n64621 , n64226 , n64302 );
and ( n64622 , n30349 , n64410 );
and ( n64623 , n64621 , n64622 );
xor ( n64624 , n64621 , n64622 );
xor ( n64625 , n64230 , n64300 );
and ( n64626 , n30354 , n64410 );
and ( n64627 , n64625 , n64626 );
xor ( n64628 , n64625 , n64626 );
xor ( n64629 , n64234 , n64298 );
and ( n64630 , n30359 , n64410 );
and ( n64631 , n64629 , n64630 );
xor ( n64632 , n64629 , n64630 );
xor ( n64633 , n64238 , n64296 );
and ( n64634 , n30364 , n64410 );
and ( n64635 , n64633 , n64634 );
xor ( n64636 , n64633 , n64634 );
xor ( n64637 , n64242 , n64294 );
and ( n64638 , n30369 , n64410 );
and ( n64639 , n64637 , n64638 );
xor ( n64640 , n64637 , n64638 );
xor ( n64641 , n64246 , n64292 );
and ( n64642 , n30374 , n64410 );
and ( n64643 , n64641 , n64642 );
xor ( n64644 , n64641 , n64642 );
xor ( n64645 , n64250 , n64290 );
and ( n64646 , n30379 , n64410 );
and ( n64647 , n64645 , n64646 );
xor ( n64648 , n64645 , n64646 );
xor ( n64649 , n64254 , n64288 );
and ( n64650 , n30384 , n64410 );
and ( n64651 , n64649 , n64650 );
xor ( n64652 , n64649 , n64650 );
xor ( n64653 , n64258 , n64286 );
and ( n64654 , n30389 , n64410 );
and ( n64655 , n64653 , n64654 );
xor ( n64656 , n64653 , n64654 );
xor ( n64657 , n64262 , n64284 );
and ( n64658 , n30394 , n64410 );
and ( n64659 , n64657 , n64658 );
xor ( n64660 , n64657 , n64658 );
xor ( n64661 , n64266 , n64282 );
and ( n64662 , n30399 , n64410 );
and ( n64663 , n64661 , n64662 );
xor ( n64664 , n64661 , n64662 );
xor ( n64665 , n64270 , n64280 );
and ( n64666 , n30404 , n64410 );
and ( n64667 , n64665 , n64666 );
xor ( n64668 , n64665 , n64666 );
xor ( n64669 , n64274 , n64278 );
and ( n64670 , n30409 , n64410 );
and ( n64671 , n64669 , n64670 );
buf ( n64672 , n64671 );
and ( n64673 , n64668 , n64672 );
or ( n64674 , n64667 , n64673 );
and ( n64675 , n64664 , n64674 );
or ( n64676 , n64663 , n64675 );
and ( n64677 , n64660 , n64676 );
or ( n64678 , n64659 , n64677 );
and ( n64679 , n64656 , n64678 );
or ( n64680 , n64655 , n64679 );
and ( n64681 , n64652 , n64680 );
or ( n64682 , n64651 , n64681 );
and ( n64683 , n64648 , n64682 );
or ( n64684 , n64647 , n64683 );
and ( n64685 , n64644 , n64684 );
or ( n64686 , n64643 , n64685 );
and ( n64687 , n64640 , n64686 );
or ( n64688 , n64639 , n64687 );
and ( n64689 , n64636 , n64688 );
or ( n64690 , n64635 , n64689 );
and ( n64691 , n64632 , n64690 );
or ( n64692 , n64631 , n64691 );
and ( n64693 , n64628 , n64692 );
or ( n64694 , n64627 , n64693 );
and ( n64695 , n64624 , n64694 );
or ( n64696 , n64623 , n64695 );
and ( n64697 , n64620 , n64696 );
or ( n64698 , n64619 , n64697 );
and ( n64699 , n64616 , n64698 );
or ( n64700 , n64615 , n64699 );
and ( n64701 , n64612 , n64700 );
or ( n64702 , n64611 , n64701 );
and ( n64703 , n64608 , n64702 );
or ( n64704 , n64607 , n64703 );
and ( n64705 , n64604 , n64704 );
or ( n64706 , n64603 , n64705 );
and ( n64707 , n64600 , n64706 );
or ( n64708 , n64599 , n64707 );
and ( n64709 , n64596 , n64708 );
or ( n64710 , n64595 , n64709 );
and ( n64711 , n64592 , n64710 );
or ( n64712 , n64591 , n64711 );
and ( n64713 , n64588 , n64712 );
or ( n64714 , n64587 , n64713 );
and ( n64715 , n64584 , n64714 );
or ( n64716 , n64583 , n64715 );
and ( n64717 , n64580 , n64716 );
or ( n64718 , n64579 , n64717 );
and ( n64719 , n64576 , n64718 );
or ( n64720 , n64575 , n64719 );
and ( n64721 , n64572 , n64720 );
or ( n64722 , n64571 , n64721 );
and ( n64723 , n64568 , n64722 );
or ( n64724 , n64567 , n64723 );
and ( n64725 , n64564 , n64724 );
or ( n64726 , n64563 , n64725 );
and ( n64727 , n64560 , n64726 );
or ( n64728 , n64559 , n64727 );
and ( n64729 , n64556 , n64728 );
or ( n64730 , n64555 , n64729 );
and ( n64731 , n64552 , n64730 );
or ( n64732 , n64551 , n64731 );
and ( n64733 , n64548 , n64732 );
or ( n64734 , n64547 , n64733 );
and ( n64735 , n64544 , n64734 );
or ( n64736 , n64543 , n64735 );
and ( n64737 , n64540 , n64736 );
or ( n64738 , n64539 , n64737 );
and ( n64739 , n64536 , n64738 );
or ( n64740 , n64535 , n64739 );
and ( n64741 , n64532 , n64740 );
or ( n64742 , n64531 , n64741 );
and ( n64743 , n64528 , n64742 );
or ( n64744 , n64527 , n64743 );
and ( n64745 , n64524 , n64744 );
or ( n64746 , n64523 , n64745 );
and ( n64747 , n64520 , n64746 );
or ( n64748 , n64519 , n64747 );
and ( n64749 , n64516 , n64748 );
or ( n64750 , n64515 , n64749 );
and ( n64751 , n64512 , n64750 );
or ( n64752 , n64511 , n64751 );
and ( n64753 , n64508 , n64752 );
or ( n64754 , n64507 , n64753 );
and ( n64755 , n64504 , n64754 );
or ( n64756 , n64503 , n64755 );
and ( n64757 , n64500 , n64756 );
or ( n64758 , n64499 , n64757 );
and ( n64759 , n64496 , n64758 );
or ( n64760 , n64495 , n64759 );
and ( n64761 , n64492 , n64760 );
or ( n64762 , n64491 , n64761 );
and ( n64763 , n64488 , n64762 );
or ( n64764 , n64487 , n64763 );
and ( n64765 , n64484 , n64764 );
or ( n64766 , n64483 , n64765 );
and ( n64767 , n64480 , n64766 );
or ( n64768 , n64479 , n64767 );
and ( n64769 , n64476 , n64768 );
or ( n64770 , n64475 , n64769 );
and ( n64771 , n64472 , n64770 );
or ( n64772 , n64471 , n64771 );
and ( n64773 , n64468 , n64772 );
or ( n64774 , n64467 , n64773 );
and ( n64775 , n64464 , n64774 );
or ( n64776 , n64463 , n64775 );
and ( n64777 , n64460 , n64776 );
or ( n64778 , n64459 , n64777 );
and ( n64779 , n64456 , n64778 );
or ( n64780 , n64455 , n64779 );
and ( n64781 , n64452 , n64780 );
or ( n64782 , n64451 , n64781 );
and ( n64783 , n64448 , n64782 );
or ( n64784 , n64447 , n64783 );
and ( n64785 , n64444 , n64784 );
or ( n64786 , n64443 , n64785 );
and ( n64787 , n64440 , n64786 );
or ( n64788 , n64439 , n64787 );
and ( n64789 , n64436 , n64788 );
or ( n64790 , n64435 , n64789 );
and ( n64791 , n64432 , n64790 );
or ( n64792 , n64431 , n64791 );
and ( n64793 , n64428 , n64792 );
or ( n64794 , n64427 , n64793 );
and ( n64795 , n64424 , n64794 );
or ( n64796 , n64423 , n64795 );
and ( n64797 , n64420 , n64796 );
or ( n64798 , n64419 , n64797 );
and ( n64799 , n64416 , n64798 );
or ( n64800 , n64415 , n64799 );
xor ( n64801 , n64412 , n64800 );
buf ( n64802 , n17982 );
and ( n64803 , n30089 , n64802 );
xor ( n64804 , n64801 , n64803 );
xor ( n64805 , n64416 , n64798 );
and ( n64806 , n30094 , n64802 );
and ( n64807 , n64805 , n64806 );
xor ( n64808 , n64805 , n64806 );
xor ( n64809 , n64420 , n64796 );
and ( n64810 , n30099 , n64802 );
and ( n64811 , n64809 , n64810 );
xor ( n64812 , n64809 , n64810 );
xor ( n64813 , n64424 , n64794 );
and ( n64814 , n30104 , n64802 );
and ( n64815 , n64813 , n64814 );
xor ( n64816 , n64813 , n64814 );
xor ( n64817 , n64428 , n64792 );
and ( n64818 , n30109 , n64802 );
and ( n64819 , n64817 , n64818 );
xor ( n64820 , n64817 , n64818 );
xor ( n64821 , n64432 , n64790 );
and ( n64822 , n30114 , n64802 );
and ( n64823 , n64821 , n64822 );
xor ( n64824 , n64821 , n64822 );
xor ( n64825 , n64436 , n64788 );
and ( n64826 , n30119 , n64802 );
and ( n64827 , n64825 , n64826 );
xor ( n64828 , n64825 , n64826 );
xor ( n64829 , n64440 , n64786 );
and ( n64830 , n30124 , n64802 );
and ( n64831 , n64829 , n64830 );
xor ( n64832 , n64829 , n64830 );
xor ( n64833 , n64444 , n64784 );
and ( n64834 , n30129 , n64802 );
and ( n64835 , n64833 , n64834 );
xor ( n64836 , n64833 , n64834 );
xor ( n64837 , n64448 , n64782 );
and ( n64838 , n30134 , n64802 );
and ( n64839 , n64837 , n64838 );
xor ( n64840 , n64837 , n64838 );
xor ( n64841 , n64452 , n64780 );
and ( n64842 , n30139 , n64802 );
and ( n64843 , n64841 , n64842 );
xor ( n64844 , n64841 , n64842 );
xor ( n64845 , n64456 , n64778 );
and ( n64846 , n30144 , n64802 );
and ( n64847 , n64845 , n64846 );
xor ( n64848 , n64845 , n64846 );
xor ( n64849 , n64460 , n64776 );
and ( n64850 , n30149 , n64802 );
and ( n64851 , n64849 , n64850 );
xor ( n64852 , n64849 , n64850 );
xor ( n64853 , n64464 , n64774 );
and ( n64854 , n30154 , n64802 );
and ( n64855 , n64853 , n64854 );
xor ( n64856 , n64853 , n64854 );
xor ( n64857 , n64468 , n64772 );
and ( n64858 , n30159 , n64802 );
and ( n64859 , n64857 , n64858 );
xor ( n64860 , n64857 , n64858 );
xor ( n64861 , n64472 , n64770 );
and ( n64862 , n30164 , n64802 );
and ( n64863 , n64861 , n64862 );
xor ( n64864 , n64861 , n64862 );
xor ( n64865 , n64476 , n64768 );
and ( n64866 , n30169 , n64802 );
and ( n64867 , n64865 , n64866 );
xor ( n64868 , n64865 , n64866 );
xor ( n64869 , n64480 , n64766 );
and ( n64870 , n30174 , n64802 );
and ( n64871 , n64869 , n64870 );
xor ( n64872 , n64869 , n64870 );
xor ( n64873 , n64484 , n64764 );
and ( n64874 , n30179 , n64802 );
and ( n64875 , n64873 , n64874 );
xor ( n64876 , n64873 , n64874 );
xor ( n64877 , n64488 , n64762 );
and ( n64878 , n30184 , n64802 );
and ( n64879 , n64877 , n64878 );
xor ( n64880 , n64877 , n64878 );
xor ( n64881 , n64492 , n64760 );
and ( n64882 , n30189 , n64802 );
and ( n64883 , n64881 , n64882 );
xor ( n64884 , n64881 , n64882 );
xor ( n64885 , n64496 , n64758 );
and ( n64886 , n30194 , n64802 );
and ( n64887 , n64885 , n64886 );
xor ( n64888 , n64885 , n64886 );
xor ( n64889 , n64500 , n64756 );
and ( n64890 , n30199 , n64802 );
and ( n64891 , n64889 , n64890 );
xor ( n64892 , n64889 , n64890 );
xor ( n64893 , n64504 , n64754 );
and ( n64894 , n30204 , n64802 );
and ( n64895 , n64893 , n64894 );
xor ( n64896 , n64893 , n64894 );
xor ( n64897 , n64508 , n64752 );
and ( n64898 , n30209 , n64802 );
and ( n64899 , n64897 , n64898 );
xor ( n64900 , n64897 , n64898 );
xor ( n64901 , n64512 , n64750 );
and ( n64902 , n30214 , n64802 );
and ( n64903 , n64901 , n64902 );
xor ( n64904 , n64901 , n64902 );
xor ( n64905 , n64516 , n64748 );
and ( n64906 , n30219 , n64802 );
and ( n64907 , n64905 , n64906 );
xor ( n64908 , n64905 , n64906 );
xor ( n64909 , n64520 , n64746 );
and ( n64910 , n30224 , n64802 );
and ( n64911 , n64909 , n64910 );
xor ( n64912 , n64909 , n64910 );
xor ( n64913 , n64524 , n64744 );
and ( n64914 , n30229 , n64802 );
and ( n64915 , n64913 , n64914 );
xor ( n64916 , n64913 , n64914 );
xor ( n64917 , n64528 , n64742 );
and ( n64918 , n30234 , n64802 );
and ( n64919 , n64917 , n64918 );
xor ( n64920 , n64917 , n64918 );
xor ( n64921 , n64532 , n64740 );
and ( n64922 , n30239 , n64802 );
and ( n64923 , n64921 , n64922 );
xor ( n64924 , n64921 , n64922 );
xor ( n64925 , n64536 , n64738 );
and ( n64926 , n30244 , n64802 );
and ( n64927 , n64925 , n64926 );
xor ( n64928 , n64925 , n64926 );
xor ( n64929 , n64540 , n64736 );
and ( n64930 , n30249 , n64802 );
and ( n64931 , n64929 , n64930 );
xor ( n64932 , n64929 , n64930 );
xor ( n64933 , n64544 , n64734 );
and ( n64934 , n30254 , n64802 );
and ( n64935 , n64933 , n64934 );
xor ( n64936 , n64933 , n64934 );
xor ( n64937 , n64548 , n64732 );
and ( n64938 , n30259 , n64802 );
and ( n64939 , n64937 , n64938 );
xor ( n64940 , n64937 , n64938 );
xor ( n64941 , n64552 , n64730 );
and ( n64942 , n30264 , n64802 );
and ( n64943 , n64941 , n64942 );
xor ( n64944 , n64941 , n64942 );
xor ( n64945 , n64556 , n64728 );
and ( n64946 , n30269 , n64802 );
and ( n64947 , n64945 , n64946 );
xor ( n64948 , n64945 , n64946 );
xor ( n64949 , n64560 , n64726 );
and ( n64950 , n30274 , n64802 );
and ( n64951 , n64949 , n64950 );
xor ( n64952 , n64949 , n64950 );
xor ( n64953 , n64564 , n64724 );
and ( n64954 , n30279 , n64802 );
and ( n64955 , n64953 , n64954 );
xor ( n64956 , n64953 , n64954 );
xor ( n64957 , n64568 , n64722 );
and ( n64958 , n30284 , n64802 );
and ( n64959 , n64957 , n64958 );
xor ( n64960 , n64957 , n64958 );
xor ( n64961 , n64572 , n64720 );
and ( n64962 , n30289 , n64802 );
and ( n64963 , n64961 , n64962 );
xor ( n64964 , n64961 , n64962 );
xor ( n64965 , n64576 , n64718 );
and ( n64966 , n30294 , n64802 );
and ( n64967 , n64965 , n64966 );
xor ( n64968 , n64965 , n64966 );
xor ( n64969 , n64580 , n64716 );
and ( n64970 , n30299 , n64802 );
and ( n64971 , n64969 , n64970 );
xor ( n64972 , n64969 , n64970 );
xor ( n64973 , n64584 , n64714 );
and ( n64974 , n30304 , n64802 );
and ( n64975 , n64973 , n64974 );
xor ( n64976 , n64973 , n64974 );
xor ( n64977 , n64588 , n64712 );
and ( n64978 , n30309 , n64802 );
and ( n64979 , n64977 , n64978 );
xor ( n64980 , n64977 , n64978 );
xor ( n64981 , n64592 , n64710 );
and ( n64982 , n30314 , n64802 );
and ( n64983 , n64981 , n64982 );
xor ( n64984 , n64981 , n64982 );
xor ( n64985 , n64596 , n64708 );
and ( n64986 , n30319 , n64802 );
and ( n64987 , n64985 , n64986 );
xor ( n64988 , n64985 , n64986 );
xor ( n64989 , n64600 , n64706 );
and ( n64990 , n30324 , n64802 );
and ( n64991 , n64989 , n64990 );
xor ( n64992 , n64989 , n64990 );
xor ( n64993 , n64604 , n64704 );
and ( n64994 , n30329 , n64802 );
and ( n64995 , n64993 , n64994 );
xor ( n64996 , n64993 , n64994 );
xor ( n64997 , n64608 , n64702 );
and ( n64998 , n30334 , n64802 );
and ( n64999 , n64997 , n64998 );
xor ( n65000 , n64997 , n64998 );
xor ( n65001 , n64612 , n64700 );
and ( n65002 , n30339 , n64802 );
and ( n65003 , n65001 , n65002 );
xor ( n65004 , n65001 , n65002 );
xor ( n65005 , n64616 , n64698 );
and ( n65006 , n30344 , n64802 );
and ( n65007 , n65005 , n65006 );
xor ( n65008 , n65005 , n65006 );
xor ( n65009 , n64620 , n64696 );
and ( n65010 , n30349 , n64802 );
and ( n65011 , n65009 , n65010 );
xor ( n65012 , n65009 , n65010 );
xor ( n65013 , n64624 , n64694 );
and ( n65014 , n30354 , n64802 );
and ( n65015 , n65013 , n65014 );
xor ( n65016 , n65013 , n65014 );
xor ( n65017 , n64628 , n64692 );
and ( n65018 , n30359 , n64802 );
and ( n65019 , n65017 , n65018 );
xor ( n65020 , n65017 , n65018 );
xor ( n65021 , n64632 , n64690 );
and ( n65022 , n30364 , n64802 );
and ( n65023 , n65021 , n65022 );
xor ( n65024 , n65021 , n65022 );
xor ( n65025 , n64636 , n64688 );
and ( n65026 , n30369 , n64802 );
and ( n65027 , n65025 , n65026 );
xor ( n65028 , n65025 , n65026 );
xor ( n65029 , n64640 , n64686 );
and ( n65030 , n30374 , n64802 );
and ( n65031 , n65029 , n65030 );
xor ( n65032 , n65029 , n65030 );
xor ( n65033 , n64644 , n64684 );
and ( n65034 , n30379 , n64802 );
and ( n65035 , n65033 , n65034 );
xor ( n65036 , n65033 , n65034 );
xor ( n65037 , n64648 , n64682 );
and ( n65038 , n30384 , n64802 );
and ( n65039 , n65037 , n65038 );
xor ( n65040 , n65037 , n65038 );
xor ( n65041 , n64652 , n64680 );
and ( n65042 , n30389 , n64802 );
and ( n65043 , n65041 , n65042 );
xor ( n65044 , n65041 , n65042 );
xor ( n65045 , n64656 , n64678 );
and ( n65046 , n30394 , n64802 );
and ( n65047 , n65045 , n65046 );
xor ( n65048 , n65045 , n65046 );
xor ( n65049 , n64660 , n64676 );
and ( n65050 , n30399 , n64802 );
and ( n65051 , n65049 , n65050 );
xor ( n65052 , n65049 , n65050 );
xor ( n65053 , n64664 , n64674 );
and ( n65054 , n30404 , n64802 );
and ( n65055 , n65053 , n65054 );
xor ( n65056 , n65053 , n65054 );
xor ( n65057 , n64668 , n64672 );
and ( n65058 , n30409 , n64802 );
and ( n65059 , n65057 , n65058 );
buf ( n65060 , n65059 );
and ( n65061 , n65056 , n65060 );
or ( n65062 , n65055 , n65061 );
and ( n65063 , n65052 , n65062 );
or ( n65064 , n65051 , n65063 );
and ( n65065 , n65048 , n65064 );
or ( n65066 , n65047 , n65065 );
and ( n65067 , n65044 , n65066 );
or ( n65068 , n65043 , n65067 );
and ( n65069 , n65040 , n65068 );
or ( n65070 , n65039 , n65069 );
and ( n65071 , n65036 , n65070 );
or ( n65072 , n65035 , n65071 );
and ( n65073 , n65032 , n65072 );
or ( n65074 , n65031 , n65073 );
and ( n65075 , n65028 , n65074 );
or ( n65076 , n65027 , n65075 );
and ( n65077 , n65024 , n65076 );
or ( n65078 , n65023 , n65077 );
and ( n65079 , n65020 , n65078 );
or ( n65080 , n65019 , n65079 );
and ( n65081 , n65016 , n65080 );
or ( n65082 , n65015 , n65081 );
and ( n65083 , n65012 , n65082 );
or ( n65084 , n65011 , n65083 );
and ( n65085 , n65008 , n65084 );
or ( n65086 , n65007 , n65085 );
and ( n65087 , n65004 , n65086 );
or ( n65088 , n65003 , n65087 );
and ( n65089 , n65000 , n65088 );
or ( n65090 , n64999 , n65089 );
and ( n65091 , n64996 , n65090 );
or ( n65092 , n64995 , n65091 );
and ( n65093 , n64992 , n65092 );
or ( n65094 , n64991 , n65093 );
and ( n65095 , n64988 , n65094 );
or ( n65096 , n64987 , n65095 );
and ( n65097 , n64984 , n65096 );
or ( n65098 , n64983 , n65097 );
and ( n65099 , n64980 , n65098 );
or ( n65100 , n64979 , n65099 );
and ( n65101 , n64976 , n65100 );
or ( n65102 , n64975 , n65101 );
and ( n65103 , n64972 , n65102 );
or ( n65104 , n64971 , n65103 );
and ( n65105 , n64968 , n65104 );
or ( n65106 , n64967 , n65105 );
and ( n65107 , n64964 , n65106 );
or ( n65108 , n64963 , n65107 );
and ( n65109 , n64960 , n65108 );
or ( n65110 , n64959 , n65109 );
and ( n65111 , n64956 , n65110 );
or ( n65112 , n64955 , n65111 );
and ( n65113 , n64952 , n65112 );
or ( n65114 , n64951 , n65113 );
and ( n65115 , n64948 , n65114 );
or ( n65116 , n64947 , n65115 );
and ( n65117 , n64944 , n65116 );
or ( n65118 , n64943 , n65117 );
and ( n65119 , n64940 , n65118 );
or ( n65120 , n64939 , n65119 );
and ( n65121 , n64936 , n65120 );
or ( n65122 , n64935 , n65121 );
and ( n65123 , n64932 , n65122 );
or ( n65124 , n64931 , n65123 );
and ( n65125 , n64928 , n65124 );
or ( n65126 , n64927 , n65125 );
and ( n65127 , n64924 , n65126 );
or ( n65128 , n64923 , n65127 );
and ( n65129 , n64920 , n65128 );
or ( n65130 , n64919 , n65129 );
and ( n65131 , n64916 , n65130 );
or ( n65132 , n64915 , n65131 );
and ( n65133 , n64912 , n65132 );
or ( n65134 , n64911 , n65133 );
and ( n65135 , n64908 , n65134 );
or ( n65136 , n64907 , n65135 );
and ( n65137 , n64904 , n65136 );
or ( n65138 , n64903 , n65137 );
and ( n65139 , n64900 , n65138 );
or ( n65140 , n64899 , n65139 );
and ( n65141 , n64896 , n65140 );
or ( n65142 , n64895 , n65141 );
and ( n65143 , n64892 , n65142 );
or ( n65144 , n64891 , n65143 );
and ( n65145 , n64888 , n65144 );
or ( n65146 , n64887 , n65145 );
and ( n65147 , n64884 , n65146 );
or ( n65148 , n64883 , n65147 );
and ( n65149 , n64880 , n65148 );
or ( n65150 , n64879 , n65149 );
and ( n65151 , n64876 , n65150 );
or ( n65152 , n64875 , n65151 );
and ( n65153 , n64872 , n65152 );
or ( n65154 , n64871 , n65153 );
and ( n65155 , n64868 , n65154 );
or ( n65156 , n64867 , n65155 );
and ( n65157 , n64864 , n65156 );
or ( n65158 , n64863 , n65157 );
and ( n65159 , n64860 , n65158 );
or ( n65160 , n64859 , n65159 );
and ( n65161 , n64856 , n65160 );
or ( n65162 , n64855 , n65161 );
and ( n65163 , n64852 , n65162 );
or ( n65164 , n64851 , n65163 );
and ( n65165 , n64848 , n65164 );
or ( n65166 , n64847 , n65165 );
and ( n65167 , n64844 , n65166 );
or ( n65168 , n64843 , n65167 );
and ( n65169 , n64840 , n65168 );
or ( n65170 , n64839 , n65169 );
and ( n65171 , n64836 , n65170 );
or ( n65172 , n64835 , n65171 );
and ( n65173 , n64832 , n65172 );
or ( n65174 , n64831 , n65173 );
and ( n65175 , n64828 , n65174 );
or ( n65176 , n64827 , n65175 );
and ( n65177 , n64824 , n65176 );
or ( n65178 , n64823 , n65177 );
and ( n65179 , n64820 , n65178 );
or ( n65180 , n64819 , n65179 );
and ( n65181 , n64816 , n65180 );
or ( n65182 , n64815 , n65181 );
and ( n65183 , n64812 , n65182 );
or ( n65184 , n64811 , n65183 );
and ( n65185 , n64808 , n65184 );
or ( n65186 , n64807 , n65185 );
xor ( n65187 , n64804 , n65186 );
buf ( n65188 , n17980 );
and ( n65189 , n30094 , n65188 );
xor ( n65190 , n65187 , n65189 );
xor ( n65191 , n64808 , n65184 );
and ( n65192 , n30099 , n65188 );
and ( n65193 , n65191 , n65192 );
xor ( n65194 , n65191 , n65192 );
xor ( n65195 , n64812 , n65182 );
and ( n65196 , n30104 , n65188 );
and ( n65197 , n65195 , n65196 );
xor ( n65198 , n65195 , n65196 );
xor ( n65199 , n64816 , n65180 );
and ( n65200 , n30109 , n65188 );
and ( n65201 , n65199 , n65200 );
xor ( n65202 , n65199 , n65200 );
xor ( n65203 , n64820 , n65178 );
and ( n65204 , n30114 , n65188 );
and ( n65205 , n65203 , n65204 );
xor ( n65206 , n65203 , n65204 );
xor ( n65207 , n64824 , n65176 );
and ( n65208 , n30119 , n65188 );
and ( n65209 , n65207 , n65208 );
xor ( n65210 , n65207 , n65208 );
xor ( n65211 , n64828 , n65174 );
and ( n65212 , n30124 , n65188 );
and ( n65213 , n65211 , n65212 );
xor ( n65214 , n65211 , n65212 );
xor ( n65215 , n64832 , n65172 );
and ( n65216 , n30129 , n65188 );
and ( n65217 , n65215 , n65216 );
xor ( n65218 , n65215 , n65216 );
xor ( n65219 , n64836 , n65170 );
and ( n65220 , n30134 , n65188 );
and ( n65221 , n65219 , n65220 );
xor ( n65222 , n65219 , n65220 );
xor ( n65223 , n64840 , n65168 );
and ( n65224 , n30139 , n65188 );
and ( n65225 , n65223 , n65224 );
xor ( n65226 , n65223 , n65224 );
xor ( n65227 , n64844 , n65166 );
and ( n65228 , n30144 , n65188 );
and ( n65229 , n65227 , n65228 );
xor ( n65230 , n65227 , n65228 );
xor ( n65231 , n64848 , n65164 );
and ( n65232 , n30149 , n65188 );
and ( n65233 , n65231 , n65232 );
xor ( n65234 , n65231 , n65232 );
xor ( n65235 , n64852 , n65162 );
and ( n65236 , n30154 , n65188 );
and ( n65237 , n65235 , n65236 );
xor ( n65238 , n65235 , n65236 );
xor ( n65239 , n64856 , n65160 );
and ( n65240 , n30159 , n65188 );
and ( n65241 , n65239 , n65240 );
xor ( n65242 , n65239 , n65240 );
xor ( n65243 , n64860 , n65158 );
and ( n65244 , n30164 , n65188 );
and ( n65245 , n65243 , n65244 );
xor ( n65246 , n65243 , n65244 );
xor ( n65247 , n64864 , n65156 );
and ( n65248 , n30169 , n65188 );
and ( n65249 , n65247 , n65248 );
xor ( n65250 , n65247 , n65248 );
xor ( n65251 , n64868 , n65154 );
and ( n65252 , n30174 , n65188 );
and ( n65253 , n65251 , n65252 );
xor ( n65254 , n65251 , n65252 );
xor ( n65255 , n64872 , n65152 );
and ( n65256 , n30179 , n65188 );
and ( n65257 , n65255 , n65256 );
xor ( n65258 , n65255 , n65256 );
xor ( n65259 , n64876 , n65150 );
and ( n65260 , n30184 , n65188 );
and ( n65261 , n65259 , n65260 );
xor ( n65262 , n65259 , n65260 );
xor ( n65263 , n64880 , n65148 );
and ( n65264 , n30189 , n65188 );
and ( n65265 , n65263 , n65264 );
xor ( n65266 , n65263 , n65264 );
xor ( n65267 , n64884 , n65146 );
and ( n65268 , n30194 , n65188 );
and ( n65269 , n65267 , n65268 );
xor ( n65270 , n65267 , n65268 );
xor ( n65271 , n64888 , n65144 );
and ( n65272 , n30199 , n65188 );
and ( n65273 , n65271 , n65272 );
xor ( n65274 , n65271 , n65272 );
xor ( n65275 , n64892 , n65142 );
and ( n65276 , n30204 , n65188 );
and ( n65277 , n65275 , n65276 );
xor ( n65278 , n65275 , n65276 );
xor ( n65279 , n64896 , n65140 );
and ( n65280 , n30209 , n65188 );
and ( n65281 , n65279 , n65280 );
xor ( n65282 , n65279 , n65280 );
xor ( n65283 , n64900 , n65138 );
and ( n65284 , n30214 , n65188 );
and ( n65285 , n65283 , n65284 );
xor ( n65286 , n65283 , n65284 );
xor ( n65287 , n64904 , n65136 );
and ( n65288 , n30219 , n65188 );
and ( n65289 , n65287 , n65288 );
xor ( n65290 , n65287 , n65288 );
xor ( n65291 , n64908 , n65134 );
and ( n65292 , n30224 , n65188 );
and ( n65293 , n65291 , n65292 );
xor ( n65294 , n65291 , n65292 );
xor ( n65295 , n64912 , n65132 );
and ( n65296 , n30229 , n65188 );
and ( n65297 , n65295 , n65296 );
xor ( n65298 , n65295 , n65296 );
xor ( n65299 , n64916 , n65130 );
and ( n65300 , n30234 , n65188 );
and ( n65301 , n65299 , n65300 );
xor ( n65302 , n65299 , n65300 );
xor ( n65303 , n64920 , n65128 );
and ( n65304 , n30239 , n65188 );
and ( n65305 , n65303 , n65304 );
xor ( n65306 , n65303 , n65304 );
xor ( n65307 , n64924 , n65126 );
and ( n65308 , n30244 , n65188 );
and ( n65309 , n65307 , n65308 );
xor ( n65310 , n65307 , n65308 );
xor ( n65311 , n64928 , n65124 );
and ( n65312 , n30249 , n65188 );
and ( n65313 , n65311 , n65312 );
xor ( n65314 , n65311 , n65312 );
xor ( n65315 , n64932 , n65122 );
and ( n65316 , n30254 , n65188 );
and ( n65317 , n65315 , n65316 );
xor ( n65318 , n65315 , n65316 );
xor ( n65319 , n64936 , n65120 );
and ( n65320 , n30259 , n65188 );
and ( n65321 , n65319 , n65320 );
xor ( n65322 , n65319 , n65320 );
xor ( n65323 , n64940 , n65118 );
and ( n65324 , n30264 , n65188 );
and ( n65325 , n65323 , n65324 );
xor ( n65326 , n65323 , n65324 );
xor ( n65327 , n64944 , n65116 );
and ( n65328 , n30269 , n65188 );
and ( n65329 , n65327 , n65328 );
xor ( n65330 , n65327 , n65328 );
xor ( n65331 , n64948 , n65114 );
and ( n65332 , n30274 , n65188 );
and ( n65333 , n65331 , n65332 );
xor ( n65334 , n65331 , n65332 );
xor ( n65335 , n64952 , n65112 );
and ( n65336 , n30279 , n65188 );
and ( n65337 , n65335 , n65336 );
xor ( n65338 , n65335 , n65336 );
xor ( n65339 , n64956 , n65110 );
and ( n65340 , n30284 , n65188 );
and ( n65341 , n65339 , n65340 );
xor ( n65342 , n65339 , n65340 );
xor ( n65343 , n64960 , n65108 );
and ( n65344 , n30289 , n65188 );
and ( n65345 , n65343 , n65344 );
xor ( n65346 , n65343 , n65344 );
xor ( n65347 , n64964 , n65106 );
and ( n65348 , n30294 , n65188 );
and ( n65349 , n65347 , n65348 );
xor ( n65350 , n65347 , n65348 );
xor ( n65351 , n64968 , n65104 );
and ( n65352 , n30299 , n65188 );
and ( n65353 , n65351 , n65352 );
xor ( n65354 , n65351 , n65352 );
xor ( n65355 , n64972 , n65102 );
and ( n65356 , n30304 , n65188 );
and ( n65357 , n65355 , n65356 );
xor ( n65358 , n65355 , n65356 );
xor ( n65359 , n64976 , n65100 );
and ( n65360 , n30309 , n65188 );
and ( n65361 , n65359 , n65360 );
xor ( n65362 , n65359 , n65360 );
xor ( n65363 , n64980 , n65098 );
and ( n65364 , n30314 , n65188 );
and ( n65365 , n65363 , n65364 );
xor ( n65366 , n65363 , n65364 );
xor ( n65367 , n64984 , n65096 );
and ( n65368 , n30319 , n65188 );
and ( n65369 , n65367 , n65368 );
xor ( n65370 , n65367 , n65368 );
xor ( n65371 , n64988 , n65094 );
and ( n65372 , n30324 , n65188 );
and ( n65373 , n65371 , n65372 );
xor ( n65374 , n65371 , n65372 );
xor ( n65375 , n64992 , n65092 );
and ( n65376 , n30329 , n65188 );
and ( n65377 , n65375 , n65376 );
xor ( n65378 , n65375 , n65376 );
xor ( n65379 , n64996 , n65090 );
and ( n65380 , n30334 , n65188 );
and ( n65381 , n65379 , n65380 );
xor ( n65382 , n65379 , n65380 );
xor ( n65383 , n65000 , n65088 );
and ( n65384 , n30339 , n65188 );
and ( n65385 , n65383 , n65384 );
xor ( n65386 , n65383 , n65384 );
xor ( n65387 , n65004 , n65086 );
and ( n65388 , n30344 , n65188 );
and ( n65389 , n65387 , n65388 );
xor ( n65390 , n65387 , n65388 );
xor ( n65391 , n65008 , n65084 );
and ( n65392 , n30349 , n65188 );
and ( n65393 , n65391 , n65392 );
xor ( n65394 , n65391 , n65392 );
xor ( n65395 , n65012 , n65082 );
and ( n65396 , n30354 , n65188 );
and ( n65397 , n65395 , n65396 );
xor ( n65398 , n65395 , n65396 );
xor ( n65399 , n65016 , n65080 );
and ( n65400 , n30359 , n65188 );
and ( n65401 , n65399 , n65400 );
xor ( n65402 , n65399 , n65400 );
xor ( n65403 , n65020 , n65078 );
and ( n65404 , n30364 , n65188 );
and ( n65405 , n65403 , n65404 );
xor ( n65406 , n65403 , n65404 );
xor ( n65407 , n65024 , n65076 );
and ( n65408 , n30369 , n65188 );
and ( n65409 , n65407 , n65408 );
xor ( n65410 , n65407 , n65408 );
xor ( n65411 , n65028 , n65074 );
and ( n65412 , n30374 , n65188 );
and ( n65413 , n65411 , n65412 );
xor ( n65414 , n65411 , n65412 );
xor ( n65415 , n65032 , n65072 );
and ( n65416 , n30379 , n65188 );
and ( n65417 , n65415 , n65416 );
xor ( n65418 , n65415 , n65416 );
xor ( n65419 , n65036 , n65070 );
and ( n65420 , n30384 , n65188 );
and ( n65421 , n65419 , n65420 );
xor ( n65422 , n65419 , n65420 );
xor ( n65423 , n65040 , n65068 );
and ( n65424 , n30389 , n65188 );
and ( n65425 , n65423 , n65424 );
xor ( n65426 , n65423 , n65424 );
xor ( n65427 , n65044 , n65066 );
and ( n65428 , n30394 , n65188 );
and ( n65429 , n65427 , n65428 );
xor ( n65430 , n65427 , n65428 );
xor ( n65431 , n65048 , n65064 );
and ( n65432 , n30399 , n65188 );
and ( n65433 , n65431 , n65432 );
xor ( n65434 , n65431 , n65432 );
xor ( n65435 , n65052 , n65062 );
and ( n65436 , n30404 , n65188 );
and ( n65437 , n65435 , n65436 );
xor ( n65438 , n65435 , n65436 );
xor ( n65439 , n65056 , n65060 );
and ( n65440 , n30409 , n65188 );
and ( n65441 , n65439 , n65440 );
buf ( n65442 , n65441 );
and ( n65443 , n65438 , n65442 );
or ( n65444 , n65437 , n65443 );
and ( n65445 , n65434 , n65444 );
or ( n65446 , n65433 , n65445 );
and ( n65447 , n65430 , n65446 );
or ( n65448 , n65429 , n65447 );
and ( n65449 , n65426 , n65448 );
or ( n65450 , n65425 , n65449 );
and ( n65451 , n65422 , n65450 );
or ( n65452 , n65421 , n65451 );
and ( n65453 , n65418 , n65452 );
or ( n65454 , n65417 , n65453 );
and ( n65455 , n65414 , n65454 );
or ( n65456 , n65413 , n65455 );
and ( n65457 , n65410 , n65456 );
or ( n65458 , n65409 , n65457 );
and ( n65459 , n65406 , n65458 );
or ( n65460 , n65405 , n65459 );
and ( n65461 , n65402 , n65460 );
or ( n65462 , n65401 , n65461 );
and ( n65463 , n65398 , n65462 );
or ( n65464 , n65397 , n65463 );
and ( n65465 , n65394 , n65464 );
or ( n65466 , n65393 , n65465 );
and ( n65467 , n65390 , n65466 );
or ( n65468 , n65389 , n65467 );
and ( n65469 , n65386 , n65468 );
or ( n65470 , n65385 , n65469 );
and ( n65471 , n65382 , n65470 );
or ( n65472 , n65381 , n65471 );
and ( n65473 , n65378 , n65472 );
or ( n65474 , n65377 , n65473 );
and ( n65475 , n65374 , n65474 );
or ( n65476 , n65373 , n65475 );
and ( n65477 , n65370 , n65476 );
or ( n65478 , n65369 , n65477 );
and ( n65479 , n65366 , n65478 );
or ( n65480 , n65365 , n65479 );
and ( n65481 , n65362 , n65480 );
or ( n65482 , n65361 , n65481 );
and ( n65483 , n65358 , n65482 );
or ( n65484 , n65357 , n65483 );
and ( n65485 , n65354 , n65484 );
or ( n65486 , n65353 , n65485 );
and ( n65487 , n65350 , n65486 );
or ( n65488 , n65349 , n65487 );
and ( n65489 , n65346 , n65488 );
or ( n65490 , n65345 , n65489 );
and ( n65491 , n65342 , n65490 );
or ( n65492 , n65341 , n65491 );
and ( n65493 , n65338 , n65492 );
or ( n65494 , n65337 , n65493 );
and ( n65495 , n65334 , n65494 );
or ( n65496 , n65333 , n65495 );
and ( n65497 , n65330 , n65496 );
or ( n65498 , n65329 , n65497 );
and ( n65499 , n65326 , n65498 );
or ( n65500 , n65325 , n65499 );
and ( n65501 , n65322 , n65500 );
or ( n65502 , n65321 , n65501 );
and ( n65503 , n65318 , n65502 );
or ( n65504 , n65317 , n65503 );
and ( n65505 , n65314 , n65504 );
or ( n65506 , n65313 , n65505 );
and ( n65507 , n65310 , n65506 );
or ( n65508 , n65309 , n65507 );
and ( n65509 , n65306 , n65508 );
or ( n65510 , n65305 , n65509 );
and ( n65511 , n65302 , n65510 );
or ( n65512 , n65301 , n65511 );
and ( n65513 , n65298 , n65512 );
or ( n65514 , n65297 , n65513 );
and ( n65515 , n65294 , n65514 );
or ( n65516 , n65293 , n65515 );
and ( n65517 , n65290 , n65516 );
or ( n65518 , n65289 , n65517 );
and ( n65519 , n65286 , n65518 );
or ( n65520 , n65285 , n65519 );
and ( n65521 , n65282 , n65520 );
or ( n65522 , n65281 , n65521 );
and ( n65523 , n65278 , n65522 );
or ( n65524 , n65277 , n65523 );
and ( n65525 , n65274 , n65524 );
or ( n65526 , n65273 , n65525 );
and ( n65527 , n65270 , n65526 );
or ( n65528 , n65269 , n65527 );
and ( n65529 , n65266 , n65528 );
or ( n65530 , n65265 , n65529 );
and ( n65531 , n65262 , n65530 );
or ( n65532 , n65261 , n65531 );
and ( n65533 , n65258 , n65532 );
or ( n65534 , n65257 , n65533 );
and ( n65535 , n65254 , n65534 );
or ( n65536 , n65253 , n65535 );
and ( n65537 , n65250 , n65536 );
or ( n65538 , n65249 , n65537 );
and ( n65539 , n65246 , n65538 );
or ( n65540 , n65245 , n65539 );
and ( n65541 , n65242 , n65540 );
or ( n65542 , n65241 , n65541 );
and ( n65543 , n65238 , n65542 );
or ( n65544 , n65237 , n65543 );
and ( n65545 , n65234 , n65544 );
or ( n65546 , n65233 , n65545 );
and ( n65547 , n65230 , n65546 );
or ( n65548 , n65229 , n65547 );
and ( n65549 , n65226 , n65548 );
or ( n65550 , n65225 , n65549 );
and ( n65551 , n65222 , n65550 );
or ( n65552 , n65221 , n65551 );
and ( n65553 , n65218 , n65552 );
or ( n65554 , n65217 , n65553 );
and ( n65555 , n65214 , n65554 );
or ( n65556 , n65213 , n65555 );
and ( n65557 , n65210 , n65556 );
or ( n65558 , n65209 , n65557 );
and ( n65559 , n65206 , n65558 );
or ( n65560 , n65205 , n65559 );
and ( n65561 , n65202 , n65560 );
or ( n65562 , n65201 , n65561 );
and ( n65563 , n65198 , n65562 );
or ( n65564 , n65197 , n65563 );
and ( n65565 , n65194 , n65564 );
or ( n65566 , n65193 , n65565 );
xor ( n65567 , n65190 , n65566 );
buf ( n65568 , n17978 );
and ( n65569 , n30099 , n65568 );
xor ( n65570 , n65567 , n65569 );
xor ( n65571 , n65194 , n65564 );
and ( n65572 , n30104 , n65568 );
and ( n65573 , n65571 , n65572 );
xor ( n65574 , n65571 , n65572 );
xor ( n65575 , n65198 , n65562 );
and ( n65576 , n30109 , n65568 );
and ( n65577 , n65575 , n65576 );
xor ( n65578 , n65575 , n65576 );
xor ( n65579 , n65202 , n65560 );
and ( n65580 , n30114 , n65568 );
and ( n65581 , n65579 , n65580 );
xor ( n65582 , n65579 , n65580 );
xor ( n65583 , n65206 , n65558 );
and ( n65584 , n30119 , n65568 );
and ( n65585 , n65583 , n65584 );
xor ( n65586 , n65583 , n65584 );
xor ( n65587 , n65210 , n65556 );
and ( n65588 , n30124 , n65568 );
and ( n65589 , n65587 , n65588 );
xor ( n65590 , n65587 , n65588 );
xor ( n65591 , n65214 , n65554 );
and ( n65592 , n30129 , n65568 );
and ( n65593 , n65591 , n65592 );
xor ( n65594 , n65591 , n65592 );
xor ( n65595 , n65218 , n65552 );
and ( n65596 , n30134 , n65568 );
and ( n65597 , n65595 , n65596 );
xor ( n65598 , n65595 , n65596 );
xor ( n65599 , n65222 , n65550 );
and ( n65600 , n30139 , n65568 );
and ( n65601 , n65599 , n65600 );
xor ( n65602 , n65599 , n65600 );
xor ( n65603 , n65226 , n65548 );
and ( n65604 , n30144 , n65568 );
and ( n65605 , n65603 , n65604 );
xor ( n65606 , n65603 , n65604 );
xor ( n65607 , n65230 , n65546 );
and ( n65608 , n30149 , n65568 );
and ( n65609 , n65607 , n65608 );
xor ( n65610 , n65607 , n65608 );
xor ( n65611 , n65234 , n65544 );
and ( n65612 , n30154 , n65568 );
and ( n65613 , n65611 , n65612 );
xor ( n65614 , n65611 , n65612 );
xor ( n65615 , n65238 , n65542 );
and ( n65616 , n30159 , n65568 );
and ( n65617 , n65615 , n65616 );
xor ( n65618 , n65615 , n65616 );
xor ( n65619 , n65242 , n65540 );
and ( n65620 , n30164 , n65568 );
and ( n65621 , n65619 , n65620 );
xor ( n65622 , n65619 , n65620 );
xor ( n65623 , n65246 , n65538 );
and ( n65624 , n30169 , n65568 );
and ( n65625 , n65623 , n65624 );
xor ( n65626 , n65623 , n65624 );
xor ( n65627 , n65250 , n65536 );
and ( n65628 , n30174 , n65568 );
and ( n65629 , n65627 , n65628 );
xor ( n65630 , n65627 , n65628 );
xor ( n65631 , n65254 , n65534 );
and ( n65632 , n30179 , n65568 );
and ( n65633 , n65631 , n65632 );
xor ( n65634 , n65631 , n65632 );
xor ( n65635 , n65258 , n65532 );
and ( n65636 , n30184 , n65568 );
and ( n65637 , n65635 , n65636 );
xor ( n65638 , n65635 , n65636 );
xor ( n65639 , n65262 , n65530 );
and ( n65640 , n30189 , n65568 );
and ( n65641 , n65639 , n65640 );
xor ( n65642 , n65639 , n65640 );
xor ( n65643 , n65266 , n65528 );
and ( n65644 , n30194 , n65568 );
and ( n65645 , n65643 , n65644 );
xor ( n65646 , n65643 , n65644 );
xor ( n65647 , n65270 , n65526 );
and ( n65648 , n30199 , n65568 );
and ( n65649 , n65647 , n65648 );
xor ( n65650 , n65647 , n65648 );
xor ( n65651 , n65274 , n65524 );
and ( n65652 , n30204 , n65568 );
and ( n65653 , n65651 , n65652 );
xor ( n65654 , n65651 , n65652 );
xor ( n65655 , n65278 , n65522 );
and ( n65656 , n30209 , n65568 );
and ( n65657 , n65655 , n65656 );
xor ( n65658 , n65655 , n65656 );
xor ( n65659 , n65282 , n65520 );
and ( n65660 , n30214 , n65568 );
and ( n65661 , n65659 , n65660 );
xor ( n65662 , n65659 , n65660 );
xor ( n65663 , n65286 , n65518 );
and ( n65664 , n30219 , n65568 );
and ( n65665 , n65663 , n65664 );
xor ( n65666 , n65663 , n65664 );
xor ( n65667 , n65290 , n65516 );
and ( n65668 , n30224 , n65568 );
and ( n65669 , n65667 , n65668 );
xor ( n65670 , n65667 , n65668 );
xor ( n65671 , n65294 , n65514 );
and ( n65672 , n30229 , n65568 );
and ( n65673 , n65671 , n65672 );
xor ( n65674 , n65671 , n65672 );
xor ( n65675 , n65298 , n65512 );
and ( n65676 , n30234 , n65568 );
and ( n65677 , n65675 , n65676 );
xor ( n65678 , n65675 , n65676 );
xor ( n65679 , n65302 , n65510 );
and ( n65680 , n30239 , n65568 );
and ( n65681 , n65679 , n65680 );
xor ( n65682 , n65679 , n65680 );
xor ( n65683 , n65306 , n65508 );
and ( n65684 , n30244 , n65568 );
and ( n65685 , n65683 , n65684 );
xor ( n65686 , n65683 , n65684 );
xor ( n65687 , n65310 , n65506 );
and ( n65688 , n30249 , n65568 );
and ( n65689 , n65687 , n65688 );
xor ( n65690 , n65687 , n65688 );
xor ( n65691 , n65314 , n65504 );
and ( n65692 , n30254 , n65568 );
and ( n65693 , n65691 , n65692 );
xor ( n65694 , n65691 , n65692 );
xor ( n65695 , n65318 , n65502 );
and ( n65696 , n30259 , n65568 );
and ( n65697 , n65695 , n65696 );
xor ( n65698 , n65695 , n65696 );
xor ( n65699 , n65322 , n65500 );
and ( n65700 , n30264 , n65568 );
and ( n65701 , n65699 , n65700 );
xor ( n65702 , n65699 , n65700 );
xor ( n65703 , n65326 , n65498 );
and ( n65704 , n30269 , n65568 );
and ( n65705 , n65703 , n65704 );
xor ( n65706 , n65703 , n65704 );
xor ( n65707 , n65330 , n65496 );
and ( n65708 , n30274 , n65568 );
and ( n65709 , n65707 , n65708 );
xor ( n65710 , n65707 , n65708 );
xor ( n65711 , n65334 , n65494 );
and ( n65712 , n30279 , n65568 );
and ( n65713 , n65711 , n65712 );
xor ( n65714 , n65711 , n65712 );
xor ( n65715 , n65338 , n65492 );
and ( n65716 , n30284 , n65568 );
and ( n65717 , n65715 , n65716 );
xor ( n65718 , n65715 , n65716 );
xor ( n65719 , n65342 , n65490 );
and ( n65720 , n30289 , n65568 );
and ( n65721 , n65719 , n65720 );
xor ( n65722 , n65719 , n65720 );
xor ( n65723 , n65346 , n65488 );
and ( n65724 , n30294 , n65568 );
and ( n65725 , n65723 , n65724 );
xor ( n65726 , n65723 , n65724 );
xor ( n65727 , n65350 , n65486 );
and ( n65728 , n30299 , n65568 );
and ( n65729 , n65727 , n65728 );
xor ( n65730 , n65727 , n65728 );
xor ( n65731 , n65354 , n65484 );
and ( n65732 , n30304 , n65568 );
and ( n65733 , n65731 , n65732 );
xor ( n65734 , n65731 , n65732 );
xor ( n65735 , n65358 , n65482 );
and ( n65736 , n30309 , n65568 );
and ( n65737 , n65735 , n65736 );
xor ( n65738 , n65735 , n65736 );
xor ( n65739 , n65362 , n65480 );
and ( n65740 , n30314 , n65568 );
and ( n65741 , n65739 , n65740 );
xor ( n65742 , n65739 , n65740 );
xor ( n65743 , n65366 , n65478 );
and ( n65744 , n30319 , n65568 );
and ( n65745 , n65743 , n65744 );
xor ( n65746 , n65743 , n65744 );
xor ( n65747 , n65370 , n65476 );
and ( n65748 , n30324 , n65568 );
and ( n65749 , n65747 , n65748 );
xor ( n65750 , n65747 , n65748 );
xor ( n65751 , n65374 , n65474 );
and ( n65752 , n30329 , n65568 );
and ( n65753 , n65751 , n65752 );
xor ( n65754 , n65751 , n65752 );
xor ( n65755 , n65378 , n65472 );
and ( n65756 , n30334 , n65568 );
and ( n65757 , n65755 , n65756 );
xor ( n65758 , n65755 , n65756 );
xor ( n65759 , n65382 , n65470 );
and ( n65760 , n30339 , n65568 );
and ( n65761 , n65759 , n65760 );
xor ( n65762 , n65759 , n65760 );
xor ( n65763 , n65386 , n65468 );
and ( n65764 , n30344 , n65568 );
and ( n65765 , n65763 , n65764 );
xor ( n65766 , n65763 , n65764 );
xor ( n65767 , n65390 , n65466 );
and ( n65768 , n30349 , n65568 );
and ( n65769 , n65767 , n65768 );
xor ( n65770 , n65767 , n65768 );
xor ( n65771 , n65394 , n65464 );
and ( n65772 , n30354 , n65568 );
and ( n65773 , n65771 , n65772 );
xor ( n65774 , n65771 , n65772 );
xor ( n65775 , n65398 , n65462 );
and ( n65776 , n30359 , n65568 );
and ( n65777 , n65775 , n65776 );
xor ( n65778 , n65775 , n65776 );
xor ( n65779 , n65402 , n65460 );
and ( n65780 , n30364 , n65568 );
and ( n65781 , n65779 , n65780 );
xor ( n65782 , n65779 , n65780 );
xor ( n65783 , n65406 , n65458 );
and ( n65784 , n30369 , n65568 );
and ( n65785 , n65783 , n65784 );
xor ( n65786 , n65783 , n65784 );
xor ( n65787 , n65410 , n65456 );
and ( n65788 , n30374 , n65568 );
and ( n65789 , n65787 , n65788 );
xor ( n65790 , n65787 , n65788 );
xor ( n65791 , n65414 , n65454 );
and ( n65792 , n30379 , n65568 );
and ( n65793 , n65791 , n65792 );
xor ( n65794 , n65791 , n65792 );
xor ( n65795 , n65418 , n65452 );
and ( n65796 , n30384 , n65568 );
and ( n65797 , n65795 , n65796 );
xor ( n65798 , n65795 , n65796 );
xor ( n65799 , n65422 , n65450 );
and ( n65800 , n30389 , n65568 );
and ( n65801 , n65799 , n65800 );
xor ( n65802 , n65799 , n65800 );
xor ( n65803 , n65426 , n65448 );
and ( n65804 , n30394 , n65568 );
and ( n65805 , n65803 , n65804 );
xor ( n65806 , n65803 , n65804 );
xor ( n65807 , n65430 , n65446 );
and ( n65808 , n30399 , n65568 );
and ( n65809 , n65807 , n65808 );
xor ( n65810 , n65807 , n65808 );
xor ( n65811 , n65434 , n65444 );
and ( n65812 , n30404 , n65568 );
and ( n65813 , n65811 , n65812 );
xor ( n65814 , n65811 , n65812 );
xor ( n65815 , n65438 , n65442 );
and ( n65816 , n30409 , n65568 );
and ( n65817 , n65815 , n65816 );
buf ( n65818 , n65817 );
and ( n65819 , n65814 , n65818 );
or ( n65820 , n65813 , n65819 );
and ( n65821 , n65810 , n65820 );
or ( n65822 , n65809 , n65821 );
and ( n65823 , n65806 , n65822 );
or ( n65824 , n65805 , n65823 );
and ( n65825 , n65802 , n65824 );
or ( n65826 , n65801 , n65825 );
and ( n65827 , n65798 , n65826 );
or ( n65828 , n65797 , n65827 );
and ( n65829 , n65794 , n65828 );
or ( n65830 , n65793 , n65829 );
and ( n65831 , n65790 , n65830 );
or ( n65832 , n65789 , n65831 );
and ( n65833 , n65786 , n65832 );
or ( n65834 , n65785 , n65833 );
and ( n65835 , n65782 , n65834 );
or ( n65836 , n65781 , n65835 );
and ( n65837 , n65778 , n65836 );
or ( n65838 , n65777 , n65837 );
and ( n65839 , n65774 , n65838 );
or ( n65840 , n65773 , n65839 );
and ( n65841 , n65770 , n65840 );
or ( n65842 , n65769 , n65841 );
and ( n65843 , n65766 , n65842 );
or ( n65844 , n65765 , n65843 );
and ( n65845 , n65762 , n65844 );
or ( n65846 , n65761 , n65845 );
and ( n65847 , n65758 , n65846 );
or ( n65848 , n65757 , n65847 );
and ( n65849 , n65754 , n65848 );
or ( n65850 , n65753 , n65849 );
and ( n65851 , n65750 , n65850 );
or ( n65852 , n65749 , n65851 );
and ( n65853 , n65746 , n65852 );
or ( n65854 , n65745 , n65853 );
and ( n65855 , n65742 , n65854 );
or ( n65856 , n65741 , n65855 );
and ( n65857 , n65738 , n65856 );
or ( n65858 , n65737 , n65857 );
and ( n65859 , n65734 , n65858 );
or ( n65860 , n65733 , n65859 );
and ( n65861 , n65730 , n65860 );
or ( n65862 , n65729 , n65861 );
and ( n65863 , n65726 , n65862 );
or ( n65864 , n65725 , n65863 );
and ( n65865 , n65722 , n65864 );
or ( n65866 , n65721 , n65865 );
and ( n65867 , n65718 , n65866 );
or ( n65868 , n65717 , n65867 );
and ( n65869 , n65714 , n65868 );
or ( n65870 , n65713 , n65869 );
and ( n65871 , n65710 , n65870 );
or ( n65872 , n65709 , n65871 );
and ( n65873 , n65706 , n65872 );
or ( n65874 , n65705 , n65873 );
and ( n65875 , n65702 , n65874 );
or ( n65876 , n65701 , n65875 );
and ( n65877 , n65698 , n65876 );
or ( n65878 , n65697 , n65877 );
and ( n65879 , n65694 , n65878 );
or ( n65880 , n65693 , n65879 );
and ( n65881 , n65690 , n65880 );
or ( n65882 , n65689 , n65881 );
and ( n65883 , n65686 , n65882 );
or ( n65884 , n65685 , n65883 );
and ( n65885 , n65682 , n65884 );
or ( n65886 , n65681 , n65885 );
and ( n65887 , n65678 , n65886 );
or ( n65888 , n65677 , n65887 );
and ( n65889 , n65674 , n65888 );
or ( n65890 , n65673 , n65889 );
and ( n65891 , n65670 , n65890 );
or ( n65892 , n65669 , n65891 );
and ( n65893 , n65666 , n65892 );
or ( n65894 , n65665 , n65893 );
and ( n65895 , n65662 , n65894 );
or ( n65896 , n65661 , n65895 );
and ( n65897 , n65658 , n65896 );
or ( n65898 , n65657 , n65897 );
and ( n65899 , n65654 , n65898 );
or ( n65900 , n65653 , n65899 );
and ( n65901 , n65650 , n65900 );
or ( n65902 , n65649 , n65901 );
and ( n65903 , n65646 , n65902 );
or ( n65904 , n65645 , n65903 );
and ( n65905 , n65642 , n65904 );
or ( n65906 , n65641 , n65905 );
and ( n65907 , n65638 , n65906 );
or ( n65908 , n65637 , n65907 );
and ( n65909 , n65634 , n65908 );
or ( n65910 , n65633 , n65909 );
and ( n65911 , n65630 , n65910 );
or ( n65912 , n65629 , n65911 );
and ( n65913 , n65626 , n65912 );
or ( n65914 , n65625 , n65913 );
and ( n65915 , n65622 , n65914 );
or ( n65916 , n65621 , n65915 );
and ( n65917 , n65618 , n65916 );
or ( n65918 , n65617 , n65917 );
and ( n65919 , n65614 , n65918 );
or ( n65920 , n65613 , n65919 );
and ( n65921 , n65610 , n65920 );
or ( n65922 , n65609 , n65921 );
and ( n65923 , n65606 , n65922 );
or ( n65924 , n65605 , n65923 );
and ( n65925 , n65602 , n65924 );
or ( n65926 , n65601 , n65925 );
and ( n65927 , n65598 , n65926 );
or ( n65928 , n65597 , n65927 );
and ( n65929 , n65594 , n65928 );
or ( n65930 , n65593 , n65929 );
and ( n65931 , n65590 , n65930 );
or ( n65932 , n65589 , n65931 );
and ( n65933 , n65586 , n65932 );
or ( n65934 , n65585 , n65933 );
and ( n65935 , n65582 , n65934 );
or ( n65936 , n65581 , n65935 );
and ( n65937 , n65578 , n65936 );
or ( n65938 , n65577 , n65937 );
and ( n65939 , n65574 , n65938 );
or ( n65940 , n65573 , n65939 );
xor ( n65941 , n65570 , n65940 );
buf ( n65942 , n17976 );
and ( n65943 , n30104 , n65942 );
xor ( n65944 , n65941 , n65943 );
xor ( n65945 , n65574 , n65938 );
and ( n65946 , n30109 , n65942 );
and ( n65947 , n65945 , n65946 );
xor ( n65948 , n65945 , n65946 );
xor ( n65949 , n65578 , n65936 );
and ( n65950 , n30114 , n65942 );
and ( n65951 , n65949 , n65950 );
xor ( n65952 , n65949 , n65950 );
xor ( n65953 , n65582 , n65934 );
and ( n65954 , n30119 , n65942 );
and ( n65955 , n65953 , n65954 );
xor ( n65956 , n65953 , n65954 );
xor ( n65957 , n65586 , n65932 );
and ( n65958 , n30124 , n65942 );
and ( n65959 , n65957 , n65958 );
xor ( n65960 , n65957 , n65958 );
xor ( n65961 , n65590 , n65930 );
and ( n65962 , n30129 , n65942 );
and ( n65963 , n65961 , n65962 );
xor ( n65964 , n65961 , n65962 );
xor ( n65965 , n65594 , n65928 );
and ( n65966 , n30134 , n65942 );
and ( n65967 , n65965 , n65966 );
xor ( n65968 , n65965 , n65966 );
xor ( n65969 , n65598 , n65926 );
and ( n65970 , n30139 , n65942 );
and ( n65971 , n65969 , n65970 );
xor ( n65972 , n65969 , n65970 );
xor ( n65973 , n65602 , n65924 );
and ( n65974 , n30144 , n65942 );
and ( n65975 , n65973 , n65974 );
xor ( n65976 , n65973 , n65974 );
xor ( n65977 , n65606 , n65922 );
and ( n65978 , n30149 , n65942 );
and ( n65979 , n65977 , n65978 );
xor ( n65980 , n65977 , n65978 );
xor ( n65981 , n65610 , n65920 );
and ( n65982 , n30154 , n65942 );
and ( n65983 , n65981 , n65982 );
xor ( n65984 , n65981 , n65982 );
xor ( n65985 , n65614 , n65918 );
and ( n65986 , n30159 , n65942 );
and ( n65987 , n65985 , n65986 );
xor ( n65988 , n65985 , n65986 );
xor ( n65989 , n65618 , n65916 );
and ( n65990 , n30164 , n65942 );
and ( n65991 , n65989 , n65990 );
xor ( n65992 , n65989 , n65990 );
xor ( n65993 , n65622 , n65914 );
and ( n65994 , n30169 , n65942 );
and ( n65995 , n65993 , n65994 );
xor ( n65996 , n65993 , n65994 );
xor ( n65997 , n65626 , n65912 );
and ( n65998 , n30174 , n65942 );
and ( n65999 , n65997 , n65998 );
xor ( n66000 , n65997 , n65998 );
xor ( n66001 , n65630 , n65910 );
and ( n66002 , n30179 , n65942 );
and ( n66003 , n66001 , n66002 );
xor ( n66004 , n66001 , n66002 );
xor ( n66005 , n65634 , n65908 );
and ( n66006 , n30184 , n65942 );
and ( n66007 , n66005 , n66006 );
xor ( n66008 , n66005 , n66006 );
xor ( n66009 , n65638 , n65906 );
and ( n66010 , n30189 , n65942 );
and ( n66011 , n66009 , n66010 );
xor ( n66012 , n66009 , n66010 );
xor ( n66013 , n65642 , n65904 );
and ( n66014 , n30194 , n65942 );
and ( n66015 , n66013 , n66014 );
xor ( n66016 , n66013 , n66014 );
xor ( n66017 , n65646 , n65902 );
and ( n66018 , n30199 , n65942 );
and ( n66019 , n66017 , n66018 );
xor ( n66020 , n66017 , n66018 );
xor ( n66021 , n65650 , n65900 );
and ( n66022 , n30204 , n65942 );
and ( n66023 , n66021 , n66022 );
xor ( n66024 , n66021 , n66022 );
xor ( n66025 , n65654 , n65898 );
and ( n66026 , n30209 , n65942 );
and ( n66027 , n66025 , n66026 );
xor ( n66028 , n66025 , n66026 );
xor ( n66029 , n65658 , n65896 );
and ( n66030 , n30214 , n65942 );
and ( n66031 , n66029 , n66030 );
xor ( n66032 , n66029 , n66030 );
xor ( n66033 , n65662 , n65894 );
and ( n66034 , n30219 , n65942 );
and ( n66035 , n66033 , n66034 );
xor ( n66036 , n66033 , n66034 );
xor ( n66037 , n65666 , n65892 );
and ( n66038 , n30224 , n65942 );
and ( n66039 , n66037 , n66038 );
xor ( n66040 , n66037 , n66038 );
xor ( n66041 , n65670 , n65890 );
and ( n66042 , n30229 , n65942 );
and ( n66043 , n66041 , n66042 );
xor ( n66044 , n66041 , n66042 );
xor ( n66045 , n65674 , n65888 );
and ( n66046 , n30234 , n65942 );
and ( n66047 , n66045 , n66046 );
xor ( n66048 , n66045 , n66046 );
xor ( n66049 , n65678 , n65886 );
and ( n66050 , n30239 , n65942 );
and ( n66051 , n66049 , n66050 );
xor ( n66052 , n66049 , n66050 );
xor ( n66053 , n65682 , n65884 );
and ( n66054 , n30244 , n65942 );
and ( n66055 , n66053 , n66054 );
xor ( n66056 , n66053 , n66054 );
xor ( n66057 , n65686 , n65882 );
and ( n66058 , n30249 , n65942 );
and ( n66059 , n66057 , n66058 );
xor ( n66060 , n66057 , n66058 );
xor ( n66061 , n65690 , n65880 );
and ( n66062 , n30254 , n65942 );
and ( n66063 , n66061 , n66062 );
xor ( n66064 , n66061 , n66062 );
xor ( n66065 , n65694 , n65878 );
and ( n66066 , n30259 , n65942 );
and ( n66067 , n66065 , n66066 );
xor ( n66068 , n66065 , n66066 );
xor ( n66069 , n65698 , n65876 );
and ( n66070 , n30264 , n65942 );
and ( n66071 , n66069 , n66070 );
xor ( n66072 , n66069 , n66070 );
xor ( n66073 , n65702 , n65874 );
and ( n66074 , n30269 , n65942 );
and ( n66075 , n66073 , n66074 );
xor ( n66076 , n66073 , n66074 );
xor ( n66077 , n65706 , n65872 );
and ( n66078 , n30274 , n65942 );
and ( n66079 , n66077 , n66078 );
xor ( n66080 , n66077 , n66078 );
xor ( n66081 , n65710 , n65870 );
and ( n66082 , n30279 , n65942 );
and ( n66083 , n66081 , n66082 );
xor ( n66084 , n66081 , n66082 );
xor ( n66085 , n65714 , n65868 );
and ( n66086 , n30284 , n65942 );
and ( n66087 , n66085 , n66086 );
xor ( n66088 , n66085 , n66086 );
xor ( n66089 , n65718 , n65866 );
and ( n66090 , n30289 , n65942 );
and ( n66091 , n66089 , n66090 );
xor ( n66092 , n66089 , n66090 );
xor ( n66093 , n65722 , n65864 );
and ( n66094 , n30294 , n65942 );
and ( n66095 , n66093 , n66094 );
xor ( n66096 , n66093 , n66094 );
xor ( n66097 , n65726 , n65862 );
and ( n66098 , n30299 , n65942 );
and ( n66099 , n66097 , n66098 );
xor ( n66100 , n66097 , n66098 );
xor ( n66101 , n65730 , n65860 );
and ( n66102 , n30304 , n65942 );
and ( n66103 , n66101 , n66102 );
xor ( n66104 , n66101 , n66102 );
xor ( n66105 , n65734 , n65858 );
and ( n66106 , n30309 , n65942 );
and ( n66107 , n66105 , n66106 );
xor ( n66108 , n66105 , n66106 );
xor ( n66109 , n65738 , n65856 );
and ( n66110 , n30314 , n65942 );
and ( n66111 , n66109 , n66110 );
xor ( n66112 , n66109 , n66110 );
xor ( n66113 , n65742 , n65854 );
and ( n66114 , n30319 , n65942 );
and ( n66115 , n66113 , n66114 );
xor ( n66116 , n66113 , n66114 );
xor ( n66117 , n65746 , n65852 );
and ( n66118 , n30324 , n65942 );
and ( n66119 , n66117 , n66118 );
xor ( n66120 , n66117 , n66118 );
xor ( n66121 , n65750 , n65850 );
and ( n66122 , n30329 , n65942 );
and ( n66123 , n66121 , n66122 );
xor ( n66124 , n66121 , n66122 );
xor ( n66125 , n65754 , n65848 );
and ( n66126 , n30334 , n65942 );
and ( n66127 , n66125 , n66126 );
xor ( n66128 , n66125 , n66126 );
xor ( n66129 , n65758 , n65846 );
and ( n66130 , n30339 , n65942 );
and ( n66131 , n66129 , n66130 );
xor ( n66132 , n66129 , n66130 );
xor ( n66133 , n65762 , n65844 );
and ( n66134 , n30344 , n65942 );
and ( n66135 , n66133 , n66134 );
xor ( n66136 , n66133 , n66134 );
xor ( n66137 , n65766 , n65842 );
and ( n66138 , n30349 , n65942 );
and ( n66139 , n66137 , n66138 );
xor ( n66140 , n66137 , n66138 );
xor ( n66141 , n65770 , n65840 );
and ( n66142 , n30354 , n65942 );
and ( n66143 , n66141 , n66142 );
xor ( n66144 , n66141 , n66142 );
xor ( n66145 , n65774 , n65838 );
and ( n66146 , n30359 , n65942 );
and ( n66147 , n66145 , n66146 );
xor ( n66148 , n66145 , n66146 );
xor ( n66149 , n65778 , n65836 );
and ( n66150 , n30364 , n65942 );
and ( n66151 , n66149 , n66150 );
xor ( n66152 , n66149 , n66150 );
xor ( n66153 , n65782 , n65834 );
and ( n66154 , n30369 , n65942 );
and ( n66155 , n66153 , n66154 );
xor ( n66156 , n66153 , n66154 );
xor ( n66157 , n65786 , n65832 );
and ( n66158 , n30374 , n65942 );
and ( n66159 , n66157 , n66158 );
xor ( n66160 , n66157 , n66158 );
xor ( n66161 , n65790 , n65830 );
and ( n66162 , n30379 , n65942 );
and ( n66163 , n66161 , n66162 );
xor ( n66164 , n66161 , n66162 );
xor ( n66165 , n65794 , n65828 );
and ( n66166 , n30384 , n65942 );
and ( n66167 , n66165 , n66166 );
xor ( n66168 , n66165 , n66166 );
xor ( n66169 , n65798 , n65826 );
and ( n66170 , n30389 , n65942 );
and ( n66171 , n66169 , n66170 );
xor ( n66172 , n66169 , n66170 );
xor ( n66173 , n65802 , n65824 );
and ( n66174 , n30394 , n65942 );
and ( n66175 , n66173 , n66174 );
xor ( n66176 , n66173 , n66174 );
xor ( n66177 , n65806 , n65822 );
and ( n66178 , n30399 , n65942 );
and ( n66179 , n66177 , n66178 );
xor ( n66180 , n66177 , n66178 );
xor ( n66181 , n65810 , n65820 );
and ( n66182 , n30404 , n65942 );
and ( n66183 , n66181 , n66182 );
xor ( n66184 , n66181 , n66182 );
xor ( n66185 , n65814 , n65818 );
and ( n66186 , n30409 , n65942 );
and ( n66187 , n66185 , n66186 );
buf ( n66188 , n66187 );
and ( n66189 , n66184 , n66188 );
or ( n66190 , n66183 , n66189 );
and ( n66191 , n66180 , n66190 );
or ( n66192 , n66179 , n66191 );
and ( n66193 , n66176 , n66192 );
or ( n66194 , n66175 , n66193 );
and ( n66195 , n66172 , n66194 );
or ( n66196 , n66171 , n66195 );
and ( n66197 , n66168 , n66196 );
or ( n66198 , n66167 , n66197 );
and ( n66199 , n66164 , n66198 );
or ( n66200 , n66163 , n66199 );
and ( n66201 , n66160 , n66200 );
or ( n66202 , n66159 , n66201 );
and ( n66203 , n66156 , n66202 );
or ( n66204 , n66155 , n66203 );
and ( n66205 , n66152 , n66204 );
or ( n66206 , n66151 , n66205 );
and ( n66207 , n66148 , n66206 );
or ( n66208 , n66147 , n66207 );
and ( n66209 , n66144 , n66208 );
or ( n66210 , n66143 , n66209 );
and ( n66211 , n66140 , n66210 );
or ( n66212 , n66139 , n66211 );
and ( n66213 , n66136 , n66212 );
or ( n66214 , n66135 , n66213 );
and ( n66215 , n66132 , n66214 );
or ( n66216 , n66131 , n66215 );
and ( n66217 , n66128 , n66216 );
or ( n66218 , n66127 , n66217 );
and ( n66219 , n66124 , n66218 );
or ( n66220 , n66123 , n66219 );
and ( n66221 , n66120 , n66220 );
or ( n66222 , n66119 , n66221 );
and ( n66223 , n66116 , n66222 );
or ( n66224 , n66115 , n66223 );
and ( n66225 , n66112 , n66224 );
or ( n66226 , n66111 , n66225 );
and ( n66227 , n66108 , n66226 );
or ( n66228 , n66107 , n66227 );
and ( n66229 , n66104 , n66228 );
or ( n66230 , n66103 , n66229 );
and ( n66231 , n66100 , n66230 );
or ( n66232 , n66099 , n66231 );
and ( n66233 , n66096 , n66232 );
or ( n66234 , n66095 , n66233 );
and ( n66235 , n66092 , n66234 );
or ( n66236 , n66091 , n66235 );
and ( n66237 , n66088 , n66236 );
or ( n66238 , n66087 , n66237 );
and ( n66239 , n66084 , n66238 );
or ( n66240 , n66083 , n66239 );
and ( n66241 , n66080 , n66240 );
or ( n66242 , n66079 , n66241 );
and ( n66243 , n66076 , n66242 );
or ( n66244 , n66075 , n66243 );
and ( n66245 , n66072 , n66244 );
or ( n66246 , n66071 , n66245 );
and ( n66247 , n66068 , n66246 );
or ( n66248 , n66067 , n66247 );
and ( n66249 , n66064 , n66248 );
or ( n66250 , n66063 , n66249 );
and ( n66251 , n66060 , n66250 );
or ( n66252 , n66059 , n66251 );
and ( n66253 , n66056 , n66252 );
or ( n66254 , n66055 , n66253 );
and ( n66255 , n66052 , n66254 );
or ( n66256 , n66051 , n66255 );
and ( n66257 , n66048 , n66256 );
or ( n66258 , n66047 , n66257 );
and ( n66259 , n66044 , n66258 );
or ( n66260 , n66043 , n66259 );
and ( n66261 , n66040 , n66260 );
or ( n66262 , n66039 , n66261 );
and ( n66263 , n66036 , n66262 );
or ( n66264 , n66035 , n66263 );
and ( n66265 , n66032 , n66264 );
or ( n66266 , n66031 , n66265 );
and ( n66267 , n66028 , n66266 );
or ( n66268 , n66027 , n66267 );
and ( n66269 , n66024 , n66268 );
or ( n66270 , n66023 , n66269 );
and ( n66271 , n66020 , n66270 );
or ( n66272 , n66019 , n66271 );
and ( n66273 , n66016 , n66272 );
or ( n66274 , n66015 , n66273 );
and ( n66275 , n66012 , n66274 );
or ( n66276 , n66011 , n66275 );
and ( n66277 , n66008 , n66276 );
or ( n66278 , n66007 , n66277 );
and ( n66279 , n66004 , n66278 );
or ( n66280 , n66003 , n66279 );
and ( n66281 , n66000 , n66280 );
or ( n66282 , n65999 , n66281 );
and ( n66283 , n65996 , n66282 );
or ( n66284 , n65995 , n66283 );
and ( n66285 , n65992 , n66284 );
or ( n66286 , n65991 , n66285 );
and ( n66287 , n65988 , n66286 );
or ( n66288 , n65987 , n66287 );
and ( n66289 , n65984 , n66288 );
or ( n66290 , n65983 , n66289 );
and ( n66291 , n65980 , n66290 );
or ( n66292 , n65979 , n66291 );
and ( n66293 , n65976 , n66292 );
or ( n66294 , n65975 , n66293 );
and ( n66295 , n65972 , n66294 );
or ( n66296 , n65971 , n66295 );
and ( n66297 , n65968 , n66296 );
or ( n66298 , n65967 , n66297 );
and ( n66299 , n65964 , n66298 );
or ( n66300 , n65963 , n66299 );
and ( n66301 , n65960 , n66300 );
or ( n66302 , n65959 , n66301 );
and ( n66303 , n65956 , n66302 );
or ( n66304 , n65955 , n66303 );
and ( n66305 , n65952 , n66304 );
or ( n66306 , n65951 , n66305 );
and ( n66307 , n65948 , n66306 );
or ( n66308 , n65947 , n66307 );
xor ( n66309 , n65944 , n66308 );
buf ( n66310 , n17974 );
and ( n66311 , n30109 , n66310 );
xor ( n66312 , n66309 , n66311 );
xor ( n66313 , n65948 , n66306 );
and ( n66314 , n30114 , n66310 );
and ( n66315 , n66313 , n66314 );
xor ( n66316 , n66313 , n66314 );
xor ( n66317 , n65952 , n66304 );
and ( n66318 , n30119 , n66310 );
and ( n66319 , n66317 , n66318 );
xor ( n66320 , n66317 , n66318 );
xor ( n66321 , n65956 , n66302 );
and ( n66322 , n30124 , n66310 );
and ( n66323 , n66321 , n66322 );
xor ( n66324 , n66321 , n66322 );
xor ( n66325 , n65960 , n66300 );
and ( n66326 , n30129 , n66310 );
and ( n66327 , n66325 , n66326 );
xor ( n66328 , n66325 , n66326 );
xor ( n66329 , n65964 , n66298 );
and ( n66330 , n30134 , n66310 );
and ( n66331 , n66329 , n66330 );
xor ( n66332 , n66329 , n66330 );
xor ( n66333 , n65968 , n66296 );
and ( n66334 , n30139 , n66310 );
and ( n66335 , n66333 , n66334 );
xor ( n66336 , n66333 , n66334 );
xor ( n66337 , n65972 , n66294 );
and ( n66338 , n30144 , n66310 );
and ( n66339 , n66337 , n66338 );
xor ( n66340 , n66337 , n66338 );
xor ( n66341 , n65976 , n66292 );
and ( n66342 , n30149 , n66310 );
and ( n66343 , n66341 , n66342 );
xor ( n66344 , n66341 , n66342 );
xor ( n66345 , n65980 , n66290 );
and ( n66346 , n30154 , n66310 );
and ( n66347 , n66345 , n66346 );
xor ( n66348 , n66345 , n66346 );
xor ( n66349 , n65984 , n66288 );
and ( n66350 , n30159 , n66310 );
and ( n66351 , n66349 , n66350 );
xor ( n66352 , n66349 , n66350 );
xor ( n66353 , n65988 , n66286 );
and ( n66354 , n30164 , n66310 );
and ( n66355 , n66353 , n66354 );
xor ( n66356 , n66353 , n66354 );
xor ( n66357 , n65992 , n66284 );
and ( n66358 , n30169 , n66310 );
and ( n66359 , n66357 , n66358 );
xor ( n66360 , n66357 , n66358 );
xor ( n66361 , n65996 , n66282 );
and ( n66362 , n30174 , n66310 );
and ( n66363 , n66361 , n66362 );
xor ( n66364 , n66361 , n66362 );
xor ( n66365 , n66000 , n66280 );
and ( n66366 , n30179 , n66310 );
and ( n66367 , n66365 , n66366 );
xor ( n66368 , n66365 , n66366 );
xor ( n66369 , n66004 , n66278 );
and ( n66370 , n30184 , n66310 );
and ( n66371 , n66369 , n66370 );
xor ( n66372 , n66369 , n66370 );
xor ( n66373 , n66008 , n66276 );
and ( n66374 , n30189 , n66310 );
and ( n66375 , n66373 , n66374 );
xor ( n66376 , n66373 , n66374 );
xor ( n66377 , n66012 , n66274 );
and ( n66378 , n30194 , n66310 );
and ( n66379 , n66377 , n66378 );
xor ( n66380 , n66377 , n66378 );
xor ( n66381 , n66016 , n66272 );
and ( n66382 , n30199 , n66310 );
and ( n66383 , n66381 , n66382 );
xor ( n66384 , n66381 , n66382 );
xor ( n66385 , n66020 , n66270 );
and ( n66386 , n30204 , n66310 );
and ( n66387 , n66385 , n66386 );
xor ( n66388 , n66385 , n66386 );
xor ( n66389 , n66024 , n66268 );
and ( n66390 , n30209 , n66310 );
and ( n66391 , n66389 , n66390 );
xor ( n66392 , n66389 , n66390 );
xor ( n66393 , n66028 , n66266 );
and ( n66394 , n30214 , n66310 );
and ( n66395 , n66393 , n66394 );
xor ( n66396 , n66393 , n66394 );
xor ( n66397 , n66032 , n66264 );
and ( n66398 , n30219 , n66310 );
and ( n66399 , n66397 , n66398 );
xor ( n66400 , n66397 , n66398 );
xor ( n66401 , n66036 , n66262 );
and ( n66402 , n30224 , n66310 );
and ( n66403 , n66401 , n66402 );
xor ( n66404 , n66401 , n66402 );
xor ( n66405 , n66040 , n66260 );
and ( n66406 , n30229 , n66310 );
and ( n66407 , n66405 , n66406 );
xor ( n66408 , n66405 , n66406 );
xor ( n66409 , n66044 , n66258 );
and ( n66410 , n30234 , n66310 );
and ( n66411 , n66409 , n66410 );
xor ( n66412 , n66409 , n66410 );
xor ( n66413 , n66048 , n66256 );
and ( n66414 , n30239 , n66310 );
and ( n66415 , n66413 , n66414 );
xor ( n66416 , n66413 , n66414 );
xor ( n66417 , n66052 , n66254 );
and ( n66418 , n30244 , n66310 );
and ( n66419 , n66417 , n66418 );
xor ( n66420 , n66417 , n66418 );
xor ( n66421 , n66056 , n66252 );
and ( n66422 , n30249 , n66310 );
and ( n66423 , n66421 , n66422 );
xor ( n66424 , n66421 , n66422 );
xor ( n66425 , n66060 , n66250 );
and ( n66426 , n30254 , n66310 );
and ( n66427 , n66425 , n66426 );
xor ( n66428 , n66425 , n66426 );
xor ( n66429 , n66064 , n66248 );
and ( n66430 , n30259 , n66310 );
and ( n66431 , n66429 , n66430 );
xor ( n66432 , n66429 , n66430 );
xor ( n66433 , n66068 , n66246 );
and ( n66434 , n30264 , n66310 );
and ( n66435 , n66433 , n66434 );
xor ( n66436 , n66433 , n66434 );
xor ( n66437 , n66072 , n66244 );
and ( n66438 , n30269 , n66310 );
and ( n66439 , n66437 , n66438 );
xor ( n66440 , n66437 , n66438 );
xor ( n66441 , n66076 , n66242 );
and ( n66442 , n30274 , n66310 );
and ( n66443 , n66441 , n66442 );
xor ( n66444 , n66441 , n66442 );
xor ( n66445 , n66080 , n66240 );
and ( n66446 , n30279 , n66310 );
and ( n66447 , n66445 , n66446 );
xor ( n66448 , n66445 , n66446 );
xor ( n66449 , n66084 , n66238 );
and ( n66450 , n30284 , n66310 );
and ( n66451 , n66449 , n66450 );
xor ( n66452 , n66449 , n66450 );
xor ( n66453 , n66088 , n66236 );
and ( n66454 , n30289 , n66310 );
and ( n66455 , n66453 , n66454 );
xor ( n66456 , n66453 , n66454 );
xor ( n66457 , n66092 , n66234 );
and ( n66458 , n30294 , n66310 );
and ( n66459 , n66457 , n66458 );
xor ( n66460 , n66457 , n66458 );
xor ( n66461 , n66096 , n66232 );
and ( n66462 , n30299 , n66310 );
and ( n66463 , n66461 , n66462 );
xor ( n66464 , n66461 , n66462 );
xor ( n66465 , n66100 , n66230 );
and ( n66466 , n30304 , n66310 );
and ( n66467 , n66465 , n66466 );
xor ( n66468 , n66465 , n66466 );
xor ( n66469 , n66104 , n66228 );
and ( n66470 , n30309 , n66310 );
and ( n66471 , n66469 , n66470 );
xor ( n66472 , n66469 , n66470 );
xor ( n66473 , n66108 , n66226 );
and ( n66474 , n30314 , n66310 );
and ( n66475 , n66473 , n66474 );
xor ( n66476 , n66473 , n66474 );
xor ( n66477 , n66112 , n66224 );
and ( n66478 , n30319 , n66310 );
and ( n66479 , n66477 , n66478 );
xor ( n66480 , n66477 , n66478 );
xor ( n66481 , n66116 , n66222 );
and ( n66482 , n30324 , n66310 );
and ( n66483 , n66481 , n66482 );
xor ( n66484 , n66481 , n66482 );
xor ( n66485 , n66120 , n66220 );
and ( n66486 , n30329 , n66310 );
and ( n66487 , n66485 , n66486 );
xor ( n66488 , n66485 , n66486 );
xor ( n66489 , n66124 , n66218 );
and ( n66490 , n30334 , n66310 );
and ( n66491 , n66489 , n66490 );
xor ( n66492 , n66489 , n66490 );
xor ( n66493 , n66128 , n66216 );
and ( n66494 , n30339 , n66310 );
and ( n66495 , n66493 , n66494 );
xor ( n66496 , n66493 , n66494 );
xor ( n66497 , n66132 , n66214 );
and ( n66498 , n30344 , n66310 );
and ( n66499 , n66497 , n66498 );
xor ( n66500 , n66497 , n66498 );
xor ( n66501 , n66136 , n66212 );
and ( n66502 , n30349 , n66310 );
and ( n66503 , n66501 , n66502 );
xor ( n66504 , n66501 , n66502 );
xor ( n66505 , n66140 , n66210 );
and ( n66506 , n30354 , n66310 );
and ( n66507 , n66505 , n66506 );
xor ( n66508 , n66505 , n66506 );
xor ( n66509 , n66144 , n66208 );
and ( n66510 , n30359 , n66310 );
and ( n66511 , n66509 , n66510 );
xor ( n66512 , n66509 , n66510 );
xor ( n66513 , n66148 , n66206 );
and ( n66514 , n30364 , n66310 );
and ( n66515 , n66513 , n66514 );
xor ( n66516 , n66513 , n66514 );
xor ( n66517 , n66152 , n66204 );
and ( n66518 , n30369 , n66310 );
and ( n66519 , n66517 , n66518 );
xor ( n66520 , n66517 , n66518 );
xor ( n66521 , n66156 , n66202 );
and ( n66522 , n30374 , n66310 );
and ( n66523 , n66521 , n66522 );
xor ( n66524 , n66521 , n66522 );
xor ( n66525 , n66160 , n66200 );
and ( n66526 , n30379 , n66310 );
and ( n66527 , n66525 , n66526 );
xor ( n66528 , n66525 , n66526 );
xor ( n66529 , n66164 , n66198 );
and ( n66530 , n30384 , n66310 );
and ( n66531 , n66529 , n66530 );
xor ( n66532 , n66529 , n66530 );
xor ( n66533 , n66168 , n66196 );
and ( n66534 , n30389 , n66310 );
and ( n66535 , n66533 , n66534 );
xor ( n66536 , n66533 , n66534 );
xor ( n66537 , n66172 , n66194 );
and ( n66538 , n30394 , n66310 );
and ( n66539 , n66537 , n66538 );
xor ( n66540 , n66537 , n66538 );
xor ( n66541 , n66176 , n66192 );
and ( n66542 , n30399 , n66310 );
and ( n66543 , n66541 , n66542 );
xor ( n66544 , n66541 , n66542 );
xor ( n66545 , n66180 , n66190 );
and ( n66546 , n30404 , n66310 );
and ( n66547 , n66545 , n66546 );
xor ( n66548 , n66545 , n66546 );
xor ( n66549 , n66184 , n66188 );
and ( n66550 , n30409 , n66310 );
and ( n66551 , n66549 , n66550 );
buf ( n66552 , n66551 );
and ( n66553 , n66548 , n66552 );
or ( n66554 , n66547 , n66553 );
and ( n66555 , n66544 , n66554 );
or ( n66556 , n66543 , n66555 );
and ( n66557 , n66540 , n66556 );
or ( n66558 , n66539 , n66557 );
and ( n66559 , n66536 , n66558 );
or ( n66560 , n66535 , n66559 );
and ( n66561 , n66532 , n66560 );
or ( n66562 , n66531 , n66561 );
and ( n66563 , n66528 , n66562 );
or ( n66564 , n66527 , n66563 );
and ( n66565 , n66524 , n66564 );
or ( n66566 , n66523 , n66565 );
and ( n66567 , n66520 , n66566 );
or ( n66568 , n66519 , n66567 );
and ( n66569 , n66516 , n66568 );
or ( n66570 , n66515 , n66569 );
and ( n66571 , n66512 , n66570 );
or ( n66572 , n66511 , n66571 );
and ( n66573 , n66508 , n66572 );
or ( n66574 , n66507 , n66573 );
and ( n66575 , n66504 , n66574 );
or ( n66576 , n66503 , n66575 );
and ( n66577 , n66500 , n66576 );
or ( n66578 , n66499 , n66577 );
and ( n66579 , n66496 , n66578 );
or ( n66580 , n66495 , n66579 );
and ( n66581 , n66492 , n66580 );
or ( n66582 , n66491 , n66581 );
and ( n66583 , n66488 , n66582 );
or ( n66584 , n66487 , n66583 );
and ( n66585 , n66484 , n66584 );
or ( n66586 , n66483 , n66585 );
and ( n66587 , n66480 , n66586 );
or ( n66588 , n66479 , n66587 );
and ( n66589 , n66476 , n66588 );
or ( n66590 , n66475 , n66589 );
and ( n66591 , n66472 , n66590 );
or ( n66592 , n66471 , n66591 );
and ( n66593 , n66468 , n66592 );
or ( n66594 , n66467 , n66593 );
and ( n66595 , n66464 , n66594 );
or ( n66596 , n66463 , n66595 );
and ( n66597 , n66460 , n66596 );
or ( n66598 , n66459 , n66597 );
and ( n66599 , n66456 , n66598 );
or ( n66600 , n66455 , n66599 );
and ( n66601 , n66452 , n66600 );
or ( n66602 , n66451 , n66601 );
and ( n66603 , n66448 , n66602 );
or ( n66604 , n66447 , n66603 );
and ( n66605 , n66444 , n66604 );
or ( n66606 , n66443 , n66605 );
and ( n66607 , n66440 , n66606 );
or ( n66608 , n66439 , n66607 );
and ( n66609 , n66436 , n66608 );
or ( n66610 , n66435 , n66609 );
and ( n66611 , n66432 , n66610 );
or ( n66612 , n66431 , n66611 );
and ( n66613 , n66428 , n66612 );
or ( n66614 , n66427 , n66613 );
and ( n66615 , n66424 , n66614 );
or ( n66616 , n66423 , n66615 );
and ( n66617 , n66420 , n66616 );
or ( n66618 , n66419 , n66617 );
and ( n66619 , n66416 , n66618 );
or ( n66620 , n66415 , n66619 );
and ( n66621 , n66412 , n66620 );
or ( n66622 , n66411 , n66621 );
and ( n66623 , n66408 , n66622 );
or ( n66624 , n66407 , n66623 );
and ( n66625 , n66404 , n66624 );
or ( n66626 , n66403 , n66625 );
and ( n66627 , n66400 , n66626 );
or ( n66628 , n66399 , n66627 );
and ( n66629 , n66396 , n66628 );
or ( n66630 , n66395 , n66629 );
and ( n66631 , n66392 , n66630 );
or ( n66632 , n66391 , n66631 );
and ( n66633 , n66388 , n66632 );
or ( n66634 , n66387 , n66633 );
and ( n66635 , n66384 , n66634 );
or ( n66636 , n66383 , n66635 );
and ( n66637 , n66380 , n66636 );
or ( n66638 , n66379 , n66637 );
and ( n66639 , n66376 , n66638 );
or ( n66640 , n66375 , n66639 );
and ( n66641 , n66372 , n66640 );
or ( n66642 , n66371 , n66641 );
and ( n66643 , n66368 , n66642 );
or ( n66644 , n66367 , n66643 );
and ( n66645 , n66364 , n66644 );
or ( n66646 , n66363 , n66645 );
and ( n66647 , n66360 , n66646 );
or ( n66648 , n66359 , n66647 );
and ( n66649 , n66356 , n66648 );
or ( n66650 , n66355 , n66649 );
and ( n66651 , n66352 , n66650 );
or ( n66652 , n66351 , n66651 );
and ( n66653 , n66348 , n66652 );
or ( n66654 , n66347 , n66653 );
and ( n66655 , n66344 , n66654 );
or ( n66656 , n66343 , n66655 );
and ( n66657 , n66340 , n66656 );
or ( n66658 , n66339 , n66657 );
and ( n66659 , n66336 , n66658 );
or ( n66660 , n66335 , n66659 );
and ( n66661 , n66332 , n66660 );
or ( n66662 , n66331 , n66661 );
and ( n66663 , n66328 , n66662 );
or ( n66664 , n66327 , n66663 );
and ( n66665 , n66324 , n66664 );
or ( n66666 , n66323 , n66665 );
and ( n66667 , n66320 , n66666 );
or ( n66668 , n66319 , n66667 );
and ( n66669 , n66316 , n66668 );
or ( n66670 , n66315 , n66669 );
xor ( n66671 , n66312 , n66670 );
buf ( n66672 , n17972 );
and ( n66673 , n30114 , n66672 );
xor ( n66674 , n66671 , n66673 );
xor ( n66675 , n66316 , n66668 );
and ( n66676 , n30119 , n66672 );
and ( n66677 , n66675 , n66676 );
xor ( n66678 , n66675 , n66676 );
xor ( n66679 , n66320 , n66666 );
and ( n66680 , n30124 , n66672 );
and ( n66681 , n66679 , n66680 );
xor ( n66682 , n66679 , n66680 );
xor ( n66683 , n66324 , n66664 );
and ( n66684 , n30129 , n66672 );
and ( n66685 , n66683 , n66684 );
xor ( n66686 , n66683 , n66684 );
xor ( n66687 , n66328 , n66662 );
and ( n66688 , n30134 , n66672 );
and ( n66689 , n66687 , n66688 );
xor ( n66690 , n66687 , n66688 );
xor ( n66691 , n66332 , n66660 );
and ( n66692 , n30139 , n66672 );
and ( n66693 , n66691 , n66692 );
xor ( n66694 , n66691 , n66692 );
xor ( n66695 , n66336 , n66658 );
and ( n66696 , n30144 , n66672 );
and ( n66697 , n66695 , n66696 );
xor ( n66698 , n66695 , n66696 );
xor ( n66699 , n66340 , n66656 );
and ( n66700 , n30149 , n66672 );
and ( n66701 , n66699 , n66700 );
xor ( n66702 , n66699 , n66700 );
xor ( n66703 , n66344 , n66654 );
and ( n66704 , n30154 , n66672 );
and ( n66705 , n66703 , n66704 );
xor ( n66706 , n66703 , n66704 );
xor ( n66707 , n66348 , n66652 );
and ( n66708 , n30159 , n66672 );
and ( n66709 , n66707 , n66708 );
xor ( n66710 , n66707 , n66708 );
xor ( n66711 , n66352 , n66650 );
and ( n66712 , n30164 , n66672 );
and ( n66713 , n66711 , n66712 );
xor ( n66714 , n66711 , n66712 );
xor ( n66715 , n66356 , n66648 );
and ( n66716 , n30169 , n66672 );
and ( n66717 , n66715 , n66716 );
xor ( n66718 , n66715 , n66716 );
xor ( n66719 , n66360 , n66646 );
and ( n66720 , n30174 , n66672 );
and ( n66721 , n66719 , n66720 );
xor ( n66722 , n66719 , n66720 );
xor ( n66723 , n66364 , n66644 );
and ( n66724 , n30179 , n66672 );
and ( n66725 , n66723 , n66724 );
xor ( n66726 , n66723 , n66724 );
xor ( n66727 , n66368 , n66642 );
and ( n66728 , n30184 , n66672 );
and ( n66729 , n66727 , n66728 );
xor ( n66730 , n66727 , n66728 );
xor ( n66731 , n66372 , n66640 );
and ( n66732 , n30189 , n66672 );
and ( n66733 , n66731 , n66732 );
xor ( n66734 , n66731 , n66732 );
xor ( n66735 , n66376 , n66638 );
and ( n66736 , n30194 , n66672 );
and ( n66737 , n66735 , n66736 );
xor ( n66738 , n66735 , n66736 );
xor ( n66739 , n66380 , n66636 );
and ( n66740 , n30199 , n66672 );
and ( n66741 , n66739 , n66740 );
xor ( n66742 , n66739 , n66740 );
xor ( n66743 , n66384 , n66634 );
and ( n66744 , n30204 , n66672 );
and ( n66745 , n66743 , n66744 );
xor ( n66746 , n66743 , n66744 );
xor ( n66747 , n66388 , n66632 );
and ( n66748 , n30209 , n66672 );
and ( n66749 , n66747 , n66748 );
xor ( n66750 , n66747 , n66748 );
xor ( n66751 , n66392 , n66630 );
and ( n66752 , n30214 , n66672 );
and ( n66753 , n66751 , n66752 );
xor ( n66754 , n66751 , n66752 );
xor ( n66755 , n66396 , n66628 );
and ( n66756 , n30219 , n66672 );
and ( n66757 , n66755 , n66756 );
xor ( n66758 , n66755 , n66756 );
xor ( n66759 , n66400 , n66626 );
and ( n66760 , n30224 , n66672 );
and ( n66761 , n66759 , n66760 );
xor ( n66762 , n66759 , n66760 );
xor ( n66763 , n66404 , n66624 );
and ( n66764 , n30229 , n66672 );
and ( n66765 , n66763 , n66764 );
xor ( n66766 , n66763 , n66764 );
xor ( n66767 , n66408 , n66622 );
and ( n66768 , n30234 , n66672 );
and ( n66769 , n66767 , n66768 );
xor ( n66770 , n66767 , n66768 );
xor ( n66771 , n66412 , n66620 );
and ( n66772 , n30239 , n66672 );
and ( n66773 , n66771 , n66772 );
xor ( n66774 , n66771 , n66772 );
xor ( n66775 , n66416 , n66618 );
and ( n66776 , n30244 , n66672 );
and ( n66777 , n66775 , n66776 );
xor ( n66778 , n66775 , n66776 );
xor ( n66779 , n66420 , n66616 );
and ( n66780 , n30249 , n66672 );
and ( n66781 , n66779 , n66780 );
xor ( n66782 , n66779 , n66780 );
xor ( n66783 , n66424 , n66614 );
and ( n66784 , n30254 , n66672 );
and ( n66785 , n66783 , n66784 );
xor ( n66786 , n66783 , n66784 );
xor ( n66787 , n66428 , n66612 );
and ( n66788 , n30259 , n66672 );
and ( n66789 , n66787 , n66788 );
xor ( n66790 , n66787 , n66788 );
xor ( n66791 , n66432 , n66610 );
and ( n66792 , n30264 , n66672 );
and ( n66793 , n66791 , n66792 );
xor ( n66794 , n66791 , n66792 );
xor ( n66795 , n66436 , n66608 );
and ( n66796 , n30269 , n66672 );
and ( n66797 , n66795 , n66796 );
xor ( n66798 , n66795 , n66796 );
xor ( n66799 , n66440 , n66606 );
and ( n66800 , n30274 , n66672 );
and ( n66801 , n66799 , n66800 );
xor ( n66802 , n66799 , n66800 );
xor ( n66803 , n66444 , n66604 );
and ( n66804 , n30279 , n66672 );
and ( n66805 , n66803 , n66804 );
xor ( n66806 , n66803 , n66804 );
xor ( n66807 , n66448 , n66602 );
and ( n66808 , n30284 , n66672 );
and ( n66809 , n66807 , n66808 );
xor ( n66810 , n66807 , n66808 );
xor ( n66811 , n66452 , n66600 );
and ( n66812 , n30289 , n66672 );
and ( n66813 , n66811 , n66812 );
xor ( n66814 , n66811 , n66812 );
xor ( n66815 , n66456 , n66598 );
and ( n66816 , n30294 , n66672 );
and ( n66817 , n66815 , n66816 );
xor ( n66818 , n66815 , n66816 );
xor ( n66819 , n66460 , n66596 );
and ( n66820 , n30299 , n66672 );
and ( n66821 , n66819 , n66820 );
xor ( n66822 , n66819 , n66820 );
xor ( n66823 , n66464 , n66594 );
and ( n66824 , n30304 , n66672 );
and ( n66825 , n66823 , n66824 );
xor ( n66826 , n66823 , n66824 );
xor ( n66827 , n66468 , n66592 );
and ( n66828 , n30309 , n66672 );
and ( n66829 , n66827 , n66828 );
xor ( n66830 , n66827 , n66828 );
xor ( n66831 , n66472 , n66590 );
and ( n66832 , n30314 , n66672 );
and ( n66833 , n66831 , n66832 );
xor ( n66834 , n66831 , n66832 );
xor ( n66835 , n66476 , n66588 );
and ( n66836 , n30319 , n66672 );
and ( n66837 , n66835 , n66836 );
xor ( n66838 , n66835 , n66836 );
xor ( n66839 , n66480 , n66586 );
and ( n66840 , n30324 , n66672 );
and ( n66841 , n66839 , n66840 );
xor ( n66842 , n66839 , n66840 );
xor ( n66843 , n66484 , n66584 );
and ( n66844 , n30329 , n66672 );
and ( n66845 , n66843 , n66844 );
xor ( n66846 , n66843 , n66844 );
xor ( n66847 , n66488 , n66582 );
and ( n66848 , n30334 , n66672 );
and ( n66849 , n66847 , n66848 );
xor ( n66850 , n66847 , n66848 );
xor ( n66851 , n66492 , n66580 );
and ( n66852 , n30339 , n66672 );
and ( n66853 , n66851 , n66852 );
xor ( n66854 , n66851 , n66852 );
xor ( n66855 , n66496 , n66578 );
and ( n66856 , n30344 , n66672 );
and ( n66857 , n66855 , n66856 );
xor ( n66858 , n66855 , n66856 );
xor ( n66859 , n66500 , n66576 );
and ( n66860 , n30349 , n66672 );
and ( n66861 , n66859 , n66860 );
xor ( n66862 , n66859 , n66860 );
xor ( n66863 , n66504 , n66574 );
and ( n66864 , n30354 , n66672 );
and ( n66865 , n66863 , n66864 );
xor ( n66866 , n66863 , n66864 );
xor ( n66867 , n66508 , n66572 );
and ( n66868 , n30359 , n66672 );
and ( n66869 , n66867 , n66868 );
xor ( n66870 , n66867 , n66868 );
xor ( n66871 , n66512 , n66570 );
and ( n66872 , n30364 , n66672 );
and ( n66873 , n66871 , n66872 );
xor ( n66874 , n66871 , n66872 );
xor ( n66875 , n66516 , n66568 );
and ( n66876 , n30369 , n66672 );
and ( n66877 , n66875 , n66876 );
xor ( n66878 , n66875 , n66876 );
xor ( n66879 , n66520 , n66566 );
and ( n66880 , n30374 , n66672 );
and ( n66881 , n66879 , n66880 );
xor ( n66882 , n66879 , n66880 );
xor ( n66883 , n66524 , n66564 );
and ( n66884 , n30379 , n66672 );
and ( n66885 , n66883 , n66884 );
xor ( n66886 , n66883 , n66884 );
xor ( n66887 , n66528 , n66562 );
and ( n66888 , n30384 , n66672 );
and ( n66889 , n66887 , n66888 );
xor ( n66890 , n66887 , n66888 );
xor ( n66891 , n66532 , n66560 );
and ( n66892 , n30389 , n66672 );
and ( n66893 , n66891 , n66892 );
xor ( n66894 , n66891 , n66892 );
xor ( n66895 , n66536 , n66558 );
and ( n66896 , n30394 , n66672 );
and ( n66897 , n66895 , n66896 );
xor ( n66898 , n66895 , n66896 );
xor ( n66899 , n66540 , n66556 );
and ( n66900 , n30399 , n66672 );
and ( n66901 , n66899 , n66900 );
xor ( n66902 , n66899 , n66900 );
xor ( n66903 , n66544 , n66554 );
and ( n66904 , n30404 , n66672 );
and ( n66905 , n66903 , n66904 );
xor ( n66906 , n66903 , n66904 );
xor ( n66907 , n66548 , n66552 );
and ( n66908 , n30409 , n66672 );
and ( n66909 , n66907 , n66908 );
buf ( n66910 , n66909 );
and ( n66911 , n66906 , n66910 );
or ( n66912 , n66905 , n66911 );
and ( n66913 , n66902 , n66912 );
or ( n66914 , n66901 , n66913 );
and ( n66915 , n66898 , n66914 );
or ( n66916 , n66897 , n66915 );
and ( n66917 , n66894 , n66916 );
or ( n66918 , n66893 , n66917 );
and ( n66919 , n66890 , n66918 );
or ( n66920 , n66889 , n66919 );
and ( n66921 , n66886 , n66920 );
or ( n66922 , n66885 , n66921 );
and ( n66923 , n66882 , n66922 );
or ( n66924 , n66881 , n66923 );
and ( n66925 , n66878 , n66924 );
or ( n66926 , n66877 , n66925 );
and ( n66927 , n66874 , n66926 );
or ( n66928 , n66873 , n66927 );
and ( n66929 , n66870 , n66928 );
or ( n66930 , n66869 , n66929 );
and ( n66931 , n66866 , n66930 );
or ( n66932 , n66865 , n66931 );
and ( n66933 , n66862 , n66932 );
or ( n66934 , n66861 , n66933 );
and ( n66935 , n66858 , n66934 );
or ( n66936 , n66857 , n66935 );
and ( n66937 , n66854 , n66936 );
or ( n66938 , n66853 , n66937 );
and ( n66939 , n66850 , n66938 );
or ( n66940 , n66849 , n66939 );
and ( n66941 , n66846 , n66940 );
or ( n66942 , n66845 , n66941 );
and ( n66943 , n66842 , n66942 );
or ( n66944 , n66841 , n66943 );
and ( n66945 , n66838 , n66944 );
or ( n66946 , n66837 , n66945 );
and ( n66947 , n66834 , n66946 );
or ( n66948 , n66833 , n66947 );
and ( n66949 , n66830 , n66948 );
or ( n66950 , n66829 , n66949 );
and ( n66951 , n66826 , n66950 );
or ( n66952 , n66825 , n66951 );
and ( n66953 , n66822 , n66952 );
or ( n66954 , n66821 , n66953 );
and ( n66955 , n66818 , n66954 );
or ( n66956 , n66817 , n66955 );
and ( n66957 , n66814 , n66956 );
or ( n66958 , n66813 , n66957 );
and ( n66959 , n66810 , n66958 );
or ( n66960 , n66809 , n66959 );
and ( n66961 , n66806 , n66960 );
or ( n66962 , n66805 , n66961 );
and ( n66963 , n66802 , n66962 );
or ( n66964 , n66801 , n66963 );
and ( n66965 , n66798 , n66964 );
or ( n66966 , n66797 , n66965 );
and ( n66967 , n66794 , n66966 );
or ( n66968 , n66793 , n66967 );
and ( n66969 , n66790 , n66968 );
or ( n66970 , n66789 , n66969 );
and ( n66971 , n66786 , n66970 );
or ( n66972 , n66785 , n66971 );
and ( n66973 , n66782 , n66972 );
or ( n66974 , n66781 , n66973 );
and ( n66975 , n66778 , n66974 );
or ( n66976 , n66777 , n66975 );
and ( n66977 , n66774 , n66976 );
or ( n66978 , n66773 , n66977 );
and ( n66979 , n66770 , n66978 );
or ( n66980 , n66769 , n66979 );
and ( n66981 , n66766 , n66980 );
or ( n66982 , n66765 , n66981 );
and ( n66983 , n66762 , n66982 );
or ( n66984 , n66761 , n66983 );
and ( n66985 , n66758 , n66984 );
or ( n66986 , n66757 , n66985 );
and ( n66987 , n66754 , n66986 );
or ( n66988 , n66753 , n66987 );
and ( n66989 , n66750 , n66988 );
or ( n66990 , n66749 , n66989 );
and ( n66991 , n66746 , n66990 );
or ( n66992 , n66745 , n66991 );
and ( n66993 , n66742 , n66992 );
or ( n66994 , n66741 , n66993 );
and ( n66995 , n66738 , n66994 );
or ( n66996 , n66737 , n66995 );
and ( n66997 , n66734 , n66996 );
or ( n66998 , n66733 , n66997 );
and ( n66999 , n66730 , n66998 );
or ( n67000 , n66729 , n66999 );
and ( n67001 , n66726 , n67000 );
or ( n67002 , n66725 , n67001 );
and ( n67003 , n66722 , n67002 );
or ( n67004 , n66721 , n67003 );
and ( n67005 , n66718 , n67004 );
or ( n67006 , n66717 , n67005 );
and ( n67007 , n66714 , n67006 );
or ( n67008 , n66713 , n67007 );
and ( n67009 , n66710 , n67008 );
or ( n67010 , n66709 , n67009 );
and ( n67011 , n66706 , n67010 );
or ( n67012 , n66705 , n67011 );
and ( n67013 , n66702 , n67012 );
or ( n67014 , n66701 , n67013 );
and ( n67015 , n66698 , n67014 );
or ( n67016 , n66697 , n67015 );
and ( n67017 , n66694 , n67016 );
or ( n67018 , n66693 , n67017 );
and ( n67019 , n66690 , n67018 );
or ( n67020 , n66689 , n67019 );
and ( n67021 , n66686 , n67020 );
or ( n67022 , n66685 , n67021 );
and ( n67023 , n66682 , n67022 );
or ( n67024 , n66681 , n67023 );
and ( n67025 , n66678 , n67024 );
or ( n67026 , n66677 , n67025 );
xor ( n67027 , n66674 , n67026 );
buf ( n67028 , n17970 );
and ( n67029 , n30119 , n67028 );
xor ( n67030 , n67027 , n67029 );
xor ( n67031 , n66678 , n67024 );
and ( n67032 , n30124 , n67028 );
and ( n67033 , n67031 , n67032 );
xor ( n67034 , n67031 , n67032 );
xor ( n67035 , n66682 , n67022 );
and ( n67036 , n30129 , n67028 );
and ( n67037 , n67035 , n67036 );
xor ( n67038 , n67035 , n67036 );
xor ( n67039 , n66686 , n67020 );
and ( n67040 , n30134 , n67028 );
and ( n67041 , n67039 , n67040 );
xor ( n67042 , n67039 , n67040 );
xor ( n67043 , n66690 , n67018 );
and ( n67044 , n30139 , n67028 );
and ( n67045 , n67043 , n67044 );
xor ( n67046 , n67043 , n67044 );
xor ( n67047 , n66694 , n67016 );
and ( n67048 , n30144 , n67028 );
and ( n67049 , n67047 , n67048 );
xor ( n67050 , n67047 , n67048 );
xor ( n67051 , n66698 , n67014 );
and ( n67052 , n30149 , n67028 );
and ( n67053 , n67051 , n67052 );
xor ( n67054 , n67051 , n67052 );
xor ( n67055 , n66702 , n67012 );
and ( n67056 , n30154 , n67028 );
and ( n67057 , n67055 , n67056 );
xor ( n67058 , n67055 , n67056 );
xor ( n67059 , n66706 , n67010 );
and ( n67060 , n30159 , n67028 );
and ( n67061 , n67059 , n67060 );
xor ( n67062 , n67059 , n67060 );
xor ( n67063 , n66710 , n67008 );
and ( n67064 , n30164 , n67028 );
and ( n67065 , n67063 , n67064 );
xor ( n67066 , n67063 , n67064 );
xor ( n67067 , n66714 , n67006 );
and ( n67068 , n30169 , n67028 );
and ( n67069 , n67067 , n67068 );
xor ( n67070 , n67067 , n67068 );
xor ( n67071 , n66718 , n67004 );
and ( n67072 , n30174 , n67028 );
and ( n67073 , n67071 , n67072 );
xor ( n67074 , n67071 , n67072 );
xor ( n67075 , n66722 , n67002 );
and ( n67076 , n30179 , n67028 );
and ( n67077 , n67075 , n67076 );
xor ( n67078 , n67075 , n67076 );
xor ( n67079 , n66726 , n67000 );
and ( n67080 , n30184 , n67028 );
and ( n67081 , n67079 , n67080 );
xor ( n67082 , n67079 , n67080 );
xor ( n67083 , n66730 , n66998 );
and ( n67084 , n30189 , n67028 );
and ( n67085 , n67083 , n67084 );
xor ( n67086 , n67083 , n67084 );
xor ( n67087 , n66734 , n66996 );
and ( n67088 , n30194 , n67028 );
and ( n67089 , n67087 , n67088 );
xor ( n67090 , n67087 , n67088 );
xor ( n67091 , n66738 , n66994 );
and ( n67092 , n30199 , n67028 );
and ( n67093 , n67091 , n67092 );
xor ( n67094 , n67091 , n67092 );
xor ( n67095 , n66742 , n66992 );
and ( n67096 , n30204 , n67028 );
and ( n67097 , n67095 , n67096 );
xor ( n67098 , n67095 , n67096 );
xor ( n67099 , n66746 , n66990 );
and ( n67100 , n30209 , n67028 );
and ( n67101 , n67099 , n67100 );
xor ( n67102 , n67099 , n67100 );
xor ( n67103 , n66750 , n66988 );
and ( n67104 , n30214 , n67028 );
and ( n67105 , n67103 , n67104 );
xor ( n67106 , n67103 , n67104 );
xor ( n67107 , n66754 , n66986 );
and ( n67108 , n30219 , n67028 );
and ( n67109 , n67107 , n67108 );
xor ( n67110 , n67107 , n67108 );
xor ( n67111 , n66758 , n66984 );
and ( n67112 , n30224 , n67028 );
and ( n67113 , n67111 , n67112 );
xor ( n67114 , n67111 , n67112 );
xor ( n67115 , n66762 , n66982 );
and ( n67116 , n30229 , n67028 );
and ( n67117 , n67115 , n67116 );
xor ( n67118 , n67115 , n67116 );
xor ( n67119 , n66766 , n66980 );
and ( n67120 , n30234 , n67028 );
and ( n67121 , n67119 , n67120 );
xor ( n67122 , n67119 , n67120 );
xor ( n67123 , n66770 , n66978 );
and ( n67124 , n30239 , n67028 );
and ( n67125 , n67123 , n67124 );
xor ( n67126 , n67123 , n67124 );
xor ( n67127 , n66774 , n66976 );
and ( n67128 , n30244 , n67028 );
and ( n67129 , n67127 , n67128 );
xor ( n67130 , n67127 , n67128 );
xor ( n67131 , n66778 , n66974 );
and ( n67132 , n30249 , n67028 );
and ( n67133 , n67131 , n67132 );
xor ( n67134 , n67131 , n67132 );
xor ( n67135 , n66782 , n66972 );
and ( n67136 , n30254 , n67028 );
and ( n67137 , n67135 , n67136 );
xor ( n67138 , n67135 , n67136 );
xor ( n67139 , n66786 , n66970 );
and ( n67140 , n30259 , n67028 );
and ( n67141 , n67139 , n67140 );
xor ( n67142 , n67139 , n67140 );
xor ( n67143 , n66790 , n66968 );
and ( n67144 , n30264 , n67028 );
and ( n67145 , n67143 , n67144 );
xor ( n67146 , n67143 , n67144 );
xor ( n67147 , n66794 , n66966 );
and ( n67148 , n30269 , n67028 );
and ( n67149 , n67147 , n67148 );
xor ( n67150 , n67147 , n67148 );
xor ( n67151 , n66798 , n66964 );
and ( n67152 , n30274 , n67028 );
and ( n67153 , n67151 , n67152 );
xor ( n67154 , n67151 , n67152 );
xor ( n67155 , n66802 , n66962 );
and ( n67156 , n30279 , n67028 );
and ( n67157 , n67155 , n67156 );
xor ( n67158 , n67155 , n67156 );
xor ( n67159 , n66806 , n66960 );
and ( n67160 , n30284 , n67028 );
and ( n67161 , n67159 , n67160 );
xor ( n67162 , n67159 , n67160 );
xor ( n67163 , n66810 , n66958 );
and ( n67164 , n30289 , n67028 );
and ( n67165 , n67163 , n67164 );
xor ( n67166 , n67163 , n67164 );
xor ( n67167 , n66814 , n66956 );
and ( n67168 , n30294 , n67028 );
and ( n67169 , n67167 , n67168 );
xor ( n67170 , n67167 , n67168 );
xor ( n67171 , n66818 , n66954 );
and ( n67172 , n30299 , n67028 );
and ( n67173 , n67171 , n67172 );
xor ( n67174 , n67171 , n67172 );
xor ( n67175 , n66822 , n66952 );
and ( n67176 , n30304 , n67028 );
and ( n67177 , n67175 , n67176 );
xor ( n67178 , n67175 , n67176 );
xor ( n67179 , n66826 , n66950 );
and ( n67180 , n30309 , n67028 );
and ( n67181 , n67179 , n67180 );
xor ( n67182 , n67179 , n67180 );
xor ( n67183 , n66830 , n66948 );
and ( n67184 , n30314 , n67028 );
and ( n67185 , n67183 , n67184 );
xor ( n67186 , n67183 , n67184 );
xor ( n67187 , n66834 , n66946 );
and ( n67188 , n30319 , n67028 );
and ( n67189 , n67187 , n67188 );
xor ( n67190 , n67187 , n67188 );
xor ( n67191 , n66838 , n66944 );
and ( n67192 , n30324 , n67028 );
and ( n67193 , n67191 , n67192 );
xor ( n67194 , n67191 , n67192 );
xor ( n67195 , n66842 , n66942 );
and ( n67196 , n30329 , n67028 );
and ( n67197 , n67195 , n67196 );
xor ( n67198 , n67195 , n67196 );
xor ( n67199 , n66846 , n66940 );
and ( n67200 , n30334 , n67028 );
and ( n67201 , n67199 , n67200 );
xor ( n67202 , n67199 , n67200 );
xor ( n67203 , n66850 , n66938 );
and ( n67204 , n30339 , n67028 );
and ( n67205 , n67203 , n67204 );
xor ( n67206 , n67203 , n67204 );
xor ( n67207 , n66854 , n66936 );
and ( n67208 , n30344 , n67028 );
and ( n67209 , n67207 , n67208 );
xor ( n67210 , n67207 , n67208 );
xor ( n67211 , n66858 , n66934 );
and ( n67212 , n30349 , n67028 );
and ( n67213 , n67211 , n67212 );
xor ( n67214 , n67211 , n67212 );
xor ( n67215 , n66862 , n66932 );
and ( n67216 , n30354 , n67028 );
and ( n67217 , n67215 , n67216 );
xor ( n67218 , n67215 , n67216 );
xor ( n67219 , n66866 , n66930 );
and ( n67220 , n30359 , n67028 );
and ( n67221 , n67219 , n67220 );
xor ( n67222 , n67219 , n67220 );
xor ( n67223 , n66870 , n66928 );
and ( n67224 , n30364 , n67028 );
and ( n67225 , n67223 , n67224 );
xor ( n67226 , n67223 , n67224 );
xor ( n67227 , n66874 , n66926 );
and ( n67228 , n30369 , n67028 );
and ( n67229 , n67227 , n67228 );
xor ( n67230 , n67227 , n67228 );
xor ( n67231 , n66878 , n66924 );
and ( n67232 , n30374 , n67028 );
and ( n67233 , n67231 , n67232 );
xor ( n67234 , n67231 , n67232 );
xor ( n67235 , n66882 , n66922 );
and ( n67236 , n30379 , n67028 );
and ( n67237 , n67235 , n67236 );
xor ( n67238 , n67235 , n67236 );
xor ( n67239 , n66886 , n66920 );
and ( n67240 , n30384 , n67028 );
and ( n67241 , n67239 , n67240 );
xor ( n67242 , n67239 , n67240 );
xor ( n67243 , n66890 , n66918 );
and ( n67244 , n30389 , n67028 );
and ( n67245 , n67243 , n67244 );
xor ( n67246 , n67243 , n67244 );
xor ( n67247 , n66894 , n66916 );
and ( n67248 , n30394 , n67028 );
and ( n67249 , n67247 , n67248 );
xor ( n67250 , n67247 , n67248 );
xor ( n67251 , n66898 , n66914 );
and ( n67252 , n30399 , n67028 );
and ( n67253 , n67251 , n67252 );
xor ( n67254 , n67251 , n67252 );
xor ( n67255 , n66902 , n66912 );
and ( n67256 , n30404 , n67028 );
and ( n67257 , n67255 , n67256 );
xor ( n67258 , n67255 , n67256 );
xor ( n67259 , n66906 , n66910 );
and ( n67260 , n30409 , n67028 );
and ( n67261 , n67259 , n67260 );
buf ( n67262 , n67261 );
and ( n67263 , n67258 , n67262 );
or ( n67264 , n67257 , n67263 );
and ( n67265 , n67254 , n67264 );
or ( n67266 , n67253 , n67265 );
and ( n67267 , n67250 , n67266 );
or ( n67268 , n67249 , n67267 );
and ( n67269 , n67246 , n67268 );
or ( n67270 , n67245 , n67269 );
and ( n67271 , n67242 , n67270 );
or ( n67272 , n67241 , n67271 );
and ( n67273 , n67238 , n67272 );
or ( n67274 , n67237 , n67273 );
and ( n67275 , n67234 , n67274 );
or ( n67276 , n67233 , n67275 );
and ( n67277 , n67230 , n67276 );
or ( n67278 , n67229 , n67277 );
and ( n67279 , n67226 , n67278 );
or ( n67280 , n67225 , n67279 );
and ( n67281 , n67222 , n67280 );
or ( n67282 , n67221 , n67281 );
and ( n67283 , n67218 , n67282 );
or ( n67284 , n67217 , n67283 );
and ( n67285 , n67214 , n67284 );
or ( n67286 , n67213 , n67285 );
and ( n67287 , n67210 , n67286 );
or ( n67288 , n67209 , n67287 );
and ( n67289 , n67206 , n67288 );
or ( n67290 , n67205 , n67289 );
and ( n67291 , n67202 , n67290 );
or ( n67292 , n67201 , n67291 );
and ( n67293 , n67198 , n67292 );
or ( n67294 , n67197 , n67293 );
and ( n67295 , n67194 , n67294 );
or ( n67296 , n67193 , n67295 );
and ( n67297 , n67190 , n67296 );
or ( n67298 , n67189 , n67297 );
and ( n67299 , n67186 , n67298 );
or ( n67300 , n67185 , n67299 );
and ( n67301 , n67182 , n67300 );
or ( n67302 , n67181 , n67301 );
and ( n67303 , n67178 , n67302 );
or ( n67304 , n67177 , n67303 );
and ( n67305 , n67174 , n67304 );
or ( n67306 , n67173 , n67305 );
and ( n67307 , n67170 , n67306 );
or ( n67308 , n67169 , n67307 );
and ( n67309 , n67166 , n67308 );
or ( n67310 , n67165 , n67309 );
and ( n67311 , n67162 , n67310 );
or ( n67312 , n67161 , n67311 );
and ( n67313 , n67158 , n67312 );
or ( n67314 , n67157 , n67313 );
and ( n67315 , n67154 , n67314 );
or ( n67316 , n67153 , n67315 );
and ( n67317 , n67150 , n67316 );
or ( n67318 , n67149 , n67317 );
and ( n67319 , n67146 , n67318 );
or ( n67320 , n67145 , n67319 );
and ( n67321 , n67142 , n67320 );
or ( n67322 , n67141 , n67321 );
and ( n67323 , n67138 , n67322 );
or ( n67324 , n67137 , n67323 );
and ( n67325 , n67134 , n67324 );
or ( n67326 , n67133 , n67325 );
and ( n67327 , n67130 , n67326 );
or ( n67328 , n67129 , n67327 );
and ( n67329 , n67126 , n67328 );
or ( n67330 , n67125 , n67329 );
and ( n67331 , n67122 , n67330 );
or ( n67332 , n67121 , n67331 );
and ( n67333 , n67118 , n67332 );
or ( n67334 , n67117 , n67333 );
and ( n67335 , n67114 , n67334 );
or ( n67336 , n67113 , n67335 );
and ( n67337 , n67110 , n67336 );
or ( n67338 , n67109 , n67337 );
and ( n67339 , n67106 , n67338 );
or ( n67340 , n67105 , n67339 );
and ( n67341 , n67102 , n67340 );
or ( n67342 , n67101 , n67341 );
and ( n67343 , n67098 , n67342 );
or ( n67344 , n67097 , n67343 );
and ( n67345 , n67094 , n67344 );
or ( n67346 , n67093 , n67345 );
and ( n67347 , n67090 , n67346 );
or ( n67348 , n67089 , n67347 );
and ( n67349 , n67086 , n67348 );
or ( n67350 , n67085 , n67349 );
and ( n67351 , n67082 , n67350 );
or ( n67352 , n67081 , n67351 );
and ( n67353 , n67078 , n67352 );
or ( n67354 , n67077 , n67353 );
and ( n67355 , n67074 , n67354 );
or ( n67356 , n67073 , n67355 );
and ( n67357 , n67070 , n67356 );
or ( n67358 , n67069 , n67357 );
and ( n67359 , n67066 , n67358 );
or ( n67360 , n67065 , n67359 );
and ( n67361 , n67062 , n67360 );
or ( n67362 , n67061 , n67361 );
and ( n67363 , n67058 , n67362 );
or ( n67364 , n67057 , n67363 );
and ( n67365 , n67054 , n67364 );
or ( n67366 , n67053 , n67365 );
and ( n67367 , n67050 , n67366 );
or ( n67368 , n67049 , n67367 );
and ( n67369 , n67046 , n67368 );
or ( n67370 , n67045 , n67369 );
and ( n67371 , n67042 , n67370 );
or ( n67372 , n67041 , n67371 );
and ( n67373 , n67038 , n67372 );
or ( n67374 , n67037 , n67373 );
and ( n67375 , n67034 , n67374 );
or ( n67376 , n67033 , n67375 );
xor ( n67377 , n67030 , n67376 );
buf ( n67378 , n17968 );
and ( n67379 , n30124 , n67378 );
xor ( n67380 , n67377 , n67379 );
xor ( n67381 , n67034 , n67374 );
and ( n67382 , n30129 , n67378 );
and ( n67383 , n67381 , n67382 );
xor ( n67384 , n67381 , n67382 );
xor ( n67385 , n67038 , n67372 );
and ( n67386 , n30134 , n67378 );
and ( n67387 , n67385 , n67386 );
xor ( n67388 , n67385 , n67386 );
xor ( n67389 , n67042 , n67370 );
and ( n67390 , n30139 , n67378 );
and ( n67391 , n67389 , n67390 );
xor ( n67392 , n67389 , n67390 );
xor ( n67393 , n67046 , n67368 );
and ( n67394 , n30144 , n67378 );
and ( n67395 , n67393 , n67394 );
xor ( n67396 , n67393 , n67394 );
xor ( n67397 , n67050 , n67366 );
and ( n67398 , n30149 , n67378 );
and ( n67399 , n67397 , n67398 );
xor ( n67400 , n67397 , n67398 );
xor ( n67401 , n67054 , n67364 );
and ( n67402 , n30154 , n67378 );
and ( n67403 , n67401 , n67402 );
xor ( n67404 , n67401 , n67402 );
xor ( n67405 , n67058 , n67362 );
and ( n67406 , n30159 , n67378 );
and ( n67407 , n67405 , n67406 );
xor ( n67408 , n67405 , n67406 );
xor ( n67409 , n67062 , n67360 );
and ( n67410 , n30164 , n67378 );
and ( n67411 , n67409 , n67410 );
xor ( n67412 , n67409 , n67410 );
xor ( n67413 , n67066 , n67358 );
and ( n67414 , n30169 , n67378 );
and ( n67415 , n67413 , n67414 );
xor ( n67416 , n67413 , n67414 );
xor ( n67417 , n67070 , n67356 );
and ( n67418 , n30174 , n67378 );
and ( n67419 , n67417 , n67418 );
xor ( n67420 , n67417 , n67418 );
xor ( n67421 , n67074 , n67354 );
and ( n67422 , n30179 , n67378 );
and ( n67423 , n67421 , n67422 );
xor ( n67424 , n67421 , n67422 );
xor ( n67425 , n67078 , n67352 );
and ( n67426 , n30184 , n67378 );
and ( n67427 , n67425 , n67426 );
xor ( n67428 , n67425 , n67426 );
xor ( n67429 , n67082 , n67350 );
and ( n67430 , n30189 , n67378 );
and ( n67431 , n67429 , n67430 );
xor ( n67432 , n67429 , n67430 );
xor ( n67433 , n67086 , n67348 );
and ( n67434 , n30194 , n67378 );
and ( n67435 , n67433 , n67434 );
xor ( n67436 , n67433 , n67434 );
xor ( n67437 , n67090 , n67346 );
and ( n67438 , n30199 , n67378 );
and ( n67439 , n67437 , n67438 );
xor ( n67440 , n67437 , n67438 );
xor ( n67441 , n67094 , n67344 );
and ( n67442 , n30204 , n67378 );
and ( n67443 , n67441 , n67442 );
xor ( n67444 , n67441 , n67442 );
xor ( n67445 , n67098 , n67342 );
and ( n67446 , n30209 , n67378 );
and ( n67447 , n67445 , n67446 );
xor ( n67448 , n67445 , n67446 );
xor ( n67449 , n67102 , n67340 );
and ( n67450 , n30214 , n67378 );
and ( n67451 , n67449 , n67450 );
xor ( n67452 , n67449 , n67450 );
xor ( n67453 , n67106 , n67338 );
and ( n67454 , n30219 , n67378 );
and ( n67455 , n67453 , n67454 );
xor ( n67456 , n67453 , n67454 );
xor ( n67457 , n67110 , n67336 );
and ( n67458 , n30224 , n67378 );
and ( n67459 , n67457 , n67458 );
xor ( n67460 , n67457 , n67458 );
xor ( n67461 , n67114 , n67334 );
and ( n67462 , n30229 , n67378 );
and ( n67463 , n67461 , n67462 );
xor ( n67464 , n67461 , n67462 );
xor ( n67465 , n67118 , n67332 );
and ( n67466 , n30234 , n67378 );
and ( n67467 , n67465 , n67466 );
xor ( n67468 , n67465 , n67466 );
xor ( n67469 , n67122 , n67330 );
and ( n67470 , n30239 , n67378 );
and ( n67471 , n67469 , n67470 );
xor ( n67472 , n67469 , n67470 );
xor ( n67473 , n67126 , n67328 );
and ( n67474 , n30244 , n67378 );
and ( n67475 , n67473 , n67474 );
xor ( n67476 , n67473 , n67474 );
xor ( n67477 , n67130 , n67326 );
and ( n67478 , n30249 , n67378 );
and ( n67479 , n67477 , n67478 );
xor ( n67480 , n67477 , n67478 );
xor ( n67481 , n67134 , n67324 );
and ( n67482 , n30254 , n67378 );
and ( n67483 , n67481 , n67482 );
xor ( n67484 , n67481 , n67482 );
xor ( n67485 , n67138 , n67322 );
and ( n67486 , n30259 , n67378 );
and ( n67487 , n67485 , n67486 );
xor ( n67488 , n67485 , n67486 );
xor ( n67489 , n67142 , n67320 );
and ( n67490 , n30264 , n67378 );
and ( n67491 , n67489 , n67490 );
xor ( n67492 , n67489 , n67490 );
xor ( n67493 , n67146 , n67318 );
and ( n67494 , n30269 , n67378 );
and ( n67495 , n67493 , n67494 );
xor ( n67496 , n67493 , n67494 );
xor ( n67497 , n67150 , n67316 );
and ( n67498 , n30274 , n67378 );
and ( n67499 , n67497 , n67498 );
xor ( n67500 , n67497 , n67498 );
xor ( n67501 , n67154 , n67314 );
and ( n67502 , n30279 , n67378 );
and ( n67503 , n67501 , n67502 );
xor ( n67504 , n67501 , n67502 );
xor ( n67505 , n67158 , n67312 );
and ( n67506 , n30284 , n67378 );
and ( n67507 , n67505 , n67506 );
xor ( n67508 , n67505 , n67506 );
xor ( n67509 , n67162 , n67310 );
and ( n67510 , n30289 , n67378 );
and ( n67511 , n67509 , n67510 );
xor ( n67512 , n67509 , n67510 );
xor ( n67513 , n67166 , n67308 );
and ( n67514 , n30294 , n67378 );
and ( n67515 , n67513 , n67514 );
xor ( n67516 , n67513 , n67514 );
xor ( n67517 , n67170 , n67306 );
and ( n67518 , n30299 , n67378 );
and ( n67519 , n67517 , n67518 );
xor ( n67520 , n67517 , n67518 );
xor ( n67521 , n67174 , n67304 );
and ( n67522 , n30304 , n67378 );
and ( n67523 , n67521 , n67522 );
xor ( n67524 , n67521 , n67522 );
xor ( n67525 , n67178 , n67302 );
and ( n67526 , n30309 , n67378 );
and ( n67527 , n67525 , n67526 );
xor ( n67528 , n67525 , n67526 );
xor ( n67529 , n67182 , n67300 );
and ( n67530 , n30314 , n67378 );
and ( n67531 , n67529 , n67530 );
xor ( n67532 , n67529 , n67530 );
xor ( n67533 , n67186 , n67298 );
and ( n67534 , n30319 , n67378 );
and ( n67535 , n67533 , n67534 );
xor ( n67536 , n67533 , n67534 );
xor ( n67537 , n67190 , n67296 );
and ( n67538 , n30324 , n67378 );
and ( n67539 , n67537 , n67538 );
xor ( n67540 , n67537 , n67538 );
xor ( n67541 , n67194 , n67294 );
and ( n67542 , n30329 , n67378 );
and ( n67543 , n67541 , n67542 );
xor ( n67544 , n67541 , n67542 );
xor ( n67545 , n67198 , n67292 );
and ( n67546 , n30334 , n67378 );
and ( n67547 , n67545 , n67546 );
xor ( n67548 , n67545 , n67546 );
xor ( n67549 , n67202 , n67290 );
and ( n67550 , n30339 , n67378 );
and ( n67551 , n67549 , n67550 );
xor ( n67552 , n67549 , n67550 );
xor ( n67553 , n67206 , n67288 );
and ( n67554 , n30344 , n67378 );
and ( n67555 , n67553 , n67554 );
xor ( n67556 , n67553 , n67554 );
xor ( n67557 , n67210 , n67286 );
and ( n67558 , n30349 , n67378 );
and ( n67559 , n67557 , n67558 );
xor ( n67560 , n67557 , n67558 );
xor ( n67561 , n67214 , n67284 );
and ( n67562 , n30354 , n67378 );
and ( n67563 , n67561 , n67562 );
xor ( n67564 , n67561 , n67562 );
xor ( n67565 , n67218 , n67282 );
and ( n67566 , n30359 , n67378 );
and ( n67567 , n67565 , n67566 );
xor ( n67568 , n67565 , n67566 );
xor ( n67569 , n67222 , n67280 );
and ( n67570 , n30364 , n67378 );
and ( n67571 , n67569 , n67570 );
xor ( n67572 , n67569 , n67570 );
xor ( n67573 , n67226 , n67278 );
and ( n67574 , n30369 , n67378 );
and ( n67575 , n67573 , n67574 );
xor ( n67576 , n67573 , n67574 );
xor ( n67577 , n67230 , n67276 );
and ( n67578 , n30374 , n67378 );
and ( n67579 , n67577 , n67578 );
xor ( n67580 , n67577 , n67578 );
xor ( n67581 , n67234 , n67274 );
and ( n67582 , n30379 , n67378 );
and ( n67583 , n67581 , n67582 );
xor ( n67584 , n67581 , n67582 );
xor ( n67585 , n67238 , n67272 );
and ( n67586 , n30384 , n67378 );
and ( n67587 , n67585 , n67586 );
xor ( n67588 , n67585 , n67586 );
xor ( n67589 , n67242 , n67270 );
and ( n67590 , n30389 , n67378 );
and ( n67591 , n67589 , n67590 );
xor ( n67592 , n67589 , n67590 );
xor ( n67593 , n67246 , n67268 );
and ( n67594 , n30394 , n67378 );
and ( n67595 , n67593 , n67594 );
xor ( n67596 , n67593 , n67594 );
xor ( n67597 , n67250 , n67266 );
and ( n67598 , n30399 , n67378 );
and ( n67599 , n67597 , n67598 );
xor ( n67600 , n67597 , n67598 );
xor ( n67601 , n67254 , n67264 );
and ( n67602 , n30404 , n67378 );
and ( n67603 , n67601 , n67602 );
xor ( n67604 , n67601 , n67602 );
xor ( n67605 , n67258 , n67262 );
and ( n67606 , n30409 , n67378 );
and ( n67607 , n67605 , n67606 );
buf ( n67608 , n67607 );
and ( n67609 , n67604 , n67608 );
or ( n67610 , n67603 , n67609 );
and ( n67611 , n67600 , n67610 );
or ( n67612 , n67599 , n67611 );
and ( n67613 , n67596 , n67612 );
or ( n67614 , n67595 , n67613 );
and ( n67615 , n67592 , n67614 );
or ( n67616 , n67591 , n67615 );
and ( n67617 , n67588 , n67616 );
or ( n67618 , n67587 , n67617 );
and ( n67619 , n67584 , n67618 );
or ( n67620 , n67583 , n67619 );
and ( n67621 , n67580 , n67620 );
or ( n67622 , n67579 , n67621 );
and ( n67623 , n67576 , n67622 );
or ( n67624 , n67575 , n67623 );
and ( n67625 , n67572 , n67624 );
or ( n67626 , n67571 , n67625 );
and ( n67627 , n67568 , n67626 );
or ( n67628 , n67567 , n67627 );
and ( n67629 , n67564 , n67628 );
or ( n67630 , n67563 , n67629 );
and ( n67631 , n67560 , n67630 );
or ( n67632 , n67559 , n67631 );
and ( n67633 , n67556 , n67632 );
or ( n67634 , n67555 , n67633 );
and ( n67635 , n67552 , n67634 );
or ( n67636 , n67551 , n67635 );
and ( n67637 , n67548 , n67636 );
or ( n67638 , n67547 , n67637 );
and ( n67639 , n67544 , n67638 );
or ( n67640 , n67543 , n67639 );
and ( n67641 , n67540 , n67640 );
or ( n67642 , n67539 , n67641 );
and ( n67643 , n67536 , n67642 );
or ( n67644 , n67535 , n67643 );
and ( n67645 , n67532 , n67644 );
or ( n67646 , n67531 , n67645 );
and ( n67647 , n67528 , n67646 );
or ( n67648 , n67527 , n67647 );
and ( n67649 , n67524 , n67648 );
or ( n67650 , n67523 , n67649 );
and ( n67651 , n67520 , n67650 );
or ( n67652 , n67519 , n67651 );
and ( n67653 , n67516 , n67652 );
or ( n67654 , n67515 , n67653 );
and ( n67655 , n67512 , n67654 );
or ( n67656 , n67511 , n67655 );
and ( n67657 , n67508 , n67656 );
or ( n67658 , n67507 , n67657 );
and ( n67659 , n67504 , n67658 );
or ( n67660 , n67503 , n67659 );
and ( n67661 , n67500 , n67660 );
or ( n67662 , n67499 , n67661 );
and ( n67663 , n67496 , n67662 );
or ( n67664 , n67495 , n67663 );
and ( n67665 , n67492 , n67664 );
or ( n67666 , n67491 , n67665 );
and ( n67667 , n67488 , n67666 );
or ( n67668 , n67487 , n67667 );
and ( n67669 , n67484 , n67668 );
or ( n67670 , n67483 , n67669 );
and ( n67671 , n67480 , n67670 );
or ( n67672 , n67479 , n67671 );
and ( n67673 , n67476 , n67672 );
or ( n67674 , n67475 , n67673 );
and ( n67675 , n67472 , n67674 );
or ( n67676 , n67471 , n67675 );
and ( n67677 , n67468 , n67676 );
or ( n67678 , n67467 , n67677 );
and ( n67679 , n67464 , n67678 );
or ( n67680 , n67463 , n67679 );
and ( n67681 , n67460 , n67680 );
or ( n67682 , n67459 , n67681 );
and ( n67683 , n67456 , n67682 );
or ( n67684 , n67455 , n67683 );
and ( n67685 , n67452 , n67684 );
or ( n67686 , n67451 , n67685 );
and ( n67687 , n67448 , n67686 );
or ( n67688 , n67447 , n67687 );
and ( n67689 , n67444 , n67688 );
or ( n67690 , n67443 , n67689 );
and ( n67691 , n67440 , n67690 );
or ( n67692 , n67439 , n67691 );
and ( n67693 , n67436 , n67692 );
or ( n67694 , n67435 , n67693 );
and ( n67695 , n67432 , n67694 );
or ( n67696 , n67431 , n67695 );
and ( n67697 , n67428 , n67696 );
or ( n67698 , n67427 , n67697 );
and ( n67699 , n67424 , n67698 );
or ( n67700 , n67423 , n67699 );
and ( n67701 , n67420 , n67700 );
or ( n67702 , n67419 , n67701 );
and ( n67703 , n67416 , n67702 );
or ( n67704 , n67415 , n67703 );
and ( n67705 , n67412 , n67704 );
or ( n67706 , n67411 , n67705 );
and ( n67707 , n67408 , n67706 );
or ( n67708 , n67407 , n67707 );
and ( n67709 , n67404 , n67708 );
or ( n67710 , n67403 , n67709 );
and ( n67711 , n67400 , n67710 );
or ( n67712 , n67399 , n67711 );
and ( n67713 , n67396 , n67712 );
or ( n67714 , n67395 , n67713 );
and ( n67715 , n67392 , n67714 );
or ( n67716 , n67391 , n67715 );
and ( n67717 , n67388 , n67716 );
or ( n67718 , n67387 , n67717 );
and ( n67719 , n67384 , n67718 );
or ( n67720 , n67383 , n67719 );
xor ( n67721 , n67380 , n67720 );
buf ( n67722 , n17966 );
and ( n67723 , n30129 , n67722 );
xor ( n67724 , n67721 , n67723 );
xor ( n67725 , n67384 , n67718 );
and ( n67726 , n30134 , n67722 );
and ( n67727 , n67725 , n67726 );
xor ( n67728 , n67725 , n67726 );
xor ( n67729 , n67388 , n67716 );
and ( n67730 , n30139 , n67722 );
and ( n67731 , n67729 , n67730 );
xor ( n67732 , n67729 , n67730 );
xor ( n67733 , n67392 , n67714 );
and ( n67734 , n30144 , n67722 );
and ( n67735 , n67733 , n67734 );
xor ( n67736 , n67733 , n67734 );
xor ( n67737 , n67396 , n67712 );
and ( n67738 , n30149 , n67722 );
and ( n67739 , n67737 , n67738 );
xor ( n67740 , n67737 , n67738 );
xor ( n67741 , n67400 , n67710 );
and ( n67742 , n30154 , n67722 );
and ( n67743 , n67741 , n67742 );
xor ( n67744 , n67741 , n67742 );
xor ( n67745 , n67404 , n67708 );
and ( n67746 , n30159 , n67722 );
and ( n67747 , n67745 , n67746 );
xor ( n67748 , n67745 , n67746 );
xor ( n67749 , n67408 , n67706 );
and ( n67750 , n30164 , n67722 );
and ( n67751 , n67749 , n67750 );
xor ( n67752 , n67749 , n67750 );
xor ( n67753 , n67412 , n67704 );
and ( n67754 , n30169 , n67722 );
and ( n67755 , n67753 , n67754 );
xor ( n67756 , n67753 , n67754 );
xor ( n67757 , n67416 , n67702 );
and ( n67758 , n30174 , n67722 );
and ( n67759 , n67757 , n67758 );
xor ( n67760 , n67757 , n67758 );
xor ( n67761 , n67420 , n67700 );
and ( n67762 , n30179 , n67722 );
and ( n67763 , n67761 , n67762 );
xor ( n67764 , n67761 , n67762 );
xor ( n67765 , n67424 , n67698 );
and ( n67766 , n30184 , n67722 );
and ( n67767 , n67765 , n67766 );
xor ( n67768 , n67765 , n67766 );
xor ( n67769 , n67428 , n67696 );
and ( n67770 , n30189 , n67722 );
and ( n67771 , n67769 , n67770 );
xor ( n67772 , n67769 , n67770 );
xor ( n67773 , n67432 , n67694 );
and ( n67774 , n30194 , n67722 );
and ( n67775 , n67773 , n67774 );
xor ( n67776 , n67773 , n67774 );
xor ( n67777 , n67436 , n67692 );
and ( n67778 , n30199 , n67722 );
and ( n67779 , n67777 , n67778 );
xor ( n67780 , n67777 , n67778 );
xor ( n67781 , n67440 , n67690 );
and ( n67782 , n30204 , n67722 );
and ( n67783 , n67781 , n67782 );
xor ( n67784 , n67781 , n67782 );
xor ( n67785 , n67444 , n67688 );
and ( n67786 , n30209 , n67722 );
and ( n67787 , n67785 , n67786 );
xor ( n67788 , n67785 , n67786 );
xor ( n67789 , n67448 , n67686 );
and ( n67790 , n30214 , n67722 );
and ( n67791 , n67789 , n67790 );
xor ( n67792 , n67789 , n67790 );
xor ( n67793 , n67452 , n67684 );
and ( n67794 , n30219 , n67722 );
and ( n67795 , n67793 , n67794 );
xor ( n67796 , n67793 , n67794 );
xor ( n67797 , n67456 , n67682 );
and ( n67798 , n30224 , n67722 );
and ( n67799 , n67797 , n67798 );
xor ( n67800 , n67797 , n67798 );
xor ( n67801 , n67460 , n67680 );
and ( n67802 , n30229 , n67722 );
and ( n67803 , n67801 , n67802 );
xor ( n67804 , n67801 , n67802 );
xor ( n67805 , n67464 , n67678 );
and ( n67806 , n30234 , n67722 );
and ( n67807 , n67805 , n67806 );
xor ( n67808 , n67805 , n67806 );
xor ( n67809 , n67468 , n67676 );
and ( n67810 , n30239 , n67722 );
and ( n67811 , n67809 , n67810 );
xor ( n67812 , n67809 , n67810 );
xor ( n67813 , n67472 , n67674 );
and ( n67814 , n30244 , n67722 );
and ( n67815 , n67813 , n67814 );
xor ( n67816 , n67813 , n67814 );
xor ( n67817 , n67476 , n67672 );
and ( n67818 , n30249 , n67722 );
and ( n67819 , n67817 , n67818 );
xor ( n67820 , n67817 , n67818 );
xor ( n67821 , n67480 , n67670 );
and ( n67822 , n30254 , n67722 );
and ( n67823 , n67821 , n67822 );
xor ( n67824 , n67821 , n67822 );
xor ( n67825 , n67484 , n67668 );
and ( n67826 , n30259 , n67722 );
and ( n67827 , n67825 , n67826 );
xor ( n67828 , n67825 , n67826 );
xor ( n67829 , n67488 , n67666 );
and ( n67830 , n30264 , n67722 );
and ( n67831 , n67829 , n67830 );
xor ( n67832 , n67829 , n67830 );
xor ( n67833 , n67492 , n67664 );
and ( n67834 , n30269 , n67722 );
and ( n67835 , n67833 , n67834 );
xor ( n67836 , n67833 , n67834 );
xor ( n67837 , n67496 , n67662 );
and ( n67838 , n30274 , n67722 );
and ( n67839 , n67837 , n67838 );
xor ( n67840 , n67837 , n67838 );
xor ( n67841 , n67500 , n67660 );
and ( n67842 , n30279 , n67722 );
and ( n67843 , n67841 , n67842 );
xor ( n67844 , n67841 , n67842 );
xor ( n67845 , n67504 , n67658 );
and ( n67846 , n30284 , n67722 );
and ( n67847 , n67845 , n67846 );
xor ( n67848 , n67845 , n67846 );
xor ( n67849 , n67508 , n67656 );
and ( n67850 , n30289 , n67722 );
and ( n67851 , n67849 , n67850 );
xor ( n67852 , n67849 , n67850 );
xor ( n67853 , n67512 , n67654 );
and ( n67854 , n30294 , n67722 );
and ( n67855 , n67853 , n67854 );
xor ( n67856 , n67853 , n67854 );
xor ( n67857 , n67516 , n67652 );
and ( n67858 , n30299 , n67722 );
and ( n67859 , n67857 , n67858 );
xor ( n67860 , n67857 , n67858 );
xor ( n67861 , n67520 , n67650 );
and ( n67862 , n30304 , n67722 );
and ( n67863 , n67861 , n67862 );
xor ( n67864 , n67861 , n67862 );
xor ( n67865 , n67524 , n67648 );
and ( n67866 , n30309 , n67722 );
and ( n67867 , n67865 , n67866 );
xor ( n67868 , n67865 , n67866 );
xor ( n67869 , n67528 , n67646 );
and ( n67870 , n30314 , n67722 );
and ( n67871 , n67869 , n67870 );
xor ( n67872 , n67869 , n67870 );
xor ( n67873 , n67532 , n67644 );
and ( n67874 , n30319 , n67722 );
and ( n67875 , n67873 , n67874 );
xor ( n67876 , n67873 , n67874 );
xor ( n67877 , n67536 , n67642 );
and ( n67878 , n30324 , n67722 );
and ( n67879 , n67877 , n67878 );
xor ( n67880 , n67877 , n67878 );
xor ( n67881 , n67540 , n67640 );
and ( n67882 , n30329 , n67722 );
and ( n67883 , n67881 , n67882 );
xor ( n67884 , n67881 , n67882 );
xor ( n67885 , n67544 , n67638 );
and ( n67886 , n30334 , n67722 );
and ( n67887 , n67885 , n67886 );
xor ( n67888 , n67885 , n67886 );
xor ( n67889 , n67548 , n67636 );
and ( n67890 , n30339 , n67722 );
and ( n67891 , n67889 , n67890 );
xor ( n67892 , n67889 , n67890 );
xor ( n67893 , n67552 , n67634 );
and ( n67894 , n30344 , n67722 );
and ( n67895 , n67893 , n67894 );
xor ( n67896 , n67893 , n67894 );
xor ( n67897 , n67556 , n67632 );
and ( n67898 , n30349 , n67722 );
and ( n67899 , n67897 , n67898 );
xor ( n67900 , n67897 , n67898 );
xor ( n67901 , n67560 , n67630 );
and ( n67902 , n30354 , n67722 );
and ( n67903 , n67901 , n67902 );
xor ( n67904 , n67901 , n67902 );
xor ( n67905 , n67564 , n67628 );
and ( n67906 , n30359 , n67722 );
and ( n67907 , n67905 , n67906 );
xor ( n67908 , n67905 , n67906 );
xor ( n67909 , n67568 , n67626 );
and ( n67910 , n30364 , n67722 );
and ( n67911 , n67909 , n67910 );
xor ( n67912 , n67909 , n67910 );
xor ( n67913 , n67572 , n67624 );
and ( n67914 , n30369 , n67722 );
and ( n67915 , n67913 , n67914 );
xor ( n67916 , n67913 , n67914 );
xor ( n67917 , n67576 , n67622 );
and ( n67918 , n30374 , n67722 );
and ( n67919 , n67917 , n67918 );
xor ( n67920 , n67917 , n67918 );
xor ( n67921 , n67580 , n67620 );
and ( n67922 , n30379 , n67722 );
and ( n67923 , n67921 , n67922 );
xor ( n67924 , n67921 , n67922 );
xor ( n67925 , n67584 , n67618 );
and ( n67926 , n30384 , n67722 );
and ( n67927 , n67925 , n67926 );
xor ( n67928 , n67925 , n67926 );
xor ( n67929 , n67588 , n67616 );
and ( n67930 , n30389 , n67722 );
and ( n67931 , n67929 , n67930 );
xor ( n67932 , n67929 , n67930 );
xor ( n67933 , n67592 , n67614 );
and ( n67934 , n30394 , n67722 );
and ( n67935 , n67933 , n67934 );
xor ( n67936 , n67933 , n67934 );
xor ( n67937 , n67596 , n67612 );
and ( n67938 , n30399 , n67722 );
and ( n67939 , n67937 , n67938 );
xor ( n67940 , n67937 , n67938 );
xor ( n67941 , n67600 , n67610 );
and ( n67942 , n30404 , n67722 );
and ( n67943 , n67941 , n67942 );
xor ( n67944 , n67941 , n67942 );
xor ( n67945 , n67604 , n67608 );
and ( n67946 , n30409 , n67722 );
and ( n67947 , n67945 , n67946 );
buf ( n67948 , n67947 );
and ( n67949 , n67944 , n67948 );
or ( n67950 , n67943 , n67949 );
and ( n67951 , n67940 , n67950 );
or ( n67952 , n67939 , n67951 );
and ( n67953 , n67936 , n67952 );
or ( n67954 , n67935 , n67953 );
and ( n67955 , n67932 , n67954 );
or ( n67956 , n67931 , n67955 );
and ( n67957 , n67928 , n67956 );
or ( n67958 , n67927 , n67957 );
and ( n67959 , n67924 , n67958 );
or ( n67960 , n67923 , n67959 );
and ( n67961 , n67920 , n67960 );
or ( n67962 , n67919 , n67961 );
and ( n67963 , n67916 , n67962 );
or ( n67964 , n67915 , n67963 );
and ( n67965 , n67912 , n67964 );
or ( n67966 , n67911 , n67965 );
and ( n67967 , n67908 , n67966 );
or ( n67968 , n67907 , n67967 );
and ( n67969 , n67904 , n67968 );
or ( n67970 , n67903 , n67969 );
and ( n67971 , n67900 , n67970 );
or ( n67972 , n67899 , n67971 );
and ( n67973 , n67896 , n67972 );
or ( n67974 , n67895 , n67973 );
and ( n67975 , n67892 , n67974 );
or ( n67976 , n67891 , n67975 );
and ( n67977 , n67888 , n67976 );
or ( n67978 , n67887 , n67977 );
and ( n67979 , n67884 , n67978 );
or ( n67980 , n67883 , n67979 );
and ( n67981 , n67880 , n67980 );
or ( n67982 , n67879 , n67981 );
and ( n67983 , n67876 , n67982 );
or ( n67984 , n67875 , n67983 );
and ( n67985 , n67872 , n67984 );
or ( n67986 , n67871 , n67985 );
and ( n67987 , n67868 , n67986 );
or ( n67988 , n67867 , n67987 );
and ( n67989 , n67864 , n67988 );
or ( n67990 , n67863 , n67989 );
and ( n67991 , n67860 , n67990 );
or ( n67992 , n67859 , n67991 );
and ( n67993 , n67856 , n67992 );
or ( n67994 , n67855 , n67993 );
and ( n67995 , n67852 , n67994 );
or ( n67996 , n67851 , n67995 );
and ( n67997 , n67848 , n67996 );
or ( n67998 , n67847 , n67997 );
and ( n67999 , n67844 , n67998 );
or ( n68000 , n67843 , n67999 );
and ( n68001 , n67840 , n68000 );
or ( n68002 , n67839 , n68001 );
and ( n68003 , n67836 , n68002 );
or ( n68004 , n67835 , n68003 );
and ( n68005 , n67832 , n68004 );
or ( n68006 , n67831 , n68005 );
and ( n68007 , n67828 , n68006 );
or ( n68008 , n67827 , n68007 );
and ( n68009 , n67824 , n68008 );
or ( n68010 , n67823 , n68009 );
and ( n68011 , n67820 , n68010 );
or ( n68012 , n67819 , n68011 );
and ( n68013 , n67816 , n68012 );
or ( n68014 , n67815 , n68013 );
and ( n68015 , n67812 , n68014 );
or ( n68016 , n67811 , n68015 );
and ( n68017 , n67808 , n68016 );
or ( n68018 , n67807 , n68017 );
and ( n68019 , n67804 , n68018 );
or ( n68020 , n67803 , n68019 );
and ( n68021 , n67800 , n68020 );
or ( n68022 , n67799 , n68021 );
and ( n68023 , n67796 , n68022 );
or ( n68024 , n67795 , n68023 );
and ( n68025 , n67792 , n68024 );
or ( n68026 , n67791 , n68025 );
and ( n68027 , n67788 , n68026 );
or ( n68028 , n67787 , n68027 );
and ( n68029 , n67784 , n68028 );
or ( n68030 , n67783 , n68029 );
and ( n68031 , n67780 , n68030 );
or ( n68032 , n67779 , n68031 );
and ( n68033 , n67776 , n68032 );
or ( n68034 , n67775 , n68033 );
and ( n68035 , n67772 , n68034 );
or ( n68036 , n67771 , n68035 );
and ( n68037 , n67768 , n68036 );
or ( n68038 , n67767 , n68037 );
and ( n68039 , n67764 , n68038 );
or ( n68040 , n67763 , n68039 );
and ( n68041 , n67760 , n68040 );
or ( n68042 , n67759 , n68041 );
and ( n68043 , n67756 , n68042 );
or ( n68044 , n67755 , n68043 );
and ( n68045 , n67752 , n68044 );
or ( n68046 , n67751 , n68045 );
and ( n68047 , n67748 , n68046 );
or ( n68048 , n67747 , n68047 );
and ( n68049 , n67744 , n68048 );
or ( n68050 , n67743 , n68049 );
and ( n68051 , n67740 , n68050 );
or ( n68052 , n67739 , n68051 );
and ( n68053 , n67736 , n68052 );
or ( n68054 , n67735 , n68053 );
and ( n68055 , n67732 , n68054 );
or ( n68056 , n67731 , n68055 );
and ( n68057 , n67728 , n68056 );
or ( n68058 , n67727 , n68057 );
xor ( n68059 , n67724 , n68058 );
buf ( n68060 , n17964 );
and ( n68061 , n30134 , n68060 );
xor ( n68062 , n68059 , n68061 );
xor ( n68063 , n67728 , n68056 );
and ( n68064 , n30139 , n68060 );
and ( n68065 , n68063 , n68064 );
xor ( n68066 , n68063 , n68064 );
xor ( n68067 , n67732 , n68054 );
and ( n68068 , n30144 , n68060 );
and ( n68069 , n68067 , n68068 );
xor ( n68070 , n68067 , n68068 );
xor ( n68071 , n67736 , n68052 );
and ( n68072 , n30149 , n68060 );
and ( n68073 , n68071 , n68072 );
xor ( n68074 , n68071 , n68072 );
xor ( n68075 , n67740 , n68050 );
and ( n68076 , n30154 , n68060 );
and ( n68077 , n68075 , n68076 );
xor ( n68078 , n68075 , n68076 );
xor ( n68079 , n67744 , n68048 );
and ( n68080 , n30159 , n68060 );
and ( n68081 , n68079 , n68080 );
xor ( n68082 , n68079 , n68080 );
xor ( n68083 , n67748 , n68046 );
and ( n68084 , n30164 , n68060 );
and ( n68085 , n68083 , n68084 );
xor ( n68086 , n68083 , n68084 );
xor ( n68087 , n67752 , n68044 );
and ( n68088 , n30169 , n68060 );
and ( n68089 , n68087 , n68088 );
xor ( n68090 , n68087 , n68088 );
xor ( n68091 , n67756 , n68042 );
and ( n68092 , n30174 , n68060 );
and ( n68093 , n68091 , n68092 );
xor ( n68094 , n68091 , n68092 );
xor ( n68095 , n67760 , n68040 );
and ( n68096 , n30179 , n68060 );
and ( n68097 , n68095 , n68096 );
xor ( n68098 , n68095 , n68096 );
xor ( n68099 , n67764 , n68038 );
and ( n68100 , n30184 , n68060 );
and ( n68101 , n68099 , n68100 );
xor ( n68102 , n68099 , n68100 );
xor ( n68103 , n67768 , n68036 );
and ( n68104 , n30189 , n68060 );
and ( n68105 , n68103 , n68104 );
xor ( n68106 , n68103 , n68104 );
xor ( n68107 , n67772 , n68034 );
and ( n68108 , n30194 , n68060 );
and ( n68109 , n68107 , n68108 );
xor ( n68110 , n68107 , n68108 );
xor ( n68111 , n67776 , n68032 );
and ( n68112 , n30199 , n68060 );
and ( n68113 , n68111 , n68112 );
xor ( n68114 , n68111 , n68112 );
xor ( n68115 , n67780 , n68030 );
and ( n68116 , n30204 , n68060 );
and ( n68117 , n68115 , n68116 );
xor ( n68118 , n68115 , n68116 );
xor ( n68119 , n67784 , n68028 );
and ( n68120 , n30209 , n68060 );
and ( n68121 , n68119 , n68120 );
xor ( n68122 , n68119 , n68120 );
xor ( n68123 , n67788 , n68026 );
and ( n68124 , n30214 , n68060 );
and ( n68125 , n68123 , n68124 );
xor ( n68126 , n68123 , n68124 );
xor ( n68127 , n67792 , n68024 );
and ( n68128 , n30219 , n68060 );
and ( n68129 , n68127 , n68128 );
xor ( n68130 , n68127 , n68128 );
xor ( n68131 , n67796 , n68022 );
and ( n68132 , n30224 , n68060 );
and ( n68133 , n68131 , n68132 );
xor ( n68134 , n68131 , n68132 );
xor ( n68135 , n67800 , n68020 );
and ( n68136 , n30229 , n68060 );
and ( n68137 , n68135 , n68136 );
xor ( n68138 , n68135 , n68136 );
xor ( n68139 , n67804 , n68018 );
and ( n68140 , n30234 , n68060 );
and ( n68141 , n68139 , n68140 );
xor ( n68142 , n68139 , n68140 );
xor ( n68143 , n67808 , n68016 );
and ( n68144 , n30239 , n68060 );
and ( n68145 , n68143 , n68144 );
xor ( n68146 , n68143 , n68144 );
xor ( n68147 , n67812 , n68014 );
and ( n68148 , n30244 , n68060 );
and ( n68149 , n68147 , n68148 );
xor ( n68150 , n68147 , n68148 );
xor ( n68151 , n67816 , n68012 );
and ( n68152 , n30249 , n68060 );
and ( n68153 , n68151 , n68152 );
xor ( n68154 , n68151 , n68152 );
xor ( n68155 , n67820 , n68010 );
and ( n68156 , n30254 , n68060 );
and ( n68157 , n68155 , n68156 );
xor ( n68158 , n68155 , n68156 );
xor ( n68159 , n67824 , n68008 );
and ( n68160 , n30259 , n68060 );
and ( n68161 , n68159 , n68160 );
xor ( n68162 , n68159 , n68160 );
xor ( n68163 , n67828 , n68006 );
and ( n68164 , n30264 , n68060 );
and ( n68165 , n68163 , n68164 );
xor ( n68166 , n68163 , n68164 );
xor ( n68167 , n67832 , n68004 );
and ( n68168 , n30269 , n68060 );
and ( n68169 , n68167 , n68168 );
xor ( n68170 , n68167 , n68168 );
xor ( n68171 , n67836 , n68002 );
and ( n68172 , n30274 , n68060 );
and ( n68173 , n68171 , n68172 );
xor ( n68174 , n68171 , n68172 );
xor ( n68175 , n67840 , n68000 );
and ( n68176 , n30279 , n68060 );
and ( n68177 , n68175 , n68176 );
xor ( n68178 , n68175 , n68176 );
xor ( n68179 , n67844 , n67998 );
and ( n68180 , n30284 , n68060 );
and ( n68181 , n68179 , n68180 );
xor ( n68182 , n68179 , n68180 );
xor ( n68183 , n67848 , n67996 );
and ( n68184 , n30289 , n68060 );
and ( n68185 , n68183 , n68184 );
xor ( n68186 , n68183 , n68184 );
xor ( n68187 , n67852 , n67994 );
and ( n68188 , n30294 , n68060 );
and ( n68189 , n68187 , n68188 );
xor ( n68190 , n68187 , n68188 );
xor ( n68191 , n67856 , n67992 );
and ( n68192 , n30299 , n68060 );
and ( n68193 , n68191 , n68192 );
xor ( n68194 , n68191 , n68192 );
xor ( n68195 , n67860 , n67990 );
and ( n68196 , n30304 , n68060 );
and ( n68197 , n68195 , n68196 );
xor ( n68198 , n68195 , n68196 );
xor ( n68199 , n67864 , n67988 );
and ( n68200 , n30309 , n68060 );
and ( n68201 , n68199 , n68200 );
xor ( n68202 , n68199 , n68200 );
xor ( n68203 , n67868 , n67986 );
and ( n68204 , n30314 , n68060 );
and ( n68205 , n68203 , n68204 );
xor ( n68206 , n68203 , n68204 );
xor ( n68207 , n67872 , n67984 );
and ( n68208 , n30319 , n68060 );
and ( n68209 , n68207 , n68208 );
xor ( n68210 , n68207 , n68208 );
xor ( n68211 , n67876 , n67982 );
and ( n68212 , n30324 , n68060 );
and ( n68213 , n68211 , n68212 );
xor ( n68214 , n68211 , n68212 );
xor ( n68215 , n67880 , n67980 );
and ( n68216 , n30329 , n68060 );
and ( n68217 , n68215 , n68216 );
xor ( n68218 , n68215 , n68216 );
xor ( n68219 , n67884 , n67978 );
and ( n68220 , n30334 , n68060 );
and ( n68221 , n68219 , n68220 );
xor ( n68222 , n68219 , n68220 );
xor ( n68223 , n67888 , n67976 );
and ( n68224 , n30339 , n68060 );
and ( n68225 , n68223 , n68224 );
xor ( n68226 , n68223 , n68224 );
xor ( n68227 , n67892 , n67974 );
and ( n68228 , n30344 , n68060 );
and ( n68229 , n68227 , n68228 );
xor ( n68230 , n68227 , n68228 );
xor ( n68231 , n67896 , n67972 );
and ( n68232 , n30349 , n68060 );
and ( n68233 , n68231 , n68232 );
xor ( n68234 , n68231 , n68232 );
xor ( n68235 , n67900 , n67970 );
and ( n68236 , n30354 , n68060 );
and ( n68237 , n68235 , n68236 );
xor ( n68238 , n68235 , n68236 );
xor ( n68239 , n67904 , n67968 );
and ( n68240 , n30359 , n68060 );
and ( n68241 , n68239 , n68240 );
xor ( n68242 , n68239 , n68240 );
xor ( n68243 , n67908 , n67966 );
and ( n68244 , n30364 , n68060 );
and ( n68245 , n68243 , n68244 );
xor ( n68246 , n68243 , n68244 );
xor ( n68247 , n67912 , n67964 );
and ( n68248 , n30369 , n68060 );
and ( n68249 , n68247 , n68248 );
xor ( n68250 , n68247 , n68248 );
xor ( n68251 , n67916 , n67962 );
and ( n68252 , n30374 , n68060 );
and ( n68253 , n68251 , n68252 );
xor ( n68254 , n68251 , n68252 );
xor ( n68255 , n67920 , n67960 );
and ( n68256 , n30379 , n68060 );
and ( n68257 , n68255 , n68256 );
xor ( n68258 , n68255 , n68256 );
xor ( n68259 , n67924 , n67958 );
and ( n68260 , n30384 , n68060 );
and ( n68261 , n68259 , n68260 );
xor ( n68262 , n68259 , n68260 );
xor ( n68263 , n67928 , n67956 );
and ( n68264 , n30389 , n68060 );
and ( n68265 , n68263 , n68264 );
xor ( n68266 , n68263 , n68264 );
xor ( n68267 , n67932 , n67954 );
and ( n68268 , n30394 , n68060 );
and ( n68269 , n68267 , n68268 );
xor ( n68270 , n68267 , n68268 );
xor ( n68271 , n67936 , n67952 );
and ( n68272 , n30399 , n68060 );
and ( n68273 , n68271 , n68272 );
xor ( n68274 , n68271 , n68272 );
xor ( n68275 , n67940 , n67950 );
and ( n68276 , n30404 , n68060 );
and ( n68277 , n68275 , n68276 );
xor ( n68278 , n68275 , n68276 );
xor ( n68279 , n67944 , n67948 );
and ( n68280 , n30409 , n68060 );
and ( n68281 , n68279 , n68280 );
buf ( n68282 , n68281 );
and ( n68283 , n68278 , n68282 );
or ( n68284 , n68277 , n68283 );
and ( n68285 , n68274 , n68284 );
or ( n68286 , n68273 , n68285 );
and ( n68287 , n68270 , n68286 );
or ( n68288 , n68269 , n68287 );
and ( n68289 , n68266 , n68288 );
or ( n68290 , n68265 , n68289 );
and ( n68291 , n68262 , n68290 );
or ( n68292 , n68261 , n68291 );
and ( n68293 , n68258 , n68292 );
or ( n68294 , n68257 , n68293 );
and ( n68295 , n68254 , n68294 );
or ( n68296 , n68253 , n68295 );
and ( n68297 , n68250 , n68296 );
or ( n68298 , n68249 , n68297 );
and ( n68299 , n68246 , n68298 );
or ( n68300 , n68245 , n68299 );
and ( n68301 , n68242 , n68300 );
or ( n68302 , n68241 , n68301 );
and ( n68303 , n68238 , n68302 );
or ( n68304 , n68237 , n68303 );
and ( n68305 , n68234 , n68304 );
or ( n68306 , n68233 , n68305 );
and ( n68307 , n68230 , n68306 );
or ( n68308 , n68229 , n68307 );
and ( n68309 , n68226 , n68308 );
or ( n68310 , n68225 , n68309 );
and ( n68311 , n68222 , n68310 );
or ( n68312 , n68221 , n68311 );
and ( n68313 , n68218 , n68312 );
or ( n68314 , n68217 , n68313 );
and ( n68315 , n68214 , n68314 );
or ( n68316 , n68213 , n68315 );
and ( n68317 , n68210 , n68316 );
or ( n68318 , n68209 , n68317 );
and ( n68319 , n68206 , n68318 );
or ( n68320 , n68205 , n68319 );
and ( n68321 , n68202 , n68320 );
or ( n68322 , n68201 , n68321 );
and ( n68323 , n68198 , n68322 );
or ( n68324 , n68197 , n68323 );
and ( n68325 , n68194 , n68324 );
or ( n68326 , n68193 , n68325 );
and ( n68327 , n68190 , n68326 );
or ( n68328 , n68189 , n68327 );
and ( n68329 , n68186 , n68328 );
or ( n68330 , n68185 , n68329 );
and ( n68331 , n68182 , n68330 );
or ( n68332 , n68181 , n68331 );
and ( n68333 , n68178 , n68332 );
or ( n68334 , n68177 , n68333 );
and ( n68335 , n68174 , n68334 );
or ( n68336 , n68173 , n68335 );
and ( n68337 , n68170 , n68336 );
or ( n68338 , n68169 , n68337 );
and ( n68339 , n68166 , n68338 );
or ( n68340 , n68165 , n68339 );
and ( n68341 , n68162 , n68340 );
or ( n68342 , n68161 , n68341 );
and ( n68343 , n68158 , n68342 );
or ( n68344 , n68157 , n68343 );
and ( n68345 , n68154 , n68344 );
or ( n68346 , n68153 , n68345 );
and ( n68347 , n68150 , n68346 );
or ( n68348 , n68149 , n68347 );
and ( n68349 , n68146 , n68348 );
or ( n68350 , n68145 , n68349 );
and ( n68351 , n68142 , n68350 );
or ( n68352 , n68141 , n68351 );
and ( n68353 , n68138 , n68352 );
or ( n68354 , n68137 , n68353 );
and ( n68355 , n68134 , n68354 );
or ( n68356 , n68133 , n68355 );
and ( n68357 , n68130 , n68356 );
or ( n68358 , n68129 , n68357 );
and ( n68359 , n68126 , n68358 );
or ( n68360 , n68125 , n68359 );
and ( n68361 , n68122 , n68360 );
or ( n68362 , n68121 , n68361 );
and ( n68363 , n68118 , n68362 );
or ( n68364 , n68117 , n68363 );
and ( n68365 , n68114 , n68364 );
or ( n68366 , n68113 , n68365 );
and ( n68367 , n68110 , n68366 );
or ( n68368 , n68109 , n68367 );
and ( n68369 , n68106 , n68368 );
or ( n68370 , n68105 , n68369 );
and ( n68371 , n68102 , n68370 );
or ( n68372 , n68101 , n68371 );
and ( n68373 , n68098 , n68372 );
or ( n68374 , n68097 , n68373 );
and ( n68375 , n68094 , n68374 );
or ( n68376 , n68093 , n68375 );
and ( n68377 , n68090 , n68376 );
or ( n68378 , n68089 , n68377 );
and ( n68379 , n68086 , n68378 );
or ( n68380 , n68085 , n68379 );
and ( n68381 , n68082 , n68380 );
or ( n68382 , n68081 , n68381 );
and ( n68383 , n68078 , n68382 );
or ( n68384 , n68077 , n68383 );
and ( n68385 , n68074 , n68384 );
or ( n68386 , n68073 , n68385 );
and ( n68387 , n68070 , n68386 );
or ( n68388 , n68069 , n68387 );
and ( n68389 , n68066 , n68388 );
or ( n68390 , n68065 , n68389 );
xor ( n68391 , n68062 , n68390 );
buf ( n68392 , n17962 );
and ( n68393 , n30139 , n68392 );
xor ( n68394 , n68391 , n68393 );
xor ( n68395 , n68066 , n68388 );
and ( n68396 , n30144 , n68392 );
and ( n68397 , n68395 , n68396 );
xor ( n68398 , n68395 , n68396 );
xor ( n68399 , n68070 , n68386 );
and ( n68400 , n30149 , n68392 );
and ( n68401 , n68399 , n68400 );
xor ( n68402 , n68399 , n68400 );
xor ( n68403 , n68074 , n68384 );
and ( n68404 , n30154 , n68392 );
and ( n68405 , n68403 , n68404 );
xor ( n68406 , n68403 , n68404 );
xor ( n68407 , n68078 , n68382 );
and ( n68408 , n30159 , n68392 );
and ( n68409 , n68407 , n68408 );
xor ( n68410 , n68407 , n68408 );
xor ( n68411 , n68082 , n68380 );
and ( n68412 , n30164 , n68392 );
and ( n68413 , n68411 , n68412 );
xor ( n68414 , n68411 , n68412 );
xor ( n68415 , n68086 , n68378 );
and ( n68416 , n30169 , n68392 );
and ( n68417 , n68415 , n68416 );
xor ( n68418 , n68415 , n68416 );
xor ( n68419 , n68090 , n68376 );
and ( n68420 , n30174 , n68392 );
and ( n68421 , n68419 , n68420 );
xor ( n68422 , n68419 , n68420 );
xor ( n68423 , n68094 , n68374 );
and ( n68424 , n30179 , n68392 );
and ( n68425 , n68423 , n68424 );
xor ( n68426 , n68423 , n68424 );
xor ( n68427 , n68098 , n68372 );
and ( n68428 , n30184 , n68392 );
and ( n68429 , n68427 , n68428 );
xor ( n68430 , n68427 , n68428 );
xor ( n68431 , n68102 , n68370 );
and ( n68432 , n30189 , n68392 );
and ( n68433 , n68431 , n68432 );
xor ( n68434 , n68431 , n68432 );
xor ( n68435 , n68106 , n68368 );
and ( n68436 , n30194 , n68392 );
and ( n68437 , n68435 , n68436 );
xor ( n68438 , n68435 , n68436 );
xor ( n68439 , n68110 , n68366 );
and ( n68440 , n30199 , n68392 );
and ( n68441 , n68439 , n68440 );
xor ( n68442 , n68439 , n68440 );
xor ( n68443 , n68114 , n68364 );
and ( n68444 , n30204 , n68392 );
and ( n68445 , n68443 , n68444 );
xor ( n68446 , n68443 , n68444 );
xor ( n68447 , n68118 , n68362 );
and ( n68448 , n30209 , n68392 );
and ( n68449 , n68447 , n68448 );
xor ( n68450 , n68447 , n68448 );
xor ( n68451 , n68122 , n68360 );
and ( n68452 , n30214 , n68392 );
and ( n68453 , n68451 , n68452 );
xor ( n68454 , n68451 , n68452 );
xor ( n68455 , n68126 , n68358 );
and ( n68456 , n30219 , n68392 );
and ( n68457 , n68455 , n68456 );
xor ( n68458 , n68455 , n68456 );
xor ( n68459 , n68130 , n68356 );
and ( n68460 , n30224 , n68392 );
and ( n68461 , n68459 , n68460 );
xor ( n68462 , n68459 , n68460 );
xor ( n68463 , n68134 , n68354 );
and ( n68464 , n30229 , n68392 );
and ( n68465 , n68463 , n68464 );
xor ( n68466 , n68463 , n68464 );
xor ( n68467 , n68138 , n68352 );
and ( n68468 , n30234 , n68392 );
and ( n68469 , n68467 , n68468 );
xor ( n68470 , n68467 , n68468 );
xor ( n68471 , n68142 , n68350 );
and ( n68472 , n30239 , n68392 );
and ( n68473 , n68471 , n68472 );
xor ( n68474 , n68471 , n68472 );
xor ( n68475 , n68146 , n68348 );
and ( n68476 , n30244 , n68392 );
and ( n68477 , n68475 , n68476 );
xor ( n68478 , n68475 , n68476 );
xor ( n68479 , n68150 , n68346 );
and ( n68480 , n30249 , n68392 );
and ( n68481 , n68479 , n68480 );
xor ( n68482 , n68479 , n68480 );
xor ( n68483 , n68154 , n68344 );
and ( n68484 , n30254 , n68392 );
and ( n68485 , n68483 , n68484 );
xor ( n68486 , n68483 , n68484 );
xor ( n68487 , n68158 , n68342 );
and ( n68488 , n30259 , n68392 );
and ( n68489 , n68487 , n68488 );
xor ( n68490 , n68487 , n68488 );
xor ( n68491 , n68162 , n68340 );
and ( n68492 , n30264 , n68392 );
and ( n68493 , n68491 , n68492 );
xor ( n68494 , n68491 , n68492 );
xor ( n68495 , n68166 , n68338 );
and ( n68496 , n30269 , n68392 );
and ( n68497 , n68495 , n68496 );
xor ( n68498 , n68495 , n68496 );
xor ( n68499 , n68170 , n68336 );
and ( n68500 , n30274 , n68392 );
and ( n68501 , n68499 , n68500 );
xor ( n68502 , n68499 , n68500 );
xor ( n68503 , n68174 , n68334 );
and ( n68504 , n30279 , n68392 );
and ( n68505 , n68503 , n68504 );
xor ( n68506 , n68503 , n68504 );
xor ( n68507 , n68178 , n68332 );
and ( n68508 , n30284 , n68392 );
and ( n68509 , n68507 , n68508 );
xor ( n68510 , n68507 , n68508 );
xor ( n68511 , n68182 , n68330 );
and ( n68512 , n30289 , n68392 );
and ( n68513 , n68511 , n68512 );
xor ( n68514 , n68511 , n68512 );
xor ( n68515 , n68186 , n68328 );
and ( n68516 , n30294 , n68392 );
and ( n68517 , n68515 , n68516 );
xor ( n68518 , n68515 , n68516 );
xor ( n68519 , n68190 , n68326 );
and ( n68520 , n30299 , n68392 );
and ( n68521 , n68519 , n68520 );
xor ( n68522 , n68519 , n68520 );
xor ( n68523 , n68194 , n68324 );
and ( n68524 , n30304 , n68392 );
and ( n68525 , n68523 , n68524 );
xor ( n68526 , n68523 , n68524 );
xor ( n68527 , n68198 , n68322 );
and ( n68528 , n30309 , n68392 );
and ( n68529 , n68527 , n68528 );
xor ( n68530 , n68527 , n68528 );
xor ( n68531 , n68202 , n68320 );
and ( n68532 , n30314 , n68392 );
and ( n68533 , n68531 , n68532 );
xor ( n68534 , n68531 , n68532 );
xor ( n68535 , n68206 , n68318 );
and ( n68536 , n30319 , n68392 );
and ( n68537 , n68535 , n68536 );
xor ( n68538 , n68535 , n68536 );
xor ( n68539 , n68210 , n68316 );
and ( n68540 , n30324 , n68392 );
and ( n68541 , n68539 , n68540 );
xor ( n68542 , n68539 , n68540 );
xor ( n68543 , n68214 , n68314 );
and ( n68544 , n30329 , n68392 );
and ( n68545 , n68543 , n68544 );
xor ( n68546 , n68543 , n68544 );
xor ( n68547 , n68218 , n68312 );
and ( n68548 , n30334 , n68392 );
and ( n68549 , n68547 , n68548 );
xor ( n68550 , n68547 , n68548 );
xor ( n68551 , n68222 , n68310 );
and ( n68552 , n30339 , n68392 );
and ( n68553 , n68551 , n68552 );
xor ( n68554 , n68551 , n68552 );
xor ( n68555 , n68226 , n68308 );
and ( n68556 , n30344 , n68392 );
and ( n68557 , n68555 , n68556 );
xor ( n68558 , n68555 , n68556 );
xor ( n68559 , n68230 , n68306 );
and ( n68560 , n30349 , n68392 );
and ( n68561 , n68559 , n68560 );
xor ( n68562 , n68559 , n68560 );
xor ( n68563 , n68234 , n68304 );
and ( n68564 , n30354 , n68392 );
and ( n68565 , n68563 , n68564 );
xor ( n68566 , n68563 , n68564 );
xor ( n68567 , n68238 , n68302 );
and ( n68568 , n30359 , n68392 );
and ( n68569 , n68567 , n68568 );
xor ( n68570 , n68567 , n68568 );
xor ( n68571 , n68242 , n68300 );
and ( n68572 , n30364 , n68392 );
and ( n68573 , n68571 , n68572 );
xor ( n68574 , n68571 , n68572 );
xor ( n68575 , n68246 , n68298 );
and ( n68576 , n30369 , n68392 );
and ( n68577 , n68575 , n68576 );
xor ( n68578 , n68575 , n68576 );
xor ( n68579 , n68250 , n68296 );
and ( n68580 , n30374 , n68392 );
and ( n68581 , n68579 , n68580 );
xor ( n68582 , n68579 , n68580 );
xor ( n68583 , n68254 , n68294 );
and ( n68584 , n30379 , n68392 );
and ( n68585 , n68583 , n68584 );
xor ( n68586 , n68583 , n68584 );
xor ( n68587 , n68258 , n68292 );
and ( n68588 , n30384 , n68392 );
and ( n68589 , n68587 , n68588 );
xor ( n68590 , n68587 , n68588 );
xor ( n68591 , n68262 , n68290 );
and ( n68592 , n30389 , n68392 );
and ( n68593 , n68591 , n68592 );
xor ( n68594 , n68591 , n68592 );
xor ( n68595 , n68266 , n68288 );
and ( n68596 , n30394 , n68392 );
and ( n68597 , n68595 , n68596 );
xor ( n68598 , n68595 , n68596 );
xor ( n68599 , n68270 , n68286 );
and ( n68600 , n30399 , n68392 );
and ( n68601 , n68599 , n68600 );
xor ( n68602 , n68599 , n68600 );
xor ( n68603 , n68274 , n68284 );
and ( n68604 , n30404 , n68392 );
and ( n68605 , n68603 , n68604 );
xor ( n68606 , n68603 , n68604 );
xor ( n68607 , n68278 , n68282 );
and ( n68608 , n30409 , n68392 );
and ( n68609 , n68607 , n68608 );
buf ( n68610 , n68609 );
and ( n68611 , n68606 , n68610 );
or ( n68612 , n68605 , n68611 );
and ( n68613 , n68602 , n68612 );
or ( n68614 , n68601 , n68613 );
and ( n68615 , n68598 , n68614 );
or ( n68616 , n68597 , n68615 );
and ( n68617 , n68594 , n68616 );
or ( n68618 , n68593 , n68617 );
and ( n68619 , n68590 , n68618 );
or ( n68620 , n68589 , n68619 );
and ( n68621 , n68586 , n68620 );
or ( n68622 , n68585 , n68621 );
and ( n68623 , n68582 , n68622 );
or ( n68624 , n68581 , n68623 );
and ( n68625 , n68578 , n68624 );
or ( n68626 , n68577 , n68625 );
and ( n68627 , n68574 , n68626 );
or ( n68628 , n68573 , n68627 );
and ( n68629 , n68570 , n68628 );
or ( n68630 , n68569 , n68629 );
and ( n68631 , n68566 , n68630 );
or ( n68632 , n68565 , n68631 );
and ( n68633 , n68562 , n68632 );
or ( n68634 , n68561 , n68633 );
and ( n68635 , n68558 , n68634 );
or ( n68636 , n68557 , n68635 );
and ( n68637 , n68554 , n68636 );
or ( n68638 , n68553 , n68637 );
and ( n68639 , n68550 , n68638 );
or ( n68640 , n68549 , n68639 );
and ( n68641 , n68546 , n68640 );
or ( n68642 , n68545 , n68641 );
and ( n68643 , n68542 , n68642 );
or ( n68644 , n68541 , n68643 );
and ( n68645 , n68538 , n68644 );
or ( n68646 , n68537 , n68645 );
and ( n68647 , n68534 , n68646 );
or ( n68648 , n68533 , n68647 );
and ( n68649 , n68530 , n68648 );
or ( n68650 , n68529 , n68649 );
and ( n68651 , n68526 , n68650 );
or ( n68652 , n68525 , n68651 );
and ( n68653 , n68522 , n68652 );
or ( n68654 , n68521 , n68653 );
and ( n68655 , n68518 , n68654 );
or ( n68656 , n68517 , n68655 );
and ( n68657 , n68514 , n68656 );
or ( n68658 , n68513 , n68657 );
and ( n68659 , n68510 , n68658 );
or ( n68660 , n68509 , n68659 );
and ( n68661 , n68506 , n68660 );
or ( n68662 , n68505 , n68661 );
and ( n68663 , n68502 , n68662 );
or ( n68664 , n68501 , n68663 );
and ( n68665 , n68498 , n68664 );
or ( n68666 , n68497 , n68665 );
and ( n68667 , n68494 , n68666 );
or ( n68668 , n68493 , n68667 );
and ( n68669 , n68490 , n68668 );
or ( n68670 , n68489 , n68669 );
and ( n68671 , n68486 , n68670 );
or ( n68672 , n68485 , n68671 );
and ( n68673 , n68482 , n68672 );
or ( n68674 , n68481 , n68673 );
and ( n68675 , n68478 , n68674 );
or ( n68676 , n68477 , n68675 );
and ( n68677 , n68474 , n68676 );
or ( n68678 , n68473 , n68677 );
and ( n68679 , n68470 , n68678 );
or ( n68680 , n68469 , n68679 );
and ( n68681 , n68466 , n68680 );
or ( n68682 , n68465 , n68681 );
and ( n68683 , n68462 , n68682 );
or ( n68684 , n68461 , n68683 );
and ( n68685 , n68458 , n68684 );
or ( n68686 , n68457 , n68685 );
and ( n68687 , n68454 , n68686 );
or ( n68688 , n68453 , n68687 );
and ( n68689 , n68450 , n68688 );
or ( n68690 , n68449 , n68689 );
and ( n68691 , n68446 , n68690 );
or ( n68692 , n68445 , n68691 );
and ( n68693 , n68442 , n68692 );
or ( n68694 , n68441 , n68693 );
and ( n68695 , n68438 , n68694 );
or ( n68696 , n68437 , n68695 );
and ( n68697 , n68434 , n68696 );
or ( n68698 , n68433 , n68697 );
and ( n68699 , n68430 , n68698 );
or ( n68700 , n68429 , n68699 );
and ( n68701 , n68426 , n68700 );
or ( n68702 , n68425 , n68701 );
and ( n68703 , n68422 , n68702 );
or ( n68704 , n68421 , n68703 );
and ( n68705 , n68418 , n68704 );
or ( n68706 , n68417 , n68705 );
and ( n68707 , n68414 , n68706 );
or ( n68708 , n68413 , n68707 );
and ( n68709 , n68410 , n68708 );
or ( n68710 , n68409 , n68709 );
and ( n68711 , n68406 , n68710 );
or ( n68712 , n68405 , n68711 );
and ( n68713 , n68402 , n68712 );
or ( n68714 , n68401 , n68713 );
and ( n68715 , n68398 , n68714 );
or ( n68716 , n68397 , n68715 );
xor ( n68717 , n68394 , n68716 );
buf ( n68718 , n17960 );
and ( n68719 , n30144 , n68718 );
xor ( n68720 , n68717 , n68719 );
xor ( n68721 , n68398 , n68714 );
and ( n68722 , n30149 , n68718 );
and ( n68723 , n68721 , n68722 );
xor ( n68724 , n68721 , n68722 );
xor ( n68725 , n68402 , n68712 );
and ( n68726 , n30154 , n68718 );
and ( n68727 , n68725 , n68726 );
xor ( n68728 , n68725 , n68726 );
xor ( n68729 , n68406 , n68710 );
and ( n68730 , n30159 , n68718 );
and ( n68731 , n68729 , n68730 );
xor ( n68732 , n68729 , n68730 );
xor ( n68733 , n68410 , n68708 );
and ( n68734 , n30164 , n68718 );
and ( n68735 , n68733 , n68734 );
xor ( n68736 , n68733 , n68734 );
xor ( n68737 , n68414 , n68706 );
and ( n68738 , n30169 , n68718 );
and ( n68739 , n68737 , n68738 );
xor ( n68740 , n68737 , n68738 );
xor ( n68741 , n68418 , n68704 );
and ( n68742 , n30174 , n68718 );
and ( n68743 , n68741 , n68742 );
xor ( n68744 , n68741 , n68742 );
xor ( n68745 , n68422 , n68702 );
and ( n68746 , n30179 , n68718 );
and ( n68747 , n68745 , n68746 );
xor ( n68748 , n68745 , n68746 );
xor ( n68749 , n68426 , n68700 );
and ( n68750 , n30184 , n68718 );
and ( n68751 , n68749 , n68750 );
xor ( n68752 , n68749 , n68750 );
xor ( n68753 , n68430 , n68698 );
and ( n68754 , n30189 , n68718 );
and ( n68755 , n68753 , n68754 );
xor ( n68756 , n68753 , n68754 );
xor ( n68757 , n68434 , n68696 );
and ( n68758 , n30194 , n68718 );
and ( n68759 , n68757 , n68758 );
xor ( n68760 , n68757 , n68758 );
xor ( n68761 , n68438 , n68694 );
and ( n68762 , n30199 , n68718 );
and ( n68763 , n68761 , n68762 );
xor ( n68764 , n68761 , n68762 );
xor ( n68765 , n68442 , n68692 );
and ( n68766 , n30204 , n68718 );
and ( n68767 , n68765 , n68766 );
xor ( n68768 , n68765 , n68766 );
xor ( n68769 , n68446 , n68690 );
and ( n68770 , n30209 , n68718 );
and ( n68771 , n68769 , n68770 );
xor ( n68772 , n68769 , n68770 );
xor ( n68773 , n68450 , n68688 );
and ( n68774 , n30214 , n68718 );
and ( n68775 , n68773 , n68774 );
xor ( n68776 , n68773 , n68774 );
xor ( n68777 , n68454 , n68686 );
and ( n68778 , n30219 , n68718 );
and ( n68779 , n68777 , n68778 );
xor ( n68780 , n68777 , n68778 );
xor ( n68781 , n68458 , n68684 );
and ( n68782 , n30224 , n68718 );
and ( n68783 , n68781 , n68782 );
xor ( n68784 , n68781 , n68782 );
xor ( n68785 , n68462 , n68682 );
and ( n68786 , n30229 , n68718 );
and ( n68787 , n68785 , n68786 );
xor ( n68788 , n68785 , n68786 );
xor ( n68789 , n68466 , n68680 );
and ( n68790 , n30234 , n68718 );
and ( n68791 , n68789 , n68790 );
xor ( n68792 , n68789 , n68790 );
xor ( n68793 , n68470 , n68678 );
and ( n68794 , n30239 , n68718 );
and ( n68795 , n68793 , n68794 );
xor ( n68796 , n68793 , n68794 );
xor ( n68797 , n68474 , n68676 );
and ( n68798 , n30244 , n68718 );
and ( n68799 , n68797 , n68798 );
xor ( n68800 , n68797 , n68798 );
xor ( n68801 , n68478 , n68674 );
and ( n68802 , n30249 , n68718 );
and ( n68803 , n68801 , n68802 );
xor ( n68804 , n68801 , n68802 );
xor ( n68805 , n68482 , n68672 );
and ( n68806 , n30254 , n68718 );
and ( n68807 , n68805 , n68806 );
xor ( n68808 , n68805 , n68806 );
xor ( n68809 , n68486 , n68670 );
and ( n68810 , n30259 , n68718 );
and ( n68811 , n68809 , n68810 );
xor ( n68812 , n68809 , n68810 );
xor ( n68813 , n68490 , n68668 );
and ( n68814 , n30264 , n68718 );
and ( n68815 , n68813 , n68814 );
xor ( n68816 , n68813 , n68814 );
xor ( n68817 , n68494 , n68666 );
and ( n68818 , n30269 , n68718 );
and ( n68819 , n68817 , n68818 );
xor ( n68820 , n68817 , n68818 );
xor ( n68821 , n68498 , n68664 );
and ( n68822 , n30274 , n68718 );
and ( n68823 , n68821 , n68822 );
xor ( n68824 , n68821 , n68822 );
xor ( n68825 , n68502 , n68662 );
and ( n68826 , n30279 , n68718 );
and ( n68827 , n68825 , n68826 );
xor ( n68828 , n68825 , n68826 );
xor ( n68829 , n68506 , n68660 );
and ( n68830 , n30284 , n68718 );
and ( n68831 , n68829 , n68830 );
xor ( n68832 , n68829 , n68830 );
xor ( n68833 , n68510 , n68658 );
and ( n68834 , n30289 , n68718 );
and ( n68835 , n68833 , n68834 );
xor ( n68836 , n68833 , n68834 );
xor ( n68837 , n68514 , n68656 );
and ( n68838 , n30294 , n68718 );
and ( n68839 , n68837 , n68838 );
xor ( n68840 , n68837 , n68838 );
xor ( n68841 , n68518 , n68654 );
and ( n68842 , n30299 , n68718 );
and ( n68843 , n68841 , n68842 );
xor ( n68844 , n68841 , n68842 );
xor ( n68845 , n68522 , n68652 );
and ( n68846 , n30304 , n68718 );
and ( n68847 , n68845 , n68846 );
xor ( n68848 , n68845 , n68846 );
xor ( n68849 , n68526 , n68650 );
and ( n68850 , n30309 , n68718 );
and ( n68851 , n68849 , n68850 );
xor ( n68852 , n68849 , n68850 );
xor ( n68853 , n68530 , n68648 );
and ( n68854 , n30314 , n68718 );
and ( n68855 , n68853 , n68854 );
xor ( n68856 , n68853 , n68854 );
xor ( n68857 , n68534 , n68646 );
and ( n68858 , n30319 , n68718 );
and ( n68859 , n68857 , n68858 );
xor ( n68860 , n68857 , n68858 );
xor ( n68861 , n68538 , n68644 );
and ( n68862 , n30324 , n68718 );
and ( n68863 , n68861 , n68862 );
xor ( n68864 , n68861 , n68862 );
xor ( n68865 , n68542 , n68642 );
and ( n68866 , n30329 , n68718 );
and ( n68867 , n68865 , n68866 );
xor ( n68868 , n68865 , n68866 );
xor ( n68869 , n68546 , n68640 );
and ( n68870 , n30334 , n68718 );
and ( n68871 , n68869 , n68870 );
xor ( n68872 , n68869 , n68870 );
xor ( n68873 , n68550 , n68638 );
and ( n68874 , n30339 , n68718 );
and ( n68875 , n68873 , n68874 );
xor ( n68876 , n68873 , n68874 );
xor ( n68877 , n68554 , n68636 );
and ( n68878 , n30344 , n68718 );
and ( n68879 , n68877 , n68878 );
xor ( n68880 , n68877 , n68878 );
xor ( n68881 , n68558 , n68634 );
and ( n68882 , n30349 , n68718 );
and ( n68883 , n68881 , n68882 );
xor ( n68884 , n68881 , n68882 );
xor ( n68885 , n68562 , n68632 );
and ( n68886 , n30354 , n68718 );
and ( n68887 , n68885 , n68886 );
xor ( n68888 , n68885 , n68886 );
xor ( n68889 , n68566 , n68630 );
and ( n68890 , n30359 , n68718 );
and ( n68891 , n68889 , n68890 );
xor ( n68892 , n68889 , n68890 );
xor ( n68893 , n68570 , n68628 );
and ( n68894 , n30364 , n68718 );
and ( n68895 , n68893 , n68894 );
xor ( n68896 , n68893 , n68894 );
xor ( n68897 , n68574 , n68626 );
and ( n68898 , n30369 , n68718 );
and ( n68899 , n68897 , n68898 );
xor ( n68900 , n68897 , n68898 );
xor ( n68901 , n68578 , n68624 );
and ( n68902 , n30374 , n68718 );
and ( n68903 , n68901 , n68902 );
xor ( n68904 , n68901 , n68902 );
xor ( n68905 , n68582 , n68622 );
and ( n68906 , n30379 , n68718 );
and ( n68907 , n68905 , n68906 );
xor ( n68908 , n68905 , n68906 );
xor ( n68909 , n68586 , n68620 );
and ( n68910 , n30384 , n68718 );
and ( n68911 , n68909 , n68910 );
xor ( n68912 , n68909 , n68910 );
xor ( n68913 , n68590 , n68618 );
and ( n68914 , n30389 , n68718 );
and ( n68915 , n68913 , n68914 );
xor ( n68916 , n68913 , n68914 );
xor ( n68917 , n68594 , n68616 );
and ( n68918 , n30394 , n68718 );
and ( n68919 , n68917 , n68918 );
xor ( n68920 , n68917 , n68918 );
xor ( n68921 , n68598 , n68614 );
and ( n68922 , n30399 , n68718 );
and ( n68923 , n68921 , n68922 );
xor ( n68924 , n68921 , n68922 );
xor ( n68925 , n68602 , n68612 );
and ( n68926 , n30404 , n68718 );
and ( n68927 , n68925 , n68926 );
xor ( n68928 , n68925 , n68926 );
xor ( n68929 , n68606 , n68610 );
and ( n68930 , n30409 , n68718 );
and ( n68931 , n68929 , n68930 );
buf ( n68932 , n68931 );
and ( n68933 , n68928 , n68932 );
or ( n68934 , n68927 , n68933 );
and ( n68935 , n68924 , n68934 );
or ( n68936 , n68923 , n68935 );
and ( n68937 , n68920 , n68936 );
or ( n68938 , n68919 , n68937 );
and ( n68939 , n68916 , n68938 );
or ( n68940 , n68915 , n68939 );
and ( n68941 , n68912 , n68940 );
or ( n68942 , n68911 , n68941 );
and ( n68943 , n68908 , n68942 );
or ( n68944 , n68907 , n68943 );
and ( n68945 , n68904 , n68944 );
or ( n68946 , n68903 , n68945 );
and ( n68947 , n68900 , n68946 );
or ( n68948 , n68899 , n68947 );
and ( n68949 , n68896 , n68948 );
or ( n68950 , n68895 , n68949 );
and ( n68951 , n68892 , n68950 );
or ( n68952 , n68891 , n68951 );
and ( n68953 , n68888 , n68952 );
or ( n68954 , n68887 , n68953 );
and ( n68955 , n68884 , n68954 );
or ( n68956 , n68883 , n68955 );
and ( n68957 , n68880 , n68956 );
or ( n68958 , n68879 , n68957 );
and ( n68959 , n68876 , n68958 );
or ( n68960 , n68875 , n68959 );
and ( n68961 , n68872 , n68960 );
or ( n68962 , n68871 , n68961 );
and ( n68963 , n68868 , n68962 );
or ( n68964 , n68867 , n68963 );
and ( n68965 , n68864 , n68964 );
or ( n68966 , n68863 , n68965 );
and ( n68967 , n68860 , n68966 );
or ( n68968 , n68859 , n68967 );
and ( n68969 , n68856 , n68968 );
or ( n68970 , n68855 , n68969 );
and ( n68971 , n68852 , n68970 );
or ( n68972 , n68851 , n68971 );
and ( n68973 , n68848 , n68972 );
or ( n68974 , n68847 , n68973 );
and ( n68975 , n68844 , n68974 );
or ( n68976 , n68843 , n68975 );
and ( n68977 , n68840 , n68976 );
or ( n68978 , n68839 , n68977 );
and ( n68979 , n68836 , n68978 );
or ( n68980 , n68835 , n68979 );
and ( n68981 , n68832 , n68980 );
or ( n68982 , n68831 , n68981 );
and ( n68983 , n68828 , n68982 );
or ( n68984 , n68827 , n68983 );
and ( n68985 , n68824 , n68984 );
or ( n68986 , n68823 , n68985 );
and ( n68987 , n68820 , n68986 );
or ( n68988 , n68819 , n68987 );
and ( n68989 , n68816 , n68988 );
or ( n68990 , n68815 , n68989 );
and ( n68991 , n68812 , n68990 );
or ( n68992 , n68811 , n68991 );
and ( n68993 , n68808 , n68992 );
or ( n68994 , n68807 , n68993 );
and ( n68995 , n68804 , n68994 );
or ( n68996 , n68803 , n68995 );
and ( n68997 , n68800 , n68996 );
or ( n68998 , n68799 , n68997 );
and ( n68999 , n68796 , n68998 );
or ( n69000 , n68795 , n68999 );
and ( n69001 , n68792 , n69000 );
or ( n69002 , n68791 , n69001 );
and ( n69003 , n68788 , n69002 );
or ( n69004 , n68787 , n69003 );
and ( n69005 , n68784 , n69004 );
or ( n69006 , n68783 , n69005 );
and ( n69007 , n68780 , n69006 );
or ( n69008 , n68779 , n69007 );
and ( n69009 , n68776 , n69008 );
or ( n69010 , n68775 , n69009 );
and ( n69011 , n68772 , n69010 );
or ( n69012 , n68771 , n69011 );
and ( n69013 , n68768 , n69012 );
or ( n69014 , n68767 , n69013 );
and ( n69015 , n68764 , n69014 );
or ( n69016 , n68763 , n69015 );
and ( n69017 , n68760 , n69016 );
or ( n69018 , n68759 , n69017 );
and ( n69019 , n68756 , n69018 );
or ( n69020 , n68755 , n69019 );
and ( n69021 , n68752 , n69020 );
or ( n69022 , n68751 , n69021 );
and ( n69023 , n68748 , n69022 );
or ( n69024 , n68747 , n69023 );
and ( n69025 , n68744 , n69024 );
or ( n69026 , n68743 , n69025 );
and ( n69027 , n68740 , n69026 );
or ( n69028 , n68739 , n69027 );
and ( n69029 , n68736 , n69028 );
or ( n69030 , n68735 , n69029 );
and ( n69031 , n68732 , n69030 );
or ( n69032 , n68731 , n69031 );
and ( n69033 , n68728 , n69032 );
or ( n69034 , n68727 , n69033 );
and ( n69035 , n68724 , n69034 );
or ( n69036 , n68723 , n69035 );
xor ( n69037 , n68720 , n69036 );
buf ( n69038 , n17958 );
and ( n69039 , n30149 , n69038 );
xor ( n69040 , n69037 , n69039 );
xor ( n69041 , n68724 , n69034 );
and ( n69042 , n30154 , n69038 );
and ( n69043 , n69041 , n69042 );
xor ( n69044 , n69041 , n69042 );
xor ( n69045 , n68728 , n69032 );
and ( n69046 , n30159 , n69038 );
and ( n69047 , n69045 , n69046 );
xor ( n69048 , n69045 , n69046 );
xor ( n69049 , n68732 , n69030 );
and ( n69050 , n30164 , n69038 );
and ( n69051 , n69049 , n69050 );
xor ( n69052 , n69049 , n69050 );
xor ( n69053 , n68736 , n69028 );
and ( n69054 , n30169 , n69038 );
and ( n69055 , n69053 , n69054 );
xor ( n69056 , n69053 , n69054 );
xor ( n69057 , n68740 , n69026 );
and ( n69058 , n30174 , n69038 );
and ( n69059 , n69057 , n69058 );
xor ( n69060 , n69057 , n69058 );
xor ( n69061 , n68744 , n69024 );
and ( n69062 , n30179 , n69038 );
and ( n69063 , n69061 , n69062 );
xor ( n69064 , n69061 , n69062 );
xor ( n69065 , n68748 , n69022 );
and ( n69066 , n30184 , n69038 );
and ( n69067 , n69065 , n69066 );
xor ( n69068 , n69065 , n69066 );
xor ( n69069 , n68752 , n69020 );
and ( n69070 , n30189 , n69038 );
and ( n69071 , n69069 , n69070 );
xor ( n69072 , n69069 , n69070 );
xor ( n69073 , n68756 , n69018 );
and ( n69074 , n30194 , n69038 );
and ( n69075 , n69073 , n69074 );
xor ( n69076 , n69073 , n69074 );
xor ( n69077 , n68760 , n69016 );
and ( n69078 , n30199 , n69038 );
and ( n69079 , n69077 , n69078 );
xor ( n69080 , n69077 , n69078 );
xor ( n69081 , n68764 , n69014 );
and ( n69082 , n30204 , n69038 );
and ( n69083 , n69081 , n69082 );
xor ( n69084 , n69081 , n69082 );
xor ( n69085 , n68768 , n69012 );
and ( n69086 , n30209 , n69038 );
and ( n69087 , n69085 , n69086 );
xor ( n69088 , n69085 , n69086 );
xor ( n69089 , n68772 , n69010 );
and ( n69090 , n30214 , n69038 );
and ( n69091 , n69089 , n69090 );
xor ( n69092 , n69089 , n69090 );
xor ( n69093 , n68776 , n69008 );
and ( n69094 , n30219 , n69038 );
and ( n69095 , n69093 , n69094 );
xor ( n69096 , n69093 , n69094 );
xor ( n69097 , n68780 , n69006 );
and ( n69098 , n30224 , n69038 );
and ( n69099 , n69097 , n69098 );
xor ( n69100 , n69097 , n69098 );
xor ( n69101 , n68784 , n69004 );
and ( n69102 , n30229 , n69038 );
and ( n69103 , n69101 , n69102 );
xor ( n69104 , n69101 , n69102 );
xor ( n69105 , n68788 , n69002 );
and ( n69106 , n30234 , n69038 );
and ( n69107 , n69105 , n69106 );
xor ( n69108 , n69105 , n69106 );
xor ( n69109 , n68792 , n69000 );
and ( n69110 , n30239 , n69038 );
and ( n69111 , n69109 , n69110 );
xor ( n69112 , n69109 , n69110 );
xor ( n69113 , n68796 , n68998 );
and ( n69114 , n30244 , n69038 );
and ( n69115 , n69113 , n69114 );
xor ( n69116 , n69113 , n69114 );
xor ( n69117 , n68800 , n68996 );
and ( n69118 , n30249 , n69038 );
and ( n69119 , n69117 , n69118 );
xor ( n69120 , n69117 , n69118 );
xor ( n69121 , n68804 , n68994 );
and ( n69122 , n30254 , n69038 );
and ( n69123 , n69121 , n69122 );
xor ( n69124 , n69121 , n69122 );
xor ( n69125 , n68808 , n68992 );
and ( n69126 , n30259 , n69038 );
and ( n69127 , n69125 , n69126 );
xor ( n69128 , n69125 , n69126 );
xor ( n69129 , n68812 , n68990 );
and ( n69130 , n30264 , n69038 );
and ( n69131 , n69129 , n69130 );
xor ( n69132 , n69129 , n69130 );
xor ( n69133 , n68816 , n68988 );
and ( n69134 , n30269 , n69038 );
and ( n69135 , n69133 , n69134 );
xor ( n69136 , n69133 , n69134 );
xor ( n69137 , n68820 , n68986 );
and ( n69138 , n30274 , n69038 );
and ( n69139 , n69137 , n69138 );
xor ( n69140 , n69137 , n69138 );
xor ( n69141 , n68824 , n68984 );
and ( n69142 , n30279 , n69038 );
and ( n69143 , n69141 , n69142 );
xor ( n69144 , n69141 , n69142 );
xor ( n69145 , n68828 , n68982 );
and ( n69146 , n30284 , n69038 );
and ( n69147 , n69145 , n69146 );
xor ( n69148 , n69145 , n69146 );
xor ( n69149 , n68832 , n68980 );
and ( n69150 , n30289 , n69038 );
and ( n69151 , n69149 , n69150 );
xor ( n69152 , n69149 , n69150 );
xor ( n69153 , n68836 , n68978 );
and ( n69154 , n30294 , n69038 );
and ( n69155 , n69153 , n69154 );
xor ( n69156 , n69153 , n69154 );
xor ( n69157 , n68840 , n68976 );
and ( n69158 , n30299 , n69038 );
and ( n69159 , n69157 , n69158 );
xor ( n69160 , n69157 , n69158 );
xor ( n69161 , n68844 , n68974 );
and ( n69162 , n30304 , n69038 );
and ( n69163 , n69161 , n69162 );
xor ( n69164 , n69161 , n69162 );
xor ( n69165 , n68848 , n68972 );
and ( n69166 , n30309 , n69038 );
and ( n69167 , n69165 , n69166 );
xor ( n69168 , n69165 , n69166 );
xor ( n69169 , n68852 , n68970 );
and ( n69170 , n30314 , n69038 );
and ( n69171 , n69169 , n69170 );
xor ( n69172 , n69169 , n69170 );
xor ( n69173 , n68856 , n68968 );
and ( n69174 , n30319 , n69038 );
and ( n69175 , n69173 , n69174 );
xor ( n69176 , n69173 , n69174 );
xor ( n69177 , n68860 , n68966 );
and ( n69178 , n30324 , n69038 );
and ( n69179 , n69177 , n69178 );
xor ( n69180 , n69177 , n69178 );
xor ( n69181 , n68864 , n68964 );
and ( n69182 , n30329 , n69038 );
and ( n69183 , n69181 , n69182 );
xor ( n69184 , n69181 , n69182 );
xor ( n69185 , n68868 , n68962 );
and ( n69186 , n30334 , n69038 );
and ( n69187 , n69185 , n69186 );
xor ( n69188 , n69185 , n69186 );
xor ( n69189 , n68872 , n68960 );
and ( n69190 , n30339 , n69038 );
and ( n69191 , n69189 , n69190 );
xor ( n69192 , n69189 , n69190 );
xor ( n69193 , n68876 , n68958 );
and ( n69194 , n30344 , n69038 );
and ( n69195 , n69193 , n69194 );
xor ( n69196 , n69193 , n69194 );
xor ( n69197 , n68880 , n68956 );
and ( n69198 , n30349 , n69038 );
and ( n69199 , n69197 , n69198 );
xor ( n69200 , n69197 , n69198 );
xor ( n69201 , n68884 , n68954 );
and ( n69202 , n30354 , n69038 );
and ( n69203 , n69201 , n69202 );
xor ( n69204 , n69201 , n69202 );
xor ( n69205 , n68888 , n68952 );
and ( n69206 , n30359 , n69038 );
and ( n69207 , n69205 , n69206 );
xor ( n69208 , n69205 , n69206 );
xor ( n69209 , n68892 , n68950 );
and ( n69210 , n30364 , n69038 );
and ( n69211 , n69209 , n69210 );
xor ( n69212 , n69209 , n69210 );
xor ( n69213 , n68896 , n68948 );
and ( n69214 , n30369 , n69038 );
and ( n69215 , n69213 , n69214 );
xor ( n69216 , n69213 , n69214 );
xor ( n69217 , n68900 , n68946 );
and ( n69218 , n30374 , n69038 );
and ( n69219 , n69217 , n69218 );
xor ( n69220 , n69217 , n69218 );
xor ( n69221 , n68904 , n68944 );
and ( n69222 , n30379 , n69038 );
and ( n69223 , n69221 , n69222 );
xor ( n69224 , n69221 , n69222 );
xor ( n69225 , n68908 , n68942 );
and ( n69226 , n30384 , n69038 );
and ( n69227 , n69225 , n69226 );
xor ( n69228 , n69225 , n69226 );
xor ( n69229 , n68912 , n68940 );
and ( n69230 , n30389 , n69038 );
and ( n69231 , n69229 , n69230 );
xor ( n69232 , n69229 , n69230 );
xor ( n69233 , n68916 , n68938 );
and ( n69234 , n30394 , n69038 );
and ( n69235 , n69233 , n69234 );
xor ( n69236 , n69233 , n69234 );
xor ( n69237 , n68920 , n68936 );
and ( n69238 , n30399 , n69038 );
and ( n69239 , n69237 , n69238 );
xor ( n69240 , n69237 , n69238 );
xor ( n69241 , n68924 , n68934 );
and ( n69242 , n30404 , n69038 );
and ( n69243 , n69241 , n69242 );
xor ( n69244 , n69241 , n69242 );
xor ( n69245 , n68928 , n68932 );
and ( n69246 , n30409 , n69038 );
and ( n69247 , n69245 , n69246 );
buf ( n69248 , n69247 );
and ( n69249 , n69244 , n69248 );
or ( n69250 , n69243 , n69249 );
and ( n69251 , n69240 , n69250 );
or ( n69252 , n69239 , n69251 );
and ( n69253 , n69236 , n69252 );
or ( n69254 , n69235 , n69253 );
and ( n69255 , n69232 , n69254 );
or ( n69256 , n69231 , n69255 );
and ( n69257 , n69228 , n69256 );
or ( n69258 , n69227 , n69257 );
and ( n69259 , n69224 , n69258 );
or ( n69260 , n69223 , n69259 );
and ( n69261 , n69220 , n69260 );
or ( n69262 , n69219 , n69261 );
and ( n69263 , n69216 , n69262 );
or ( n69264 , n69215 , n69263 );
and ( n69265 , n69212 , n69264 );
or ( n69266 , n69211 , n69265 );
and ( n69267 , n69208 , n69266 );
or ( n69268 , n69207 , n69267 );
and ( n69269 , n69204 , n69268 );
or ( n69270 , n69203 , n69269 );
and ( n69271 , n69200 , n69270 );
or ( n69272 , n69199 , n69271 );
and ( n69273 , n69196 , n69272 );
or ( n69274 , n69195 , n69273 );
and ( n69275 , n69192 , n69274 );
or ( n69276 , n69191 , n69275 );
and ( n69277 , n69188 , n69276 );
or ( n69278 , n69187 , n69277 );
and ( n69279 , n69184 , n69278 );
or ( n69280 , n69183 , n69279 );
and ( n69281 , n69180 , n69280 );
or ( n69282 , n69179 , n69281 );
and ( n69283 , n69176 , n69282 );
or ( n69284 , n69175 , n69283 );
and ( n69285 , n69172 , n69284 );
or ( n69286 , n69171 , n69285 );
and ( n69287 , n69168 , n69286 );
or ( n69288 , n69167 , n69287 );
and ( n69289 , n69164 , n69288 );
or ( n69290 , n69163 , n69289 );
and ( n69291 , n69160 , n69290 );
or ( n69292 , n69159 , n69291 );
and ( n69293 , n69156 , n69292 );
or ( n69294 , n69155 , n69293 );
and ( n69295 , n69152 , n69294 );
or ( n69296 , n69151 , n69295 );
and ( n69297 , n69148 , n69296 );
or ( n69298 , n69147 , n69297 );
and ( n69299 , n69144 , n69298 );
or ( n69300 , n69143 , n69299 );
and ( n69301 , n69140 , n69300 );
or ( n69302 , n69139 , n69301 );
and ( n69303 , n69136 , n69302 );
or ( n69304 , n69135 , n69303 );
and ( n69305 , n69132 , n69304 );
or ( n69306 , n69131 , n69305 );
and ( n69307 , n69128 , n69306 );
or ( n69308 , n69127 , n69307 );
and ( n69309 , n69124 , n69308 );
or ( n69310 , n69123 , n69309 );
and ( n69311 , n69120 , n69310 );
or ( n69312 , n69119 , n69311 );
and ( n69313 , n69116 , n69312 );
or ( n69314 , n69115 , n69313 );
and ( n69315 , n69112 , n69314 );
or ( n69316 , n69111 , n69315 );
and ( n69317 , n69108 , n69316 );
or ( n69318 , n69107 , n69317 );
and ( n69319 , n69104 , n69318 );
or ( n69320 , n69103 , n69319 );
and ( n69321 , n69100 , n69320 );
or ( n69322 , n69099 , n69321 );
and ( n69323 , n69096 , n69322 );
or ( n69324 , n69095 , n69323 );
and ( n69325 , n69092 , n69324 );
or ( n69326 , n69091 , n69325 );
and ( n69327 , n69088 , n69326 );
or ( n69328 , n69087 , n69327 );
and ( n69329 , n69084 , n69328 );
or ( n69330 , n69083 , n69329 );
and ( n69331 , n69080 , n69330 );
or ( n69332 , n69079 , n69331 );
and ( n69333 , n69076 , n69332 );
or ( n69334 , n69075 , n69333 );
and ( n69335 , n69072 , n69334 );
or ( n69336 , n69071 , n69335 );
and ( n69337 , n69068 , n69336 );
or ( n69338 , n69067 , n69337 );
and ( n69339 , n69064 , n69338 );
or ( n69340 , n69063 , n69339 );
and ( n69341 , n69060 , n69340 );
or ( n69342 , n69059 , n69341 );
and ( n69343 , n69056 , n69342 );
or ( n69344 , n69055 , n69343 );
and ( n69345 , n69052 , n69344 );
or ( n69346 , n69051 , n69345 );
and ( n69347 , n69048 , n69346 );
or ( n69348 , n69047 , n69347 );
and ( n69349 , n69044 , n69348 );
or ( n69350 , n69043 , n69349 );
xor ( n69351 , n69040 , n69350 );
buf ( n69352 , n17956 );
and ( n69353 , n30154 , n69352 );
xor ( n69354 , n69351 , n69353 );
xor ( n69355 , n69044 , n69348 );
and ( n69356 , n30159 , n69352 );
and ( n69357 , n69355 , n69356 );
xor ( n69358 , n69355 , n69356 );
xor ( n69359 , n69048 , n69346 );
and ( n69360 , n30164 , n69352 );
and ( n69361 , n69359 , n69360 );
xor ( n69362 , n69359 , n69360 );
xor ( n69363 , n69052 , n69344 );
and ( n69364 , n30169 , n69352 );
and ( n69365 , n69363 , n69364 );
xor ( n69366 , n69363 , n69364 );
xor ( n69367 , n69056 , n69342 );
and ( n69368 , n30174 , n69352 );
and ( n69369 , n69367 , n69368 );
xor ( n69370 , n69367 , n69368 );
xor ( n69371 , n69060 , n69340 );
and ( n69372 , n30179 , n69352 );
and ( n69373 , n69371 , n69372 );
xor ( n69374 , n69371 , n69372 );
xor ( n69375 , n69064 , n69338 );
and ( n69376 , n30184 , n69352 );
and ( n69377 , n69375 , n69376 );
xor ( n69378 , n69375 , n69376 );
xor ( n69379 , n69068 , n69336 );
and ( n69380 , n30189 , n69352 );
and ( n69381 , n69379 , n69380 );
xor ( n69382 , n69379 , n69380 );
xor ( n69383 , n69072 , n69334 );
and ( n69384 , n30194 , n69352 );
and ( n69385 , n69383 , n69384 );
xor ( n69386 , n69383 , n69384 );
xor ( n69387 , n69076 , n69332 );
and ( n69388 , n30199 , n69352 );
and ( n69389 , n69387 , n69388 );
xor ( n69390 , n69387 , n69388 );
xor ( n69391 , n69080 , n69330 );
and ( n69392 , n30204 , n69352 );
and ( n69393 , n69391 , n69392 );
xor ( n69394 , n69391 , n69392 );
xor ( n69395 , n69084 , n69328 );
and ( n69396 , n30209 , n69352 );
and ( n69397 , n69395 , n69396 );
xor ( n69398 , n69395 , n69396 );
xor ( n69399 , n69088 , n69326 );
and ( n69400 , n30214 , n69352 );
and ( n69401 , n69399 , n69400 );
xor ( n69402 , n69399 , n69400 );
xor ( n69403 , n69092 , n69324 );
and ( n69404 , n30219 , n69352 );
and ( n69405 , n69403 , n69404 );
xor ( n69406 , n69403 , n69404 );
xor ( n69407 , n69096 , n69322 );
and ( n69408 , n30224 , n69352 );
and ( n69409 , n69407 , n69408 );
xor ( n69410 , n69407 , n69408 );
xor ( n69411 , n69100 , n69320 );
and ( n69412 , n30229 , n69352 );
and ( n69413 , n69411 , n69412 );
xor ( n69414 , n69411 , n69412 );
xor ( n69415 , n69104 , n69318 );
and ( n69416 , n30234 , n69352 );
and ( n69417 , n69415 , n69416 );
xor ( n69418 , n69415 , n69416 );
xor ( n69419 , n69108 , n69316 );
and ( n69420 , n30239 , n69352 );
and ( n69421 , n69419 , n69420 );
xor ( n69422 , n69419 , n69420 );
xor ( n69423 , n69112 , n69314 );
and ( n69424 , n30244 , n69352 );
and ( n69425 , n69423 , n69424 );
xor ( n69426 , n69423 , n69424 );
xor ( n69427 , n69116 , n69312 );
and ( n69428 , n30249 , n69352 );
and ( n69429 , n69427 , n69428 );
xor ( n69430 , n69427 , n69428 );
xor ( n69431 , n69120 , n69310 );
and ( n69432 , n30254 , n69352 );
and ( n69433 , n69431 , n69432 );
xor ( n69434 , n69431 , n69432 );
xor ( n69435 , n69124 , n69308 );
and ( n69436 , n30259 , n69352 );
and ( n69437 , n69435 , n69436 );
xor ( n69438 , n69435 , n69436 );
xor ( n69439 , n69128 , n69306 );
and ( n69440 , n30264 , n69352 );
and ( n69441 , n69439 , n69440 );
xor ( n69442 , n69439 , n69440 );
xor ( n69443 , n69132 , n69304 );
and ( n69444 , n30269 , n69352 );
and ( n69445 , n69443 , n69444 );
xor ( n69446 , n69443 , n69444 );
xor ( n69447 , n69136 , n69302 );
and ( n69448 , n30274 , n69352 );
and ( n69449 , n69447 , n69448 );
xor ( n69450 , n69447 , n69448 );
xor ( n69451 , n69140 , n69300 );
and ( n69452 , n30279 , n69352 );
and ( n69453 , n69451 , n69452 );
xor ( n69454 , n69451 , n69452 );
xor ( n69455 , n69144 , n69298 );
and ( n69456 , n30284 , n69352 );
and ( n69457 , n69455 , n69456 );
xor ( n69458 , n69455 , n69456 );
xor ( n69459 , n69148 , n69296 );
and ( n69460 , n30289 , n69352 );
and ( n69461 , n69459 , n69460 );
xor ( n69462 , n69459 , n69460 );
xor ( n69463 , n69152 , n69294 );
and ( n69464 , n30294 , n69352 );
and ( n69465 , n69463 , n69464 );
xor ( n69466 , n69463 , n69464 );
xor ( n69467 , n69156 , n69292 );
and ( n69468 , n30299 , n69352 );
and ( n69469 , n69467 , n69468 );
xor ( n69470 , n69467 , n69468 );
xor ( n69471 , n69160 , n69290 );
and ( n69472 , n30304 , n69352 );
and ( n69473 , n69471 , n69472 );
xor ( n69474 , n69471 , n69472 );
xor ( n69475 , n69164 , n69288 );
and ( n69476 , n30309 , n69352 );
and ( n69477 , n69475 , n69476 );
xor ( n69478 , n69475 , n69476 );
xor ( n69479 , n69168 , n69286 );
and ( n69480 , n30314 , n69352 );
and ( n69481 , n69479 , n69480 );
xor ( n69482 , n69479 , n69480 );
xor ( n69483 , n69172 , n69284 );
and ( n69484 , n30319 , n69352 );
and ( n69485 , n69483 , n69484 );
xor ( n69486 , n69483 , n69484 );
xor ( n69487 , n69176 , n69282 );
and ( n69488 , n30324 , n69352 );
and ( n69489 , n69487 , n69488 );
xor ( n69490 , n69487 , n69488 );
xor ( n69491 , n69180 , n69280 );
and ( n69492 , n30329 , n69352 );
and ( n69493 , n69491 , n69492 );
xor ( n69494 , n69491 , n69492 );
xor ( n69495 , n69184 , n69278 );
and ( n69496 , n30334 , n69352 );
and ( n69497 , n69495 , n69496 );
xor ( n69498 , n69495 , n69496 );
xor ( n69499 , n69188 , n69276 );
and ( n69500 , n30339 , n69352 );
and ( n69501 , n69499 , n69500 );
xor ( n69502 , n69499 , n69500 );
xor ( n69503 , n69192 , n69274 );
and ( n69504 , n30344 , n69352 );
and ( n69505 , n69503 , n69504 );
xor ( n69506 , n69503 , n69504 );
xor ( n69507 , n69196 , n69272 );
and ( n69508 , n30349 , n69352 );
and ( n69509 , n69507 , n69508 );
xor ( n69510 , n69507 , n69508 );
xor ( n69511 , n69200 , n69270 );
and ( n69512 , n30354 , n69352 );
and ( n69513 , n69511 , n69512 );
xor ( n69514 , n69511 , n69512 );
xor ( n69515 , n69204 , n69268 );
and ( n69516 , n30359 , n69352 );
and ( n69517 , n69515 , n69516 );
xor ( n69518 , n69515 , n69516 );
xor ( n69519 , n69208 , n69266 );
and ( n69520 , n30364 , n69352 );
and ( n69521 , n69519 , n69520 );
xor ( n69522 , n69519 , n69520 );
xor ( n69523 , n69212 , n69264 );
and ( n69524 , n30369 , n69352 );
and ( n69525 , n69523 , n69524 );
xor ( n69526 , n69523 , n69524 );
xor ( n69527 , n69216 , n69262 );
and ( n69528 , n30374 , n69352 );
and ( n69529 , n69527 , n69528 );
xor ( n69530 , n69527 , n69528 );
xor ( n69531 , n69220 , n69260 );
and ( n69532 , n30379 , n69352 );
and ( n69533 , n69531 , n69532 );
xor ( n69534 , n69531 , n69532 );
xor ( n69535 , n69224 , n69258 );
and ( n69536 , n30384 , n69352 );
and ( n69537 , n69535 , n69536 );
xor ( n69538 , n69535 , n69536 );
xor ( n69539 , n69228 , n69256 );
and ( n69540 , n30389 , n69352 );
and ( n69541 , n69539 , n69540 );
xor ( n69542 , n69539 , n69540 );
xor ( n69543 , n69232 , n69254 );
and ( n69544 , n30394 , n69352 );
and ( n69545 , n69543 , n69544 );
xor ( n69546 , n69543 , n69544 );
xor ( n69547 , n69236 , n69252 );
and ( n69548 , n30399 , n69352 );
and ( n69549 , n69547 , n69548 );
xor ( n69550 , n69547 , n69548 );
xor ( n69551 , n69240 , n69250 );
and ( n69552 , n30404 , n69352 );
and ( n69553 , n69551 , n69552 );
xor ( n69554 , n69551 , n69552 );
xor ( n69555 , n69244 , n69248 );
and ( n69556 , n30409 , n69352 );
and ( n69557 , n69555 , n69556 );
buf ( n69558 , n69557 );
and ( n69559 , n69554 , n69558 );
or ( n69560 , n69553 , n69559 );
and ( n69561 , n69550 , n69560 );
or ( n69562 , n69549 , n69561 );
and ( n69563 , n69546 , n69562 );
or ( n69564 , n69545 , n69563 );
and ( n69565 , n69542 , n69564 );
or ( n69566 , n69541 , n69565 );
and ( n69567 , n69538 , n69566 );
or ( n69568 , n69537 , n69567 );
and ( n69569 , n69534 , n69568 );
or ( n69570 , n69533 , n69569 );
and ( n69571 , n69530 , n69570 );
or ( n69572 , n69529 , n69571 );
and ( n69573 , n69526 , n69572 );
or ( n69574 , n69525 , n69573 );
and ( n69575 , n69522 , n69574 );
or ( n69576 , n69521 , n69575 );
and ( n69577 , n69518 , n69576 );
or ( n69578 , n69517 , n69577 );
and ( n69579 , n69514 , n69578 );
or ( n69580 , n69513 , n69579 );
and ( n69581 , n69510 , n69580 );
or ( n69582 , n69509 , n69581 );
and ( n69583 , n69506 , n69582 );
or ( n69584 , n69505 , n69583 );
and ( n69585 , n69502 , n69584 );
or ( n69586 , n69501 , n69585 );
and ( n69587 , n69498 , n69586 );
or ( n69588 , n69497 , n69587 );
and ( n69589 , n69494 , n69588 );
or ( n69590 , n69493 , n69589 );
and ( n69591 , n69490 , n69590 );
or ( n69592 , n69489 , n69591 );
and ( n69593 , n69486 , n69592 );
or ( n69594 , n69485 , n69593 );
and ( n69595 , n69482 , n69594 );
or ( n69596 , n69481 , n69595 );
and ( n69597 , n69478 , n69596 );
or ( n69598 , n69477 , n69597 );
and ( n69599 , n69474 , n69598 );
or ( n69600 , n69473 , n69599 );
and ( n69601 , n69470 , n69600 );
or ( n69602 , n69469 , n69601 );
and ( n69603 , n69466 , n69602 );
or ( n69604 , n69465 , n69603 );
and ( n69605 , n69462 , n69604 );
or ( n69606 , n69461 , n69605 );
and ( n69607 , n69458 , n69606 );
or ( n69608 , n69457 , n69607 );
and ( n69609 , n69454 , n69608 );
or ( n69610 , n69453 , n69609 );
and ( n69611 , n69450 , n69610 );
or ( n69612 , n69449 , n69611 );
and ( n69613 , n69446 , n69612 );
or ( n69614 , n69445 , n69613 );
and ( n69615 , n69442 , n69614 );
or ( n69616 , n69441 , n69615 );
and ( n69617 , n69438 , n69616 );
or ( n69618 , n69437 , n69617 );
and ( n69619 , n69434 , n69618 );
or ( n69620 , n69433 , n69619 );
and ( n69621 , n69430 , n69620 );
or ( n69622 , n69429 , n69621 );
and ( n69623 , n69426 , n69622 );
or ( n69624 , n69425 , n69623 );
and ( n69625 , n69422 , n69624 );
or ( n69626 , n69421 , n69625 );
and ( n69627 , n69418 , n69626 );
or ( n69628 , n69417 , n69627 );
and ( n69629 , n69414 , n69628 );
or ( n69630 , n69413 , n69629 );
and ( n69631 , n69410 , n69630 );
or ( n69632 , n69409 , n69631 );
and ( n69633 , n69406 , n69632 );
or ( n69634 , n69405 , n69633 );
and ( n69635 , n69402 , n69634 );
or ( n69636 , n69401 , n69635 );
and ( n69637 , n69398 , n69636 );
or ( n69638 , n69397 , n69637 );
and ( n69639 , n69394 , n69638 );
or ( n69640 , n69393 , n69639 );
and ( n69641 , n69390 , n69640 );
or ( n69642 , n69389 , n69641 );
and ( n69643 , n69386 , n69642 );
or ( n69644 , n69385 , n69643 );
and ( n69645 , n69382 , n69644 );
or ( n69646 , n69381 , n69645 );
and ( n69647 , n69378 , n69646 );
or ( n69648 , n69377 , n69647 );
and ( n69649 , n69374 , n69648 );
or ( n69650 , n69373 , n69649 );
and ( n69651 , n69370 , n69650 );
or ( n69652 , n69369 , n69651 );
and ( n69653 , n69366 , n69652 );
or ( n69654 , n69365 , n69653 );
and ( n69655 , n69362 , n69654 );
or ( n69656 , n69361 , n69655 );
and ( n69657 , n69358 , n69656 );
or ( n69658 , n69357 , n69657 );
xor ( n69659 , n69354 , n69658 );
buf ( n69660 , n17954 );
and ( n69661 , n30159 , n69660 );
xor ( n69662 , n69659 , n69661 );
xor ( n69663 , n69358 , n69656 );
and ( n69664 , n30164 , n69660 );
and ( n69665 , n69663 , n69664 );
xor ( n69666 , n69663 , n69664 );
xor ( n69667 , n69362 , n69654 );
and ( n69668 , n30169 , n69660 );
and ( n69669 , n69667 , n69668 );
xor ( n69670 , n69667 , n69668 );
xor ( n69671 , n69366 , n69652 );
and ( n69672 , n30174 , n69660 );
and ( n69673 , n69671 , n69672 );
xor ( n69674 , n69671 , n69672 );
xor ( n69675 , n69370 , n69650 );
and ( n69676 , n30179 , n69660 );
and ( n69677 , n69675 , n69676 );
xor ( n69678 , n69675 , n69676 );
xor ( n69679 , n69374 , n69648 );
and ( n69680 , n30184 , n69660 );
and ( n69681 , n69679 , n69680 );
xor ( n69682 , n69679 , n69680 );
xor ( n69683 , n69378 , n69646 );
and ( n69684 , n30189 , n69660 );
and ( n69685 , n69683 , n69684 );
xor ( n69686 , n69683 , n69684 );
xor ( n69687 , n69382 , n69644 );
and ( n69688 , n30194 , n69660 );
and ( n69689 , n69687 , n69688 );
xor ( n69690 , n69687 , n69688 );
xor ( n69691 , n69386 , n69642 );
and ( n69692 , n30199 , n69660 );
and ( n69693 , n69691 , n69692 );
xor ( n69694 , n69691 , n69692 );
xor ( n69695 , n69390 , n69640 );
and ( n69696 , n30204 , n69660 );
and ( n69697 , n69695 , n69696 );
xor ( n69698 , n69695 , n69696 );
xor ( n69699 , n69394 , n69638 );
and ( n69700 , n30209 , n69660 );
and ( n69701 , n69699 , n69700 );
xor ( n69702 , n69699 , n69700 );
xor ( n69703 , n69398 , n69636 );
and ( n69704 , n30214 , n69660 );
and ( n69705 , n69703 , n69704 );
xor ( n69706 , n69703 , n69704 );
xor ( n69707 , n69402 , n69634 );
and ( n69708 , n30219 , n69660 );
and ( n69709 , n69707 , n69708 );
xor ( n69710 , n69707 , n69708 );
xor ( n69711 , n69406 , n69632 );
and ( n69712 , n30224 , n69660 );
and ( n69713 , n69711 , n69712 );
xor ( n69714 , n69711 , n69712 );
xor ( n69715 , n69410 , n69630 );
and ( n69716 , n30229 , n69660 );
and ( n69717 , n69715 , n69716 );
xor ( n69718 , n69715 , n69716 );
xor ( n69719 , n69414 , n69628 );
and ( n69720 , n30234 , n69660 );
and ( n69721 , n69719 , n69720 );
xor ( n69722 , n69719 , n69720 );
xor ( n69723 , n69418 , n69626 );
and ( n69724 , n30239 , n69660 );
and ( n69725 , n69723 , n69724 );
xor ( n69726 , n69723 , n69724 );
xor ( n69727 , n69422 , n69624 );
and ( n69728 , n30244 , n69660 );
and ( n69729 , n69727 , n69728 );
xor ( n69730 , n69727 , n69728 );
xor ( n69731 , n69426 , n69622 );
and ( n69732 , n30249 , n69660 );
and ( n69733 , n69731 , n69732 );
xor ( n69734 , n69731 , n69732 );
xor ( n69735 , n69430 , n69620 );
and ( n69736 , n30254 , n69660 );
and ( n69737 , n69735 , n69736 );
xor ( n69738 , n69735 , n69736 );
xor ( n69739 , n69434 , n69618 );
and ( n69740 , n30259 , n69660 );
and ( n69741 , n69739 , n69740 );
xor ( n69742 , n69739 , n69740 );
xor ( n69743 , n69438 , n69616 );
and ( n69744 , n30264 , n69660 );
and ( n69745 , n69743 , n69744 );
xor ( n69746 , n69743 , n69744 );
xor ( n69747 , n69442 , n69614 );
and ( n69748 , n30269 , n69660 );
and ( n69749 , n69747 , n69748 );
xor ( n69750 , n69747 , n69748 );
xor ( n69751 , n69446 , n69612 );
and ( n69752 , n30274 , n69660 );
and ( n69753 , n69751 , n69752 );
xor ( n69754 , n69751 , n69752 );
xor ( n69755 , n69450 , n69610 );
and ( n69756 , n30279 , n69660 );
and ( n69757 , n69755 , n69756 );
xor ( n69758 , n69755 , n69756 );
xor ( n69759 , n69454 , n69608 );
and ( n69760 , n30284 , n69660 );
and ( n69761 , n69759 , n69760 );
xor ( n69762 , n69759 , n69760 );
xor ( n69763 , n69458 , n69606 );
and ( n69764 , n30289 , n69660 );
and ( n69765 , n69763 , n69764 );
xor ( n69766 , n69763 , n69764 );
xor ( n69767 , n69462 , n69604 );
and ( n69768 , n30294 , n69660 );
and ( n69769 , n69767 , n69768 );
xor ( n69770 , n69767 , n69768 );
xor ( n69771 , n69466 , n69602 );
and ( n69772 , n30299 , n69660 );
and ( n69773 , n69771 , n69772 );
xor ( n69774 , n69771 , n69772 );
xor ( n69775 , n69470 , n69600 );
and ( n69776 , n30304 , n69660 );
and ( n69777 , n69775 , n69776 );
xor ( n69778 , n69775 , n69776 );
xor ( n69779 , n69474 , n69598 );
and ( n69780 , n30309 , n69660 );
and ( n69781 , n69779 , n69780 );
xor ( n69782 , n69779 , n69780 );
xor ( n69783 , n69478 , n69596 );
and ( n69784 , n30314 , n69660 );
and ( n69785 , n69783 , n69784 );
xor ( n69786 , n69783 , n69784 );
xor ( n69787 , n69482 , n69594 );
and ( n69788 , n30319 , n69660 );
and ( n69789 , n69787 , n69788 );
xor ( n69790 , n69787 , n69788 );
xor ( n69791 , n69486 , n69592 );
and ( n69792 , n30324 , n69660 );
and ( n69793 , n69791 , n69792 );
xor ( n69794 , n69791 , n69792 );
xor ( n69795 , n69490 , n69590 );
and ( n69796 , n30329 , n69660 );
and ( n69797 , n69795 , n69796 );
xor ( n69798 , n69795 , n69796 );
xor ( n69799 , n69494 , n69588 );
and ( n69800 , n30334 , n69660 );
and ( n69801 , n69799 , n69800 );
xor ( n69802 , n69799 , n69800 );
xor ( n69803 , n69498 , n69586 );
and ( n69804 , n30339 , n69660 );
and ( n69805 , n69803 , n69804 );
xor ( n69806 , n69803 , n69804 );
xor ( n69807 , n69502 , n69584 );
and ( n69808 , n30344 , n69660 );
and ( n69809 , n69807 , n69808 );
xor ( n69810 , n69807 , n69808 );
xor ( n69811 , n69506 , n69582 );
and ( n69812 , n30349 , n69660 );
and ( n69813 , n69811 , n69812 );
xor ( n69814 , n69811 , n69812 );
xor ( n69815 , n69510 , n69580 );
and ( n69816 , n30354 , n69660 );
and ( n69817 , n69815 , n69816 );
xor ( n69818 , n69815 , n69816 );
xor ( n69819 , n69514 , n69578 );
and ( n69820 , n30359 , n69660 );
and ( n69821 , n69819 , n69820 );
xor ( n69822 , n69819 , n69820 );
xor ( n69823 , n69518 , n69576 );
and ( n69824 , n30364 , n69660 );
and ( n69825 , n69823 , n69824 );
xor ( n69826 , n69823 , n69824 );
xor ( n69827 , n69522 , n69574 );
and ( n69828 , n30369 , n69660 );
and ( n69829 , n69827 , n69828 );
xor ( n69830 , n69827 , n69828 );
xor ( n69831 , n69526 , n69572 );
and ( n69832 , n30374 , n69660 );
and ( n69833 , n69831 , n69832 );
xor ( n69834 , n69831 , n69832 );
xor ( n69835 , n69530 , n69570 );
and ( n69836 , n30379 , n69660 );
and ( n69837 , n69835 , n69836 );
xor ( n69838 , n69835 , n69836 );
xor ( n69839 , n69534 , n69568 );
and ( n69840 , n30384 , n69660 );
and ( n69841 , n69839 , n69840 );
xor ( n69842 , n69839 , n69840 );
xor ( n69843 , n69538 , n69566 );
and ( n69844 , n30389 , n69660 );
and ( n69845 , n69843 , n69844 );
xor ( n69846 , n69843 , n69844 );
xor ( n69847 , n69542 , n69564 );
and ( n69848 , n30394 , n69660 );
and ( n69849 , n69847 , n69848 );
xor ( n69850 , n69847 , n69848 );
xor ( n69851 , n69546 , n69562 );
and ( n69852 , n30399 , n69660 );
and ( n69853 , n69851 , n69852 );
xor ( n69854 , n69851 , n69852 );
xor ( n69855 , n69550 , n69560 );
and ( n69856 , n30404 , n69660 );
and ( n69857 , n69855 , n69856 );
xor ( n69858 , n69855 , n69856 );
xor ( n69859 , n69554 , n69558 );
and ( n69860 , n30409 , n69660 );
and ( n69861 , n69859 , n69860 );
buf ( n69862 , n69861 );
and ( n69863 , n69858 , n69862 );
or ( n69864 , n69857 , n69863 );
and ( n69865 , n69854 , n69864 );
or ( n69866 , n69853 , n69865 );
and ( n69867 , n69850 , n69866 );
or ( n69868 , n69849 , n69867 );
and ( n69869 , n69846 , n69868 );
or ( n69870 , n69845 , n69869 );
and ( n69871 , n69842 , n69870 );
or ( n69872 , n69841 , n69871 );
and ( n69873 , n69838 , n69872 );
or ( n69874 , n69837 , n69873 );
and ( n69875 , n69834 , n69874 );
or ( n69876 , n69833 , n69875 );
and ( n69877 , n69830 , n69876 );
or ( n69878 , n69829 , n69877 );
and ( n69879 , n69826 , n69878 );
or ( n69880 , n69825 , n69879 );
and ( n69881 , n69822 , n69880 );
or ( n69882 , n69821 , n69881 );
and ( n69883 , n69818 , n69882 );
or ( n69884 , n69817 , n69883 );
and ( n69885 , n69814 , n69884 );
or ( n69886 , n69813 , n69885 );
and ( n69887 , n69810 , n69886 );
or ( n69888 , n69809 , n69887 );
and ( n69889 , n69806 , n69888 );
or ( n69890 , n69805 , n69889 );
and ( n69891 , n69802 , n69890 );
or ( n69892 , n69801 , n69891 );
and ( n69893 , n69798 , n69892 );
or ( n69894 , n69797 , n69893 );
and ( n69895 , n69794 , n69894 );
or ( n69896 , n69793 , n69895 );
and ( n69897 , n69790 , n69896 );
or ( n69898 , n69789 , n69897 );
and ( n69899 , n69786 , n69898 );
or ( n69900 , n69785 , n69899 );
and ( n69901 , n69782 , n69900 );
or ( n69902 , n69781 , n69901 );
and ( n69903 , n69778 , n69902 );
or ( n69904 , n69777 , n69903 );
and ( n69905 , n69774 , n69904 );
or ( n69906 , n69773 , n69905 );
and ( n69907 , n69770 , n69906 );
or ( n69908 , n69769 , n69907 );
and ( n69909 , n69766 , n69908 );
or ( n69910 , n69765 , n69909 );
and ( n69911 , n69762 , n69910 );
or ( n69912 , n69761 , n69911 );
and ( n69913 , n69758 , n69912 );
or ( n69914 , n69757 , n69913 );
and ( n69915 , n69754 , n69914 );
or ( n69916 , n69753 , n69915 );
and ( n69917 , n69750 , n69916 );
or ( n69918 , n69749 , n69917 );
and ( n69919 , n69746 , n69918 );
or ( n69920 , n69745 , n69919 );
and ( n69921 , n69742 , n69920 );
or ( n69922 , n69741 , n69921 );
and ( n69923 , n69738 , n69922 );
or ( n69924 , n69737 , n69923 );
and ( n69925 , n69734 , n69924 );
or ( n69926 , n69733 , n69925 );
and ( n69927 , n69730 , n69926 );
or ( n69928 , n69729 , n69927 );
and ( n69929 , n69726 , n69928 );
or ( n69930 , n69725 , n69929 );
and ( n69931 , n69722 , n69930 );
or ( n69932 , n69721 , n69931 );
and ( n69933 , n69718 , n69932 );
or ( n69934 , n69717 , n69933 );
and ( n69935 , n69714 , n69934 );
or ( n69936 , n69713 , n69935 );
and ( n69937 , n69710 , n69936 );
or ( n69938 , n69709 , n69937 );
and ( n69939 , n69706 , n69938 );
or ( n69940 , n69705 , n69939 );
and ( n69941 , n69702 , n69940 );
or ( n69942 , n69701 , n69941 );
and ( n69943 , n69698 , n69942 );
or ( n69944 , n69697 , n69943 );
and ( n69945 , n69694 , n69944 );
or ( n69946 , n69693 , n69945 );
and ( n69947 , n69690 , n69946 );
or ( n69948 , n69689 , n69947 );
and ( n69949 , n69686 , n69948 );
or ( n69950 , n69685 , n69949 );
and ( n69951 , n69682 , n69950 );
or ( n69952 , n69681 , n69951 );
and ( n69953 , n69678 , n69952 );
or ( n69954 , n69677 , n69953 );
and ( n69955 , n69674 , n69954 );
or ( n69956 , n69673 , n69955 );
and ( n69957 , n69670 , n69956 );
or ( n69958 , n69669 , n69957 );
and ( n69959 , n69666 , n69958 );
or ( n69960 , n69665 , n69959 );
xor ( n69961 , n69662 , n69960 );
buf ( n69962 , n17952 );
and ( n69963 , n30164 , n69962 );
xor ( n69964 , n69961 , n69963 );
xor ( n69965 , n69666 , n69958 );
and ( n69966 , n30169 , n69962 );
and ( n69967 , n69965 , n69966 );
xor ( n69968 , n69965 , n69966 );
xor ( n69969 , n69670 , n69956 );
and ( n69970 , n30174 , n69962 );
and ( n69971 , n69969 , n69970 );
xor ( n69972 , n69969 , n69970 );
xor ( n69973 , n69674 , n69954 );
and ( n69974 , n30179 , n69962 );
and ( n69975 , n69973 , n69974 );
xor ( n69976 , n69973 , n69974 );
xor ( n69977 , n69678 , n69952 );
and ( n69978 , n30184 , n69962 );
and ( n69979 , n69977 , n69978 );
xor ( n69980 , n69977 , n69978 );
xor ( n69981 , n69682 , n69950 );
and ( n69982 , n30189 , n69962 );
and ( n69983 , n69981 , n69982 );
xor ( n69984 , n69981 , n69982 );
xor ( n69985 , n69686 , n69948 );
and ( n69986 , n30194 , n69962 );
and ( n69987 , n69985 , n69986 );
xor ( n69988 , n69985 , n69986 );
xor ( n69989 , n69690 , n69946 );
and ( n69990 , n30199 , n69962 );
and ( n69991 , n69989 , n69990 );
xor ( n69992 , n69989 , n69990 );
xor ( n69993 , n69694 , n69944 );
and ( n69994 , n30204 , n69962 );
and ( n69995 , n69993 , n69994 );
xor ( n69996 , n69993 , n69994 );
xor ( n69997 , n69698 , n69942 );
and ( n69998 , n30209 , n69962 );
and ( n69999 , n69997 , n69998 );
xor ( n70000 , n69997 , n69998 );
xor ( n70001 , n69702 , n69940 );
and ( n70002 , n30214 , n69962 );
and ( n70003 , n70001 , n70002 );
xor ( n70004 , n70001 , n70002 );
xor ( n70005 , n69706 , n69938 );
and ( n70006 , n30219 , n69962 );
and ( n70007 , n70005 , n70006 );
xor ( n70008 , n70005 , n70006 );
xor ( n70009 , n69710 , n69936 );
and ( n70010 , n30224 , n69962 );
and ( n70011 , n70009 , n70010 );
xor ( n70012 , n70009 , n70010 );
xor ( n70013 , n69714 , n69934 );
and ( n70014 , n30229 , n69962 );
and ( n70015 , n70013 , n70014 );
xor ( n70016 , n70013 , n70014 );
xor ( n70017 , n69718 , n69932 );
and ( n70018 , n30234 , n69962 );
and ( n70019 , n70017 , n70018 );
xor ( n70020 , n70017 , n70018 );
xor ( n70021 , n69722 , n69930 );
and ( n70022 , n30239 , n69962 );
and ( n70023 , n70021 , n70022 );
xor ( n70024 , n70021 , n70022 );
xor ( n70025 , n69726 , n69928 );
and ( n70026 , n30244 , n69962 );
and ( n70027 , n70025 , n70026 );
xor ( n70028 , n70025 , n70026 );
xor ( n70029 , n69730 , n69926 );
and ( n70030 , n30249 , n69962 );
and ( n70031 , n70029 , n70030 );
xor ( n70032 , n70029 , n70030 );
xor ( n70033 , n69734 , n69924 );
and ( n70034 , n30254 , n69962 );
and ( n70035 , n70033 , n70034 );
xor ( n70036 , n70033 , n70034 );
xor ( n70037 , n69738 , n69922 );
and ( n70038 , n30259 , n69962 );
and ( n70039 , n70037 , n70038 );
xor ( n70040 , n70037 , n70038 );
xor ( n70041 , n69742 , n69920 );
and ( n70042 , n30264 , n69962 );
and ( n70043 , n70041 , n70042 );
xor ( n70044 , n70041 , n70042 );
xor ( n70045 , n69746 , n69918 );
and ( n70046 , n30269 , n69962 );
and ( n70047 , n70045 , n70046 );
xor ( n70048 , n70045 , n70046 );
xor ( n70049 , n69750 , n69916 );
and ( n70050 , n30274 , n69962 );
and ( n70051 , n70049 , n70050 );
xor ( n70052 , n70049 , n70050 );
xor ( n70053 , n69754 , n69914 );
and ( n70054 , n30279 , n69962 );
and ( n70055 , n70053 , n70054 );
xor ( n70056 , n70053 , n70054 );
xor ( n70057 , n69758 , n69912 );
and ( n70058 , n30284 , n69962 );
and ( n70059 , n70057 , n70058 );
xor ( n70060 , n70057 , n70058 );
xor ( n70061 , n69762 , n69910 );
and ( n70062 , n30289 , n69962 );
and ( n70063 , n70061 , n70062 );
xor ( n70064 , n70061 , n70062 );
xor ( n70065 , n69766 , n69908 );
and ( n70066 , n30294 , n69962 );
and ( n70067 , n70065 , n70066 );
xor ( n70068 , n70065 , n70066 );
xor ( n70069 , n69770 , n69906 );
and ( n70070 , n30299 , n69962 );
and ( n70071 , n70069 , n70070 );
xor ( n70072 , n70069 , n70070 );
xor ( n70073 , n69774 , n69904 );
and ( n70074 , n30304 , n69962 );
and ( n70075 , n70073 , n70074 );
xor ( n70076 , n70073 , n70074 );
xor ( n70077 , n69778 , n69902 );
and ( n70078 , n30309 , n69962 );
and ( n70079 , n70077 , n70078 );
xor ( n70080 , n70077 , n70078 );
xor ( n70081 , n69782 , n69900 );
and ( n70082 , n30314 , n69962 );
and ( n70083 , n70081 , n70082 );
xor ( n70084 , n70081 , n70082 );
xor ( n70085 , n69786 , n69898 );
and ( n70086 , n30319 , n69962 );
and ( n70087 , n70085 , n70086 );
xor ( n70088 , n70085 , n70086 );
xor ( n70089 , n69790 , n69896 );
and ( n70090 , n30324 , n69962 );
and ( n70091 , n70089 , n70090 );
xor ( n70092 , n70089 , n70090 );
xor ( n70093 , n69794 , n69894 );
and ( n70094 , n30329 , n69962 );
and ( n70095 , n70093 , n70094 );
xor ( n70096 , n70093 , n70094 );
xor ( n70097 , n69798 , n69892 );
and ( n70098 , n30334 , n69962 );
and ( n70099 , n70097 , n70098 );
xor ( n70100 , n70097 , n70098 );
xor ( n70101 , n69802 , n69890 );
and ( n70102 , n30339 , n69962 );
and ( n70103 , n70101 , n70102 );
xor ( n70104 , n70101 , n70102 );
xor ( n70105 , n69806 , n69888 );
and ( n70106 , n30344 , n69962 );
and ( n70107 , n70105 , n70106 );
xor ( n70108 , n70105 , n70106 );
xor ( n70109 , n69810 , n69886 );
and ( n70110 , n30349 , n69962 );
and ( n70111 , n70109 , n70110 );
xor ( n70112 , n70109 , n70110 );
xor ( n70113 , n69814 , n69884 );
and ( n70114 , n30354 , n69962 );
and ( n70115 , n70113 , n70114 );
xor ( n70116 , n70113 , n70114 );
xor ( n70117 , n69818 , n69882 );
and ( n70118 , n30359 , n69962 );
and ( n70119 , n70117 , n70118 );
xor ( n70120 , n70117 , n70118 );
xor ( n70121 , n69822 , n69880 );
and ( n70122 , n30364 , n69962 );
and ( n70123 , n70121 , n70122 );
xor ( n70124 , n70121 , n70122 );
xor ( n70125 , n69826 , n69878 );
and ( n70126 , n30369 , n69962 );
and ( n70127 , n70125 , n70126 );
xor ( n70128 , n70125 , n70126 );
xor ( n70129 , n69830 , n69876 );
and ( n70130 , n30374 , n69962 );
and ( n70131 , n70129 , n70130 );
xor ( n70132 , n70129 , n70130 );
xor ( n70133 , n69834 , n69874 );
and ( n70134 , n30379 , n69962 );
and ( n70135 , n70133 , n70134 );
xor ( n70136 , n70133 , n70134 );
xor ( n70137 , n69838 , n69872 );
and ( n70138 , n30384 , n69962 );
and ( n70139 , n70137 , n70138 );
xor ( n70140 , n70137 , n70138 );
xor ( n70141 , n69842 , n69870 );
and ( n70142 , n30389 , n69962 );
and ( n70143 , n70141 , n70142 );
xor ( n70144 , n70141 , n70142 );
xor ( n70145 , n69846 , n69868 );
and ( n70146 , n30394 , n69962 );
and ( n70147 , n70145 , n70146 );
xor ( n70148 , n70145 , n70146 );
xor ( n70149 , n69850 , n69866 );
and ( n70150 , n30399 , n69962 );
and ( n70151 , n70149 , n70150 );
xor ( n70152 , n70149 , n70150 );
xor ( n70153 , n69854 , n69864 );
and ( n70154 , n30404 , n69962 );
and ( n70155 , n70153 , n70154 );
xor ( n70156 , n70153 , n70154 );
xor ( n70157 , n69858 , n69862 );
and ( n70158 , n30409 , n69962 );
and ( n70159 , n70157 , n70158 );
buf ( n70160 , n70159 );
and ( n70161 , n70156 , n70160 );
or ( n70162 , n70155 , n70161 );
and ( n70163 , n70152 , n70162 );
or ( n70164 , n70151 , n70163 );
and ( n70165 , n70148 , n70164 );
or ( n70166 , n70147 , n70165 );
and ( n70167 , n70144 , n70166 );
or ( n70168 , n70143 , n70167 );
and ( n70169 , n70140 , n70168 );
or ( n70170 , n70139 , n70169 );
and ( n70171 , n70136 , n70170 );
or ( n70172 , n70135 , n70171 );
and ( n70173 , n70132 , n70172 );
or ( n70174 , n70131 , n70173 );
and ( n70175 , n70128 , n70174 );
or ( n70176 , n70127 , n70175 );
and ( n70177 , n70124 , n70176 );
or ( n70178 , n70123 , n70177 );
and ( n70179 , n70120 , n70178 );
or ( n70180 , n70119 , n70179 );
and ( n70181 , n70116 , n70180 );
or ( n70182 , n70115 , n70181 );
and ( n70183 , n70112 , n70182 );
or ( n70184 , n70111 , n70183 );
and ( n70185 , n70108 , n70184 );
or ( n70186 , n70107 , n70185 );
and ( n70187 , n70104 , n70186 );
or ( n70188 , n70103 , n70187 );
and ( n70189 , n70100 , n70188 );
or ( n70190 , n70099 , n70189 );
and ( n70191 , n70096 , n70190 );
or ( n70192 , n70095 , n70191 );
and ( n70193 , n70092 , n70192 );
or ( n70194 , n70091 , n70193 );
and ( n70195 , n70088 , n70194 );
or ( n70196 , n70087 , n70195 );
and ( n70197 , n70084 , n70196 );
or ( n70198 , n70083 , n70197 );
and ( n70199 , n70080 , n70198 );
or ( n70200 , n70079 , n70199 );
and ( n70201 , n70076 , n70200 );
or ( n70202 , n70075 , n70201 );
and ( n70203 , n70072 , n70202 );
or ( n70204 , n70071 , n70203 );
and ( n70205 , n70068 , n70204 );
or ( n70206 , n70067 , n70205 );
and ( n70207 , n70064 , n70206 );
or ( n70208 , n70063 , n70207 );
and ( n70209 , n70060 , n70208 );
or ( n70210 , n70059 , n70209 );
and ( n70211 , n70056 , n70210 );
or ( n70212 , n70055 , n70211 );
and ( n70213 , n70052 , n70212 );
or ( n70214 , n70051 , n70213 );
and ( n70215 , n70048 , n70214 );
or ( n70216 , n70047 , n70215 );
and ( n70217 , n70044 , n70216 );
or ( n70218 , n70043 , n70217 );
and ( n70219 , n70040 , n70218 );
or ( n70220 , n70039 , n70219 );
and ( n70221 , n70036 , n70220 );
or ( n70222 , n70035 , n70221 );
and ( n70223 , n70032 , n70222 );
or ( n70224 , n70031 , n70223 );
and ( n70225 , n70028 , n70224 );
or ( n70226 , n70027 , n70225 );
and ( n70227 , n70024 , n70226 );
or ( n70228 , n70023 , n70227 );
and ( n70229 , n70020 , n70228 );
or ( n70230 , n70019 , n70229 );
and ( n70231 , n70016 , n70230 );
or ( n70232 , n70015 , n70231 );
and ( n70233 , n70012 , n70232 );
or ( n70234 , n70011 , n70233 );
and ( n70235 , n70008 , n70234 );
or ( n70236 , n70007 , n70235 );
and ( n70237 , n70004 , n70236 );
or ( n70238 , n70003 , n70237 );
and ( n70239 , n70000 , n70238 );
or ( n70240 , n69999 , n70239 );
and ( n70241 , n69996 , n70240 );
or ( n70242 , n69995 , n70241 );
and ( n70243 , n69992 , n70242 );
or ( n70244 , n69991 , n70243 );
and ( n70245 , n69988 , n70244 );
or ( n70246 , n69987 , n70245 );
and ( n70247 , n69984 , n70246 );
or ( n70248 , n69983 , n70247 );
and ( n70249 , n69980 , n70248 );
or ( n70250 , n69979 , n70249 );
and ( n70251 , n69976 , n70250 );
or ( n70252 , n69975 , n70251 );
and ( n70253 , n69972 , n70252 );
or ( n70254 , n69971 , n70253 );
and ( n70255 , n69968 , n70254 );
or ( n70256 , n69967 , n70255 );
xor ( n70257 , n69964 , n70256 );
buf ( n70258 , n17950 );
and ( n70259 , n30169 , n70258 );
xor ( n70260 , n70257 , n70259 );
xor ( n70261 , n69968 , n70254 );
and ( n70262 , n30174 , n70258 );
and ( n70263 , n70261 , n70262 );
xor ( n70264 , n70261 , n70262 );
xor ( n70265 , n69972 , n70252 );
and ( n70266 , n30179 , n70258 );
and ( n70267 , n70265 , n70266 );
xor ( n70268 , n70265 , n70266 );
xor ( n70269 , n69976 , n70250 );
and ( n70270 , n30184 , n70258 );
and ( n70271 , n70269 , n70270 );
xor ( n70272 , n70269 , n70270 );
xor ( n70273 , n69980 , n70248 );
and ( n70274 , n30189 , n70258 );
and ( n70275 , n70273 , n70274 );
xor ( n70276 , n70273 , n70274 );
xor ( n70277 , n69984 , n70246 );
and ( n70278 , n30194 , n70258 );
and ( n70279 , n70277 , n70278 );
xor ( n70280 , n70277 , n70278 );
xor ( n70281 , n69988 , n70244 );
and ( n70282 , n30199 , n70258 );
and ( n70283 , n70281 , n70282 );
xor ( n70284 , n70281 , n70282 );
xor ( n70285 , n69992 , n70242 );
and ( n70286 , n30204 , n70258 );
and ( n70287 , n70285 , n70286 );
xor ( n70288 , n70285 , n70286 );
xor ( n70289 , n69996 , n70240 );
and ( n70290 , n30209 , n70258 );
and ( n70291 , n70289 , n70290 );
xor ( n70292 , n70289 , n70290 );
xor ( n70293 , n70000 , n70238 );
and ( n70294 , n30214 , n70258 );
and ( n70295 , n70293 , n70294 );
xor ( n70296 , n70293 , n70294 );
xor ( n70297 , n70004 , n70236 );
and ( n70298 , n30219 , n70258 );
and ( n70299 , n70297 , n70298 );
xor ( n70300 , n70297 , n70298 );
xor ( n70301 , n70008 , n70234 );
and ( n70302 , n30224 , n70258 );
and ( n70303 , n70301 , n70302 );
xor ( n70304 , n70301 , n70302 );
xor ( n70305 , n70012 , n70232 );
and ( n70306 , n30229 , n70258 );
and ( n70307 , n70305 , n70306 );
xor ( n70308 , n70305 , n70306 );
xor ( n70309 , n70016 , n70230 );
and ( n70310 , n30234 , n70258 );
and ( n70311 , n70309 , n70310 );
xor ( n70312 , n70309 , n70310 );
xor ( n70313 , n70020 , n70228 );
and ( n70314 , n30239 , n70258 );
and ( n70315 , n70313 , n70314 );
xor ( n70316 , n70313 , n70314 );
xor ( n70317 , n70024 , n70226 );
and ( n70318 , n30244 , n70258 );
and ( n70319 , n70317 , n70318 );
xor ( n70320 , n70317 , n70318 );
xor ( n70321 , n70028 , n70224 );
and ( n70322 , n30249 , n70258 );
and ( n70323 , n70321 , n70322 );
xor ( n70324 , n70321 , n70322 );
xor ( n70325 , n70032 , n70222 );
and ( n70326 , n30254 , n70258 );
and ( n70327 , n70325 , n70326 );
xor ( n70328 , n70325 , n70326 );
xor ( n70329 , n70036 , n70220 );
and ( n70330 , n30259 , n70258 );
and ( n70331 , n70329 , n70330 );
xor ( n70332 , n70329 , n70330 );
xor ( n70333 , n70040 , n70218 );
and ( n70334 , n30264 , n70258 );
and ( n70335 , n70333 , n70334 );
xor ( n70336 , n70333 , n70334 );
xor ( n70337 , n70044 , n70216 );
and ( n70338 , n30269 , n70258 );
and ( n70339 , n70337 , n70338 );
xor ( n70340 , n70337 , n70338 );
xor ( n70341 , n70048 , n70214 );
and ( n70342 , n30274 , n70258 );
and ( n70343 , n70341 , n70342 );
xor ( n70344 , n70341 , n70342 );
xor ( n70345 , n70052 , n70212 );
and ( n70346 , n30279 , n70258 );
and ( n70347 , n70345 , n70346 );
xor ( n70348 , n70345 , n70346 );
xor ( n70349 , n70056 , n70210 );
and ( n70350 , n30284 , n70258 );
and ( n70351 , n70349 , n70350 );
xor ( n70352 , n70349 , n70350 );
xor ( n70353 , n70060 , n70208 );
and ( n70354 , n30289 , n70258 );
and ( n70355 , n70353 , n70354 );
xor ( n70356 , n70353 , n70354 );
xor ( n70357 , n70064 , n70206 );
and ( n70358 , n30294 , n70258 );
and ( n70359 , n70357 , n70358 );
xor ( n70360 , n70357 , n70358 );
xor ( n70361 , n70068 , n70204 );
and ( n70362 , n30299 , n70258 );
and ( n70363 , n70361 , n70362 );
xor ( n70364 , n70361 , n70362 );
xor ( n70365 , n70072 , n70202 );
and ( n70366 , n30304 , n70258 );
and ( n70367 , n70365 , n70366 );
xor ( n70368 , n70365 , n70366 );
xor ( n70369 , n70076 , n70200 );
and ( n70370 , n30309 , n70258 );
and ( n70371 , n70369 , n70370 );
xor ( n70372 , n70369 , n70370 );
xor ( n70373 , n70080 , n70198 );
and ( n70374 , n30314 , n70258 );
and ( n70375 , n70373 , n70374 );
xor ( n70376 , n70373 , n70374 );
xor ( n70377 , n70084 , n70196 );
and ( n70378 , n30319 , n70258 );
and ( n70379 , n70377 , n70378 );
xor ( n70380 , n70377 , n70378 );
xor ( n70381 , n70088 , n70194 );
and ( n70382 , n30324 , n70258 );
and ( n70383 , n70381 , n70382 );
xor ( n70384 , n70381 , n70382 );
xor ( n70385 , n70092 , n70192 );
and ( n70386 , n30329 , n70258 );
and ( n70387 , n70385 , n70386 );
xor ( n70388 , n70385 , n70386 );
xor ( n70389 , n70096 , n70190 );
and ( n70390 , n30334 , n70258 );
and ( n70391 , n70389 , n70390 );
xor ( n70392 , n70389 , n70390 );
xor ( n70393 , n70100 , n70188 );
and ( n70394 , n30339 , n70258 );
and ( n70395 , n70393 , n70394 );
xor ( n70396 , n70393 , n70394 );
xor ( n70397 , n70104 , n70186 );
and ( n70398 , n30344 , n70258 );
and ( n70399 , n70397 , n70398 );
xor ( n70400 , n70397 , n70398 );
xor ( n70401 , n70108 , n70184 );
and ( n70402 , n30349 , n70258 );
and ( n70403 , n70401 , n70402 );
xor ( n70404 , n70401 , n70402 );
xor ( n70405 , n70112 , n70182 );
and ( n70406 , n30354 , n70258 );
and ( n70407 , n70405 , n70406 );
xor ( n70408 , n70405 , n70406 );
xor ( n70409 , n70116 , n70180 );
and ( n70410 , n30359 , n70258 );
and ( n70411 , n70409 , n70410 );
xor ( n70412 , n70409 , n70410 );
xor ( n70413 , n70120 , n70178 );
and ( n70414 , n30364 , n70258 );
and ( n70415 , n70413 , n70414 );
xor ( n70416 , n70413 , n70414 );
xor ( n70417 , n70124 , n70176 );
and ( n70418 , n30369 , n70258 );
and ( n70419 , n70417 , n70418 );
xor ( n70420 , n70417 , n70418 );
xor ( n70421 , n70128 , n70174 );
and ( n70422 , n30374 , n70258 );
and ( n70423 , n70421 , n70422 );
xor ( n70424 , n70421 , n70422 );
xor ( n70425 , n70132 , n70172 );
and ( n70426 , n30379 , n70258 );
and ( n70427 , n70425 , n70426 );
xor ( n70428 , n70425 , n70426 );
xor ( n70429 , n70136 , n70170 );
and ( n70430 , n30384 , n70258 );
and ( n70431 , n70429 , n70430 );
xor ( n70432 , n70429 , n70430 );
xor ( n70433 , n70140 , n70168 );
and ( n70434 , n30389 , n70258 );
and ( n70435 , n70433 , n70434 );
xor ( n70436 , n70433 , n70434 );
xor ( n70437 , n70144 , n70166 );
and ( n70438 , n30394 , n70258 );
and ( n70439 , n70437 , n70438 );
xor ( n70440 , n70437 , n70438 );
xor ( n70441 , n70148 , n70164 );
and ( n70442 , n30399 , n70258 );
and ( n70443 , n70441 , n70442 );
xor ( n70444 , n70441 , n70442 );
xor ( n70445 , n70152 , n70162 );
and ( n70446 , n30404 , n70258 );
and ( n70447 , n70445 , n70446 );
xor ( n70448 , n70445 , n70446 );
xor ( n70449 , n70156 , n70160 );
and ( n70450 , n30409 , n70258 );
and ( n70451 , n70449 , n70450 );
buf ( n70452 , n70451 );
and ( n70453 , n70448 , n70452 );
or ( n70454 , n70447 , n70453 );
and ( n70455 , n70444 , n70454 );
or ( n70456 , n70443 , n70455 );
and ( n70457 , n70440 , n70456 );
or ( n70458 , n70439 , n70457 );
and ( n70459 , n70436 , n70458 );
or ( n70460 , n70435 , n70459 );
and ( n70461 , n70432 , n70460 );
or ( n70462 , n70431 , n70461 );
and ( n70463 , n70428 , n70462 );
or ( n70464 , n70427 , n70463 );
and ( n70465 , n70424 , n70464 );
or ( n70466 , n70423 , n70465 );
and ( n70467 , n70420 , n70466 );
or ( n70468 , n70419 , n70467 );
and ( n70469 , n70416 , n70468 );
or ( n70470 , n70415 , n70469 );
and ( n70471 , n70412 , n70470 );
or ( n70472 , n70411 , n70471 );
and ( n70473 , n70408 , n70472 );
or ( n70474 , n70407 , n70473 );
and ( n70475 , n70404 , n70474 );
or ( n70476 , n70403 , n70475 );
and ( n70477 , n70400 , n70476 );
or ( n70478 , n70399 , n70477 );
and ( n70479 , n70396 , n70478 );
or ( n70480 , n70395 , n70479 );
and ( n70481 , n70392 , n70480 );
or ( n70482 , n70391 , n70481 );
and ( n70483 , n70388 , n70482 );
or ( n70484 , n70387 , n70483 );
and ( n70485 , n70384 , n70484 );
or ( n70486 , n70383 , n70485 );
and ( n70487 , n70380 , n70486 );
or ( n70488 , n70379 , n70487 );
and ( n70489 , n70376 , n70488 );
or ( n70490 , n70375 , n70489 );
and ( n70491 , n70372 , n70490 );
or ( n70492 , n70371 , n70491 );
and ( n70493 , n70368 , n70492 );
or ( n70494 , n70367 , n70493 );
and ( n70495 , n70364 , n70494 );
or ( n70496 , n70363 , n70495 );
and ( n70497 , n70360 , n70496 );
or ( n70498 , n70359 , n70497 );
and ( n70499 , n70356 , n70498 );
or ( n70500 , n70355 , n70499 );
and ( n70501 , n70352 , n70500 );
or ( n70502 , n70351 , n70501 );
and ( n70503 , n70348 , n70502 );
or ( n70504 , n70347 , n70503 );
and ( n70505 , n70344 , n70504 );
or ( n70506 , n70343 , n70505 );
and ( n70507 , n70340 , n70506 );
or ( n70508 , n70339 , n70507 );
and ( n70509 , n70336 , n70508 );
or ( n70510 , n70335 , n70509 );
and ( n70511 , n70332 , n70510 );
or ( n70512 , n70331 , n70511 );
and ( n70513 , n70328 , n70512 );
or ( n70514 , n70327 , n70513 );
and ( n70515 , n70324 , n70514 );
or ( n70516 , n70323 , n70515 );
and ( n70517 , n70320 , n70516 );
or ( n70518 , n70319 , n70517 );
and ( n70519 , n70316 , n70518 );
or ( n70520 , n70315 , n70519 );
and ( n70521 , n70312 , n70520 );
or ( n70522 , n70311 , n70521 );
and ( n70523 , n70308 , n70522 );
or ( n70524 , n70307 , n70523 );
and ( n70525 , n70304 , n70524 );
or ( n70526 , n70303 , n70525 );
and ( n70527 , n70300 , n70526 );
or ( n70528 , n70299 , n70527 );
and ( n70529 , n70296 , n70528 );
or ( n70530 , n70295 , n70529 );
and ( n70531 , n70292 , n70530 );
or ( n70532 , n70291 , n70531 );
and ( n70533 , n70288 , n70532 );
or ( n70534 , n70287 , n70533 );
and ( n70535 , n70284 , n70534 );
or ( n70536 , n70283 , n70535 );
and ( n70537 , n70280 , n70536 );
or ( n70538 , n70279 , n70537 );
and ( n70539 , n70276 , n70538 );
or ( n70540 , n70275 , n70539 );
and ( n70541 , n70272 , n70540 );
or ( n70542 , n70271 , n70541 );
and ( n70543 , n70268 , n70542 );
or ( n70544 , n70267 , n70543 );
and ( n70545 , n70264 , n70544 );
or ( n70546 , n70263 , n70545 );
xor ( n70547 , n70260 , n70546 );
buf ( n70548 , n17948 );
and ( n70549 , n30174 , n70548 );
xor ( n70550 , n70547 , n70549 );
xor ( n70551 , n70264 , n70544 );
and ( n70552 , n30179 , n70548 );
and ( n70553 , n70551 , n70552 );
xor ( n70554 , n70551 , n70552 );
xor ( n70555 , n70268 , n70542 );
and ( n70556 , n30184 , n70548 );
and ( n70557 , n70555 , n70556 );
xor ( n70558 , n70555 , n70556 );
xor ( n70559 , n70272 , n70540 );
and ( n70560 , n30189 , n70548 );
and ( n70561 , n70559 , n70560 );
xor ( n70562 , n70559 , n70560 );
xor ( n70563 , n70276 , n70538 );
and ( n70564 , n30194 , n70548 );
and ( n70565 , n70563 , n70564 );
xor ( n70566 , n70563 , n70564 );
xor ( n70567 , n70280 , n70536 );
and ( n70568 , n30199 , n70548 );
and ( n70569 , n70567 , n70568 );
xor ( n70570 , n70567 , n70568 );
xor ( n70571 , n70284 , n70534 );
and ( n70572 , n30204 , n70548 );
and ( n70573 , n70571 , n70572 );
xor ( n70574 , n70571 , n70572 );
xor ( n70575 , n70288 , n70532 );
and ( n70576 , n30209 , n70548 );
and ( n70577 , n70575 , n70576 );
xor ( n70578 , n70575 , n70576 );
xor ( n70579 , n70292 , n70530 );
and ( n70580 , n30214 , n70548 );
and ( n70581 , n70579 , n70580 );
xor ( n70582 , n70579 , n70580 );
xor ( n70583 , n70296 , n70528 );
and ( n70584 , n30219 , n70548 );
and ( n70585 , n70583 , n70584 );
xor ( n70586 , n70583 , n70584 );
xor ( n70587 , n70300 , n70526 );
and ( n70588 , n30224 , n70548 );
and ( n70589 , n70587 , n70588 );
xor ( n70590 , n70587 , n70588 );
xor ( n70591 , n70304 , n70524 );
and ( n70592 , n30229 , n70548 );
and ( n70593 , n70591 , n70592 );
xor ( n70594 , n70591 , n70592 );
xor ( n70595 , n70308 , n70522 );
and ( n70596 , n30234 , n70548 );
and ( n70597 , n70595 , n70596 );
xor ( n70598 , n70595 , n70596 );
xor ( n70599 , n70312 , n70520 );
and ( n70600 , n30239 , n70548 );
and ( n70601 , n70599 , n70600 );
xor ( n70602 , n70599 , n70600 );
xor ( n70603 , n70316 , n70518 );
and ( n70604 , n30244 , n70548 );
and ( n70605 , n70603 , n70604 );
xor ( n70606 , n70603 , n70604 );
xor ( n70607 , n70320 , n70516 );
and ( n70608 , n30249 , n70548 );
and ( n70609 , n70607 , n70608 );
xor ( n70610 , n70607 , n70608 );
xor ( n70611 , n70324 , n70514 );
and ( n70612 , n30254 , n70548 );
and ( n70613 , n70611 , n70612 );
xor ( n70614 , n70611 , n70612 );
xor ( n70615 , n70328 , n70512 );
and ( n70616 , n30259 , n70548 );
and ( n70617 , n70615 , n70616 );
xor ( n70618 , n70615 , n70616 );
xor ( n70619 , n70332 , n70510 );
and ( n70620 , n30264 , n70548 );
and ( n70621 , n70619 , n70620 );
xor ( n70622 , n70619 , n70620 );
xor ( n70623 , n70336 , n70508 );
and ( n70624 , n30269 , n70548 );
and ( n70625 , n70623 , n70624 );
xor ( n70626 , n70623 , n70624 );
xor ( n70627 , n70340 , n70506 );
and ( n70628 , n30274 , n70548 );
and ( n70629 , n70627 , n70628 );
xor ( n70630 , n70627 , n70628 );
xor ( n70631 , n70344 , n70504 );
and ( n70632 , n30279 , n70548 );
and ( n70633 , n70631 , n70632 );
xor ( n70634 , n70631 , n70632 );
xor ( n70635 , n70348 , n70502 );
and ( n70636 , n30284 , n70548 );
and ( n70637 , n70635 , n70636 );
xor ( n70638 , n70635 , n70636 );
xor ( n70639 , n70352 , n70500 );
and ( n70640 , n30289 , n70548 );
and ( n70641 , n70639 , n70640 );
xor ( n70642 , n70639 , n70640 );
xor ( n70643 , n70356 , n70498 );
and ( n70644 , n30294 , n70548 );
and ( n70645 , n70643 , n70644 );
xor ( n70646 , n70643 , n70644 );
xor ( n70647 , n70360 , n70496 );
and ( n70648 , n30299 , n70548 );
and ( n70649 , n70647 , n70648 );
xor ( n70650 , n70647 , n70648 );
xor ( n70651 , n70364 , n70494 );
and ( n70652 , n30304 , n70548 );
and ( n70653 , n70651 , n70652 );
xor ( n70654 , n70651 , n70652 );
xor ( n70655 , n70368 , n70492 );
and ( n70656 , n30309 , n70548 );
and ( n70657 , n70655 , n70656 );
xor ( n70658 , n70655 , n70656 );
xor ( n70659 , n70372 , n70490 );
and ( n70660 , n30314 , n70548 );
and ( n70661 , n70659 , n70660 );
xor ( n70662 , n70659 , n70660 );
xor ( n70663 , n70376 , n70488 );
and ( n70664 , n30319 , n70548 );
and ( n70665 , n70663 , n70664 );
xor ( n70666 , n70663 , n70664 );
xor ( n70667 , n70380 , n70486 );
and ( n70668 , n30324 , n70548 );
and ( n70669 , n70667 , n70668 );
xor ( n70670 , n70667 , n70668 );
xor ( n70671 , n70384 , n70484 );
and ( n70672 , n30329 , n70548 );
and ( n70673 , n70671 , n70672 );
xor ( n70674 , n70671 , n70672 );
xor ( n70675 , n70388 , n70482 );
and ( n70676 , n30334 , n70548 );
and ( n70677 , n70675 , n70676 );
xor ( n70678 , n70675 , n70676 );
xor ( n70679 , n70392 , n70480 );
and ( n70680 , n30339 , n70548 );
and ( n70681 , n70679 , n70680 );
xor ( n70682 , n70679 , n70680 );
xor ( n70683 , n70396 , n70478 );
and ( n70684 , n30344 , n70548 );
and ( n70685 , n70683 , n70684 );
xor ( n70686 , n70683 , n70684 );
xor ( n70687 , n70400 , n70476 );
and ( n70688 , n30349 , n70548 );
and ( n70689 , n70687 , n70688 );
xor ( n70690 , n70687 , n70688 );
xor ( n70691 , n70404 , n70474 );
and ( n70692 , n30354 , n70548 );
and ( n70693 , n70691 , n70692 );
xor ( n70694 , n70691 , n70692 );
xor ( n70695 , n70408 , n70472 );
and ( n70696 , n30359 , n70548 );
and ( n70697 , n70695 , n70696 );
xor ( n70698 , n70695 , n70696 );
xor ( n70699 , n70412 , n70470 );
and ( n70700 , n30364 , n70548 );
and ( n70701 , n70699 , n70700 );
xor ( n70702 , n70699 , n70700 );
xor ( n70703 , n70416 , n70468 );
and ( n70704 , n30369 , n70548 );
and ( n70705 , n70703 , n70704 );
xor ( n70706 , n70703 , n70704 );
xor ( n70707 , n70420 , n70466 );
and ( n70708 , n30374 , n70548 );
and ( n70709 , n70707 , n70708 );
xor ( n70710 , n70707 , n70708 );
xor ( n70711 , n70424 , n70464 );
and ( n70712 , n30379 , n70548 );
and ( n70713 , n70711 , n70712 );
xor ( n70714 , n70711 , n70712 );
xor ( n70715 , n70428 , n70462 );
and ( n70716 , n30384 , n70548 );
and ( n70717 , n70715 , n70716 );
xor ( n70718 , n70715 , n70716 );
xor ( n70719 , n70432 , n70460 );
and ( n70720 , n30389 , n70548 );
and ( n70721 , n70719 , n70720 );
xor ( n70722 , n70719 , n70720 );
xor ( n70723 , n70436 , n70458 );
and ( n70724 , n30394 , n70548 );
and ( n70725 , n70723 , n70724 );
xor ( n70726 , n70723 , n70724 );
xor ( n70727 , n70440 , n70456 );
and ( n70728 , n30399 , n70548 );
and ( n70729 , n70727 , n70728 );
xor ( n70730 , n70727 , n70728 );
xor ( n70731 , n70444 , n70454 );
and ( n70732 , n30404 , n70548 );
and ( n70733 , n70731 , n70732 );
xor ( n70734 , n70731 , n70732 );
xor ( n70735 , n70448 , n70452 );
and ( n70736 , n30409 , n70548 );
and ( n70737 , n70735 , n70736 );
buf ( n70738 , n70737 );
and ( n70739 , n70734 , n70738 );
or ( n70740 , n70733 , n70739 );
and ( n70741 , n70730 , n70740 );
or ( n70742 , n70729 , n70741 );
and ( n70743 , n70726 , n70742 );
or ( n70744 , n70725 , n70743 );
and ( n70745 , n70722 , n70744 );
or ( n70746 , n70721 , n70745 );
and ( n70747 , n70718 , n70746 );
or ( n70748 , n70717 , n70747 );
and ( n70749 , n70714 , n70748 );
or ( n70750 , n70713 , n70749 );
and ( n70751 , n70710 , n70750 );
or ( n70752 , n70709 , n70751 );
and ( n70753 , n70706 , n70752 );
or ( n70754 , n70705 , n70753 );
and ( n70755 , n70702 , n70754 );
or ( n70756 , n70701 , n70755 );
and ( n70757 , n70698 , n70756 );
or ( n70758 , n70697 , n70757 );
and ( n70759 , n70694 , n70758 );
or ( n70760 , n70693 , n70759 );
and ( n70761 , n70690 , n70760 );
or ( n70762 , n70689 , n70761 );
and ( n70763 , n70686 , n70762 );
or ( n70764 , n70685 , n70763 );
and ( n70765 , n70682 , n70764 );
or ( n70766 , n70681 , n70765 );
and ( n70767 , n70678 , n70766 );
or ( n70768 , n70677 , n70767 );
and ( n70769 , n70674 , n70768 );
or ( n70770 , n70673 , n70769 );
and ( n70771 , n70670 , n70770 );
or ( n70772 , n70669 , n70771 );
and ( n70773 , n70666 , n70772 );
or ( n70774 , n70665 , n70773 );
and ( n70775 , n70662 , n70774 );
or ( n70776 , n70661 , n70775 );
and ( n70777 , n70658 , n70776 );
or ( n70778 , n70657 , n70777 );
and ( n70779 , n70654 , n70778 );
or ( n70780 , n70653 , n70779 );
and ( n70781 , n70650 , n70780 );
or ( n70782 , n70649 , n70781 );
and ( n70783 , n70646 , n70782 );
or ( n70784 , n70645 , n70783 );
and ( n70785 , n70642 , n70784 );
or ( n70786 , n70641 , n70785 );
and ( n70787 , n70638 , n70786 );
or ( n70788 , n70637 , n70787 );
and ( n70789 , n70634 , n70788 );
or ( n70790 , n70633 , n70789 );
and ( n70791 , n70630 , n70790 );
or ( n70792 , n70629 , n70791 );
and ( n70793 , n70626 , n70792 );
or ( n70794 , n70625 , n70793 );
and ( n70795 , n70622 , n70794 );
or ( n70796 , n70621 , n70795 );
and ( n70797 , n70618 , n70796 );
or ( n70798 , n70617 , n70797 );
and ( n70799 , n70614 , n70798 );
or ( n70800 , n70613 , n70799 );
and ( n70801 , n70610 , n70800 );
or ( n70802 , n70609 , n70801 );
and ( n70803 , n70606 , n70802 );
or ( n70804 , n70605 , n70803 );
and ( n70805 , n70602 , n70804 );
or ( n70806 , n70601 , n70805 );
and ( n70807 , n70598 , n70806 );
or ( n70808 , n70597 , n70807 );
and ( n70809 , n70594 , n70808 );
or ( n70810 , n70593 , n70809 );
and ( n70811 , n70590 , n70810 );
or ( n70812 , n70589 , n70811 );
and ( n70813 , n70586 , n70812 );
or ( n70814 , n70585 , n70813 );
and ( n70815 , n70582 , n70814 );
or ( n70816 , n70581 , n70815 );
and ( n70817 , n70578 , n70816 );
or ( n70818 , n70577 , n70817 );
and ( n70819 , n70574 , n70818 );
or ( n70820 , n70573 , n70819 );
and ( n70821 , n70570 , n70820 );
or ( n70822 , n70569 , n70821 );
and ( n70823 , n70566 , n70822 );
or ( n70824 , n70565 , n70823 );
and ( n70825 , n70562 , n70824 );
or ( n70826 , n70561 , n70825 );
and ( n70827 , n70558 , n70826 );
or ( n70828 , n70557 , n70827 );
and ( n70829 , n70554 , n70828 );
or ( n70830 , n70553 , n70829 );
xor ( n70831 , n70550 , n70830 );
buf ( n70832 , n17946 );
and ( n70833 , n30179 , n70832 );
xor ( n70834 , n70831 , n70833 );
xor ( n70835 , n70554 , n70828 );
and ( n70836 , n30184 , n70832 );
and ( n70837 , n70835 , n70836 );
xor ( n70838 , n70835 , n70836 );
xor ( n70839 , n70558 , n70826 );
and ( n70840 , n30189 , n70832 );
and ( n70841 , n70839 , n70840 );
xor ( n70842 , n70839 , n70840 );
xor ( n70843 , n70562 , n70824 );
and ( n70844 , n30194 , n70832 );
and ( n70845 , n70843 , n70844 );
xor ( n70846 , n70843 , n70844 );
xor ( n70847 , n70566 , n70822 );
and ( n70848 , n30199 , n70832 );
and ( n70849 , n70847 , n70848 );
xor ( n70850 , n70847 , n70848 );
xor ( n70851 , n70570 , n70820 );
and ( n70852 , n30204 , n70832 );
and ( n70853 , n70851 , n70852 );
xor ( n70854 , n70851 , n70852 );
xor ( n70855 , n70574 , n70818 );
and ( n70856 , n30209 , n70832 );
and ( n70857 , n70855 , n70856 );
xor ( n70858 , n70855 , n70856 );
xor ( n70859 , n70578 , n70816 );
and ( n70860 , n30214 , n70832 );
and ( n70861 , n70859 , n70860 );
xor ( n70862 , n70859 , n70860 );
xor ( n70863 , n70582 , n70814 );
and ( n70864 , n30219 , n70832 );
and ( n70865 , n70863 , n70864 );
xor ( n70866 , n70863 , n70864 );
xor ( n70867 , n70586 , n70812 );
and ( n70868 , n30224 , n70832 );
and ( n70869 , n70867 , n70868 );
xor ( n70870 , n70867 , n70868 );
xor ( n70871 , n70590 , n70810 );
and ( n70872 , n30229 , n70832 );
and ( n70873 , n70871 , n70872 );
xor ( n70874 , n70871 , n70872 );
xor ( n70875 , n70594 , n70808 );
and ( n70876 , n30234 , n70832 );
and ( n70877 , n70875 , n70876 );
xor ( n70878 , n70875 , n70876 );
xor ( n70879 , n70598 , n70806 );
and ( n70880 , n30239 , n70832 );
and ( n70881 , n70879 , n70880 );
xor ( n70882 , n70879 , n70880 );
xor ( n70883 , n70602 , n70804 );
and ( n70884 , n30244 , n70832 );
and ( n70885 , n70883 , n70884 );
xor ( n70886 , n70883 , n70884 );
xor ( n70887 , n70606 , n70802 );
and ( n70888 , n30249 , n70832 );
and ( n70889 , n70887 , n70888 );
xor ( n70890 , n70887 , n70888 );
xor ( n70891 , n70610 , n70800 );
and ( n70892 , n30254 , n70832 );
and ( n70893 , n70891 , n70892 );
xor ( n70894 , n70891 , n70892 );
xor ( n70895 , n70614 , n70798 );
and ( n70896 , n30259 , n70832 );
and ( n70897 , n70895 , n70896 );
xor ( n70898 , n70895 , n70896 );
xor ( n70899 , n70618 , n70796 );
and ( n70900 , n30264 , n70832 );
and ( n70901 , n70899 , n70900 );
xor ( n70902 , n70899 , n70900 );
xor ( n70903 , n70622 , n70794 );
and ( n70904 , n30269 , n70832 );
and ( n70905 , n70903 , n70904 );
xor ( n70906 , n70903 , n70904 );
xor ( n70907 , n70626 , n70792 );
and ( n70908 , n30274 , n70832 );
and ( n70909 , n70907 , n70908 );
xor ( n70910 , n70907 , n70908 );
xor ( n70911 , n70630 , n70790 );
and ( n70912 , n30279 , n70832 );
and ( n70913 , n70911 , n70912 );
xor ( n70914 , n70911 , n70912 );
xor ( n70915 , n70634 , n70788 );
and ( n70916 , n30284 , n70832 );
and ( n70917 , n70915 , n70916 );
xor ( n70918 , n70915 , n70916 );
xor ( n70919 , n70638 , n70786 );
and ( n70920 , n30289 , n70832 );
and ( n70921 , n70919 , n70920 );
xor ( n70922 , n70919 , n70920 );
xor ( n70923 , n70642 , n70784 );
and ( n70924 , n30294 , n70832 );
and ( n70925 , n70923 , n70924 );
xor ( n70926 , n70923 , n70924 );
xor ( n70927 , n70646 , n70782 );
and ( n70928 , n30299 , n70832 );
and ( n70929 , n70927 , n70928 );
xor ( n70930 , n70927 , n70928 );
xor ( n70931 , n70650 , n70780 );
and ( n70932 , n30304 , n70832 );
and ( n70933 , n70931 , n70932 );
xor ( n70934 , n70931 , n70932 );
xor ( n70935 , n70654 , n70778 );
and ( n70936 , n30309 , n70832 );
and ( n70937 , n70935 , n70936 );
xor ( n70938 , n70935 , n70936 );
xor ( n70939 , n70658 , n70776 );
and ( n70940 , n30314 , n70832 );
and ( n70941 , n70939 , n70940 );
xor ( n70942 , n70939 , n70940 );
xor ( n70943 , n70662 , n70774 );
and ( n70944 , n30319 , n70832 );
and ( n70945 , n70943 , n70944 );
xor ( n70946 , n70943 , n70944 );
xor ( n70947 , n70666 , n70772 );
and ( n70948 , n30324 , n70832 );
and ( n70949 , n70947 , n70948 );
xor ( n70950 , n70947 , n70948 );
xor ( n70951 , n70670 , n70770 );
and ( n70952 , n30329 , n70832 );
and ( n70953 , n70951 , n70952 );
xor ( n70954 , n70951 , n70952 );
xor ( n70955 , n70674 , n70768 );
and ( n70956 , n30334 , n70832 );
and ( n70957 , n70955 , n70956 );
xor ( n70958 , n70955 , n70956 );
xor ( n70959 , n70678 , n70766 );
and ( n70960 , n30339 , n70832 );
and ( n70961 , n70959 , n70960 );
xor ( n70962 , n70959 , n70960 );
xor ( n70963 , n70682 , n70764 );
and ( n70964 , n30344 , n70832 );
and ( n70965 , n70963 , n70964 );
xor ( n70966 , n70963 , n70964 );
xor ( n70967 , n70686 , n70762 );
and ( n70968 , n30349 , n70832 );
and ( n70969 , n70967 , n70968 );
xor ( n70970 , n70967 , n70968 );
xor ( n70971 , n70690 , n70760 );
and ( n70972 , n30354 , n70832 );
and ( n70973 , n70971 , n70972 );
xor ( n70974 , n70971 , n70972 );
xor ( n70975 , n70694 , n70758 );
and ( n70976 , n30359 , n70832 );
and ( n70977 , n70975 , n70976 );
xor ( n70978 , n70975 , n70976 );
xor ( n70979 , n70698 , n70756 );
and ( n70980 , n30364 , n70832 );
and ( n70981 , n70979 , n70980 );
xor ( n70982 , n70979 , n70980 );
xor ( n70983 , n70702 , n70754 );
and ( n70984 , n30369 , n70832 );
and ( n70985 , n70983 , n70984 );
xor ( n70986 , n70983 , n70984 );
xor ( n70987 , n70706 , n70752 );
and ( n70988 , n30374 , n70832 );
and ( n70989 , n70987 , n70988 );
xor ( n70990 , n70987 , n70988 );
xor ( n70991 , n70710 , n70750 );
and ( n70992 , n30379 , n70832 );
and ( n70993 , n70991 , n70992 );
xor ( n70994 , n70991 , n70992 );
xor ( n70995 , n70714 , n70748 );
and ( n70996 , n30384 , n70832 );
and ( n70997 , n70995 , n70996 );
xor ( n70998 , n70995 , n70996 );
xor ( n70999 , n70718 , n70746 );
and ( n71000 , n30389 , n70832 );
and ( n71001 , n70999 , n71000 );
xor ( n71002 , n70999 , n71000 );
xor ( n71003 , n70722 , n70744 );
and ( n71004 , n30394 , n70832 );
and ( n71005 , n71003 , n71004 );
xor ( n71006 , n71003 , n71004 );
xor ( n71007 , n70726 , n70742 );
and ( n71008 , n30399 , n70832 );
and ( n71009 , n71007 , n71008 );
xor ( n71010 , n71007 , n71008 );
xor ( n71011 , n70730 , n70740 );
and ( n71012 , n30404 , n70832 );
and ( n71013 , n71011 , n71012 );
xor ( n71014 , n71011 , n71012 );
xor ( n71015 , n70734 , n70738 );
and ( n71016 , n30409 , n70832 );
and ( n71017 , n71015 , n71016 );
buf ( n71018 , n71017 );
and ( n71019 , n71014 , n71018 );
or ( n71020 , n71013 , n71019 );
and ( n71021 , n71010 , n71020 );
or ( n71022 , n71009 , n71021 );
and ( n71023 , n71006 , n71022 );
or ( n71024 , n71005 , n71023 );
and ( n71025 , n71002 , n71024 );
or ( n71026 , n71001 , n71025 );
and ( n71027 , n70998 , n71026 );
or ( n71028 , n70997 , n71027 );
and ( n71029 , n70994 , n71028 );
or ( n71030 , n70993 , n71029 );
and ( n71031 , n70990 , n71030 );
or ( n71032 , n70989 , n71031 );
and ( n71033 , n70986 , n71032 );
or ( n71034 , n70985 , n71033 );
and ( n71035 , n70982 , n71034 );
or ( n71036 , n70981 , n71035 );
and ( n71037 , n70978 , n71036 );
or ( n71038 , n70977 , n71037 );
and ( n71039 , n70974 , n71038 );
or ( n71040 , n70973 , n71039 );
and ( n71041 , n70970 , n71040 );
or ( n71042 , n70969 , n71041 );
and ( n71043 , n70966 , n71042 );
or ( n71044 , n70965 , n71043 );
and ( n71045 , n70962 , n71044 );
or ( n71046 , n70961 , n71045 );
and ( n71047 , n70958 , n71046 );
or ( n71048 , n70957 , n71047 );
and ( n71049 , n70954 , n71048 );
or ( n71050 , n70953 , n71049 );
and ( n71051 , n70950 , n71050 );
or ( n71052 , n70949 , n71051 );
and ( n71053 , n70946 , n71052 );
or ( n71054 , n70945 , n71053 );
and ( n71055 , n70942 , n71054 );
or ( n71056 , n70941 , n71055 );
and ( n71057 , n70938 , n71056 );
or ( n71058 , n70937 , n71057 );
and ( n71059 , n70934 , n71058 );
or ( n71060 , n70933 , n71059 );
and ( n71061 , n70930 , n71060 );
or ( n71062 , n70929 , n71061 );
and ( n71063 , n70926 , n71062 );
or ( n71064 , n70925 , n71063 );
and ( n71065 , n70922 , n71064 );
or ( n71066 , n70921 , n71065 );
and ( n71067 , n70918 , n71066 );
or ( n71068 , n70917 , n71067 );
and ( n71069 , n70914 , n71068 );
or ( n71070 , n70913 , n71069 );
and ( n71071 , n70910 , n71070 );
or ( n71072 , n70909 , n71071 );
and ( n71073 , n70906 , n71072 );
or ( n71074 , n70905 , n71073 );
and ( n71075 , n70902 , n71074 );
or ( n71076 , n70901 , n71075 );
and ( n71077 , n70898 , n71076 );
or ( n71078 , n70897 , n71077 );
and ( n71079 , n70894 , n71078 );
or ( n71080 , n70893 , n71079 );
and ( n71081 , n70890 , n71080 );
or ( n71082 , n70889 , n71081 );
and ( n71083 , n70886 , n71082 );
or ( n71084 , n70885 , n71083 );
and ( n71085 , n70882 , n71084 );
or ( n71086 , n70881 , n71085 );
and ( n71087 , n70878 , n71086 );
or ( n71088 , n70877 , n71087 );
and ( n71089 , n70874 , n71088 );
or ( n71090 , n70873 , n71089 );
and ( n71091 , n70870 , n71090 );
or ( n71092 , n70869 , n71091 );
and ( n71093 , n70866 , n71092 );
or ( n71094 , n70865 , n71093 );
and ( n71095 , n70862 , n71094 );
or ( n71096 , n70861 , n71095 );
and ( n71097 , n70858 , n71096 );
or ( n71098 , n70857 , n71097 );
and ( n71099 , n70854 , n71098 );
or ( n71100 , n70853 , n71099 );
and ( n71101 , n70850 , n71100 );
or ( n71102 , n70849 , n71101 );
and ( n71103 , n70846 , n71102 );
or ( n71104 , n70845 , n71103 );
and ( n71105 , n70842 , n71104 );
or ( n71106 , n70841 , n71105 );
and ( n71107 , n70838 , n71106 );
or ( n71108 , n70837 , n71107 );
xor ( n71109 , n70834 , n71108 );
buf ( n71110 , n17944 );
and ( n71111 , n30184 , n71110 );
xor ( n71112 , n71109 , n71111 );
xor ( n71113 , n70838 , n71106 );
and ( n71114 , n30189 , n71110 );
and ( n71115 , n71113 , n71114 );
xor ( n71116 , n71113 , n71114 );
xor ( n71117 , n70842 , n71104 );
and ( n71118 , n30194 , n71110 );
and ( n71119 , n71117 , n71118 );
xor ( n71120 , n71117 , n71118 );
xor ( n71121 , n70846 , n71102 );
and ( n71122 , n30199 , n71110 );
and ( n71123 , n71121 , n71122 );
xor ( n71124 , n71121 , n71122 );
xor ( n71125 , n70850 , n71100 );
and ( n71126 , n30204 , n71110 );
and ( n71127 , n71125 , n71126 );
xor ( n71128 , n71125 , n71126 );
xor ( n71129 , n70854 , n71098 );
and ( n71130 , n30209 , n71110 );
and ( n71131 , n71129 , n71130 );
xor ( n71132 , n71129 , n71130 );
xor ( n71133 , n70858 , n71096 );
and ( n71134 , n30214 , n71110 );
and ( n71135 , n71133 , n71134 );
xor ( n71136 , n71133 , n71134 );
xor ( n71137 , n70862 , n71094 );
and ( n71138 , n30219 , n71110 );
and ( n71139 , n71137 , n71138 );
xor ( n71140 , n71137 , n71138 );
xor ( n71141 , n70866 , n71092 );
and ( n71142 , n30224 , n71110 );
and ( n71143 , n71141 , n71142 );
xor ( n71144 , n71141 , n71142 );
xor ( n71145 , n70870 , n71090 );
and ( n71146 , n30229 , n71110 );
and ( n71147 , n71145 , n71146 );
xor ( n71148 , n71145 , n71146 );
xor ( n71149 , n70874 , n71088 );
and ( n71150 , n30234 , n71110 );
and ( n71151 , n71149 , n71150 );
xor ( n71152 , n71149 , n71150 );
xor ( n71153 , n70878 , n71086 );
and ( n71154 , n30239 , n71110 );
and ( n71155 , n71153 , n71154 );
xor ( n71156 , n71153 , n71154 );
xor ( n71157 , n70882 , n71084 );
and ( n71158 , n30244 , n71110 );
and ( n71159 , n71157 , n71158 );
xor ( n71160 , n71157 , n71158 );
xor ( n71161 , n70886 , n71082 );
and ( n71162 , n30249 , n71110 );
and ( n71163 , n71161 , n71162 );
xor ( n71164 , n71161 , n71162 );
xor ( n71165 , n70890 , n71080 );
and ( n71166 , n30254 , n71110 );
and ( n71167 , n71165 , n71166 );
xor ( n71168 , n71165 , n71166 );
xor ( n71169 , n70894 , n71078 );
and ( n71170 , n30259 , n71110 );
and ( n71171 , n71169 , n71170 );
xor ( n71172 , n71169 , n71170 );
xor ( n71173 , n70898 , n71076 );
and ( n71174 , n30264 , n71110 );
and ( n71175 , n71173 , n71174 );
xor ( n71176 , n71173 , n71174 );
xor ( n71177 , n70902 , n71074 );
and ( n71178 , n30269 , n71110 );
and ( n71179 , n71177 , n71178 );
xor ( n71180 , n71177 , n71178 );
xor ( n71181 , n70906 , n71072 );
and ( n71182 , n30274 , n71110 );
and ( n71183 , n71181 , n71182 );
xor ( n71184 , n71181 , n71182 );
xor ( n71185 , n70910 , n71070 );
and ( n71186 , n30279 , n71110 );
and ( n71187 , n71185 , n71186 );
xor ( n71188 , n71185 , n71186 );
xor ( n71189 , n70914 , n71068 );
and ( n71190 , n30284 , n71110 );
and ( n71191 , n71189 , n71190 );
xor ( n71192 , n71189 , n71190 );
xor ( n71193 , n70918 , n71066 );
and ( n71194 , n30289 , n71110 );
and ( n71195 , n71193 , n71194 );
xor ( n71196 , n71193 , n71194 );
xor ( n71197 , n70922 , n71064 );
and ( n71198 , n30294 , n71110 );
and ( n71199 , n71197 , n71198 );
xor ( n71200 , n71197 , n71198 );
xor ( n71201 , n70926 , n71062 );
and ( n71202 , n30299 , n71110 );
and ( n71203 , n71201 , n71202 );
xor ( n71204 , n71201 , n71202 );
xor ( n71205 , n70930 , n71060 );
and ( n71206 , n30304 , n71110 );
and ( n71207 , n71205 , n71206 );
xor ( n71208 , n71205 , n71206 );
xor ( n71209 , n70934 , n71058 );
and ( n71210 , n30309 , n71110 );
and ( n71211 , n71209 , n71210 );
xor ( n71212 , n71209 , n71210 );
xor ( n71213 , n70938 , n71056 );
and ( n71214 , n30314 , n71110 );
and ( n71215 , n71213 , n71214 );
xor ( n71216 , n71213 , n71214 );
xor ( n71217 , n70942 , n71054 );
and ( n71218 , n30319 , n71110 );
and ( n71219 , n71217 , n71218 );
xor ( n71220 , n71217 , n71218 );
xor ( n71221 , n70946 , n71052 );
and ( n71222 , n30324 , n71110 );
and ( n71223 , n71221 , n71222 );
xor ( n71224 , n71221 , n71222 );
xor ( n71225 , n70950 , n71050 );
and ( n71226 , n30329 , n71110 );
and ( n71227 , n71225 , n71226 );
xor ( n71228 , n71225 , n71226 );
xor ( n71229 , n70954 , n71048 );
and ( n71230 , n30334 , n71110 );
and ( n71231 , n71229 , n71230 );
xor ( n71232 , n71229 , n71230 );
xor ( n71233 , n70958 , n71046 );
and ( n71234 , n30339 , n71110 );
and ( n71235 , n71233 , n71234 );
xor ( n71236 , n71233 , n71234 );
xor ( n71237 , n70962 , n71044 );
and ( n71238 , n30344 , n71110 );
and ( n71239 , n71237 , n71238 );
xor ( n71240 , n71237 , n71238 );
xor ( n71241 , n70966 , n71042 );
and ( n71242 , n30349 , n71110 );
and ( n71243 , n71241 , n71242 );
xor ( n71244 , n71241 , n71242 );
xor ( n71245 , n70970 , n71040 );
and ( n71246 , n30354 , n71110 );
and ( n71247 , n71245 , n71246 );
xor ( n71248 , n71245 , n71246 );
xor ( n71249 , n70974 , n71038 );
and ( n71250 , n30359 , n71110 );
and ( n71251 , n71249 , n71250 );
xor ( n71252 , n71249 , n71250 );
xor ( n71253 , n70978 , n71036 );
and ( n71254 , n30364 , n71110 );
and ( n71255 , n71253 , n71254 );
xor ( n71256 , n71253 , n71254 );
xor ( n71257 , n70982 , n71034 );
and ( n71258 , n30369 , n71110 );
and ( n71259 , n71257 , n71258 );
xor ( n71260 , n71257 , n71258 );
xor ( n71261 , n70986 , n71032 );
and ( n71262 , n30374 , n71110 );
and ( n71263 , n71261 , n71262 );
xor ( n71264 , n71261 , n71262 );
xor ( n71265 , n70990 , n71030 );
and ( n71266 , n30379 , n71110 );
and ( n71267 , n71265 , n71266 );
xor ( n71268 , n71265 , n71266 );
xor ( n71269 , n70994 , n71028 );
and ( n71270 , n30384 , n71110 );
and ( n71271 , n71269 , n71270 );
xor ( n71272 , n71269 , n71270 );
xor ( n71273 , n70998 , n71026 );
and ( n71274 , n30389 , n71110 );
and ( n71275 , n71273 , n71274 );
xor ( n71276 , n71273 , n71274 );
xor ( n71277 , n71002 , n71024 );
and ( n71278 , n30394 , n71110 );
and ( n71279 , n71277 , n71278 );
xor ( n71280 , n71277 , n71278 );
xor ( n71281 , n71006 , n71022 );
and ( n71282 , n30399 , n71110 );
and ( n71283 , n71281 , n71282 );
xor ( n71284 , n71281 , n71282 );
xor ( n71285 , n71010 , n71020 );
and ( n71286 , n30404 , n71110 );
and ( n71287 , n71285 , n71286 );
xor ( n71288 , n71285 , n71286 );
xor ( n71289 , n71014 , n71018 );
and ( n71290 , n30409 , n71110 );
and ( n71291 , n71289 , n71290 );
buf ( n71292 , n71291 );
and ( n71293 , n71288 , n71292 );
or ( n71294 , n71287 , n71293 );
and ( n71295 , n71284 , n71294 );
or ( n71296 , n71283 , n71295 );
and ( n71297 , n71280 , n71296 );
or ( n71298 , n71279 , n71297 );
and ( n71299 , n71276 , n71298 );
or ( n71300 , n71275 , n71299 );
and ( n71301 , n71272 , n71300 );
or ( n71302 , n71271 , n71301 );
and ( n71303 , n71268 , n71302 );
or ( n71304 , n71267 , n71303 );
and ( n71305 , n71264 , n71304 );
or ( n71306 , n71263 , n71305 );
and ( n71307 , n71260 , n71306 );
or ( n71308 , n71259 , n71307 );
and ( n71309 , n71256 , n71308 );
or ( n71310 , n71255 , n71309 );
and ( n71311 , n71252 , n71310 );
or ( n71312 , n71251 , n71311 );
and ( n71313 , n71248 , n71312 );
or ( n71314 , n71247 , n71313 );
and ( n71315 , n71244 , n71314 );
or ( n71316 , n71243 , n71315 );
and ( n71317 , n71240 , n71316 );
or ( n71318 , n71239 , n71317 );
and ( n71319 , n71236 , n71318 );
or ( n71320 , n71235 , n71319 );
and ( n71321 , n71232 , n71320 );
or ( n71322 , n71231 , n71321 );
and ( n71323 , n71228 , n71322 );
or ( n71324 , n71227 , n71323 );
and ( n71325 , n71224 , n71324 );
or ( n71326 , n71223 , n71325 );
and ( n71327 , n71220 , n71326 );
or ( n71328 , n71219 , n71327 );
and ( n71329 , n71216 , n71328 );
or ( n71330 , n71215 , n71329 );
and ( n71331 , n71212 , n71330 );
or ( n71332 , n71211 , n71331 );
and ( n71333 , n71208 , n71332 );
or ( n71334 , n71207 , n71333 );
and ( n71335 , n71204 , n71334 );
or ( n71336 , n71203 , n71335 );
and ( n71337 , n71200 , n71336 );
or ( n71338 , n71199 , n71337 );
and ( n71339 , n71196 , n71338 );
or ( n71340 , n71195 , n71339 );
and ( n71341 , n71192 , n71340 );
or ( n71342 , n71191 , n71341 );
and ( n71343 , n71188 , n71342 );
or ( n71344 , n71187 , n71343 );
and ( n71345 , n71184 , n71344 );
or ( n71346 , n71183 , n71345 );
and ( n71347 , n71180 , n71346 );
or ( n71348 , n71179 , n71347 );
and ( n71349 , n71176 , n71348 );
or ( n71350 , n71175 , n71349 );
and ( n71351 , n71172 , n71350 );
or ( n71352 , n71171 , n71351 );
and ( n71353 , n71168 , n71352 );
or ( n71354 , n71167 , n71353 );
and ( n71355 , n71164 , n71354 );
or ( n71356 , n71163 , n71355 );
and ( n71357 , n71160 , n71356 );
or ( n71358 , n71159 , n71357 );
and ( n71359 , n71156 , n71358 );
or ( n71360 , n71155 , n71359 );
and ( n71361 , n71152 , n71360 );
or ( n71362 , n71151 , n71361 );
and ( n71363 , n71148 , n71362 );
or ( n71364 , n71147 , n71363 );
and ( n71365 , n71144 , n71364 );
or ( n71366 , n71143 , n71365 );
and ( n71367 , n71140 , n71366 );
or ( n71368 , n71139 , n71367 );
and ( n71369 , n71136 , n71368 );
or ( n71370 , n71135 , n71369 );
and ( n71371 , n71132 , n71370 );
or ( n71372 , n71131 , n71371 );
and ( n71373 , n71128 , n71372 );
or ( n71374 , n71127 , n71373 );
and ( n71375 , n71124 , n71374 );
or ( n71376 , n71123 , n71375 );
and ( n71377 , n71120 , n71376 );
or ( n71378 , n71119 , n71377 );
and ( n71379 , n71116 , n71378 );
or ( n71380 , n71115 , n71379 );
xor ( n71381 , n71112 , n71380 );
buf ( n71382 , n17942 );
and ( n71383 , n30189 , n71382 );
xor ( n71384 , n71381 , n71383 );
xor ( n71385 , n71116 , n71378 );
and ( n71386 , n30194 , n71382 );
and ( n71387 , n71385 , n71386 );
xor ( n71388 , n71385 , n71386 );
xor ( n71389 , n71120 , n71376 );
and ( n71390 , n30199 , n71382 );
and ( n71391 , n71389 , n71390 );
xor ( n71392 , n71389 , n71390 );
xor ( n71393 , n71124 , n71374 );
and ( n71394 , n30204 , n71382 );
and ( n71395 , n71393 , n71394 );
xor ( n71396 , n71393 , n71394 );
xor ( n71397 , n71128 , n71372 );
and ( n71398 , n30209 , n71382 );
and ( n71399 , n71397 , n71398 );
xor ( n71400 , n71397 , n71398 );
xor ( n71401 , n71132 , n71370 );
and ( n71402 , n30214 , n71382 );
and ( n71403 , n71401 , n71402 );
xor ( n71404 , n71401 , n71402 );
xor ( n71405 , n71136 , n71368 );
and ( n71406 , n30219 , n71382 );
and ( n71407 , n71405 , n71406 );
xor ( n71408 , n71405 , n71406 );
xor ( n71409 , n71140 , n71366 );
and ( n71410 , n30224 , n71382 );
and ( n71411 , n71409 , n71410 );
xor ( n71412 , n71409 , n71410 );
xor ( n71413 , n71144 , n71364 );
and ( n71414 , n30229 , n71382 );
and ( n71415 , n71413 , n71414 );
xor ( n71416 , n71413 , n71414 );
xor ( n71417 , n71148 , n71362 );
and ( n71418 , n30234 , n71382 );
and ( n71419 , n71417 , n71418 );
xor ( n71420 , n71417 , n71418 );
xor ( n71421 , n71152 , n71360 );
and ( n71422 , n30239 , n71382 );
and ( n71423 , n71421 , n71422 );
xor ( n71424 , n71421 , n71422 );
xor ( n71425 , n71156 , n71358 );
and ( n71426 , n30244 , n71382 );
and ( n71427 , n71425 , n71426 );
xor ( n71428 , n71425 , n71426 );
xor ( n71429 , n71160 , n71356 );
and ( n71430 , n30249 , n71382 );
and ( n71431 , n71429 , n71430 );
xor ( n71432 , n71429 , n71430 );
xor ( n71433 , n71164 , n71354 );
and ( n71434 , n30254 , n71382 );
and ( n71435 , n71433 , n71434 );
xor ( n71436 , n71433 , n71434 );
xor ( n71437 , n71168 , n71352 );
and ( n71438 , n30259 , n71382 );
and ( n71439 , n71437 , n71438 );
xor ( n71440 , n71437 , n71438 );
xor ( n71441 , n71172 , n71350 );
and ( n71442 , n30264 , n71382 );
and ( n71443 , n71441 , n71442 );
xor ( n71444 , n71441 , n71442 );
xor ( n71445 , n71176 , n71348 );
and ( n71446 , n30269 , n71382 );
and ( n71447 , n71445 , n71446 );
xor ( n71448 , n71445 , n71446 );
xor ( n71449 , n71180 , n71346 );
and ( n71450 , n30274 , n71382 );
and ( n71451 , n71449 , n71450 );
xor ( n71452 , n71449 , n71450 );
xor ( n71453 , n71184 , n71344 );
and ( n71454 , n30279 , n71382 );
and ( n71455 , n71453 , n71454 );
xor ( n71456 , n71453 , n71454 );
xor ( n71457 , n71188 , n71342 );
and ( n71458 , n30284 , n71382 );
and ( n71459 , n71457 , n71458 );
xor ( n71460 , n71457 , n71458 );
xor ( n71461 , n71192 , n71340 );
and ( n71462 , n30289 , n71382 );
and ( n71463 , n71461 , n71462 );
xor ( n71464 , n71461 , n71462 );
xor ( n71465 , n71196 , n71338 );
and ( n71466 , n30294 , n71382 );
and ( n71467 , n71465 , n71466 );
xor ( n71468 , n71465 , n71466 );
xor ( n71469 , n71200 , n71336 );
and ( n71470 , n30299 , n71382 );
and ( n71471 , n71469 , n71470 );
xor ( n71472 , n71469 , n71470 );
xor ( n71473 , n71204 , n71334 );
and ( n71474 , n30304 , n71382 );
and ( n71475 , n71473 , n71474 );
xor ( n71476 , n71473 , n71474 );
xor ( n71477 , n71208 , n71332 );
and ( n71478 , n30309 , n71382 );
and ( n71479 , n71477 , n71478 );
xor ( n71480 , n71477 , n71478 );
xor ( n71481 , n71212 , n71330 );
and ( n71482 , n30314 , n71382 );
and ( n71483 , n71481 , n71482 );
xor ( n71484 , n71481 , n71482 );
xor ( n71485 , n71216 , n71328 );
and ( n71486 , n30319 , n71382 );
and ( n71487 , n71485 , n71486 );
xor ( n71488 , n71485 , n71486 );
xor ( n71489 , n71220 , n71326 );
and ( n71490 , n30324 , n71382 );
and ( n71491 , n71489 , n71490 );
xor ( n71492 , n71489 , n71490 );
xor ( n71493 , n71224 , n71324 );
and ( n71494 , n30329 , n71382 );
and ( n71495 , n71493 , n71494 );
xor ( n71496 , n71493 , n71494 );
xor ( n71497 , n71228 , n71322 );
and ( n71498 , n30334 , n71382 );
and ( n71499 , n71497 , n71498 );
xor ( n71500 , n71497 , n71498 );
xor ( n71501 , n71232 , n71320 );
and ( n71502 , n30339 , n71382 );
and ( n71503 , n71501 , n71502 );
xor ( n71504 , n71501 , n71502 );
xor ( n71505 , n71236 , n71318 );
and ( n71506 , n30344 , n71382 );
and ( n71507 , n71505 , n71506 );
xor ( n71508 , n71505 , n71506 );
xor ( n71509 , n71240 , n71316 );
and ( n71510 , n30349 , n71382 );
and ( n71511 , n71509 , n71510 );
xor ( n71512 , n71509 , n71510 );
xor ( n71513 , n71244 , n71314 );
and ( n71514 , n30354 , n71382 );
and ( n71515 , n71513 , n71514 );
xor ( n71516 , n71513 , n71514 );
xor ( n71517 , n71248 , n71312 );
and ( n71518 , n30359 , n71382 );
and ( n71519 , n71517 , n71518 );
xor ( n71520 , n71517 , n71518 );
xor ( n71521 , n71252 , n71310 );
and ( n71522 , n30364 , n71382 );
and ( n71523 , n71521 , n71522 );
xor ( n71524 , n71521 , n71522 );
xor ( n71525 , n71256 , n71308 );
and ( n71526 , n30369 , n71382 );
and ( n71527 , n71525 , n71526 );
xor ( n71528 , n71525 , n71526 );
xor ( n71529 , n71260 , n71306 );
and ( n71530 , n30374 , n71382 );
and ( n71531 , n71529 , n71530 );
xor ( n71532 , n71529 , n71530 );
xor ( n71533 , n71264 , n71304 );
and ( n71534 , n30379 , n71382 );
and ( n71535 , n71533 , n71534 );
xor ( n71536 , n71533 , n71534 );
xor ( n71537 , n71268 , n71302 );
and ( n71538 , n30384 , n71382 );
and ( n71539 , n71537 , n71538 );
xor ( n71540 , n71537 , n71538 );
xor ( n71541 , n71272 , n71300 );
and ( n71542 , n30389 , n71382 );
and ( n71543 , n71541 , n71542 );
xor ( n71544 , n71541 , n71542 );
xor ( n71545 , n71276 , n71298 );
and ( n71546 , n30394 , n71382 );
and ( n71547 , n71545 , n71546 );
xor ( n71548 , n71545 , n71546 );
xor ( n71549 , n71280 , n71296 );
and ( n71550 , n30399 , n71382 );
and ( n71551 , n71549 , n71550 );
xor ( n71552 , n71549 , n71550 );
xor ( n71553 , n71284 , n71294 );
and ( n71554 , n30404 , n71382 );
and ( n71555 , n71553 , n71554 );
xor ( n71556 , n71553 , n71554 );
xor ( n71557 , n71288 , n71292 );
and ( n71558 , n30409 , n71382 );
and ( n71559 , n71557 , n71558 );
buf ( n71560 , n71559 );
and ( n71561 , n71556 , n71560 );
or ( n71562 , n71555 , n71561 );
and ( n71563 , n71552 , n71562 );
or ( n71564 , n71551 , n71563 );
and ( n71565 , n71548 , n71564 );
or ( n71566 , n71547 , n71565 );
and ( n71567 , n71544 , n71566 );
or ( n71568 , n71543 , n71567 );
and ( n71569 , n71540 , n71568 );
or ( n71570 , n71539 , n71569 );
and ( n71571 , n71536 , n71570 );
or ( n71572 , n71535 , n71571 );
and ( n71573 , n71532 , n71572 );
or ( n71574 , n71531 , n71573 );
and ( n71575 , n71528 , n71574 );
or ( n71576 , n71527 , n71575 );
and ( n71577 , n71524 , n71576 );
or ( n71578 , n71523 , n71577 );
and ( n71579 , n71520 , n71578 );
or ( n71580 , n71519 , n71579 );
and ( n71581 , n71516 , n71580 );
or ( n71582 , n71515 , n71581 );
and ( n71583 , n71512 , n71582 );
or ( n71584 , n71511 , n71583 );
and ( n71585 , n71508 , n71584 );
or ( n71586 , n71507 , n71585 );
and ( n71587 , n71504 , n71586 );
or ( n71588 , n71503 , n71587 );
and ( n71589 , n71500 , n71588 );
or ( n71590 , n71499 , n71589 );
and ( n71591 , n71496 , n71590 );
or ( n71592 , n71495 , n71591 );
and ( n71593 , n71492 , n71592 );
or ( n71594 , n71491 , n71593 );
and ( n71595 , n71488 , n71594 );
or ( n71596 , n71487 , n71595 );
and ( n71597 , n71484 , n71596 );
or ( n71598 , n71483 , n71597 );
and ( n71599 , n71480 , n71598 );
or ( n71600 , n71479 , n71599 );
and ( n71601 , n71476 , n71600 );
or ( n71602 , n71475 , n71601 );
and ( n71603 , n71472 , n71602 );
or ( n71604 , n71471 , n71603 );
and ( n71605 , n71468 , n71604 );
or ( n71606 , n71467 , n71605 );
and ( n71607 , n71464 , n71606 );
or ( n71608 , n71463 , n71607 );
and ( n71609 , n71460 , n71608 );
or ( n71610 , n71459 , n71609 );
and ( n71611 , n71456 , n71610 );
or ( n71612 , n71455 , n71611 );
and ( n71613 , n71452 , n71612 );
or ( n71614 , n71451 , n71613 );
and ( n71615 , n71448 , n71614 );
or ( n71616 , n71447 , n71615 );
and ( n71617 , n71444 , n71616 );
or ( n71618 , n71443 , n71617 );
and ( n71619 , n71440 , n71618 );
or ( n71620 , n71439 , n71619 );
and ( n71621 , n71436 , n71620 );
or ( n71622 , n71435 , n71621 );
and ( n71623 , n71432 , n71622 );
or ( n71624 , n71431 , n71623 );
and ( n71625 , n71428 , n71624 );
or ( n71626 , n71427 , n71625 );
and ( n71627 , n71424 , n71626 );
or ( n71628 , n71423 , n71627 );
and ( n71629 , n71420 , n71628 );
or ( n71630 , n71419 , n71629 );
and ( n71631 , n71416 , n71630 );
or ( n71632 , n71415 , n71631 );
and ( n71633 , n71412 , n71632 );
or ( n71634 , n71411 , n71633 );
and ( n71635 , n71408 , n71634 );
or ( n71636 , n71407 , n71635 );
and ( n71637 , n71404 , n71636 );
or ( n71638 , n71403 , n71637 );
and ( n71639 , n71400 , n71638 );
or ( n71640 , n71399 , n71639 );
and ( n71641 , n71396 , n71640 );
or ( n71642 , n71395 , n71641 );
and ( n71643 , n71392 , n71642 );
or ( n71644 , n71391 , n71643 );
and ( n71645 , n71388 , n71644 );
or ( n71646 , n71387 , n71645 );
xor ( n71647 , n71384 , n71646 );
buf ( n71648 , n17940 );
and ( n71649 , n30194 , n71648 );
xor ( n71650 , n71647 , n71649 );
xor ( n71651 , n71388 , n71644 );
and ( n71652 , n30199 , n71648 );
and ( n71653 , n71651 , n71652 );
xor ( n71654 , n71651 , n71652 );
xor ( n71655 , n71392 , n71642 );
and ( n71656 , n30204 , n71648 );
and ( n71657 , n71655 , n71656 );
xor ( n71658 , n71655 , n71656 );
xor ( n71659 , n71396 , n71640 );
and ( n71660 , n30209 , n71648 );
and ( n71661 , n71659 , n71660 );
xor ( n71662 , n71659 , n71660 );
xor ( n71663 , n71400 , n71638 );
and ( n71664 , n30214 , n71648 );
and ( n71665 , n71663 , n71664 );
xor ( n71666 , n71663 , n71664 );
xor ( n71667 , n71404 , n71636 );
and ( n71668 , n30219 , n71648 );
and ( n71669 , n71667 , n71668 );
xor ( n71670 , n71667 , n71668 );
xor ( n71671 , n71408 , n71634 );
and ( n71672 , n30224 , n71648 );
and ( n71673 , n71671 , n71672 );
xor ( n71674 , n71671 , n71672 );
xor ( n71675 , n71412 , n71632 );
and ( n71676 , n30229 , n71648 );
and ( n71677 , n71675 , n71676 );
xor ( n71678 , n71675 , n71676 );
xor ( n71679 , n71416 , n71630 );
and ( n71680 , n30234 , n71648 );
and ( n71681 , n71679 , n71680 );
xor ( n71682 , n71679 , n71680 );
xor ( n71683 , n71420 , n71628 );
and ( n71684 , n30239 , n71648 );
and ( n71685 , n71683 , n71684 );
xor ( n71686 , n71683 , n71684 );
xor ( n71687 , n71424 , n71626 );
and ( n71688 , n30244 , n71648 );
and ( n71689 , n71687 , n71688 );
xor ( n71690 , n71687 , n71688 );
xor ( n71691 , n71428 , n71624 );
and ( n71692 , n30249 , n71648 );
and ( n71693 , n71691 , n71692 );
xor ( n71694 , n71691 , n71692 );
xor ( n71695 , n71432 , n71622 );
and ( n71696 , n30254 , n71648 );
and ( n71697 , n71695 , n71696 );
xor ( n71698 , n71695 , n71696 );
xor ( n71699 , n71436 , n71620 );
and ( n71700 , n30259 , n71648 );
and ( n71701 , n71699 , n71700 );
xor ( n71702 , n71699 , n71700 );
xor ( n71703 , n71440 , n71618 );
and ( n71704 , n30264 , n71648 );
and ( n71705 , n71703 , n71704 );
xor ( n71706 , n71703 , n71704 );
xor ( n71707 , n71444 , n71616 );
and ( n71708 , n30269 , n71648 );
and ( n71709 , n71707 , n71708 );
xor ( n71710 , n71707 , n71708 );
xor ( n71711 , n71448 , n71614 );
and ( n71712 , n30274 , n71648 );
and ( n71713 , n71711 , n71712 );
xor ( n71714 , n71711 , n71712 );
xor ( n71715 , n71452 , n71612 );
and ( n71716 , n30279 , n71648 );
and ( n71717 , n71715 , n71716 );
xor ( n71718 , n71715 , n71716 );
xor ( n71719 , n71456 , n71610 );
and ( n71720 , n30284 , n71648 );
and ( n71721 , n71719 , n71720 );
xor ( n71722 , n71719 , n71720 );
xor ( n71723 , n71460 , n71608 );
and ( n71724 , n30289 , n71648 );
and ( n71725 , n71723 , n71724 );
xor ( n71726 , n71723 , n71724 );
xor ( n71727 , n71464 , n71606 );
and ( n71728 , n30294 , n71648 );
and ( n71729 , n71727 , n71728 );
xor ( n71730 , n71727 , n71728 );
xor ( n71731 , n71468 , n71604 );
and ( n71732 , n30299 , n71648 );
and ( n71733 , n71731 , n71732 );
xor ( n71734 , n71731 , n71732 );
xor ( n71735 , n71472 , n71602 );
and ( n71736 , n30304 , n71648 );
and ( n71737 , n71735 , n71736 );
xor ( n71738 , n71735 , n71736 );
xor ( n71739 , n71476 , n71600 );
and ( n71740 , n30309 , n71648 );
and ( n71741 , n71739 , n71740 );
xor ( n71742 , n71739 , n71740 );
xor ( n71743 , n71480 , n71598 );
and ( n71744 , n30314 , n71648 );
and ( n71745 , n71743 , n71744 );
xor ( n71746 , n71743 , n71744 );
xor ( n71747 , n71484 , n71596 );
and ( n71748 , n30319 , n71648 );
and ( n71749 , n71747 , n71748 );
xor ( n71750 , n71747 , n71748 );
xor ( n71751 , n71488 , n71594 );
and ( n71752 , n30324 , n71648 );
and ( n71753 , n71751 , n71752 );
xor ( n71754 , n71751 , n71752 );
xor ( n71755 , n71492 , n71592 );
and ( n71756 , n30329 , n71648 );
and ( n71757 , n71755 , n71756 );
xor ( n71758 , n71755 , n71756 );
xor ( n71759 , n71496 , n71590 );
and ( n71760 , n30334 , n71648 );
and ( n71761 , n71759 , n71760 );
xor ( n71762 , n71759 , n71760 );
xor ( n71763 , n71500 , n71588 );
and ( n71764 , n30339 , n71648 );
and ( n71765 , n71763 , n71764 );
xor ( n71766 , n71763 , n71764 );
xor ( n71767 , n71504 , n71586 );
and ( n71768 , n30344 , n71648 );
and ( n71769 , n71767 , n71768 );
xor ( n71770 , n71767 , n71768 );
xor ( n71771 , n71508 , n71584 );
and ( n71772 , n30349 , n71648 );
and ( n71773 , n71771 , n71772 );
xor ( n71774 , n71771 , n71772 );
xor ( n71775 , n71512 , n71582 );
and ( n71776 , n30354 , n71648 );
and ( n71777 , n71775 , n71776 );
xor ( n71778 , n71775 , n71776 );
xor ( n71779 , n71516 , n71580 );
and ( n71780 , n30359 , n71648 );
and ( n71781 , n71779 , n71780 );
xor ( n71782 , n71779 , n71780 );
xor ( n71783 , n71520 , n71578 );
and ( n71784 , n30364 , n71648 );
and ( n71785 , n71783 , n71784 );
xor ( n71786 , n71783 , n71784 );
xor ( n71787 , n71524 , n71576 );
and ( n71788 , n30369 , n71648 );
and ( n71789 , n71787 , n71788 );
xor ( n71790 , n71787 , n71788 );
xor ( n71791 , n71528 , n71574 );
and ( n71792 , n30374 , n71648 );
and ( n71793 , n71791 , n71792 );
xor ( n71794 , n71791 , n71792 );
xor ( n71795 , n71532 , n71572 );
and ( n71796 , n30379 , n71648 );
and ( n71797 , n71795 , n71796 );
xor ( n71798 , n71795 , n71796 );
xor ( n71799 , n71536 , n71570 );
and ( n71800 , n30384 , n71648 );
and ( n71801 , n71799 , n71800 );
xor ( n71802 , n71799 , n71800 );
xor ( n71803 , n71540 , n71568 );
and ( n71804 , n30389 , n71648 );
and ( n71805 , n71803 , n71804 );
xor ( n71806 , n71803 , n71804 );
xor ( n71807 , n71544 , n71566 );
and ( n71808 , n30394 , n71648 );
and ( n71809 , n71807 , n71808 );
xor ( n71810 , n71807 , n71808 );
xor ( n71811 , n71548 , n71564 );
and ( n71812 , n30399 , n71648 );
and ( n71813 , n71811 , n71812 );
xor ( n71814 , n71811 , n71812 );
xor ( n71815 , n71552 , n71562 );
and ( n71816 , n30404 , n71648 );
and ( n71817 , n71815 , n71816 );
xor ( n71818 , n71815 , n71816 );
xor ( n71819 , n71556 , n71560 );
and ( n71820 , n30409 , n71648 );
and ( n71821 , n71819 , n71820 );
buf ( n71822 , n71821 );
and ( n71823 , n71818 , n71822 );
or ( n71824 , n71817 , n71823 );
and ( n71825 , n71814 , n71824 );
or ( n71826 , n71813 , n71825 );
and ( n71827 , n71810 , n71826 );
or ( n71828 , n71809 , n71827 );
and ( n71829 , n71806 , n71828 );
or ( n71830 , n71805 , n71829 );
and ( n71831 , n71802 , n71830 );
or ( n71832 , n71801 , n71831 );
and ( n71833 , n71798 , n71832 );
or ( n71834 , n71797 , n71833 );
and ( n71835 , n71794 , n71834 );
or ( n71836 , n71793 , n71835 );
and ( n71837 , n71790 , n71836 );
or ( n71838 , n71789 , n71837 );
and ( n71839 , n71786 , n71838 );
or ( n71840 , n71785 , n71839 );
and ( n71841 , n71782 , n71840 );
or ( n71842 , n71781 , n71841 );
and ( n71843 , n71778 , n71842 );
or ( n71844 , n71777 , n71843 );
and ( n71845 , n71774 , n71844 );
or ( n71846 , n71773 , n71845 );
and ( n71847 , n71770 , n71846 );
or ( n71848 , n71769 , n71847 );
and ( n71849 , n71766 , n71848 );
or ( n71850 , n71765 , n71849 );
and ( n71851 , n71762 , n71850 );
or ( n71852 , n71761 , n71851 );
and ( n71853 , n71758 , n71852 );
or ( n71854 , n71757 , n71853 );
and ( n71855 , n71754 , n71854 );
or ( n71856 , n71753 , n71855 );
and ( n71857 , n71750 , n71856 );
or ( n71858 , n71749 , n71857 );
and ( n71859 , n71746 , n71858 );
or ( n71860 , n71745 , n71859 );
and ( n71861 , n71742 , n71860 );
or ( n71862 , n71741 , n71861 );
and ( n71863 , n71738 , n71862 );
or ( n71864 , n71737 , n71863 );
and ( n71865 , n71734 , n71864 );
or ( n71866 , n71733 , n71865 );
and ( n71867 , n71730 , n71866 );
or ( n71868 , n71729 , n71867 );
and ( n71869 , n71726 , n71868 );
or ( n71870 , n71725 , n71869 );
and ( n71871 , n71722 , n71870 );
or ( n71872 , n71721 , n71871 );
and ( n71873 , n71718 , n71872 );
or ( n71874 , n71717 , n71873 );
and ( n71875 , n71714 , n71874 );
or ( n71876 , n71713 , n71875 );
and ( n71877 , n71710 , n71876 );
or ( n71878 , n71709 , n71877 );
and ( n71879 , n71706 , n71878 );
or ( n71880 , n71705 , n71879 );
and ( n71881 , n71702 , n71880 );
or ( n71882 , n71701 , n71881 );
and ( n71883 , n71698 , n71882 );
or ( n71884 , n71697 , n71883 );
and ( n71885 , n71694 , n71884 );
or ( n71886 , n71693 , n71885 );
and ( n71887 , n71690 , n71886 );
or ( n71888 , n71689 , n71887 );
and ( n71889 , n71686 , n71888 );
or ( n71890 , n71685 , n71889 );
and ( n71891 , n71682 , n71890 );
or ( n71892 , n71681 , n71891 );
and ( n71893 , n71678 , n71892 );
or ( n71894 , n71677 , n71893 );
and ( n71895 , n71674 , n71894 );
or ( n71896 , n71673 , n71895 );
and ( n71897 , n71670 , n71896 );
or ( n71898 , n71669 , n71897 );
and ( n71899 , n71666 , n71898 );
or ( n71900 , n71665 , n71899 );
and ( n71901 , n71662 , n71900 );
or ( n71902 , n71661 , n71901 );
and ( n71903 , n71658 , n71902 );
or ( n71904 , n71657 , n71903 );
and ( n71905 , n71654 , n71904 );
or ( n71906 , n71653 , n71905 );
xor ( n71907 , n71650 , n71906 );
buf ( n71908 , n17938 );
and ( n71909 , n30199 , n71908 );
xor ( n71910 , n71907 , n71909 );
xor ( n71911 , n71654 , n71904 );
and ( n71912 , n30204 , n71908 );
and ( n71913 , n71911 , n71912 );
xor ( n71914 , n71911 , n71912 );
xor ( n71915 , n71658 , n71902 );
and ( n71916 , n30209 , n71908 );
and ( n71917 , n71915 , n71916 );
xor ( n71918 , n71915 , n71916 );
xor ( n71919 , n71662 , n71900 );
and ( n71920 , n30214 , n71908 );
and ( n71921 , n71919 , n71920 );
xor ( n71922 , n71919 , n71920 );
xor ( n71923 , n71666 , n71898 );
and ( n71924 , n30219 , n71908 );
and ( n71925 , n71923 , n71924 );
xor ( n71926 , n71923 , n71924 );
xor ( n71927 , n71670 , n71896 );
and ( n71928 , n30224 , n71908 );
and ( n71929 , n71927 , n71928 );
xor ( n71930 , n71927 , n71928 );
xor ( n71931 , n71674 , n71894 );
and ( n71932 , n30229 , n71908 );
and ( n71933 , n71931 , n71932 );
xor ( n71934 , n71931 , n71932 );
xor ( n71935 , n71678 , n71892 );
and ( n71936 , n30234 , n71908 );
and ( n71937 , n71935 , n71936 );
xor ( n71938 , n71935 , n71936 );
xor ( n71939 , n71682 , n71890 );
and ( n71940 , n30239 , n71908 );
and ( n71941 , n71939 , n71940 );
xor ( n71942 , n71939 , n71940 );
xor ( n71943 , n71686 , n71888 );
and ( n71944 , n30244 , n71908 );
and ( n71945 , n71943 , n71944 );
xor ( n71946 , n71943 , n71944 );
xor ( n71947 , n71690 , n71886 );
and ( n71948 , n30249 , n71908 );
and ( n71949 , n71947 , n71948 );
xor ( n71950 , n71947 , n71948 );
xor ( n71951 , n71694 , n71884 );
and ( n71952 , n30254 , n71908 );
and ( n71953 , n71951 , n71952 );
xor ( n71954 , n71951 , n71952 );
xor ( n71955 , n71698 , n71882 );
and ( n71956 , n30259 , n71908 );
and ( n71957 , n71955 , n71956 );
xor ( n71958 , n71955 , n71956 );
xor ( n71959 , n71702 , n71880 );
and ( n71960 , n30264 , n71908 );
and ( n71961 , n71959 , n71960 );
xor ( n71962 , n71959 , n71960 );
xor ( n71963 , n71706 , n71878 );
and ( n71964 , n30269 , n71908 );
and ( n71965 , n71963 , n71964 );
xor ( n71966 , n71963 , n71964 );
xor ( n71967 , n71710 , n71876 );
and ( n71968 , n30274 , n71908 );
and ( n71969 , n71967 , n71968 );
xor ( n71970 , n71967 , n71968 );
xor ( n71971 , n71714 , n71874 );
and ( n71972 , n30279 , n71908 );
and ( n71973 , n71971 , n71972 );
xor ( n71974 , n71971 , n71972 );
xor ( n71975 , n71718 , n71872 );
and ( n71976 , n30284 , n71908 );
and ( n71977 , n71975 , n71976 );
xor ( n71978 , n71975 , n71976 );
xor ( n71979 , n71722 , n71870 );
and ( n71980 , n30289 , n71908 );
and ( n71981 , n71979 , n71980 );
xor ( n71982 , n71979 , n71980 );
xor ( n71983 , n71726 , n71868 );
and ( n71984 , n30294 , n71908 );
and ( n71985 , n71983 , n71984 );
xor ( n71986 , n71983 , n71984 );
xor ( n71987 , n71730 , n71866 );
and ( n71988 , n30299 , n71908 );
and ( n71989 , n71987 , n71988 );
xor ( n71990 , n71987 , n71988 );
xor ( n71991 , n71734 , n71864 );
and ( n71992 , n30304 , n71908 );
and ( n71993 , n71991 , n71992 );
xor ( n71994 , n71991 , n71992 );
xor ( n71995 , n71738 , n71862 );
and ( n71996 , n30309 , n71908 );
and ( n71997 , n71995 , n71996 );
xor ( n71998 , n71995 , n71996 );
xor ( n71999 , n71742 , n71860 );
and ( n72000 , n30314 , n71908 );
and ( n72001 , n71999 , n72000 );
xor ( n72002 , n71999 , n72000 );
xor ( n72003 , n71746 , n71858 );
and ( n72004 , n30319 , n71908 );
and ( n72005 , n72003 , n72004 );
xor ( n72006 , n72003 , n72004 );
xor ( n72007 , n71750 , n71856 );
and ( n72008 , n30324 , n71908 );
and ( n72009 , n72007 , n72008 );
xor ( n72010 , n72007 , n72008 );
xor ( n72011 , n71754 , n71854 );
and ( n72012 , n30329 , n71908 );
and ( n72013 , n72011 , n72012 );
xor ( n72014 , n72011 , n72012 );
xor ( n72015 , n71758 , n71852 );
and ( n72016 , n30334 , n71908 );
and ( n72017 , n72015 , n72016 );
xor ( n72018 , n72015 , n72016 );
xor ( n72019 , n71762 , n71850 );
and ( n72020 , n30339 , n71908 );
and ( n72021 , n72019 , n72020 );
xor ( n72022 , n72019 , n72020 );
xor ( n72023 , n71766 , n71848 );
and ( n72024 , n30344 , n71908 );
and ( n72025 , n72023 , n72024 );
xor ( n72026 , n72023 , n72024 );
xor ( n72027 , n71770 , n71846 );
and ( n72028 , n30349 , n71908 );
and ( n72029 , n72027 , n72028 );
xor ( n72030 , n72027 , n72028 );
xor ( n72031 , n71774 , n71844 );
and ( n72032 , n30354 , n71908 );
and ( n72033 , n72031 , n72032 );
xor ( n72034 , n72031 , n72032 );
xor ( n72035 , n71778 , n71842 );
and ( n72036 , n30359 , n71908 );
and ( n72037 , n72035 , n72036 );
xor ( n72038 , n72035 , n72036 );
xor ( n72039 , n71782 , n71840 );
and ( n72040 , n30364 , n71908 );
and ( n72041 , n72039 , n72040 );
xor ( n72042 , n72039 , n72040 );
xor ( n72043 , n71786 , n71838 );
and ( n72044 , n30369 , n71908 );
and ( n72045 , n72043 , n72044 );
xor ( n72046 , n72043 , n72044 );
xor ( n72047 , n71790 , n71836 );
and ( n72048 , n30374 , n71908 );
and ( n72049 , n72047 , n72048 );
xor ( n72050 , n72047 , n72048 );
xor ( n72051 , n71794 , n71834 );
and ( n72052 , n30379 , n71908 );
and ( n72053 , n72051 , n72052 );
xor ( n72054 , n72051 , n72052 );
xor ( n72055 , n71798 , n71832 );
and ( n72056 , n30384 , n71908 );
and ( n72057 , n72055 , n72056 );
xor ( n72058 , n72055 , n72056 );
xor ( n72059 , n71802 , n71830 );
and ( n72060 , n30389 , n71908 );
and ( n72061 , n72059 , n72060 );
xor ( n72062 , n72059 , n72060 );
xor ( n72063 , n71806 , n71828 );
and ( n72064 , n30394 , n71908 );
and ( n72065 , n72063 , n72064 );
xor ( n72066 , n72063 , n72064 );
xor ( n72067 , n71810 , n71826 );
and ( n72068 , n30399 , n71908 );
and ( n72069 , n72067 , n72068 );
xor ( n72070 , n72067 , n72068 );
xor ( n72071 , n71814 , n71824 );
and ( n72072 , n30404 , n71908 );
and ( n72073 , n72071 , n72072 );
xor ( n72074 , n72071 , n72072 );
xor ( n72075 , n71818 , n71822 );
and ( n72076 , n30409 , n71908 );
and ( n72077 , n72075 , n72076 );
buf ( n72078 , n72077 );
and ( n72079 , n72074 , n72078 );
or ( n72080 , n72073 , n72079 );
and ( n72081 , n72070 , n72080 );
or ( n72082 , n72069 , n72081 );
and ( n72083 , n72066 , n72082 );
or ( n72084 , n72065 , n72083 );
and ( n72085 , n72062 , n72084 );
or ( n72086 , n72061 , n72085 );
and ( n72087 , n72058 , n72086 );
or ( n72088 , n72057 , n72087 );
and ( n72089 , n72054 , n72088 );
or ( n72090 , n72053 , n72089 );
and ( n72091 , n72050 , n72090 );
or ( n72092 , n72049 , n72091 );
and ( n72093 , n72046 , n72092 );
or ( n72094 , n72045 , n72093 );
and ( n72095 , n72042 , n72094 );
or ( n72096 , n72041 , n72095 );
and ( n72097 , n72038 , n72096 );
or ( n72098 , n72037 , n72097 );
and ( n72099 , n72034 , n72098 );
or ( n72100 , n72033 , n72099 );
and ( n72101 , n72030 , n72100 );
or ( n72102 , n72029 , n72101 );
and ( n72103 , n72026 , n72102 );
or ( n72104 , n72025 , n72103 );
and ( n72105 , n72022 , n72104 );
or ( n72106 , n72021 , n72105 );
and ( n72107 , n72018 , n72106 );
or ( n72108 , n72017 , n72107 );
and ( n72109 , n72014 , n72108 );
or ( n72110 , n72013 , n72109 );
and ( n72111 , n72010 , n72110 );
or ( n72112 , n72009 , n72111 );
and ( n72113 , n72006 , n72112 );
or ( n72114 , n72005 , n72113 );
and ( n72115 , n72002 , n72114 );
or ( n72116 , n72001 , n72115 );
and ( n72117 , n71998 , n72116 );
or ( n72118 , n71997 , n72117 );
and ( n72119 , n71994 , n72118 );
or ( n72120 , n71993 , n72119 );
and ( n72121 , n71990 , n72120 );
or ( n72122 , n71989 , n72121 );
and ( n72123 , n71986 , n72122 );
or ( n72124 , n71985 , n72123 );
and ( n72125 , n71982 , n72124 );
or ( n72126 , n71981 , n72125 );
and ( n72127 , n71978 , n72126 );
or ( n72128 , n71977 , n72127 );
and ( n72129 , n71974 , n72128 );
or ( n72130 , n71973 , n72129 );
and ( n72131 , n71970 , n72130 );
or ( n72132 , n71969 , n72131 );
and ( n72133 , n71966 , n72132 );
or ( n72134 , n71965 , n72133 );
and ( n72135 , n71962 , n72134 );
or ( n72136 , n71961 , n72135 );
and ( n72137 , n71958 , n72136 );
or ( n72138 , n71957 , n72137 );
and ( n72139 , n71954 , n72138 );
or ( n72140 , n71953 , n72139 );
and ( n72141 , n71950 , n72140 );
or ( n72142 , n71949 , n72141 );
and ( n72143 , n71946 , n72142 );
or ( n72144 , n71945 , n72143 );
and ( n72145 , n71942 , n72144 );
or ( n72146 , n71941 , n72145 );
and ( n72147 , n71938 , n72146 );
or ( n72148 , n71937 , n72147 );
and ( n72149 , n71934 , n72148 );
or ( n72150 , n71933 , n72149 );
and ( n72151 , n71930 , n72150 );
or ( n72152 , n71929 , n72151 );
and ( n72153 , n71926 , n72152 );
or ( n72154 , n71925 , n72153 );
and ( n72155 , n71922 , n72154 );
or ( n72156 , n71921 , n72155 );
and ( n72157 , n71918 , n72156 );
or ( n72158 , n71917 , n72157 );
and ( n72159 , n71914 , n72158 );
or ( n72160 , n71913 , n72159 );
xor ( n72161 , n71910 , n72160 );
buf ( n72162 , n17936 );
and ( n72163 , n30204 , n72162 );
xor ( n72164 , n72161 , n72163 );
xor ( n72165 , n71914 , n72158 );
and ( n72166 , n30209 , n72162 );
and ( n72167 , n72165 , n72166 );
xor ( n72168 , n72165 , n72166 );
xor ( n72169 , n71918 , n72156 );
and ( n72170 , n30214 , n72162 );
and ( n72171 , n72169 , n72170 );
xor ( n72172 , n72169 , n72170 );
xor ( n72173 , n71922 , n72154 );
and ( n72174 , n30219 , n72162 );
and ( n72175 , n72173 , n72174 );
xor ( n72176 , n72173 , n72174 );
xor ( n72177 , n71926 , n72152 );
and ( n72178 , n30224 , n72162 );
and ( n72179 , n72177 , n72178 );
xor ( n72180 , n72177 , n72178 );
xor ( n72181 , n71930 , n72150 );
and ( n72182 , n30229 , n72162 );
and ( n72183 , n72181 , n72182 );
xor ( n72184 , n72181 , n72182 );
xor ( n72185 , n71934 , n72148 );
and ( n72186 , n30234 , n72162 );
and ( n72187 , n72185 , n72186 );
xor ( n72188 , n72185 , n72186 );
xor ( n72189 , n71938 , n72146 );
and ( n72190 , n30239 , n72162 );
and ( n72191 , n72189 , n72190 );
xor ( n72192 , n72189 , n72190 );
xor ( n72193 , n71942 , n72144 );
and ( n72194 , n30244 , n72162 );
and ( n72195 , n72193 , n72194 );
xor ( n72196 , n72193 , n72194 );
xor ( n72197 , n71946 , n72142 );
and ( n72198 , n30249 , n72162 );
and ( n72199 , n72197 , n72198 );
xor ( n72200 , n72197 , n72198 );
xor ( n72201 , n71950 , n72140 );
and ( n72202 , n30254 , n72162 );
and ( n72203 , n72201 , n72202 );
xor ( n72204 , n72201 , n72202 );
xor ( n72205 , n71954 , n72138 );
and ( n72206 , n30259 , n72162 );
and ( n72207 , n72205 , n72206 );
xor ( n72208 , n72205 , n72206 );
xor ( n72209 , n71958 , n72136 );
and ( n72210 , n30264 , n72162 );
and ( n72211 , n72209 , n72210 );
xor ( n72212 , n72209 , n72210 );
xor ( n72213 , n71962 , n72134 );
and ( n72214 , n30269 , n72162 );
and ( n72215 , n72213 , n72214 );
xor ( n72216 , n72213 , n72214 );
xor ( n72217 , n71966 , n72132 );
and ( n72218 , n30274 , n72162 );
and ( n72219 , n72217 , n72218 );
xor ( n72220 , n72217 , n72218 );
xor ( n72221 , n71970 , n72130 );
and ( n72222 , n30279 , n72162 );
and ( n72223 , n72221 , n72222 );
xor ( n72224 , n72221 , n72222 );
xor ( n72225 , n71974 , n72128 );
and ( n72226 , n30284 , n72162 );
and ( n72227 , n72225 , n72226 );
xor ( n72228 , n72225 , n72226 );
xor ( n72229 , n71978 , n72126 );
and ( n72230 , n30289 , n72162 );
and ( n72231 , n72229 , n72230 );
xor ( n72232 , n72229 , n72230 );
xor ( n72233 , n71982 , n72124 );
and ( n72234 , n30294 , n72162 );
and ( n72235 , n72233 , n72234 );
xor ( n72236 , n72233 , n72234 );
xor ( n72237 , n71986 , n72122 );
and ( n72238 , n30299 , n72162 );
and ( n72239 , n72237 , n72238 );
xor ( n72240 , n72237 , n72238 );
xor ( n72241 , n71990 , n72120 );
and ( n72242 , n30304 , n72162 );
and ( n72243 , n72241 , n72242 );
xor ( n72244 , n72241 , n72242 );
xor ( n72245 , n71994 , n72118 );
and ( n72246 , n30309 , n72162 );
and ( n72247 , n72245 , n72246 );
xor ( n72248 , n72245 , n72246 );
xor ( n72249 , n71998 , n72116 );
and ( n72250 , n30314 , n72162 );
and ( n72251 , n72249 , n72250 );
xor ( n72252 , n72249 , n72250 );
xor ( n72253 , n72002 , n72114 );
and ( n72254 , n30319 , n72162 );
and ( n72255 , n72253 , n72254 );
xor ( n72256 , n72253 , n72254 );
xor ( n72257 , n72006 , n72112 );
and ( n72258 , n30324 , n72162 );
and ( n72259 , n72257 , n72258 );
xor ( n72260 , n72257 , n72258 );
xor ( n72261 , n72010 , n72110 );
and ( n72262 , n30329 , n72162 );
and ( n72263 , n72261 , n72262 );
xor ( n72264 , n72261 , n72262 );
xor ( n72265 , n72014 , n72108 );
and ( n72266 , n30334 , n72162 );
and ( n72267 , n72265 , n72266 );
xor ( n72268 , n72265 , n72266 );
xor ( n72269 , n72018 , n72106 );
and ( n72270 , n30339 , n72162 );
and ( n72271 , n72269 , n72270 );
xor ( n72272 , n72269 , n72270 );
xor ( n72273 , n72022 , n72104 );
and ( n72274 , n30344 , n72162 );
and ( n72275 , n72273 , n72274 );
xor ( n72276 , n72273 , n72274 );
xor ( n72277 , n72026 , n72102 );
and ( n72278 , n30349 , n72162 );
and ( n72279 , n72277 , n72278 );
xor ( n72280 , n72277 , n72278 );
xor ( n72281 , n72030 , n72100 );
and ( n72282 , n30354 , n72162 );
and ( n72283 , n72281 , n72282 );
xor ( n72284 , n72281 , n72282 );
xor ( n72285 , n72034 , n72098 );
and ( n72286 , n30359 , n72162 );
and ( n72287 , n72285 , n72286 );
xor ( n72288 , n72285 , n72286 );
xor ( n72289 , n72038 , n72096 );
and ( n72290 , n30364 , n72162 );
and ( n72291 , n72289 , n72290 );
xor ( n72292 , n72289 , n72290 );
xor ( n72293 , n72042 , n72094 );
and ( n72294 , n30369 , n72162 );
and ( n72295 , n72293 , n72294 );
xor ( n72296 , n72293 , n72294 );
xor ( n72297 , n72046 , n72092 );
and ( n72298 , n30374 , n72162 );
and ( n72299 , n72297 , n72298 );
xor ( n72300 , n72297 , n72298 );
xor ( n72301 , n72050 , n72090 );
and ( n72302 , n30379 , n72162 );
and ( n72303 , n72301 , n72302 );
xor ( n72304 , n72301 , n72302 );
xor ( n72305 , n72054 , n72088 );
and ( n72306 , n30384 , n72162 );
and ( n72307 , n72305 , n72306 );
xor ( n72308 , n72305 , n72306 );
xor ( n72309 , n72058 , n72086 );
and ( n72310 , n30389 , n72162 );
and ( n72311 , n72309 , n72310 );
xor ( n72312 , n72309 , n72310 );
xor ( n72313 , n72062 , n72084 );
and ( n72314 , n30394 , n72162 );
and ( n72315 , n72313 , n72314 );
xor ( n72316 , n72313 , n72314 );
xor ( n72317 , n72066 , n72082 );
and ( n72318 , n30399 , n72162 );
and ( n72319 , n72317 , n72318 );
xor ( n72320 , n72317 , n72318 );
xor ( n72321 , n72070 , n72080 );
and ( n72322 , n30404 , n72162 );
and ( n72323 , n72321 , n72322 );
xor ( n72324 , n72321 , n72322 );
xor ( n72325 , n72074 , n72078 );
and ( n72326 , n30409 , n72162 );
and ( n72327 , n72325 , n72326 );
buf ( n72328 , n72327 );
and ( n72329 , n72324 , n72328 );
or ( n72330 , n72323 , n72329 );
and ( n72331 , n72320 , n72330 );
or ( n72332 , n72319 , n72331 );
and ( n72333 , n72316 , n72332 );
or ( n72334 , n72315 , n72333 );
and ( n72335 , n72312 , n72334 );
or ( n72336 , n72311 , n72335 );
and ( n72337 , n72308 , n72336 );
or ( n72338 , n72307 , n72337 );
and ( n72339 , n72304 , n72338 );
or ( n72340 , n72303 , n72339 );
and ( n72341 , n72300 , n72340 );
or ( n72342 , n72299 , n72341 );
and ( n72343 , n72296 , n72342 );
or ( n72344 , n72295 , n72343 );
and ( n72345 , n72292 , n72344 );
or ( n72346 , n72291 , n72345 );
and ( n72347 , n72288 , n72346 );
or ( n72348 , n72287 , n72347 );
and ( n72349 , n72284 , n72348 );
or ( n72350 , n72283 , n72349 );
and ( n72351 , n72280 , n72350 );
or ( n72352 , n72279 , n72351 );
and ( n72353 , n72276 , n72352 );
or ( n72354 , n72275 , n72353 );
and ( n72355 , n72272 , n72354 );
or ( n72356 , n72271 , n72355 );
and ( n72357 , n72268 , n72356 );
or ( n72358 , n72267 , n72357 );
and ( n72359 , n72264 , n72358 );
or ( n72360 , n72263 , n72359 );
and ( n72361 , n72260 , n72360 );
or ( n72362 , n72259 , n72361 );
and ( n72363 , n72256 , n72362 );
or ( n72364 , n72255 , n72363 );
and ( n72365 , n72252 , n72364 );
or ( n72366 , n72251 , n72365 );
and ( n72367 , n72248 , n72366 );
or ( n72368 , n72247 , n72367 );
and ( n72369 , n72244 , n72368 );
or ( n72370 , n72243 , n72369 );
and ( n72371 , n72240 , n72370 );
or ( n72372 , n72239 , n72371 );
and ( n72373 , n72236 , n72372 );
or ( n72374 , n72235 , n72373 );
and ( n72375 , n72232 , n72374 );
or ( n72376 , n72231 , n72375 );
and ( n72377 , n72228 , n72376 );
or ( n72378 , n72227 , n72377 );
and ( n72379 , n72224 , n72378 );
or ( n72380 , n72223 , n72379 );
and ( n72381 , n72220 , n72380 );
or ( n72382 , n72219 , n72381 );
and ( n72383 , n72216 , n72382 );
or ( n72384 , n72215 , n72383 );
and ( n72385 , n72212 , n72384 );
or ( n72386 , n72211 , n72385 );
and ( n72387 , n72208 , n72386 );
or ( n72388 , n72207 , n72387 );
and ( n72389 , n72204 , n72388 );
or ( n72390 , n72203 , n72389 );
and ( n72391 , n72200 , n72390 );
or ( n72392 , n72199 , n72391 );
and ( n72393 , n72196 , n72392 );
or ( n72394 , n72195 , n72393 );
and ( n72395 , n72192 , n72394 );
or ( n72396 , n72191 , n72395 );
and ( n72397 , n72188 , n72396 );
or ( n72398 , n72187 , n72397 );
and ( n72399 , n72184 , n72398 );
or ( n72400 , n72183 , n72399 );
and ( n72401 , n72180 , n72400 );
or ( n72402 , n72179 , n72401 );
and ( n72403 , n72176 , n72402 );
or ( n72404 , n72175 , n72403 );
and ( n72405 , n72172 , n72404 );
or ( n72406 , n72171 , n72405 );
and ( n72407 , n72168 , n72406 );
or ( n72408 , n72167 , n72407 );
xor ( n72409 , n72164 , n72408 );
buf ( n72410 , n17934 );
and ( n72411 , n30209 , n72410 );
xor ( n72412 , n72409 , n72411 );
xor ( n72413 , n72168 , n72406 );
and ( n72414 , n30214 , n72410 );
and ( n72415 , n72413 , n72414 );
xor ( n72416 , n72413 , n72414 );
xor ( n72417 , n72172 , n72404 );
and ( n72418 , n30219 , n72410 );
and ( n72419 , n72417 , n72418 );
xor ( n72420 , n72417 , n72418 );
xor ( n72421 , n72176 , n72402 );
and ( n72422 , n30224 , n72410 );
and ( n72423 , n72421 , n72422 );
xor ( n72424 , n72421 , n72422 );
xor ( n72425 , n72180 , n72400 );
and ( n72426 , n30229 , n72410 );
and ( n72427 , n72425 , n72426 );
xor ( n72428 , n72425 , n72426 );
xor ( n72429 , n72184 , n72398 );
and ( n72430 , n30234 , n72410 );
and ( n72431 , n72429 , n72430 );
xor ( n72432 , n72429 , n72430 );
xor ( n72433 , n72188 , n72396 );
and ( n72434 , n30239 , n72410 );
and ( n72435 , n72433 , n72434 );
xor ( n72436 , n72433 , n72434 );
xor ( n72437 , n72192 , n72394 );
and ( n72438 , n30244 , n72410 );
and ( n72439 , n72437 , n72438 );
xor ( n72440 , n72437 , n72438 );
xor ( n72441 , n72196 , n72392 );
and ( n72442 , n30249 , n72410 );
and ( n72443 , n72441 , n72442 );
xor ( n72444 , n72441 , n72442 );
xor ( n72445 , n72200 , n72390 );
and ( n72446 , n30254 , n72410 );
and ( n72447 , n72445 , n72446 );
xor ( n72448 , n72445 , n72446 );
xor ( n72449 , n72204 , n72388 );
and ( n72450 , n30259 , n72410 );
and ( n72451 , n72449 , n72450 );
xor ( n72452 , n72449 , n72450 );
xor ( n72453 , n72208 , n72386 );
and ( n72454 , n30264 , n72410 );
and ( n72455 , n72453 , n72454 );
xor ( n72456 , n72453 , n72454 );
xor ( n72457 , n72212 , n72384 );
and ( n72458 , n30269 , n72410 );
and ( n72459 , n72457 , n72458 );
xor ( n72460 , n72457 , n72458 );
xor ( n72461 , n72216 , n72382 );
and ( n72462 , n30274 , n72410 );
and ( n72463 , n72461 , n72462 );
xor ( n72464 , n72461 , n72462 );
xor ( n72465 , n72220 , n72380 );
and ( n72466 , n30279 , n72410 );
and ( n72467 , n72465 , n72466 );
xor ( n72468 , n72465 , n72466 );
xor ( n72469 , n72224 , n72378 );
and ( n72470 , n30284 , n72410 );
and ( n72471 , n72469 , n72470 );
xor ( n72472 , n72469 , n72470 );
xor ( n72473 , n72228 , n72376 );
and ( n72474 , n30289 , n72410 );
and ( n72475 , n72473 , n72474 );
xor ( n72476 , n72473 , n72474 );
xor ( n72477 , n72232 , n72374 );
and ( n72478 , n30294 , n72410 );
and ( n72479 , n72477 , n72478 );
xor ( n72480 , n72477 , n72478 );
xor ( n72481 , n72236 , n72372 );
and ( n72482 , n30299 , n72410 );
and ( n72483 , n72481 , n72482 );
xor ( n72484 , n72481 , n72482 );
xor ( n72485 , n72240 , n72370 );
and ( n72486 , n30304 , n72410 );
and ( n72487 , n72485 , n72486 );
xor ( n72488 , n72485 , n72486 );
xor ( n72489 , n72244 , n72368 );
and ( n72490 , n30309 , n72410 );
and ( n72491 , n72489 , n72490 );
xor ( n72492 , n72489 , n72490 );
xor ( n72493 , n72248 , n72366 );
and ( n72494 , n30314 , n72410 );
and ( n72495 , n72493 , n72494 );
xor ( n72496 , n72493 , n72494 );
xor ( n72497 , n72252 , n72364 );
and ( n72498 , n30319 , n72410 );
and ( n72499 , n72497 , n72498 );
xor ( n72500 , n72497 , n72498 );
xor ( n72501 , n72256 , n72362 );
and ( n72502 , n30324 , n72410 );
and ( n72503 , n72501 , n72502 );
xor ( n72504 , n72501 , n72502 );
xor ( n72505 , n72260 , n72360 );
and ( n72506 , n30329 , n72410 );
and ( n72507 , n72505 , n72506 );
xor ( n72508 , n72505 , n72506 );
xor ( n72509 , n72264 , n72358 );
and ( n72510 , n30334 , n72410 );
and ( n72511 , n72509 , n72510 );
xor ( n72512 , n72509 , n72510 );
xor ( n72513 , n72268 , n72356 );
and ( n72514 , n30339 , n72410 );
and ( n72515 , n72513 , n72514 );
xor ( n72516 , n72513 , n72514 );
xor ( n72517 , n72272 , n72354 );
and ( n72518 , n30344 , n72410 );
and ( n72519 , n72517 , n72518 );
xor ( n72520 , n72517 , n72518 );
xor ( n72521 , n72276 , n72352 );
and ( n72522 , n30349 , n72410 );
and ( n72523 , n72521 , n72522 );
xor ( n72524 , n72521 , n72522 );
xor ( n72525 , n72280 , n72350 );
and ( n72526 , n30354 , n72410 );
and ( n72527 , n72525 , n72526 );
xor ( n72528 , n72525 , n72526 );
xor ( n72529 , n72284 , n72348 );
and ( n72530 , n30359 , n72410 );
and ( n72531 , n72529 , n72530 );
xor ( n72532 , n72529 , n72530 );
xor ( n72533 , n72288 , n72346 );
and ( n72534 , n30364 , n72410 );
and ( n72535 , n72533 , n72534 );
xor ( n72536 , n72533 , n72534 );
xor ( n72537 , n72292 , n72344 );
and ( n72538 , n30369 , n72410 );
and ( n72539 , n72537 , n72538 );
xor ( n72540 , n72537 , n72538 );
xor ( n72541 , n72296 , n72342 );
and ( n72542 , n30374 , n72410 );
and ( n72543 , n72541 , n72542 );
xor ( n72544 , n72541 , n72542 );
xor ( n72545 , n72300 , n72340 );
and ( n72546 , n30379 , n72410 );
and ( n72547 , n72545 , n72546 );
xor ( n72548 , n72545 , n72546 );
xor ( n72549 , n72304 , n72338 );
and ( n72550 , n30384 , n72410 );
and ( n72551 , n72549 , n72550 );
xor ( n72552 , n72549 , n72550 );
xor ( n72553 , n72308 , n72336 );
and ( n72554 , n30389 , n72410 );
and ( n72555 , n72553 , n72554 );
xor ( n72556 , n72553 , n72554 );
xor ( n72557 , n72312 , n72334 );
and ( n72558 , n30394 , n72410 );
and ( n72559 , n72557 , n72558 );
xor ( n72560 , n72557 , n72558 );
xor ( n72561 , n72316 , n72332 );
and ( n72562 , n30399 , n72410 );
and ( n72563 , n72561 , n72562 );
xor ( n72564 , n72561 , n72562 );
xor ( n72565 , n72320 , n72330 );
and ( n72566 , n30404 , n72410 );
and ( n72567 , n72565 , n72566 );
xor ( n72568 , n72565 , n72566 );
xor ( n72569 , n72324 , n72328 );
and ( n72570 , n30409 , n72410 );
and ( n72571 , n72569 , n72570 );
buf ( n72572 , n72571 );
and ( n72573 , n72568 , n72572 );
or ( n72574 , n72567 , n72573 );
and ( n72575 , n72564 , n72574 );
or ( n72576 , n72563 , n72575 );
and ( n72577 , n72560 , n72576 );
or ( n72578 , n72559 , n72577 );
and ( n72579 , n72556 , n72578 );
or ( n72580 , n72555 , n72579 );
and ( n72581 , n72552 , n72580 );
or ( n72582 , n72551 , n72581 );
and ( n72583 , n72548 , n72582 );
or ( n72584 , n72547 , n72583 );
and ( n72585 , n72544 , n72584 );
or ( n72586 , n72543 , n72585 );
and ( n72587 , n72540 , n72586 );
or ( n72588 , n72539 , n72587 );
and ( n72589 , n72536 , n72588 );
or ( n72590 , n72535 , n72589 );
and ( n72591 , n72532 , n72590 );
or ( n72592 , n72531 , n72591 );
and ( n72593 , n72528 , n72592 );
or ( n72594 , n72527 , n72593 );
and ( n72595 , n72524 , n72594 );
or ( n72596 , n72523 , n72595 );
and ( n72597 , n72520 , n72596 );
or ( n72598 , n72519 , n72597 );
and ( n72599 , n72516 , n72598 );
or ( n72600 , n72515 , n72599 );
and ( n72601 , n72512 , n72600 );
or ( n72602 , n72511 , n72601 );
and ( n72603 , n72508 , n72602 );
or ( n72604 , n72507 , n72603 );
and ( n72605 , n72504 , n72604 );
or ( n72606 , n72503 , n72605 );
and ( n72607 , n72500 , n72606 );
or ( n72608 , n72499 , n72607 );
and ( n72609 , n72496 , n72608 );
or ( n72610 , n72495 , n72609 );
and ( n72611 , n72492 , n72610 );
or ( n72612 , n72491 , n72611 );
and ( n72613 , n72488 , n72612 );
or ( n72614 , n72487 , n72613 );
and ( n72615 , n72484 , n72614 );
or ( n72616 , n72483 , n72615 );
and ( n72617 , n72480 , n72616 );
or ( n72618 , n72479 , n72617 );
and ( n72619 , n72476 , n72618 );
or ( n72620 , n72475 , n72619 );
and ( n72621 , n72472 , n72620 );
or ( n72622 , n72471 , n72621 );
and ( n72623 , n72468 , n72622 );
or ( n72624 , n72467 , n72623 );
and ( n72625 , n72464 , n72624 );
or ( n72626 , n72463 , n72625 );
and ( n72627 , n72460 , n72626 );
or ( n72628 , n72459 , n72627 );
and ( n72629 , n72456 , n72628 );
or ( n72630 , n72455 , n72629 );
and ( n72631 , n72452 , n72630 );
or ( n72632 , n72451 , n72631 );
and ( n72633 , n72448 , n72632 );
or ( n72634 , n72447 , n72633 );
and ( n72635 , n72444 , n72634 );
or ( n72636 , n72443 , n72635 );
and ( n72637 , n72440 , n72636 );
or ( n72638 , n72439 , n72637 );
and ( n72639 , n72436 , n72638 );
or ( n72640 , n72435 , n72639 );
and ( n72641 , n72432 , n72640 );
or ( n72642 , n72431 , n72641 );
and ( n72643 , n72428 , n72642 );
or ( n72644 , n72427 , n72643 );
and ( n72645 , n72424 , n72644 );
or ( n72646 , n72423 , n72645 );
and ( n72647 , n72420 , n72646 );
or ( n72648 , n72419 , n72647 );
and ( n72649 , n72416 , n72648 );
or ( n72650 , n72415 , n72649 );
xor ( n72651 , n72412 , n72650 );
buf ( n72652 , n17932 );
and ( n72653 , n30214 , n72652 );
xor ( n72654 , n72651 , n72653 );
xor ( n72655 , n72416 , n72648 );
and ( n72656 , n30219 , n72652 );
and ( n72657 , n72655 , n72656 );
xor ( n72658 , n72655 , n72656 );
xor ( n72659 , n72420 , n72646 );
and ( n72660 , n30224 , n72652 );
and ( n72661 , n72659 , n72660 );
xor ( n72662 , n72659 , n72660 );
xor ( n72663 , n72424 , n72644 );
and ( n72664 , n30229 , n72652 );
and ( n72665 , n72663 , n72664 );
xor ( n72666 , n72663 , n72664 );
xor ( n72667 , n72428 , n72642 );
and ( n72668 , n30234 , n72652 );
and ( n72669 , n72667 , n72668 );
xor ( n72670 , n72667 , n72668 );
xor ( n72671 , n72432 , n72640 );
and ( n72672 , n30239 , n72652 );
and ( n72673 , n72671 , n72672 );
xor ( n72674 , n72671 , n72672 );
xor ( n72675 , n72436 , n72638 );
and ( n72676 , n30244 , n72652 );
and ( n72677 , n72675 , n72676 );
xor ( n72678 , n72675 , n72676 );
xor ( n72679 , n72440 , n72636 );
and ( n72680 , n30249 , n72652 );
and ( n72681 , n72679 , n72680 );
xor ( n72682 , n72679 , n72680 );
xor ( n72683 , n72444 , n72634 );
and ( n72684 , n30254 , n72652 );
and ( n72685 , n72683 , n72684 );
xor ( n72686 , n72683 , n72684 );
xor ( n72687 , n72448 , n72632 );
and ( n72688 , n30259 , n72652 );
and ( n72689 , n72687 , n72688 );
xor ( n72690 , n72687 , n72688 );
xor ( n72691 , n72452 , n72630 );
and ( n72692 , n30264 , n72652 );
and ( n72693 , n72691 , n72692 );
xor ( n72694 , n72691 , n72692 );
xor ( n72695 , n72456 , n72628 );
and ( n72696 , n30269 , n72652 );
and ( n72697 , n72695 , n72696 );
xor ( n72698 , n72695 , n72696 );
xor ( n72699 , n72460 , n72626 );
and ( n72700 , n30274 , n72652 );
and ( n72701 , n72699 , n72700 );
xor ( n72702 , n72699 , n72700 );
xor ( n72703 , n72464 , n72624 );
and ( n72704 , n30279 , n72652 );
and ( n72705 , n72703 , n72704 );
xor ( n72706 , n72703 , n72704 );
xor ( n72707 , n72468 , n72622 );
and ( n72708 , n30284 , n72652 );
and ( n72709 , n72707 , n72708 );
xor ( n72710 , n72707 , n72708 );
xor ( n72711 , n72472 , n72620 );
and ( n72712 , n30289 , n72652 );
and ( n72713 , n72711 , n72712 );
xor ( n72714 , n72711 , n72712 );
xor ( n72715 , n72476 , n72618 );
and ( n72716 , n30294 , n72652 );
and ( n72717 , n72715 , n72716 );
xor ( n72718 , n72715 , n72716 );
xor ( n72719 , n72480 , n72616 );
and ( n72720 , n30299 , n72652 );
and ( n72721 , n72719 , n72720 );
xor ( n72722 , n72719 , n72720 );
xor ( n72723 , n72484 , n72614 );
and ( n72724 , n30304 , n72652 );
and ( n72725 , n72723 , n72724 );
xor ( n72726 , n72723 , n72724 );
xor ( n72727 , n72488 , n72612 );
and ( n72728 , n30309 , n72652 );
and ( n72729 , n72727 , n72728 );
xor ( n72730 , n72727 , n72728 );
xor ( n72731 , n72492 , n72610 );
and ( n72732 , n30314 , n72652 );
and ( n72733 , n72731 , n72732 );
xor ( n72734 , n72731 , n72732 );
xor ( n72735 , n72496 , n72608 );
and ( n72736 , n30319 , n72652 );
and ( n72737 , n72735 , n72736 );
xor ( n72738 , n72735 , n72736 );
xor ( n72739 , n72500 , n72606 );
and ( n72740 , n30324 , n72652 );
and ( n72741 , n72739 , n72740 );
xor ( n72742 , n72739 , n72740 );
xor ( n72743 , n72504 , n72604 );
and ( n72744 , n30329 , n72652 );
and ( n72745 , n72743 , n72744 );
xor ( n72746 , n72743 , n72744 );
xor ( n72747 , n72508 , n72602 );
and ( n72748 , n30334 , n72652 );
and ( n72749 , n72747 , n72748 );
xor ( n72750 , n72747 , n72748 );
xor ( n72751 , n72512 , n72600 );
and ( n72752 , n30339 , n72652 );
and ( n72753 , n72751 , n72752 );
xor ( n72754 , n72751 , n72752 );
xor ( n72755 , n72516 , n72598 );
and ( n72756 , n30344 , n72652 );
and ( n72757 , n72755 , n72756 );
xor ( n72758 , n72755 , n72756 );
xor ( n72759 , n72520 , n72596 );
and ( n72760 , n30349 , n72652 );
and ( n72761 , n72759 , n72760 );
xor ( n72762 , n72759 , n72760 );
xor ( n72763 , n72524 , n72594 );
and ( n72764 , n30354 , n72652 );
and ( n72765 , n72763 , n72764 );
xor ( n72766 , n72763 , n72764 );
xor ( n72767 , n72528 , n72592 );
and ( n72768 , n30359 , n72652 );
and ( n72769 , n72767 , n72768 );
xor ( n72770 , n72767 , n72768 );
xor ( n72771 , n72532 , n72590 );
and ( n72772 , n30364 , n72652 );
and ( n72773 , n72771 , n72772 );
xor ( n72774 , n72771 , n72772 );
xor ( n72775 , n72536 , n72588 );
and ( n72776 , n30369 , n72652 );
and ( n72777 , n72775 , n72776 );
xor ( n72778 , n72775 , n72776 );
xor ( n72779 , n72540 , n72586 );
and ( n72780 , n30374 , n72652 );
and ( n72781 , n72779 , n72780 );
xor ( n72782 , n72779 , n72780 );
xor ( n72783 , n72544 , n72584 );
and ( n72784 , n30379 , n72652 );
and ( n72785 , n72783 , n72784 );
xor ( n72786 , n72783 , n72784 );
xor ( n72787 , n72548 , n72582 );
and ( n72788 , n30384 , n72652 );
and ( n72789 , n72787 , n72788 );
xor ( n72790 , n72787 , n72788 );
xor ( n72791 , n72552 , n72580 );
and ( n72792 , n30389 , n72652 );
and ( n72793 , n72791 , n72792 );
xor ( n72794 , n72791 , n72792 );
xor ( n72795 , n72556 , n72578 );
and ( n72796 , n30394 , n72652 );
and ( n72797 , n72795 , n72796 );
xor ( n72798 , n72795 , n72796 );
xor ( n72799 , n72560 , n72576 );
and ( n72800 , n30399 , n72652 );
and ( n72801 , n72799 , n72800 );
xor ( n72802 , n72799 , n72800 );
xor ( n72803 , n72564 , n72574 );
and ( n72804 , n30404 , n72652 );
and ( n72805 , n72803 , n72804 );
xor ( n72806 , n72803 , n72804 );
xor ( n72807 , n72568 , n72572 );
and ( n72808 , n30409 , n72652 );
and ( n72809 , n72807 , n72808 );
buf ( n72810 , n72809 );
and ( n72811 , n72806 , n72810 );
or ( n72812 , n72805 , n72811 );
and ( n72813 , n72802 , n72812 );
or ( n72814 , n72801 , n72813 );
and ( n72815 , n72798 , n72814 );
or ( n72816 , n72797 , n72815 );
and ( n72817 , n72794 , n72816 );
or ( n72818 , n72793 , n72817 );
and ( n72819 , n72790 , n72818 );
or ( n72820 , n72789 , n72819 );
and ( n72821 , n72786 , n72820 );
or ( n72822 , n72785 , n72821 );
and ( n72823 , n72782 , n72822 );
or ( n72824 , n72781 , n72823 );
and ( n72825 , n72778 , n72824 );
or ( n72826 , n72777 , n72825 );
and ( n72827 , n72774 , n72826 );
or ( n72828 , n72773 , n72827 );
and ( n72829 , n72770 , n72828 );
or ( n72830 , n72769 , n72829 );
and ( n72831 , n72766 , n72830 );
or ( n72832 , n72765 , n72831 );
and ( n72833 , n72762 , n72832 );
or ( n72834 , n72761 , n72833 );
and ( n72835 , n72758 , n72834 );
or ( n72836 , n72757 , n72835 );
and ( n72837 , n72754 , n72836 );
or ( n72838 , n72753 , n72837 );
and ( n72839 , n72750 , n72838 );
or ( n72840 , n72749 , n72839 );
and ( n72841 , n72746 , n72840 );
or ( n72842 , n72745 , n72841 );
and ( n72843 , n72742 , n72842 );
or ( n72844 , n72741 , n72843 );
and ( n72845 , n72738 , n72844 );
or ( n72846 , n72737 , n72845 );
and ( n72847 , n72734 , n72846 );
or ( n72848 , n72733 , n72847 );
and ( n72849 , n72730 , n72848 );
or ( n72850 , n72729 , n72849 );
and ( n72851 , n72726 , n72850 );
or ( n72852 , n72725 , n72851 );
and ( n72853 , n72722 , n72852 );
or ( n72854 , n72721 , n72853 );
and ( n72855 , n72718 , n72854 );
or ( n72856 , n72717 , n72855 );
and ( n72857 , n72714 , n72856 );
or ( n72858 , n72713 , n72857 );
and ( n72859 , n72710 , n72858 );
or ( n72860 , n72709 , n72859 );
and ( n72861 , n72706 , n72860 );
or ( n72862 , n72705 , n72861 );
and ( n72863 , n72702 , n72862 );
or ( n72864 , n72701 , n72863 );
and ( n72865 , n72698 , n72864 );
or ( n72866 , n72697 , n72865 );
and ( n72867 , n72694 , n72866 );
or ( n72868 , n72693 , n72867 );
and ( n72869 , n72690 , n72868 );
or ( n72870 , n72689 , n72869 );
and ( n72871 , n72686 , n72870 );
or ( n72872 , n72685 , n72871 );
and ( n72873 , n72682 , n72872 );
or ( n72874 , n72681 , n72873 );
and ( n72875 , n72678 , n72874 );
or ( n72876 , n72677 , n72875 );
and ( n72877 , n72674 , n72876 );
or ( n72878 , n72673 , n72877 );
and ( n72879 , n72670 , n72878 );
or ( n72880 , n72669 , n72879 );
and ( n72881 , n72666 , n72880 );
or ( n72882 , n72665 , n72881 );
and ( n72883 , n72662 , n72882 );
or ( n72884 , n72661 , n72883 );
and ( n72885 , n72658 , n72884 );
or ( n72886 , n72657 , n72885 );
xor ( n72887 , n72654 , n72886 );
buf ( n72888 , n17930 );
and ( n72889 , n30219 , n72888 );
xor ( n72890 , n72887 , n72889 );
xor ( n72891 , n72658 , n72884 );
and ( n72892 , n30224 , n72888 );
and ( n72893 , n72891 , n72892 );
xor ( n72894 , n72891 , n72892 );
xor ( n72895 , n72662 , n72882 );
and ( n72896 , n30229 , n72888 );
and ( n72897 , n72895 , n72896 );
xor ( n72898 , n72895 , n72896 );
xor ( n72899 , n72666 , n72880 );
and ( n72900 , n30234 , n72888 );
and ( n72901 , n72899 , n72900 );
xor ( n72902 , n72899 , n72900 );
xor ( n72903 , n72670 , n72878 );
and ( n72904 , n30239 , n72888 );
and ( n72905 , n72903 , n72904 );
xor ( n72906 , n72903 , n72904 );
xor ( n72907 , n72674 , n72876 );
and ( n72908 , n30244 , n72888 );
and ( n72909 , n72907 , n72908 );
xor ( n72910 , n72907 , n72908 );
xor ( n72911 , n72678 , n72874 );
and ( n72912 , n30249 , n72888 );
and ( n72913 , n72911 , n72912 );
xor ( n72914 , n72911 , n72912 );
xor ( n72915 , n72682 , n72872 );
and ( n72916 , n30254 , n72888 );
and ( n72917 , n72915 , n72916 );
xor ( n72918 , n72915 , n72916 );
xor ( n72919 , n72686 , n72870 );
and ( n72920 , n30259 , n72888 );
and ( n72921 , n72919 , n72920 );
xor ( n72922 , n72919 , n72920 );
xor ( n72923 , n72690 , n72868 );
and ( n72924 , n30264 , n72888 );
and ( n72925 , n72923 , n72924 );
xor ( n72926 , n72923 , n72924 );
xor ( n72927 , n72694 , n72866 );
and ( n72928 , n30269 , n72888 );
and ( n72929 , n72927 , n72928 );
xor ( n72930 , n72927 , n72928 );
xor ( n72931 , n72698 , n72864 );
and ( n72932 , n30274 , n72888 );
and ( n72933 , n72931 , n72932 );
xor ( n72934 , n72931 , n72932 );
xor ( n72935 , n72702 , n72862 );
and ( n72936 , n30279 , n72888 );
and ( n72937 , n72935 , n72936 );
xor ( n72938 , n72935 , n72936 );
xor ( n72939 , n72706 , n72860 );
and ( n72940 , n30284 , n72888 );
and ( n72941 , n72939 , n72940 );
xor ( n72942 , n72939 , n72940 );
xor ( n72943 , n72710 , n72858 );
and ( n72944 , n30289 , n72888 );
and ( n72945 , n72943 , n72944 );
xor ( n72946 , n72943 , n72944 );
xor ( n72947 , n72714 , n72856 );
and ( n72948 , n30294 , n72888 );
and ( n72949 , n72947 , n72948 );
xor ( n72950 , n72947 , n72948 );
xor ( n72951 , n72718 , n72854 );
and ( n72952 , n30299 , n72888 );
and ( n72953 , n72951 , n72952 );
xor ( n72954 , n72951 , n72952 );
xor ( n72955 , n72722 , n72852 );
and ( n72956 , n30304 , n72888 );
and ( n72957 , n72955 , n72956 );
xor ( n72958 , n72955 , n72956 );
xor ( n72959 , n72726 , n72850 );
and ( n72960 , n30309 , n72888 );
and ( n72961 , n72959 , n72960 );
xor ( n72962 , n72959 , n72960 );
xor ( n72963 , n72730 , n72848 );
and ( n72964 , n30314 , n72888 );
and ( n72965 , n72963 , n72964 );
xor ( n72966 , n72963 , n72964 );
xor ( n72967 , n72734 , n72846 );
and ( n72968 , n30319 , n72888 );
and ( n72969 , n72967 , n72968 );
xor ( n72970 , n72967 , n72968 );
xor ( n72971 , n72738 , n72844 );
and ( n72972 , n30324 , n72888 );
and ( n72973 , n72971 , n72972 );
xor ( n72974 , n72971 , n72972 );
xor ( n72975 , n72742 , n72842 );
and ( n72976 , n30329 , n72888 );
and ( n72977 , n72975 , n72976 );
xor ( n72978 , n72975 , n72976 );
xor ( n72979 , n72746 , n72840 );
and ( n72980 , n30334 , n72888 );
and ( n72981 , n72979 , n72980 );
xor ( n72982 , n72979 , n72980 );
xor ( n72983 , n72750 , n72838 );
and ( n72984 , n30339 , n72888 );
and ( n72985 , n72983 , n72984 );
xor ( n72986 , n72983 , n72984 );
xor ( n72987 , n72754 , n72836 );
and ( n72988 , n30344 , n72888 );
and ( n72989 , n72987 , n72988 );
xor ( n72990 , n72987 , n72988 );
xor ( n72991 , n72758 , n72834 );
and ( n72992 , n30349 , n72888 );
and ( n72993 , n72991 , n72992 );
xor ( n72994 , n72991 , n72992 );
xor ( n72995 , n72762 , n72832 );
and ( n72996 , n30354 , n72888 );
and ( n72997 , n72995 , n72996 );
xor ( n72998 , n72995 , n72996 );
xor ( n72999 , n72766 , n72830 );
and ( n73000 , n30359 , n72888 );
and ( n73001 , n72999 , n73000 );
xor ( n73002 , n72999 , n73000 );
xor ( n73003 , n72770 , n72828 );
and ( n73004 , n30364 , n72888 );
and ( n73005 , n73003 , n73004 );
xor ( n73006 , n73003 , n73004 );
xor ( n73007 , n72774 , n72826 );
and ( n73008 , n30369 , n72888 );
and ( n73009 , n73007 , n73008 );
xor ( n73010 , n73007 , n73008 );
xor ( n73011 , n72778 , n72824 );
and ( n73012 , n30374 , n72888 );
and ( n73013 , n73011 , n73012 );
xor ( n73014 , n73011 , n73012 );
xor ( n73015 , n72782 , n72822 );
and ( n73016 , n30379 , n72888 );
and ( n73017 , n73015 , n73016 );
xor ( n73018 , n73015 , n73016 );
xor ( n73019 , n72786 , n72820 );
and ( n73020 , n30384 , n72888 );
and ( n73021 , n73019 , n73020 );
xor ( n73022 , n73019 , n73020 );
xor ( n73023 , n72790 , n72818 );
and ( n73024 , n30389 , n72888 );
and ( n73025 , n73023 , n73024 );
xor ( n73026 , n73023 , n73024 );
xor ( n73027 , n72794 , n72816 );
and ( n73028 , n30394 , n72888 );
and ( n73029 , n73027 , n73028 );
xor ( n73030 , n73027 , n73028 );
xor ( n73031 , n72798 , n72814 );
and ( n73032 , n30399 , n72888 );
and ( n73033 , n73031 , n73032 );
xor ( n73034 , n73031 , n73032 );
xor ( n73035 , n72802 , n72812 );
and ( n73036 , n30404 , n72888 );
and ( n73037 , n73035 , n73036 );
xor ( n73038 , n73035 , n73036 );
xor ( n73039 , n72806 , n72810 );
and ( n73040 , n30409 , n72888 );
and ( n73041 , n73039 , n73040 );
buf ( n73042 , n73041 );
and ( n73043 , n73038 , n73042 );
or ( n73044 , n73037 , n73043 );
and ( n73045 , n73034 , n73044 );
or ( n73046 , n73033 , n73045 );
and ( n73047 , n73030 , n73046 );
or ( n73048 , n73029 , n73047 );
and ( n73049 , n73026 , n73048 );
or ( n73050 , n73025 , n73049 );
and ( n73051 , n73022 , n73050 );
or ( n73052 , n73021 , n73051 );
and ( n73053 , n73018 , n73052 );
or ( n73054 , n73017 , n73053 );
and ( n73055 , n73014 , n73054 );
or ( n73056 , n73013 , n73055 );
and ( n73057 , n73010 , n73056 );
or ( n73058 , n73009 , n73057 );
and ( n73059 , n73006 , n73058 );
or ( n73060 , n73005 , n73059 );
and ( n73061 , n73002 , n73060 );
or ( n73062 , n73001 , n73061 );
and ( n73063 , n72998 , n73062 );
or ( n73064 , n72997 , n73063 );
and ( n73065 , n72994 , n73064 );
or ( n73066 , n72993 , n73065 );
and ( n73067 , n72990 , n73066 );
or ( n73068 , n72989 , n73067 );
and ( n73069 , n72986 , n73068 );
or ( n73070 , n72985 , n73069 );
and ( n73071 , n72982 , n73070 );
or ( n73072 , n72981 , n73071 );
and ( n73073 , n72978 , n73072 );
or ( n73074 , n72977 , n73073 );
and ( n73075 , n72974 , n73074 );
or ( n73076 , n72973 , n73075 );
and ( n73077 , n72970 , n73076 );
or ( n73078 , n72969 , n73077 );
and ( n73079 , n72966 , n73078 );
or ( n73080 , n72965 , n73079 );
and ( n73081 , n72962 , n73080 );
or ( n73082 , n72961 , n73081 );
and ( n73083 , n72958 , n73082 );
or ( n73084 , n72957 , n73083 );
and ( n73085 , n72954 , n73084 );
or ( n73086 , n72953 , n73085 );
and ( n73087 , n72950 , n73086 );
or ( n73088 , n72949 , n73087 );
and ( n73089 , n72946 , n73088 );
or ( n73090 , n72945 , n73089 );
and ( n73091 , n72942 , n73090 );
or ( n73092 , n72941 , n73091 );
and ( n73093 , n72938 , n73092 );
or ( n73094 , n72937 , n73093 );
and ( n73095 , n72934 , n73094 );
or ( n73096 , n72933 , n73095 );
and ( n73097 , n72930 , n73096 );
or ( n73098 , n72929 , n73097 );
and ( n73099 , n72926 , n73098 );
or ( n73100 , n72925 , n73099 );
and ( n73101 , n72922 , n73100 );
or ( n73102 , n72921 , n73101 );
and ( n73103 , n72918 , n73102 );
or ( n73104 , n72917 , n73103 );
and ( n73105 , n72914 , n73104 );
or ( n73106 , n72913 , n73105 );
and ( n73107 , n72910 , n73106 );
or ( n73108 , n72909 , n73107 );
and ( n73109 , n72906 , n73108 );
or ( n73110 , n72905 , n73109 );
and ( n73111 , n72902 , n73110 );
or ( n73112 , n72901 , n73111 );
and ( n73113 , n72898 , n73112 );
or ( n73114 , n72897 , n73113 );
and ( n73115 , n72894 , n73114 );
or ( n73116 , n72893 , n73115 );
xor ( n73117 , n72890 , n73116 );
buf ( n73118 , n17928 );
and ( n73119 , n30224 , n73118 );
xor ( n73120 , n73117 , n73119 );
xor ( n73121 , n72894 , n73114 );
and ( n73122 , n30229 , n73118 );
and ( n73123 , n73121 , n73122 );
xor ( n73124 , n73121 , n73122 );
xor ( n73125 , n72898 , n73112 );
and ( n73126 , n30234 , n73118 );
and ( n73127 , n73125 , n73126 );
xor ( n73128 , n73125 , n73126 );
xor ( n73129 , n72902 , n73110 );
and ( n73130 , n30239 , n73118 );
and ( n73131 , n73129 , n73130 );
xor ( n73132 , n73129 , n73130 );
xor ( n73133 , n72906 , n73108 );
and ( n73134 , n30244 , n73118 );
and ( n73135 , n73133 , n73134 );
xor ( n73136 , n73133 , n73134 );
xor ( n73137 , n72910 , n73106 );
and ( n73138 , n30249 , n73118 );
and ( n73139 , n73137 , n73138 );
xor ( n73140 , n73137 , n73138 );
xor ( n73141 , n72914 , n73104 );
and ( n73142 , n30254 , n73118 );
and ( n73143 , n73141 , n73142 );
xor ( n73144 , n73141 , n73142 );
xor ( n73145 , n72918 , n73102 );
and ( n73146 , n30259 , n73118 );
and ( n73147 , n73145 , n73146 );
xor ( n73148 , n73145 , n73146 );
xor ( n73149 , n72922 , n73100 );
and ( n73150 , n30264 , n73118 );
and ( n73151 , n73149 , n73150 );
xor ( n73152 , n73149 , n73150 );
xor ( n73153 , n72926 , n73098 );
and ( n73154 , n30269 , n73118 );
and ( n73155 , n73153 , n73154 );
xor ( n73156 , n73153 , n73154 );
xor ( n73157 , n72930 , n73096 );
and ( n73158 , n30274 , n73118 );
and ( n73159 , n73157 , n73158 );
xor ( n73160 , n73157 , n73158 );
xor ( n73161 , n72934 , n73094 );
and ( n73162 , n30279 , n73118 );
and ( n73163 , n73161 , n73162 );
xor ( n73164 , n73161 , n73162 );
xor ( n73165 , n72938 , n73092 );
and ( n73166 , n30284 , n73118 );
and ( n73167 , n73165 , n73166 );
xor ( n73168 , n73165 , n73166 );
xor ( n73169 , n72942 , n73090 );
and ( n73170 , n30289 , n73118 );
and ( n73171 , n73169 , n73170 );
xor ( n73172 , n73169 , n73170 );
xor ( n73173 , n72946 , n73088 );
and ( n73174 , n30294 , n73118 );
and ( n73175 , n73173 , n73174 );
xor ( n73176 , n73173 , n73174 );
xor ( n73177 , n72950 , n73086 );
and ( n73178 , n30299 , n73118 );
and ( n73179 , n73177 , n73178 );
xor ( n73180 , n73177 , n73178 );
xor ( n73181 , n72954 , n73084 );
and ( n73182 , n30304 , n73118 );
and ( n73183 , n73181 , n73182 );
xor ( n73184 , n73181 , n73182 );
xor ( n73185 , n72958 , n73082 );
and ( n73186 , n30309 , n73118 );
and ( n73187 , n73185 , n73186 );
xor ( n73188 , n73185 , n73186 );
xor ( n73189 , n72962 , n73080 );
and ( n73190 , n30314 , n73118 );
and ( n73191 , n73189 , n73190 );
xor ( n73192 , n73189 , n73190 );
xor ( n73193 , n72966 , n73078 );
and ( n73194 , n30319 , n73118 );
and ( n73195 , n73193 , n73194 );
xor ( n73196 , n73193 , n73194 );
xor ( n73197 , n72970 , n73076 );
and ( n73198 , n30324 , n73118 );
and ( n73199 , n73197 , n73198 );
xor ( n73200 , n73197 , n73198 );
xor ( n73201 , n72974 , n73074 );
and ( n73202 , n30329 , n73118 );
and ( n73203 , n73201 , n73202 );
xor ( n73204 , n73201 , n73202 );
xor ( n73205 , n72978 , n73072 );
and ( n73206 , n30334 , n73118 );
and ( n73207 , n73205 , n73206 );
xor ( n73208 , n73205 , n73206 );
xor ( n73209 , n72982 , n73070 );
and ( n73210 , n30339 , n73118 );
and ( n73211 , n73209 , n73210 );
xor ( n73212 , n73209 , n73210 );
xor ( n73213 , n72986 , n73068 );
and ( n73214 , n30344 , n73118 );
and ( n73215 , n73213 , n73214 );
xor ( n73216 , n73213 , n73214 );
xor ( n73217 , n72990 , n73066 );
and ( n73218 , n30349 , n73118 );
and ( n73219 , n73217 , n73218 );
xor ( n73220 , n73217 , n73218 );
xor ( n73221 , n72994 , n73064 );
and ( n73222 , n30354 , n73118 );
and ( n73223 , n73221 , n73222 );
xor ( n73224 , n73221 , n73222 );
xor ( n73225 , n72998 , n73062 );
and ( n73226 , n30359 , n73118 );
and ( n73227 , n73225 , n73226 );
xor ( n73228 , n73225 , n73226 );
xor ( n73229 , n73002 , n73060 );
and ( n73230 , n30364 , n73118 );
and ( n73231 , n73229 , n73230 );
xor ( n73232 , n73229 , n73230 );
xor ( n73233 , n73006 , n73058 );
and ( n73234 , n30369 , n73118 );
and ( n73235 , n73233 , n73234 );
xor ( n73236 , n73233 , n73234 );
xor ( n73237 , n73010 , n73056 );
and ( n73238 , n30374 , n73118 );
and ( n73239 , n73237 , n73238 );
xor ( n73240 , n73237 , n73238 );
xor ( n73241 , n73014 , n73054 );
and ( n73242 , n30379 , n73118 );
and ( n73243 , n73241 , n73242 );
xor ( n73244 , n73241 , n73242 );
xor ( n73245 , n73018 , n73052 );
and ( n73246 , n30384 , n73118 );
and ( n73247 , n73245 , n73246 );
xor ( n73248 , n73245 , n73246 );
xor ( n73249 , n73022 , n73050 );
and ( n73250 , n30389 , n73118 );
and ( n73251 , n73249 , n73250 );
xor ( n73252 , n73249 , n73250 );
xor ( n73253 , n73026 , n73048 );
and ( n73254 , n30394 , n73118 );
and ( n73255 , n73253 , n73254 );
xor ( n73256 , n73253 , n73254 );
xor ( n73257 , n73030 , n73046 );
and ( n73258 , n30399 , n73118 );
and ( n73259 , n73257 , n73258 );
xor ( n73260 , n73257 , n73258 );
xor ( n73261 , n73034 , n73044 );
and ( n73262 , n30404 , n73118 );
and ( n73263 , n73261 , n73262 );
xor ( n73264 , n73261 , n73262 );
xor ( n73265 , n73038 , n73042 );
and ( n73266 , n30409 , n73118 );
and ( n73267 , n73265 , n73266 );
buf ( n73268 , n73267 );
and ( n73269 , n73264 , n73268 );
or ( n73270 , n73263 , n73269 );
and ( n73271 , n73260 , n73270 );
or ( n73272 , n73259 , n73271 );
and ( n73273 , n73256 , n73272 );
or ( n73274 , n73255 , n73273 );
and ( n73275 , n73252 , n73274 );
or ( n73276 , n73251 , n73275 );
and ( n73277 , n73248 , n73276 );
or ( n73278 , n73247 , n73277 );
and ( n73279 , n73244 , n73278 );
or ( n73280 , n73243 , n73279 );
and ( n73281 , n73240 , n73280 );
or ( n73282 , n73239 , n73281 );
and ( n73283 , n73236 , n73282 );
or ( n73284 , n73235 , n73283 );
and ( n73285 , n73232 , n73284 );
or ( n73286 , n73231 , n73285 );
and ( n73287 , n73228 , n73286 );
or ( n73288 , n73227 , n73287 );
and ( n73289 , n73224 , n73288 );
or ( n73290 , n73223 , n73289 );
and ( n73291 , n73220 , n73290 );
or ( n73292 , n73219 , n73291 );
and ( n73293 , n73216 , n73292 );
or ( n73294 , n73215 , n73293 );
and ( n73295 , n73212 , n73294 );
or ( n73296 , n73211 , n73295 );
and ( n73297 , n73208 , n73296 );
or ( n73298 , n73207 , n73297 );
and ( n73299 , n73204 , n73298 );
or ( n73300 , n73203 , n73299 );
and ( n73301 , n73200 , n73300 );
or ( n73302 , n73199 , n73301 );
and ( n73303 , n73196 , n73302 );
or ( n73304 , n73195 , n73303 );
and ( n73305 , n73192 , n73304 );
or ( n73306 , n73191 , n73305 );
and ( n73307 , n73188 , n73306 );
or ( n73308 , n73187 , n73307 );
and ( n73309 , n73184 , n73308 );
or ( n73310 , n73183 , n73309 );
and ( n73311 , n73180 , n73310 );
or ( n73312 , n73179 , n73311 );
and ( n73313 , n73176 , n73312 );
or ( n73314 , n73175 , n73313 );
and ( n73315 , n73172 , n73314 );
or ( n73316 , n73171 , n73315 );
and ( n73317 , n73168 , n73316 );
or ( n73318 , n73167 , n73317 );
and ( n73319 , n73164 , n73318 );
or ( n73320 , n73163 , n73319 );
and ( n73321 , n73160 , n73320 );
or ( n73322 , n73159 , n73321 );
and ( n73323 , n73156 , n73322 );
or ( n73324 , n73155 , n73323 );
and ( n73325 , n73152 , n73324 );
or ( n73326 , n73151 , n73325 );
and ( n73327 , n73148 , n73326 );
or ( n73328 , n73147 , n73327 );
and ( n73329 , n73144 , n73328 );
or ( n73330 , n73143 , n73329 );
and ( n73331 , n73140 , n73330 );
or ( n73332 , n73139 , n73331 );
and ( n73333 , n73136 , n73332 );
or ( n73334 , n73135 , n73333 );
and ( n73335 , n73132 , n73334 );
or ( n73336 , n73131 , n73335 );
and ( n73337 , n73128 , n73336 );
or ( n73338 , n73127 , n73337 );
and ( n73339 , n73124 , n73338 );
or ( n73340 , n73123 , n73339 );
xor ( n73341 , n73120 , n73340 );
buf ( n73342 , n17926 );
and ( n73343 , n30229 , n73342 );
xor ( n73344 , n73341 , n73343 );
xor ( n73345 , n73124 , n73338 );
and ( n73346 , n30234 , n73342 );
and ( n73347 , n73345 , n73346 );
xor ( n73348 , n73345 , n73346 );
xor ( n73349 , n73128 , n73336 );
and ( n73350 , n30239 , n73342 );
and ( n73351 , n73349 , n73350 );
xor ( n73352 , n73349 , n73350 );
xor ( n73353 , n73132 , n73334 );
and ( n73354 , n30244 , n73342 );
and ( n73355 , n73353 , n73354 );
xor ( n73356 , n73353 , n73354 );
xor ( n73357 , n73136 , n73332 );
and ( n73358 , n30249 , n73342 );
and ( n73359 , n73357 , n73358 );
xor ( n73360 , n73357 , n73358 );
xor ( n73361 , n73140 , n73330 );
and ( n73362 , n30254 , n73342 );
and ( n73363 , n73361 , n73362 );
xor ( n73364 , n73361 , n73362 );
xor ( n73365 , n73144 , n73328 );
and ( n73366 , n30259 , n73342 );
and ( n73367 , n73365 , n73366 );
xor ( n73368 , n73365 , n73366 );
xor ( n73369 , n73148 , n73326 );
and ( n73370 , n30264 , n73342 );
and ( n73371 , n73369 , n73370 );
xor ( n73372 , n73369 , n73370 );
xor ( n73373 , n73152 , n73324 );
and ( n73374 , n30269 , n73342 );
and ( n73375 , n73373 , n73374 );
xor ( n73376 , n73373 , n73374 );
xor ( n73377 , n73156 , n73322 );
and ( n73378 , n30274 , n73342 );
and ( n73379 , n73377 , n73378 );
xor ( n73380 , n73377 , n73378 );
xor ( n73381 , n73160 , n73320 );
and ( n73382 , n30279 , n73342 );
and ( n73383 , n73381 , n73382 );
xor ( n73384 , n73381 , n73382 );
xor ( n73385 , n73164 , n73318 );
and ( n73386 , n30284 , n73342 );
and ( n73387 , n73385 , n73386 );
xor ( n73388 , n73385 , n73386 );
xor ( n73389 , n73168 , n73316 );
and ( n73390 , n30289 , n73342 );
and ( n73391 , n73389 , n73390 );
xor ( n73392 , n73389 , n73390 );
xor ( n73393 , n73172 , n73314 );
and ( n73394 , n30294 , n73342 );
and ( n73395 , n73393 , n73394 );
xor ( n73396 , n73393 , n73394 );
xor ( n73397 , n73176 , n73312 );
and ( n73398 , n30299 , n73342 );
and ( n73399 , n73397 , n73398 );
xor ( n73400 , n73397 , n73398 );
xor ( n73401 , n73180 , n73310 );
and ( n73402 , n30304 , n73342 );
and ( n73403 , n73401 , n73402 );
xor ( n73404 , n73401 , n73402 );
xor ( n73405 , n73184 , n73308 );
and ( n73406 , n30309 , n73342 );
and ( n73407 , n73405 , n73406 );
xor ( n73408 , n73405 , n73406 );
xor ( n73409 , n73188 , n73306 );
and ( n73410 , n30314 , n73342 );
and ( n73411 , n73409 , n73410 );
xor ( n73412 , n73409 , n73410 );
xor ( n73413 , n73192 , n73304 );
and ( n73414 , n30319 , n73342 );
and ( n73415 , n73413 , n73414 );
xor ( n73416 , n73413 , n73414 );
xor ( n73417 , n73196 , n73302 );
and ( n73418 , n30324 , n73342 );
and ( n73419 , n73417 , n73418 );
xor ( n73420 , n73417 , n73418 );
xor ( n73421 , n73200 , n73300 );
and ( n73422 , n30329 , n73342 );
and ( n73423 , n73421 , n73422 );
xor ( n73424 , n73421 , n73422 );
xor ( n73425 , n73204 , n73298 );
and ( n73426 , n30334 , n73342 );
and ( n73427 , n73425 , n73426 );
xor ( n73428 , n73425 , n73426 );
xor ( n73429 , n73208 , n73296 );
and ( n73430 , n30339 , n73342 );
and ( n73431 , n73429 , n73430 );
xor ( n73432 , n73429 , n73430 );
xor ( n73433 , n73212 , n73294 );
and ( n73434 , n30344 , n73342 );
and ( n73435 , n73433 , n73434 );
xor ( n73436 , n73433 , n73434 );
xor ( n73437 , n73216 , n73292 );
and ( n73438 , n30349 , n73342 );
and ( n73439 , n73437 , n73438 );
xor ( n73440 , n73437 , n73438 );
xor ( n73441 , n73220 , n73290 );
and ( n73442 , n30354 , n73342 );
and ( n73443 , n73441 , n73442 );
xor ( n73444 , n73441 , n73442 );
xor ( n73445 , n73224 , n73288 );
and ( n73446 , n30359 , n73342 );
and ( n73447 , n73445 , n73446 );
xor ( n73448 , n73445 , n73446 );
xor ( n73449 , n73228 , n73286 );
and ( n73450 , n30364 , n73342 );
and ( n73451 , n73449 , n73450 );
xor ( n73452 , n73449 , n73450 );
xor ( n73453 , n73232 , n73284 );
and ( n73454 , n30369 , n73342 );
and ( n73455 , n73453 , n73454 );
xor ( n73456 , n73453 , n73454 );
xor ( n73457 , n73236 , n73282 );
and ( n73458 , n30374 , n73342 );
and ( n73459 , n73457 , n73458 );
xor ( n73460 , n73457 , n73458 );
xor ( n73461 , n73240 , n73280 );
and ( n73462 , n30379 , n73342 );
and ( n73463 , n73461 , n73462 );
xor ( n73464 , n73461 , n73462 );
xor ( n73465 , n73244 , n73278 );
and ( n73466 , n30384 , n73342 );
and ( n73467 , n73465 , n73466 );
xor ( n73468 , n73465 , n73466 );
xor ( n73469 , n73248 , n73276 );
and ( n73470 , n30389 , n73342 );
and ( n73471 , n73469 , n73470 );
xor ( n73472 , n73469 , n73470 );
xor ( n73473 , n73252 , n73274 );
and ( n73474 , n30394 , n73342 );
and ( n73475 , n73473 , n73474 );
xor ( n73476 , n73473 , n73474 );
xor ( n73477 , n73256 , n73272 );
and ( n73478 , n30399 , n73342 );
and ( n73479 , n73477 , n73478 );
xor ( n73480 , n73477 , n73478 );
xor ( n73481 , n73260 , n73270 );
and ( n73482 , n30404 , n73342 );
and ( n73483 , n73481 , n73482 );
xor ( n73484 , n73481 , n73482 );
xor ( n73485 , n73264 , n73268 );
and ( n73486 , n30409 , n73342 );
and ( n73487 , n73485 , n73486 );
buf ( n73488 , n73487 );
and ( n73489 , n73484 , n73488 );
or ( n73490 , n73483 , n73489 );
and ( n73491 , n73480 , n73490 );
or ( n73492 , n73479 , n73491 );
and ( n73493 , n73476 , n73492 );
or ( n73494 , n73475 , n73493 );
and ( n73495 , n73472 , n73494 );
or ( n73496 , n73471 , n73495 );
and ( n73497 , n73468 , n73496 );
or ( n73498 , n73467 , n73497 );
and ( n73499 , n73464 , n73498 );
or ( n73500 , n73463 , n73499 );
and ( n73501 , n73460 , n73500 );
or ( n73502 , n73459 , n73501 );
and ( n73503 , n73456 , n73502 );
or ( n73504 , n73455 , n73503 );
and ( n73505 , n73452 , n73504 );
or ( n73506 , n73451 , n73505 );
and ( n73507 , n73448 , n73506 );
or ( n73508 , n73447 , n73507 );
and ( n73509 , n73444 , n73508 );
or ( n73510 , n73443 , n73509 );
and ( n73511 , n73440 , n73510 );
or ( n73512 , n73439 , n73511 );
and ( n73513 , n73436 , n73512 );
or ( n73514 , n73435 , n73513 );
and ( n73515 , n73432 , n73514 );
or ( n73516 , n73431 , n73515 );
and ( n73517 , n73428 , n73516 );
or ( n73518 , n73427 , n73517 );
and ( n73519 , n73424 , n73518 );
or ( n73520 , n73423 , n73519 );
and ( n73521 , n73420 , n73520 );
or ( n73522 , n73419 , n73521 );
and ( n73523 , n73416 , n73522 );
or ( n73524 , n73415 , n73523 );
and ( n73525 , n73412 , n73524 );
or ( n73526 , n73411 , n73525 );
and ( n73527 , n73408 , n73526 );
or ( n73528 , n73407 , n73527 );
and ( n73529 , n73404 , n73528 );
or ( n73530 , n73403 , n73529 );
and ( n73531 , n73400 , n73530 );
or ( n73532 , n73399 , n73531 );
and ( n73533 , n73396 , n73532 );
or ( n73534 , n73395 , n73533 );
and ( n73535 , n73392 , n73534 );
or ( n73536 , n73391 , n73535 );
and ( n73537 , n73388 , n73536 );
or ( n73538 , n73387 , n73537 );
and ( n73539 , n73384 , n73538 );
or ( n73540 , n73383 , n73539 );
and ( n73541 , n73380 , n73540 );
or ( n73542 , n73379 , n73541 );
and ( n73543 , n73376 , n73542 );
or ( n73544 , n73375 , n73543 );
and ( n73545 , n73372 , n73544 );
or ( n73546 , n73371 , n73545 );
and ( n73547 , n73368 , n73546 );
or ( n73548 , n73367 , n73547 );
and ( n73549 , n73364 , n73548 );
or ( n73550 , n73363 , n73549 );
and ( n73551 , n73360 , n73550 );
or ( n73552 , n73359 , n73551 );
and ( n73553 , n73356 , n73552 );
or ( n73554 , n73355 , n73553 );
and ( n73555 , n73352 , n73554 );
or ( n73556 , n73351 , n73555 );
and ( n73557 , n73348 , n73556 );
or ( n73558 , n73347 , n73557 );
xor ( n73559 , n73344 , n73558 );
buf ( n73560 , n17924 );
and ( n73561 , n30234 , n73560 );
xor ( n73562 , n73559 , n73561 );
xor ( n73563 , n73348 , n73556 );
and ( n73564 , n30239 , n73560 );
and ( n73565 , n73563 , n73564 );
xor ( n73566 , n73563 , n73564 );
xor ( n73567 , n73352 , n73554 );
and ( n73568 , n30244 , n73560 );
and ( n73569 , n73567 , n73568 );
xor ( n73570 , n73567 , n73568 );
xor ( n73571 , n73356 , n73552 );
and ( n73572 , n30249 , n73560 );
and ( n73573 , n73571 , n73572 );
xor ( n73574 , n73571 , n73572 );
xor ( n73575 , n73360 , n73550 );
and ( n73576 , n30254 , n73560 );
and ( n73577 , n73575 , n73576 );
xor ( n73578 , n73575 , n73576 );
xor ( n73579 , n73364 , n73548 );
and ( n73580 , n30259 , n73560 );
and ( n73581 , n73579 , n73580 );
xor ( n73582 , n73579 , n73580 );
xor ( n73583 , n73368 , n73546 );
and ( n73584 , n30264 , n73560 );
and ( n73585 , n73583 , n73584 );
xor ( n73586 , n73583 , n73584 );
xor ( n73587 , n73372 , n73544 );
and ( n73588 , n30269 , n73560 );
and ( n73589 , n73587 , n73588 );
xor ( n73590 , n73587 , n73588 );
xor ( n73591 , n73376 , n73542 );
and ( n73592 , n30274 , n73560 );
and ( n73593 , n73591 , n73592 );
xor ( n73594 , n73591 , n73592 );
xor ( n73595 , n73380 , n73540 );
and ( n73596 , n30279 , n73560 );
and ( n73597 , n73595 , n73596 );
xor ( n73598 , n73595 , n73596 );
xor ( n73599 , n73384 , n73538 );
and ( n73600 , n30284 , n73560 );
and ( n73601 , n73599 , n73600 );
xor ( n73602 , n73599 , n73600 );
xor ( n73603 , n73388 , n73536 );
and ( n73604 , n30289 , n73560 );
and ( n73605 , n73603 , n73604 );
xor ( n73606 , n73603 , n73604 );
xor ( n73607 , n73392 , n73534 );
and ( n73608 , n30294 , n73560 );
and ( n73609 , n73607 , n73608 );
xor ( n73610 , n73607 , n73608 );
xor ( n73611 , n73396 , n73532 );
and ( n73612 , n30299 , n73560 );
and ( n73613 , n73611 , n73612 );
xor ( n73614 , n73611 , n73612 );
xor ( n73615 , n73400 , n73530 );
and ( n73616 , n30304 , n73560 );
and ( n73617 , n73615 , n73616 );
xor ( n73618 , n73615 , n73616 );
xor ( n73619 , n73404 , n73528 );
and ( n73620 , n30309 , n73560 );
and ( n73621 , n73619 , n73620 );
xor ( n73622 , n73619 , n73620 );
xor ( n73623 , n73408 , n73526 );
and ( n73624 , n30314 , n73560 );
and ( n73625 , n73623 , n73624 );
xor ( n73626 , n73623 , n73624 );
xor ( n73627 , n73412 , n73524 );
and ( n73628 , n30319 , n73560 );
and ( n73629 , n73627 , n73628 );
xor ( n73630 , n73627 , n73628 );
xor ( n73631 , n73416 , n73522 );
and ( n73632 , n30324 , n73560 );
and ( n73633 , n73631 , n73632 );
xor ( n73634 , n73631 , n73632 );
xor ( n73635 , n73420 , n73520 );
and ( n73636 , n30329 , n73560 );
and ( n73637 , n73635 , n73636 );
xor ( n73638 , n73635 , n73636 );
xor ( n73639 , n73424 , n73518 );
and ( n73640 , n30334 , n73560 );
and ( n73641 , n73639 , n73640 );
xor ( n73642 , n73639 , n73640 );
xor ( n73643 , n73428 , n73516 );
and ( n73644 , n30339 , n73560 );
and ( n73645 , n73643 , n73644 );
xor ( n73646 , n73643 , n73644 );
xor ( n73647 , n73432 , n73514 );
and ( n73648 , n30344 , n73560 );
and ( n73649 , n73647 , n73648 );
xor ( n73650 , n73647 , n73648 );
xor ( n73651 , n73436 , n73512 );
and ( n73652 , n30349 , n73560 );
and ( n73653 , n73651 , n73652 );
xor ( n73654 , n73651 , n73652 );
xor ( n73655 , n73440 , n73510 );
and ( n73656 , n30354 , n73560 );
and ( n73657 , n73655 , n73656 );
xor ( n73658 , n73655 , n73656 );
xor ( n73659 , n73444 , n73508 );
and ( n73660 , n30359 , n73560 );
and ( n73661 , n73659 , n73660 );
xor ( n73662 , n73659 , n73660 );
xor ( n73663 , n73448 , n73506 );
and ( n73664 , n30364 , n73560 );
and ( n73665 , n73663 , n73664 );
xor ( n73666 , n73663 , n73664 );
xor ( n73667 , n73452 , n73504 );
and ( n73668 , n30369 , n73560 );
and ( n73669 , n73667 , n73668 );
xor ( n73670 , n73667 , n73668 );
xor ( n73671 , n73456 , n73502 );
and ( n73672 , n30374 , n73560 );
and ( n73673 , n73671 , n73672 );
xor ( n73674 , n73671 , n73672 );
xor ( n73675 , n73460 , n73500 );
and ( n73676 , n30379 , n73560 );
and ( n73677 , n73675 , n73676 );
xor ( n73678 , n73675 , n73676 );
xor ( n73679 , n73464 , n73498 );
and ( n73680 , n30384 , n73560 );
and ( n73681 , n73679 , n73680 );
xor ( n73682 , n73679 , n73680 );
xor ( n73683 , n73468 , n73496 );
and ( n73684 , n30389 , n73560 );
and ( n73685 , n73683 , n73684 );
xor ( n73686 , n73683 , n73684 );
xor ( n73687 , n73472 , n73494 );
and ( n73688 , n30394 , n73560 );
and ( n73689 , n73687 , n73688 );
xor ( n73690 , n73687 , n73688 );
xor ( n73691 , n73476 , n73492 );
and ( n73692 , n30399 , n73560 );
and ( n73693 , n73691 , n73692 );
xor ( n73694 , n73691 , n73692 );
xor ( n73695 , n73480 , n73490 );
and ( n73696 , n30404 , n73560 );
and ( n73697 , n73695 , n73696 );
xor ( n73698 , n73695 , n73696 );
xor ( n73699 , n73484 , n73488 );
and ( n73700 , n30409 , n73560 );
and ( n73701 , n73699 , n73700 );
buf ( n73702 , n73701 );
and ( n73703 , n73698 , n73702 );
or ( n73704 , n73697 , n73703 );
and ( n73705 , n73694 , n73704 );
or ( n73706 , n73693 , n73705 );
and ( n73707 , n73690 , n73706 );
or ( n73708 , n73689 , n73707 );
and ( n73709 , n73686 , n73708 );
or ( n73710 , n73685 , n73709 );
and ( n73711 , n73682 , n73710 );
or ( n73712 , n73681 , n73711 );
and ( n73713 , n73678 , n73712 );
or ( n73714 , n73677 , n73713 );
and ( n73715 , n73674 , n73714 );
or ( n73716 , n73673 , n73715 );
and ( n73717 , n73670 , n73716 );
or ( n73718 , n73669 , n73717 );
and ( n73719 , n73666 , n73718 );
or ( n73720 , n73665 , n73719 );
and ( n73721 , n73662 , n73720 );
or ( n73722 , n73661 , n73721 );
and ( n73723 , n73658 , n73722 );
or ( n73724 , n73657 , n73723 );
and ( n73725 , n73654 , n73724 );
or ( n73726 , n73653 , n73725 );
and ( n73727 , n73650 , n73726 );
or ( n73728 , n73649 , n73727 );
and ( n73729 , n73646 , n73728 );
or ( n73730 , n73645 , n73729 );
and ( n73731 , n73642 , n73730 );
or ( n73732 , n73641 , n73731 );
and ( n73733 , n73638 , n73732 );
or ( n73734 , n73637 , n73733 );
and ( n73735 , n73634 , n73734 );
or ( n73736 , n73633 , n73735 );
and ( n73737 , n73630 , n73736 );
or ( n73738 , n73629 , n73737 );
and ( n73739 , n73626 , n73738 );
or ( n73740 , n73625 , n73739 );
and ( n73741 , n73622 , n73740 );
or ( n73742 , n73621 , n73741 );
and ( n73743 , n73618 , n73742 );
or ( n73744 , n73617 , n73743 );
and ( n73745 , n73614 , n73744 );
or ( n73746 , n73613 , n73745 );
and ( n73747 , n73610 , n73746 );
or ( n73748 , n73609 , n73747 );
and ( n73749 , n73606 , n73748 );
or ( n73750 , n73605 , n73749 );
and ( n73751 , n73602 , n73750 );
or ( n73752 , n73601 , n73751 );
and ( n73753 , n73598 , n73752 );
or ( n73754 , n73597 , n73753 );
and ( n73755 , n73594 , n73754 );
or ( n73756 , n73593 , n73755 );
and ( n73757 , n73590 , n73756 );
or ( n73758 , n73589 , n73757 );
and ( n73759 , n73586 , n73758 );
or ( n73760 , n73585 , n73759 );
and ( n73761 , n73582 , n73760 );
or ( n73762 , n73581 , n73761 );
and ( n73763 , n73578 , n73762 );
or ( n73764 , n73577 , n73763 );
and ( n73765 , n73574 , n73764 );
or ( n73766 , n73573 , n73765 );
and ( n73767 , n73570 , n73766 );
or ( n73768 , n73569 , n73767 );
and ( n73769 , n73566 , n73768 );
or ( n73770 , n73565 , n73769 );
xor ( n73771 , n73562 , n73770 );
buf ( n73772 , n17922 );
and ( n73773 , n30239 , n73772 );
xor ( n73774 , n73771 , n73773 );
xor ( n73775 , n73566 , n73768 );
and ( n73776 , n30244 , n73772 );
and ( n73777 , n73775 , n73776 );
xor ( n73778 , n73775 , n73776 );
xor ( n73779 , n73570 , n73766 );
and ( n73780 , n30249 , n73772 );
and ( n73781 , n73779 , n73780 );
xor ( n73782 , n73779 , n73780 );
xor ( n73783 , n73574 , n73764 );
and ( n73784 , n30254 , n73772 );
and ( n73785 , n73783 , n73784 );
xor ( n73786 , n73783 , n73784 );
xor ( n73787 , n73578 , n73762 );
and ( n73788 , n30259 , n73772 );
and ( n73789 , n73787 , n73788 );
xor ( n73790 , n73787 , n73788 );
xor ( n73791 , n73582 , n73760 );
and ( n73792 , n30264 , n73772 );
and ( n73793 , n73791 , n73792 );
xor ( n73794 , n73791 , n73792 );
xor ( n73795 , n73586 , n73758 );
and ( n73796 , n30269 , n73772 );
and ( n73797 , n73795 , n73796 );
xor ( n73798 , n73795 , n73796 );
xor ( n73799 , n73590 , n73756 );
and ( n73800 , n30274 , n73772 );
and ( n73801 , n73799 , n73800 );
xor ( n73802 , n73799 , n73800 );
xor ( n73803 , n73594 , n73754 );
and ( n73804 , n30279 , n73772 );
and ( n73805 , n73803 , n73804 );
xor ( n73806 , n73803 , n73804 );
xor ( n73807 , n73598 , n73752 );
and ( n73808 , n30284 , n73772 );
and ( n73809 , n73807 , n73808 );
xor ( n73810 , n73807 , n73808 );
xor ( n73811 , n73602 , n73750 );
and ( n73812 , n30289 , n73772 );
and ( n73813 , n73811 , n73812 );
xor ( n73814 , n73811 , n73812 );
xor ( n73815 , n73606 , n73748 );
and ( n73816 , n30294 , n73772 );
and ( n73817 , n73815 , n73816 );
xor ( n73818 , n73815 , n73816 );
xor ( n73819 , n73610 , n73746 );
and ( n73820 , n30299 , n73772 );
and ( n73821 , n73819 , n73820 );
xor ( n73822 , n73819 , n73820 );
xor ( n73823 , n73614 , n73744 );
and ( n73824 , n30304 , n73772 );
and ( n73825 , n73823 , n73824 );
xor ( n73826 , n73823 , n73824 );
xor ( n73827 , n73618 , n73742 );
and ( n73828 , n30309 , n73772 );
and ( n73829 , n73827 , n73828 );
xor ( n73830 , n73827 , n73828 );
xor ( n73831 , n73622 , n73740 );
and ( n73832 , n30314 , n73772 );
and ( n73833 , n73831 , n73832 );
xor ( n73834 , n73831 , n73832 );
xor ( n73835 , n73626 , n73738 );
and ( n73836 , n30319 , n73772 );
and ( n73837 , n73835 , n73836 );
xor ( n73838 , n73835 , n73836 );
xor ( n73839 , n73630 , n73736 );
and ( n73840 , n30324 , n73772 );
and ( n73841 , n73839 , n73840 );
xor ( n73842 , n73839 , n73840 );
xor ( n73843 , n73634 , n73734 );
and ( n73844 , n30329 , n73772 );
and ( n73845 , n73843 , n73844 );
xor ( n73846 , n73843 , n73844 );
xor ( n73847 , n73638 , n73732 );
and ( n73848 , n30334 , n73772 );
and ( n73849 , n73847 , n73848 );
xor ( n73850 , n73847 , n73848 );
xor ( n73851 , n73642 , n73730 );
and ( n73852 , n30339 , n73772 );
and ( n73853 , n73851 , n73852 );
xor ( n73854 , n73851 , n73852 );
xor ( n73855 , n73646 , n73728 );
and ( n73856 , n30344 , n73772 );
and ( n73857 , n73855 , n73856 );
xor ( n73858 , n73855 , n73856 );
xor ( n73859 , n73650 , n73726 );
and ( n73860 , n30349 , n73772 );
and ( n73861 , n73859 , n73860 );
xor ( n73862 , n73859 , n73860 );
xor ( n73863 , n73654 , n73724 );
and ( n73864 , n30354 , n73772 );
and ( n73865 , n73863 , n73864 );
xor ( n73866 , n73863 , n73864 );
xor ( n73867 , n73658 , n73722 );
and ( n73868 , n30359 , n73772 );
and ( n73869 , n73867 , n73868 );
xor ( n73870 , n73867 , n73868 );
xor ( n73871 , n73662 , n73720 );
and ( n73872 , n30364 , n73772 );
and ( n73873 , n73871 , n73872 );
xor ( n73874 , n73871 , n73872 );
xor ( n73875 , n73666 , n73718 );
and ( n73876 , n30369 , n73772 );
and ( n73877 , n73875 , n73876 );
xor ( n73878 , n73875 , n73876 );
xor ( n73879 , n73670 , n73716 );
and ( n73880 , n30374 , n73772 );
and ( n73881 , n73879 , n73880 );
xor ( n73882 , n73879 , n73880 );
xor ( n73883 , n73674 , n73714 );
and ( n73884 , n30379 , n73772 );
and ( n73885 , n73883 , n73884 );
xor ( n73886 , n73883 , n73884 );
xor ( n73887 , n73678 , n73712 );
and ( n73888 , n30384 , n73772 );
and ( n73889 , n73887 , n73888 );
xor ( n73890 , n73887 , n73888 );
xor ( n73891 , n73682 , n73710 );
and ( n73892 , n30389 , n73772 );
and ( n73893 , n73891 , n73892 );
xor ( n73894 , n73891 , n73892 );
xor ( n73895 , n73686 , n73708 );
and ( n73896 , n30394 , n73772 );
and ( n73897 , n73895 , n73896 );
xor ( n73898 , n73895 , n73896 );
xor ( n73899 , n73690 , n73706 );
and ( n73900 , n30399 , n73772 );
and ( n73901 , n73899 , n73900 );
xor ( n73902 , n73899 , n73900 );
xor ( n73903 , n73694 , n73704 );
and ( n73904 , n30404 , n73772 );
and ( n73905 , n73903 , n73904 );
xor ( n73906 , n73903 , n73904 );
xor ( n73907 , n73698 , n73702 );
and ( n73908 , n30409 , n73772 );
and ( n73909 , n73907 , n73908 );
buf ( n73910 , n73909 );
and ( n73911 , n73906 , n73910 );
or ( n73912 , n73905 , n73911 );
and ( n73913 , n73902 , n73912 );
or ( n73914 , n73901 , n73913 );
and ( n73915 , n73898 , n73914 );
or ( n73916 , n73897 , n73915 );
and ( n73917 , n73894 , n73916 );
or ( n73918 , n73893 , n73917 );
and ( n73919 , n73890 , n73918 );
or ( n73920 , n73889 , n73919 );
and ( n73921 , n73886 , n73920 );
or ( n73922 , n73885 , n73921 );
and ( n73923 , n73882 , n73922 );
or ( n73924 , n73881 , n73923 );
and ( n73925 , n73878 , n73924 );
or ( n73926 , n73877 , n73925 );
and ( n73927 , n73874 , n73926 );
or ( n73928 , n73873 , n73927 );
and ( n73929 , n73870 , n73928 );
or ( n73930 , n73869 , n73929 );
and ( n73931 , n73866 , n73930 );
or ( n73932 , n73865 , n73931 );
and ( n73933 , n73862 , n73932 );
or ( n73934 , n73861 , n73933 );
and ( n73935 , n73858 , n73934 );
or ( n73936 , n73857 , n73935 );
and ( n73937 , n73854 , n73936 );
or ( n73938 , n73853 , n73937 );
and ( n73939 , n73850 , n73938 );
or ( n73940 , n73849 , n73939 );
and ( n73941 , n73846 , n73940 );
or ( n73942 , n73845 , n73941 );
and ( n73943 , n73842 , n73942 );
or ( n73944 , n73841 , n73943 );
and ( n73945 , n73838 , n73944 );
or ( n73946 , n73837 , n73945 );
and ( n73947 , n73834 , n73946 );
or ( n73948 , n73833 , n73947 );
and ( n73949 , n73830 , n73948 );
or ( n73950 , n73829 , n73949 );
and ( n73951 , n73826 , n73950 );
or ( n73952 , n73825 , n73951 );
and ( n73953 , n73822 , n73952 );
or ( n73954 , n73821 , n73953 );
and ( n73955 , n73818 , n73954 );
or ( n73956 , n73817 , n73955 );
and ( n73957 , n73814 , n73956 );
or ( n73958 , n73813 , n73957 );
and ( n73959 , n73810 , n73958 );
or ( n73960 , n73809 , n73959 );
and ( n73961 , n73806 , n73960 );
or ( n73962 , n73805 , n73961 );
and ( n73963 , n73802 , n73962 );
or ( n73964 , n73801 , n73963 );
and ( n73965 , n73798 , n73964 );
or ( n73966 , n73797 , n73965 );
and ( n73967 , n73794 , n73966 );
or ( n73968 , n73793 , n73967 );
and ( n73969 , n73790 , n73968 );
or ( n73970 , n73789 , n73969 );
and ( n73971 , n73786 , n73970 );
or ( n73972 , n73785 , n73971 );
and ( n73973 , n73782 , n73972 );
or ( n73974 , n73781 , n73973 );
and ( n73975 , n73778 , n73974 );
or ( n73976 , n73777 , n73975 );
xor ( n73977 , n73774 , n73976 );
buf ( n73978 , n17920 );
and ( n73979 , n30244 , n73978 );
xor ( n73980 , n73977 , n73979 );
xor ( n73981 , n73778 , n73974 );
and ( n73982 , n30249 , n73978 );
and ( n73983 , n73981 , n73982 );
xor ( n73984 , n73981 , n73982 );
xor ( n73985 , n73782 , n73972 );
and ( n73986 , n30254 , n73978 );
and ( n73987 , n73985 , n73986 );
xor ( n73988 , n73985 , n73986 );
xor ( n73989 , n73786 , n73970 );
and ( n73990 , n30259 , n73978 );
and ( n73991 , n73989 , n73990 );
xor ( n73992 , n73989 , n73990 );
xor ( n73993 , n73790 , n73968 );
and ( n73994 , n30264 , n73978 );
and ( n73995 , n73993 , n73994 );
xor ( n73996 , n73993 , n73994 );
xor ( n73997 , n73794 , n73966 );
and ( n73998 , n30269 , n73978 );
and ( n73999 , n73997 , n73998 );
xor ( n74000 , n73997 , n73998 );
xor ( n74001 , n73798 , n73964 );
and ( n74002 , n30274 , n73978 );
and ( n74003 , n74001 , n74002 );
xor ( n74004 , n74001 , n74002 );
xor ( n74005 , n73802 , n73962 );
and ( n74006 , n30279 , n73978 );
and ( n74007 , n74005 , n74006 );
xor ( n74008 , n74005 , n74006 );
xor ( n74009 , n73806 , n73960 );
and ( n74010 , n30284 , n73978 );
and ( n74011 , n74009 , n74010 );
xor ( n74012 , n74009 , n74010 );
xor ( n74013 , n73810 , n73958 );
and ( n74014 , n30289 , n73978 );
and ( n74015 , n74013 , n74014 );
xor ( n74016 , n74013 , n74014 );
xor ( n74017 , n73814 , n73956 );
and ( n74018 , n30294 , n73978 );
and ( n74019 , n74017 , n74018 );
xor ( n74020 , n74017 , n74018 );
xor ( n74021 , n73818 , n73954 );
and ( n74022 , n30299 , n73978 );
and ( n74023 , n74021 , n74022 );
xor ( n74024 , n74021 , n74022 );
xor ( n74025 , n73822 , n73952 );
and ( n74026 , n30304 , n73978 );
and ( n74027 , n74025 , n74026 );
xor ( n74028 , n74025 , n74026 );
xor ( n74029 , n73826 , n73950 );
and ( n74030 , n30309 , n73978 );
and ( n74031 , n74029 , n74030 );
xor ( n74032 , n74029 , n74030 );
xor ( n74033 , n73830 , n73948 );
and ( n74034 , n30314 , n73978 );
and ( n74035 , n74033 , n74034 );
xor ( n74036 , n74033 , n74034 );
xor ( n74037 , n73834 , n73946 );
and ( n74038 , n30319 , n73978 );
and ( n74039 , n74037 , n74038 );
xor ( n74040 , n74037 , n74038 );
xor ( n74041 , n73838 , n73944 );
and ( n74042 , n30324 , n73978 );
and ( n74043 , n74041 , n74042 );
xor ( n74044 , n74041 , n74042 );
xor ( n74045 , n73842 , n73942 );
and ( n74046 , n30329 , n73978 );
and ( n74047 , n74045 , n74046 );
xor ( n74048 , n74045 , n74046 );
xor ( n74049 , n73846 , n73940 );
and ( n74050 , n30334 , n73978 );
and ( n74051 , n74049 , n74050 );
xor ( n74052 , n74049 , n74050 );
xor ( n74053 , n73850 , n73938 );
and ( n74054 , n30339 , n73978 );
and ( n74055 , n74053 , n74054 );
xor ( n74056 , n74053 , n74054 );
xor ( n74057 , n73854 , n73936 );
and ( n74058 , n30344 , n73978 );
and ( n74059 , n74057 , n74058 );
xor ( n74060 , n74057 , n74058 );
xor ( n74061 , n73858 , n73934 );
and ( n74062 , n30349 , n73978 );
and ( n74063 , n74061 , n74062 );
xor ( n74064 , n74061 , n74062 );
xor ( n74065 , n73862 , n73932 );
and ( n74066 , n30354 , n73978 );
and ( n74067 , n74065 , n74066 );
xor ( n74068 , n74065 , n74066 );
xor ( n74069 , n73866 , n73930 );
and ( n74070 , n30359 , n73978 );
and ( n74071 , n74069 , n74070 );
xor ( n74072 , n74069 , n74070 );
xor ( n74073 , n73870 , n73928 );
and ( n74074 , n30364 , n73978 );
and ( n74075 , n74073 , n74074 );
xor ( n74076 , n74073 , n74074 );
xor ( n74077 , n73874 , n73926 );
and ( n74078 , n30369 , n73978 );
and ( n74079 , n74077 , n74078 );
xor ( n74080 , n74077 , n74078 );
xor ( n74081 , n73878 , n73924 );
and ( n74082 , n30374 , n73978 );
and ( n74083 , n74081 , n74082 );
xor ( n74084 , n74081 , n74082 );
xor ( n74085 , n73882 , n73922 );
and ( n74086 , n30379 , n73978 );
and ( n74087 , n74085 , n74086 );
xor ( n74088 , n74085 , n74086 );
xor ( n74089 , n73886 , n73920 );
and ( n74090 , n30384 , n73978 );
and ( n74091 , n74089 , n74090 );
xor ( n74092 , n74089 , n74090 );
xor ( n74093 , n73890 , n73918 );
and ( n74094 , n30389 , n73978 );
and ( n74095 , n74093 , n74094 );
xor ( n74096 , n74093 , n74094 );
xor ( n74097 , n73894 , n73916 );
and ( n74098 , n30394 , n73978 );
and ( n74099 , n74097 , n74098 );
xor ( n74100 , n74097 , n74098 );
xor ( n74101 , n73898 , n73914 );
and ( n74102 , n30399 , n73978 );
and ( n74103 , n74101 , n74102 );
xor ( n74104 , n74101 , n74102 );
xor ( n74105 , n73902 , n73912 );
and ( n74106 , n30404 , n73978 );
and ( n74107 , n74105 , n74106 );
xor ( n74108 , n74105 , n74106 );
xor ( n74109 , n73906 , n73910 );
and ( n74110 , n30409 , n73978 );
and ( n74111 , n74109 , n74110 );
buf ( n74112 , n74111 );
and ( n74113 , n74108 , n74112 );
or ( n74114 , n74107 , n74113 );
and ( n74115 , n74104 , n74114 );
or ( n74116 , n74103 , n74115 );
and ( n74117 , n74100 , n74116 );
or ( n74118 , n74099 , n74117 );
and ( n74119 , n74096 , n74118 );
or ( n74120 , n74095 , n74119 );
and ( n74121 , n74092 , n74120 );
or ( n74122 , n74091 , n74121 );
and ( n74123 , n74088 , n74122 );
or ( n74124 , n74087 , n74123 );
and ( n74125 , n74084 , n74124 );
or ( n74126 , n74083 , n74125 );
and ( n74127 , n74080 , n74126 );
or ( n74128 , n74079 , n74127 );
and ( n74129 , n74076 , n74128 );
or ( n74130 , n74075 , n74129 );
and ( n74131 , n74072 , n74130 );
or ( n74132 , n74071 , n74131 );
and ( n74133 , n74068 , n74132 );
or ( n74134 , n74067 , n74133 );
and ( n74135 , n74064 , n74134 );
or ( n74136 , n74063 , n74135 );
and ( n74137 , n74060 , n74136 );
or ( n74138 , n74059 , n74137 );
and ( n74139 , n74056 , n74138 );
or ( n74140 , n74055 , n74139 );
and ( n74141 , n74052 , n74140 );
or ( n74142 , n74051 , n74141 );
and ( n74143 , n74048 , n74142 );
or ( n74144 , n74047 , n74143 );
and ( n74145 , n74044 , n74144 );
or ( n74146 , n74043 , n74145 );
and ( n74147 , n74040 , n74146 );
or ( n74148 , n74039 , n74147 );
and ( n74149 , n74036 , n74148 );
or ( n74150 , n74035 , n74149 );
and ( n74151 , n74032 , n74150 );
or ( n74152 , n74031 , n74151 );
and ( n74153 , n74028 , n74152 );
or ( n74154 , n74027 , n74153 );
and ( n74155 , n74024 , n74154 );
or ( n74156 , n74023 , n74155 );
and ( n74157 , n74020 , n74156 );
or ( n74158 , n74019 , n74157 );
and ( n74159 , n74016 , n74158 );
or ( n74160 , n74015 , n74159 );
and ( n74161 , n74012 , n74160 );
or ( n74162 , n74011 , n74161 );
and ( n74163 , n74008 , n74162 );
or ( n74164 , n74007 , n74163 );
and ( n74165 , n74004 , n74164 );
or ( n74166 , n74003 , n74165 );
and ( n74167 , n74000 , n74166 );
or ( n74168 , n73999 , n74167 );
and ( n74169 , n73996 , n74168 );
or ( n74170 , n73995 , n74169 );
and ( n74171 , n73992 , n74170 );
or ( n74172 , n73991 , n74171 );
and ( n74173 , n73988 , n74172 );
or ( n74174 , n73987 , n74173 );
and ( n74175 , n73984 , n74174 );
or ( n74176 , n73983 , n74175 );
xor ( n74177 , n73980 , n74176 );
buf ( n74178 , n17918 );
and ( n74179 , n30249 , n74178 );
xor ( n74180 , n74177 , n74179 );
xor ( n74181 , n73984 , n74174 );
and ( n74182 , n30254 , n74178 );
and ( n74183 , n74181 , n74182 );
xor ( n74184 , n74181 , n74182 );
xor ( n74185 , n73988 , n74172 );
and ( n74186 , n30259 , n74178 );
and ( n74187 , n74185 , n74186 );
xor ( n74188 , n74185 , n74186 );
xor ( n74189 , n73992 , n74170 );
and ( n74190 , n30264 , n74178 );
and ( n74191 , n74189 , n74190 );
xor ( n74192 , n74189 , n74190 );
xor ( n74193 , n73996 , n74168 );
and ( n74194 , n30269 , n74178 );
and ( n74195 , n74193 , n74194 );
xor ( n74196 , n74193 , n74194 );
xor ( n74197 , n74000 , n74166 );
and ( n74198 , n30274 , n74178 );
and ( n74199 , n74197 , n74198 );
xor ( n74200 , n74197 , n74198 );
xor ( n74201 , n74004 , n74164 );
and ( n74202 , n30279 , n74178 );
and ( n74203 , n74201 , n74202 );
xor ( n74204 , n74201 , n74202 );
xor ( n74205 , n74008 , n74162 );
and ( n74206 , n30284 , n74178 );
and ( n74207 , n74205 , n74206 );
xor ( n74208 , n74205 , n74206 );
xor ( n74209 , n74012 , n74160 );
and ( n74210 , n30289 , n74178 );
and ( n74211 , n74209 , n74210 );
xor ( n74212 , n74209 , n74210 );
xor ( n74213 , n74016 , n74158 );
and ( n74214 , n30294 , n74178 );
and ( n74215 , n74213 , n74214 );
xor ( n74216 , n74213 , n74214 );
xor ( n74217 , n74020 , n74156 );
and ( n74218 , n30299 , n74178 );
and ( n74219 , n74217 , n74218 );
xor ( n74220 , n74217 , n74218 );
xor ( n74221 , n74024 , n74154 );
and ( n74222 , n30304 , n74178 );
and ( n74223 , n74221 , n74222 );
xor ( n74224 , n74221 , n74222 );
xor ( n74225 , n74028 , n74152 );
and ( n74226 , n30309 , n74178 );
and ( n74227 , n74225 , n74226 );
xor ( n74228 , n74225 , n74226 );
xor ( n74229 , n74032 , n74150 );
and ( n74230 , n30314 , n74178 );
and ( n74231 , n74229 , n74230 );
xor ( n74232 , n74229 , n74230 );
xor ( n74233 , n74036 , n74148 );
and ( n74234 , n30319 , n74178 );
and ( n74235 , n74233 , n74234 );
xor ( n74236 , n74233 , n74234 );
xor ( n74237 , n74040 , n74146 );
and ( n74238 , n30324 , n74178 );
and ( n74239 , n74237 , n74238 );
xor ( n74240 , n74237 , n74238 );
xor ( n74241 , n74044 , n74144 );
and ( n74242 , n30329 , n74178 );
and ( n74243 , n74241 , n74242 );
xor ( n74244 , n74241 , n74242 );
xor ( n74245 , n74048 , n74142 );
and ( n74246 , n30334 , n74178 );
and ( n74247 , n74245 , n74246 );
xor ( n74248 , n74245 , n74246 );
xor ( n74249 , n74052 , n74140 );
and ( n74250 , n30339 , n74178 );
and ( n74251 , n74249 , n74250 );
xor ( n74252 , n74249 , n74250 );
xor ( n74253 , n74056 , n74138 );
and ( n74254 , n30344 , n74178 );
and ( n74255 , n74253 , n74254 );
xor ( n74256 , n74253 , n74254 );
xor ( n74257 , n74060 , n74136 );
and ( n74258 , n30349 , n74178 );
and ( n74259 , n74257 , n74258 );
xor ( n74260 , n74257 , n74258 );
xor ( n74261 , n74064 , n74134 );
and ( n74262 , n30354 , n74178 );
and ( n74263 , n74261 , n74262 );
xor ( n74264 , n74261 , n74262 );
xor ( n74265 , n74068 , n74132 );
and ( n74266 , n30359 , n74178 );
and ( n74267 , n74265 , n74266 );
xor ( n74268 , n74265 , n74266 );
xor ( n74269 , n74072 , n74130 );
and ( n74270 , n30364 , n74178 );
and ( n74271 , n74269 , n74270 );
xor ( n74272 , n74269 , n74270 );
xor ( n74273 , n74076 , n74128 );
and ( n74274 , n30369 , n74178 );
and ( n74275 , n74273 , n74274 );
xor ( n74276 , n74273 , n74274 );
xor ( n74277 , n74080 , n74126 );
and ( n74278 , n30374 , n74178 );
and ( n74279 , n74277 , n74278 );
xor ( n74280 , n74277 , n74278 );
xor ( n74281 , n74084 , n74124 );
and ( n74282 , n30379 , n74178 );
and ( n74283 , n74281 , n74282 );
xor ( n74284 , n74281 , n74282 );
xor ( n74285 , n74088 , n74122 );
and ( n74286 , n30384 , n74178 );
and ( n74287 , n74285 , n74286 );
xor ( n74288 , n74285 , n74286 );
xor ( n74289 , n74092 , n74120 );
and ( n74290 , n30389 , n74178 );
and ( n74291 , n74289 , n74290 );
xor ( n74292 , n74289 , n74290 );
xor ( n74293 , n74096 , n74118 );
and ( n74294 , n30394 , n74178 );
and ( n74295 , n74293 , n74294 );
xor ( n74296 , n74293 , n74294 );
xor ( n74297 , n74100 , n74116 );
and ( n74298 , n30399 , n74178 );
and ( n74299 , n74297 , n74298 );
xor ( n74300 , n74297 , n74298 );
xor ( n74301 , n74104 , n74114 );
and ( n74302 , n30404 , n74178 );
and ( n74303 , n74301 , n74302 );
xor ( n74304 , n74301 , n74302 );
xor ( n74305 , n74108 , n74112 );
and ( n74306 , n30409 , n74178 );
and ( n74307 , n74305 , n74306 );
buf ( n74308 , n74307 );
and ( n74309 , n74304 , n74308 );
or ( n74310 , n74303 , n74309 );
and ( n74311 , n74300 , n74310 );
or ( n74312 , n74299 , n74311 );
and ( n74313 , n74296 , n74312 );
or ( n74314 , n74295 , n74313 );
and ( n74315 , n74292 , n74314 );
or ( n74316 , n74291 , n74315 );
and ( n74317 , n74288 , n74316 );
or ( n74318 , n74287 , n74317 );
and ( n74319 , n74284 , n74318 );
or ( n74320 , n74283 , n74319 );
and ( n74321 , n74280 , n74320 );
or ( n74322 , n74279 , n74321 );
and ( n74323 , n74276 , n74322 );
or ( n74324 , n74275 , n74323 );
and ( n74325 , n74272 , n74324 );
or ( n74326 , n74271 , n74325 );
and ( n74327 , n74268 , n74326 );
or ( n74328 , n74267 , n74327 );
and ( n74329 , n74264 , n74328 );
or ( n74330 , n74263 , n74329 );
and ( n74331 , n74260 , n74330 );
or ( n74332 , n74259 , n74331 );
and ( n74333 , n74256 , n74332 );
or ( n74334 , n74255 , n74333 );
and ( n74335 , n74252 , n74334 );
or ( n74336 , n74251 , n74335 );
and ( n74337 , n74248 , n74336 );
or ( n74338 , n74247 , n74337 );
and ( n74339 , n74244 , n74338 );
or ( n74340 , n74243 , n74339 );
and ( n74341 , n74240 , n74340 );
or ( n74342 , n74239 , n74341 );
and ( n74343 , n74236 , n74342 );
or ( n74344 , n74235 , n74343 );
and ( n74345 , n74232 , n74344 );
or ( n74346 , n74231 , n74345 );
and ( n74347 , n74228 , n74346 );
or ( n74348 , n74227 , n74347 );
and ( n74349 , n74224 , n74348 );
or ( n74350 , n74223 , n74349 );
and ( n74351 , n74220 , n74350 );
or ( n74352 , n74219 , n74351 );
and ( n74353 , n74216 , n74352 );
or ( n74354 , n74215 , n74353 );
and ( n74355 , n74212 , n74354 );
or ( n74356 , n74211 , n74355 );
and ( n74357 , n74208 , n74356 );
or ( n74358 , n74207 , n74357 );
and ( n74359 , n74204 , n74358 );
or ( n74360 , n74203 , n74359 );
and ( n74361 , n74200 , n74360 );
or ( n74362 , n74199 , n74361 );
and ( n74363 , n74196 , n74362 );
or ( n74364 , n74195 , n74363 );
and ( n74365 , n74192 , n74364 );
or ( n74366 , n74191 , n74365 );
and ( n74367 , n74188 , n74366 );
or ( n74368 , n74187 , n74367 );
and ( n74369 , n74184 , n74368 );
or ( n74370 , n74183 , n74369 );
xor ( n74371 , n74180 , n74370 );
buf ( n74372 , n17916 );
and ( n74373 , n30254 , n74372 );
xor ( n74374 , n74371 , n74373 );
xor ( n74375 , n74184 , n74368 );
and ( n74376 , n30259 , n74372 );
and ( n74377 , n74375 , n74376 );
xor ( n74378 , n74375 , n74376 );
xor ( n74379 , n74188 , n74366 );
and ( n74380 , n30264 , n74372 );
and ( n74381 , n74379 , n74380 );
xor ( n74382 , n74379 , n74380 );
xor ( n74383 , n74192 , n74364 );
and ( n74384 , n30269 , n74372 );
and ( n74385 , n74383 , n74384 );
xor ( n74386 , n74383 , n74384 );
xor ( n74387 , n74196 , n74362 );
and ( n74388 , n30274 , n74372 );
and ( n74389 , n74387 , n74388 );
xor ( n74390 , n74387 , n74388 );
xor ( n74391 , n74200 , n74360 );
and ( n74392 , n30279 , n74372 );
and ( n74393 , n74391 , n74392 );
xor ( n74394 , n74391 , n74392 );
xor ( n74395 , n74204 , n74358 );
and ( n74396 , n30284 , n74372 );
and ( n74397 , n74395 , n74396 );
xor ( n74398 , n74395 , n74396 );
xor ( n74399 , n74208 , n74356 );
and ( n74400 , n30289 , n74372 );
and ( n74401 , n74399 , n74400 );
xor ( n74402 , n74399 , n74400 );
xor ( n74403 , n74212 , n74354 );
and ( n74404 , n30294 , n74372 );
and ( n74405 , n74403 , n74404 );
xor ( n74406 , n74403 , n74404 );
xor ( n74407 , n74216 , n74352 );
and ( n74408 , n30299 , n74372 );
and ( n74409 , n74407 , n74408 );
xor ( n74410 , n74407 , n74408 );
xor ( n74411 , n74220 , n74350 );
and ( n74412 , n30304 , n74372 );
and ( n74413 , n74411 , n74412 );
xor ( n74414 , n74411 , n74412 );
xor ( n74415 , n74224 , n74348 );
and ( n74416 , n30309 , n74372 );
and ( n74417 , n74415 , n74416 );
xor ( n74418 , n74415 , n74416 );
xor ( n74419 , n74228 , n74346 );
and ( n74420 , n30314 , n74372 );
and ( n74421 , n74419 , n74420 );
xor ( n74422 , n74419 , n74420 );
xor ( n74423 , n74232 , n74344 );
and ( n74424 , n30319 , n74372 );
and ( n74425 , n74423 , n74424 );
xor ( n74426 , n74423 , n74424 );
xor ( n74427 , n74236 , n74342 );
and ( n74428 , n30324 , n74372 );
and ( n74429 , n74427 , n74428 );
xor ( n74430 , n74427 , n74428 );
xor ( n74431 , n74240 , n74340 );
and ( n74432 , n30329 , n74372 );
and ( n74433 , n74431 , n74432 );
xor ( n74434 , n74431 , n74432 );
xor ( n74435 , n74244 , n74338 );
and ( n74436 , n30334 , n74372 );
and ( n74437 , n74435 , n74436 );
xor ( n74438 , n74435 , n74436 );
xor ( n74439 , n74248 , n74336 );
and ( n74440 , n30339 , n74372 );
and ( n74441 , n74439 , n74440 );
xor ( n74442 , n74439 , n74440 );
xor ( n74443 , n74252 , n74334 );
and ( n74444 , n30344 , n74372 );
and ( n74445 , n74443 , n74444 );
xor ( n74446 , n74443 , n74444 );
xor ( n74447 , n74256 , n74332 );
and ( n74448 , n30349 , n74372 );
and ( n74449 , n74447 , n74448 );
xor ( n74450 , n74447 , n74448 );
xor ( n74451 , n74260 , n74330 );
and ( n74452 , n30354 , n74372 );
and ( n74453 , n74451 , n74452 );
xor ( n74454 , n74451 , n74452 );
xor ( n74455 , n74264 , n74328 );
and ( n74456 , n30359 , n74372 );
and ( n74457 , n74455 , n74456 );
xor ( n74458 , n74455 , n74456 );
xor ( n74459 , n74268 , n74326 );
and ( n74460 , n30364 , n74372 );
and ( n74461 , n74459 , n74460 );
xor ( n74462 , n74459 , n74460 );
xor ( n74463 , n74272 , n74324 );
and ( n74464 , n30369 , n74372 );
and ( n74465 , n74463 , n74464 );
xor ( n74466 , n74463 , n74464 );
xor ( n74467 , n74276 , n74322 );
and ( n74468 , n30374 , n74372 );
and ( n74469 , n74467 , n74468 );
xor ( n74470 , n74467 , n74468 );
xor ( n74471 , n74280 , n74320 );
and ( n74472 , n30379 , n74372 );
and ( n74473 , n74471 , n74472 );
xor ( n74474 , n74471 , n74472 );
xor ( n74475 , n74284 , n74318 );
and ( n74476 , n30384 , n74372 );
and ( n74477 , n74475 , n74476 );
xor ( n74478 , n74475 , n74476 );
xor ( n74479 , n74288 , n74316 );
and ( n74480 , n30389 , n74372 );
and ( n74481 , n74479 , n74480 );
xor ( n74482 , n74479 , n74480 );
xor ( n74483 , n74292 , n74314 );
and ( n74484 , n30394 , n74372 );
and ( n74485 , n74483 , n74484 );
xor ( n74486 , n74483 , n74484 );
xor ( n74487 , n74296 , n74312 );
and ( n74488 , n30399 , n74372 );
and ( n74489 , n74487 , n74488 );
xor ( n74490 , n74487 , n74488 );
xor ( n74491 , n74300 , n74310 );
and ( n74492 , n30404 , n74372 );
and ( n74493 , n74491 , n74492 );
xor ( n74494 , n74491 , n74492 );
xor ( n74495 , n74304 , n74308 );
and ( n74496 , n30409 , n74372 );
and ( n74497 , n74495 , n74496 );
buf ( n74498 , n74497 );
and ( n74499 , n74494 , n74498 );
or ( n74500 , n74493 , n74499 );
and ( n74501 , n74490 , n74500 );
or ( n74502 , n74489 , n74501 );
and ( n74503 , n74486 , n74502 );
or ( n74504 , n74485 , n74503 );
and ( n74505 , n74482 , n74504 );
or ( n74506 , n74481 , n74505 );
and ( n74507 , n74478 , n74506 );
or ( n74508 , n74477 , n74507 );
and ( n74509 , n74474 , n74508 );
or ( n74510 , n74473 , n74509 );
and ( n74511 , n74470 , n74510 );
or ( n74512 , n74469 , n74511 );
and ( n74513 , n74466 , n74512 );
or ( n74514 , n74465 , n74513 );
and ( n74515 , n74462 , n74514 );
or ( n74516 , n74461 , n74515 );
and ( n74517 , n74458 , n74516 );
or ( n74518 , n74457 , n74517 );
and ( n74519 , n74454 , n74518 );
or ( n74520 , n74453 , n74519 );
and ( n74521 , n74450 , n74520 );
or ( n74522 , n74449 , n74521 );
and ( n74523 , n74446 , n74522 );
or ( n74524 , n74445 , n74523 );
and ( n74525 , n74442 , n74524 );
or ( n74526 , n74441 , n74525 );
and ( n74527 , n74438 , n74526 );
or ( n74528 , n74437 , n74527 );
and ( n74529 , n74434 , n74528 );
or ( n74530 , n74433 , n74529 );
and ( n74531 , n74430 , n74530 );
or ( n74532 , n74429 , n74531 );
and ( n74533 , n74426 , n74532 );
or ( n74534 , n74425 , n74533 );
and ( n74535 , n74422 , n74534 );
or ( n74536 , n74421 , n74535 );
and ( n74537 , n74418 , n74536 );
or ( n74538 , n74417 , n74537 );
and ( n74539 , n74414 , n74538 );
or ( n74540 , n74413 , n74539 );
and ( n74541 , n74410 , n74540 );
or ( n74542 , n74409 , n74541 );
and ( n74543 , n74406 , n74542 );
or ( n74544 , n74405 , n74543 );
and ( n74545 , n74402 , n74544 );
or ( n74546 , n74401 , n74545 );
and ( n74547 , n74398 , n74546 );
or ( n74548 , n74397 , n74547 );
and ( n74549 , n74394 , n74548 );
or ( n74550 , n74393 , n74549 );
and ( n74551 , n74390 , n74550 );
or ( n74552 , n74389 , n74551 );
and ( n74553 , n74386 , n74552 );
or ( n74554 , n74385 , n74553 );
and ( n74555 , n74382 , n74554 );
or ( n74556 , n74381 , n74555 );
and ( n74557 , n74378 , n74556 );
or ( n74558 , n74377 , n74557 );
xor ( n74559 , n74374 , n74558 );
buf ( n74560 , n17914 );
and ( n74561 , n30259 , n74560 );
xor ( n74562 , n74559 , n74561 );
xor ( n74563 , n74378 , n74556 );
and ( n74564 , n30264 , n74560 );
and ( n74565 , n74563 , n74564 );
xor ( n74566 , n74563 , n74564 );
xor ( n74567 , n74382 , n74554 );
and ( n74568 , n30269 , n74560 );
and ( n74569 , n74567 , n74568 );
xor ( n74570 , n74567 , n74568 );
xor ( n74571 , n74386 , n74552 );
and ( n74572 , n30274 , n74560 );
and ( n74573 , n74571 , n74572 );
xor ( n74574 , n74571 , n74572 );
xor ( n74575 , n74390 , n74550 );
and ( n74576 , n30279 , n74560 );
and ( n74577 , n74575 , n74576 );
xor ( n74578 , n74575 , n74576 );
xor ( n74579 , n74394 , n74548 );
and ( n74580 , n30284 , n74560 );
and ( n74581 , n74579 , n74580 );
xor ( n74582 , n74579 , n74580 );
xor ( n74583 , n74398 , n74546 );
and ( n74584 , n30289 , n74560 );
and ( n74585 , n74583 , n74584 );
xor ( n74586 , n74583 , n74584 );
xor ( n74587 , n74402 , n74544 );
and ( n74588 , n30294 , n74560 );
and ( n74589 , n74587 , n74588 );
xor ( n74590 , n74587 , n74588 );
xor ( n74591 , n74406 , n74542 );
and ( n74592 , n30299 , n74560 );
and ( n74593 , n74591 , n74592 );
xor ( n74594 , n74591 , n74592 );
xor ( n74595 , n74410 , n74540 );
and ( n74596 , n30304 , n74560 );
and ( n74597 , n74595 , n74596 );
xor ( n74598 , n74595 , n74596 );
xor ( n74599 , n74414 , n74538 );
and ( n74600 , n30309 , n74560 );
and ( n74601 , n74599 , n74600 );
xor ( n74602 , n74599 , n74600 );
xor ( n74603 , n74418 , n74536 );
and ( n74604 , n30314 , n74560 );
and ( n74605 , n74603 , n74604 );
xor ( n74606 , n74603 , n74604 );
xor ( n74607 , n74422 , n74534 );
and ( n74608 , n30319 , n74560 );
and ( n74609 , n74607 , n74608 );
xor ( n74610 , n74607 , n74608 );
xor ( n74611 , n74426 , n74532 );
and ( n74612 , n30324 , n74560 );
and ( n74613 , n74611 , n74612 );
xor ( n74614 , n74611 , n74612 );
xor ( n74615 , n74430 , n74530 );
and ( n74616 , n30329 , n74560 );
and ( n74617 , n74615 , n74616 );
xor ( n74618 , n74615 , n74616 );
xor ( n74619 , n74434 , n74528 );
and ( n74620 , n30334 , n74560 );
and ( n74621 , n74619 , n74620 );
xor ( n74622 , n74619 , n74620 );
xor ( n74623 , n74438 , n74526 );
and ( n74624 , n30339 , n74560 );
and ( n74625 , n74623 , n74624 );
xor ( n74626 , n74623 , n74624 );
xor ( n74627 , n74442 , n74524 );
and ( n74628 , n30344 , n74560 );
and ( n74629 , n74627 , n74628 );
xor ( n74630 , n74627 , n74628 );
xor ( n74631 , n74446 , n74522 );
and ( n74632 , n30349 , n74560 );
and ( n74633 , n74631 , n74632 );
xor ( n74634 , n74631 , n74632 );
xor ( n74635 , n74450 , n74520 );
and ( n74636 , n30354 , n74560 );
and ( n74637 , n74635 , n74636 );
xor ( n74638 , n74635 , n74636 );
xor ( n74639 , n74454 , n74518 );
and ( n74640 , n30359 , n74560 );
and ( n74641 , n74639 , n74640 );
xor ( n74642 , n74639 , n74640 );
xor ( n74643 , n74458 , n74516 );
and ( n74644 , n30364 , n74560 );
and ( n74645 , n74643 , n74644 );
xor ( n74646 , n74643 , n74644 );
xor ( n74647 , n74462 , n74514 );
and ( n74648 , n30369 , n74560 );
and ( n74649 , n74647 , n74648 );
xor ( n74650 , n74647 , n74648 );
xor ( n74651 , n74466 , n74512 );
and ( n74652 , n30374 , n74560 );
and ( n74653 , n74651 , n74652 );
xor ( n74654 , n74651 , n74652 );
xor ( n74655 , n74470 , n74510 );
and ( n74656 , n30379 , n74560 );
and ( n74657 , n74655 , n74656 );
xor ( n74658 , n74655 , n74656 );
xor ( n74659 , n74474 , n74508 );
and ( n74660 , n30384 , n74560 );
and ( n74661 , n74659 , n74660 );
xor ( n74662 , n74659 , n74660 );
xor ( n74663 , n74478 , n74506 );
and ( n74664 , n30389 , n74560 );
and ( n74665 , n74663 , n74664 );
xor ( n74666 , n74663 , n74664 );
xor ( n74667 , n74482 , n74504 );
and ( n74668 , n30394 , n74560 );
and ( n74669 , n74667 , n74668 );
xor ( n74670 , n74667 , n74668 );
xor ( n74671 , n74486 , n74502 );
and ( n74672 , n30399 , n74560 );
and ( n74673 , n74671 , n74672 );
xor ( n74674 , n74671 , n74672 );
xor ( n74675 , n74490 , n74500 );
and ( n74676 , n30404 , n74560 );
and ( n74677 , n74675 , n74676 );
xor ( n74678 , n74675 , n74676 );
xor ( n74679 , n74494 , n74498 );
and ( n74680 , n30409 , n74560 );
and ( n74681 , n74679 , n74680 );
buf ( n74682 , n74681 );
and ( n74683 , n74678 , n74682 );
or ( n74684 , n74677 , n74683 );
and ( n74685 , n74674 , n74684 );
or ( n74686 , n74673 , n74685 );
and ( n74687 , n74670 , n74686 );
or ( n74688 , n74669 , n74687 );
and ( n74689 , n74666 , n74688 );
or ( n74690 , n74665 , n74689 );
and ( n74691 , n74662 , n74690 );
or ( n74692 , n74661 , n74691 );
and ( n74693 , n74658 , n74692 );
or ( n74694 , n74657 , n74693 );
and ( n74695 , n74654 , n74694 );
or ( n74696 , n74653 , n74695 );
and ( n74697 , n74650 , n74696 );
or ( n74698 , n74649 , n74697 );
and ( n74699 , n74646 , n74698 );
or ( n74700 , n74645 , n74699 );
and ( n74701 , n74642 , n74700 );
or ( n74702 , n74641 , n74701 );
and ( n74703 , n74638 , n74702 );
or ( n74704 , n74637 , n74703 );
and ( n74705 , n74634 , n74704 );
or ( n74706 , n74633 , n74705 );
and ( n74707 , n74630 , n74706 );
or ( n74708 , n74629 , n74707 );
and ( n74709 , n74626 , n74708 );
or ( n74710 , n74625 , n74709 );
and ( n74711 , n74622 , n74710 );
or ( n74712 , n74621 , n74711 );
and ( n74713 , n74618 , n74712 );
or ( n74714 , n74617 , n74713 );
and ( n74715 , n74614 , n74714 );
or ( n74716 , n74613 , n74715 );
and ( n74717 , n74610 , n74716 );
or ( n74718 , n74609 , n74717 );
and ( n74719 , n74606 , n74718 );
or ( n74720 , n74605 , n74719 );
and ( n74721 , n74602 , n74720 );
or ( n74722 , n74601 , n74721 );
and ( n74723 , n74598 , n74722 );
or ( n74724 , n74597 , n74723 );
and ( n74725 , n74594 , n74724 );
or ( n74726 , n74593 , n74725 );
and ( n74727 , n74590 , n74726 );
or ( n74728 , n74589 , n74727 );
and ( n74729 , n74586 , n74728 );
or ( n74730 , n74585 , n74729 );
and ( n74731 , n74582 , n74730 );
or ( n74732 , n74581 , n74731 );
and ( n74733 , n74578 , n74732 );
or ( n74734 , n74577 , n74733 );
and ( n74735 , n74574 , n74734 );
or ( n74736 , n74573 , n74735 );
and ( n74737 , n74570 , n74736 );
or ( n74738 , n74569 , n74737 );
and ( n74739 , n74566 , n74738 );
or ( n74740 , n74565 , n74739 );
xor ( n74741 , n74562 , n74740 );
buf ( n74742 , n17912 );
and ( n74743 , n30264 , n74742 );
xor ( n74744 , n74741 , n74743 );
xor ( n74745 , n74566 , n74738 );
and ( n74746 , n30269 , n74742 );
and ( n74747 , n74745 , n74746 );
xor ( n74748 , n74745 , n74746 );
xor ( n74749 , n74570 , n74736 );
and ( n74750 , n30274 , n74742 );
and ( n74751 , n74749 , n74750 );
xor ( n74752 , n74749 , n74750 );
xor ( n74753 , n74574 , n74734 );
and ( n74754 , n30279 , n74742 );
and ( n74755 , n74753 , n74754 );
xor ( n74756 , n74753 , n74754 );
xor ( n74757 , n74578 , n74732 );
and ( n74758 , n30284 , n74742 );
and ( n74759 , n74757 , n74758 );
xor ( n74760 , n74757 , n74758 );
xor ( n74761 , n74582 , n74730 );
and ( n74762 , n30289 , n74742 );
and ( n74763 , n74761 , n74762 );
xor ( n74764 , n74761 , n74762 );
xor ( n74765 , n74586 , n74728 );
and ( n74766 , n30294 , n74742 );
and ( n74767 , n74765 , n74766 );
xor ( n74768 , n74765 , n74766 );
xor ( n74769 , n74590 , n74726 );
and ( n74770 , n30299 , n74742 );
and ( n74771 , n74769 , n74770 );
xor ( n74772 , n74769 , n74770 );
xor ( n74773 , n74594 , n74724 );
and ( n74774 , n30304 , n74742 );
and ( n74775 , n74773 , n74774 );
xor ( n74776 , n74773 , n74774 );
xor ( n74777 , n74598 , n74722 );
and ( n74778 , n30309 , n74742 );
and ( n74779 , n74777 , n74778 );
xor ( n74780 , n74777 , n74778 );
xor ( n74781 , n74602 , n74720 );
and ( n74782 , n30314 , n74742 );
and ( n74783 , n74781 , n74782 );
xor ( n74784 , n74781 , n74782 );
xor ( n74785 , n74606 , n74718 );
and ( n74786 , n30319 , n74742 );
and ( n74787 , n74785 , n74786 );
xor ( n74788 , n74785 , n74786 );
xor ( n74789 , n74610 , n74716 );
and ( n74790 , n30324 , n74742 );
and ( n74791 , n74789 , n74790 );
xor ( n74792 , n74789 , n74790 );
xor ( n74793 , n74614 , n74714 );
and ( n74794 , n30329 , n74742 );
and ( n74795 , n74793 , n74794 );
xor ( n74796 , n74793 , n74794 );
xor ( n74797 , n74618 , n74712 );
and ( n74798 , n30334 , n74742 );
and ( n74799 , n74797 , n74798 );
xor ( n74800 , n74797 , n74798 );
xor ( n74801 , n74622 , n74710 );
and ( n74802 , n30339 , n74742 );
and ( n74803 , n74801 , n74802 );
xor ( n74804 , n74801 , n74802 );
xor ( n74805 , n74626 , n74708 );
and ( n74806 , n30344 , n74742 );
and ( n74807 , n74805 , n74806 );
xor ( n74808 , n74805 , n74806 );
xor ( n74809 , n74630 , n74706 );
and ( n74810 , n30349 , n74742 );
and ( n74811 , n74809 , n74810 );
xor ( n74812 , n74809 , n74810 );
xor ( n74813 , n74634 , n74704 );
and ( n74814 , n30354 , n74742 );
and ( n74815 , n74813 , n74814 );
xor ( n74816 , n74813 , n74814 );
xor ( n74817 , n74638 , n74702 );
and ( n74818 , n30359 , n74742 );
and ( n74819 , n74817 , n74818 );
xor ( n74820 , n74817 , n74818 );
xor ( n74821 , n74642 , n74700 );
and ( n74822 , n30364 , n74742 );
and ( n74823 , n74821 , n74822 );
xor ( n74824 , n74821 , n74822 );
xor ( n74825 , n74646 , n74698 );
and ( n74826 , n30369 , n74742 );
and ( n74827 , n74825 , n74826 );
xor ( n74828 , n74825 , n74826 );
xor ( n74829 , n74650 , n74696 );
and ( n74830 , n30374 , n74742 );
and ( n74831 , n74829 , n74830 );
xor ( n74832 , n74829 , n74830 );
xor ( n74833 , n74654 , n74694 );
and ( n74834 , n30379 , n74742 );
and ( n74835 , n74833 , n74834 );
xor ( n74836 , n74833 , n74834 );
xor ( n74837 , n74658 , n74692 );
and ( n74838 , n30384 , n74742 );
and ( n74839 , n74837 , n74838 );
xor ( n74840 , n74837 , n74838 );
xor ( n74841 , n74662 , n74690 );
and ( n74842 , n30389 , n74742 );
and ( n74843 , n74841 , n74842 );
xor ( n74844 , n74841 , n74842 );
xor ( n74845 , n74666 , n74688 );
and ( n74846 , n30394 , n74742 );
and ( n74847 , n74845 , n74846 );
xor ( n74848 , n74845 , n74846 );
xor ( n74849 , n74670 , n74686 );
and ( n74850 , n30399 , n74742 );
and ( n74851 , n74849 , n74850 );
xor ( n74852 , n74849 , n74850 );
xor ( n74853 , n74674 , n74684 );
and ( n74854 , n30404 , n74742 );
and ( n74855 , n74853 , n74854 );
xor ( n74856 , n74853 , n74854 );
xor ( n74857 , n74678 , n74682 );
and ( n74858 , n30409 , n74742 );
and ( n74859 , n74857 , n74858 );
buf ( n74860 , n74859 );
and ( n74861 , n74856 , n74860 );
or ( n74862 , n74855 , n74861 );
and ( n74863 , n74852 , n74862 );
or ( n74864 , n74851 , n74863 );
and ( n74865 , n74848 , n74864 );
or ( n74866 , n74847 , n74865 );
and ( n74867 , n74844 , n74866 );
or ( n74868 , n74843 , n74867 );
and ( n74869 , n74840 , n74868 );
or ( n74870 , n74839 , n74869 );
and ( n74871 , n74836 , n74870 );
or ( n74872 , n74835 , n74871 );
and ( n74873 , n74832 , n74872 );
or ( n74874 , n74831 , n74873 );
and ( n74875 , n74828 , n74874 );
or ( n74876 , n74827 , n74875 );
and ( n74877 , n74824 , n74876 );
or ( n74878 , n74823 , n74877 );
and ( n74879 , n74820 , n74878 );
or ( n74880 , n74819 , n74879 );
and ( n74881 , n74816 , n74880 );
or ( n74882 , n74815 , n74881 );
and ( n74883 , n74812 , n74882 );
or ( n74884 , n74811 , n74883 );
and ( n74885 , n74808 , n74884 );
or ( n74886 , n74807 , n74885 );
and ( n74887 , n74804 , n74886 );
or ( n74888 , n74803 , n74887 );
and ( n74889 , n74800 , n74888 );
or ( n74890 , n74799 , n74889 );
and ( n74891 , n74796 , n74890 );
or ( n74892 , n74795 , n74891 );
and ( n74893 , n74792 , n74892 );
or ( n74894 , n74791 , n74893 );
and ( n74895 , n74788 , n74894 );
or ( n74896 , n74787 , n74895 );
and ( n74897 , n74784 , n74896 );
or ( n74898 , n74783 , n74897 );
and ( n74899 , n74780 , n74898 );
or ( n74900 , n74779 , n74899 );
and ( n74901 , n74776 , n74900 );
or ( n74902 , n74775 , n74901 );
and ( n74903 , n74772 , n74902 );
or ( n74904 , n74771 , n74903 );
and ( n74905 , n74768 , n74904 );
or ( n74906 , n74767 , n74905 );
and ( n74907 , n74764 , n74906 );
or ( n74908 , n74763 , n74907 );
and ( n74909 , n74760 , n74908 );
or ( n74910 , n74759 , n74909 );
and ( n74911 , n74756 , n74910 );
or ( n74912 , n74755 , n74911 );
and ( n74913 , n74752 , n74912 );
or ( n74914 , n74751 , n74913 );
and ( n74915 , n74748 , n74914 );
or ( n74916 , n74747 , n74915 );
xor ( n74917 , n74744 , n74916 );
buf ( n74918 , n17910 );
and ( n74919 , n30269 , n74918 );
xor ( n74920 , n74917 , n74919 );
xor ( n74921 , n74748 , n74914 );
and ( n74922 , n30274 , n74918 );
and ( n74923 , n74921 , n74922 );
xor ( n74924 , n74921 , n74922 );
xor ( n74925 , n74752 , n74912 );
and ( n74926 , n30279 , n74918 );
and ( n74927 , n74925 , n74926 );
xor ( n74928 , n74925 , n74926 );
xor ( n74929 , n74756 , n74910 );
and ( n74930 , n30284 , n74918 );
and ( n74931 , n74929 , n74930 );
xor ( n74932 , n74929 , n74930 );
xor ( n74933 , n74760 , n74908 );
and ( n74934 , n30289 , n74918 );
and ( n74935 , n74933 , n74934 );
xor ( n74936 , n74933 , n74934 );
xor ( n74937 , n74764 , n74906 );
and ( n74938 , n30294 , n74918 );
and ( n74939 , n74937 , n74938 );
xor ( n74940 , n74937 , n74938 );
xor ( n74941 , n74768 , n74904 );
and ( n74942 , n30299 , n74918 );
and ( n74943 , n74941 , n74942 );
xor ( n74944 , n74941 , n74942 );
xor ( n74945 , n74772 , n74902 );
and ( n74946 , n30304 , n74918 );
and ( n74947 , n74945 , n74946 );
xor ( n74948 , n74945 , n74946 );
xor ( n74949 , n74776 , n74900 );
and ( n74950 , n30309 , n74918 );
and ( n74951 , n74949 , n74950 );
xor ( n74952 , n74949 , n74950 );
xor ( n74953 , n74780 , n74898 );
and ( n74954 , n30314 , n74918 );
and ( n74955 , n74953 , n74954 );
xor ( n74956 , n74953 , n74954 );
xor ( n74957 , n74784 , n74896 );
and ( n74958 , n30319 , n74918 );
and ( n74959 , n74957 , n74958 );
xor ( n74960 , n74957 , n74958 );
xor ( n74961 , n74788 , n74894 );
and ( n74962 , n30324 , n74918 );
and ( n74963 , n74961 , n74962 );
xor ( n74964 , n74961 , n74962 );
xor ( n74965 , n74792 , n74892 );
and ( n74966 , n30329 , n74918 );
and ( n74967 , n74965 , n74966 );
xor ( n74968 , n74965 , n74966 );
xor ( n74969 , n74796 , n74890 );
and ( n74970 , n30334 , n74918 );
and ( n74971 , n74969 , n74970 );
xor ( n74972 , n74969 , n74970 );
xor ( n74973 , n74800 , n74888 );
and ( n74974 , n30339 , n74918 );
and ( n74975 , n74973 , n74974 );
xor ( n74976 , n74973 , n74974 );
xor ( n74977 , n74804 , n74886 );
and ( n74978 , n30344 , n74918 );
and ( n74979 , n74977 , n74978 );
xor ( n74980 , n74977 , n74978 );
xor ( n74981 , n74808 , n74884 );
and ( n74982 , n30349 , n74918 );
and ( n74983 , n74981 , n74982 );
xor ( n74984 , n74981 , n74982 );
xor ( n74985 , n74812 , n74882 );
and ( n74986 , n30354 , n74918 );
and ( n74987 , n74985 , n74986 );
xor ( n74988 , n74985 , n74986 );
xor ( n74989 , n74816 , n74880 );
and ( n74990 , n30359 , n74918 );
and ( n74991 , n74989 , n74990 );
xor ( n74992 , n74989 , n74990 );
xor ( n74993 , n74820 , n74878 );
and ( n74994 , n30364 , n74918 );
and ( n74995 , n74993 , n74994 );
xor ( n74996 , n74993 , n74994 );
xor ( n74997 , n74824 , n74876 );
and ( n74998 , n30369 , n74918 );
and ( n74999 , n74997 , n74998 );
xor ( n75000 , n74997 , n74998 );
xor ( n75001 , n74828 , n74874 );
and ( n75002 , n30374 , n74918 );
and ( n75003 , n75001 , n75002 );
xor ( n75004 , n75001 , n75002 );
xor ( n75005 , n74832 , n74872 );
and ( n75006 , n30379 , n74918 );
and ( n75007 , n75005 , n75006 );
xor ( n75008 , n75005 , n75006 );
xor ( n75009 , n74836 , n74870 );
and ( n75010 , n30384 , n74918 );
and ( n75011 , n75009 , n75010 );
xor ( n75012 , n75009 , n75010 );
xor ( n75013 , n74840 , n74868 );
and ( n75014 , n30389 , n74918 );
and ( n75015 , n75013 , n75014 );
xor ( n75016 , n75013 , n75014 );
xor ( n75017 , n74844 , n74866 );
and ( n75018 , n30394 , n74918 );
and ( n75019 , n75017 , n75018 );
xor ( n75020 , n75017 , n75018 );
xor ( n75021 , n74848 , n74864 );
and ( n75022 , n30399 , n74918 );
and ( n75023 , n75021 , n75022 );
xor ( n75024 , n75021 , n75022 );
xor ( n75025 , n74852 , n74862 );
and ( n75026 , n30404 , n74918 );
and ( n75027 , n75025 , n75026 );
xor ( n75028 , n75025 , n75026 );
xor ( n75029 , n74856 , n74860 );
and ( n75030 , n30409 , n74918 );
and ( n75031 , n75029 , n75030 );
buf ( n75032 , n75031 );
and ( n75033 , n75028 , n75032 );
or ( n75034 , n75027 , n75033 );
and ( n75035 , n75024 , n75034 );
or ( n75036 , n75023 , n75035 );
and ( n75037 , n75020 , n75036 );
or ( n75038 , n75019 , n75037 );
and ( n75039 , n75016 , n75038 );
or ( n75040 , n75015 , n75039 );
and ( n75041 , n75012 , n75040 );
or ( n75042 , n75011 , n75041 );
and ( n75043 , n75008 , n75042 );
or ( n75044 , n75007 , n75043 );
and ( n75045 , n75004 , n75044 );
or ( n75046 , n75003 , n75045 );
and ( n75047 , n75000 , n75046 );
or ( n75048 , n74999 , n75047 );
and ( n75049 , n74996 , n75048 );
or ( n75050 , n74995 , n75049 );
and ( n75051 , n74992 , n75050 );
or ( n75052 , n74991 , n75051 );
and ( n75053 , n74988 , n75052 );
or ( n75054 , n74987 , n75053 );
and ( n75055 , n74984 , n75054 );
or ( n75056 , n74983 , n75055 );
and ( n75057 , n74980 , n75056 );
or ( n75058 , n74979 , n75057 );
and ( n75059 , n74976 , n75058 );
or ( n75060 , n74975 , n75059 );
and ( n75061 , n74972 , n75060 );
or ( n75062 , n74971 , n75061 );
and ( n75063 , n74968 , n75062 );
or ( n75064 , n74967 , n75063 );
and ( n75065 , n74964 , n75064 );
or ( n75066 , n74963 , n75065 );
and ( n75067 , n74960 , n75066 );
or ( n75068 , n74959 , n75067 );
and ( n75069 , n74956 , n75068 );
or ( n75070 , n74955 , n75069 );
and ( n75071 , n74952 , n75070 );
or ( n75072 , n74951 , n75071 );
and ( n75073 , n74948 , n75072 );
or ( n75074 , n74947 , n75073 );
and ( n75075 , n74944 , n75074 );
or ( n75076 , n74943 , n75075 );
and ( n75077 , n74940 , n75076 );
or ( n75078 , n74939 , n75077 );
and ( n75079 , n74936 , n75078 );
or ( n75080 , n74935 , n75079 );
and ( n75081 , n74932 , n75080 );
or ( n75082 , n74931 , n75081 );
and ( n75083 , n74928 , n75082 );
or ( n75084 , n74927 , n75083 );
and ( n75085 , n74924 , n75084 );
or ( n75086 , n74923 , n75085 );
xor ( n75087 , n74920 , n75086 );
buf ( n75088 , n17908 );
and ( n75089 , n30274 , n75088 );
xor ( n75090 , n75087 , n75089 );
xor ( n75091 , n74924 , n75084 );
and ( n75092 , n30279 , n75088 );
and ( n75093 , n75091 , n75092 );
xor ( n75094 , n75091 , n75092 );
xor ( n75095 , n74928 , n75082 );
and ( n75096 , n30284 , n75088 );
and ( n75097 , n75095 , n75096 );
xor ( n75098 , n75095 , n75096 );
xor ( n75099 , n74932 , n75080 );
and ( n75100 , n30289 , n75088 );
and ( n75101 , n75099 , n75100 );
xor ( n75102 , n75099 , n75100 );
xor ( n75103 , n74936 , n75078 );
and ( n75104 , n30294 , n75088 );
and ( n75105 , n75103 , n75104 );
xor ( n75106 , n75103 , n75104 );
xor ( n75107 , n74940 , n75076 );
and ( n75108 , n30299 , n75088 );
and ( n75109 , n75107 , n75108 );
xor ( n75110 , n75107 , n75108 );
xor ( n75111 , n74944 , n75074 );
and ( n75112 , n30304 , n75088 );
and ( n75113 , n75111 , n75112 );
xor ( n75114 , n75111 , n75112 );
xor ( n75115 , n74948 , n75072 );
and ( n75116 , n30309 , n75088 );
and ( n75117 , n75115 , n75116 );
xor ( n75118 , n75115 , n75116 );
xor ( n75119 , n74952 , n75070 );
and ( n75120 , n30314 , n75088 );
and ( n75121 , n75119 , n75120 );
xor ( n75122 , n75119 , n75120 );
xor ( n75123 , n74956 , n75068 );
and ( n75124 , n30319 , n75088 );
and ( n75125 , n75123 , n75124 );
xor ( n75126 , n75123 , n75124 );
xor ( n75127 , n74960 , n75066 );
and ( n75128 , n30324 , n75088 );
and ( n75129 , n75127 , n75128 );
xor ( n75130 , n75127 , n75128 );
xor ( n75131 , n74964 , n75064 );
and ( n75132 , n30329 , n75088 );
and ( n75133 , n75131 , n75132 );
xor ( n75134 , n75131 , n75132 );
xor ( n75135 , n74968 , n75062 );
and ( n75136 , n30334 , n75088 );
and ( n75137 , n75135 , n75136 );
xor ( n75138 , n75135 , n75136 );
xor ( n75139 , n74972 , n75060 );
and ( n75140 , n30339 , n75088 );
and ( n75141 , n75139 , n75140 );
xor ( n75142 , n75139 , n75140 );
xor ( n75143 , n74976 , n75058 );
and ( n75144 , n30344 , n75088 );
and ( n75145 , n75143 , n75144 );
xor ( n75146 , n75143 , n75144 );
xor ( n75147 , n74980 , n75056 );
and ( n75148 , n30349 , n75088 );
and ( n75149 , n75147 , n75148 );
xor ( n75150 , n75147 , n75148 );
xor ( n75151 , n74984 , n75054 );
and ( n75152 , n30354 , n75088 );
and ( n75153 , n75151 , n75152 );
xor ( n75154 , n75151 , n75152 );
xor ( n75155 , n74988 , n75052 );
and ( n75156 , n30359 , n75088 );
and ( n75157 , n75155 , n75156 );
xor ( n75158 , n75155 , n75156 );
xor ( n75159 , n74992 , n75050 );
and ( n75160 , n30364 , n75088 );
and ( n75161 , n75159 , n75160 );
xor ( n75162 , n75159 , n75160 );
xor ( n75163 , n74996 , n75048 );
and ( n75164 , n30369 , n75088 );
and ( n75165 , n75163 , n75164 );
xor ( n75166 , n75163 , n75164 );
xor ( n75167 , n75000 , n75046 );
and ( n75168 , n30374 , n75088 );
and ( n75169 , n75167 , n75168 );
xor ( n75170 , n75167 , n75168 );
xor ( n75171 , n75004 , n75044 );
and ( n75172 , n30379 , n75088 );
and ( n75173 , n75171 , n75172 );
xor ( n75174 , n75171 , n75172 );
xor ( n75175 , n75008 , n75042 );
and ( n75176 , n30384 , n75088 );
and ( n75177 , n75175 , n75176 );
xor ( n75178 , n75175 , n75176 );
xor ( n75179 , n75012 , n75040 );
and ( n75180 , n30389 , n75088 );
and ( n75181 , n75179 , n75180 );
xor ( n75182 , n75179 , n75180 );
xor ( n75183 , n75016 , n75038 );
and ( n75184 , n30394 , n75088 );
and ( n75185 , n75183 , n75184 );
xor ( n75186 , n75183 , n75184 );
xor ( n75187 , n75020 , n75036 );
and ( n75188 , n30399 , n75088 );
and ( n75189 , n75187 , n75188 );
xor ( n75190 , n75187 , n75188 );
xor ( n75191 , n75024 , n75034 );
and ( n75192 , n30404 , n75088 );
and ( n75193 , n75191 , n75192 );
xor ( n75194 , n75191 , n75192 );
xor ( n75195 , n75028 , n75032 );
and ( n75196 , n30409 , n75088 );
and ( n75197 , n75195 , n75196 );
buf ( n75198 , n75197 );
and ( n75199 , n75194 , n75198 );
or ( n75200 , n75193 , n75199 );
and ( n75201 , n75190 , n75200 );
or ( n75202 , n75189 , n75201 );
and ( n75203 , n75186 , n75202 );
or ( n75204 , n75185 , n75203 );
and ( n75205 , n75182 , n75204 );
or ( n75206 , n75181 , n75205 );
and ( n75207 , n75178 , n75206 );
or ( n75208 , n75177 , n75207 );
and ( n75209 , n75174 , n75208 );
or ( n75210 , n75173 , n75209 );
and ( n75211 , n75170 , n75210 );
or ( n75212 , n75169 , n75211 );
and ( n75213 , n75166 , n75212 );
or ( n75214 , n75165 , n75213 );
and ( n75215 , n75162 , n75214 );
or ( n75216 , n75161 , n75215 );
and ( n75217 , n75158 , n75216 );
or ( n75218 , n75157 , n75217 );
and ( n75219 , n75154 , n75218 );
or ( n75220 , n75153 , n75219 );
and ( n75221 , n75150 , n75220 );
or ( n75222 , n75149 , n75221 );
and ( n75223 , n75146 , n75222 );
or ( n75224 , n75145 , n75223 );
and ( n75225 , n75142 , n75224 );
or ( n75226 , n75141 , n75225 );
and ( n75227 , n75138 , n75226 );
or ( n75228 , n75137 , n75227 );
and ( n75229 , n75134 , n75228 );
or ( n75230 , n75133 , n75229 );
and ( n75231 , n75130 , n75230 );
or ( n75232 , n75129 , n75231 );
and ( n75233 , n75126 , n75232 );
or ( n75234 , n75125 , n75233 );
and ( n75235 , n75122 , n75234 );
or ( n75236 , n75121 , n75235 );
and ( n75237 , n75118 , n75236 );
or ( n75238 , n75117 , n75237 );
and ( n75239 , n75114 , n75238 );
or ( n75240 , n75113 , n75239 );
and ( n75241 , n75110 , n75240 );
or ( n75242 , n75109 , n75241 );
and ( n75243 , n75106 , n75242 );
or ( n75244 , n75105 , n75243 );
and ( n75245 , n75102 , n75244 );
or ( n75246 , n75101 , n75245 );
and ( n75247 , n75098 , n75246 );
or ( n75248 , n75097 , n75247 );
and ( n75249 , n75094 , n75248 );
or ( n75250 , n75093 , n75249 );
xor ( n75251 , n75090 , n75250 );
buf ( n75252 , n17906 );
and ( n75253 , n30279 , n75252 );
xor ( n75254 , n75251 , n75253 );
xor ( n75255 , n75094 , n75248 );
and ( n75256 , n30284 , n75252 );
and ( n75257 , n75255 , n75256 );
xor ( n75258 , n75255 , n75256 );
xor ( n75259 , n75098 , n75246 );
and ( n75260 , n30289 , n75252 );
and ( n75261 , n75259 , n75260 );
xor ( n75262 , n75259 , n75260 );
xor ( n75263 , n75102 , n75244 );
and ( n75264 , n30294 , n75252 );
and ( n75265 , n75263 , n75264 );
xor ( n75266 , n75263 , n75264 );
xor ( n75267 , n75106 , n75242 );
and ( n75268 , n30299 , n75252 );
and ( n75269 , n75267 , n75268 );
xor ( n75270 , n75267 , n75268 );
xor ( n75271 , n75110 , n75240 );
and ( n75272 , n30304 , n75252 );
and ( n75273 , n75271 , n75272 );
xor ( n75274 , n75271 , n75272 );
xor ( n75275 , n75114 , n75238 );
and ( n75276 , n30309 , n75252 );
and ( n75277 , n75275 , n75276 );
xor ( n75278 , n75275 , n75276 );
xor ( n75279 , n75118 , n75236 );
and ( n75280 , n30314 , n75252 );
and ( n75281 , n75279 , n75280 );
xor ( n75282 , n75279 , n75280 );
xor ( n75283 , n75122 , n75234 );
and ( n75284 , n30319 , n75252 );
and ( n75285 , n75283 , n75284 );
xor ( n75286 , n75283 , n75284 );
xor ( n75287 , n75126 , n75232 );
and ( n75288 , n30324 , n75252 );
and ( n75289 , n75287 , n75288 );
xor ( n75290 , n75287 , n75288 );
xor ( n75291 , n75130 , n75230 );
and ( n75292 , n30329 , n75252 );
and ( n75293 , n75291 , n75292 );
xor ( n75294 , n75291 , n75292 );
xor ( n75295 , n75134 , n75228 );
and ( n75296 , n30334 , n75252 );
and ( n75297 , n75295 , n75296 );
xor ( n75298 , n75295 , n75296 );
xor ( n75299 , n75138 , n75226 );
and ( n75300 , n30339 , n75252 );
and ( n75301 , n75299 , n75300 );
xor ( n75302 , n75299 , n75300 );
xor ( n75303 , n75142 , n75224 );
and ( n75304 , n30344 , n75252 );
and ( n75305 , n75303 , n75304 );
xor ( n75306 , n75303 , n75304 );
xor ( n75307 , n75146 , n75222 );
and ( n75308 , n30349 , n75252 );
and ( n75309 , n75307 , n75308 );
xor ( n75310 , n75307 , n75308 );
xor ( n75311 , n75150 , n75220 );
and ( n75312 , n30354 , n75252 );
and ( n75313 , n75311 , n75312 );
xor ( n75314 , n75311 , n75312 );
xor ( n75315 , n75154 , n75218 );
and ( n75316 , n30359 , n75252 );
and ( n75317 , n75315 , n75316 );
xor ( n75318 , n75315 , n75316 );
xor ( n75319 , n75158 , n75216 );
and ( n75320 , n30364 , n75252 );
and ( n75321 , n75319 , n75320 );
xor ( n75322 , n75319 , n75320 );
xor ( n75323 , n75162 , n75214 );
and ( n75324 , n30369 , n75252 );
and ( n75325 , n75323 , n75324 );
xor ( n75326 , n75323 , n75324 );
xor ( n75327 , n75166 , n75212 );
and ( n75328 , n30374 , n75252 );
and ( n75329 , n75327 , n75328 );
xor ( n75330 , n75327 , n75328 );
xor ( n75331 , n75170 , n75210 );
and ( n75332 , n30379 , n75252 );
and ( n75333 , n75331 , n75332 );
xor ( n75334 , n75331 , n75332 );
xor ( n75335 , n75174 , n75208 );
and ( n75336 , n30384 , n75252 );
and ( n75337 , n75335 , n75336 );
xor ( n75338 , n75335 , n75336 );
xor ( n75339 , n75178 , n75206 );
and ( n75340 , n30389 , n75252 );
and ( n75341 , n75339 , n75340 );
xor ( n75342 , n75339 , n75340 );
xor ( n75343 , n75182 , n75204 );
and ( n75344 , n30394 , n75252 );
and ( n75345 , n75343 , n75344 );
xor ( n75346 , n75343 , n75344 );
xor ( n75347 , n75186 , n75202 );
and ( n75348 , n30399 , n75252 );
and ( n75349 , n75347 , n75348 );
xor ( n75350 , n75347 , n75348 );
xor ( n75351 , n75190 , n75200 );
and ( n75352 , n30404 , n75252 );
and ( n75353 , n75351 , n75352 );
xor ( n75354 , n75351 , n75352 );
xor ( n75355 , n75194 , n75198 );
and ( n75356 , n30409 , n75252 );
and ( n75357 , n75355 , n75356 );
buf ( n75358 , n75357 );
and ( n75359 , n75354 , n75358 );
or ( n75360 , n75353 , n75359 );
and ( n75361 , n75350 , n75360 );
or ( n75362 , n75349 , n75361 );
and ( n75363 , n75346 , n75362 );
or ( n75364 , n75345 , n75363 );
and ( n75365 , n75342 , n75364 );
or ( n75366 , n75341 , n75365 );
and ( n75367 , n75338 , n75366 );
or ( n75368 , n75337 , n75367 );
and ( n75369 , n75334 , n75368 );
or ( n75370 , n75333 , n75369 );
and ( n75371 , n75330 , n75370 );
or ( n75372 , n75329 , n75371 );
and ( n75373 , n75326 , n75372 );
or ( n75374 , n75325 , n75373 );
and ( n75375 , n75322 , n75374 );
or ( n75376 , n75321 , n75375 );
and ( n75377 , n75318 , n75376 );
or ( n75378 , n75317 , n75377 );
and ( n75379 , n75314 , n75378 );
or ( n75380 , n75313 , n75379 );
and ( n75381 , n75310 , n75380 );
or ( n75382 , n75309 , n75381 );
and ( n75383 , n75306 , n75382 );
or ( n75384 , n75305 , n75383 );
and ( n75385 , n75302 , n75384 );
or ( n75386 , n75301 , n75385 );
and ( n75387 , n75298 , n75386 );
or ( n75388 , n75297 , n75387 );
and ( n75389 , n75294 , n75388 );
or ( n75390 , n75293 , n75389 );
and ( n75391 , n75290 , n75390 );
or ( n75392 , n75289 , n75391 );
and ( n75393 , n75286 , n75392 );
or ( n75394 , n75285 , n75393 );
and ( n75395 , n75282 , n75394 );
or ( n75396 , n75281 , n75395 );
and ( n75397 , n75278 , n75396 );
or ( n75398 , n75277 , n75397 );
and ( n75399 , n75274 , n75398 );
or ( n75400 , n75273 , n75399 );
and ( n75401 , n75270 , n75400 );
or ( n75402 , n75269 , n75401 );
and ( n75403 , n75266 , n75402 );
or ( n75404 , n75265 , n75403 );
and ( n75405 , n75262 , n75404 );
or ( n75406 , n75261 , n75405 );
and ( n75407 , n75258 , n75406 );
or ( n75408 , n75257 , n75407 );
xor ( n75409 , n75254 , n75408 );
buf ( n75410 , n17904 );
and ( n75411 , n30284 , n75410 );
xor ( n75412 , n75409 , n75411 );
xor ( n75413 , n75258 , n75406 );
and ( n75414 , n30289 , n75410 );
and ( n75415 , n75413 , n75414 );
xor ( n75416 , n75413 , n75414 );
xor ( n75417 , n75262 , n75404 );
and ( n75418 , n30294 , n75410 );
and ( n75419 , n75417 , n75418 );
xor ( n75420 , n75417 , n75418 );
xor ( n75421 , n75266 , n75402 );
and ( n75422 , n30299 , n75410 );
and ( n75423 , n75421 , n75422 );
xor ( n75424 , n75421 , n75422 );
xor ( n75425 , n75270 , n75400 );
and ( n75426 , n30304 , n75410 );
and ( n75427 , n75425 , n75426 );
xor ( n75428 , n75425 , n75426 );
xor ( n75429 , n75274 , n75398 );
and ( n75430 , n30309 , n75410 );
and ( n75431 , n75429 , n75430 );
xor ( n75432 , n75429 , n75430 );
xor ( n75433 , n75278 , n75396 );
and ( n75434 , n30314 , n75410 );
and ( n75435 , n75433 , n75434 );
xor ( n75436 , n75433 , n75434 );
xor ( n75437 , n75282 , n75394 );
and ( n75438 , n30319 , n75410 );
and ( n75439 , n75437 , n75438 );
xor ( n75440 , n75437 , n75438 );
xor ( n75441 , n75286 , n75392 );
and ( n75442 , n30324 , n75410 );
and ( n75443 , n75441 , n75442 );
xor ( n75444 , n75441 , n75442 );
xor ( n75445 , n75290 , n75390 );
and ( n75446 , n30329 , n75410 );
and ( n75447 , n75445 , n75446 );
xor ( n75448 , n75445 , n75446 );
xor ( n75449 , n75294 , n75388 );
and ( n75450 , n30334 , n75410 );
and ( n75451 , n75449 , n75450 );
xor ( n75452 , n75449 , n75450 );
xor ( n75453 , n75298 , n75386 );
and ( n75454 , n30339 , n75410 );
and ( n75455 , n75453 , n75454 );
xor ( n75456 , n75453 , n75454 );
xor ( n75457 , n75302 , n75384 );
and ( n75458 , n30344 , n75410 );
and ( n75459 , n75457 , n75458 );
xor ( n75460 , n75457 , n75458 );
xor ( n75461 , n75306 , n75382 );
and ( n75462 , n30349 , n75410 );
and ( n75463 , n75461 , n75462 );
xor ( n75464 , n75461 , n75462 );
xor ( n75465 , n75310 , n75380 );
and ( n75466 , n30354 , n75410 );
and ( n75467 , n75465 , n75466 );
xor ( n75468 , n75465 , n75466 );
xor ( n75469 , n75314 , n75378 );
and ( n75470 , n30359 , n75410 );
and ( n75471 , n75469 , n75470 );
xor ( n75472 , n75469 , n75470 );
xor ( n75473 , n75318 , n75376 );
and ( n75474 , n30364 , n75410 );
and ( n75475 , n75473 , n75474 );
xor ( n75476 , n75473 , n75474 );
xor ( n75477 , n75322 , n75374 );
and ( n75478 , n30369 , n75410 );
and ( n75479 , n75477 , n75478 );
xor ( n75480 , n75477 , n75478 );
xor ( n75481 , n75326 , n75372 );
and ( n75482 , n30374 , n75410 );
and ( n75483 , n75481 , n75482 );
xor ( n75484 , n75481 , n75482 );
xor ( n75485 , n75330 , n75370 );
and ( n75486 , n30379 , n75410 );
and ( n75487 , n75485 , n75486 );
xor ( n75488 , n75485 , n75486 );
xor ( n75489 , n75334 , n75368 );
and ( n75490 , n30384 , n75410 );
and ( n75491 , n75489 , n75490 );
xor ( n75492 , n75489 , n75490 );
xor ( n75493 , n75338 , n75366 );
and ( n75494 , n30389 , n75410 );
and ( n75495 , n75493 , n75494 );
xor ( n75496 , n75493 , n75494 );
xor ( n75497 , n75342 , n75364 );
and ( n75498 , n30394 , n75410 );
and ( n75499 , n75497 , n75498 );
xor ( n75500 , n75497 , n75498 );
xor ( n75501 , n75346 , n75362 );
and ( n75502 , n30399 , n75410 );
and ( n75503 , n75501 , n75502 );
xor ( n75504 , n75501 , n75502 );
xor ( n75505 , n75350 , n75360 );
and ( n75506 , n30404 , n75410 );
and ( n75507 , n75505 , n75506 );
xor ( n75508 , n75505 , n75506 );
xor ( n75509 , n75354 , n75358 );
and ( n75510 , n30409 , n75410 );
and ( n75511 , n75509 , n75510 );
buf ( n75512 , n75511 );
and ( n75513 , n75508 , n75512 );
or ( n75514 , n75507 , n75513 );
and ( n75515 , n75504 , n75514 );
or ( n75516 , n75503 , n75515 );
and ( n75517 , n75500 , n75516 );
or ( n75518 , n75499 , n75517 );
and ( n75519 , n75496 , n75518 );
or ( n75520 , n75495 , n75519 );
and ( n75521 , n75492 , n75520 );
or ( n75522 , n75491 , n75521 );
and ( n75523 , n75488 , n75522 );
or ( n75524 , n75487 , n75523 );
and ( n75525 , n75484 , n75524 );
or ( n75526 , n75483 , n75525 );
and ( n75527 , n75480 , n75526 );
or ( n75528 , n75479 , n75527 );
and ( n75529 , n75476 , n75528 );
or ( n75530 , n75475 , n75529 );
and ( n75531 , n75472 , n75530 );
or ( n75532 , n75471 , n75531 );
and ( n75533 , n75468 , n75532 );
or ( n75534 , n75467 , n75533 );
and ( n75535 , n75464 , n75534 );
or ( n75536 , n75463 , n75535 );
and ( n75537 , n75460 , n75536 );
or ( n75538 , n75459 , n75537 );
and ( n75539 , n75456 , n75538 );
or ( n75540 , n75455 , n75539 );
and ( n75541 , n75452 , n75540 );
or ( n75542 , n75451 , n75541 );
and ( n75543 , n75448 , n75542 );
or ( n75544 , n75447 , n75543 );
and ( n75545 , n75444 , n75544 );
or ( n75546 , n75443 , n75545 );
and ( n75547 , n75440 , n75546 );
or ( n75548 , n75439 , n75547 );
and ( n75549 , n75436 , n75548 );
or ( n75550 , n75435 , n75549 );
and ( n75551 , n75432 , n75550 );
or ( n75552 , n75431 , n75551 );
and ( n75553 , n75428 , n75552 );
or ( n75554 , n75427 , n75553 );
and ( n75555 , n75424 , n75554 );
or ( n75556 , n75423 , n75555 );
and ( n75557 , n75420 , n75556 );
or ( n75558 , n75419 , n75557 );
and ( n75559 , n75416 , n75558 );
or ( n75560 , n75415 , n75559 );
xor ( n75561 , n75412 , n75560 );
buf ( n75562 , n17902 );
and ( n75563 , n30289 , n75562 );
xor ( n75564 , n75561 , n75563 );
xor ( n75565 , n75416 , n75558 );
and ( n75566 , n30294 , n75562 );
and ( n75567 , n75565 , n75566 );
xor ( n75568 , n75565 , n75566 );
xor ( n75569 , n75420 , n75556 );
and ( n75570 , n30299 , n75562 );
and ( n75571 , n75569 , n75570 );
xor ( n75572 , n75569 , n75570 );
xor ( n75573 , n75424 , n75554 );
and ( n75574 , n30304 , n75562 );
and ( n75575 , n75573 , n75574 );
xor ( n75576 , n75573 , n75574 );
xor ( n75577 , n75428 , n75552 );
and ( n75578 , n30309 , n75562 );
and ( n75579 , n75577 , n75578 );
xor ( n75580 , n75577 , n75578 );
xor ( n75581 , n75432 , n75550 );
and ( n75582 , n30314 , n75562 );
and ( n75583 , n75581 , n75582 );
xor ( n75584 , n75581 , n75582 );
xor ( n75585 , n75436 , n75548 );
and ( n75586 , n30319 , n75562 );
and ( n75587 , n75585 , n75586 );
xor ( n75588 , n75585 , n75586 );
xor ( n75589 , n75440 , n75546 );
and ( n75590 , n30324 , n75562 );
and ( n75591 , n75589 , n75590 );
xor ( n75592 , n75589 , n75590 );
xor ( n75593 , n75444 , n75544 );
and ( n75594 , n30329 , n75562 );
and ( n75595 , n75593 , n75594 );
xor ( n75596 , n75593 , n75594 );
xor ( n75597 , n75448 , n75542 );
and ( n75598 , n30334 , n75562 );
and ( n75599 , n75597 , n75598 );
xor ( n75600 , n75597 , n75598 );
xor ( n75601 , n75452 , n75540 );
and ( n75602 , n30339 , n75562 );
and ( n75603 , n75601 , n75602 );
xor ( n75604 , n75601 , n75602 );
xor ( n75605 , n75456 , n75538 );
and ( n75606 , n30344 , n75562 );
and ( n75607 , n75605 , n75606 );
xor ( n75608 , n75605 , n75606 );
xor ( n75609 , n75460 , n75536 );
and ( n75610 , n30349 , n75562 );
and ( n75611 , n75609 , n75610 );
xor ( n75612 , n75609 , n75610 );
xor ( n75613 , n75464 , n75534 );
and ( n75614 , n30354 , n75562 );
and ( n75615 , n75613 , n75614 );
xor ( n75616 , n75613 , n75614 );
xor ( n75617 , n75468 , n75532 );
and ( n75618 , n30359 , n75562 );
and ( n75619 , n75617 , n75618 );
xor ( n75620 , n75617 , n75618 );
xor ( n75621 , n75472 , n75530 );
and ( n75622 , n30364 , n75562 );
and ( n75623 , n75621 , n75622 );
xor ( n75624 , n75621 , n75622 );
xor ( n75625 , n75476 , n75528 );
and ( n75626 , n30369 , n75562 );
and ( n75627 , n75625 , n75626 );
xor ( n75628 , n75625 , n75626 );
xor ( n75629 , n75480 , n75526 );
and ( n75630 , n30374 , n75562 );
and ( n75631 , n75629 , n75630 );
xor ( n75632 , n75629 , n75630 );
xor ( n75633 , n75484 , n75524 );
and ( n75634 , n30379 , n75562 );
and ( n75635 , n75633 , n75634 );
xor ( n75636 , n75633 , n75634 );
xor ( n75637 , n75488 , n75522 );
and ( n75638 , n30384 , n75562 );
and ( n75639 , n75637 , n75638 );
xor ( n75640 , n75637 , n75638 );
xor ( n75641 , n75492 , n75520 );
and ( n75642 , n30389 , n75562 );
and ( n75643 , n75641 , n75642 );
xor ( n75644 , n75641 , n75642 );
xor ( n75645 , n75496 , n75518 );
and ( n75646 , n30394 , n75562 );
and ( n75647 , n75645 , n75646 );
xor ( n75648 , n75645 , n75646 );
xor ( n75649 , n75500 , n75516 );
and ( n75650 , n30399 , n75562 );
and ( n75651 , n75649 , n75650 );
xor ( n75652 , n75649 , n75650 );
xor ( n75653 , n75504 , n75514 );
and ( n75654 , n30404 , n75562 );
and ( n75655 , n75653 , n75654 );
xor ( n75656 , n75653 , n75654 );
xor ( n75657 , n75508 , n75512 );
and ( n75658 , n30409 , n75562 );
and ( n75659 , n75657 , n75658 );
buf ( n75660 , n75659 );
and ( n75661 , n75656 , n75660 );
or ( n75662 , n75655 , n75661 );
and ( n75663 , n75652 , n75662 );
or ( n75664 , n75651 , n75663 );
and ( n75665 , n75648 , n75664 );
or ( n75666 , n75647 , n75665 );
and ( n75667 , n75644 , n75666 );
or ( n75668 , n75643 , n75667 );
and ( n75669 , n75640 , n75668 );
or ( n75670 , n75639 , n75669 );
and ( n75671 , n75636 , n75670 );
or ( n75672 , n75635 , n75671 );
and ( n75673 , n75632 , n75672 );
or ( n75674 , n75631 , n75673 );
and ( n75675 , n75628 , n75674 );
or ( n75676 , n75627 , n75675 );
and ( n75677 , n75624 , n75676 );
or ( n75678 , n75623 , n75677 );
and ( n75679 , n75620 , n75678 );
or ( n75680 , n75619 , n75679 );
and ( n75681 , n75616 , n75680 );
or ( n75682 , n75615 , n75681 );
and ( n75683 , n75612 , n75682 );
or ( n75684 , n75611 , n75683 );
and ( n75685 , n75608 , n75684 );
or ( n75686 , n75607 , n75685 );
and ( n75687 , n75604 , n75686 );
or ( n75688 , n75603 , n75687 );
and ( n75689 , n75600 , n75688 );
or ( n75690 , n75599 , n75689 );
and ( n75691 , n75596 , n75690 );
or ( n75692 , n75595 , n75691 );
and ( n75693 , n75592 , n75692 );
or ( n75694 , n75591 , n75693 );
and ( n75695 , n75588 , n75694 );
or ( n75696 , n75587 , n75695 );
and ( n75697 , n75584 , n75696 );
or ( n75698 , n75583 , n75697 );
and ( n75699 , n75580 , n75698 );
or ( n75700 , n75579 , n75699 );
and ( n75701 , n75576 , n75700 );
or ( n75702 , n75575 , n75701 );
and ( n75703 , n75572 , n75702 );
or ( n75704 , n75571 , n75703 );
and ( n75705 , n75568 , n75704 );
or ( n75706 , n75567 , n75705 );
xor ( n75707 , n75564 , n75706 );
buf ( n75708 , n17900 );
and ( n75709 , n30294 , n75708 );
xor ( n75710 , n75707 , n75709 );
xor ( n75711 , n75568 , n75704 );
and ( n75712 , n30299 , n75708 );
and ( n75713 , n75711 , n75712 );
xor ( n75714 , n75711 , n75712 );
xor ( n75715 , n75572 , n75702 );
and ( n75716 , n30304 , n75708 );
and ( n75717 , n75715 , n75716 );
xor ( n75718 , n75715 , n75716 );
xor ( n75719 , n75576 , n75700 );
and ( n75720 , n30309 , n75708 );
and ( n75721 , n75719 , n75720 );
xor ( n75722 , n75719 , n75720 );
xor ( n75723 , n75580 , n75698 );
and ( n75724 , n30314 , n75708 );
and ( n75725 , n75723 , n75724 );
xor ( n75726 , n75723 , n75724 );
xor ( n75727 , n75584 , n75696 );
and ( n75728 , n30319 , n75708 );
and ( n75729 , n75727 , n75728 );
xor ( n75730 , n75727 , n75728 );
xor ( n75731 , n75588 , n75694 );
and ( n75732 , n30324 , n75708 );
and ( n75733 , n75731 , n75732 );
xor ( n75734 , n75731 , n75732 );
xor ( n75735 , n75592 , n75692 );
and ( n75736 , n30329 , n75708 );
and ( n75737 , n75735 , n75736 );
xor ( n75738 , n75735 , n75736 );
xor ( n75739 , n75596 , n75690 );
and ( n75740 , n30334 , n75708 );
and ( n75741 , n75739 , n75740 );
xor ( n75742 , n75739 , n75740 );
xor ( n75743 , n75600 , n75688 );
and ( n75744 , n30339 , n75708 );
and ( n75745 , n75743 , n75744 );
xor ( n75746 , n75743 , n75744 );
xor ( n75747 , n75604 , n75686 );
and ( n75748 , n30344 , n75708 );
and ( n75749 , n75747 , n75748 );
xor ( n75750 , n75747 , n75748 );
xor ( n75751 , n75608 , n75684 );
and ( n75752 , n30349 , n75708 );
and ( n75753 , n75751 , n75752 );
xor ( n75754 , n75751 , n75752 );
xor ( n75755 , n75612 , n75682 );
and ( n75756 , n30354 , n75708 );
and ( n75757 , n75755 , n75756 );
xor ( n75758 , n75755 , n75756 );
xor ( n75759 , n75616 , n75680 );
and ( n75760 , n30359 , n75708 );
and ( n75761 , n75759 , n75760 );
xor ( n75762 , n75759 , n75760 );
xor ( n75763 , n75620 , n75678 );
and ( n75764 , n30364 , n75708 );
and ( n75765 , n75763 , n75764 );
xor ( n75766 , n75763 , n75764 );
xor ( n75767 , n75624 , n75676 );
and ( n75768 , n30369 , n75708 );
and ( n75769 , n75767 , n75768 );
xor ( n75770 , n75767 , n75768 );
xor ( n75771 , n75628 , n75674 );
and ( n75772 , n30374 , n75708 );
and ( n75773 , n75771 , n75772 );
xor ( n75774 , n75771 , n75772 );
xor ( n75775 , n75632 , n75672 );
and ( n75776 , n30379 , n75708 );
and ( n75777 , n75775 , n75776 );
xor ( n75778 , n75775 , n75776 );
xor ( n75779 , n75636 , n75670 );
and ( n75780 , n30384 , n75708 );
and ( n75781 , n75779 , n75780 );
xor ( n75782 , n75779 , n75780 );
xor ( n75783 , n75640 , n75668 );
and ( n75784 , n30389 , n75708 );
and ( n75785 , n75783 , n75784 );
xor ( n75786 , n75783 , n75784 );
xor ( n75787 , n75644 , n75666 );
and ( n75788 , n30394 , n75708 );
and ( n75789 , n75787 , n75788 );
xor ( n75790 , n75787 , n75788 );
xor ( n75791 , n75648 , n75664 );
and ( n75792 , n30399 , n75708 );
and ( n75793 , n75791 , n75792 );
xor ( n75794 , n75791 , n75792 );
xor ( n75795 , n75652 , n75662 );
and ( n75796 , n30404 , n75708 );
and ( n75797 , n75795 , n75796 );
xor ( n75798 , n75795 , n75796 );
xor ( n75799 , n75656 , n75660 );
and ( n75800 , n30409 , n75708 );
and ( n75801 , n75799 , n75800 );
buf ( n75802 , n75801 );
and ( n75803 , n75798 , n75802 );
or ( n75804 , n75797 , n75803 );
and ( n75805 , n75794 , n75804 );
or ( n75806 , n75793 , n75805 );
and ( n75807 , n75790 , n75806 );
or ( n75808 , n75789 , n75807 );
and ( n75809 , n75786 , n75808 );
or ( n75810 , n75785 , n75809 );
and ( n75811 , n75782 , n75810 );
or ( n75812 , n75781 , n75811 );
and ( n75813 , n75778 , n75812 );
or ( n75814 , n75777 , n75813 );
and ( n75815 , n75774 , n75814 );
or ( n75816 , n75773 , n75815 );
and ( n75817 , n75770 , n75816 );
or ( n75818 , n75769 , n75817 );
and ( n75819 , n75766 , n75818 );
or ( n75820 , n75765 , n75819 );
and ( n75821 , n75762 , n75820 );
or ( n75822 , n75761 , n75821 );
and ( n75823 , n75758 , n75822 );
or ( n75824 , n75757 , n75823 );
and ( n75825 , n75754 , n75824 );
or ( n75826 , n75753 , n75825 );
and ( n75827 , n75750 , n75826 );
or ( n75828 , n75749 , n75827 );
and ( n75829 , n75746 , n75828 );
or ( n75830 , n75745 , n75829 );
and ( n75831 , n75742 , n75830 );
or ( n75832 , n75741 , n75831 );
and ( n75833 , n75738 , n75832 );
or ( n75834 , n75737 , n75833 );
and ( n75835 , n75734 , n75834 );
or ( n75836 , n75733 , n75835 );
and ( n75837 , n75730 , n75836 );
or ( n75838 , n75729 , n75837 );
and ( n75839 , n75726 , n75838 );
or ( n75840 , n75725 , n75839 );
and ( n75841 , n75722 , n75840 );
or ( n75842 , n75721 , n75841 );
and ( n75843 , n75718 , n75842 );
or ( n75844 , n75717 , n75843 );
and ( n75845 , n75714 , n75844 );
or ( n75846 , n75713 , n75845 );
xor ( n75847 , n75710 , n75846 );
buf ( n75848 , n17898 );
and ( n75849 , n30299 , n75848 );
xor ( n75850 , n75847 , n75849 );
xor ( n75851 , n75714 , n75844 );
and ( n75852 , n30304 , n75848 );
and ( n75853 , n75851 , n75852 );
xor ( n75854 , n75851 , n75852 );
xor ( n75855 , n75718 , n75842 );
and ( n75856 , n30309 , n75848 );
and ( n75857 , n75855 , n75856 );
xor ( n75858 , n75855 , n75856 );
xor ( n75859 , n75722 , n75840 );
and ( n75860 , n30314 , n75848 );
and ( n75861 , n75859 , n75860 );
xor ( n75862 , n75859 , n75860 );
xor ( n75863 , n75726 , n75838 );
and ( n75864 , n30319 , n75848 );
and ( n75865 , n75863 , n75864 );
xor ( n75866 , n75863 , n75864 );
xor ( n75867 , n75730 , n75836 );
and ( n75868 , n30324 , n75848 );
and ( n75869 , n75867 , n75868 );
xor ( n75870 , n75867 , n75868 );
xor ( n75871 , n75734 , n75834 );
and ( n75872 , n30329 , n75848 );
and ( n75873 , n75871 , n75872 );
xor ( n75874 , n75871 , n75872 );
xor ( n75875 , n75738 , n75832 );
and ( n75876 , n30334 , n75848 );
and ( n75877 , n75875 , n75876 );
xor ( n75878 , n75875 , n75876 );
xor ( n75879 , n75742 , n75830 );
and ( n75880 , n30339 , n75848 );
and ( n75881 , n75879 , n75880 );
xor ( n75882 , n75879 , n75880 );
xor ( n75883 , n75746 , n75828 );
and ( n75884 , n30344 , n75848 );
and ( n75885 , n75883 , n75884 );
xor ( n75886 , n75883 , n75884 );
xor ( n75887 , n75750 , n75826 );
and ( n75888 , n30349 , n75848 );
and ( n75889 , n75887 , n75888 );
xor ( n75890 , n75887 , n75888 );
xor ( n75891 , n75754 , n75824 );
and ( n75892 , n30354 , n75848 );
and ( n75893 , n75891 , n75892 );
xor ( n75894 , n75891 , n75892 );
xor ( n75895 , n75758 , n75822 );
and ( n75896 , n30359 , n75848 );
and ( n75897 , n75895 , n75896 );
xor ( n75898 , n75895 , n75896 );
xor ( n75899 , n75762 , n75820 );
and ( n75900 , n30364 , n75848 );
and ( n75901 , n75899 , n75900 );
xor ( n75902 , n75899 , n75900 );
xor ( n75903 , n75766 , n75818 );
and ( n75904 , n30369 , n75848 );
and ( n75905 , n75903 , n75904 );
xor ( n75906 , n75903 , n75904 );
xor ( n75907 , n75770 , n75816 );
and ( n75908 , n30374 , n75848 );
and ( n75909 , n75907 , n75908 );
xor ( n75910 , n75907 , n75908 );
xor ( n75911 , n75774 , n75814 );
and ( n75912 , n30379 , n75848 );
and ( n75913 , n75911 , n75912 );
xor ( n75914 , n75911 , n75912 );
xor ( n75915 , n75778 , n75812 );
and ( n75916 , n30384 , n75848 );
and ( n75917 , n75915 , n75916 );
xor ( n75918 , n75915 , n75916 );
xor ( n75919 , n75782 , n75810 );
and ( n75920 , n30389 , n75848 );
and ( n75921 , n75919 , n75920 );
xor ( n75922 , n75919 , n75920 );
xor ( n75923 , n75786 , n75808 );
and ( n75924 , n30394 , n75848 );
and ( n75925 , n75923 , n75924 );
xor ( n75926 , n75923 , n75924 );
xor ( n75927 , n75790 , n75806 );
and ( n75928 , n30399 , n75848 );
and ( n75929 , n75927 , n75928 );
xor ( n75930 , n75927 , n75928 );
xor ( n75931 , n75794 , n75804 );
and ( n75932 , n30404 , n75848 );
and ( n75933 , n75931 , n75932 );
xor ( n75934 , n75931 , n75932 );
xor ( n75935 , n75798 , n75802 );
and ( n75936 , n30409 , n75848 );
and ( n75937 , n75935 , n75936 );
buf ( n75938 , n75937 );
and ( n75939 , n75934 , n75938 );
or ( n75940 , n75933 , n75939 );
and ( n75941 , n75930 , n75940 );
or ( n75942 , n75929 , n75941 );
and ( n75943 , n75926 , n75942 );
or ( n75944 , n75925 , n75943 );
and ( n75945 , n75922 , n75944 );
or ( n75946 , n75921 , n75945 );
and ( n75947 , n75918 , n75946 );
or ( n75948 , n75917 , n75947 );
and ( n75949 , n75914 , n75948 );
or ( n75950 , n75913 , n75949 );
and ( n75951 , n75910 , n75950 );
or ( n75952 , n75909 , n75951 );
and ( n75953 , n75906 , n75952 );
or ( n75954 , n75905 , n75953 );
and ( n75955 , n75902 , n75954 );
or ( n75956 , n75901 , n75955 );
and ( n75957 , n75898 , n75956 );
or ( n75958 , n75897 , n75957 );
and ( n75959 , n75894 , n75958 );
or ( n75960 , n75893 , n75959 );
and ( n75961 , n75890 , n75960 );
or ( n75962 , n75889 , n75961 );
and ( n75963 , n75886 , n75962 );
or ( n75964 , n75885 , n75963 );
and ( n75965 , n75882 , n75964 );
or ( n75966 , n75881 , n75965 );
and ( n75967 , n75878 , n75966 );
or ( n75968 , n75877 , n75967 );
and ( n75969 , n75874 , n75968 );
or ( n75970 , n75873 , n75969 );
and ( n75971 , n75870 , n75970 );
or ( n75972 , n75869 , n75971 );
and ( n75973 , n75866 , n75972 );
or ( n75974 , n75865 , n75973 );
and ( n75975 , n75862 , n75974 );
or ( n75976 , n75861 , n75975 );
and ( n75977 , n75858 , n75976 );
or ( n75978 , n75857 , n75977 );
and ( n75979 , n75854 , n75978 );
or ( n75980 , n75853 , n75979 );
xor ( n75981 , n75850 , n75980 );
buf ( n75982 , n17896 );
and ( n75983 , n30304 , n75982 );
xor ( n75984 , n75981 , n75983 );
xor ( n75985 , n75854 , n75978 );
and ( n75986 , n30309 , n75982 );
and ( n75987 , n75985 , n75986 );
xor ( n75988 , n75985 , n75986 );
xor ( n75989 , n75858 , n75976 );
and ( n75990 , n30314 , n75982 );
and ( n75991 , n75989 , n75990 );
xor ( n75992 , n75989 , n75990 );
xor ( n75993 , n75862 , n75974 );
and ( n75994 , n30319 , n75982 );
and ( n75995 , n75993 , n75994 );
xor ( n75996 , n75993 , n75994 );
xor ( n75997 , n75866 , n75972 );
and ( n75998 , n30324 , n75982 );
and ( n75999 , n75997 , n75998 );
xor ( n76000 , n75997 , n75998 );
xor ( n76001 , n75870 , n75970 );
and ( n76002 , n30329 , n75982 );
and ( n76003 , n76001 , n76002 );
xor ( n76004 , n76001 , n76002 );
xor ( n76005 , n75874 , n75968 );
and ( n76006 , n30334 , n75982 );
and ( n76007 , n76005 , n76006 );
xor ( n76008 , n76005 , n76006 );
xor ( n76009 , n75878 , n75966 );
and ( n76010 , n30339 , n75982 );
and ( n76011 , n76009 , n76010 );
xor ( n76012 , n76009 , n76010 );
xor ( n76013 , n75882 , n75964 );
and ( n76014 , n30344 , n75982 );
and ( n76015 , n76013 , n76014 );
xor ( n76016 , n76013 , n76014 );
xor ( n76017 , n75886 , n75962 );
and ( n76018 , n30349 , n75982 );
and ( n76019 , n76017 , n76018 );
xor ( n76020 , n76017 , n76018 );
xor ( n76021 , n75890 , n75960 );
and ( n76022 , n30354 , n75982 );
and ( n76023 , n76021 , n76022 );
xor ( n76024 , n76021 , n76022 );
xor ( n76025 , n75894 , n75958 );
and ( n76026 , n30359 , n75982 );
and ( n76027 , n76025 , n76026 );
xor ( n76028 , n76025 , n76026 );
xor ( n76029 , n75898 , n75956 );
and ( n76030 , n30364 , n75982 );
and ( n76031 , n76029 , n76030 );
xor ( n76032 , n76029 , n76030 );
xor ( n76033 , n75902 , n75954 );
and ( n76034 , n30369 , n75982 );
and ( n76035 , n76033 , n76034 );
xor ( n76036 , n76033 , n76034 );
xor ( n76037 , n75906 , n75952 );
and ( n76038 , n30374 , n75982 );
and ( n76039 , n76037 , n76038 );
xor ( n76040 , n76037 , n76038 );
xor ( n76041 , n75910 , n75950 );
and ( n76042 , n30379 , n75982 );
and ( n76043 , n76041 , n76042 );
xor ( n76044 , n76041 , n76042 );
xor ( n76045 , n75914 , n75948 );
and ( n76046 , n30384 , n75982 );
and ( n76047 , n76045 , n76046 );
xor ( n76048 , n76045 , n76046 );
xor ( n76049 , n75918 , n75946 );
and ( n76050 , n30389 , n75982 );
and ( n76051 , n76049 , n76050 );
xor ( n76052 , n76049 , n76050 );
xor ( n76053 , n75922 , n75944 );
and ( n76054 , n30394 , n75982 );
and ( n76055 , n76053 , n76054 );
xor ( n76056 , n76053 , n76054 );
xor ( n76057 , n75926 , n75942 );
and ( n76058 , n30399 , n75982 );
and ( n76059 , n76057 , n76058 );
xor ( n76060 , n76057 , n76058 );
xor ( n76061 , n75930 , n75940 );
and ( n76062 , n30404 , n75982 );
and ( n76063 , n76061 , n76062 );
xor ( n76064 , n76061 , n76062 );
xor ( n76065 , n75934 , n75938 );
and ( n76066 , n30409 , n75982 );
and ( n76067 , n76065 , n76066 );
buf ( n76068 , n76067 );
and ( n76069 , n76064 , n76068 );
or ( n76070 , n76063 , n76069 );
and ( n76071 , n76060 , n76070 );
or ( n76072 , n76059 , n76071 );
and ( n76073 , n76056 , n76072 );
or ( n76074 , n76055 , n76073 );
and ( n76075 , n76052 , n76074 );
or ( n76076 , n76051 , n76075 );
and ( n76077 , n76048 , n76076 );
or ( n76078 , n76047 , n76077 );
and ( n76079 , n76044 , n76078 );
or ( n76080 , n76043 , n76079 );
and ( n76081 , n76040 , n76080 );
or ( n76082 , n76039 , n76081 );
and ( n76083 , n76036 , n76082 );
or ( n76084 , n76035 , n76083 );
and ( n76085 , n76032 , n76084 );
or ( n76086 , n76031 , n76085 );
and ( n76087 , n76028 , n76086 );
or ( n76088 , n76027 , n76087 );
and ( n76089 , n76024 , n76088 );
or ( n76090 , n76023 , n76089 );
and ( n76091 , n76020 , n76090 );
or ( n76092 , n76019 , n76091 );
and ( n76093 , n76016 , n76092 );
or ( n76094 , n76015 , n76093 );
and ( n76095 , n76012 , n76094 );
or ( n76096 , n76011 , n76095 );
and ( n76097 , n76008 , n76096 );
or ( n76098 , n76007 , n76097 );
and ( n76099 , n76004 , n76098 );
or ( n76100 , n76003 , n76099 );
and ( n76101 , n76000 , n76100 );
or ( n76102 , n75999 , n76101 );
and ( n76103 , n75996 , n76102 );
or ( n76104 , n75995 , n76103 );
and ( n76105 , n75992 , n76104 );
or ( n76106 , n75991 , n76105 );
and ( n76107 , n75988 , n76106 );
or ( n76108 , n75987 , n76107 );
xor ( n76109 , n75984 , n76108 );
buf ( n76110 , n17894 );
and ( n76111 , n30309 , n76110 );
xor ( n76112 , n76109 , n76111 );
xor ( n76113 , n75988 , n76106 );
and ( n76114 , n30314 , n76110 );
and ( n76115 , n76113 , n76114 );
xor ( n76116 , n76113 , n76114 );
xor ( n76117 , n75992 , n76104 );
and ( n76118 , n30319 , n76110 );
and ( n76119 , n76117 , n76118 );
xor ( n76120 , n76117 , n76118 );
xor ( n76121 , n75996 , n76102 );
and ( n76122 , n30324 , n76110 );
and ( n76123 , n76121 , n76122 );
xor ( n76124 , n76121 , n76122 );
xor ( n76125 , n76000 , n76100 );
and ( n76126 , n30329 , n76110 );
and ( n76127 , n76125 , n76126 );
xor ( n76128 , n76125 , n76126 );
xor ( n76129 , n76004 , n76098 );
and ( n76130 , n30334 , n76110 );
and ( n76131 , n76129 , n76130 );
xor ( n76132 , n76129 , n76130 );
xor ( n76133 , n76008 , n76096 );
and ( n76134 , n30339 , n76110 );
and ( n76135 , n76133 , n76134 );
xor ( n76136 , n76133 , n76134 );
xor ( n76137 , n76012 , n76094 );
and ( n76138 , n30344 , n76110 );
and ( n76139 , n76137 , n76138 );
xor ( n76140 , n76137 , n76138 );
xor ( n76141 , n76016 , n76092 );
and ( n76142 , n30349 , n76110 );
and ( n76143 , n76141 , n76142 );
xor ( n76144 , n76141 , n76142 );
xor ( n76145 , n76020 , n76090 );
and ( n76146 , n30354 , n76110 );
and ( n76147 , n76145 , n76146 );
xor ( n76148 , n76145 , n76146 );
xor ( n76149 , n76024 , n76088 );
and ( n76150 , n30359 , n76110 );
and ( n76151 , n76149 , n76150 );
xor ( n76152 , n76149 , n76150 );
xor ( n76153 , n76028 , n76086 );
and ( n76154 , n30364 , n76110 );
and ( n76155 , n76153 , n76154 );
xor ( n76156 , n76153 , n76154 );
xor ( n76157 , n76032 , n76084 );
and ( n76158 , n30369 , n76110 );
and ( n76159 , n76157 , n76158 );
xor ( n76160 , n76157 , n76158 );
xor ( n76161 , n76036 , n76082 );
and ( n76162 , n30374 , n76110 );
and ( n76163 , n76161 , n76162 );
xor ( n76164 , n76161 , n76162 );
xor ( n76165 , n76040 , n76080 );
and ( n76166 , n30379 , n76110 );
and ( n76167 , n76165 , n76166 );
xor ( n76168 , n76165 , n76166 );
xor ( n76169 , n76044 , n76078 );
and ( n76170 , n30384 , n76110 );
and ( n76171 , n76169 , n76170 );
xor ( n76172 , n76169 , n76170 );
xor ( n76173 , n76048 , n76076 );
and ( n76174 , n30389 , n76110 );
and ( n76175 , n76173 , n76174 );
xor ( n76176 , n76173 , n76174 );
xor ( n76177 , n76052 , n76074 );
and ( n76178 , n30394 , n76110 );
and ( n76179 , n76177 , n76178 );
xor ( n76180 , n76177 , n76178 );
xor ( n76181 , n76056 , n76072 );
and ( n76182 , n30399 , n76110 );
and ( n76183 , n76181 , n76182 );
xor ( n76184 , n76181 , n76182 );
xor ( n76185 , n76060 , n76070 );
and ( n76186 , n30404 , n76110 );
and ( n76187 , n76185 , n76186 );
xor ( n76188 , n76185 , n76186 );
xor ( n76189 , n76064 , n76068 );
and ( n76190 , n30409 , n76110 );
and ( n76191 , n76189 , n76190 );
buf ( n76192 , n76191 );
and ( n76193 , n76188 , n76192 );
or ( n76194 , n76187 , n76193 );
and ( n76195 , n76184 , n76194 );
or ( n76196 , n76183 , n76195 );
and ( n76197 , n76180 , n76196 );
or ( n76198 , n76179 , n76197 );
and ( n76199 , n76176 , n76198 );
or ( n76200 , n76175 , n76199 );
and ( n76201 , n76172 , n76200 );
or ( n76202 , n76171 , n76201 );
and ( n76203 , n76168 , n76202 );
or ( n76204 , n76167 , n76203 );
and ( n76205 , n76164 , n76204 );
or ( n76206 , n76163 , n76205 );
and ( n76207 , n76160 , n76206 );
or ( n76208 , n76159 , n76207 );
and ( n76209 , n76156 , n76208 );
or ( n76210 , n76155 , n76209 );
and ( n76211 , n76152 , n76210 );
or ( n76212 , n76151 , n76211 );
and ( n76213 , n76148 , n76212 );
or ( n76214 , n76147 , n76213 );
and ( n76215 , n76144 , n76214 );
or ( n76216 , n76143 , n76215 );
and ( n76217 , n76140 , n76216 );
or ( n76218 , n76139 , n76217 );
and ( n76219 , n76136 , n76218 );
or ( n76220 , n76135 , n76219 );
and ( n76221 , n76132 , n76220 );
or ( n76222 , n76131 , n76221 );
and ( n76223 , n76128 , n76222 );
or ( n76224 , n76127 , n76223 );
and ( n76225 , n76124 , n76224 );
or ( n76226 , n76123 , n76225 );
and ( n76227 , n76120 , n76226 );
or ( n76228 , n76119 , n76227 );
and ( n76229 , n76116 , n76228 );
or ( n76230 , n76115 , n76229 );
xor ( n76231 , n76112 , n76230 );
buf ( n76232 , n17892 );
and ( n76233 , n30314 , n76232 );
xor ( n76234 , n76231 , n76233 );
xor ( n76235 , n76116 , n76228 );
and ( n76236 , n30319 , n76232 );
and ( n76237 , n76235 , n76236 );
xor ( n76238 , n76235 , n76236 );
xor ( n76239 , n76120 , n76226 );
and ( n76240 , n30324 , n76232 );
and ( n76241 , n76239 , n76240 );
xor ( n76242 , n76239 , n76240 );
xor ( n76243 , n76124 , n76224 );
and ( n76244 , n30329 , n76232 );
and ( n76245 , n76243 , n76244 );
xor ( n76246 , n76243 , n76244 );
xor ( n76247 , n76128 , n76222 );
and ( n76248 , n30334 , n76232 );
and ( n76249 , n76247 , n76248 );
xor ( n76250 , n76247 , n76248 );
xor ( n76251 , n76132 , n76220 );
and ( n76252 , n30339 , n76232 );
and ( n76253 , n76251 , n76252 );
xor ( n76254 , n76251 , n76252 );
xor ( n76255 , n76136 , n76218 );
and ( n76256 , n30344 , n76232 );
and ( n76257 , n76255 , n76256 );
xor ( n76258 , n76255 , n76256 );
xor ( n76259 , n76140 , n76216 );
and ( n76260 , n30349 , n76232 );
and ( n76261 , n76259 , n76260 );
xor ( n76262 , n76259 , n76260 );
xor ( n76263 , n76144 , n76214 );
and ( n76264 , n30354 , n76232 );
and ( n76265 , n76263 , n76264 );
xor ( n76266 , n76263 , n76264 );
xor ( n76267 , n76148 , n76212 );
and ( n76268 , n30359 , n76232 );
and ( n76269 , n76267 , n76268 );
xor ( n76270 , n76267 , n76268 );
xor ( n76271 , n76152 , n76210 );
and ( n76272 , n30364 , n76232 );
and ( n76273 , n76271 , n76272 );
xor ( n76274 , n76271 , n76272 );
xor ( n76275 , n76156 , n76208 );
and ( n76276 , n30369 , n76232 );
and ( n76277 , n76275 , n76276 );
xor ( n76278 , n76275 , n76276 );
xor ( n76279 , n76160 , n76206 );
and ( n76280 , n30374 , n76232 );
and ( n76281 , n76279 , n76280 );
xor ( n76282 , n76279 , n76280 );
xor ( n76283 , n76164 , n76204 );
and ( n76284 , n30379 , n76232 );
and ( n76285 , n76283 , n76284 );
xor ( n76286 , n76283 , n76284 );
xor ( n76287 , n76168 , n76202 );
and ( n76288 , n30384 , n76232 );
and ( n76289 , n76287 , n76288 );
xor ( n76290 , n76287 , n76288 );
xor ( n76291 , n76172 , n76200 );
and ( n76292 , n30389 , n76232 );
and ( n76293 , n76291 , n76292 );
xor ( n76294 , n76291 , n76292 );
xor ( n76295 , n76176 , n76198 );
and ( n76296 , n30394 , n76232 );
and ( n76297 , n76295 , n76296 );
xor ( n76298 , n76295 , n76296 );
xor ( n76299 , n76180 , n76196 );
and ( n76300 , n30399 , n76232 );
and ( n76301 , n76299 , n76300 );
xor ( n76302 , n76299 , n76300 );
xor ( n76303 , n76184 , n76194 );
and ( n76304 , n30404 , n76232 );
and ( n76305 , n76303 , n76304 );
xor ( n76306 , n76303 , n76304 );
xor ( n76307 , n76188 , n76192 );
and ( n76308 , n30409 , n76232 );
and ( n76309 , n76307 , n76308 );
buf ( n76310 , n76309 );
and ( n76311 , n76306 , n76310 );
or ( n76312 , n76305 , n76311 );
and ( n76313 , n76302 , n76312 );
or ( n76314 , n76301 , n76313 );
and ( n76315 , n76298 , n76314 );
or ( n76316 , n76297 , n76315 );
and ( n76317 , n76294 , n76316 );
or ( n76318 , n76293 , n76317 );
and ( n76319 , n76290 , n76318 );
or ( n76320 , n76289 , n76319 );
and ( n76321 , n76286 , n76320 );
or ( n76322 , n76285 , n76321 );
and ( n76323 , n76282 , n76322 );
or ( n76324 , n76281 , n76323 );
and ( n76325 , n76278 , n76324 );
or ( n76326 , n76277 , n76325 );
and ( n76327 , n76274 , n76326 );
or ( n76328 , n76273 , n76327 );
and ( n76329 , n76270 , n76328 );
or ( n76330 , n76269 , n76329 );
and ( n76331 , n76266 , n76330 );
or ( n76332 , n76265 , n76331 );
and ( n76333 , n76262 , n76332 );
or ( n76334 , n76261 , n76333 );
and ( n76335 , n76258 , n76334 );
or ( n76336 , n76257 , n76335 );
and ( n76337 , n76254 , n76336 );
or ( n76338 , n76253 , n76337 );
and ( n76339 , n76250 , n76338 );
or ( n76340 , n76249 , n76339 );
and ( n76341 , n76246 , n76340 );
or ( n76342 , n76245 , n76341 );
and ( n76343 , n76242 , n76342 );
or ( n76344 , n76241 , n76343 );
and ( n76345 , n76238 , n76344 );
or ( n76346 , n76237 , n76345 );
xor ( n76347 , n76234 , n76346 );
buf ( n76348 , n17890 );
and ( n76349 , n30319 , n76348 );
xor ( n76350 , n76347 , n76349 );
xor ( n76351 , n76238 , n76344 );
and ( n76352 , n30324 , n76348 );
and ( n76353 , n76351 , n76352 );
xor ( n76354 , n76351 , n76352 );
xor ( n76355 , n76242 , n76342 );
and ( n76356 , n30329 , n76348 );
and ( n76357 , n76355 , n76356 );
xor ( n76358 , n76355 , n76356 );
xor ( n76359 , n76246 , n76340 );
and ( n76360 , n30334 , n76348 );
and ( n76361 , n76359 , n76360 );
xor ( n76362 , n76359 , n76360 );
xor ( n76363 , n76250 , n76338 );
and ( n76364 , n30339 , n76348 );
and ( n76365 , n76363 , n76364 );
xor ( n76366 , n76363 , n76364 );
xor ( n76367 , n76254 , n76336 );
and ( n76368 , n30344 , n76348 );
and ( n76369 , n76367 , n76368 );
xor ( n76370 , n76367 , n76368 );
xor ( n76371 , n76258 , n76334 );
and ( n76372 , n30349 , n76348 );
and ( n76373 , n76371 , n76372 );
xor ( n76374 , n76371 , n76372 );
xor ( n76375 , n76262 , n76332 );
and ( n76376 , n30354 , n76348 );
and ( n76377 , n76375 , n76376 );
xor ( n76378 , n76375 , n76376 );
xor ( n76379 , n76266 , n76330 );
and ( n76380 , n30359 , n76348 );
and ( n76381 , n76379 , n76380 );
xor ( n76382 , n76379 , n76380 );
xor ( n76383 , n76270 , n76328 );
and ( n76384 , n30364 , n76348 );
and ( n76385 , n76383 , n76384 );
xor ( n76386 , n76383 , n76384 );
xor ( n76387 , n76274 , n76326 );
and ( n76388 , n30369 , n76348 );
and ( n76389 , n76387 , n76388 );
xor ( n76390 , n76387 , n76388 );
xor ( n76391 , n76278 , n76324 );
and ( n76392 , n30374 , n76348 );
and ( n76393 , n76391 , n76392 );
xor ( n76394 , n76391 , n76392 );
xor ( n76395 , n76282 , n76322 );
and ( n76396 , n30379 , n76348 );
and ( n76397 , n76395 , n76396 );
xor ( n76398 , n76395 , n76396 );
xor ( n76399 , n76286 , n76320 );
and ( n76400 , n30384 , n76348 );
and ( n76401 , n76399 , n76400 );
xor ( n76402 , n76399 , n76400 );
xor ( n76403 , n76290 , n76318 );
and ( n76404 , n30389 , n76348 );
and ( n76405 , n76403 , n76404 );
xor ( n76406 , n76403 , n76404 );
xor ( n76407 , n76294 , n76316 );
and ( n76408 , n30394 , n76348 );
and ( n76409 , n76407 , n76408 );
xor ( n76410 , n76407 , n76408 );
xor ( n76411 , n76298 , n76314 );
and ( n76412 , n30399 , n76348 );
and ( n76413 , n76411 , n76412 );
xor ( n76414 , n76411 , n76412 );
xor ( n76415 , n76302 , n76312 );
and ( n76416 , n30404 , n76348 );
and ( n76417 , n76415 , n76416 );
xor ( n76418 , n76415 , n76416 );
xor ( n76419 , n76306 , n76310 );
and ( n76420 , n30409 , n76348 );
and ( n76421 , n76419 , n76420 );
buf ( n76422 , n76421 );
and ( n76423 , n76418 , n76422 );
or ( n76424 , n76417 , n76423 );
and ( n76425 , n76414 , n76424 );
or ( n76426 , n76413 , n76425 );
and ( n76427 , n76410 , n76426 );
or ( n76428 , n76409 , n76427 );
and ( n76429 , n76406 , n76428 );
or ( n76430 , n76405 , n76429 );
and ( n76431 , n76402 , n76430 );
or ( n76432 , n76401 , n76431 );
and ( n76433 , n76398 , n76432 );
or ( n76434 , n76397 , n76433 );
and ( n76435 , n76394 , n76434 );
or ( n76436 , n76393 , n76435 );
and ( n76437 , n76390 , n76436 );
or ( n76438 , n76389 , n76437 );
and ( n76439 , n76386 , n76438 );
or ( n76440 , n76385 , n76439 );
and ( n76441 , n76382 , n76440 );
or ( n76442 , n76381 , n76441 );
and ( n76443 , n76378 , n76442 );
or ( n76444 , n76377 , n76443 );
and ( n76445 , n76374 , n76444 );
or ( n76446 , n76373 , n76445 );
and ( n76447 , n76370 , n76446 );
or ( n76448 , n76369 , n76447 );
and ( n76449 , n76366 , n76448 );
or ( n76450 , n76365 , n76449 );
and ( n76451 , n76362 , n76450 );
or ( n76452 , n76361 , n76451 );
and ( n76453 , n76358 , n76452 );
or ( n76454 , n76357 , n76453 );
and ( n76455 , n76354 , n76454 );
or ( n76456 , n76353 , n76455 );
xor ( n76457 , n76350 , n76456 );
buf ( n76458 , n17888 );
and ( n76459 , n30324 , n76458 );
xor ( n76460 , n76457 , n76459 );
xor ( n76461 , n76354 , n76454 );
and ( n76462 , n30329 , n76458 );
and ( n76463 , n76461 , n76462 );
xor ( n76464 , n76461 , n76462 );
xor ( n76465 , n76358 , n76452 );
and ( n76466 , n30334 , n76458 );
and ( n76467 , n76465 , n76466 );
xor ( n76468 , n76465 , n76466 );
xor ( n76469 , n76362 , n76450 );
and ( n76470 , n30339 , n76458 );
and ( n76471 , n76469 , n76470 );
xor ( n76472 , n76469 , n76470 );
xor ( n76473 , n76366 , n76448 );
and ( n76474 , n30344 , n76458 );
and ( n76475 , n76473 , n76474 );
xor ( n76476 , n76473 , n76474 );
xor ( n76477 , n76370 , n76446 );
and ( n76478 , n30349 , n76458 );
and ( n76479 , n76477 , n76478 );
xor ( n76480 , n76477 , n76478 );
xor ( n76481 , n76374 , n76444 );
and ( n76482 , n30354 , n76458 );
and ( n76483 , n76481 , n76482 );
xor ( n76484 , n76481 , n76482 );
xor ( n76485 , n76378 , n76442 );
and ( n76486 , n30359 , n76458 );
and ( n76487 , n76485 , n76486 );
xor ( n76488 , n76485 , n76486 );
xor ( n76489 , n76382 , n76440 );
and ( n76490 , n30364 , n76458 );
and ( n76491 , n76489 , n76490 );
xor ( n76492 , n76489 , n76490 );
xor ( n76493 , n76386 , n76438 );
and ( n76494 , n30369 , n76458 );
and ( n76495 , n76493 , n76494 );
xor ( n76496 , n76493 , n76494 );
xor ( n76497 , n76390 , n76436 );
and ( n76498 , n30374 , n76458 );
and ( n76499 , n76497 , n76498 );
xor ( n76500 , n76497 , n76498 );
xor ( n76501 , n76394 , n76434 );
and ( n76502 , n30379 , n76458 );
and ( n76503 , n76501 , n76502 );
xor ( n76504 , n76501 , n76502 );
xor ( n76505 , n76398 , n76432 );
and ( n76506 , n30384 , n76458 );
and ( n76507 , n76505 , n76506 );
xor ( n76508 , n76505 , n76506 );
xor ( n76509 , n76402 , n76430 );
and ( n76510 , n30389 , n76458 );
and ( n76511 , n76509 , n76510 );
xor ( n76512 , n76509 , n76510 );
xor ( n76513 , n76406 , n76428 );
and ( n76514 , n30394 , n76458 );
and ( n76515 , n76513 , n76514 );
xor ( n76516 , n76513 , n76514 );
xor ( n76517 , n76410 , n76426 );
and ( n76518 , n30399 , n76458 );
and ( n76519 , n76517 , n76518 );
xor ( n76520 , n76517 , n76518 );
xor ( n76521 , n76414 , n76424 );
and ( n76522 , n30404 , n76458 );
and ( n76523 , n76521 , n76522 );
xor ( n76524 , n76521 , n76522 );
xor ( n76525 , n76418 , n76422 );
and ( n76526 , n30409 , n76458 );
and ( n76527 , n76525 , n76526 );
buf ( n76528 , n76527 );
and ( n76529 , n76524 , n76528 );
or ( n76530 , n76523 , n76529 );
and ( n76531 , n76520 , n76530 );
or ( n76532 , n76519 , n76531 );
and ( n76533 , n76516 , n76532 );
or ( n76534 , n76515 , n76533 );
and ( n76535 , n76512 , n76534 );
or ( n76536 , n76511 , n76535 );
and ( n76537 , n76508 , n76536 );
or ( n76538 , n76507 , n76537 );
and ( n76539 , n76504 , n76538 );
or ( n76540 , n76503 , n76539 );
and ( n76541 , n76500 , n76540 );
or ( n76542 , n76499 , n76541 );
and ( n76543 , n76496 , n76542 );
or ( n76544 , n76495 , n76543 );
and ( n76545 , n76492 , n76544 );
or ( n76546 , n76491 , n76545 );
and ( n76547 , n76488 , n76546 );
or ( n76548 , n76487 , n76547 );
and ( n76549 , n76484 , n76548 );
or ( n76550 , n76483 , n76549 );
and ( n76551 , n76480 , n76550 );
or ( n76552 , n76479 , n76551 );
and ( n76553 , n76476 , n76552 );
or ( n76554 , n76475 , n76553 );
and ( n76555 , n76472 , n76554 );
or ( n76556 , n76471 , n76555 );
and ( n76557 , n76468 , n76556 );
or ( n76558 , n76467 , n76557 );
and ( n76559 , n76464 , n76558 );
or ( n76560 , n76463 , n76559 );
xor ( n76561 , n76460 , n76560 );
buf ( n76562 , n17886 );
and ( n76563 , n30329 , n76562 );
xor ( n76564 , n76561 , n76563 );
xor ( n76565 , n76464 , n76558 );
and ( n76566 , n30334 , n76562 );
and ( n76567 , n76565 , n76566 );
xor ( n76568 , n76565 , n76566 );
xor ( n76569 , n76468 , n76556 );
and ( n76570 , n30339 , n76562 );
and ( n76571 , n76569 , n76570 );
xor ( n76572 , n76569 , n76570 );
xor ( n76573 , n76472 , n76554 );
and ( n76574 , n30344 , n76562 );
and ( n76575 , n76573 , n76574 );
xor ( n76576 , n76573 , n76574 );
xor ( n76577 , n76476 , n76552 );
and ( n76578 , n30349 , n76562 );
and ( n76579 , n76577 , n76578 );
xor ( n76580 , n76577 , n76578 );
xor ( n76581 , n76480 , n76550 );
and ( n76582 , n30354 , n76562 );
and ( n76583 , n76581 , n76582 );
xor ( n76584 , n76581 , n76582 );
xor ( n76585 , n76484 , n76548 );
and ( n76586 , n30359 , n76562 );
and ( n76587 , n76585 , n76586 );
xor ( n76588 , n76585 , n76586 );
xor ( n76589 , n76488 , n76546 );
and ( n76590 , n30364 , n76562 );
and ( n76591 , n76589 , n76590 );
xor ( n76592 , n76589 , n76590 );
xor ( n76593 , n76492 , n76544 );
and ( n76594 , n30369 , n76562 );
and ( n76595 , n76593 , n76594 );
xor ( n76596 , n76593 , n76594 );
xor ( n76597 , n76496 , n76542 );
and ( n76598 , n30374 , n76562 );
and ( n76599 , n76597 , n76598 );
xor ( n76600 , n76597 , n76598 );
xor ( n76601 , n76500 , n76540 );
and ( n76602 , n30379 , n76562 );
and ( n76603 , n76601 , n76602 );
xor ( n76604 , n76601 , n76602 );
xor ( n76605 , n76504 , n76538 );
and ( n76606 , n30384 , n76562 );
and ( n76607 , n76605 , n76606 );
xor ( n76608 , n76605 , n76606 );
xor ( n76609 , n76508 , n76536 );
and ( n76610 , n30389 , n76562 );
and ( n76611 , n76609 , n76610 );
xor ( n76612 , n76609 , n76610 );
xor ( n76613 , n76512 , n76534 );
and ( n76614 , n30394 , n76562 );
and ( n76615 , n76613 , n76614 );
xor ( n76616 , n76613 , n76614 );
xor ( n76617 , n76516 , n76532 );
and ( n76618 , n30399 , n76562 );
and ( n76619 , n76617 , n76618 );
xor ( n76620 , n76617 , n76618 );
xor ( n76621 , n76520 , n76530 );
and ( n76622 , n30404 , n76562 );
and ( n76623 , n76621 , n76622 );
xor ( n76624 , n76621 , n76622 );
xor ( n76625 , n76524 , n76528 );
and ( n76626 , n30409 , n76562 );
and ( n76627 , n76625 , n76626 );
buf ( n76628 , n76627 );
and ( n76629 , n76624 , n76628 );
or ( n76630 , n76623 , n76629 );
and ( n76631 , n76620 , n76630 );
or ( n76632 , n76619 , n76631 );
and ( n76633 , n76616 , n76632 );
or ( n76634 , n76615 , n76633 );
and ( n76635 , n76612 , n76634 );
or ( n76636 , n76611 , n76635 );
and ( n76637 , n76608 , n76636 );
or ( n76638 , n76607 , n76637 );
and ( n76639 , n76604 , n76638 );
or ( n76640 , n76603 , n76639 );
and ( n76641 , n76600 , n76640 );
or ( n76642 , n76599 , n76641 );
and ( n76643 , n76596 , n76642 );
or ( n76644 , n76595 , n76643 );
and ( n76645 , n76592 , n76644 );
or ( n76646 , n76591 , n76645 );
and ( n76647 , n76588 , n76646 );
or ( n76648 , n76587 , n76647 );
and ( n76649 , n76584 , n76648 );
or ( n76650 , n76583 , n76649 );
and ( n76651 , n76580 , n76650 );
or ( n76652 , n76579 , n76651 );
and ( n76653 , n76576 , n76652 );
or ( n76654 , n76575 , n76653 );
and ( n76655 , n76572 , n76654 );
or ( n76656 , n76571 , n76655 );
and ( n76657 , n76568 , n76656 );
or ( n76658 , n76567 , n76657 );
xor ( n76659 , n76564 , n76658 );
buf ( n76660 , n17884 );
and ( n76661 , n30334 , n76660 );
xor ( n76662 , n76659 , n76661 );
xor ( n76663 , n76568 , n76656 );
and ( n76664 , n30339 , n76660 );
and ( n76665 , n76663 , n76664 );
xor ( n76666 , n76663 , n76664 );
xor ( n76667 , n76572 , n76654 );
and ( n76668 , n30344 , n76660 );
and ( n76669 , n76667 , n76668 );
xor ( n76670 , n76667 , n76668 );
xor ( n76671 , n76576 , n76652 );
and ( n76672 , n30349 , n76660 );
and ( n76673 , n76671 , n76672 );
xor ( n76674 , n76671 , n76672 );
xor ( n76675 , n76580 , n76650 );
and ( n76676 , n30354 , n76660 );
and ( n76677 , n76675 , n76676 );
xor ( n76678 , n76675 , n76676 );
xor ( n76679 , n76584 , n76648 );
and ( n76680 , n30359 , n76660 );
and ( n76681 , n76679 , n76680 );
xor ( n76682 , n76679 , n76680 );
xor ( n76683 , n76588 , n76646 );
and ( n76684 , n30364 , n76660 );
and ( n76685 , n76683 , n76684 );
xor ( n76686 , n76683 , n76684 );
xor ( n76687 , n76592 , n76644 );
and ( n76688 , n30369 , n76660 );
and ( n76689 , n76687 , n76688 );
xor ( n76690 , n76687 , n76688 );
xor ( n76691 , n76596 , n76642 );
and ( n76692 , n30374 , n76660 );
and ( n76693 , n76691 , n76692 );
xor ( n76694 , n76691 , n76692 );
xor ( n76695 , n76600 , n76640 );
and ( n76696 , n30379 , n76660 );
and ( n76697 , n76695 , n76696 );
xor ( n76698 , n76695 , n76696 );
xor ( n76699 , n76604 , n76638 );
and ( n76700 , n30384 , n76660 );
and ( n76701 , n76699 , n76700 );
xor ( n76702 , n76699 , n76700 );
xor ( n76703 , n76608 , n76636 );
and ( n76704 , n30389 , n76660 );
and ( n76705 , n76703 , n76704 );
xor ( n76706 , n76703 , n76704 );
xor ( n76707 , n76612 , n76634 );
and ( n76708 , n30394 , n76660 );
and ( n76709 , n76707 , n76708 );
xor ( n76710 , n76707 , n76708 );
xor ( n76711 , n76616 , n76632 );
and ( n76712 , n30399 , n76660 );
and ( n76713 , n76711 , n76712 );
xor ( n76714 , n76711 , n76712 );
xor ( n76715 , n76620 , n76630 );
and ( n76716 , n30404 , n76660 );
and ( n76717 , n76715 , n76716 );
xor ( n76718 , n76715 , n76716 );
xor ( n76719 , n76624 , n76628 );
and ( n76720 , n30409 , n76660 );
and ( n76721 , n76719 , n76720 );
buf ( n76722 , n76721 );
and ( n76723 , n76718 , n76722 );
or ( n76724 , n76717 , n76723 );
and ( n76725 , n76714 , n76724 );
or ( n76726 , n76713 , n76725 );
and ( n76727 , n76710 , n76726 );
or ( n76728 , n76709 , n76727 );
and ( n76729 , n76706 , n76728 );
or ( n76730 , n76705 , n76729 );
and ( n76731 , n76702 , n76730 );
or ( n76732 , n76701 , n76731 );
and ( n76733 , n76698 , n76732 );
or ( n76734 , n76697 , n76733 );
and ( n76735 , n76694 , n76734 );
or ( n76736 , n76693 , n76735 );
and ( n76737 , n76690 , n76736 );
or ( n76738 , n76689 , n76737 );
and ( n76739 , n76686 , n76738 );
or ( n76740 , n76685 , n76739 );
and ( n76741 , n76682 , n76740 );
or ( n76742 , n76681 , n76741 );
and ( n76743 , n76678 , n76742 );
or ( n76744 , n76677 , n76743 );
and ( n76745 , n76674 , n76744 );
or ( n76746 , n76673 , n76745 );
and ( n76747 , n76670 , n76746 );
or ( n76748 , n76669 , n76747 );
and ( n76749 , n76666 , n76748 );
or ( n76750 , n76665 , n76749 );
xor ( n76751 , n76662 , n76750 );
buf ( n76752 , n17882 );
and ( n76753 , n30339 , n76752 );
xor ( n76754 , n76751 , n76753 );
xor ( n76755 , n76666 , n76748 );
and ( n76756 , n30344 , n76752 );
and ( n76757 , n76755 , n76756 );
xor ( n76758 , n76755 , n76756 );
xor ( n76759 , n76670 , n76746 );
and ( n76760 , n30349 , n76752 );
and ( n76761 , n76759 , n76760 );
xor ( n76762 , n76759 , n76760 );
xor ( n76763 , n76674 , n76744 );
and ( n76764 , n30354 , n76752 );
and ( n76765 , n76763 , n76764 );
xor ( n76766 , n76763 , n76764 );
xor ( n76767 , n76678 , n76742 );
and ( n76768 , n30359 , n76752 );
and ( n76769 , n76767 , n76768 );
xor ( n76770 , n76767 , n76768 );
xor ( n76771 , n76682 , n76740 );
and ( n76772 , n30364 , n76752 );
and ( n76773 , n76771 , n76772 );
xor ( n76774 , n76771 , n76772 );
xor ( n76775 , n76686 , n76738 );
and ( n76776 , n30369 , n76752 );
and ( n76777 , n76775 , n76776 );
xor ( n76778 , n76775 , n76776 );
xor ( n76779 , n76690 , n76736 );
and ( n76780 , n30374 , n76752 );
and ( n76781 , n76779 , n76780 );
xor ( n76782 , n76779 , n76780 );
xor ( n76783 , n76694 , n76734 );
and ( n76784 , n30379 , n76752 );
and ( n76785 , n76783 , n76784 );
xor ( n76786 , n76783 , n76784 );
xor ( n76787 , n76698 , n76732 );
and ( n76788 , n30384 , n76752 );
and ( n76789 , n76787 , n76788 );
xor ( n76790 , n76787 , n76788 );
xor ( n76791 , n76702 , n76730 );
and ( n76792 , n30389 , n76752 );
and ( n76793 , n76791 , n76792 );
xor ( n76794 , n76791 , n76792 );
xor ( n76795 , n76706 , n76728 );
and ( n76796 , n30394 , n76752 );
and ( n76797 , n76795 , n76796 );
xor ( n76798 , n76795 , n76796 );
xor ( n76799 , n76710 , n76726 );
and ( n76800 , n30399 , n76752 );
and ( n76801 , n76799 , n76800 );
xor ( n76802 , n76799 , n76800 );
xor ( n76803 , n76714 , n76724 );
and ( n76804 , n30404 , n76752 );
and ( n76805 , n76803 , n76804 );
xor ( n76806 , n76803 , n76804 );
xor ( n76807 , n76718 , n76722 );
and ( n76808 , n30409 , n76752 );
and ( n76809 , n76807 , n76808 );
buf ( n76810 , n76809 );
and ( n76811 , n76806 , n76810 );
or ( n76812 , n76805 , n76811 );
and ( n76813 , n76802 , n76812 );
or ( n76814 , n76801 , n76813 );
and ( n76815 , n76798 , n76814 );
or ( n76816 , n76797 , n76815 );
and ( n76817 , n76794 , n76816 );
or ( n76818 , n76793 , n76817 );
and ( n76819 , n76790 , n76818 );
or ( n76820 , n76789 , n76819 );
and ( n76821 , n76786 , n76820 );
or ( n76822 , n76785 , n76821 );
and ( n76823 , n76782 , n76822 );
or ( n76824 , n76781 , n76823 );
and ( n76825 , n76778 , n76824 );
or ( n76826 , n76777 , n76825 );
and ( n76827 , n76774 , n76826 );
or ( n76828 , n76773 , n76827 );
and ( n76829 , n76770 , n76828 );
or ( n76830 , n76769 , n76829 );
and ( n76831 , n76766 , n76830 );
or ( n76832 , n76765 , n76831 );
and ( n76833 , n76762 , n76832 );
or ( n76834 , n76761 , n76833 );
and ( n76835 , n76758 , n76834 );
or ( n76836 , n76757 , n76835 );
xor ( n76837 , n76754 , n76836 );
buf ( n76838 , n17880 );
and ( n76839 , n30344 , n76838 );
xor ( n76840 , n76837 , n76839 );
xor ( n76841 , n76758 , n76834 );
and ( n76842 , n30349 , n76838 );
and ( n76843 , n76841 , n76842 );
xor ( n76844 , n76841 , n76842 );
xor ( n76845 , n76762 , n76832 );
and ( n76846 , n30354 , n76838 );
and ( n76847 , n76845 , n76846 );
xor ( n76848 , n76845 , n76846 );
xor ( n76849 , n76766 , n76830 );
and ( n76850 , n30359 , n76838 );
and ( n76851 , n76849 , n76850 );
xor ( n76852 , n76849 , n76850 );
xor ( n76853 , n76770 , n76828 );
and ( n76854 , n30364 , n76838 );
and ( n76855 , n76853 , n76854 );
xor ( n76856 , n76853 , n76854 );
xor ( n76857 , n76774 , n76826 );
and ( n76858 , n30369 , n76838 );
and ( n76859 , n76857 , n76858 );
xor ( n76860 , n76857 , n76858 );
xor ( n76861 , n76778 , n76824 );
and ( n76862 , n30374 , n76838 );
and ( n76863 , n76861 , n76862 );
xor ( n76864 , n76861 , n76862 );
xor ( n76865 , n76782 , n76822 );
and ( n76866 , n30379 , n76838 );
and ( n76867 , n76865 , n76866 );
xor ( n76868 , n76865 , n76866 );
xor ( n76869 , n76786 , n76820 );
and ( n76870 , n30384 , n76838 );
and ( n76871 , n76869 , n76870 );
xor ( n76872 , n76869 , n76870 );
xor ( n76873 , n76790 , n76818 );
and ( n76874 , n30389 , n76838 );
and ( n76875 , n76873 , n76874 );
xor ( n76876 , n76873 , n76874 );
xor ( n76877 , n76794 , n76816 );
and ( n76878 , n30394 , n76838 );
and ( n76879 , n76877 , n76878 );
xor ( n76880 , n76877 , n76878 );
xor ( n76881 , n76798 , n76814 );
and ( n76882 , n30399 , n76838 );
and ( n76883 , n76881 , n76882 );
xor ( n76884 , n76881 , n76882 );
xor ( n76885 , n76802 , n76812 );
and ( n76886 , n30404 , n76838 );
and ( n76887 , n76885 , n76886 );
xor ( n76888 , n76885 , n76886 );
xor ( n76889 , n76806 , n76810 );
and ( n76890 , n30409 , n76838 );
and ( n76891 , n76889 , n76890 );
buf ( n76892 , n76891 );
and ( n76893 , n76888 , n76892 );
or ( n76894 , n76887 , n76893 );
and ( n76895 , n76884 , n76894 );
or ( n76896 , n76883 , n76895 );
and ( n76897 , n76880 , n76896 );
or ( n76898 , n76879 , n76897 );
and ( n76899 , n76876 , n76898 );
or ( n76900 , n76875 , n76899 );
and ( n76901 , n76872 , n76900 );
or ( n76902 , n76871 , n76901 );
and ( n76903 , n76868 , n76902 );
or ( n76904 , n76867 , n76903 );
and ( n76905 , n76864 , n76904 );
or ( n76906 , n76863 , n76905 );
and ( n76907 , n76860 , n76906 );
or ( n76908 , n76859 , n76907 );
and ( n76909 , n76856 , n76908 );
or ( n76910 , n76855 , n76909 );
and ( n76911 , n76852 , n76910 );
or ( n76912 , n76851 , n76911 );
and ( n76913 , n76848 , n76912 );
or ( n76914 , n76847 , n76913 );
and ( n76915 , n76844 , n76914 );
or ( n76916 , n76843 , n76915 );
xor ( n76917 , n76840 , n76916 );
buf ( n76918 , n17878 );
and ( n76919 , n30349 , n76918 );
xor ( n76920 , n76917 , n76919 );
xor ( n76921 , n76844 , n76914 );
and ( n76922 , n30354 , n76918 );
and ( n76923 , n76921 , n76922 );
xor ( n76924 , n76921 , n76922 );
xor ( n76925 , n76848 , n76912 );
and ( n76926 , n30359 , n76918 );
and ( n76927 , n76925 , n76926 );
xor ( n76928 , n76925 , n76926 );
xor ( n76929 , n76852 , n76910 );
and ( n76930 , n30364 , n76918 );
and ( n76931 , n76929 , n76930 );
xor ( n76932 , n76929 , n76930 );
xor ( n76933 , n76856 , n76908 );
and ( n76934 , n30369 , n76918 );
and ( n76935 , n76933 , n76934 );
xor ( n76936 , n76933 , n76934 );
xor ( n76937 , n76860 , n76906 );
and ( n76938 , n30374 , n76918 );
and ( n76939 , n76937 , n76938 );
xor ( n76940 , n76937 , n76938 );
xor ( n76941 , n76864 , n76904 );
and ( n76942 , n30379 , n76918 );
and ( n76943 , n76941 , n76942 );
xor ( n76944 , n76941 , n76942 );
xor ( n76945 , n76868 , n76902 );
and ( n76946 , n30384 , n76918 );
and ( n76947 , n76945 , n76946 );
xor ( n76948 , n76945 , n76946 );
xor ( n76949 , n76872 , n76900 );
and ( n76950 , n30389 , n76918 );
and ( n76951 , n76949 , n76950 );
xor ( n76952 , n76949 , n76950 );
xor ( n76953 , n76876 , n76898 );
and ( n76954 , n30394 , n76918 );
and ( n76955 , n76953 , n76954 );
xor ( n76956 , n76953 , n76954 );
xor ( n76957 , n76880 , n76896 );
and ( n76958 , n30399 , n76918 );
and ( n76959 , n76957 , n76958 );
xor ( n76960 , n76957 , n76958 );
xor ( n76961 , n76884 , n76894 );
and ( n76962 , n30404 , n76918 );
and ( n76963 , n76961 , n76962 );
xor ( n76964 , n76961 , n76962 );
xor ( n76965 , n76888 , n76892 );
and ( n76966 , n30409 , n76918 );
and ( n76967 , n76965 , n76966 );
buf ( n76968 , n76967 );
and ( n76969 , n76964 , n76968 );
or ( n76970 , n76963 , n76969 );
and ( n76971 , n76960 , n76970 );
or ( n76972 , n76959 , n76971 );
and ( n76973 , n76956 , n76972 );
or ( n76974 , n76955 , n76973 );
and ( n76975 , n76952 , n76974 );
or ( n76976 , n76951 , n76975 );
and ( n76977 , n76948 , n76976 );
or ( n76978 , n76947 , n76977 );
and ( n76979 , n76944 , n76978 );
or ( n76980 , n76943 , n76979 );
and ( n76981 , n76940 , n76980 );
or ( n76982 , n76939 , n76981 );
and ( n76983 , n76936 , n76982 );
or ( n76984 , n76935 , n76983 );
and ( n76985 , n76932 , n76984 );
or ( n76986 , n76931 , n76985 );
and ( n76987 , n76928 , n76986 );
or ( n76988 , n76927 , n76987 );
and ( n76989 , n76924 , n76988 );
or ( n76990 , n76923 , n76989 );
xor ( n76991 , n76920 , n76990 );
buf ( n76992 , n17876 );
and ( n76993 , n30354 , n76992 );
xor ( n76994 , n76991 , n76993 );
xor ( n76995 , n76924 , n76988 );
and ( n76996 , n30359 , n76992 );
and ( n76997 , n76995 , n76996 );
xor ( n76998 , n76995 , n76996 );
xor ( n76999 , n76928 , n76986 );
and ( n77000 , n30364 , n76992 );
and ( n77001 , n76999 , n77000 );
xor ( n77002 , n76999 , n77000 );
xor ( n77003 , n76932 , n76984 );
and ( n77004 , n30369 , n76992 );
and ( n77005 , n77003 , n77004 );
xor ( n77006 , n77003 , n77004 );
xor ( n77007 , n76936 , n76982 );
and ( n77008 , n30374 , n76992 );
and ( n77009 , n77007 , n77008 );
xor ( n77010 , n77007 , n77008 );
xor ( n77011 , n76940 , n76980 );
and ( n77012 , n30379 , n76992 );
and ( n77013 , n77011 , n77012 );
xor ( n77014 , n77011 , n77012 );
xor ( n77015 , n76944 , n76978 );
and ( n77016 , n30384 , n76992 );
and ( n77017 , n77015 , n77016 );
xor ( n77018 , n77015 , n77016 );
xor ( n77019 , n76948 , n76976 );
and ( n77020 , n30389 , n76992 );
and ( n77021 , n77019 , n77020 );
xor ( n77022 , n77019 , n77020 );
xor ( n77023 , n76952 , n76974 );
and ( n77024 , n30394 , n76992 );
and ( n77025 , n77023 , n77024 );
xor ( n77026 , n77023 , n77024 );
xor ( n77027 , n76956 , n76972 );
and ( n77028 , n30399 , n76992 );
and ( n77029 , n77027 , n77028 );
xor ( n77030 , n77027 , n77028 );
xor ( n77031 , n76960 , n76970 );
and ( n77032 , n30404 , n76992 );
and ( n77033 , n77031 , n77032 );
xor ( n77034 , n77031 , n77032 );
xor ( n77035 , n76964 , n76968 );
and ( n77036 , n30409 , n76992 );
and ( n77037 , n77035 , n77036 );
buf ( n77038 , n77037 );
and ( n77039 , n77034 , n77038 );
or ( n77040 , n77033 , n77039 );
and ( n77041 , n77030 , n77040 );
or ( n77042 , n77029 , n77041 );
and ( n77043 , n77026 , n77042 );
or ( n77044 , n77025 , n77043 );
and ( n77045 , n77022 , n77044 );
or ( n77046 , n77021 , n77045 );
and ( n77047 , n77018 , n77046 );
or ( n77048 , n77017 , n77047 );
and ( n77049 , n77014 , n77048 );
or ( n77050 , n77013 , n77049 );
and ( n77051 , n77010 , n77050 );
or ( n77052 , n77009 , n77051 );
and ( n77053 , n77006 , n77052 );
or ( n77054 , n77005 , n77053 );
and ( n77055 , n77002 , n77054 );
or ( n77056 , n77001 , n77055 );
and ( n77057 , n76998 , n77056 );
or ( n77058 , n76997 , n77057 );
xor ( n77059 , n76994 , n77058 );
buf ( n77060 , n17874 );
and ( n77061 , n30359 , n77060 );
xor ( n77062 , n77059 , n77061 );
xor ( n77063 , n76998 , n77056 );
and ( n77064 , n30364 , n77060 );
and ( n77065 , n77063 , n77064 );
xor ( n77066 , n77063 , n77064 );
xor ( n77067 , n77002 , n77054 );
and ( n77068 , n30369 , n77060 );
and ( n77069 , n77067 , n77068 );
xor ( n77070 , n77067 , n77068 );
xor ( n77071 , n77006 , n77052 );
and ( n77072 , n30374 , n77060 );
and ( n77073 , n77071 , n77072 );
xor ( n77074 , n77071 , n77072 );
xor ( n77075 , n77010 , n77050 );
and ( n77076 , n30379 , n77060 );
and ( n77077 , n77075 , n77076 );
xor ( n77078 , n77075 , n77076 );
xor ( n77079 , n77014 , n77048 );
and ( n77080 , n30384 , n77060 );
and ( n77081 , n77079 , n77080 );
xor ( n77082 , n77079 , n77080 );
xor ( n77083 , n77018 , n77046 );
and ( n77084 , n30389 , n77060 );
and ( n77085 , n77083 , n77084 );
xor ( n77086 , n77083 , n77084 );
xor ( n77087 , n77022 , n77044 );
and ( n77088 , n30394 , n77060 );
and ( n77089 , n77087 , n77088 );
xor ( n77090 , n77087 , n77088 );
xor ( n77091 , n77026 , n77042 );
and ( n77092 , n30399 , n77060 );
and ( n77093 , n77091 , n77092 );
xor ( n77094 , n77091 , n77092 );
xor ( n77095 , n77030 , n77040 );
and ( n77096 , n30404 , n77060 );
and ( n77097 , n77095 , n77096 );
xor ( n77098 , n77095 , n77096 );
xor ( n77099 , n77034 , n77038 );
and ( n77100 , n30409 , n77060 );
and ( n77101 , n77099 , n77100 );
buf ( n77102 , n77101 );
and ( n77103 , n77098 , n77102 );
or ( n77104 , n77097 , n77103 );
and ( n77105 , n77094 , n77104 );
or ( n77106 , n77093 , n77105 );
and ( n77107 , n77090 , n77106 );
or ( n77108 , n77089 , n77107 );
and ( n77109 , n77086 , n77108 );
or ( n77110 , n77085 , n77109 );
and ( n77111 , n77082 , n77110 );
or ( n77112 , n77081 , n77111 );
and ( n77113 , n77078 , n77112 );
or ( n77114 , n77077 , n77113 );
and ( n77115 , n77074 , n77114 );
or ( n77116 , n77073 , n77115 );
and ( n77117 , n77070 , n77116 );
or ( n77118 , n77069 , n77117 );
and ( n77119 , n77066 , n77118 );
or ( n77120 , n77065 , n77119 );
xor ( n77121 , n77062 , n77120 );
buf ( n77122 , n17872 );
and ( n77123 , n30364 , n77122 );
xor ( n77124 , n77121 , n77123 );
xor ( n77125 , n77066 , n77118 );
and ( n77126 , n30369 , n77122 );
and ( n77127 , n77125 , n77126 );
xor ( n77128 , n77125 , n77126 );
xor ( n77129 , n77070 , n77116 );
and ( n77130 , n30374 , n77122 );
and ( n77131 , n77129 , n77130 );
xor ( n77132 , n77129 , n77130 );
xor ( n77133 , n77074 , n77114 );
and ( n77134 , n30379 , n77122 );
and ( n77135 , n77133 , n77134 );
xor ( n77136 , n77133 , n77134 );
xor ( n77137 , n77078 , n77112 );
and ( n77138 , n30384 , n77122 );
and ( n77139 , n77137 , n77138 );
xor ( n77140 , n77137 , n77138 );
xor ( n77141 , n77082 , n77110 );
and ( n77142 , n30389 , n77122 );
and ( n77143 , n77141 , n77142 );
xor ( n77144 , n77141 , n77142 );
xor ( n77145 , n77086 , n77108 );
and ( n77146 , n30394 , n77122 );
and ( n77147 , n77145 , n77146 );
xor ( n77148 , n77145 , n77146 );
xor ( n77149 , n77090 , n77106 );
and ( n77150 , n30399 , n77122 );
and ( n77151 , n77149 , n77150 );
xor ( n77152 , n77149 , n77150 );
xor ( n77153 , n77094 , n77104 );
and ( n77154 , n30404 , n77122 );
and ( n77155 , n77153 , n77154 );
xor ( n77156 , n77153 , n77154 );
xor ( n77157 , n77098 , n77102 );
and ( n77158 , n30409 , n77122 );
and ( n77159 , n77157 , n77158 );
buf ( n77160 , n77159 );
and ( n77161 , n77156 , n77160 );
or ( n77162 , n77155 , n77161 );
and ( n77163 , n77152 , n77162 );
or ( n77164 , n77151 , n77163 );
and ( n77165 , n77148 , n77164 );
or ( n77166 , n77147 , n77165 );
and ( n77167 , n77144 , n77166 );
or ( n77168 , n77143 , n77167 );
and ( n77169 , n77140 , n77168 );
or ( n77170 , n77139 , n77169 );
and ( n77171 , n77136 , n77170 );
or ( n77172 , n77135 , n77171 );
and ( n77173 , n77132 , n77172 );
or ( n77174 , n77131 , n77173 );
and ( n77175 , n77128 , n77174 );
or ( n77176 , n77127 , n77175 );
xor ( n77177 , n77124 , n77176 );
buf ( n77178 , n17870 );
and ( n77179 , n30369 , n77178 );
xor ( n77180 , n77177 , n77179 );
xor ( n77181 , n77128 , n77174 );
and ( n77182 , n30374 , n77178 );
and ( n77183 , n77181 , n77182 );
xor ( n77184 , n77181 , n77182 );
xor ( n77185 , n77132 , n77172 );
and ( n77186 , n30379 , n77178 );
and ( n77187 , n77185 , n77186 );
xor ( n77188 , n77185 , n77186 );
xor ( n77189 , n77136 , n77170 );
and ( n77190 , n30384 , n77178 );
and ( n77191 , n77189 , n77190 );
xor ( n77192 , n77189 , n77190 );
xor ( n77193 , n77140 , n77168 );
and ( n77194 , n30389 , n77178 );
and ( n77195 , n77193 , n77194 );
xor ( n77196 , n77193 , n77194 );
xor ( n77197 , n77144 , n77166 );
and ( n77198 , n30394 , n77178 );
and ( n77199 , n77197 , n77198 );
xor ( n77200 , n77197 , n77198 );
xor ( n77201 , n77148 , n77164 );
and ( n77202 , n30399 , n77178 );
and ( n77203 , n77201 , n77202 );
xor ( n77204 , n77201 , n77202 );
xor ( n77205 , n77152 , n77162 );
and ( n77206 , n30404 , n77178 );
and ( n77207 , n77205 , n77206 );
xor ( n77208 , n77205 , n77206 );
xor ( n77209 , n77156 , n77160 );
and ( n77210 , n30409 , n77178 );
and ( n77211 , n77209 , n77210 );
buf ( n77212 , n77211 );
and ( n77213 , n77208 , n77212 );
or ( n77214 , n77207 , n77213 );
and ( n77215 , n77204 , n77214 );
or ( n77216 , n77203 , n77215 );
and ( n77217 , n77200 , n77216 );
or ( n77218 , n77199 , n77217 );
and ( n77219 , n77196 , n77218 );
or ( n77220 , n77195 , n77219 );
and ( n77221 , n77192 , n77220 );
or ( n77222 , n77191 , n77221 );
and ( n77223 , n77188 , n77222 );
or ( n77224 , n77187 , n77223 );
and ( n77225 , n77184 , n77224 );
or ( n77226 , n77183 , n77225 );
xor ( n77227 , n77180 , n77226 );
buf ( n77228 , n17868 );
and ( n77229 , n30374 , n77228 );
xor ( n77230 , n77227 , n77229 );
xor ( n77231 , n77184 , n77224 );
and ( n77232 , n30379 , n77228 );
and ( n77233 , n77231 , n77232 );
xor ( n77234 , n77231 , n77232 );
xor ( n77235 , n77188 , n77222 );
and ( n77236 , n30384 , n77228 );
and ( n77237 , n77235 , n77236 );
xor ( n77238 , n77235 , n77236 );
xor ( n77239 , n77192 , n77220 );
and ( n77240 , n30389 , n77228 );
and ( n77241 , n77239 , n77240 );
xor ( n77242 , n77239 , n77240 );
xor ( n77243 , n77196 , n77218 );
and ( n77244 , n30394 , n77228 );
and ( n77245 , n77243 , n77244 );
xor ( n77246 , n77243 , n77244 );
xor ( n77247 , n77200 , n77216 );
and ( n77248 , n30399 , n77228 );
and ( n77249 , n77247 , n77248 );
xor ( n77250 , n77247 , n77248 );
xor ( n77251 , n77204 , n77214 );
and ( n77252 , n30404 , n77228 );
and ( n77253 , n77251 , n77252 );
xor ( n77254 , n77251 , n77252 );
xor ( n77255 , n77208 , n77212 );
and ( n77256 , n30409 , n77228 );
and ( n77257 , n77255 , n77256 );
buf ( n77258 , n77257 );
and ( n77259 , n77254 , n77258 );
or ( n77260 , n77253 , n77259 );
and ( n77261 , n77250 , n77260 );
or ( n77262 , n77249 , n77261 );
and ( n77263 , n77246 , n77262 );
or ( n77264 , n77245 , n77263 );
and ( n77265 , n77242 , n77264 );
or ( n77266 , n77241 , n77265 );
and ( n77267 , n77238 , n77266 );
or ( n77268 , n77237 , n77267 );
and ( n77269 , n77234 , n77268 );
or ( n77270 , n77233 , n77269 );
xor ( n77271 , n77230 , n77270 );
buf ( n77272 , n17866 );
and ( n77273 , n30379 , n77272 );
xor ( n77274 , n77271 , n77273 );
xor ( n77275 , n77234 , n77268 );
and ( n77276 , n30384 , n77272 );
and ( n77277 , n77275 , n77276 );
xor ( n77278 , n77275 , n77276 );
xor ( n77279 , n77238 , n77266 );
and ( n77280 , n30389 , n77272 );
and ( n77281 , n77279 , n77280 );
xor ( n77282 , n77279 , n77280 );
xor ( n77283 , n77242 , n77264 );
and ( n77284 , n30394 , n77272 );
and ( n77285 , n77283 , n77284 );
xor ( n77286 , n77283 , n77284 );
xor ( n77287 , n77246 , n77262 );
and ( n77288 , n30399 , n77272 );
and ( n77289 , n77287 , n77288 );
xor ( n77290 , n77287 , n77288 );
xor ( n77291 , n77250 , n77260 );
and ( n77292 , n30404 , n77272 );
and ( n77293 , n77291 , n77292 );
xor ( n77294 , n77291 , n77292 );
xor ( n77295 , n77254 , n77258 );
and ( n77296 , n30409 , n77272 );
and ( n77297 , n77295 , n77296 );
buf ( n77298 , n77297 );
and ( n77299 , n77294 , n77298 );
or ( n77300 , n77293 , n77299 );
and ( n77301 , n77290 , n77300 );
or ( n77302 , n77289 , n77301 );
and ( n77303 , n77286 , n77302 );
or ( n77304 , n77285 , n77303 );
and ( n77305 , n77282 , n77304 );
or ( n77306 , n77281 , n77305 );
and ( n77307 , n77278 , n77306 );
or ( n77308 , n77277 , n77307 );
xor ( n77309 , n77274 , n77308 );
buf ( n77310 , n17864 );
and ( n77311 , n30384 , n77310 );
xor ( n77312 , n77309 , n77311 );
xor ( n77313 , n77278 , n77306 );
and ( n77314 , n30389 , n77310 );
and ( n77315 , n77313 , n77314 );
xor ( n77316 , n77313 , n77314 );
xor ( n77317 , n77282 , n77304 );
and ( n77318 , n30394 , n77310 );
and ( n77319 , n77317 , n77318 );
xor ( n77320 , n77317 , n77318 );
xor ( n77321 , n77286 , n77302 );
and ( n77322 , n30399 , n77310 );
and ( n77323 , n77321 , n77322 );
xor ( n77324 , n77321 , n77322 );
xor ( n77325 , n77290 , n77300 );
and ( n77326 , n30404 , n77310 );
and ( n77327 , n77325 , n77326 );
xor ( n77328 , n77325 , n77326 );
xor ( n77329 , n77294 , n77298 );
and ( n77330 , n30409 , n77310 );
and ( n77331 , n77329 , n77330 );
buf ( n77332 , n77331 );
and ( n77333 , n77328 , n77332 );
or ( n77334 , n77327 , n77333 );
and ( n77335 , n77324 , n77334 );
or ( n77336 , n77323 , n77335 );
and ( n77337 , n77320 , n77336 );
or ( n77338 , n77319 , n77337 );
and ( n77339 , n77316 , n77338 );
or ( n77340 , n77315 , n77339 );
xor ( n77341 , n77312 , n77340 );
buf ( n77342 , n17862 );
and ( n77343 , n30389 , n77342 );
xor ( n77344 , n77341 , n77343 );
xor ( n77345 , n77316 , n77338 );
and ( n77346 , n30394 , n77342 );
and ( n77347 , n77345 , n77346 );
xor ( n77348 , n77345 , n77346 );
xor ( n77349 , n77320 , n77336 );
and ( n77350 , n30399 , n77342 );
and ( n77351 , n77349 , n77350 );
xor ( n77352 , n77349 , n77350 );
xor ( n77353 , n77324 , n77334 );
and ( n77354 , n30404 , n77342 );
and ( n77355 , n77353 , n77354 );
xor ( n77356 , n77353 , n77354 );
xor ( n77357 , n77328 , n77332 );
and ( n77358 , n30409 , n77342 );
and ( n77359 , n77357 , n77358 );
buf ( n77360 , n77359 );
and ( n77361 , n77356 , n77360 );
or ( n77362 , n77355 , n77361 );
and ( n77363 , n77352 , n77362 );
or ( n77364 , n77351 , n77363 );
and ( n77365 , n77348 , n77364 );
or ( n77366 , n77347 , n77365 );
xor ( n77367 , n77344 , n77366 );
buf ( n77368 , n17860 );
and ( n77369 , n30394 , n77368 );
xor ( n77370 , n77367 , n77369 );
xor ( n77371 , n77348 , n77364 );
and ( n77372 , n30399 , n77368 );
and ( n77373 , n77371 , n77372 );
xor ( n77374 , n77371 , n77372 );
xor ( n77375 , n77352 , n77362 );
and ( n77376 , n30404 , n77368 );
and ( n77377 , n77375 , n77376 );
xor ( n77378 , n77375 , n77376 );
xor ( n77379 , n77356 , n77360 );
and ( n77380 , n30409 , n77368 );
and ( n77381 , n77379 , n77380 );
buf ( n77382 , n77381 );
and ( n77383 , n77378 , n77382 );
or ( n77384 , n77377 , n77383 );
and ( n77385 , n77374 , n77384 );
or ( n77386 , n77373 , n77385 );
xor ( n77387 , n77370 , n77386 );
buf ( n77388 , n17858 );
and ( n77389 , n30399 , n77388 );
xor ( n77390 , n77387 , n77389 );
xor ( n77391 , n77374 , n77384 );
and ( n77392 , n30404 , n77388 );
and ( n77393 , n77391 , n77392 );
xor ( n77394 , n77391 , n77392 );
xor ( n77395 , n77378 , n77382 );
and ( n77396 , n30409 , n77388 );
and ( n77397 , n77395 , n77396 );
buf ( n77398 , n77397 );
and ( n77399 , n77394 , n77398 );
or ( n77400 , n77393 , n77399 );
xor ( n77401 , n77390 , n77400 );
buf ( n77402 , n17856 );
and ( n77403 , n30404 , n77402 );
xor ( n77404 , n77401 , n77403 );
xor ( n77405 , n77394 , n77398 );
and ( n77406 , n30409 , n77402 );
and ( n77407 , n77405 , n77406 );
buf ( n77408 , n77407 );
xor ( n77409 , n77404 , n77408 );
buf ( n77410 , n17854 );
and ( n77411 , n30409 , n77410 );
xor ( n77412 , n77409 , n77411 );
buf ( n77413 , n77412 );
buf ( n77414 , n77413 );
buf ( n77415 , n77414 );
buf ( n77416 , n77415 );
xor ( n77417 , n77405 , n77406 );
buf ( n77418 , n77417 );
buf ( n77419 , n77418 );
buf ( n77420 , n77419 );
buf ( n77421 , n77420 );
xor ( n77422 , n77395 , n77396 );
buf ( n77423 , n77422 );
buf ( n77424 , n77423 );
buf ( n77425 , n77424 );
buf ( n77426 , n77425 );
xor ( n77427 , n77379 , n77380 );
buf ( n77428 , n77427 );
buf ( n77429 , n77428 );
buf ( n77430 , n77429 );
buf ( n77431 , n77430 );
xor ( n77432 , n77357 , n77358 );
buf ( n77433 , n77432 );
buf ( n77434 , n77433 );
buf ( n77435 , n77434 );
buf ( n77436 , n77435 );
xor ( n77437 , n77329 , n77330 );
buf ( n77438 , n77437 );
buf ( n77439 , n77438 );
buf ( n77440 , n77439 );
buf ( n77441 , n77440 );
xor ( n77442 , n77295 , n77296 );
buf ( n77443 , n77442 );
buf ( n77444 , n77443 );
buf ( n77445 , n77444 );
buf ( n77446 , n77445 );
xor ( n77447 , n77255 , n77256 );
buf ( n77448 , n77447 );
buf ( n77449 , n77448 );
buf ( n77450 , n77449 );
buf ( n77451 , n77450 );
xor ( n77452 , n77209 , n77210 );
buf ( n77453 , n77452 );
buf ( n77454 , n77453 );
buf ( n77455 , n77454 );
buf ( n77456 , n77455 );
xor ( n77457 , n77157 , n77158 );
buf ( n77458 , n77457 );
buf ( n77459 , n77458 );
buf ( n77460 , n77459 );
buf ( n77461 , n77460 );
xor ( n77462 , n77099 , n77100 );
buf ( n77463 , n77462 );
buf ( n77464 , n77463 );
buf ( n77465 , n77464 );
buf ( n77466 , n77465 );
xor ( n77467 , n77035 , n77036 );
buf ( n77468 , n77467 );
buf ( n77469 , n77468 );
buf ( n77470 , n77469 );
buf ( n77471 , n77470 );
xor ( n77472 , n76965 , n76966 );
buf ( n77473 , n77472 );
buf ( n77474 , n77473 );
buf ( n77475 , n77474 );
buf ( n77476 , n77475 );
xor ( n77477 , n76889 , n76890 );
buf ( n77478 , n77477 );
buf ( n77479 , n77478 );
buf ( n77480 , n77479 );
buf ( n77481 , n77480 );
xor ( n77482 , n76807 , n76808 );
buf ( n77483 , n77482 );
buf ( n77484 , n77483 );
buf ( n77485 , n77484 );
buf ( n77486 , n77485 );
xor ( n77487 , n76719 , n76720 );
buf ( n77488 , n77487 );
buf ( n77489 , n77488 );
buf ( n77490 , n77489 );
buf ( n77491 , n77490 );
xor ( n77492 , n76625 , n76626 );
buf ( n77493 , n77492 );
buf ( n77494 , n77493 );
buf ( n77495 , n77494 );
buf ( n77496 , n77495 );
xor ( n77497 , n76525 , n76526 );
buf ( n77498 , n77497 );
buf ( n77499 , n77498 );
buf ( n77500 , n77499 );
buf ( n77501 , n77500 );
xor ( n77502 , n76419 , n76420 );
buf ( n77503 , n77502 );
buf ( n77504 , n77503 );
buf ( n77505 , n77504 );
buf ( n77506 , n77505 );
xor ( n77507 , n76307 , n76308 );
buf ( n77508 , n77507 );
buf ( n77509 , n77508 );
buf ( n77510 , n77509 );
buf ( n77511 , n77510 );
xor ( n77512 , n76189 , n76190 );
buf ( n77513 , n77512 );
buf ( n77514 , n77513 );
buf ( n77515 , n77514 );
buf ( n77516 , n77515 );
xor ( n77517 , n76065 , n76066 );
buf ( n77518 , n77517 );
buf ( n77519 , n77518 );
buf ( n77520 , n77519 );
buf ( n77521 , n77520 );
xor ( n77522 , n75935 , n75936 );
buf ( n77523 , n77522 );
buf ( n77524 , n77523 );
buf ( n77525 , n77524 );
buf ( n77526 , n77525 );
xor ( n77527 , n75799 , n75800 );
buf ( n77528 , n77527 );
buf ( n77529 , n77528 );
buf ( n77530 , n77529 );
buf ( n77531 , n77530 );
xor ( n77532 , n75657 , n75658 );
buf ( n77533 , n77532 );
buf ( n77534 , n77533 );
buf ( n77535 , n77534 );
buf ( n77536 , n77535 );
xor ( n77537 , n75509 , n75510 );
buf ( n77538 , n77537 );
buf ( n77539 , n77538 );
buf ( n77540 , n77539 );
buf ( n77541 , n77540 );
xor ( n77542 , n75355 , n75356 );
buf ( n77543 , n77542 );
buf ( n77544 , n77543 );
buf ( n77545 , n77544 );
buf ( n77546 , n77545 );
xor ( n77547 , n75195 , n75196 );
buf ( n77548 , n77547 );
buf ( n77549 , n77548 );
buf ( n77550 , n77549 );
buf ( n77551 , n77550 );
xor ( n77552 , n75029 , n75030 );
buf ( n77553 , n77552 );
buf ( n77554 , n77553 );
buf ( n77555 , n77554 );
buf ( n77556 , n77555 );
xor ( n77557 , n74857 , n74858 );
buf ( n77558 , n77557 );
buf ( n77559 , n77558 );
buf ( n77560 , n77559 );
buf ( n77561 , n77560 );
xor ( n77562 , n74679 , n74680 );
buf ( n77563 , n77562 );
buf ( n77564 , n77563 );
buf ( n77565 , n77564 );
buf ( n77566 , n77565 );
xor ( n77567 , n74495 , n74496 );
buf ( n77568 , n77567 );
buf ( n77569 , n77568 );
buf ( n77570 , n77569 );
buf ( n77571 , n77570 );
xor ( n77572 , n74305 , n74306 );
buf ( n77573 , n77572 );
buf ( n77574 , n77573 );
buf ( n77575 , n77574 );
buf ( n77576 , n77575 );
xor ( n77577 , n74109 , n74110 );
buf ( n77578 , n77577 );
buf ( n77579 , n77578 );
buf ( n77580 , n77579 );
buf ( n77581 , n77580 );
xor ( n77582 , n73907 , n73908 );
buf ( n77583 , n77582 );
buf ( n77584 , n77583 );
buf ( n77585 , n77584 );
buf ( n77586 , n77585 );
xor ( n77587 , n73699 , n73700 );
buf ( n77588 , n77587 );
buf ( n77589 , n77588 );
buf ( n77590 , n77589 );
buf ( n77591 , n77590 );
xor ( n77592 , n73485 , n73486 );
buf ( n77593 , n77592 );
buf ( n77594 , n77593 );
buf ( n77595 , n77594 );
buf ( n77596 , n77595 );
xor ( n77597 , n73265 , n73266 );
buf ( n77598 , n77597 );
buf ( n77599 , n77598 );
buf ( n77600 , n77599 );
buf ( n77601 , n77600 );
xor ( n77602 , n73039 , n73040 );
buf ( n77603 , n77602 );
buf ( n77604 , n77603 );
buf ( n77605 , n77604 );
buf ( n77606 , n77605 );
xor ( n77607 , n72807 , n72808 );
buf ( n77608 , n77607 );
buf ( n77609 , n77608 );
buf ( n77610 , n77609 );
buf ( n77611 , n77610 );
xor ( n77612 , n72569 , n72570 );
buf ( n77613 , n77612 );
buf ( n77614 , n77613 );
buf ( n77615 , n77614 );
buf ( n77616 , n77615 );
xor ( n77617 , n72325 , n72326 );
buf ( n77618 , n77617 );
buf ( n77619 , n77618 );
buf ( n77620 , n77619 );
buf ( n77621 , n77620 );
xor ( n77622 , n72075 , n72076 );
buf ( n77623 , n77622 );
buf ( n77624 , n77623 );
buf ( n77625 , n77624 );
buf ( n77626 , n77625 );
xor ( n77627 , n71819 , n71820 );
buf ( n77628 , n77627 );
buf ( n77629 , n77628 );
buf ( n77630 , n77629 );
buf ( n77631 , n77630 );
xor ( n77632 , n71557 , n71558 );
buf ( n77633 , n77632 );
buf ( n77634 , n77633 );
buf ( n77635 , n77634 );
buf ( n77636 , n77635 );
xor ( n77637 , n71289 , n71290 );
buf ( n77638 , n77637 );
buf ( n77639 , n77638 );
buf ( n77640 , n77639 );
buf ( n77641 , n77640 );
xor ( n77642 , n71015 , n71016 );
buf ( n77643 , n77642 );
buf ( n77644 , n77643 );
buf ( n77645 , n77644 );
buf ( n77646 , n77645 );
xor ( n77647 , n70735 , n70736 );
buf ( n77648 , n77647 );
buf ( n77649 , n77648 );
buf ( n77650 , n77649 );
buf ( n77651 , n77650 );
xor ( n77652 , n70449 , n70450 );
buf ( n77653 , n77652 );
buf ( n77654 , n77653 );
buf ( n77655 , n77654 );
buf ( n77656 , n77655 );
xor ( n77657 , n70157 , n70158 );
buf ( n77658 , n77657 );
buf ( n77659 , n77658 );
buf ( n77660 , n77659 );
buf ( n77661 , n77660 );
xor ( n77662 , n69859 , n69860 );
buf ( n77663 , n77662 );
buf ( n77664 , n77663 );
buf ( n77665 , n77664 );
buf ( n77666 , n77665 );
xor ( n77667 , n69555 , n69556 );
buf ( n77668 , n77667 );
buf ( n77669 , n77668 );
buf ( n77670 , n77669 );
buf ( n77671 , n77670 );
xor ( n77672 , n69245 , n69246 );
buf ( n77673 , n77672 );
buf ( n77674 , n77673 );
buf ( n77675 , n77674 );
buf ( n77676 , n77675 );
xor ( n77677 , n68929 , n68930 );
buf ( n77678 , n77677 );
buf ( n77679 , n77678 );
buf ( n77680 , n77679 );
buf ( n77681 , n77680 );
xor ( n77682 , n68607 , n68608 );
buf ( n77683 , n77682 );
buf ( n77684 , n77683 );
buf ( n77685 , n77684 );
buf ( n77686 , n77685 );
xor ( n77687 , n68279 , n68280 );
buf ( n77688 , n77687 );
buf ( n77689 , n77688 );
buf ( n77690 , n77689 );
buf ( n77691 , n77690 );
xor ( n77692 , n67945 , n67946 );
buf ( n77693 , n77692 );
buf ( n77694 , n77693 );
buf ( n77695 , n77694 );
buf ( n77696 , n77695 );
xor ( n77697 , n67605 , n67606 );
buf ( n77698 , n77697 );
buf ( n77699 , n77698 );
buf ( n77700 , n77699 );
buf ( n77701 , n77700 );
xor ( n77702 , n67259 , n67260 );
buf ( n77703 , n77702 );
buf ( n77704 , n77703 );
buf ( n77705 , n77704 );
buf ( n77706 , n77705 );
xor ( n77707 , n66907 , n66908 );
buf ( n77708 , n77707 );
buf ( n77709 , n77708 );
buf ( n77710 , n77709 );
buf ( n77711 , n77710 );
xor ( n77712 , n66549 , n66550 );
buf ( n77713 , n77712 );
buf ( n77714 , n77713 );
buf ( n77715 , n77714 );
buf ( n77716 , n77715 );
xor ( n77717 , n66185 , n66186 );
buf ( n77718 , n77717 );
buf ( n77719 , n77718 );
buf ( n77720 , n77719 );
buf ( n77721 , n77720 );
xor ( n77722 , n65815 , n65816 );
buf ( n77723 , n77722 );
buf ( n77724 , n77723 );
buf ( n77725 , n77724 );
buf ( n77726 , n77725 );
xor ( n77727 , n65439 , n65440 );
buf ( n77728 , n77727 );
buf ( n77729 , n77728 );
buf ( n77730 , n77729 );
buf ( n77731 , n77730 );
xor ( n77732 , n65057 , n65058 );
buf ( n77733 , n77732 );
buf ( n77734 , n77733 );
buf ( n77735 , n77734 );
buf ( n77736 , n77735 );
xor ( n77737 , n64669 , n64670 );
buf ( n77738 , n77737 );
buf ( n77739 , n77738 );
buf ( n77740 , n77739 );
buf ( n77741 , n77740 );
xor ( n77742 , n64275 , n64276 );
buf ( n77743 , n77742 );
buf ( n77744 , n77743 );
buf ( n77745 , n77744 );
buf ( n77746 , n77745 );
xor ( n77747 , n63875 , n63876 );
buf ( n77748 , n77747 );
buf ( n77749 , n77748 );
buf ( n77750 , n77749 );
buf ( n77751 , n77750 );
xor ( n77752 , n63469 , n63470 );
buf ( n77753 , n77752 );
buf ( n77754 , n77753 );
buf ( n77755 , n77754 );
buf ( n77756 , n77755 );
xor ( n77757 , n63057 , n63058 );
buf ( n77758 , n77757 );
buf ( n77759 , n77758 );
buf ( n77760 , n77759 );
buf ( n77761 , n77760 );
xor ( n77762 , n62639 , n62640 );
buf ( n77763 , n77762 );
buf ( n77764 , n77763 );
buf ( n77765 , n77764 );
buf ( n77766 , n77765 );
xor ( n77767 , n62215 , n62216 );
buf ( n77768 , n77767 );
buf ( n77769 , n77768 );
buf ( n77770 , n77769 );
buf ( n77771 , n77770 );
xor ( n77772 , n61785 , n61786 );
buf ( n77773 , n77772 );
buf ( n77774 , n77773 );
buf ( n77775 , n77774 );
buf ( n77776 , n77775 );
xor ( n77777 , n61349 , n61350 );
buf ( n77778 , n77777 );
buf ( n77779 , n77778 );
buf ( n77780 , n77779 );
buf ( n77781 , n77780 );
xor ( n77782 , n60907 , n60908 );
buf ( n77783 , n77782 );
buf ( n77784 , n77783 );
buf ( n77785 , n77784 );
buf ( n77786 , n77785 );
xor ( n77787 , n60459 , n60460 );
buf ( n77788 , n77787 );
buf ( n77789 , n77788 );
buf ( n77790 , n77789 );
buf ( n77791 , n77790 );
xor ( n77792 , n60005 , n60006 );
buf ( n77793 , n77792 );
buf ( n77794 , n77793 );
buf ( n77795 , n77794 );
buf ( n77796 , n77795 );
xor ( n77797 , n59545 , n59546 );
buf ( n77798 , n77797 );
buf ( n77799 , n77798 );
buf ( n77800 , n77799 );
buf ( n77801 , n77800 );
xor ( n77802 , n59079 , n59080 );
buf ( n77803 , n77802 );
buf ( n77804 , n77803 );
buf ( n77805 , n77804 );
buf ( n77806 , n77805 );
xor ( n77807 , n58607 , n58608 );
buf ( n77808 , n77807 );
buf ( n77809 , n77808 );
buf ( n77810 , n77809 );
buf ( n77811 , n77810 );
xor ( n77812 , n58129 , n58130 );
buf ( n77813 , n77812 );
buf ( n77814 , n77813 );
buf ( n77815 , n77814 );
buf ( n77816 , n77815 );
xor ( n77817 , n57645 , n57646 );
buf ( n77818 , n77817 );
buf ( n77819 , n77818 );
buf ( n77820 , n77819 );
buf ( n77821 , n77820 );
xor ( n77822 , n57155 , n57156 );
buf ( n77823 , n77822 );
buf ( n77824 , n77823 );
buf ( n77825 , n77824 );
buf ( n77826 , n77825 );
xor ( n77827 , n56659 , n56660 );
buf ( n77828 , n77827 );
buf ( n77829 , n77828 );
buf ( n77830 , n77829 );
buf ( n77831 , n77830 );
xor ( n77832 , n56157 , n56158 );
buf ( n77833 , n77832 );
buf ( n77834 , n77833 );
buf ( n77835 , n77834 );
buf ( n77836 , n77835 );
xor ( n77837 , n55649 , n55650 );
buf ( n77838 , n77837 );
buf ( n77839 , n77838 );
buf ( n77840 , n77839 );
buf ( n77841 , n77840 );
xor ( n77842 , n55135 , n55136 );
buf ( n77843 , n77842 );
buf ( n77844 , n77843 );
buf ( n77845 , n77844 );
buf ( n77846 , n77845 );
xor ( n77847 , n54615 , n54616 );
buf ( n77848 , n77847 );
buf ( n77849 , n77848 );
buf ( n77850 , n77849 );
buf ( n77851 , n77850 );
xor ( n77852 , n54089 , n54090 );
buf ( n77853 , n77852 );
buf ( n77854 , n77853 );
buf ( n77855 , n77854 );
buf ( n77856 , n77855 );
xor ( n77857 , n53557 , n53558 );
buf ( n77858 , n77857 );
buf ( n77859 , n77858 );
buf ( n77860 , n77859 );
buf ( n77861 , n77860 );
xor ( n77862 , n53019 , n53020 );
buf ( n77863 , n77862 );
buf ( n77864 , n77863 );
buf ( n77865 , n77864 );
buf ( n77866 , n77865 );
xor ( n77867 , n52475 , n52476 );
buf ( n77868 , n77867 );
buf ( n77869 , n77868 );
buf ( n77870 , n77869 );
buf ( n77871 , n77870 );
xor ( n77872 , n51925 , n51926 );
buf ( n77873 , n77872 );
buf ( n77874 , n77873 );
buf ( n77875 , n77874 );
buf ( n77876 , n77875 );
xor ( n77877 , n51369 , n51370 );
buf ( n77878 , n77877 );
buf ( n77879 , n77878 );
buf ( n77880 , n77879 );
buf ( n77881 , n77880 );
xor ( n77882 , n50807 , n50808 );
buf ( n77883 , n77882 );
buf ( n77884 , n77883 );
buf ( n77885 , n77884 );
buf ( n77886 , n77885 );
xor ( n77887 , n50239 , n50240 );
buf ( n77888 , n77887 );
buf ( n77889 , n77888 );
buf ( n77890 , n77889 );
buf ( n77891 , n77890 );
xor ( n77892 , n49665 , n49666 );
buf ( n77893 , n77892 );
buf ( n77894 , n77893 );
buf ( n77895 , n77894 );
buf ( n77896 , n77895 );
xor ( n77897 , n49085 , n49086 );
buf ( n77898 , n77897 );
buf ( n77899 , n77898 );
buf ( n77900 , n77899 );
buf ( n77901 , n77900 );
xor ( n77902 , n48499 , n48500 );
buf ( n77903 , n77902 );
buf ( n77904 , n77903 );
buf ( n77905 , n77904 );
buf ( n77906 , n77905 );
xor ( n77907 , n47907 , n47908 );
buf ( n77908 , n77907 );
buf ( n77909 , n77908 );
buf ( n77910 , n77909 );
buf ( n77911 , n77910 );
xor ( n77912 , n47309 , n47310 );
buf ( n77913 , n77912 );
buf ( n77914 , n77913 );
buf ( n77915 , n77914 );
buf ( n77916 , n77915 );
xor ( n77917 , n46705 , n46706 );
buf ( n77918 , n77917 );
buf ( n77919 , n77918 );
buf ( n77920 , n77919 );
buf ( n77921 , n77920 );
xor ( n77922 , n46095 , n46096 );
buf ( n77923 , n77922 );
buf ( n77924 , n77923 );
buf ( n77925 , n77924 );
buf ( n77926 , n77925 );
xor ( n77927 , n45479 , n45480 );
buf ( n77928 , n77927 );
buf ( n77929 , n77928 );
buf ( n77930 , n77929 );
buf ( n77931 , n77930 );
xor ( n77932 , n44857 , n44858 );
buf ( n77933 , n77932 );
buf ( n77934 , n77933 );
buf ( n77935 , n77934 );
buf ( n77936 , n77935 );
xor ( n77937 , n44229 , n44230 );
buf ( n77938 , n77937 );
buf ( n77939 , n77938 );
buf ( n77940 , n77939 );
buf ( n77941 , n77940 );
xor ( n77942 , n43595 , n43596 );
buf ( n77943 , n77942 );
buf ( n77944 , n77943 );
buf ( n77945 , n77944 );
buf ( n77946 , n77945 );
xor ( n77947 , n42955 , n42956 );
buf ( n77948 , n77947 );
buf ( n77949 , n77948 );
buf ( n77950 , n77949 );
buf ( n77951 , n77950 );
xor ( n77952 , n42309 , n42310 );
buf ( n77953 , n77952 );
buf ( n77954 , n77953 );
buf ( n77955 , n77954 );
buf ( n77956 , n77955 );
xor ( n77957 , n41657 , n41658 );
buf ( n77958 , n77957 );
buf ( n77959 , n77958 );
buf ( n77960 , n77959 );
buf ( n77961 , n77960 );
xor ( n77962 , n40999 , n41000 );
buf ( n77963 , n77962 );
buf ( n77964 , n77963 );
buf ( n77965 , n77964 );
buf ( n77966 , n77965 );
xor ( n77967 , n40335 , n40336 );
buf ( n77968 , n77967 );
buf ( n77969 , n77968 );
buf ( n77970 , n77969 );
buf ( n77971 , n77970 );
xor ( n77972 , n39665 , n39666 );
buf ( n77973 , n77972 );
buf ( n77974 , n77973 );
buf ( n77975 , n77974 );
buf ( n77976 , n77975 );
xor ( n77977 , n38989 , n38990 );
buf ( n77978 , n77977 );
buf ( n77979 , n77978 );
buf ( n77980 , n77979 );
buf ( n77981 , n77980 );
xor ( n77982 , n38307 , n38308 );
buf ( n77983 , n77982 );
buf ( n77984 , n77983 );
buf ( n77985 , n77984 );
buf ( n77986 , n77985 );
xor ( n77987 , n37619 , n37620 );
buf ( n77988 , n77987 );
buf ( n77989 , n77988 );
buf ( n77990 , n77989 );
buf ( n77991 , n77990 );
xor ( n77992 , n36925 , n36926 );
buf ( n77993 , n77992 );
buf ( n77994 , n77993 );
buf ( n77995 , n77994 );
buf ( n77996 , n77995 );
xor ( n77997 , n36225 , n36226 );
buf ( n77998 , n77997 );
buf ( n77999 , n77998 );
buf ( n78000 , n77999 );
buf ( n78001 , n78000 );
xor ( n78002 , n35519 , n35520 );
buf ( n78003 , n78002 );
buf ( n78004 , n78003 );
buf ( n78005 , n78004 );
buf ( n78006 , n78005 );
xor ( n78007 , n34807 , n34808 );
buf ( n78008 , n78007 );
buf ( n78009 , n78008 );
buf ( n78010 , n78009 );
buf ( n78011 , n78010 );
xor ( n78012 , n34089 , n34090 );
buf ( n78013 , n78012 );
buf ( n78014 , n78013 );
buf ( n78015 , n78014 );
buf ( n78016 , n78015 );
xor ( n78017 , n33365 , n33366 );
buf ( n78018 , n78017 );
buf ( n78019 , n78018 );
buf ( n78020 , n78019 );
buf ( n78021 , n78020 );
xor ( n78022 , n32635 , n32636 );
buf ( n78023 , n78022 );
buf ( n78024 , n78023 );
buf ( n78025 , n78024 );
buf ( n78026 , n78025 );
xor ( n78027 , n31899 , n31900 );
buf ( n78028 , n78027 );
buf ( n78029 , n78028 );
buf ( n78030 , n78029 );
buf ( n78031 , n78030 );
xor ( n78032 , n31157 , n31158 );
buf ( n78033 , n78032 );
buf ( n78034 , n78033 );
buf ( n78035 , n78034 );
buf ( n78036 , n78035 );
xor ( n78037 , n30408 , n30410 );
buf ( n78038 , n78037 );
buf ( n78039 , n78038 );
buf ( n78040 , n78039 );
buf ( n78041 , n78040 );
and ( n78042 , n30409 , n29782 );
buf ( n78043 , n78042 );
buf ( n78044 , n78043 );
buf ( n78045 , n78044 );
buf ( n78046 , n608 );
buf ( n78047 , n78046 );
buf ( n78048 , n78047 );
buf ( n78049 , n609 );
buf ( n78050 , n78049 );
buf ( n78051 , n608 );
buf ( n78052 , n78051 );
and ( n78053 , n78050 , n78052 );
buf ( n78054 , n609 );
buf ( n78055 , n78054 );
and ( n78056 , n78047 , n78055 );
and ( n78057 , n78053 , n78056 );
buf ( n78058 , n610 );
buf ( n78059 , n78058 );
and ( n78060 , n78047 , n78059 );
buf ( n78061 , n610 );
buf ( n78062 , n78061 );
and ( n78063 , n78062 , n78052 );
and ( n78064 , n78060 , n78063 );
and ( n78065 , n78056 , n78064 );
and ( n78066 , n78053 , n78064 );
or ( n78067 , n78057 , n78065 , n78066 );
and ( n78068 , n78048 , n78067 );
buf ( n78069 , n611 );
buf ( n78070 , n78069 );
and ( n78071 , n78070 , n78052 );
and ( n78072 , n78062 , n78055 );
or ( n78073 , n78071 , n78072 );
buf ( n78074 , n611 );
buf ( n78075 , n78074 );
and ( n78076 , n78047 , n78075 );
and ( n78077 , n78050 , n78059 );
or ( n78078 , n78076 , n78077 );
and ( n78079 , n78073 , n78078 );
xor ( n78080 , n78053 , n78056 );
xor ( n78081 , n78080 , n78064 );
and ( n78082 , n78079 , n78081 );
xnor ( n78083 , n78071 , n78072 );
xnor ( n78084 , n78076 , n78077 );
and ( n78085 , n78083 , n78084 );
buf ( n78086 , n78050 );
or ( n78087 , n78085 , n78086 );
and ( n78088 , n78081 , n78087 );
and ( n78089 , n78079 , n78087 );
or ( n78090 , n78082 , n78088 , n78089 );
and ( n78091 , n78067 , n78090 );
and ( n78092 , n78048 , n78090 );
or ( n78093 , n78068 , n78091 , n78092 );
xor ( n78094 , n78060 , n78063 );
xor ( n78095 , n78073 , n78078 );
and ( n78096 , n78094 , n78095 );
buf ( n78097 , n612 );
buf ( n78098 , n78097 );
and ( n78099 , n78098 , n78052 );
and ( n78100 , n78070 , n78055 );
or ( n78101 , n78099 , n78100 );
buf ( n78102 , n612 );
buf ( n78103 , n78102 );
and ( n78104 , n78047 , n78103 );
and ( n78105 , n78050 , n78075 );
or ( n78106 , n78104 , n78105 );
and ( n78107 , n78101 , n78106 );
and ( n78108 , n78095 , n78107 );
and ( n78109 , n78094 , n78107 );
or ( n78110 , n78096 , n78108 , n78109 );
xnor ( n78111 , n78085 , n78086 );
xor ( n78112 , n78101 , n78106 );
xor ( n78113 , n78083 , n78084 );
and ( n78114 , n78112 , n78113 );
buf ( n78115 , n613 );
buf ( n78116 , n78115 );
and ( n78117 , n78116 , n78052 );
and ( n78118 , n78070 , n78059 );
or ( n78119 , n78117 , n78118 );
buf ( n78120 , n613 );
buf ( n78121 , n78120 );
and ( n78122 , n78047 , n78121 );
and ( n78123 , n78062 , n78075 );
or ( n78124 , n78122 , n78123 );
and ( n78125 , n78119 , n78124 );
and ( n78126 , n78113 , n78125 );
and ( n78127 , n78112 , n78125 );
or ( n78128 , n78114 , n78126 , n78127 );
and ( n78129 , n78111 , n78128 );
xor ( n78130 , n78094 , n78095 );
xor ( n78131 , n78130 , n78107 );
and ( n78132 , n78128 , n78131 );
and ( n78133 , n78111 , n78131 );
or ( n78134 , n78129 , n78132 , n78133 );
and ( n78135 , n78110 , n78134 );
xor ( n78136 , n78079 , n78081 );
xor ( n78137 , n78136 , n78087 );
and ( n78138 , n78134 , n78137 );
and ( n78139 , n78110 , n78137 );
or ( n78140 , n78135 , n78138 , n78139 );
xor ( n78141 , n78048 , n78067 );
xor ( n78142 , n78141 , n78090 );
and ( n78143 , n78140 , n78142 );
xor ( n78144 , n78110 , n78134 );
xor ( n78145 , n78144 , n78137 );
xnor ( n78146 , n78099 , n78100 );
xnor ( n78147 , n78104 , n78105 );
and ( n78148 , n78146 , n78147 );
xnor ( n78149 , n78117 , n78118 );
xnor ( n78150 , n78122 , n78123 );
and ( n78151 , n78149 , n78150 );
buf ( n78152 , n78062 );
or ( n78153 , n78151 , n78152 );
and ( n78154 , n78148 , n78153 );
buf ( n78155 , n614 );
buf ( n78156 , n78155 );
and ( n78157 , n78047 , n78156 );
and ( n78158 , n78050 , n78121 );
and ( n78159 , n78157 , n78158 );
and ( n78160 , n78062 , n78103 );
and ( n78161 , n78158 , n78160 );
and ( n78162 , n78157 , n78160 );
or ( n78163 , n78159 , n78161 , n78162 );
and ( n78164 , n78098 , n78055 );
or ( n78165 , n78163 , n78164 );
buf ( n78166 , n614 );
buf ( n78167 , n78166 );
and ( n78168 , n78167 , n78052 );
and ( n78169 , n78116 , n78055 );
and ( n78170 , n78168 , n78169 );
and ( n78171 , n78098 , n78059 );
and ( n78172 , n78169 , n78171 );
and ( n78173 , n78168 , n78171 );
or ( n78174 , n78170 , n78172 , n78173 );
and ( n78175 , n78050 , n78103 );
or ( n78176 , n78174 , n78175 );
and ( n78177 , n78165 , n78176 );
and ( n78178 , n78153 , n78177 );
and ( n78179 , n78148 , n78177 );
or ( n78180 , n78154 , n78178 , n78179 );
xor ( n78181 , n78111 , n78128 );
xor ( n78182 , n78181 , n78131 );
and ( n78183 , n78180 , n78182 );
xor ( n78184 , n78112 , n78113 );
xor ( n78185 , n78184 , n78125 );
xnor ( n78186 , n78163 , n78164 );
xnor ( n78187 , n78174 , n78175 );
and ( n78188 , n78186 , n78187 );
xnor ( n78189 , n78151 , n78152 );
or ( n78190 , n78188 , n78189 );
and ( n78191 , n78185 , n78190 );
xor ( n78192 , n78119 , n78124 );
xor ( n78193 , n78146 , n78147 );
and ( n78194 , n78192 , n78193 );
xor ( n78195 , n78165 , n78176 );
and ( n78196 , n78193 , n78195 );
and ( n78197 , n78192 , n78195 );
or ( n78198 , n78194 , n78196 , n78197 );
and ( n78199 , n78190 , n78198 );
and ( n78200 , n78185 , n78198 );
or ( n78201 , n78191 , n78199 , n78200 );
and ( n78202 , n78182 , n78201 );
and ( n78203 , n78180 , n78201 );
or ( n78204 , n78183 , n78202 , n78203 );
and ( n78205 , n78145 , n78204 );
xor ( n78206 , n78148 , n78153 );
xor ( n78207 , n78206 , n78177 );
xor ( n78208 , n78149 , n78150 );
and ( n78209 , n78167 , n78055 );
and ( n78210 , n78098 , n78075 );
or ( n78211 , n78209 , n78210 );
and ( n78212 , n78050 , n78156 );
and ( n78213 , n78070 , n78103 );
or ( n78214 , n78212 , n78213 );
and ( n78215 , n78211 , n78214 );
and ( n78216 , n78208 , n78215 );
xor ( n78217 , n78168 , n78169 );
xor ( n78218 , n78217 , n78171 );
xor ( n78219 , n78157 , n78158 );
xor ( n78220 , n78219 , n78160 );
and ( n78221 , n78218 , n78220 );
and ( n78222 , n78215 , n78221 );
and ( n78223 , n78208 , n78221 );
or ( n78224 , n78216 , n78222 , n78223 );
xnor ( n78225 , n78188 , n78189 );
and ( n78226 , n78224 , n78225 );
xor ( n78227 , n78186 , n78187 );
xnor ( n78228 , n78209 , n78210 );
xnor ( n78229 , n78212 , n78213 );
and ( n78230 , n78228 , n78229 );
buf ( n78231 , n78070 );
or ( n78232 , n78230 , n78231 );
and ( n78233 , n78227 , n78232 );
buf ( n78234 , n616 );
buf ( n78235 , n78234 );
and ( n78236 , n78047 , n78235 );
and ( n78237 , n78062 , n78156 );
and ( n78238 , n78236 , n78237 );
and ( n78239 , n78070 , n78121 );
and ( n78240 , n78237 , n78239 );
and ( n78241 , n78236 , n78239 );
or ( n78242 , n78238 , n78240 , n78241 );
buf ( n78243 , n615 );
buf ( n78244 , n78243 );
and ( n78245 , n78244 , n78052 );
and ( n78246 , n78242 , n78245 );
and ( n78247 , n78116 , n78059 );
and ( n78248 , n78245 , n78247 );
and ( n78249 , n78242 , n78247 );
or ( n78250 , n78246 , n78248 , n78249 );
buf ( n78251 , n616 );
buf ( n78252 , n78251 );
and ( n78253 , n78252 , n78052 );
and ( n78254 , n78167 , n78059 );
and ( n78255 , n78253 , n78254 );
and ( n78256 , n78116 , n78075 );
and ( n78257 , n78254 , n78256 );
and ( n78258 , n78253 , n78256 );
or ( n78259 , n78255 , n78257 , n78258 );
buf ( n78260 , n615 );
buf ( n78261 , n78260 );
and ( n78262 , n78047 , n78261 );
and ( n78263 , n78259 , n78262 );
and ( n78264 , n78062 , n78121 );
and ( n78265 , n78262 , n78264 );
and ( n78266 , n78259 , n78264 );
or ( n78267 , n78263 , n78265 , n78266 );
and ( n78268 , n78250 , n78267 );
and ( n78269 , n78232 , n78268 );
and ( n78270 , n78227 , n78268 );
or ( n78271 , n78233 , n78269 , n78270 );
and ( n78272 , n78225 , n78271 );
and ( n78273 , n78224 , n78271 );
or ( n78274 , n78226 , n78272 , n78273 );
and ( n78275 , n78207 , n78274 );
xor ( n78276 , n78185 , n78190 );
xor ( n78277 , n78276 , n78198 );
and ( n78278 , n78274 , n78277 );
and ( n78279 , n78207 , n78277 );
or ( n78280 , n78275 , n78278 , n78279 );
xor ( n78281 , n78180 , n78182 );
xor ( n78282 , n78281 , n78201 );
and ( n78283 , n78280 , n78282 );
xor ( n78284 , n78192 , n78193 );
xor ( n78285 , n78284 , n78195 );
xor ( n78286 , n78208 , n78215 );
xor ( n78287 , n78286 , n78221 );
xor ( n78288 , n78211 , n78214 );
xor ( n78289 , n78218 , n78220 );
and ( n78290 , n78288 , n78289 );
xnor ( n78291 , n78230 , n78231 );
and ( n78292 , n78289 , n78291 );
and ( n78293 , n78288 , n78291 );
or ( n78294 , n78290 , n78292 , n78293 );
and ( n78295 , n78287 , n78294 );
xor ( n78296 , n78250 , n78267 );
xor ( n78297 , n78242 , n78245 );
xor ( n78298 , n78297 , n78247 );
xor ( n78299 , n78259 , n78262 );
xor ( n78300 , n78299 , n78264 );
and ( n78301 , n78298 , n78300 );
and ( n78302 , n78296 , n78301 );
and ( n78303 , n78050 , n78261 );
and ( n78304 , n78244 , n78055 );
and ( n78305 , n78303 , n78304 );
xor ( n78306 , n78228 , n78229 );
and ( n78307 , n78305 , n78306 );
and ( n78308 , n78098 , n78121 );
and ( n78309 , n78116 , n78103 );
and ( n78310 , n78308 , n78309 );
not ( n78311 , n78310 );
buf ( n78312 , n78098 );
and ( n78313 , n78311 , n78312 );
and ( n78314 , n78306 , n78313 );
and ( n78315 , n78305 , n78313 );
or ( n78316 , n78307 , n78314 , n78315 );
and ( n78317 , n78301 , n78316 );
and ( n78318 , n78296 , n78316 );
or ( n78319 , n78302 , n78317 , n78318 );
and ( n78320 , n78294 , n78319 );
and ( n78321 , n78287 , n78319 );
or ( n78322 , n78295 , n78320 , n78321 );
and ( n78323 , n78285 , n78322 );
xor ( n78324 , n78224 , n78225 );
xor ( n78325 , n78324 , n78271 );
and ( n78326 , n78322 , n78325 );
and ( n78327 , n78285 , n78325 );
or ( n78328 , n78323 , n78326 , n78327 );
xor ( n78329 , n78207 , n78274 );
xor ( n78330 , n78329 , n78277 );
and ( n78331 , n78328 , n78330 );
xor ( n78332 , n78227 , n78232 );
xor ( n78333 , n78332 , n78268 );
buf ( n78334 , n78310 );
buf ( n78335 , n617 );
buf ( n78336 , n78335 );
and ( n78337 , n78336 , n78052 );
and ( n78338 , n78252 , n78055 );
and ( n78339 , n78337 , n78338 );
and ( n78340 , n78167 , n78075 );
and ( n78341 , n78338 , n78340 );
and ( n78342 , n78337 , n78340 );
or ( n78343 , n78339 , n78341 , n78342 );
buf ( n78344 , n617 );
buf ( n78345 , n78344 );
and ( n78346 , n78047 , n78345 );
and ( n78347 , n78050 , n78235 );
and ( n78348 , n78346 , n78347 );
and ( n78349 , n78070 , n78156 );
and ( n78350 , n78347 , n78349 );
and ( n78351 , n78346 , n78349 );
or ( n78352 , n78348 , n78350 , n78351 );
and ( n78353 , n78343 , n78352 );
and ( n78354 , n78334 , n78353 );
xor ( n78355 , n78253 , n78254 );
xor ( n78356 , n78355 , n78256 );
xor ( n78357 , n78236 , n78237 );
xor ( n78358 , n78357 , n78239 );
and ( n78359 , n78356 , n78358 );
and ( n78360 , n78353 , n78359 );
and ( n78361 , n78334 , n78359 );
or ( n78362 , n78354 , n78360 , n78361 );
xor ( n78363 , n78298 , n78300 );
and ( n78364 , n78062 , n78261 );
and ( n78365 , n78244 , n78059 );
and ( n78366 , n78364 , n78365 );
xor ( n78367 , n78311 , n78312 );
or ( n78368 , n78366 , n78367 );
and ( n78369 , n78363 , n78368 );
xor ( n78370 , n78303 , n78304 );
xor ( n78371 , n78343 , n78352 );
and ( n78372 , n78370 , n78371 );
xor ( n78373 , n78356 , n78358 );
and ( n78374 , n78371 , n78373 );
and ( n78375 , n78370 , n78373 );
or ( n78376 , n78372 , n78374 , n78375 );
and ( n78377 , n78368 , n78376 );
and ( n78378 , n78363 , n78376 );
or ( n78379 , n78369 , n78377 , n78378 );
and ( n78380 , n78362 , n78379 );
xor ( n78381 , n78288 , n78289 );
xor ( n78382 , n78381 , n78291 );
and ( n78383 , n78379 , n78382 );
and ( n78384 , n78362 , n78382 );
or ( n78385 , n78380 , n78383 , n78384 );
and ( n78386 , n78333 , n78385 );
xor ( n78387 , n78287 , n78294 );
xor ( n78388 , n78387 , n78319 );
and ( n78389 , n78385 , n78388 );
and ( n78390 , n78333 , n78388 );
or ( n78391 , n78386 , n78389 , n78390 );
xor ( n78392 , n78285 , n78322 );
xor ( n78393 , n78392 , n78325 );
and ( n78394 , n78391 , n78393 );
xor ( n78395 , n78296 , n78301 );
xor ( n78396 , n78395 , n78316 );
xor ( n78397 , n78305 , n78306 );
xor ( n78398 , n78397 , n78313 );
xor ( n78399 , n78334 , n78353 );
xor ( n78400 , n78399 , n78359 );
and ( n78401 , n78398 , n78400 );
xnor ( n78402 , n78366 , n78367 );
and ( n78403 , n78336 , n78055 );
and ( n78404 , n78244 , n78075 );
and ( n78405 , n78403 , n78404 );
and ( n78406 , n78167 , n78103 );
and ( n78407 , n78404 , n78406 );
and ( n78408 , n78403 , n78406 );
or ( n78409 , n78405 , n78407 , n78408 );
and ( n78410 , n78050 , n78345 );
and ( n78411 , n78070 , n78261 );
and ( n78412 , n78410 , n78411 );
and ( n78413 , n78098 , n78156 );
and ( n78414 , n78411 , n78413 );
and ( n78415 , n78410 , n78413 );
or ( n78416 , n78412 , n78414 , n78415 );
and ( n78417 , n78409 , n78416 );
and ( n78418 , n78402 , n78417 );
xor ( n78419 , n78337 , n78338 );
xor ( n78420 , n78419 , n78340 );
xor ( n78421 , n78346 , n78347 );
xor ( n78422 , n78421 , n78349 );
and ( n78423 , n78420 , n78422 );
and ( n78424 , n78417 , n78423 );
and ( n78425 , n78402 , n78423 );
or ( n78426 , n78418 , n78424 , n78425 );
and ( n78427 , n78400 , n78426 );
and ( n78428 , n78398 , n78426 );
or ( n78429 , n78401 , n78427 , n78428 );
and ( n78430 , n78396 , n78429 );
xor ( n78431 , n78362 , n78379 );
xor ( n78432 , n78431 , n78382 );
and ( n78433 , n78429 , n78432 );
and ( n78434 , n78396 , n78432 );
or ( n78435 , n78430 , n78433 , n78434 );
xor ( n78436 , n78333 , n78385 );
xor ( n78437 , n78436 , n78388 );
and ( n78438 , n78435 , n78437 );
buf ( n78439 , n618 );
buf ( n78440 , n78439 );
and ( n78441 , n78050 , n78440 );
and ( n78442 , n78062 , n78345 );
and ( n78443 , n78441 , n78442 );
and ( n78444 , n78098 , n78261 );
and ( n78445 , n78442 , n78444 );
and ( n78446 , n78441 , n78444 );
or ( n78447 , n78443 , n78445 , n78446 );
buf ( n78448 , n618 );
buf ( n78449 , n78448 );
and ( n78450 , n78449 , n78052 );
and ( n78451 , n78447 , n78450 );
and ( n78452 , n78252 , n78059 );
and ( n78453 , n78450 , n78452 );
and ( n78454 , n78447 , n78452 );
or ( n78455 , n78451 , n78453 , n78454 );
and ( n78456 , n78449 , n78055 );
and ( n78457 , n78336 , n78059 );
and ( n78458 , n78456 , n78457 );
and ( n78459 , n78244 , n78103 );
and ( n78460 , n78457 , n78459 );
and ( n78461 , n78456 , n78459 );
or ( n78462 , n78458 , n78460 , n78461 );
and ( n78463 , n78047 , n78440 );
and ( n78464 , n78462 , n78463 );
and ( n78465 , n78062 , n78235 );
and ( n78466 , n78463 , n78465 );
and ( n78467 , n78462 , n78465 );
or ( n78468 , n78464 , n78466 , n78467 );
and ( n78469 , n78455 , n78468 );
xor ( n78470 , n78364 , n78365 );
xor ( n78471 , n78308 , n78309 );
and ( n78472 , n78470 , n78471 );
xor ( n78473 , n78409 , n78416 );
and ( n78474 , n78471 , n78473 );
and ( n78475 , n78470 , n78473 );
or ( n78476 , n78472 , n78474 , n78475 );
and ( n78477 , n78469 , n78476 );
xor ( n78478 , n78420 , n78422 );
and ( n78479 , n78116 , n78156 );
and ( n78480 , n78167 , n78121 );
and ( n78481 , n78479 , n78480 );
not ( n78482 , n78481 );
buf ( n78483 , n78116 );
and ( n78484 , n78482 , n78483 );
and ( n78485 , n78478 , n78484 );
buf ( n78486 , n78481 );
and ( n78487 , n78484 , n78486 );
and ( n78488 , n78478 , n78486 );
or ( n78489 , n78485 , n78487 , n78488 );
and ( n78490 , n78476 , n78489 );
and ( n78491 , n78469 , n78489 );
or ( n78492 , n78477 , n78490 , n78491 );
xor ( n78493 , n78363 , n78368 );
xor ( n78494 , n78493 , n78376 );
and ( n78495 , n78492 , n78494 );
xor ( n78496 , n78370 , n78371 );
xor ( n78497 , n78496 , n78373 );
xor ( n78498 , n78402 , n78417 );
xor ( n78499 , n78498 , n78423 );
and ( n78500 , n78497 , n78499 );
xor ( n78501 , n78403 , n78404 );
xor ( n78502 , n78501 , n78406 );
xor ( n78503 , n78410 , n78411 );
xor ( n78504 , n78503 , n78413 );
and ( n78505 , n78502 , n78504 );
xor ( n78506 , n78455 , n78468 );
and ( n78507 , n78505 , n78506 );
and ( n78508 , n78062 , n78440 );
and ( n78509 , n78098 , n78235 );
and ( n78510 , n78508 , n78509 );
and ( n78511 , n78116 , n78261 );
and ( n78512 , n78509 , n78511 );
and ( n78513 , n78508 , n78511 );
or ( n78514 , n78510 , n78512 , n78513 );
buf ( n78515 , n620 );
buf ( n78516 , n78515 );
and ( n78517 , n78047 , n78516 );
buf ( n78518 , n619 );
buf ( n78519 , n78518 );
and ( n78520 , n78050 , n78519 );
and ( n78521 , n78517 , n78520 );
and ( n78522 , n78070 , n78345 );
and ( n78523 , n78520 , n78522 );
and ( n78524 , n78517 , n78522 );
or ( n78525 , n78521 , n78523 , n78524 );
and ( n78526 , n78514 , n78525 );
buf ( n78527 , n619 );
buf ( n78528 , n78527 );
and ( n78529 , n78528 , n78052 );
and ( n78530 , n78525 , n78529 );
and ( n78531 , n78514 , n78529 );
or ( n78532 , n78526 , n78530 , n78531 );
and ( n78533 , n78449 , n78059 );
and ( n78534 , n78252 , n78103 );
and ( n78535 , n78533 , n78534 );
and ( n78536 , n78244 , n78121 );
and ( n78537 , n78534 , n78536 );
and ( n78538 , n78533 , n78536 );
or ( n78539 , n78535 , n78537 , n78538 );
buf ( n78540 , n620 );
buf ( n78541 , n78540 );
and ( n78542 , n78541 , n78052 );
and ( n78543 , n78528 , n78055 );
and ( n78544 , n78542 , n78543 );
and ( n78545 , n78336 , n78075 );
and ( n78546 , n78543 , n78545 );
and ( n78547 , n78542 , n78545 );
or ( n78548 , n78544 , n78546 , n78547 );
and ( n78549 , n78539 , n78548 );
and ( n78550 , n78047 , n78519 );
and ( n78551 , n78548 , n78550 );
and ( n78552 , n78539 , n78550 );
or ( n78553 , n78549 , n78551 , n78552 );
and ( n78554 , n78532 , n78553 );
and ( n78555 , n78506 , n78554 );
and ( n78556 , n78505 , n78554 );
or ( n78557 , n78507 , n78555 , n78556 );
and ( n78558 , n78499 , n78557 );
and ( n78559 , n78497 , n78557 );
or ( n78560 , n78500 , n78558 , n78559 );
and ( n78561 , n78494 , n78560 );
and ( n78562 , n78492 , n78560 );
or ( n78563 , n78495 , n78561 , n78562 );
xor ( n78564 , n78396 , n78429 );
xor ( n78565 , n78564 , n78432 );
and ( n78566 , n78563 , n78565 );
xor ( n78567 , n78398 , n78400 );
xor ( n78568 , n78567 , n78426 );
xor ( n78569 , n78447 , n78450 );
xor ( n78570 , n78569 , n78452 );
xor ( n78571 , n78462 , n78463 );
xor ( n78572 , n78571 , n78465 );
and ( n78573 , n78570 , n78572 );
and ( n78574 , n78070 , n78235 );
and ( n78575 , n78252 , n78075 );
and ( n78576 , n78574 , n78575 );
xor ( n78577 , n78482 , n78483 );
and ( n78578 , n78576 , n78577 );
xor ( n78579 , n78502 , n78504 );
and ( n78580 , n78577 , n78579 );
and ( n78581 , n78576 , n78579 );
or ( n78582 , n78578 , n78580 , n78581 );
and ( n78583 , n78573 , n78582 );
xor ( n78584 , n78470 , n78471 );
xor ( n78585 , n78584 , n78473 );
and ( n78586 , n78582 , n78585 );
and ( n78587 , n78573 , n78585 );
or ( n78588 , n78583 , n78586 , n78587 );
xor ( n78589 , n78469 , n78476 );
xor ( n78590 , n78589 , n78489 );
and ( n78591 , n78588 , n78590 );
xor ( n78592 , n78478 , n78484 );
xor ( n78593 , n78592 , n78486 );
xor ( n78594 , n78456 , n78457 );
xor ( n78595 , n78594 , n78459 );
xor ( n78596 , n78441 , n78442 );
xor ( n78597 , n78596 , n78444 );
and ( n78598 , n78595 , n78597 );
xor ( n78599 , n78532 , n78553 );
and ( n78600 , n78598 , n78599 );
xor ( n78601 , n78570 , n78572 );
and ( n78602 , n78599 , n78601 );
and ( n78603 , n78598 , n78601 );
or ( n78604 , n78600 , n78602 , n78603 );
and ( n78605 , n78593 , n78604 );
xor ( n78606 , n78514 , n78525 );
xor ( n78607 , n78606 , n78529 );
xor ( n78608 , n78539 , n78548 );
xor ( n78609 , n78608 , n78550 );
and ( n78610 , n78607 , n78609 );
xor ( n78611 , n78574 , n78575 );
xor ( n78612 , n78479 , n78480 );
and ( n78613 , n78611 , n78612 );
xor ( n78614 , n78595 , n78597 );
and ( n78615 , n78612 , n78614 );
and ( n78616 , n78611 , n78614 );
or ( n78617 , n78613 , n78615 , n78616 );
and ( n78618 , n78610 , n78617 );
buf ( n78619 , n621 );
buf ( n78620 , n78619 );
and ( n78621 , n78620 , n78052 );
and ( n78622 , n78449 , n78075 );
and ( n78623 , n78621 , n78622 );
and ( n78624 , n78252 , n78121 );
and ( n78625 , n78622 , n78624 );
and ( n78626 , n78621 , n78624 );
or ( n78627 , n78623 , n78625 , n78626 );
buf ( n78628 , n621 );
buf ( n78629 , n78628 );
and ( n78630 , n78047 , n78629 );
and ( n78631 , n78070 , n78440 );
and ( n78632 , n78630 , n78631 );
and ( n78633 , n78116 , n78235 );
and ( n78634 , n78631 , n78633 );
and ( n78635 , n78630 , n78633 );
or ( n78636 , n78632 , n78634 , n78635 );
and ( n78637 , n78627 , n78636 );
and ( n78638 , n78336 , n78103 );
and ( n78639 , n78244 , n78156 );
or ( n78640 , n78638 , n78639 );
and ( n78641 , n78098 , n78345 );
and ( n78642 , n78167 , n78261 );
or ( n78643 , n78641 , n78642 );
and ( n78644 , n78640 , n78643 );
and ( n78645 , n78637 , n78644 );
xor ( n78646 , n78533 , n78534 );
xor ( n78647 , n78646 , n78536 );
xor ( n78648 , n78508 , n78509 );
xor ( n78649 , n78648 , n78511 );
and ( n78650 , n78647 , n78649 );
and ( n78651 , n78644 , n78650 );
and ( n78652 , n78637 , n78650 );
or ( n78653 , n78645 , n78651 , n78652 );
and ( n78654 , n78617 , n78653 );
and ( n78655 , n78610 , n78653 );
or ( n78656 , n78618 , n78654 , n78655 );
and ( n78657 , n78604 , n78656 );
and ( n78658 , n78593 , n78656 );
or ( n78659 , n78605 , n78657 , n78658 );
and ( n78660 , n78590 , n78659 );
and ( n78661 , n78588 , n78659 );
or ( n78662 , n78591 , n78660 , n78661 );
and ( n78663 , n78568 , n78662 );
xor ( n78664 , n78492 , n78494 );
xor ( n78665 , n78664 , n78560 );
and ( n78666 , n78662 , n78665 );
and ( n78667 , n78568 , n78665 );
or ( n78668 , n78663 , n78666 , n78667 );
and ( n78669 , n78565 , n78668 );
and ( n78670 , n78563 , n78668 );
or ( n78671 , n78566 , n78669 , n78670 );
and ( n78672 , n78437 , n78671 );
and ( n78673 , n78435 , n78671 );
or ( n78674 , n78438 , n78672 , n78673 );
and ( n78675 , n78393 , n78674 );
and ( n78676 , n78391 , n78674 );
or ( n78677 , n78394 , n78675 , n78676 );
and ( n78678 , n78330 , n78677 );
and ( n78679 , n78328 , n78677 );
or ( n78680 , n78331 , n78678 , n78679 );
and ( n78681 , n78282 , n78680 );
and ( n78682 , n78280 , n78680 );
or ( n78683 , n78283 , n78681 , n78682 );
and ( n78684 , n78204 , n78683 );
and ( n78685 , n78145 , n78683 );
or ( n78686 , n78205 , n78684 , n78685 );
and ( n78687 , n78142 , n78686 );
and ( n78688 , n78140 , n78686 );
or ( n78689 , n78143 , n78687 , n78688 );
xnor ( n78690 , n78093 , n78689 );
xor ( n78691 , n78140 , n78142 );
xor ( n78692 , n78691 , n78686 );
not ( n78693 , n78692 );
xor ( n78694 , n78145 , n78204 );
xor ( n78695 , n78694 , n78683 );
xor ( n78696 , n78280 , n78282 );
xor ( n78697 , n78696 , n78680 );
xor ( n78698 , n78328 , n78330 );
xor ( n78699 , n78698 , n78677 );
xor ( n78700 , n78391 , n78393 );
xor ( n78701 , n78700 , n78674 );
not ( n78702 , n78701 );
xor ( n78703 , n78435 , n78437 );
xor ( n78704 , n78703 , n78671 );
xor ( n78705 , n78563 , n78565 );
xor ( n78706 , n78705 , n78668 );
xor ( n78707 , n78497 , n78499 );
xor ( n78708 , n78707 , n78557 );
xor ( n78709 , n78505 , n78506 );
xor ( n78710 , n78709 , n78554 );
xor ( n78711 , n78573 , n78582 );
xor ( n78712 , n78711 , n78585 );
and ( n78713 , n78710 , n78712 );
xor ( n78714 , n78576 , n78577 );
xor ( n78715 , n78714 , n78579 );
and ( n78716 , n78528 , n78075 );
and ( n78717 , n78336 , n78121 );
and ( n78718 , n78716 , n78717 );
and ( n78719 , n78252 , n78156 );
and ( n78720 , n78717 , n78719 );
and ( n78721 , n78716 , n78719 );
or ( n78722 , n78718 , n78720 , n78721 );
and ( n78723 , n78050 , n78516 );
and ( n78724 , n78722 , n78723 );
and ( n78725 , n78062 , n78519 );
and ( n78726 , n78723 , n78725 );
and ( n78727 , n78722 , n78725 );
or ( n78728 , n78724 , n78726 , n78727 );
xor ( n78729 , n78517 , n78520 );
xor ( n78730 , n78729 , n78522 );
or ( n78731 , n78728 , n78730 );
and ( n78732 , n78070 , n78519 );
and ( n78733 , n78116 , n78345 );
and ( n78734 , n78732 , n78733 );
and ( n78735 , n78167 , n78235 );
and ( n78736 , n78733 , n78735 );
and ( n78737 , n78732 , n78735 );
or ( n78738 , n78734 , n78736 , n78737 );
and ( n78739 , n78541 , n78055 );
and ( n78740 , n78738 , n78739 );
and ( n78741 , n78528 , n78059 );
and ( n78742 , n78739 , n78741 );
and ( n78743 , n78738 , n78741 );
or ( n78744 , n78740 , n78742 , n78743 );
xor ( n78745 , n78542 , n78543 );
xor ( n78746 , n78745 , n78545 );
or ( n78747 , n78744 , n78746 );
and ( n78748 , n78731 , n78747 );
and ( n78749 , n78715 , n78748 );
xor ( n78750 , n78607 , n78609 );
xnor ( n78751 , n78638 , n78639 );
xnor ( n78752 , n78641 , n78642 );
and ( n78753 , n78751 , n78752 );
buf ( n78754 , n78167 );
or ( n78755 , n78753 , n78754 );
and ( n78756 , n78750 , n78755 );
xor ( n78757 , n78627 , n78636 );
xor ( n78758 , n78640 , n78643 );
and ( n78759 , n78757 , n78758 );
xor ( n78760 , n78647 , n78649 );
and ( n78761 , n78758 , n78760 );
and ( n78762 , n78757 , n78760 );
or ( n78763 , n78759 , n78761 , n78762 );
and ( n78764 , n78755 , n78763 );
and ( n78765 , n78750 , n78763 );
or ( n78766 , n78756 , n78764 , n78765 );
and ( n78767 , n78748 , n78766 );
and ( n78768 , n78715 , n78766 );
or ( n78769 , n78749 , n78767 , n78768 );
and ( n78770 , n78712 , n78769 );
and ( n78771 , n78710 , n78769 );
or ( n78772 , n78713 , n78770 , n78771 );
and ( n78773 , n78708 , n78772 );
xor ( n78774 , n78588 , n78590 );
xor ( n78775 , n78774 , n78659 );
and ( n78776 , n78772 , n78775 );
and ( n78777 , n78708 , n78775 );
or ( n78778 , n78773 , n78776 , n78777 );
xor ( n78779 , n78568 , n78662 );
xor ( n78780 , n78779 , n78665 );
and ( n78781 , n78778 , n78780 );
xor ( n78782 , n78593 , n78604 );
xor ( n78783 , n78782 , n78656 );
xor ( n78784 , n78598 , n78599 );
xor ( n78785 , n78784 , n78601 );
xor ( n78786 , n78610 , n78617 );
xor ( n78787 , n78786 , n78653 );
and ( n78788 , n78785 , n78787 );
xor ( n78789 , n78611 , n78612 );
xor ( n78790 , n78789 , n78614 );
xor ( n78791 , n78637 , n78644 );
xor ( n78792 , n78791 , n78650 );
and ( n78793 , n78790 , n78792 );
xor ( n78794 , n78731 , n78747 );
and ( n78795 , n78792 , n78794 );
and ( n78796 , n78790 , n78794 );
or ( n78797 , n78793 , n78795 , n78796 );
and ( n78798 , n78787 , n78797 );
and ( n78799 , n78785 , n78797 );
or ( n78800 , n78788 , n78798 , n78799 );
and ( n78801 , n78783 , n78800 );
xor ( n78802 , n78710 , n78712 );
xor ( n78803 , n78802 , n78769 );
and ( n78804 , n78800 , n78803 );
and ( n78805 , n78783 , n78803 );
or ( n78806 , n78801 , n78804 , n78805 );
xor ( n78807 , n78708 , n78772 );
xor ( n78808 , n78807 , n78775 );
and ( n78809 , n78806 , n78808 );
xnor ( n78810 , n78753 , n78754 );
and ( n78811 , n78620 , n78055 );
and ( n78812 , n78541 , n78059 );
and ( n78813 , n78811 , n78812 );
and ( n78814 , n78449 , n78103 );
and ( n78815 , n78812 , n78814 );
and ( n78816 , n78811 , n78814 );
or ( n78817 , n78813 , n78815 , n78816 );
and ( n78818 , n78050 , n78629 );
and ( n78819 , n78062 , n78516 );
and ( n78820 , n78818 , n78819 );
and ( n78821 , n78098 , n78440 );
and ( n78822 , n78819 , n78821 );
and ( n78823 , n78818 , n78821 );
or ( n78824 , n78820 , n78822 , n78823 );
and ( n78825 , n78817 , n78824 );
and ( n78826 , n78810 , n78825 );
xor ( n78827 , n78621 , n78622 );
xor ( n78828 , n78827 , n78624 );
xor ( n78829 , n78630 , n78631 );
xor ( n78830 , n78829 , n78633 );
and ( n78831 , n78828 , n78830 );
and ( n78832 , n78825 , n78831 );
and ( n78833 , n78810 , n78831 );
or ( n78834 , n78826 , n78832 , n78833 );
xnor ( n78835 , n78728 , n78730 );
xnor ( n78836 , n78744 , n78746 );
and ( n78837 , n78835 , n78836 );
and ( n78838 , n78834 , n78837 );
buf ( n78839 , n623 );
buf ( n78840 , n78839 );
and ( n78841 , n78840 , n78052 );
buf ( n78842 , n622 );
buf ( n78843 , n78842 );
and ( n78844 , n78843 , n78055 );
and ( n78845 , n78841 , n78844 );
and ( n78846 , n78449 , n78121 );
and ( n78847 , n78844 , n78846 );
and ( n78848 , n78841 , n78846 );
or ( n78849 , n78845 , n78847 , n78848 );
and ( n78850 , n78244 , n78235 );
and ( n78851 , n78252 , n78261 );
and ( n78852 , n78850 , n78851 );
and ( n78853 , n78849 , n78852 );
buf ( n78854 , n622 );
buf ( n78855 , n78854 );
and ( n78856 , n78047 , n78855 );
and ( n78857 , n78852 , n78856 );
and ( n78858 , n78849 , n78856 );
or ( n78859 , n78853 , n78857 , n78858 );
and ( n78860 , n78070 , n78516 );
and ( n78861 , n78098 , n78519 );
and ( n78862 , n78860 , n78861 );
and ( n78863 , n78167 , n78345 );
and ( n78864 , n78861 , n78863 );
and ( n78865 , n78860 , n78863 );
or ( n78866 , n78862 , n78864 , n78865 );
xor ( n78867 , n78811 , n78812 );
xor ( n78868 , n78867 , n78814 );
and ( n78869 , n78866 , n78868 );
xor ( n78870 , n78716 , n78717 );
xor ( n78871 , n78870 , n78719 );
and ( n78872 , n78868 , n78871 );
and ( n78873 , n78866 , n78871 );
or ( n78874 , n78869 , n78872 , n78873 );
and ( n78875 , n78859 , n78874 );
xor ( n78876 , n78722 , n78723 );
xor ( n78877 , n78876 , n78725 );
and ( n78878 , n78874 , n78877 );
and ( n78879 , n78859 , n78877 );
or ( n78880 , n78875 , n78878 , n78879 );
xor ( n78881 , n78738 , n78739 );
xor ( n78882 , n78881 , n78741 );
xor ( n78883 , n78817 , n78824 );
and ( n78884 , n78882 , n78883 );
xor ( n78885 , n78828 , n78830 );
and ( n78886 , n78883 , n78885 );
and ( n78887 , n78882 , n78885 );
or ( n78888 , n78884 , n78886 , n78887 );
and ( n78889 , n78880 , n78888 );
xor ( n78890 , n78751 , n78752 );
and ( n78891 , n78541 , n78075 );
and ( n78892 , n78528 , n78103 );
and ( n78893 , n78891 , n78892 );
and ( n78894 , n78336 , n78156 );
and ( n78895 , n78892 , n78894 );
and ( n78896 , n78891 , n78894 );
or ( n78897 , n78893 , n78895 , n78896 );
xor ( n78898 , n78818 , n78819 );
xor ( n78899 , n78898 , n78821 );
and ( n78900 , n78897 , n78899 );
xor ( n78901 , n78732 , n78733 );
xor ( n78902 , n78901 , n78735 );
and ( n78903 , n78899 , n78902 );
and ( n78904 , n78897 , n78902 );
or ( n78905 , n78900 , n78903 , n78904 );
and ( n78906 , n78890 , n78905 );
and ( n78907 , n78843 , n78052 );
buf ( n78908 , n78244 );
and ( n78909 , n78907 , n78908 );
buf ( n78910 , n623 );
buf ( n78911 , n78910 );
and ( n78912 , n78047 , n78911 );
and ( n78913 , n78050 , n78855 );
and ( n78914 , n78912 , n78913 );
and ( n78915 , n78116 , n78440 );
and ( n78916 , n78913 , n78915 );
and ( n78917 , n78912 , n78915 );
or ( n78918 , n78914 , n78916 , n78917 );
and ( n78919 , n78908 , n78918 );
and ( n78920 , n78907 , n78918 );
or ( n78921 , n78909 , n78919 , n78920 );
and ( n78922 , n78905 , n78921 );
and ( n78923 , n78890 , n78921 );
or ( n78924 , n78906 , n78922 , n78923 );
and ( n78925 , n78888 , n78924 );
and ( n78926 , n78880 , n78924 );
or ( n78927 , n78889 , n78925 , n78926 );
and ( n78928 , n78837 , n78927 );
and ( n78929 , n78834 , n78927 );
or ( n78930 , n78838 , n78928 , n78929 );
xor ( n78931 , n78715 , n78748 );
xor ( n78932 , n78931 , n78766 );
and ( n78933 , n78930 , n78932 );
xor ( n78934 , n78750 , n78755 );
xor ( n78935 , n78934 , n78763 );
xor ( n78936 , n78757 , n78758 );
xor ( n78937 , n78936 , n78760 );
xor ( n78938 , n78810 , n78825 );
xor ( n78939 , n78938 , n78831 );
and ( n78940 , n78937 , n78939 );
xor ( n78941 , n78835 , n78836 );
and ( n78942 , n78939 , n78941 );
and ( n78943 , n78937 , n78941 );
or ( n78944 , n78940 , n78942 , n78943 );
and ( n78945 , n78935 , n78944 );
xor ( n78946 , n78859 , n78874 );
xor ( n78947 , n78946 , n78877 );
and ( n78948 , n78070 , n78629 );
and ( n78949 , n78098 , n78516 );
and ( n78950 , n78948 , n78949 );
and ( n78951 , n78116 , n78519 );
and ( n78952 , n78949 , n78951 );
and ( n78953 , n78948 , n78951 );
or ( n78954 , n78950 , n78952 , n78953 );
xor ( n78955 , n78891 , n78892 );
xor ( n78956 , n78955 , n78894 );
and ( n78957 , n78954 , n78956 );
xor ( n78958 , n78841 , n78844 );
xor ( n78959 , n78958 , n78846 );
and ( n78960 , n78956 , n78959 );
and ( n78961 , n78954 , n78959 );
or ( n78962 , n78957 , n78960 , n78961 );
and ( n78963 , n78620 , n78075 );
and ( n78964 , n78541 , n78103 );
and ( n78965 , n78963 , n78964 );
and ( n78966 , n78528 , n78121 );
and ( n78967 , n78964 , n78966 );
and ( n78968 , n78963 , n78966 );
or ( n78969 , n78965 , n78967 , n78968 );
xor ( n78970 , n78860 , n78861 );
xor ( n78971 , n78970 , n78863 );
and ( n78972 , n78969 , n78971 );
xor ( n78973 , n78912 , n78913 );
xor ( n78974 , n78973 , n78915 );
and ( n78975 , n78971 , n78974 );
and ( n78976 , n78969 , n78974 );
or ( n78977 , n78972 , n78975 , n78976 );
and ( n78978 , n78962 , n78977 );
and ( n78979 , n78947 , n78978 );
xor ( n78980 , n78866 , n78868 );
xor ( n78981 , n78980 , n78871 );
xor ( n78982 , n78897 , n78899 );
xor ( n78983 , n78982 , n78902 );
and ( n78984 , n78981 , n78983 );
and ( n78985 , n78978 , n78984 );
and ( n78986 , n78947 , n78984 );
or ( n78987 , n78979 , n78985 , n78986 );
and ( n78988 , n78062 , n78629 );
and ( n78989 , n78620 , n78059 );
and ( n78990 , n78988 , n78989 );
xor ( n78991 , n78849 , n78852 );
xor ( n78992 , n78991 , n78856 );
and ( n78993 , n78990 , n78992 );
and ( n78994 , n78840 , n78055 );
and ( n78995 , n78843 , n78059 );
or ( n78996 , n78994 , n78995 );
and ( n78997 , n78050 , n78911 );
and ( n78998 , n78062 , n78855 );
or ( n78999 , n78997 , n78998 );
and ( n79000 , n78996 , n78999 );
and ( n79001 , n78992 , n79000 );
and ( n79002 , n78990 , n79000 );
or ( n79003 , n78993 , n79001 , n79002 );
and ( n79004 , n78449 , n78156 );
not ( n79005 , n79004 );
and ( n79006 , n78336 , n78261 );
and ( n79007 , n79005 , n79006 );
and ( n79008 , n78167 , n78440 );
not ( n79009 , n79008 );
and ( n79010 , n78244 , n78345 );
and ( n79011 , n79009 , n79010 );
and ( n79012 , n79007 , n79011 );
buf ( n79013 , n79004 );
buf ( n79014 , n79008 );
and ( n79015 , n79013 , n79014 );
and ( n79016 , n79012 , n79015 );
xor ( n79017 , n78907 , n78908 );
xor ( n79018 , n79017 , n78918 );
and ( n79019 , n79015 , n79018 );
and ( n79020 , n79012 , n79018 );
or ( n79021 , n79016 , n79019 , n79020 );
and ( n79022 , n79003 , n79021 );
xor ( n79023 , n78882 , n78883 );
xor ( n79024 , n79023 , n78885 );
and ( n79025 , n79021 , n79024 );
and ( n79026 , n79003 , n79024 );
or ( n79027 , n79022 , n79025 , n79026 );
and ( n79028 , n78987 , n79027 );
xor ( n79029 , n78880 , n78888 );
xor ( n79030 , n79029 , n78924 );
and ( n79031 , n79027 , n79030 );
and ( n79032 , n78987 , n79030 );
or ( n79033 , n79028 , n79031 , n79032 );
and ( n79034 , n78944 , n79033 );
and ( n79035 , n78935 , n79033 );
or ( n79036 , n78945 , n79034 , n79035 );
and ( n79037 , n78932 , n79036 );
and ( n79038 , n78930 , n79036 );
or ( n79039 , n78933 , n79037 , n79038 );
xor ( n79040 , n78783 , n78800 );
xor ( n79041 , n79040 , n78803 );
and ( n79042 , n79039 , n79041 );
xor ( n79043 , n78785 , n78787 );
xor ( n79044 , n79043 , n78797 );
xor ( n79045 , n78790 , n78792 );
xor ( n79046 , n79045 , n78794 );
xor ( n79047 , n78834 , n78837 );
xor ( n79048 , n79047 , n78927 );
and ( n79049 , n79046 , n79048 );
xor ( n79050 , n78890 , n78905 );
xor ( n79051 , n79050 , n78921 );
xor ( n79052 , n78962 , n78977 );
xor ( n79053 , n78981 , n78983 );
and ( n79054 , n79052 , n79053 );
xnor ( n79055 , n78997 , n78998 );
not ( n79056 , n79055 );
xor ( n79057 , n79009 , n79010 );
and ( n79058 , n79056 , n79057 );
xnor ( n79059 , n78994 , n78995 );
not ( n79060 , n79059 );
xor ( n79061 , n79005 , n79006 );
and ( n79062 , n79060 , n79061 );
and ( n79063 , n79058 , n79062 );
and ( n79064 , n79053 , n79063 );
and ( n79065 , n79052 , n79063 );
or ( n79066 , n79054 , n79064 , n79065 );
and ( n79067 , n79051 , n79066 );
buf ( n79068 , n79055 );
buf ( n79069 , n79059 );
and ( n79070 , n79068 , n79069 );
xor ( n79071 , n78954 , n78956 );
xor ( n79072 , n79071 , n78959 );
xor ( n79073 , n78969 , n78971 );
xor ( n79074 , n79073 , n78974 );
and ( n79075 , n79072 , n79074 );
and ( n79076 , n79070 , n79075 );
xor ( n79077 , n78988 , n78989 );
xor ( n79078 , n78850 , n78851 );
and ( n79079 , n79077 , n79078 );
xor ( n79080 , n78996 , n78999 );
and ( n79081 , n79078 , n79080 );
and ( n79082 , n79077 , n79080 );
or ( n79083 , n79079 , n79081 , n79082 );
and ( n79084 , n79075 , n79083 );
and ( n79085 , n79070 , n79083 );
or ( n79086 , n79076 , n79084 , n79085 );
and ( n79087 , n79066 , n79086 );
and ( n79088 , n79051 , n79086 );
or ( n79089 , n79067 , n79087 , n79088 );
xor ( n79090 , n79007 , n79011 );
xor ( n79091 , n79013 , n79014 );
and ( n79092 , n79090 , n79091 );
and ( n79093 , n78840 , n78059 );
and ( n79094 , n78541 , n78121 );
and ( n79095 , n79093 , n79094 );
and ( n79096 , n78528 , n78156 );
and ( n79097 , n79094 , n79096 );
and ( n79098 , n79093 , n79096 );
or ( n79099 , n79095 , n79097 , n79098 );
and ( n79100 , n78843 , n78075 );
and ( n79101 , n78620 , n78103 );
and ( n79102 , n79100 , n79101 );
and ( n79103 , n78449 , n78261 );
and ( n79104 , n79101 , n79103 );
and ( n79105 , n79100 , n79103 );
or ( n79106 , n79102 , n79104 , n79105 );
and ( n79107 , n79099 , n79106 );
and ( n79108 , n78252 , n78345 );
and ( n79109 , n78336 , n78235 );
and ( n79110 , n79108 , n79109 );
and ( n79111 , n79106 , n79110 );
and ( n79112 , n79099 , n79110 );
or ( n79113 , n79107 , n79111 , n79112 );
and ( n79114 , n79091 , n79113 );
and ( n79115 , n79090 , n79113 );
or ( n79116 , n79092 , n79114 , n79115 );
xor ( n79117 , n78990 , n78992 );
xor ( n79118 , n79117 , n79000 );
and ( n79119 , n79116 , n79118 );
xor ( n79120 , n79012 , n79015 );
xor ( n79121 , n79120 , n79018 );
and ( n79122 , n79118 , n79121 );
and ( n79123 , n79116 , n79121 );
or ( n79124 , n79119 , n79122 , n79123 );
xor ( n79125 , n78947 , n78978 );
xor ( n79126 , n79125 , n78984 );
and ( n79127 , n79124 , n79126 );
xor ( n79128 , n79003 , n79021 );
xor ( n79129 , n79128 , n79024 );
and ( n79130 , n79126 , n79129 );
and ( n79131 , n79124 , n79129 );
or ( n79132 , n79127 , n79130 , n79131 );
and ( n79133 , n79089 , n79132 );
xor ( n79134 , n78937 , n78939 );
xor ( n79135 , n79134 , n78941 );
and ( n79136 , n79132 , n79135 );
and ( n79137 , n79089 , n79135 );
or ( n79138 , n79133 , n79136 , n79137 );
and ( n79139 , n79048 , n79138 );
and ( n79140 , n79046 , n79138 );
or ( n79141 , n79049 , n79139 , n79140 );
and ( n79142 , n79044 , n79141 );
xor ( n79143 , n78930 , n78932 );
xor ( n79144 , n79143 , n79036 );
and ( n79145 , n79141 , n79144 );
and ( n79146 , n79044 , n79144 );
or ( n79147 , n79142 , n79145 , n79146 );
and ( n79148 , n79041 , n79147 );
and ( n79149 , n79039 , n79147 );
or ( n79150 , n79042 , n79148 , n79149 );
and ( n79151 , n78808 , n79150 );
and ( n79152 , n78806 , n79150 );
or ( n79153 , n78809 , n79151 , n79152 );
and ( n79154 , n78780 , n79153 );
and ( n79155 , n78778 , n79153 );
or ( n79156 , n78781 , n79154 , n79155 );
or ( n79157 , n78706 , n79156 );
and ( n79158 , n78704 , n79157 );
xor ( n79159 , n78704 , n79157 );
xnor ( n79160 , n78706 , n79156 );
xor ( n79161 , n78778 , n78780 );
xor ( n79162 , n79161 , n79153 );
xor ( n79163 , n78806 , n78808 );
xor ( n79164 , n79163 , n79150 );
not ( n79165 , n79164 );
xor ( n79166 , n79039 , n79041 );
xor ( n79167 , n79166 , n79147 );
xor ( n79168 , n78935 , n78944 );
xor ( n79169 , n79168 , n79033 );
xor ( n79170 , n78987 , n79027 );
xor ( n79171 , n79170 , n79030 );
xor ( n79172 , n78963 , n78964 );
xor ( n79173 , n79172 , n78966 );
xor ( n79174 , n78948 , n78949 );
xor ( n79175 , n79174 , n78951 );
and ( n79176 , n79173 , n79175 );
buf ( n79177 , n78252 );
and ( n79178 , n78062 , n78911 );
and ( n79179 , n78116 , n78516 );
and ( n79180 , n79178 , n79179 );
and ( n79181 , n78167 , n78519 );
and ( n79182 , n79179 , n79181 );
and ( n79183 , n79178 , n79181 );
or ( n79184 , n79180 , n79182 , n79183 );
and ( n79185 , n79177 , n79184 );
and ( n79186 , n78070 , n78855 );
and ( n79187 , n78098 , n78629 );
and ( n79188 , n79186 , n79187 );
and ( n79189 , n78244 , n78440 );
and ( n79190 , n79187 , n79189 );
and ( n79191 , n79186 , n79189 );
or ( n79192 , n79188 , n79190 , n79191 );
and ( n79193 , n79184 , n79192 );
and ( n79194 , n79177 , n79192 );
or ( n79195 , n79185 , n79193 , n79194 );
and ( n79196 , n79176 , n79195 );
xor ( n79197 , n79058 , n79062 );
and ( n79198 , n79195 , n79197 );
and ( n79199 , n79176 , n79197 );
or ( n79200 , n79196 , n79198 , n79199 );
xor ( n79201 , n79068 , n79069 );
xor ( n79202 , n79072 , n79074 );
and ( n79203 , n79201 , n79202 );
xor ( n79204 , n79056 , n79057 );
xor ( n79205 , n79060 , n79061 );
and ( n79206 , n79204 , n79205 );
and ( n79207 , n79202 , n79206 );
and ( n79208 , n79201 , n79206 );
or ( n79209 , n79203 , n79207 , n79208 );
and ( n79210 , n79200 , n79209 );
xor ( n79211 , n79173 , n79175 );
xor ( n79212 , n79093 , n79094 );
xor ( n79213 , n79212 , n79096 );
xor ( n79214 , n79100 , n79101 );
xor ( n79215 , n79214 , n79103 );
or ( n79216 , n79213 , n79215 );
and ( n79217 , n79211 , n79216 );
and ( n79218 , n78843 , n78103 );
and ( n79219 , n78620 , n78121 );
and ( n79220 , n79218 , n79219 );
and ( n79221 , n78541 , n78156 );
and ( n79222 , n79219 , n79221 );
and ( n79223 , n79218 , n79221 );
or ( n79224 , n79220 , n79222 , n79223 );
and ( n79225 , n78098 , n78855 );
and ( n79226 , n78116 , n78629 );
and ( n79227 , n79225 , n79226 );
and ( n79228 , n78167 , n78516 );
and ( n79229 , n79226 , n79228 );
and ( n79230 , n79225 , n79228 );
or ( n79231 , n79227 , n79229 , n79230 );
and ( n79232 , n79224 , n79231 );
and ( n79233 , n79216 , n79232 );
and ( n79234 , n79211 , n79232 );
or ( n79235 , n79217 , n79233 , n79234 );
xor ( n79236 , n79077 , n79078 );
xor ( n79237 , n79236 , n79080 );
and ( n79238 , n79235 , n79237 );
xor ( n79239 , n79090 , n79091 );
xor ( n79240 , n79239 , n79113 );
and ( n79241 , n79237 , n79240 );
and ( n79242 , n79235 , n79240 );
or ( n79243 , n79238 , n79241 , n79242 );
and ( n79244 , n79209 , n79243 );
and ( n79245 , n79200 , n79243 );
or ( n79246 , n79210 , n79244 , n79245 );
xor ( n79247 , n79052 , n79053 );
xor ( n79248 , n79247 , n79063 );
xor ( n79249 , n79070 , n79075 );
xor ( n79250 , n79249 , n79083 );
and ( n79251 , n79248 , n79250 );
xor ( n79252 , n79116 , n79118 );
xor ( n79253 , n79252 , n79121 );
and ( n79254 , n79250 , n79253 );
and ( n79255 , n79248 , n79253 );
or ( n79256 , n79251 , n79254 , n79255 );
and ( n79257 , n79246 , n79256 );
xor ( n79258 , n79051 , n79066 );
xor ( n79259 , n79258 , n79086 );
and ( n79260 , n79256 , n79259 );
and ( n79261 , n79246 , n79259 );
or ( n79262 , n79257 , n79260 , n79261 );
and ( n79263 , n79171 , n79262 );
xor ( n79264 , n79089 , n79132 );
xor ( n79265 , n79264 , n79135 );
and ( n79266 , n79262 , n79265 );
and ( n79267 , n79171 , n79265 );
or ( n79268 , n79263 , n79266 , n79267 );
and ( n79269 , n79169 , n79268 );
xor ( n79270 , n79046 , n79048 );
xor ( n79271 , n79270 , n79138 );
and ( n79272 , n79268 , n79271 );
and ( n79273 , n79169 , n79271 );
or ( n79274 , n79269 , n79272 , n79273 );
xor ( n79275 , n79044 , n79141 );
xor ( n79276 , n79275 , n79144 );
and ( n79277 , n79274 , n79276 );
xor ( n79278 , n79169 , n79268 );
xor ( n79279 , n79278 , n79271 );
xor ( n79280 , n79124 , n79126 );
xor ( n79281 , n79280 , n79129 );
and ( n79282 , n78244 , n78519 );
and ( n79283 , n78252 , n78440 );
xor ( n79284 , n79282 , n79283 );
and ( n79285 , n78336 , n78440 );
and ( n79286 , n78449 , n78345 );
and ( n79287 , n79285 , n79286 );
and ( n79288 , n79284 , n79287 );
and ( n79289 , n78070 , n78911 );
and ( n79290 , n79287 , n79289 );
and ( n79291 , n79284 , n79289 );
or ( n79292 , n79288 , n79290 , n79291 );
xor ( n79293 , n79178 , n79179 );
xor ( n79294 , n79293 , n79181 );
and ( n79295 , n79292 , n79294 );
xor ( n79296 , n79186 , n79187 );
xor ( n79297 , n79296 , n79189 );
and ( n79298 , n79294 , n79297 );
and ( n79299 , n79292 , n79297 );
or ( n79300 , n79295 , n79298 , n79299 );
xor ( n79301 , n79099 , n79106 );
xor ( n79302 , n79301 , n79110 );
or ( n79303 , n79300 , n79302 );
and ( n79304 , n78528 , n78261 );
and ( n79305 , n78449 , n78235 );
and ( n79306 , n79304 , n79305 );
and ( n79307 , n79282 , n79283 );
and ( n79308 , n79306 , n79307 );
xor ( n79309 , n79177 , n79184 );
xor ( n79310 , n79309 , n79192 );
and ( n79311 , n79308 , n79310 );
xor ( n79312 , n79204 , n79205 );
and ( n79313 , n79310 , n79312 );
and ( n79314 , n79308 , n79312 );
or ( n79315 , n79311 , n79313 , n79314 );
and ( n79316 , n79303 , n79315 );
xor ( n79317 , n79176 , n79195 );
xor ( n79318 , n79317 , n79197 );
and ( n79319 , n79315 , n79318 );
and ( n79320 , n79303 , n79318 );
or ( n79321 , n79316 , n79319 , n79320 );
xor ( n79322 , n79200 , n79209 );
xor ( n79323 , n79322 , n79243 );
and ( n79324 , n79321 , n79323 );
xor ( n79325 , n79248 , n79250 );
xor ( n79326 , n79325 , n79253 );
and ( n79327 , n79323 , n79326 );
and ( n79328 , n79321 , n79326 );
or ( n79329 , n79324 , n79327 , n79328 );
and ( n79330 , n79281 , n79329 );
xor ( n79331 , n79246 , n79256 );
xor ( n79332 , n79331 , n79259 );
and ( n79333 , n79329 , n79332 );
and ( n79334 , n79281 , n79332 );
or ( n79335 , n79330 , n79333 , n79334 );
xor ( n79336 , n79171 , n79262 );
xor ( n79337 , n79336 , n79265 );
and ( n79338 , n79335 , n79337 );
xor ( n79339 , n79281 , n79329 );
xor ( n79340 , n79339 , n79332 );
xor ( n79341 , n79201 , n79202 );
xor ( n79342 , n79341 , n79206 );
xor ( n79343 , n79235 , n79237 );
xor ( n79344 , n79343 , n79240 );
and ( n79345 , n79342 , n79344 );
xor ( n79346 , n79108 , n79109 );
xnor ( n79347 , n79213 , n79215 );
and ( n79348 , n79346 , n79347 );
xor ( n79349 , n79224 , n79231 );
and ( n79350 , n79347 , n79349 );
and ( n79351 , n79346 , n79349 );
or ( n79352 , n79348 , n79350 , n79351 );
xor ( n79353 , n79211 , n79216 );
xor ( n79354 , n79353 , n79232 );
and ( n79355 , n79352 , n79354 );
xnor ( n79356 , n79300 , n79302 );
and ( n79357 , n79354 , n79356 );
and ( n79358 , n79352 , n79356 );
or ( n79359 , n79355 , n79357 , n79358 );
and ( n79360 , n79344 , n79359 );
and ( n79361 , n79342 , n79359 );
or ( n79362 , n79345 , n79360 , n79361 );
xor ( n79363 , n79321 , n79323 );
xor ( n79364 , n79363 , n79326 );
and ( n79365 , n79362 , n79364 );
and ( n79366 , n78167 , n78629 );
and ( n79367 , n78244 , n78516 );
and ( n79368 , n79366 , n79367 );
and ( n79369 , n78252 , n78519 );
and ( n79370 , n79367 , n79369 );
and ( n79371 , n79366 , n79369 );
or ( n79372 , n79368 , n79370 , n79371 );
and ( n79373 , n78541 , n78235 );
and ( n79374 , n78528 , n78345 );
and ( n79375 , n79373 , n79374 );
and ( n79376 , n78098 , n78911 );
and ( n79377 , n79375 , n79376 );
and ( n79378 , n78116 , n78855 );
and ( n79379 , n79376 , n79378 );
and ( n79380 , n79375 , n79378 );
or ( n79381 , n79377 , n79379 , n79380 );
and ( n79382 , n79372 , n79381 );
xor ( n79383 , n79218 , n79219 );
xor ( n79384 , n79383 , n79221 );
and ( n79385 , n79381 , n79384 );
and ( n79386 , n79372 , n79384 );
or ( n79387 , n79382 , n79385 , n79386 );
and ( n79388 , n78620 , n78156 );
and ( n79389 , n78541 , n78261 );
and ( n79390 , n79388 , n79389 );
and ( n79391 , n78528 , n78235 );
and ( n79392 , n79389 , n79391 );
and ( n79393 , n79388 , n79391 );
or ( n79394 , n79390 , n79392 , n79393 );
and ( n79395 , n78252 , n78516 );
and ( n79396 , n78336 , n78519 );
and ( n79397 , n79395 , n79396 );
and ( n79398 , n78840 , n78103 );
and ( n79399 , n79397 , n79398 );
and ( n79400 , n78843 , n78121 );
and ( n79401 , n79398 , n79400 );
and ( n79402 , n79397 , n79400 );
or ( n79403 , n79399 , n79401 , n79402 );
and ( n79404 , n79394 , n79403 );
xor ( n79405 , n79225 , n79226 );
xor ( n79406 , n79405 , n79228 );
and ( n79407 , n79403 , n79406 );
and ( n79408 , n79394 , n79406 );
or ( n79409 , n79404 , n79407 , n79408 );
and ( n79410 , n79387 , n79409 );
xor ( n79411 , n79306 , n79307 );
and ( n79412 , n78840 , n78075 );
buf ( n79413 , n78336 );
and ( n79414 , n79412 , n79413 );
xor ( n79415 , n79304 , n79305 );
and ( n79416 , n79413 , n79415 );
and ( n79417 , n79412 , n79415 );
or ( n79418 , n79414 , n79416 , n79417 );
and ( n79419 , n79411 , n79418 );
xor ( n79420 , n79292 , n79294 );
xor ( n79421 , n79420 , n79297 );
and ( n79422 , n79418 , n79421 );
and ( n79423 , n79411 , n79421 );
or ( n79424 , n79419 , n79422 , n79423 );
and ( n79425 , n79410 , n79424 );
xor ( n79426 , n79308 , n79310 );
xor ( n79427 , n79426 , n79312 );
and ( n79428 , n79424 , n79427 );
and ( n79429 , n79410 , n79427 );
or ( n79430 , n79425 , n79428 , n79429 );
xor ( n79431 , n79303 , n79315 );
xor ( n79432 , n79431 , n79318 );
and ( n79433 , n79430 , n79432 );
xor ( n79434 , n79284 , n79287 );
xor ( n79435 , n79434 , n79289 );
and ( n79436 , n78840 , n78121 );
and ( n79437 , n78843 , n78156 );
and ( n79438 , n79436 , n79437 );
and ( n79439 , n78620 , n78261 );
and ( n79440 , n79437 , n79439 );
and ( n79441 , n79436 , n79439 );
or ( n79442 , n79438 , n79440 , n79441 );
and ( n79443 , n78116 , n78911 );
and ( n79444 , n78167 , n78855 );
and ( n79445 , n79443 , n79444 );
and ( n79446 , n78244 , n78629 );
and ( n79447 , n79444 , n79446 );
and ( n79448 , n79443 , n79446 );
or ( n79449 , n79445 , n79447 , n79448 );
and ( n79450 , n79442 , n79449 );
and ( n79451 , n79435 , n79450 );
xor ( n79452 , n79388 , n79389 );
xor ( n79453 , n79452 , n79391 );
xor ( n79454 , n79366 , n79367 );
xor ( n79455 , n79454 , n79369 );
and ( n79456 , n79453 , n79455 );
and ( n79457 , n79450 , n79456 );
and ( n79458 , n79435 , n79456 );
or ( n79459 , n79451 , n79457 , n79458 );
xor ( n79460 , n79346 , n79347 );
xor ( n79461 , n79460 , n79349 );
and ( n79462 , n79459 , n79461 );
xor ( n79463 , n79387 , n79409 );
and ( n79464 , n79461 , n79463 );
and ( n79465 , n79459 , n79463 );
or ( n79466 , n79462 , n79464 , n79465 );
xor ( n79467 , n79372 , n79381 );
xor ( n79468 , n79467 , n79384 );
xor ( n79469 , n79394 , n79403 );
xor ( n79470 , n79469 , n79406 );
and ( n79471 , n79468 , n79470 );
xor ( n79472 , n79412 , n79413 );
xor ( n79473 , n79472 , n79415 );
xor ( n79474 , n79395 , n79396 );
and ( n79475 , n78843 , n78261 );
and ( n79476 , n78620 , n78235 );
and ( n79477 , n79475 , n79476 );
and ( n79478 , n78541 , n78345 );
and ( n79479 , n79476 , n79478 );
and ( n79480 , n79475 , n79478 );
or ( n79481 , n79477 , n79479 , n79480 );
and ( n79482 , n79474 , n79481 );
and ( n79483 , n78449 , n78519 );
and ( n79484 , n78528 , n78440 );
and ( n79485 , n79483 , n79484 );
and ( n79486 , n79481 , n79485 );
and ( n79487 , n79474 , n79485 );
or ( n79488 , n79482 , n79486 , n79487 );
xor ( n79489 , n79397 , n79398 );
xor ( n79490 , n79489 , n79400 );
or ( n79491 , n79488 , n79490 );
and ( n79492 , n79473 , n79491 );
xor ( n79493 , n79285 , n79286 );
xor ( n79494 , n79375 , n79376 );
xor ( n79495 , n79494 , n79378 );
and ( n79496 , n79493 , n79495 );
xor ( n79497 , n79442 , n79449 );
and ( n79498 , n79495 , n79497 );
and ( n79499 , n79493 , n79497 );
or ( n79500 , n79496 , n79498 , n79499 );
and ( n79501 , n79491 , n79500 );
and ( n79502 , n79473 , n79500 );
or ( n79503 , n79492 , n79501 , n79502 );
and ( n79504 , n79471 , n79503 );
xor ( n79505 , n79411 , n79418 );
xor ( n79506 , n79505 , n79421 );
and ( n79507 , n79503 , n79506 );
and ( n79508 , n79471 , n79506 );
or ( n79509 , n79504 , n79507 , n79508 );
and ( n79510 , n79466 , n79509 );
xor ( n79511 , n79352 , n79354 );
xor ( n79512 , n79511 , n79356 );
and ( n79513 , n79509 , n79512 );
and ( n79514 , n79466 , n79512 );
or ( n79515 , n79510 , n79513 , n79514 );
and ( n79516 , n79432 , n79515 );
and ( n79517 , n79430 , n79515 );
or ( n79518 , n79433 , n79516 , n79517 );
and ( n79519 , n79364 , n79518 );
and ( n79520 , n79362 , n79518 );
or ( n79521 , n79365 , n79519 , n79520 );
or ( n79522 , n79340 , n79521 );
and ( n79523 , n79337 , n79522 );
and ( n79524 , n79335 , n79522 );
or ( n79525 , n79338 , n79523 , n79524 );
or ( n79526 , n79279 , n79525 );
and ( n79527 , n79276 , n79526 );
and ( n79528 , n79274 , n79526 );
or ( n79529 , n79277 , n79527 , n79528 );
and ( n79530 , n79167 , n79529 );
xor ( n79531 , n79167 , n79529 );
xor ( n79532 , n79274 , n79276 );
xor ( n79533 , n79532 , n79526 );
not ( n79534 , n79533 );
xnor ( n79535 , n79279 , n79525 );
xor ( n79536 , n79335 , n79337 );
xor ( n79537 , n79536 , n79522 );
not ( n79538 , n79537 );
xnor ( n79539 , n79340 , n79521 );
xor ( n79540 , n79342 , n79344 );
xor ( n79541 , n79540 , n79359 );
xor ( n79542 , n79410 , n79424 );
xor ( n79543 , n79542 , n79427 );
xor ( n79544 , n79453 , n79455 );
xor ( n79545 , n79436 , n79437 );
xor ( n79546 , n79545 , n79439 );
xor ( n79547 , n79443 , n79444 );
xor ( n79548 , n79547 , n79446 );
and ( n79549 , n79546 , n79548 );
and ( n79550 , n79544 , n79549 );
buf ( n79551 , n78449 );
xor ( n79552 , n79373 , n79374 );
and ( n79553 , n79551 , n79552 );
and ( n79554 , n78244 , n78855 );
and ( n79555 , n78252 , n78629 );
and ( n79556 , n79554 , n79555 );
and ( n79557 , n78336 , n78516 );
and ( n79558 , n79555 , n79557 );
and ( n79559 , n79554 , n79557 );
or ( n79560 , n79556 , n79558 , n79559 );
and ( n79561 , n79552 , n79560 );
and ( n79562 , n79551 , n79560 );
or ( n79563 , n79553 , n79561 , n79562 );
and ( n79564 , n79549 , n79563 );
and ( n79565 , n79544 , n79563 );
or ( n79566 , n79550 , n79564 , n79565 );
xor ( n79567 , n79435 , n79450 );
xor ( n79568 , n79567 , n79456 );
and ( n79569 , n79566 , n79568 );
xor ( n79570 , n79468 , n79470 );
and ( n79571 , n79568 , n79570 );
and ( n79572 , n79566 , n79570 );
or ( n79573 , n79569 , n79571 , n79572 );
xor ( n79574 , n79459 , n79461 );
xor ( n79575 , n79574 , n79463 );
and ( n79576 , n79573 , n79575 );
xor ( n79577 , n79471 , n79503 );
xor ( n79578 , n79577 , n79506 );
and ( n79579 , n79575 , n79578 );
and ( n79580 , n79573 , n79578 );
or ( n79581 , n79576 , n79579 , n79580 );
and ( n79582 , n79543 , n79581 );
xor ( n79583 , n79466 , n79509 );
xor ( n79584 , n79583 , n79512 );
and ( n79585 , n79581 , n79584 );
and ( n79586 , n79543 , n79584 );
or ( n79587 , n79582 , n79585 , n79586 );
and ( n79588 , n79541 , n79587 );
xor ( n79589 , n79430 , n79432 );
xor ( n79590 , n79589 , n79515 );
and ( n79591 , n79587 , n79590 );
and ( n79592 , n79541 , n79590 );
or ( n79593 , n79588 , n79591 , n79592 );
xor ( n79594 , n79362 , n79364 );
xor ( n79595 , n79594 , n79518 );
and ( n79596 , n79593 , n79595 );
xor ( n79597 , n79593 , n79595 );
xor ( n79598 , n79541 , n79587 );
xor ( n79599 , n79598 , n79590 );
xor ( n79600 , n79543 , n79581 );
xor ( n79601 , n79600 , n79584 );
xnor ( n79602 , n79488 , n79490 );
and ( n79603 , n78336 , n78629 );
and ( n79604 , n78449 , n78516 );
and ( n79605 , n79603 , n79604 );
and ( n79606 , n78840 , n78156 );
or ( n79607 , n79605 , n79606 );
and ( n79608 , n78620 , n78345 );
and ( n79609 , n78541 , n78440 );
and ( n79610 , n79608 , n79609 );
and ( n79611 , n78167 , n78911 );
or ( n79612 , n79610 , n79611 );
and ( n79613 , n79607 , n79612 );
and ( n79614 , n79602 , n79613 );
xor ( n79615 , n79474 , n79481 );
xor ( n79616 , n79615 , n79485 );
xor ( n79617 , n79546 , n79548 );
and ( n79618 , n79616 , n79617 );
xor ( n79619 , n79554 , n79555 );
xor ( n79620 , n79619 , n79557 );
xor ( n79621 , n79483 , n79484 );
and ( n79622 , n79620 , n79621 );
and ( n79623 , n78840 , n78261 );
and ( n79624 , n78843 , n78235 );
or ( n79625 , n79623 , n79624 );
and ( n79626 , n79621 , n79625 );
and ( n79627 , n79620 , n79625 );
or ( n79628 , n79622 , n79626 , n79627 );
and ( n79629 , n79617 , n79628 );
and ( n79630 , n79616 , n79628 );
or ( n79631 , n79618 , n79629 , n79630 );
and ( n79632 , n79613 , n79631 );
and ( n79633 , n79602 , n79631 );
or ( n79634 , n79614 , n79632 , n79633 );
xor ( n79635 , n79473 , n79491 );
xor ( n79636 , n79635 , n79500 );
and ( n79637 , n79634 , n79636 );
xor ( n79638 , n79493 , n79495 );
xor ( n79639 , n79638 , n79497 );
xor ( n79640 , n79544 , n79549 );
xor ( n79641 , n79640 , n79563 );
and ( n79642 , n79639 , n79641 );
xor ( n79643 , n79551 , n79552 );
xor ( n79644 , n79643 , n79560 );
xor ( n79645 , n79607 , n79612 );
and ( n79646 , n79644 , n79645 );
and ( n79647 , n78528 , n78516 );
and ( n79648 , n78541 , n78519 );
and ( n79649 , n79647 , n79648 );
and ( n79650 , n78244 , n78911 );
and ( n79651 , n79649 , n79650 );
and ( n79652 , n78252 , n78855 );
and ( n79653 , n79650 , n79652 );
and ( n79654 , n79649 , n79652 );
or ( n79655 , n79651 , n79653 , n79654 );
xor ( n79656 , n79475 , n79476 );
xor ( n79657 , n79656 , n79478 );
or ( n79658 , n79655 , n79657 );
and ( n79659 , n79645 , n79658 );
and ( n79660 , n79644 , n79658 );
or ( n79661 , n79646 , n79659 , n79660 );
and ( n79662 , n79641 , n79661 );
and ( n79663 , n79639 , n79661 );
or ( n79664 , n79642 , n79662 , n79663 );
and ( n79665 , n79636 , n79664 );
and ( n79666 , n79634 , n79664 );
or ( n79667 , n79637 , n79665 , n79666 );
xor ( n79668 , n79573 , n79575 );
xor ( n79669 , n79668 , n79578 );
and ( n79670 , n79667 , n79669 );
xor ( n79671 , n79566 , n79568 );
xor ( n79672 , n79671 , n79570 );
xor ( n79673 , n79602 , n79613 );
xor ( n79674 , n79673 , n79631 );
xnor ( n79675 , n79605 , n79606 );
xnor ( n79676 , n79610 , n79611 );
and ( n79677 , n79675 , n79676 );
xor ( n79678 , n79616 , n79617 );
xor ( n79679 , n79678 , n79628 );
and ( n79680 , n79677 , n79679 );
and ( n79681 , n78252 , n78911 );
and ( n79682 , n78336 , n78855 );
and ( n79683 , n79681 , n79682 );
and ( n79684 , n78449 , n78629 );
and ( n79685 , n79682 , n79684 );
and ( n79686 , n79681 , n79684 );
or ( n79687 , n79683 , n79685 , n79686 );
xor ( n79688 , n79608 , n79609 );
or ( n79689 , n79687 , n79688 );
xor ( n79690 , n79620 , n79621 );
xor ( n79691 , n79690 , n79625 );
and ( n79692 , n79689 , n79691 );
xnor ( n79693 , n79655 , n79657 );
and ( n79694 , n79691 , n79693 );
and ( n79695 , n79689 , n79693 );
or ( n79696 , n79692 , n79694 , n79695 );
and ( n79697 , n79679 , n79696 );
and ( n79698 , n79677 , n79696 );
or ( n79699 , n79680 , n79697 , n79698 );
and ( n79700 , n79674 , n79699 );
xor ( n79701 , n79639 , n79641 );
xor ( n79702 , n79701 , n79661 );
and ( n79703 , n79699 , n79702 );
and ( n79704 , n79674 , n79702 );
or ( n79705 , n79700 , n79703 , n79704 );
and ( n79706 , n79672 , n79705 );
xor ( n79707 , n79634 , n79636 );
xor ( n79708 , n79707 , n79664 );
and ( n79709 , n79705 , n79708 );
and ( n79710 , n79672 , n79708 );
or ( n79711 , n79706 , n79709 , n79710 );
and ( n79712 , n79669 , n79711 );
and ( n79713 , n79667 , n79711 );
or ( n79714 , n79670 , n79712 , n79713 );
and ( n79715 , n79601 , n79714 );
xor ( n79716 , n79601 , n79714 );
xor ( n79717 , n79667 , n79669 );
xor ( n79718 , n79717 , n79711 );
xor ( n79719 , n79672 , n79705 );
xor ( n79720 , n79719 , n79708 );
xor ( n79721 , n79675 , n79676 );
xor ( n79722 , n79603 , n79604 );
and ( n79723 , n78840 , n78235 );
and ( n79724 , n78843 , n78345 );
and ( n79725 , n79723 , n79724 );
and ( n79726 , n78620 , n78440 );
and ( n79727 , n79724 , n79726 );
and ( n79728 , n79723 , n79726 );
or ( n79729 , n79725 , n79727 , n79728 );
and ( n79730 , n79722 , n79729 );
xor ( n79731 , n79649 , n79650 );
xor ( n79732 , n79731 , n79652 );
and ( n79733 , n79729 , n79732 );
and ( n79734 , n79722 , n79732 );
or ( n79735 , n79730 , n79733 , n79734 );
and ( n79736 , n79721 , n79735 );
buf ( n79737 , n78528 );
xnor ( n79738 , n79623 , n79624 );
and ( n79739 , n79737 , n79738 );
xnor ( n79740 , n79687 , n79688 );
and ( n79741 , n79738 , n79740 );
and ( n79742 , n79737 , n79740 );
or ( n79743 , n79739 , n79741 , n79742 );
and ( n79744 , n79735 , n79743 );
and ( n79745 , n79721 , n79743 );
or ( n79746 , n79736 , n79744 , n79745 );
xor ( n79747 , n79644 , n79645 );
xor ( n79748 , n79747 , n79658 );
and ( n79749 , n79746 , n79748 );
and ( n79750 , n78843 , n78440 );
and ( n79751 , n78620 , n78519 );
and ( n79752 , n79750 , n79751 );
and ( n79753 , n78449 , n78855 );
and ( n79754 , n78528 , n78629 );
and ( n79755 , n79753 , n79754 );
and ( n79756 , n79752 , n79755 );
xor ( n79757 , n79723 , n79724 );
xor ( n79758 , n79757 , n79726 );
xor ( n79759 , n79681 , n79682 );
xor ( n79760 , n79759 , n79684 );
and ( n79761 , n79758 , n79760 );
and ( n79762 , n79756 , n79761 );
xor ( n79763 , n79722 , n79729 );
xor ( n79764 , n79763 , n79732 );
and ( n79765 , n79761 , n79764 );
and ( n79766 , n79756 , n79764 );
or ( n79767 , n79762 , n79765 , n79766 );
xor ( n79768 , n79647 , n79648 );
xor ( n79769 , n79752 , n79755 );
and ( n79770 , n79768 , n79769 );
xor ( n79771 , n79758 , n79760 );
and ( n79772 , n79769 , n79771 );
and ( n79773 , n79768 , n79771 );
or ( n79774 , n79770 , n79772 , n79773 );
xor ( n79775 , n79753 , n79754 );
and ( n79776 , n78541 , n78629 );
and ( n79777 , n78620 , n78516 );
and ( n79778 , n79776 , n79777 );
and ( n79779 , n79775 , n79778 );
and ( n79780 , n78336 , n78911 );
and ( n79781 , n79778 , n79780 );
and ( n79782 , n79775 , n79780 );
or ( n79783 , n79779 , n79781 , n79782 );
and ( n79784 , n78840 , n78345 );
not ( n79785 , n79784 );
xor ( n79786 , n79750 , n79751 );
and ( n79787 , n79785 , n79786 );
and ( n79788 , n79783 , n79787 );
buf ( n79789 , n79784 );
and ( n79790 , n79787 , n79789 );
and ( n79791 , n79783 , n79789 );
or ( n79792 , n79788 , n79790 , n79791 );
and ( n79793 , n79774 , n79792 );
xor ( n79794 , n79737 , n79738 );
xor ( n79795 , n79794 , n79740 );
and ( n79796 , n79792 , n79795 );
and ( n79797 , n79774 , n79795 );
or ( n79798 , n79793 , n79796 , n79797 );
and ( n79799 , n79767 , n79798 );
xor ( n79800 , n79689 , n79691 );
xor ( n79801 , n79800 , n79693 );
and ( n79802 , n79798 , n79801 );
and ( n79803 , n79767 , n79801 );
or ( n79804 , n79799 , n79802 , n79803 );
and ( n79805 , n79748 , n79804 );
and ( n79806 , n79746 , n79804 );
or ( n79807 , n79749 , n79805 , n79806 );
xor ( n79808 , n79674 , n79699 );
xor ( n79809 , n79808 , n79702 );
and ( n79810 , n79807 , n79809 );
xor ( n79811 , n79677 , n79679 );
xor ( n79812 , n79811 , n79696 );
xor ( n79813 , n79721 , n79735 );
xor ( n79814 , n79813 , n79743 );
and ( n79815 , n78840 , n78440 );
and ( n79816 , n78843 , n78519 );
and ( n79817 , n79815 , n79816 );
and ( n79818 , n78449 , n78911 );
and ( n79819 , n78528 , n78855 );
and ( n79820 , n79818 , n79819 );
and ( n79821 , n79817 , n79820 );
buf ( n79822 , n78541 );
xor ( n79823 , n79775 , n79778 );
xor ( n79824 , n79823 , n79780 );
and ( n79825 , n79822 , n79824 );
xor ( n79826 , n79785 , n79786 );
and ( n79827 , n79824 , n79826 );
and ( n79828 , n79822 , n79826 );
or ( n79829 , n79825 , n79827 , n79828 );
and ( n79830 , n79821 , n79829 );
xor ( n79831 , n79817 , n79820 );
and ( n79832 , n78840 , n78519 );
not ( n79833 , n79832 );
and ( n79834 , n78843 , n78516 );
and ( n79835 , n79833 , n79834 );
and ( n79836 , n78528 , n78911 );
not ( n79837 , n79836 );
and ( n79838 , n78541 , n78855 );
and ( n79839 , n79837 , n79838 );
and ( n79840 , n79835 , n79839 );
and ( n79841 , n79831 , n79840 );
buf ( n79842 , n79832 );
buf ( n79843 , n79836 );
and ( n79844 , n79842 , n79843 );
and ( n79845 , n79840 , n79844 );
and ( n79846 , n79831 , n79844 );
or ( n79847 , n79841 , n79845 , n79846 );
and ( n79848 , n79829 , n79847 );
and ( n79849 , n79821 , n79847 );
or ( n79850 , n79830 , n79848 , n79849 );
xor ( n79851 , n79756 , n79761 );
xor ( n79852 , n79851 , n79764 );
and ( n79853 , n79850 , n79852 );
xor ( n79854 , n79774 , n79792 );
xor ( n79855 , n79854 , n79795 );
and ( n79856 , n79852 , n79855 );
and ( n79857 , n79850 , n79855 );
or ( n79858 , n79853 , n79856 , n79857 );
and ( n79859 , n79814 , n79858 );
xor ( n79860 , n79767 , n79798 );
xor ( n79861 , n79860 , n79801 );
and ( n79862 , n79858 , n79861 );
and ( n79863 , n79814 , n79861 );
or ( n79864 , n79859 , n79862 , n79863 );
and ( n79865 , n79812 , n79864 );
xor ( n79866 , n79746 , n79748 );
xor ( n79867 , n79866 , n79804 );
and ( n79868 , n79864 , n79867 );
and ( n79869 , n79812 , n79867 );
or ( n79870 , n79865 , n79868 , n79869 );
and ( n79871 , n79809 , n79870 );
and ( n79872 , n79807 , n79870 );
or ( n79873 , n79810 , n79871 , n79872 );
and ( n79874 , n79720 , n79873 );
xor ( n79875 , n79807 , n79809 );
xor ( n79876 , n79875 , n79870 );
xor ( n79877 , n79812 , n79864 );
xor ( n79878 , n79877 , n79867 );
xor ( n79879 , n79814 , n79858 );
xor ( n79880 , n79879 , n79861 );
xor ( n79881 , n79768 , n79769 );
xor ( n79882 , n79881 , n79771 );
xor ( n79883 , n79783 , n79787 );
xor ( n79884 , n79883 , n79789 );
and ( n79885 , n79882 , n79884 );
xor ( n79886 , n79815 , n79816 );
xor ( n79887 , n79818 , n79819 );
and ( n79888 , n79886 , n79887 );
xor ( n79889 , n79776 , n79777 );
xor ( n79890 , n79835 , n79839 );
and ( n79891 , n79889 , n79890 );
xor ( n79892 , n79842 , n79843 );
and ( n79893 , n79890 , n79892 );
and ( n79894 , n79889 , n79892 );
or ( n79895 , n79891 , n79893 , n79894 );
and ( n79896 , n79888 , n79895 );
xor ( n79897 , n79886 , n79887 );
xor ( n79898 , n79833 , n79834 );
xor ( n79899 , n79837 , n79838 );
and ( n79900 , n79898 , n79899 );
and ( n79901 , n79897 , n79900 );
buf ( n79902 , n78620 );
and ( n79903 , n78541 , n78911 );
and ( n79904 , n78840 , n78516 );
and ( n79905 , n79903 , n79904 );
and ( n79906 , n79902 , n79905 );
and ( n79907 , n78620 , n78855 );
and ( n79908 , n78843 , n78629 );
and ( n79909 , n79907 , n79908 );
and ( n79910 , n79905 , n79909 );
and ( n79911 , n79902 , n79909 );
or ( n79912 , n79906 , n79910 , n79911 );
and ( n79913 , n79900 , n79912 );
and ( n79914 , n79897 , n79912 );
or ( n79915 , n79901 , n79913 , n79914 );
and ( n79916 , n79895 , n79915 );
and ( n79917 , n79888 , n79915 );
or ( n79918 , n79896 , n79916 , n79917 );
and ( n79919 , n79884 , n79918 );
and ( n79920 , n79882 , n79918 );
or ( n79921 , n79885 , n79919 , n79920 );
xor ( n79922 , n79850 , n79852 );
xor ( n79923 , n79922 , n79855 );
and ( n79924 , n79921 , n79923 );
xor ( n79925 , n79821 , n79829 );
xor ( n79926 , n79925 , n79847 );
xor ( n79927 , n79822 , n79824 );
xor ( n79928 , n79927 , n79826 );
xor ( n79929 , n79831 , n79840 );
xor ( n79930 , n79929 , n79844 );
and ( n79931 , n79928 , n79930 );
xor ( n79932 , n79888 , n79895 );
xor ( n79933 , n79932 , n79915 );
and ( n79934 , n79930 , n79933 );
and ( n79935 , n79928 , n79933 );
or ( n79936 , n79931 , n79934 , n79935 );
or ( n79937 , n79926 , n79936 );
and ( n79938 , n79923 , n79937 );
and ( n79939 , n79921 , n79937 );
or ( n79940 , n79924 , n79938 , n79939 );
or ( n79941 , n79880 , n79940 );
or ( n79942 , n79878 , n79941 );
or ( n79943 , n79876 , n79942 );
and ( n79944 , n79873 , n79943 );
and ( n79945 , n79720 , n79943 );
or ( n79946 , n79874 , n79944 , n79945 );
and ( n79947 , n79718 , n79946 );
xor ( n79948 , n79718 , n79946 );
xor ( n79949 , n79720 , n79873 );
xor ( n79950 , n79949 , n79943 );
xnor ( n79951 , n79876 , n79942 );
xnor ( n79952 , n79878 , n79941 );
xnor ( n79953 , n79880 , n79940 );
xor ( n79954 , n79921 , n79923 );
xor ( n79955 , n79954 , n79937 );
not ( n79956 , n79955 );
xor ( n79957 , n79882 , n79884 );
xor ( n79958 , n79957 , n79918 );
xnor ( n79959 , n79926 , n79936 );
and ( n79960 , n79958 , n79959 );
xor ( n79961 , n79958 , n79959 );
xor ( n79962 , n79889 , n79890 );
xor ( n79963 , n79962 , n79892 );
xor ( n79964 , n79897 , n79900 );
xor ( n79965 , n79964 , n79912 );
and ( n79966 , n79963 , n79965 );
xor ( n79967 , n79898 , n79899 );
xor ( n79968 , n79902 , n79905 );
xor ( n79969 , n79968 , n79909 );
and ( n79970 , n79967 , n79969 );
xor ( n79971 , n79903 , n79904 );
xor ( n79972 , n79907 , n79908 );
and ( n79973 , n79971 , n79972 );
and ( n79974 , n78843 , n78911 );
and ( n79975 , n78840 , n78855 );
and ( n79976 , n79974 , n79975 );
and ( n79977 , n78620 , n78911 );
and ( n79978 , n79976 , n79977 );
and ( n79979 , n79972 , n79978 );
and ( n79980 , n79971 , n79978 );
or ( n79981 , n79973 , n79979 , n79980 );
and ( n79982 , n79969 , n79981 );
and ( n79983 , n79967 , n79981 );
or ( n79984 , n79970 , n79982 , n79983 );
and ( n79985 , n79965 , n79984 );
and ( n79986 , n79963 , n79984 );
or ( n79987 , n79966 , n79985 , n79986 );
xor ( n79988 , n79928 , n79930 );
xor ( n79989 , n79988 , n79933 );
and ( n79990 , n79987 , n79989 );
xor ( n79991 , n79987 , n79989 );
xor ( n79992 , n79963 , n79965 );
xor ( n79993 , n79992 , n79984 );
not ( n79994 , n79993 );
xor ( n79995 , n79967 , n79969 );
xor ( n79996 , n79995 , n79981 );
and ( n79997 , n78840 , n78629 );
buf ( n79998 , n78843 );
and ( n79999 , n79997 , n79998 );
xor ( n80000 , n79976 , n79977 );
and ( n80001 , n79998 , n80000 );
and ( n80002 , n79997 , n80000 );
or ( n80003 , n79999 , n80001 , n80002 );
xor ( n80004 , n79971 , n79972 );
xor ( n80005 , n80004 , n79978 );
and ( n80006 , n80003 , n80005 );
and ( n80007 , n79996 , n80006 );
and ( n80008 , n79994 , n80007 );
or ( n80009 , n79993 , n80008 );
and ( n80010 , n79991 , n80009 );
or ( n80011 , n79990 , n80010 );
and ( n80012 , n79961 , n80011 );
or ( n80013 , n79960 , n80012 );
and ( n80014 , n79956 , n80013 );
or ( n80015 , n79955 , n80014 );
and ( n80016 , n79953 , n80015 );
and ( n80017 , n79952 , n80016 );
and ( n80018 , n79951 , n80017 );
and ( n80019 , n79950 , n80018 );
and ( n80020 , n79948 , n80019 );
or ( n80021 , n79947 , n80020 );
and ( n80022 , n79716 , n80021 );
or ( n80023 , n79715 , n80022 );
and ( n80024 , n79599 , n80023 );
and ( n80025 , n79597 , n80024 );
or ( n80026 , n79596 , n80025 );
and ( n80027 , n79539 , n80026 );
and ( n80028 , n79538 , n80027 );
or ( n80029 , n79537 , n80028 );
and ( n80030 , n79535 , n80029 );
and ( n80031 , n79534 , n80030 );
or ( n80032 , n79533 , n80031 );
and ( n80033 , n79531 , n80032 );
or ( n80034 , n79530 , n80033 );
and ( n80035 , n79165 , n80034 );
or ( n80036 , n79164 , n80035 );
and ( n80037 , n79162 , n80036 );
and ( n80038 , n79160 , n80037 );
and ( n80039 , n79159 , n80038 );
or ( n80040 , n79158 , n80039 );
and ( n80041 , n78702 , n80040 );
or ( n80042 , n78701 , n80041 );
and ( n80043 , n78699 , n80042 );
and ( n80044 , n78697 , n80043 );
and ( n80045 , n78695 , n80044 );
and ( n80046 , n78693 , n80045 );
or ( n80047 , n78692 , n80046 );
xor ( n80048 , n78690 , n80047 );
buf ( n80049 , n80048 );
buf ( n80050 , n80049 );
buf ( n80051 , n80050 );
buf ( n80052 , n560 );
buf ( n80053 , n576 );
and ( n80054 , n80052 , n80053 );
buf ( n80055 , n561 );
buf ( n80056 , n577 );
and ( n80057 , n80055 , n80056 );
buf ( n80058 , n562 );
buf ( n80059 , n578 );
and ( n80060 , n80058 , n80059 );
buf ( n80061 , n563 );
buf ( n80062 , n579 );
and ( n80063 , n80061 , n80062 );
buf ( n80064 , n564 );
buf ( n80065 , n580 );
and ( n80066 , n80064 , n80065 );
buf ( n80067 , n565 );
buf ( n80068 , n581 );
and ( n80069 , n80067 , n80068 );
buf ( n80070 , n566 );
buf ( n80071 , n582 );
and ( n80072 , n80070 , n80071 );
buf ( n80073 , n567 );
buf ( n80074 , n583 );
and ( n80075 , n80073 , n80074 );
buf ( n80076 , n568 );
buf ( n80077 , n584 );
and ( n80078 , n80076 , n80077 );
buf ( n80079 , n569 );
buf ( n80080 , n585 );
and ( n80081 , n80079 , n80080 );
buf ( n80082 , n570 );
buf ( n80083 , n586 );
and ( n80084 , n80082 , n80083 );
buf ( n80085 , n571 );
buf ( n80086 , n587 );
and ( n80087 , n80085 , n80086 );
buf ( n80088 , n572 );
buf ( n80089 , n588 );
and ( n80090 , n80088 , n80089 );
buf ( n80091 , n573 );
buf ( n80092 , n589 );
and ( n80093 , n80091 , n80092 );
buf ( n80094 , n574 );
buf ( n80095 , n590 );
and ( n80096 , n80094 , n80095 );
buf ( n80097 , n575 );
buf ( n80098 , n591 );
and ( n80099 , n80097 , n80098 );
and ( n80100 , n80095 , n80099 );
and ( n80101 , n80094 , n80099 );
or ( n80102 , n80096 , n80100 , n80101 );
and ( n80103 , n80092 , n80102 );
and ( n80104 , n80091 , n80102 );
or ( n80105 , n80093 , n80103 , n80104 );
and ( n80106 , n80089 , n80105 );
and ( n80107 , n80088 , n80105 );
or ( n80108 , n80090 , n80106 , n80107 );
and ( n80109 , n80086 , n80108 );
and ( n80110 , n80085 , n80108 );
or ( n80111 , n80087 , n80109 , n80110 );
and ( n80112 , n80083 , n80111 );
and ( n80113 , n80082 , n80111 );
or ( n80114 , n80084 , n80112 , n80113 );
and ( n80115 , n80080 , n80114 );
and ( n80116 , n80079 , n80114 );
or ( n80117 , n80081 , n80115 , n80116 );
and ( n80118 , n80077 , n80117 );
and ( n80119 , n80076 , n80117 );
or ( n80120 , n80078 , n80118 , n80119 );
and ( n80121 , n80074 , n80120 );
and ( n80122 , n80073 , n80120 );
or ( n80123 , n80075 , n80121 , n80122 );
and ( n80124 , n80071 , n80123 );
and ( n80125 , n80070 , n80123 );
or ( n80126 , n80072 , n80124 , n80125 );
and ( n80127 , n80068 , n80126 );
and ( n80128 , n80067 , n80126 );
or ( n80129 , n80069 , n80127 , n80128 );
and ( n80130 , n80065 , n80129 );
and ( n80131 , n80064 , n80129 );
or ( n80132 , n80066 , n80130 , n80131 );
and ( n80133 , n80062 , n80132 );
and ( n80134 , n80061 , n80132 );
or ( n80135 , n80063 , n80133 , n80134 );
and ( n80136 , n80059 , n80135 );
and ( n80137 , n80058 , n80135 );
or ( n80138 , n80060 , n80136 , n80137 );
and ( n80139 , n80056 , n80138 );
and ( n80140 , n80055 , n80138 );
or ( n80141 , n80057 , n80139 , n80140 );
and ( n80142 , n80053 , n80141 );
and ( n80143 , n80052 , n80141 );
or ( n80144 , n80054 , n80142 , n80143 );
buf ( n80145 , n80144 );
buf ( n80146 , n80145 );
buf ( n80147 , n80146 );
xor ( n80148 , n80052 , n80053 );
xor ( n80149 , n80148 , n80141 );
buf ( n80150 , n80149 );
buf ( n80151 , n80150 );
buf ( n80152 , n80151 );
xor ( n80153 , n80147 , n80152 );
not ( n80154 , n80153 );
and ( n80155 , n80147 , n80154 );
and ( n80156 , n80051 , n80155 );
xor ( n80157 , n80055 , n80056 );
xor ( n80158 , n80157 , n80138 );
buf ( n80159 , n80158 );
buf ( n80160 , n80159 );
buf ( n80161 , n80160 );
xor ( n80162 , n80152 , n80161 );
xor ( n80163 , n80058 , n80059 );
xor ( n80164 , n80163 , n80135 );
buf ( n80165 , n80164 );
buf ( n80166 , n80165 );
buf ( n80167 , n80166 );
xor ( n80168 , n80161 , n80167 );
not ( n80169 , n80168 );
and ( n80170 , n80162 , n80169 );
and ( n80171 , n80051 , n80170 );
not ( n80172 , n80171 );
and ( n80173 , n80161 , n80167 );
not ( n80174 , n80173 );
and ( n80175 , n80152 , n80174 );
xnor ( n80176 , n80172 , n80175 );
xor ( n80177 , n78695 , n80044 );
buf ( n80178 , n80177 );
buf ( n80179 , n80178 );
buf ( n80180 , n80179 );
and ( n80181 , n80180 , n80155 );
xor ( n80182 , n78693 , n80045 );
buf ( n80183 , n80182 );
buf ( n80184 , n80183 );
buf ( n80185 , n80184 );
and ( n80186 , n80185 , n80153 );
nor ( n80187 , n80181 , n80186 );
not ( n80188 , n80187 );
or ( n80189 , n80176 , n80188 );
not ( n80190 , n80175 );
and ( n80191 , n80189 , n80190 );
and ( n80192 , n80185 , n80155 );
and ( n80193 , n80051 , n80153 );
nor ( n80194 , n80192 , n80193 );
not ( n80195 , n80194 );
and ( n80196 , n80190 , n80195 );
and ( n80197 , n80189 , n80195 );
or ( n80198 , n80191 , n80196 , n80197 );
xnor ( n80199 , n80156 , n80198 );
xor ( n80200 , n80189 , n80190 );
xor ( n80201 , n80200 , n80195 );
xnor ( n80202 , n80176 , n80188 );
xor ( n80203 , n80061 , n80062 );
xor ( n80204 , n80203 , n80132 );
buf ( n80205 , n80204 );
buf ( n80206 , n80205 );
buf ( n80207 , n80206 );
xor ( n80208 , n80064 , n80065 );
xor ( n80209 , n80208 , n80129 );
buf ( n80210 , n80209 );
buf ( n80211 , n80210 );
buf ( n80212 , n80211 );
and ( n80213 , n80207 , n80212 );
not ( n80214 , n80213 );
and ( n80215 , n80167 , n80214 );
not ( n80216 , n80215 );
and ( n80217 , n80185 , n80170 );
and ( n80218 , n80051 , n80168 );
nor ( n80219 , n80217 , n80218 );
xnor ( n80220 , n80219 , n80175 );
and ( n80221 , n80216 , n80220 );
xor ( n80222 , n78697 , n80043 );
buf ( n80223 , n80222 );
buf ( n80224 , n80223 );
buf ( n80225 , n80224 );
and ( n80226 , n80225 , n80155 );
and ( n80227 , n80180 , n80153 );
nor ( n80228 , n80226 , n80227 );
not ( n80229 , n80228 );
and ( n80230 , n80220 , n80229 );
and ( n80231 , n80216 , n80229 );
or ( n80232 , n80221 , n80230 , n80231 );
and ( n80233 , n80202 , n80232 );
xor ( n80234 , n80167 , n80207 );
xor ( n80235 , n80207 , n80212 );
not ( n80236 , n80235 );
and ( n80237 , n80234 , n80236 );
and ( n80238 , n80051 , n80237 );
not ( n80239 , n80238 );
xnor ( n80240 , n80239 , n80215 );
xor ( n80241 , n78699 , n80042 );
buf ( n80242 , n80241 );
buf ( n80243 , n80242 );
buf ( n80244 , n80243 );
and ( n80245 , n80244 , n80155 );
and ( n80246 , n80225 , n80153 );
nor ( n80247 , n80245 , n80246 );
not ( n80248 , n80247 );
or ( n80249 , n80240 , n80248 );
xnor ( n80250 , n80240 , n80248 );
xor ( n80251 , n80067 , n80068 );
xor ( n80252 , n80251 , n80126 );
buf ( n80253 , n80252 );
buf ( n80254 , n80253 );
buf ( n80255 , n80254 );
xor ( n80256 , n80070 , n80071 );
xor ( n80257 , n80256 , n80123 );
buf ( n80258 , n80257 );
buf ( n80259 , n80258 );
buf ( n80260 , n80259 );
and ( n80261 , n80255 , n80260 );
not ( n80262 , n80261 );
and ( n80263 , n80212 , n80262 );
not ( n80264 , n80263 );
and ( n80265 , n80185 , n80237 );
and ( n80266 , n80051 , n80235 );
nor ( n80267 , n80265 , n80266 );
xnor ( n80268 , n80267 , n80215 );
and ( n80269 , n80264 , n80268 );
and ( n80270 , n80225 , n80170 );
and ( n80271 , n80180 , n80168 );
nor ( n80272 , n80270 , n80271 );
xnor ( n80273 , n80272 , n80175 );
and ( n80274 , n80268 , n80273 );
and ( n80275 , n80264 , n80273 );
or ( n80276 , n80269 , n80274 , n80275 );
and ( n80277 , n80250 , n80276 );
and ( n80278 , n80180 , n80170 );
and ( n80279 , n80185 , n80168 );
nor ( n80280 , n80278 , n80279 );
xnor ( n80281 , n80280 , n80175 );
and ( n80282 , n80276 , n80281 );
and ( n80283 , n80250 , n80281 );
or ( n80284 , n80277 , n80282 , n80283 );
and ( n80285 , n80249 , n80284 );
xor ( n80286 , n80216 , n80220 );
xor ( n80287 , n80286 , n80229 );
and ( n80288 , n80284 , n80287 );
and ( n80289 , n80249 , n80287 );
or ( n80290 , n80285 , n80288 , n80289 );
and ( n80291 , n80232 , n80290 );
and ( n80292 , n80202 , n80290 );
or ( n80293 , n80233 , n80291 , n80292 );
and ( n80294 , n80201 , n80293 );
xor ( n80295 , n80201 , n80293 );
xor ( n80296 , n80202 , n80232 );
xor ( n80297 , n80296 , n80290 );
xor ( n80298 , n80249 , n80284 );
xor ( n80299 , n80298 , n80287 );
xor ( n80300 , n80212 , n80255 );
xor ( n80301 , n80255 , n80260 );
not ( n80302 , n80301 );
and ( n80303 , n80300 , n80302 );
and ( n80304 , n80051 , n80303 );
not ( n80305 , n80304 );
xnor ( n80306 , n80305 , n80263 );
and ( n80307 , n80180 , n80237 );
and ( n80308 , n80185 , n80235 );
nor ( n80309 , n80307 , n80308 );
xnor ( n80310 , n80309 , n80215 );
or ( n80311 , n80306 , n80310 );
xor ( n80312 , n78702 , n80040 );
buf ( n80313 , n80312 );
buf ( n80314 , n80313 );
buf ( n80315 , n80314 );
and ( n80316 , n80315 , n80155 );
and ( n80317 , n80244 , n80153 );
nor ( n80318 , n80316 , n80317 );
not ( n80319 , n80318 );
and ( n80320 , n80311 , n80319 );
xor ( n80321 , n80264 , n80268 );
xor ( n80322 , n80321 , n80273 );
and ( n80323 , n80319 , n80322 );
and ( n80324 , n80311 , n80322 );
or ( n80325 , n80320 , n80323 , n80324 );
xor ( n80326 , n80073 , n80074 );
xor ( n80327 , n80326 , n80120 );
buf ( n80328 , n80327 );
buf ( n80329 , n80328 );
buf ( n80330 , n80329 );
xor ( n80331 , n80076 , n80077 );
xor ( n80332 , n80331 , n80117 );
buf ( n80333 , n80332 );
buf ( n80334 , n80333 );
buf ( n80335 , n80334 );
and ( n80336 , n80330 , n80335 );
not ( n80337 , n80336 );
and ( n80338 , n80260 , n80337 );
not ( n80339 , n80338 );
and ( n80340 , n80315 , n80170 );
and ( n80341 , n80244 , n80168 );
nor ( n80342 , n80340 , n80341 );
xnor ( n80343 , n80342 , n80175 );
and ( n80344 , n80339 , n80343 );
xor ( n80345 , n79160 , n80037 );
buf ( n80346 , n80345 );
buf ( n80347 , n80346 );
buf ( n80348 , n80347 );
and ( n80349 , n80348 , n80155 );
xor ( n80350 , n79159 , n80038 );
buf ( n80351 , n80350 );
buf ( n80352 , n80351 );
buf ( n80353 , n80352 );
and ( n80354 , n80353 , n80153 );
nor ( n80355 , n80349 , n80354 );
not ( n80356 , n80355 );
and ( n80357 , n80343 , n80356 );
and ( n80358 , n80339 , n80356 );
or ( n80359 , n80344 , n80357 , n80358 );
and ( n80360 , n80244 , n80170 );
and ( n80361 , n80225 , n80168 );
nor ( n80362 , n80360 , n80361 );
xnor ( n80363 , n80362 , n80175 );
and ( n80364 , n80359 , n80363 );
and ( n80365 , n80353 , n80155 );
and ( n80366 , n80315 , n80153 );
nor ( n80367 , n80365 , n80366 );
not ( n80368 , n80367 );
and ( n80369 , n80363 , n80368 );
and ( n80370 , n80359 , n80368 );
or ( n80371 , n80364 , n80369 , n80370 );
xnor ( n80372 , n80306 , n80310 );
xor ( n80373 , n80260 , n80330 );
xor ( n80374 , n80330 , n80335 );
not ( n80375 , n80374 );
and ( n80376 , n80373 , n80375 );
and ( n80377 , n80051 , n80376 );
not ( n80378 , n80377 );
xnor ( n80379 , n80378 , n80338 );
xor ( n80380 , n79162 , n80036 );
buf ( n80381 , n80380 );
buf ( n80382 , n80381 );
buf ( n80383 , n80382 );
and ( n80384 , n80383 , n80155 );
and ( n80385 , n80348 , n80153 );
nor ( n80386 , n80384 , n80385 );
not ( n80387 , n80386 );
or ( n80388 , n80379 , n80387 );
and ( n80389 , n80185 , n80303 );
and ( n80390 , n80051 , n80301 );
nor ( n80391 , n80389 , n80390 );
xnor ( n80392 , n80391 , n80263 );
and ( n80393 , n80388 , n80392 );
and ( n80394 , n80225 , n80237 );
and ( n80395 , n80180 , n80235 );
nor ( n80396 , n80394 , n80395 );
xnor ( n80397 , n80396 , n80215 );
and ( n80398 , n80392 , n80397 );
and ( n80399 , n80388 , n80397 );
or ( n80400 , n80393 , n80398 , n80399 );
and ( n80401 , n80372 , n80400 );
xor ( n80402 , n80359 , n80363 );
xor ( n80403 , n80402 , n80368 );
and ( n80404 , n80400 , n80403 );
and ( n80405 , n80372 , n80403 );
or ( n80406 , n80401 , n80404 , n80405 );
and ( n80407 , n80371 , n80406 );
xor ( n80408 , n80311 , n80319 );
xor ( n80409 , n80408 , n80322 );
and ( n80410 , n80406 , n80409 );
and ( n80411 , n80371 , n80409 );
or ( n80412 , n80407 , n80410 , n80411 );
and ( n80413 , n80325 , n80412 );
xor ( n80414 , n80250 , n80276 );
xor ( n80415 , n80414 , n80281 );
and ( n80416 , n80412 , n80415 );
and ( n80417 , n80325 , n80415 );
or ( n80418 , n80413 , n80416 , n80417 );
and ( n80419 , n80299 , n80418 );
xor ( n80420 , n80299 , n80418 );
xor ( n80421 , n80325 , n80412 );
xor ( n80422 , n80421 , n80415 );
xor ( n80423 , n80371 , n80406 );
xor ( n80424 , n80423 , n80409 );
and ( n80425 , n80180 , n80303 );
and ( n80426 , n80185 , n80301 );
nor ( n80427 , n80425 , n80426 );
xnor ( n80428 , n80427 , n80263 );
and ( n80429 , n80244 , n80237 );
and ( n80430 , n80225 , n80235 );
nor ( n80431 , n80429 , n80430 );
xnor ( n80432 , n80431 , n80215 );
and ( n80433 , n80428 , n80432 );
and ( n80434 , n80353 , n80170 );
and ( n80435 , n80315 , n80168 );
nor ( n80436 , n80434 , n80435 );
xnor ( n80437 , n80436 , n80175 );
and ( n80438 , n80432 , n80437 );
and ( n80439 , n80428 , n80437 );
or ( n80440 , n80433 , n80438 , n80439 );
xor ( n80441 , n80339 , n80343 );
xor ( n80442 , n80441 , n80356 );
and ( n80443 , n80440 , n80442 );
xor ( n80444 , n80388 , n80392 );
xor ( n80445 , n80444 , n80397 );
and ( n80446 , n80442 , n80445 );
and ( n80447 , n80440 , n80445 );
or ( n80448 , n80443 , n80446 , n80447 );
xnor ( n80449 , n80379 , n80387 );
xor ( n80450 , n80079 , n80080 );
xor ( n80451 , n80450 , n80114 );
buf ( n80452 , n80451 );
buf ( n80453 , n80452 );
buf ( n80454 , n80453 );
xor ( n80455 , n80082 , n80083 );
xor ( n80456 , n80455 , n80111 );
buf ( n80457 , n80456 );
buf ( n80458 , n80457 );
buf ( n80459 , n80458 );
and ( n80460 , n80454 , n80459 );
not ( n80461 , n80460 );
and ( n80462 , n80335 , n80461 );
not ( n80463 , n80462 );
and ( n80464 , n80225 , n80303 );
and ( n80465 , n80180 , n80301 );
nor ( n80466 , n80464 , n80465 );
xnor ( n80467 , n80466 , n80263 );
and ( n80468 , n80463 , n80467 );
xor ( n80469 , n79165 , n80034 );
buf ( n80470 , n80469 );
buf ( n80471 , n80470 );
buf ( n80472 , n80471 );
and ( n80473 , n80472 , n80155 );
and ( n80474 , n80383 , n80153 );
nor ( n80475 , n80473 , n80474 );
not ( n80476 , n80475 );
and ( n80477 , n80467 , n80476 );
and ( n80478 , n80463 , n80476 );
or ( n80479 , n80468 , n80477 , n80478 );
and ( n80480 , n80449 , n80479 );
and ( n80481 , n80185 , n80376 );
and ( n80482 , n80051 , n80374 );
nor ( n80483 , n80481 , n80482 );
xnor ( n80484 , n80483 , n80338 );
and ( n80485 , n80315 , n80237 );
and ( n80486 , n80244 , n80235 );
nor ( n80487 , n80485 , n80486 );
xnor ( n80488 , n80487 , n80215 );
and ( n80489 , n80484 , n80488 );
and ( n80490 , n80348 , n80170 );
and ( n80491 , n80353 , n80168 );
nor ( n80492 , n80490 , n80491 );
xnor ( n80493 , n80492 , n80175 );
and ( n80494 , n80488 , n80493 );
and ( n80495 , n80484 , n80493 );
or ( n80496 , n80489 , n80494 , n80495 );
and ( n80497 , n80479 , n80496 );
and ( n80498 , n80449 , n80496 );
or ( n80499 , n80480 , n80497 , n80498 );
xor ( n80500 , n80335 , n80454 );
xor ( n80501 , n80454 , n80459 );
not ( n80502 , n80501 );
and ( n80503 , n80500 , n80502 );
and ( n80504 , n80051 , n80503 );
not ( n80505 , n80504 );
xnor ( n80506 , n80505 , n80462 );
and ( n80507 , n80180 , n80376 );
and ( n80508 , n80185 , n80374 );
nor ( n80509 , n80507 , n80508 );
xnor ( n80510 , n80509 , n80338 );
and ( n80511 , n80506 , n80510 );
and ( n80512 , n80244 , n80303 );
and ( n80513 , n80225 , n80301 );
nor ( n80514 , n80512 , n80513 );
xnor ( n80515 , n80514 , n80263 );
and ( n80516 , n80510 , n80515 );
and ( n80517 , n80506 , n80515 );
or ( n80518 , n80511 , n80516 , n80517 );
and ( n80519 , n80383 , n80170 );
and ( n80520 , n80348 , n80168 );
nor ( n80521 , n80519 , n80520 );
xnor ( n80522 , n80521 , n80175 );
xor ( n80523 , n79531 , n80032 );
buf ( n80524 , n80523 );
buf ( n80525 , n80524 );
buf ( n80526 , n80525 );
and ( n80527 , n80526 , n80155 );
and ( n80528 , n80472 , n80153 );
nor ( n80529 , n80527 , n80528 );
not ( n80530 , n80529 );
or ( n80531 , n80522 , n80530 );
and ( n80532 , n80518 , n80531 );
xor ( n80533 , n80463 , n80467 );
xor ( n80534 , n80533 , n80476 );
and ( n80535 , n80531 , n80534 );
and ( n80536 , n80518 , n80534 );
or ( n80537 , n80532 , n80535 , n80536 );
xor ( n80538 , n80428 , n80432 );
xor ( n80539 , n80538 , n80437 );
and ( n80540 , n80537 , n80539 );
xor ( n80541 , n80449 , n80479 );
xor ( n80542 , n80541 , n80496 );
and ( n80543 , n80539 , n80542 );
and ( n80544 , n80537 , n80542 );
or ( n80545 , n80540 , n80543 , n80544 );
and ( n80546 , n80499 , n80545 );
xor ( n80547 , n80440 , n80442 );
xor ( n80548 , n80547 , n80445 );
and ( n80549 , n80545 , n80548 );
and ( n80550 , n80499 , n80548 );
or ( n80551 , n80546 , n80549 , n80550 );
and ( n80552 , n80448 , n80551 );
xor ( n80553 , n80372 , n80400 );
xor ( n80554 , n80553 , n80403 );
and ( n80555 , n80551 , n80554 );
and ( n80556 , n80448 , n80554 );
or ( n80557 , n80552 , n80555 , n80556 );
and ( n80558 , n80424 , n80557 );
xor ( n80559 , n80424 , n80557 );
xor ( n80560 , n80448 , n80551 );
xor ( n80561 , n80560 , n80554 );
xor ( n80562 , n80499 , n80545 );
xor ( n80563 , n80562 , n80548 );
xnor ( n80564 , n80522 , n80530 );
xor ( n80565 , n80085 , n80086 );
xor ( n80566 , n80565 , n80108 );
buf ( n80567 , n80566 );
buf ( n80568 , n80567 );
buf ( n80569 , n80568 );
xor ( n80570 , n80088 , n80089 );
xor ( n80571 , n80570 , n80105 );
buf ( n80572 , n80571 );
buf ( n80573 , n80572 );
buf ( n80574 , n80573 );
and ( n80575 , n80569 , n80574 );
not ( n80576 , n80575 );
and ( n80577 , n80459 , n80576 );
not ( n80578 , n80577 );
and ( n80579 , n80472 , n80170 );
and ( n80580 , n80383 , n80168 );
nor ( n80581 , n80579 , n80580 );
xnor ( n80582 , n80581 , n80175 );
and ( n80583 , n80578 , n80582 );
xor ( n80584 , n79534 , n80030 );
buf ( n80585 , n80584 );
buf ( n80586 , n80585 );
buf ( n80587 , n80586 );
and ( n80588 , n80587 , n80155 );
and ( n80589 , n80526 , n80153 );
nor ( n80590 , n80588 , n80589 );
not ( n80591 , n80590 );
and ( n80592 , n80582 , n80591 );
and ( n80593 , n80578 , n80591 );
or ( n80594 , n80583 , n80592 , n80593 );
and ( n80595 , n80564 , n80594 );
and ( n80596 , n80353 , n80237 );
and ( n80597 , n80315 , n80235 );
nor ( n80598 , n80596 , n80597 );
xnor ( n80599 , n80598 , n80215 );
and ( n80600 , n80594 , n80599 );
and ( n80601 , n80564 , n80599 );
or ( n80602 , n80595 , n80600 , n80601 );
xor ( n80603 , n80484 , n80488 );
xor ( n80604 , n80603 , n80493 );
and ( n80605 , n80602 , n80604 );
xor ( n80606 , n80518 , n80531 );
xor ( n80607 , n80606 , n80534 );
and ( n80608 , n80604 , n80607 );
and ( n80609 , n80602 , n80607 );
or ( n80610 , n80605 , n80608 , n80609 );
and ( n80611 , n80526 , n80170 );
and ( n80612 , n80472 , n80168 );
nor ( n80613 , n80611 , n80612 );
xnor ( n80614 , n80613 , n80175 );
xor ( n80615 , n79535 , n80029 );
buf ( n80616 , n80615 );
buf ( n80617 , n80616 );
buf ( n80618 , n80617 );
and ( n80619 , n80618 , n80155 );
and ( n80620 , n80587 , n80153 );
nor ( n80621 , n80619 , n80620 );
not ( n80622 , n80621 );
or ( n80623 , n80614 , n80622 );
and ( n80624 , n80185 , n80503 );
and ( n80625 , n80051 , n80501 );
nor ( n80626 , n80624 , n80625 );
xnor ( n80627 , n80626 , n80462 );
and ( n80628 , n80623 , n80627 );
and ( n80629 , n80225 , n80376 );
and ( n80630 , n80180 , n80374 );
nor ( n80631 , n80629 , n80630 );
xnor ( n80632 , n80631 , n80338 );
and ( n80633 , n80627 , n80632 );
and ( n80634 , n80623 , n80632 );
or ( n80635 , n80628 , n80633 , n80634 );
and ( n80636 , n80315 , n80303 );
and ( n80637 , n80244 , n80301 );
nor ( n80638 , n80636 , n80637 );
xnor ( n80639 , n80638 , n80263 );
and ( n80640 , n80348 , n80237 );
and ( n80641 , n80353 , n80235 );
nor ( n80642 , n80640 , n80641 );
xnor ( n80643 , n80642 , n80215 );
and ( n80644 , n80639 , n80643 );
xor ( n80645 , n80578 , n80582 );
xor ( n80646 , n80645 , n80591 );
and ( n80647 , n80643 , n80646 );
and ( n80648 , n80639 , n80646 );
or ( n80649 , n80644 , n80647 , n80648 );
and ( n80650 , n80635 , n80649 );
xor ( n80651 , n80506 , n80510 );
xor ( n80652 , n80651 , n80515 );
and ( n80653 , n80649 , n80652 );
and ( n80654 , n80635 , n80652 );
or ( n80655 , n80650 , n80653 , n80654 );
and ( n80656 , n80180 , n80503 );
and ( n80657 , n80185 , n80501 );
nor ( n80658 , n80656 , n80657 );
xnor ( n80659 , n80658 , n80462 );
and ( n80660 , n80244 , n80376 );
and ( n80661 , n80225 , n80374 );
nor ( n80662 , n80660 , n80661 );
xnor ( n80663 , n80662 , n80338 );
and ( n80664 , n80659 , n80663 );
and ( n80665 , n80353 , n80303 );
and ( n80666 , n80315 , n80301 );
nor ( n80667 , n80665 , n80666 );
xnor ( n80668 , n80667 , n80263 );
and ( n80669 , n80663 , n80668 );
and ( n80670 , n80659 , n80668 );
or ( n80671 , n80664 , n80669 , n80670 );
xor ( n80672 , n80091 , n80092 );
xor ( n80673 , n80672 , n80102 );
buf ( n80674 , n80673 );
buf ( n80675 , n80674 );
buf ( n80676 , n80675 );
xor ( n80677 , n80094 , n80095 );
xor ( n80678 , n80677 , n80099 );
buf ( n80679 , n80678 );
buf ( n80680 , n80679 );
buf ( n80681 , n80680 );
and ( n80682 , n80676 , n80681 );
not ( n80683 , n80682 );
and ( n80684 , n80574 , n80683 );
not ( n80685 , n80684 );
and ( n80686 , n80587 , n80170 );
and ( n80687 , n80526 , n80168 );
nor ( n80688 , n80686 , n80687 );
xnor ( n80689 , n80688 , n80175 );
and ( n80690 , n80685 , n80689 );
xor ( n80691 , n79538 , n80027 );
buf ( n80692 , n80691 );
buf ( n80693 , n80692 );
buf ( n80694 , n80693 );
and ( n80695 , n80694 , n80155 );
and ( n80696 , n80618 , n80153 );
nor ( n80697 , n80695 , n80696 );
not ( n80698 , n80697 );
and ( n80699 , n80689 , n80698 );
and ( n80700 , n80685 , n80698 );
or ( n80701 , n80690 , n80699 , n80700 );
xor ( n80702 , n80459 , n80569 );
xor ( n80703 , n80569 , n80574 );
not ( n80704 , n80703 );
and ( n80705 , n80702 , n80704 );
and ( n80706 , n80051 , n80705 );
not ( n80707 , n80706 );
xnor ( n80708 , n80707 , n80577 );
and ( n80709 , n80701 , n80708 );
and ( n80710 , n80383 , n80237 );
and ( n80711 , n80348 , n80235 );
nor ( n80712 , n80710 , n80711 );
xnor ( n80713 , n80712 , n80215 );
and ( n80714 , n80708 , n80713 );
and ( n80715 , n80701 , n80713 );
or ( n80716 , n80709 , n80714 , n80715 );
and ( n80717 , n80671 , n80716 );
xor ( n80718 , n80623 , n80627 );
xor ( n80719 , n80718 , n80632 );
and ( n80720 , n80716 , n80719 );
and ( n80721 , n80671 , n80719 );
or ( n80722 , n80717 , n80720 , n80721 );
xor ( n80723 , n80564 , n80594 );
xor ( n80724 , n80723 , n80599 );
and ( n80725 , n80722 , n80724 );
xor ( n80726 , n80635 , n80649 );
xor ( n80727 , n80726 , n80652 );
and ( n80728 , n80724 , n80727 );
and ( n80729 , n80722 , n80727 );
or ( n80730 , n80725 , n80728 , n80729 );
and ( n80731 , n80655 , n80730 );
xor ( n80732 , n80602 , n80604 );
xor ( n80733 , n80732 , n80607 );
and ( n80734 , n80730 , n80733 );
and ( n80735 , n80655 , n80733 );
or ( n80736 , n80731 , n80734 , n80735 );
and ( n80737 , n80610 , n80736 );
xor ( n80738 , n80537 , n80539 );
xor ( n80739 , n80738 , n80542 );
and ( n80740 , n80736 , n80739 );
and ( n80741 , n80610 , n80739 );
or ( n80742 , n80737 , n80740 , n80741 );
and ( n80743 , n80563 , n80742 );
xor ( n80744 , n80563 , n80742 );
xor ( n80745 , n80610 , n80736 );
xor ( n80746 , n80745 , n80739 );
xor ( n80747 , n80655 , n80730 );
xor ( n80748 , n80747 , n80733 );
xnor ( n80749 , n80614 , n80622 );
and ( n80750 , n80185 , n80705 );
and ( n80751 , n80051 , n80703 );
nor ( n80752 , n80750 , n80751 );
xnor ( n80753 , n80752 , n80577 );
and ( n80754 , n80225 , n80503 );
and ( n80755 , n80180 , n80501 );
nor ( n80756 , n80754 , n80755 );
xnor ( n80757 , n80756 , n80462 );
and ( n80758 , n80753 , n80757 );
and ( n80759 , n80348 , n80303 );
and ( n80760 , n80353 , n80301 );
nor ( n80761 , n80759 , n80760 );
xnor ( n80762 , n80761 , n80263 );
and ( n80763 , n80757 , n80762 );
and ( n80764 , n80753 , n80762 );
or ( n80765 , n80758 , n80763 , n80764 );
and ( n80766 , n80749 , n80765 );
and ( n80767 , n80618 , n80170 );
and ( n80768 , n80587 , n80168 );
nor ( n80769 , n80767 , n80768 );
xnor ( n80770 , n80769 , n80175 );
xor ( n80771 , n79539 , n80026 );
buf ( n80772 , n80771 );
buf ( n80773 , n80772 );
buf ( n80774 , n80773 );
and ( n80775 , n80774 , n80155 );
and ( n80776 , n80694 , n80153 );
nor ( n80777 , n80775 , n80776 );
not ( n80778 , n80777 );
or ( n80779 , n80770 , n80778 );
and ( n80780 , n80315 , n80376 );
and ( n80781 , n80244 , n80374 );
nor ( n80782 , n80780 , n80781 );
xnor ( n80783 , n80782 , n80338 );
and ( n80784 , n80779 , n80783 );
and ( n80785 , n80472 , n80237 );
and ( n80786 , n80383 , n80235 );
nor ( n80787 , n80785 , n80786 );
xnor ( n80788 , n80787 , n80215 );
and ( n80789 , n80783 , n80788 );
and ( n80790 , n80779 , n80788 );
or ( n80791 , n80784 , n80789 , n80790 );
and ( n80792 , n80765 , n80791 );
and ( n80793 , n80749 , n80791 );
or ( n80794 , n80766 , n80792 , n80793 );
xor ( n80795 , n80639 , n80643 );
xor ( n80796 , n80795 , n80646 );
and ( n80797 , n80794 , n80796 );
xor ( n80798 , n80671 , n80716 );
xor ( n80799 , n80798 , n80719 );
and ( n80800 , n80796 , n80799 );
and ( n80801 , n80794 , n80799 );
or ( n80802 , n80797 , n80800 , n80801 );
xor ( n80803 , n80574 , n80676 );
xor ( n80804 , n80676 , n80681 );
not ( n80805 , n80804 );
and ( n80806 , n80803 , n80805 );
and ( n80807 , n80051 , n80806 );
not ( n80808 , n80807 );
xnor ( n80809 , n80808 , n80684 );
and ( n80810 , n80383 , n80303 );
and ( n80811 , n80348 , n80301 );
nor ( n80812 , n80810 , n80811 );
xnor ( n80813 , n80812 , n80263 );
and ( n80814 , n80809 , n80813 );
and ( n80815 , n80526 , n80237 );
and ( n80816 , n80472 , n80235 );
nor ( n80817 , n80815 , n80816 );
xnor ( n80818 , n80817 , n80215 );
and ( n80819 , n80813 , n80818 );
and ( n80820 , n80809 , n80818 );
or ( n80821 , n80814 , n80819 , n80820 );
not ( n80822 , n80681 );
xor ( n80823 , n79597 , n80024 );
buf ( n80824 , n80823 );
buf ( n80825 , n80824 );
buf ( n80826 , n80825 );
and ( n80827 , n80826 , n80155 );
and ( n80828 , n80774 , n80153 );
nor ( n80829 , n80827 , n80828 );
not ( n80830 , n80829 );
or ( n80831 , n80822 , n80830 );
and ( n80832 , n80180 , n80705 );
and ( n80833 , n80185 , n80703 );
nor ( n80834 , n80832 , n80833 );
xnor ( n80835 , n80834 , n80577 );
and ( n80836 , n80831 , n80835 );
and ( n80837 , n80353 , n80376 );
and ( n80838 , n80315 , n80374 );
nor ( n80839 , n80837 , n80838 );
xnor ( n80840 , n80839 , n80338 );
and ( n80841 , n80835 , n80840 );
and ( n80842 , n80831 , n80840 );
or ( n80843 , n80836 , n80841 , n80842 );
and ( n80844 , n80821 , n80843 );
xor ( n80845 , n80685 , n80689 );
xor ( n80846 , n80845 , n80698 );
and ( n80847 , n80843 , n80846 );
and ( n80848 , n80821 , n80846 );
or ( n80849 , n80844 , n80847 , n80848 );
xor ( n80850 , n80659 , n80663 );
xor ( n80851 , n80850 , n80668 );
and ( n80852 , n80849 , n80851 );
xor ( n80853 , n80701 , n80708 );
xor ( n80854 , n80853 , n80713 );
and ( n80855 , n80851 , n80854 );
and ( n80856 , n80849 , n80854 );
or ( n80857 , n80852 , n80855 , n80856 );
xnor ( n80858 , n80770 , n80778 );
and ( n80859 , n80472 , n80303 );
and ( n80860 , n80383 , n80301 );
nor ( n80861 , n80859 , n80860 );
xnor ( n80862 , n80861 , n80263 );
and ( n80863 , n80587 , n80237 );
and ( n80864 , n80526 , n80235 );
nor ( n80865 , n80863 , n80864 );
xnor ( n80866 , n80865 , n80215 );
and ( n80867 , n80862 , n80866 );
and ( n80868 , n80694 , n80170 );
and ( n80869 , n80618 , n80168 );
nor ( n80870 , n80868 , n80869 );
xnor ( n80871 , n80870 , n80175 );
and ( n80872 , n80866 , n80871 );
and ( n80873 , n80862 , n80871 );
or ( n80874 , n80867 , n80872 , n80873 );
and ( n80875 , n80858 , n80874 );
and ( n80876 , n80244 , n80503 );
and ( n80877 , n80225 , n80501 );
nor ( n80878 , n80876 , n80877 );
xnor ( n80879 , n80878 , n80462 );
and ( n80880 , n80874 , n80879 );
and ( n80881 , n80858 , n80879 );
or ( n80882 , n80875 , n80880 , n80881 );
xor ( n80883 , n80753 , n80757 );
xor ( n80884 , n80883 , n80762 );
and ( n80885 , n80882 , n80884 );
xor ( n80886 , n80779 , n80783 );
xor ( n80887 , n80886 , n80788 );
and ( n80888 , n80884 , n80887 );
and ( n80889 , n80882 , n80887 );
or ( n80890 , n80885 , n80888 , n80889 );
xor ( n80891 , n80749 , n80765 );
xor ( n80892 , n80891 , n80791 );
and ( n80893 , n80890 , n80892 );
xor ( n80894 , n80849 , n80851 );
xor ( n80895 , n80894 , n80854 );
and ( n80896 , n80892 , n80895 );
and ( n80897 , n80890 , n80895 );
or ( n80898 , n80893 , n80896 , n80897 );
and ( n80899 , n80857 , n80898 );
xor ( n80900 , n80794 , n80796 );
xor ( n80901 , n80900 , n80799 );
and ( n80902 , n80898 , n80901 );
and ( n80903 , n80857 , n80901 );
or ( n80904 , n80899 , n80902 , n80903 );
and ( n80905 , n80802 , n80904 );
xor ( n80906 , n80722 , n80724 );
xor ( n80907 , n80906 , n80727 );
and ( n80908 , n80904 , n80907 );
and ( n80909 , n80802 , n80907 );
or ( n80910 , n80905 , n80908 , n80909 );
and ( n80911 , n80748 , n80910 );
xor ( n80912 , n80748 , n80910 );
xor ( n80913 , n80802 , n80904 );
xor ( n80914 , n80913 , n80907 );
xor ( n80915 , n80857 , n80898 );
xor ( n80916 , n80915 , n80901 );
and ( n80917 , n80526 , n80303 );
and ( n80918 , n80472 , n80301 );
nor ( n80919 , n80917 , n80918 );
xnor ( n80920 , n80919 , n80263 );
and ( n80921 , n80774 , n80170 );
and ( n80922 , n80694 , n80168 );
nor ( n80923 , n80921 , n80922 );
xnor ( n80924 , n80923 , n80175 );
and ( n80925 , n80920 , n80924 );
xor ( n80926 , n79599 , n80023 );
buf ( n80927 , n80926 );
buf ( n80928 , n80927 );
buf ( n80929 , n80928 );
and ( n80930 , n80929 , n80155 );
and ( n80931 , n80826 , n80153 );
nor ( n80932 , n80930 , n80931 );
not ( n80933 , n80932 );
and ( n80934 , n80924 , n80933 );
and ( n80935 , n80920 , n80933 );
or ( n80936 , n80925 , n80934 , n80935 );
and ( n80937 , n80185 , n80806 );
and ( n80938 , n80051 , n80804 );
nor ( n80939 , n80937 , n80938 );
xnor ( n80940 , n80939 , n80684 );
and ( n80941 , n80936 , n80940 );
and ( n80942 , n80225 , n80705 );
and ( n80943 , n80180 , n80703 );
nor ( n80944 , n80942 , n80943 );
xnor ( n80945 , n80944 , n80577 );
and ( n80946 , n80940 , n80945 );
and ( n80947 , n80936 , n80945 );
or ( n80948 , n80941 , n80946 , n80947 );
xnor ( n80949 , n80822 , n80830 );
and ( n80950 , n80315 , n80503 );
and ( n80951 , n80244 , n80501 );
nor ( n80952 , n80950 , n80951 );
xnor ( n80953 , n80952 , n80462 );
and ( n80954 , n80949 , n80953 );
and ( n80955 , n80348 , n80376 );
and ( n80956 , n80353 , n80374 );
nor ( n80957 , n80955 , n80956 );
xnor ( n80958 , n80957 , n80338 );
and ( n80959 , n80953 , n80958 );
and ( n80960 , n80949 , n80958 );
or ( n80961 , n80954 , n80959 , n80960 );
and ( n80962 , n80948 , n80961 );
xor ( n80963 , n80809 , n80813 );
xor ( n80964 , n80963 , n80818 );
and ( n80965 , n80961 , n80964 );
and ( n80966 , n80948 , n80964 );
or ( n80967 , n80962 , n80965 , n80966 );
xor ( n80968 , n80821 , n80843 );
xor ( n80969 , n80968 , n80846 );
and ( n80970 , n80967 , n80969 );
xor ( n80971 , n80882 , n80884 );
xor ( n80972 , n80971 , n80887 );
and ( n80973 , n80969 , n80972 );
and ( n80974 , n80967 , n80972 );
or ( n80975 , n80970 , n80973 , n80974 );
and ( n80976 , n80180 , n80806 );
and ( n80977 , n80185 , n80804 );
nor ( n80978 , n80976 , n80977 );
xnor ( n80979 , n80978 , n80684 );
and ( n80980 , n80353 , n80503 );
and ( n80981 , n80315 , n80501 );
nor ( n80982 , n80980 , n80981 );
xnor ( n80983 , n80982 , n80462 );
and ( n80984 , n80979 , n80983 );
and ( n80985 , n80383 , n80376 );
and ( n80986 , n80348 , n80374 );
nor ( n80987 , n80985 , n80986 );
xnor ( n80988 , n80987 , n80338 );
and ( n80989 , n80983 , n80988 );
and ( n80990 , n80979 , n80988 );
or ( n80991 , n80984 , n80989 , n80990 );
and ( n80992 , n80826 , n80170 );
and ( n80993 , n80774 , n80168 );
nor ( n80994 , n80992 , n80993 );
xnor ( n80995 , n80994 , n80175 );
xor ( n80996 , n79716 , n80021 );
buf ( n80997 , n80996 );
buf ( n80998 , n80997 );
buf ( n80999 , n80998 );
and ( n81000 , n80999 , n80155 );
and ( n81001 , n80929 , n80153 );
nor ( n81002 , n81000 , n81001 );
not ( n81003 , n81002 );
and ( n81004 , n80995 , n81003 );
xor ( n81005 , n80097 , n80098 );
buf ( n81006 , n81005 );
buf ( n81007 , n81006 );
buf ( n81008 , n81007 );
xor ( n81009 , n80681 , n81008 );
not ( n81010 , n81008 );
and ( n81011 , n81009 , n81010 );
and ( n81012 , n80051 , n81011 );
not ( n81013 , n81012 );
xnor ( n81014 , n81013 , n80681 );
and ( n81015 , n81004 , n81014 );
and ( n81016 , n80618 , n80237 );
and ( n81017 , n80587 , n80235 );
nor ( n81018 , n81016 , n81017 );
xnor ( n81019 , n81018 , n80215 );
and ( n81020 , n81014 , n81019 );
and ( n81021 , n81004 , n81019 );
or ( n81022 , n81015 , n81020 , n81021 );
and ( n81023 , n80991 , n81022 );
xor ( n81024 , n80862 , n80866 );
xor ( n81025 , n81024 , n80871 );
and ( n81026 , n81022 , n81025 );
and ( n81027 , n80991 , n81025 );
or ( n81028 , n81023 , n81026 , n81027 );
xor ( n81029 , n80831 , n80835 );
xor ( n81030 , n81029 , n80840 );
and ( n81031 , n81028 , n81030 );
xor ( n81032 , n80858 , n80874 );
xor ( n81033 , n81032 , n80879 );
and ( n81034 , n81030 , n81033 );
and ( n81035 , n81028 , n81033 );
or ( n81036 , n81031 , n81034 , n81035 );
xor ( n81037 , n80995 , n81003 );
and ( n81038 , n80587 , n80303 );
and ( n81039 , n80526 , n80301 );
nor ( n81040 , n81038 , n81039 );
xnor ( n81041 , n81040 , n80263 );
and ( n81042 , n81037 , n81041 );
and ( n81043 , n80694 , n80237 );
and ( n81044 , n80618 , n80235 );
nor ( n81045 , n81043 , n81044 );
xnor ( n81046 , n81045 , n80215 );
and ( n81047 , n81041 , n81046 );
and ( n81048 , n81037 , n81046 );
or ( n81049 , n81042 , n81047 , n81048 );
and ( n81050 , n80244 , n80705 );
and ( n81051 , n80225 , n80703 );
nor ( n81052 , n81050 , n81051 );
xnor ( n81053 , n81052 , n80577 );
and ( n81054 , n81049 , n81053 );
xor ( n81055 , n80920 , n80924 );
xor ( n81056 , n81055 , n80933 );
and ( n81057 , n81053 , n81056 );
and ( n81058 , n81049 , n81056 );
or ( n81059 , n81054 , n81057 , n81058 );
xor ( n81060 , n80936 , n80940 );
xor ( n81061 , n81060 , n80945 );
and ( n81062 , n81059 , n81061 );
xor ( n81063 , n80949 , n80953 );
xor ( n81064 , n81063 , n80958 );
and ( n81065 , n81061 , n81064 );
and ( n81066 , n81059 , n81064 );
or ( n81067 , n81062 , n81065 , n81066 );
xor ( n81068 , n80948 , n80961 );
xor ( n81069 , n81068 , n80964 );
and ( n81070 , n81067 , n81069 );
xor ( n81071 , n81028 , n81030 );
xor ( n81072 , n81071 , n81033 );
and ( n81073 , n81069 , n81072 );
and ( n81074 , n81067 , n81072 );
or ( n81075 , n81070 , n81073 , n81074 );
and ( n81076 , n81036 , n81075 );
xor ( n81077 , n80967 , n80969 );
xor ( n81078 , n81077 , n80972 );
and ( n81079 , n81075 , n81078 );
and ( n81080 , n81036 , n81078 );
or ( n81081 , n81076 , n81079 , n81080 );
and ( n81082 , n80975 , n81081 );
xor ( n81083 , n80890 , n80892 );
xor ( n81084 , n81083 , n80895 );
and ( n81085 , n81081 , n81084 );
and ( n81086 , n80975 , n81084 );
or ( n81087 , n81082 , n81085 , n81086 );
and ( n81088 , n80916 , n81087 );
xor ( n81089 , n80916 , n81087 );
xor ( n81090 , n80975 , n81081 );
xor ( n81091 , n81090 , n81084 );
xor ( n81092 , n81036 , n81075 );
xor ( n81093 , n81092 , n81078 );
and ( n81094 , n80526 , n80376 );
and ( n81095 , n80472 , n80374 );
nor ( n81096 , n81094 , n81095 );
xnor ( n81097 , n81096 , n80338 );
and ( n81098 , n80618 , n80303 );
and ( n81099 , n80587 , n80301 );
nor ( n81100 , n81098 , n81099 );
xnor ( n81101 , n81100 , n80263 );
and ( n81102 , n81097 , n81101 );
and ( n81103 , n80774 , n80237 );
and ( n81104 , n80694 , n80235 );
nor ( n81105 , n81103 , n81104 );
xnor ( n81106 , n81105 , n80215 );
and ( n81107 , n81101 , n81106 );
and ( n81108 , n81097 , n81106 );
or ( n81109 , n81102 , n81107 , n81108 );
and ( n81110 , n80185 , n81011 );
and ( n81111 , n80051 , n81008 );
nor ( n81112 , n81110 , n81111 );
xnor ( n81113 , n81112 , n80681 );
and ( n81114 , n81109 , n81113 );
and ( n81115 , n80315 , n80705 );
and ( n81116 , n80244 , n80703 );
nor ( n81117 , n81115 , n81116 );
xnor ( n81118 , n81117 , n80577 );
and ( n81119 , n81113 , n81118 );
and ( n81120 , n81109 , n81118 );
or ( n81121 , n81114 , n81119 , n81120 );
and ( n81122 , n80999 , n80170 );
and ( n81123 , n80929 , n80168 );
nor ( n81124 , n81122 , n81123 );
xnor ( n81125 , n81124 , n80175 );
xor ( n81126 , n79950 , n80018 );
buf ( n81127 , n81126 );
buf ( n81128 , n81127 );
buf ( n81129 , n81128 );
and ( n81130 , n81129 , n80155 );
xor ( n81131 , n79948 , n80019 );
buf ( n81132 , n81131 );
buf ( n81133 , n81132 );
buf ( n81134 , n81133 );
and ( n81135 , n81134 , n80153 );
nor ( n81136 , n81130 , n81135 );
not ( n81137 , n81136 );
and ( n81138 , n81125 , n81137 );
and ( n81139 , n80929 , n80170 );
and ( n81140 , n80826 , n80168 );
nor ( n81141 , n81139 , n81140 );
xnor ( n81142 , n81141 , n80175 );
and ( n81143 , n81138 , n81142 );
and ( n81144 , n81134 , n80155 );
and ( n81145 , n80999 , n80153 );
nor ( n81146 , n81144 , n81145 );
not ( n81147 , n81146 );
and ( n81148 , n81142 , n81147 );
and ( n81149 , n81138 , n81147 );
or ( n81150 , n81143 , n81148 , n81149 );
and ( n81151 , n80225 , n80806 );
and ( n81152 , n80180 , n80804 );
nor ( n81153 , n81151 , n81152 );
xnor ( n81154 , n81153 , n80684 );
and ( n81155 , n81150 , n81154 );
and ( n81156 , n80472 , n80376 );
and ( n81157 , n80383 , n80374 );
nor ( n81158 , n81156 , n81157 );
xnor ( n81159 , n81158 , n80338 );
and ( n81160 , n81154 , n81159 );
and ( n81161 , n81150 , n81159 );
or ( n81162 , n81155 , n81160 , n81161 );
and ( n81163 , n81121 , n81162 );
xor ( n81164 , n81004 , n81014 );
xor ( n81165 , n81164 , n81019 );
and ( n81166 , n81162 , n81165 );
and ( n81167 , n81121 , n81165 );
or ( n81168 , n81163 , n81166 , n81167 );
xor ( n81169 , n80991 , n81022 );
xor ( n81170 , n81169 , n81025 );
and ( n81171 , n81168 , n81170 );
xor ( n81172 , n81059 , n81061 );
xor ( n81173 , n81172 , n81064 );
and ( n81174 , n81170 , n81173 );
and ( n81175 , n81168 , n81173 );
or ( n81176 , n81171 , n81174 , n81175 );
and ( n81177 , n80348 , n80503 );
and ( n81178 , n80353 , n80501 );
nor ( n81179 , n81177 , n81178 );
xnor ( n81180 , n81179 , n80462 );
xor ( n81181 , n81150 , n81154 );
xor ( n81182 , n81181 , n81159 );
and ( n81183 , n81180 , n81182 );
xor ( n81184 , n81037 , n81041 );
xor ( n81185 , n81184 , n81046 );
and ( n81186 , n81182 , n81185 );
and ( n81187 , n81180 , n81185 );
or ( n81188 , n81183 , n81186 , n81187 );
xor ( n81189 , n80979 , n80983 );
xor ( n81190 , n81189 , n80988 );
and ( n81191 , n81188 , n81190 );
xor ( n81192 , n81049 , n81053 );
xor ( n81193 , n81192 , n81056 );
and ( n81194 , n81190 , n81193 );
and ( n81195 , n81188 , n81193 );
or ( n81196 , n81191 , n81194 , n81195 );
xor ( n81197 , n81125 , n81137 );
and ( n81198 , n80587 , n80376 );
and ( n81199 , n80526 , n80374 );
nor ( n81200 , n81198 , n81199 );
xnor ( n81201 , n81200 , n80338 );
and ( n81202 , n81197 , n81201 );
and ( n81203 , n80826 , n80237 );
and ( n81204 , n80774 , n80235 );
nor ( n81205 , n81203 , n81204 );
xnor ( n81206 , n81205 , n80215 );
and ( n81207 , n81201 , n81206 );
and ( n81208 , n81197 , n81206 );
or ( n81209 , n81202 , n81207 , n81208 );
and ( n81210 , n80180 , n81011 );
and ( n81211 , n80185 , n81008 );
nor ( n81212 , n81210 , n81211 );
xnor ( n81213 , n81212 , n80681 );
and ( n81214 , n81209 , n81213 );
and ( n81215 , n80353 , n80705 );
and ( n81216 , n80315 , n80703 );
nor ( n81217 , n81215 , n81216 );
xnor ( n81218 , n81217 , n80577 );
and ( n81219 , n81213 , n81218 );
and ( n81220 , n81209 , n81218 );
or ( n81221 , n81214 , n81219 , n81220 );
and ( n81222 , n80244 , n80806 );
and ( n81223 , n80225 , n80804 );
nor ( n81224 , n81222 , n81223 );
xnor ( n81225 , n81224 , n80684 );
and ( n81226 , n80383 , n80503 );
and ( n81227 , n80348 , n80501 );
nor ( n81228 , n81226 , n81227 );
xnor ( n81229 , n81228 , n80462 );
and ( n81230 , n81225 , n81229 );
xor ( n81231 , n81138 , n81142 );
xor ( n81232 , n81231 , n81147 );
and ( n81233 , n81229 , n81232 );
and ( n81234 , n81225 , n81232 );
or ( n81235 , n81230 , n81233 , n81234 );
and ( n81236 , n81221 , n81235 );
xor ( n81237 , n81109 , n81113 );
xor ( n81238 , n81237 , n81118 );
and ( n81239 , n81235 , n81238 );
and ( n81240 , n81221 , n81238 );
or ( n81241 , n81236 , n81239 , n81240 );
xor ( n81242 , n81121 , n81162 );
xor ( n81243 , n81242 , n81165 );
and ( n81244 , n81241 , n81243 );
xor ( n81245 , n81188 , n81190 );
xor ( n81246 , n81245 , n81193 );
and ( n81247 , n81243 , n81246 );
and ( n81248 , n81241 , n81246 );
or ( n81249 , n81244 , n81247 , n81248 );
and ( n81250 , n81196 , n81249 );
xor ( n81251 , n81168 , n81170 );
xor ( n81252 , n81251 , n81173 );
and ( n81253 , n81249 , n81252 );
and ( n81254 , n81196 , n81252 );
or ( n81255 , n81250 , n81253 , n81254 );
and ( n81256 , n81176 , n81255 );
xor ( n81257 , n81067 , n81069 );
xor ( n81258 , n81257 , n81072 );
and ( n81259 , n81255 , n81258 );
and ( n81260 , n81176 , n81258 );
or ( n81261 , n81256 , n81259 , n81260 );
and ( n81262 , n81093 , n81261 );
xor ( n81263 , n81093 , n81261 );
xor ( n81264 , n81176 , n81255 );
xor ( n81265 , n81264 , n81258 );
xor ( n81266 , n81196 , n81249 );
xor ( n81267 , n81266 , n81252 );
and ( n81268 , n81129 , n80170 );
and ( n81269 , n81134 , n80168 );
nor ( n81270 , n81268 , n81269 );
xnor ( n81271 , n81270 , n80175 );
xor ( n81272 , n79952 , n80016 );
buf ( n81273 , n81272 );
buf ( n81274 , n81273 );
buf ( n81275 , n81274 );
and ( n81276 , n81275 , n80155 );
xor ( n81277 , n79951 , n80017 );
buf ( n81278 , n81277 );
buf ( n81279 , n81278 );
buf ( n81280 , n81279 );
and ( n81281 , n81280 , n80153 );
nor ( n81282 , n81276 , n81281 );
not ( n81283 , n81282 );
and ( n81284 , n81271 , n81283 );
and ( n81285 , n81134 , n80170 );
and ( n81286 , n80999 , n80168 );
nor ( n81287 , n81285 , n81286 );
xnor ( n81288 , n81287 , n80175 );
and ( n81289 , n81284 , n81288 );
and ( n81290 , n81280 , n80155 );
and ( n81291 , n81129 , n80153 );
nor ( n81292 , n81290 , n81291 );
not ( n81293 , n81292 );
and ( n81294 , n81288 , n81293 );
and ( n81295 , n81284 , n81293 );
or ( n81296 , n81289 , n81294 , n81295 );
and ( n81297 , n80472 , n80503 );
and ( n81298 , n80383 , n80501 );
nor ( n81299 , n81297 , n81298 );
xnor ( n81300 , n81299 , n80462 );
and ( n81301 , n81296 , n81300 );
and ( n81302 , n80694 , n80303 );
and ( n81303 , n80618 , n80301 );
nor ( n81304 , n81302 , n81303 );
xnor ( n81305 , n81304 , n80263 );
and ( n81306 , n81300 , n81305 );
and ( n81307 , n81296 , n81305 );
or ( n81308 , n81301 , n81306 , n81307 );
xor ( n81309 , n81097 , n81101 );
xor ( n81310 , n81309 , n81106 );
and ( n81311 , n81308 , n81310 );
xor ( n81312 , n81225 , n81229 );
xor ( n81313 , n81312 , n81232 );
and ( n81314 , n81310 , n81313 );
and ( n81315 , n81308 , n81313 );
or ( n81316 , n81311 , n81314 , n81315 );
xor ( n81317 , n81180 , n81182 );
xor ( n81318 , n81317 , n81185 );
and ( n81319 , n81316 , n81318 );
xor ( n81320 , n81221 , n81235 );
xor ( n81321 , n81320 , n81238 );
and ( n81322 , n81318 , n81321 );
and ( n81323 , n81316 , n81321 );
or ( n81324 , n81319 , n81322 , n81323 );
and ( n81325 , n80774 , n80303 );
and ( n81326 , n80694 , n80301 );
nor ( n81327 , n81325 , n81326 );
xnor ( n81328 , n81327 , n80263 );
and ( n81329 , n80929 , n80237 );
and ( n81330 , n80826 , n80235 );
nor ( n81331 , n81329 , n81330 );
xnor ( n81332 , n81331 , n80215 );
and ( n81333 , n81328 , n81332 );
xor ( n81334 , n81284 , n81288 );
xor ( n81335 , n81334 , n81293 );
and ( n81336 , n81332 , n81335 );
and ( n81337 , n81328 , n81335 );
or ( n81338 , n81333 , n81336 , n81337 );
and ( n81339 , n80225 , n81011 );
and ( n81340 , n80180 , n81008 );
nor ( n81341 , n81339 , n81340 );
xnor ( n81342 , n81341 , n80681 );
and ( n81343 , n81338 , n81342 );
and ( n81344 , n80315 , n80806 );
and ( n81345 , n80244 , n80804 );
nor ( n81346 , n81344 , n81345 );
xnor ( n81347 , n81346 , n80684 );
and ( n81348 , n81342 , n81347 );
and ( n81349 , n81338 , n81347 );
or ( n81350 , n81343 , n81348 , n81349 );
xor ( n81351 , n81271 , n81283 );
and ( n81352 , n81134 , n80237 );
and ( n81353 , n80999 , n80235 );
nor ( n81354 , n81352 , n81353 );
xnor ( n81355 , n81354 , n80215 );
and ( n81356 , n81280 , n80170 );
and ( n81357 , n81129 , n80168 );
nor ( n81358 , n81356 , n81357 );
xnor ( n81359 , n81358 , n80175 );
and ( n81360 , n81355 , n81359 );
xor ( n81361 , n79953 , n80015 );
buf ( n81362 , n81361 );
buf ( n81363 , n81362 );
buf ( n81364 , n81363 );
and ( n81365 , n81364 , n80155 );
and ( n81366 , n81275 , n80153 );
nor ( n81367 , n81365 , n81366 );
not ( n81368 , n81367 );
and ( n81369 , n81359 , n81368 );
and ( n81370 , n81355 , n81368 );
or ( n81371 , n81360 , n81369 , n81370 );
and ( n81372 , n81351 , n81371 );
and ( n81373 , n80999 , n80237 );
and ( n81374 , n80929 , n80235 );
nor ( n81375 , n81373 , n81374 );
xnor ( n81376 , n81375 , n80215 );
and ( n81377 , n81371 , n81376 );
and ( n81378 , n81351 , n81376 );
or ( n81379 , n81372 , n81377 , n81378 );
and ( n81380 , n80526 , n80503 );
and ( n81381 , n80472 , n80501 );
nor ( n81382 , n81380 , n81381 );
xnor ( n81383 , n81382 , n80462 );
and ( n81384 , n81379 , n81383 );
and ( n81385 , n80618 , n80376 );
and ( n81386 , n80587 , n80374 );
nor ( n81387 , n81385 , n81386 );
xnor ( n81388 , n81387 , n80338 );
and ( n81389 , n81383 , n81388 );
and ( n81390 , n81379 , n81388 );
or ( n81391 , n81384 , n81389 , n81390 );
and ( n81392 , n80348 , n80705 );
and ( n81393 , n80353 , n80703 );
nor ( n81394 , n81392 , n81393 );
xnor ( n81395 , n81394 , n80577 );
and ( n81396 , n81391 , n81395 );
xor ( n81397 , n81197 , n81201 );
xor ( n81398 , n81397 , n81206 );
and ( n81399 , n81395 , n81398 );
and ( n81400 , n81391 , n81398 );
or ( n81401 , n81396 , n81399 , n81400 );
and ( n81402 , n81350 , n81401 );
xor ( n81403 , n81209 , n81213 );
xor ( n81404 , n81403 , n81218 );
and ( n81405 , n81401 , n81404 );
and ( n81406 , n81350 , n81404 );
or ( n81407 , n81402 , n81405 , n81406 );
and ( n81408 , n80244 , n81011 );
and ( n81409 , n80225 , n81008 );
nor ( n81410 , n81408 , n81409 );
xnor ( n81411 , n81410 , n80681 );
and ( n81412 , n80383 , n80705 );
and ( n81413 , n80348 , n80703 );
nor ( n81414 , n81412 , n81413 );
xnor ( n81415 , n81414 , n80577 );
and ( n81416 , n81411 , n81415 );
xor ( n81417 , n81328 , n81332 );
xor ( n81418 , n81417 , n81335 );
and ( n81419 , n81415 , n81418 );
and ( n81420 , n81411 , n81418 );
or ( n81421 , n81416 , n81419 , n81420 );
xor ( n81422 , n81296 , n81300 );
xor ( n81423 , n81422 , n81305 );
and ( n81424 , n81421 , n81423 );
xor ( n81425 , n81338 , n81342 );
xor ( n81426 , n81425 , n81347 );
and ( n81427 , n81423 , n81426 );
and ( n81428 , n81421 , n81426 );
or ( n81429 , n81424 , n81427 , n81428 );
xor ( n81430 , n81350 , n81401 );
xor ( n81431 , n81430 , n81404 );
and ( n81432 , n81429 , n81431 );
xor ( n81433 , n81308 , n81310 );
xor ( n81434 , n81433 , n81313 );
and ( n81435 , n81431 , n81434 );
and ( n81436 , n81429 , n81434 );
or ( n81437 , n81432 , n81435 , n81436 );
and ( n81438 , n81407 , n81437 );
xor ( n81439 , n81316 , n81318 );
xor ( n81440 , n81439 , n81321 );
and ( n81441 , n81437 , n81440 );
and ( n81442 , n81407 , n81440 );
or ( n81443 , n81438 , n81441 , n81442 );
and ( n81444 , n81324 , n81443 );
xor ( n81445 , n81241 , n81243 );
xor ( n81446 , n81445 , n81246 );
and ( n81447 , n81443 , n81446 );
and ( n81448 , n81324 , n81446 );
or ( n81449 , n81444 , n81447 , n81448 );
and ( n81450 , n81267 , n81449 );
xor ( n81451 , n81267 , n81449 );
xor ( n81452 , n81324 , n81443 );
xor ( n81453 , n81452 , n81446 );
xor ( n81454 , n81407 , n81437 );
xor ( n81455 , n81454 , n81440 );
and ( n81456 , n80587 , n80503 );
and ( n81457 , n80526 , n80501 );
nor ( n81458 , n81456 , n81457 );
xnor ( n81459 , n81458 , n80462 );
and ( n81460 , n80694 , n80376 );
and ( n81461 , n80618 , n80374 );
nor ( n81462 , n81460 , n81461 );
xnor ( n81463 , n81462 , n80338 );
and ( n81464 , n81459 , n81463 );
and ( n81465 , n80826 , n80303 );
and ( n81466 , n80774 , n80301 );
nor ( n81467 , n81465 , n81466 );
xnor ( n81468 , n81467 , n80263 );
and ( n81469 , n81463 , n81468 );
and ( n81470 , n81459 , n81468 );
or ( n81471 , n81464 , n81469 , n81470 );
and ( n81472 , n80353 , n80806 );
and ( n81473 , n80315 , n80804 );
nor ( n81474 , n81472 , n81473 );
xnor ( n81475 , n81474 , n80684 );
and ( n81476 , n81471 , n81475 );
xor ( n81477 , n81379 , n81383 );
xor ( n81478 , n81477 , n81388 );
and ( n81479 , n81475 , n81478 );
and ( n81480 , n81471 , n81478 );
or ( n81481 , n81476 , n81479 , n81480 );
xor ( n81482 , n81391 , n81395 );
xor ( n81483 , n81482 , n81398 );
and ( n81484 , n81481 , n81483 );
xor ( n81485 , n81421 , n81423 );
xor ( n81486 , n81485 , n81426 );
and ( n81487 , n81483 , n81486 );
and ( n81488 , n81481 , n81486 );
or ( n81489 , n81484 , n81487 , n81488 );
and ( n81490 , n81275 , n80170 );
and ( n81491 , n81280 , n80168 );
nor ( n81492 , n81490 , n81491 );
xnor ( n81493 , n81492 , n80175 );
xor ( n81494 , n79956 , n80013 );
buf ( n81495 , n81494 );
buf ( n81496 , n81495 );
buf ( n81497 , n81496 );
and ( n81498 , n81497 , n80155 );
and ( n81499 , n81364 , n80153 );
nor ( n81500 , n81498 , n81499 );
not ( n81501 , n81500 );
xor ( n81502 , n81493 , n81501 );
and ( n81503 , n80999 , n80303 );
and ( n81504 , n80929 , n80301 );
nor ( n81505 , n81503 , n81504 );
xnor ( n81506 , n81505 , n80263 );
and ( n81507 , n81502 , n81506 );
and ( n81508 , n81129 , n80237 );
and ( n81509 , n81134 , n80235 );
nor ( n81510 , n81508 , n81509 );
xnor ( n81511 , n81510 , n80215 );
and ( n81512 , n81506 , n81511 );
and ( n81513 , n81502 , n81511 );
or ( n81514 , n81507 , n81512 , n81513 );
and ( n81515 , n80526 , n80705 );
and ( n81516 , n80472 , n80703 );
nor ( n81517 , n81515 , n81516 );
xnor ( n81518 , n81517 , n80577 );
and ( n81519 , n81514 , n81518 );
and ( n81520 , n80774 , n80376 );
and ( n81521 , n80694 , n80374 );
nor ( n81522 , n81520 , n81521 );
xnor ( n81523 , n81522 , n80338 );
and ( n81524 , n81518 , n81523 );
and ( n81525 , n81514 , n81523 );
or ( n81526 , n81519 , n81524 , n81525 );
and ( n81527 , n80315 , n81011 );
and ( n81528 , n80244 , n81008 );
nor ( n81529 , n81527 , n81528 );
xnor ( n81530 , n81529 , n80681 );
and ( n81531 , n81526 , n81530 );
and ( n81532 , n80348 , n80806 );
and ( n81533 , n80353 , n80804 );
nor ( n81534 , n81532 , n81533 );
xnor ( n81535 , n81534 , n80684 );
and ( n81536 , n81530 , n81535 );
and ( n81537 , n81526 , n81535 );
or ( n81538 , n81531 , n81536 , n81537 );
and ( n81539 , n81493 , n81501 );
and ( n81540 , n80929 , n80303 );
and ( n81541 , n80826 , n80301 );
nor ( n81542 , n81540 , n81541 );
xnor ( n81543 , n81542 , n80263 );
and ( n81544 , n81539 , n81543 );
xor ( n81545 , n81355 , n81359 );
xor ( n81546 , n81545 , n81368 );
and ( n81547 , n81543 , n81546 );
and ( n81548 , n81539 , n81546 );
or ( n81549 , n81544 , n81547 , n81548 );
and ( n81550 , n80472 , n80705 );
and ( n81551 , n80383 , n80703 );
nor ( n81552 , n81550 , n81551 );
xnor ( n81553 , n81552 , n80577 );
and ( n81554 , n81549 , n81553 );
xor ( n81555 , n81351 , n81371 );
xor ( n81556 , n81555 , n81376 );
and ( n81557 , n81553 , n81556 );
and ( n81558 , n81549 , n81556 );
or ( n81559 , n81554 , n81557 , n81558 );
and ( n81560 , n81538 , n81559 );
xor ( n81561 , n81411 , n81415 );
xor ( n81562 , n81561 , n81418 );
and ( n81563 , n81559 , n81562 );
and ( n81564 , n81538 , n81562 );
or ( n81565 , n81560 , n81563 , n81564 );
and ( n81566 , n80383 , n80806 );
and ( n81567 , n80348 , n80804 );
nor ( n81568 , n81566 , n81567 );
xnor ( n81569 , n81568 , n80684 );
and ( n81570 , n80618 , n80503 );
and ( n81571 , n80587 , n80501 );
nor ( n81572 , n81570 , n81571 );
xnor ( n81573 , n81572 , n80462 );
and ( n81574 , n81569 , n81573 );
xor ( n81575 , n81539 , n81543 );
xor ( n81576 , n81575 , n81546 );
and ( n81577 , n81573 , n81576 );
and ( n81578 , n81569 , n81576 );
or ( n81579 , n81574 , n81577 , n81578 );
xor ( n81580 , n81459 , n81463 );
xor ( n81581 , n81580 , n81468 );
and ( n81582 , n81579 , n81581 );
xor ( n81583 , n81549 , n81553 );
xor ( n81584 , n81583 , n81556 );
and ( n81585 , n81581 , n81584 );
and ( n81586 , n81579 , n81584 );
or ( n81587 , n81582 , n81585 , n81586 );
xor ( n81588 , n81471 , n81475 );
xor ( n81589 , n81588 , n81478 );
and ( n81590 , n81587 , n81589 );
xor ( n81591 , n81538 , n81559 );
xor ( n81592 , n81591 , n81562 );
and ( n81593 , n81589 , n81592 );
and ( n81594 , n81587 , n81592 );
or ( n81595 , n81590 , n81593 , n81594 );
and ( n81596 , n81565 , n81595 );
xor ( n81597 , n81481 , n81483 );
xor ( n81598 , n81597 , n81486 );
and ( n81599 , n81595 , n81598 );
and ( n81600 , n81565 , n81598 );
or ( n81601 , n81596 , n81599 , n81600 );
and ( n81602 , n81489 , n81601 );
xor ( n81603 , n81429 , n81431 );
xor ( n81604 , n81603 , n81434 );
and ( n81605 , n81601 , n81604 );
and ( n81606 , n81489 , n81604 );
or ( n81607 , n81602 , n81605 , n81606 );
and ( n81608 , n81455 , n81607 );
xor ( n81609 , n81455 , n81607 );
xor ( n81610 , n81489 , n81601 );
xor ( n81611 , n81610 , n81604 );
xor ( n81612 , n81565 , n81595 );
xor ( n81613 , n81612 , n81598 );
and ( n81614 , n81280 , n80237 );
and ( n81615 , n81129 , n80235 );
nor ( n81616 , n81614 , n81615 );
xnor ( n81617 , n81616 , n80215 );
and ( n81618 , n81364 , n80170 );
and ( n81619 , n81275 , n80168 );
nor ( n81620 , n81618 , n81619 );
xnor ( n81621 , n81620 , n80175 );
and ( n81622 , n81617 , n81621 );
xor ( n81623 , n79961 , n80011 );
buf ( n81624 , n81623 );
buf ( n81625 , n81624 );
buf ( n81626 , n81625 );
and ( n81627 , n81626 , n80155 );
and ( n81628 , n81497 , n80153 );
nor ( n81629 , n81627 , n81628 );
not ( n81630 , n81629 );
and ( n81631 , n81621 , n81630 );
and ( n81632 , n81617 , n81630 );
or ( n81633 , n81622 , n81631 , n81632 );
and ( n81634 , n81497 , n80170 );
and ( n81635 , n81364 , n80168 );
nor ( n81636 , n81634 , n81635 );
xnor ( n81637 , n81636 , n80175 );
xor ( n81638 , n79991 , n80009 );
buf ( n81639 , n81638 );
buf ( n81640 , n81639 );
buf ( n81641 , n81640 );
and ( n81642 , n81641 , n80155 );
and ( n81643 , n81626 , n80153 );
nor ( n81644 , n81642 , n81643 );
not ( n81645 , n81644 );
and ( n81646 , n81637 , n81645 );
and ( n81647 , n81134 , n80303 );
and ( n81648 , n80999 , n80301 );
nor ( n81649 , n81647 , n81648 );
xnor ( n81650 , n81649 , n80263 );
and ( n81651 , n81646 , n81650 );
xor ( n81652 , n81617 , n81621 );
xor ( n81653 , n81652 , n81630 );
and ( n81654 , n81650 , n81653 );
and ( n81655 , n81646 , n81653 );
or ( n81656 , n81651 , n81654 , n81655 );
and ( n81657 , n81633 , n81656 );
and ( n81658 , n80826 , n80376 );
and ( n81659 , n80774 , n80374 );
nor ( n81660 , n81658 , n81659 );
xnor ( n81661 , n81660 , n80338 );
and ( n81662 , n81656 , n81661 );
and ( n81663 , n81633 , n81661 );
or ( n81664 , n81657 , n81662 , n81663 );
and ( n81665 , n80587 , n80705 );
and ( n81666 , n80526 , n80703 );
nor ( n81667 , n81665 , n81666 );
xnor ( n81668 , n81667 , n80577 );
and ( n81669 , n80694 , n80503 );
and ( n81670 , n80618 , n80501 );
nor ( n81671 , n81669 , n81670 );
xnor ( n81672 , n81671 , n80462 );
and ( n81673 , n81668 , n81672 );
xor ( n81674 , n81502 , n81506 );
xor ( n81675 , n81674 , n81511 );
and ( n81676 , n81672 , n81675 );
and ( n81677 , n81668 , n81675 );
or ( n81678 , n81673 , n81676 , n81677 );
and ( n81679 , n81664 , n81678 );
and ( n81680 , n80353 , n81011 );
and ( n81681 , n80315 , n81008 );
nor ( n81682 , n81680 , n81681 );
xnor ( n81683 , n81682 , n80681 );
and ( n81684 , n81678 , n81683 );
and ( n81685 , n81664 , n81683 );
or ( n81686 , n81679 , n81684 , n81685 );
xor ( n81687 , n81526 , n81530 );
xor ( n81688 , n81687 , n81535 );
and ( n81689 , n81686 , n81688 );
xor ( n81690 , n81579 , n81581 );
xor ( n81691 , n81690 , n81584 );
and ( n81692 , n81688 , n81691 );
and ( n81693 , n81686 , n81691 );
or ( n81694 , n81689 , n81692 , n81693 );
xor ( n81695 , n81637 , n81645 );
and ( n81696 , n81641 , n80170 );
and ( n81697 , n81626 , n80168 );
nor ( n81698 , n81696 , n81697 );
xnor ( n81699 , n81698 , n80175 );
xor ( n81700 , n79996 , n80006 );
buf ( n81701 , n81700 );
buf ( n81702 , n81701 );
buf ( n81703 , n81702 );
and ( n81704 , n81703 , n80155 );
xor ( n81705 , n79994 , n80007 );
buf ( n81706 , n81705 );
buf ( n81707 , n81706 );
buf ( n81708 , n81707 );
and ( n81709 , n81708 , n80153 );
nor ( n81710 , n81704 , n81709 );
not ( n81711 , n81710 );
and ( n81712 , n81699 , n81711 );
and ( n81713 , n81626 , n80170 );
and ( n81714 , n81497 , n80168 );
nor ( n81715 , n81713 , n81714 );
xnor ( n81716 , n81715 , n80175 );
and ( n81717 , n81712 , n81716 );
and ( n81718 , n81708 , n80155 );
and ( n81719 , n81641 , n80153 );
nor ( n81720 , n81718 , n81719 );
not ( n81721 , n81720 );
and ( n81722 , n81716 , n81721 );
and ( n81723 , n81712 , n81721 );
or ( n81724 , n81717 , n81722 , n81723 );
and ( n81725 , n81695 , n81724 );
and ( n81726 , n81275 , n80237 );
and ( n81727 , n81280 , n80235 );
nor ( n81728 , n81726 , n81727 );
xnor ( n81729 , n81728 , n80215 );
and ( n81730 , n81724 , n81729 );
and ( n81731 , n81695 , n81729 );
or ( n81732 , n81725 , n81730 , n81731 );
and ( n81733 , n80774 , n80503 );
and ( n81734 , n80694 , n80501 );
nor ( n81735 , n81733 , n81734 );
xnor ( n81736 , n81735 , n80462 );
and ( n81737 , n81732 , n81736 );
and ( n81738 , n80929 , n80376 );
and ( n81739 , n80826 , n80374 );
nor ( n81740 , n81738 , n81739 );
xnor ( n81741 , n81740 , n80338 );
and ( n81742 , n81736 , n81741 );
and ( n81743 , n81732 , n81741 );
or ( n81744 , n81737 , n81742 , n81743 );
and ( n81745 , n80472 , n80806 );
and ( n81746 , n80383 , n80804 );
nor ( n81747 , n81745 , n81746 );
xnor ( n81748 , n81747 , n80684 );
and ( n81749 , n81744 , n81748 );
xor ( n81750 , n81633 , n81656 );
xor ( n81751 , n81750 , n81661 );
and ( n81752 , n81748 , n81751 );
and ( n81753 , n81744 , n81751 );
or ( n81754 , n81749 , n81752 , n81753 );
xor ( n81755 , n81514 , n81518 );
xor ( n81756 , n81755 , n81523 );
and ( n81757 , n81754 , n81756 );
xor ( n81758 , n81569 , n81573 );
xor ( n81759 , n81758 , n81576 );
and ( n81760 , n81756 , n81759 );
and ( n81761 , n81754 , n81759 );
or ( n81762 , n81757 , n81760 , n81761 );
and ( n81763 , n81280 , n80303 );
and ( n81764 , n81129 , n80301 );
nor ( n81765 , n81763 , n81764 );
xnor ( n81766 , n81765 , n80263 );
and ( n81767 , n81364 , n80237 );
and ( n81768 , n81275 , n80235 );
nor ( n81769 , n81767 , n81768 );
xnor ( n81770 , n81769 , n80215 );
and ( n81771 , n81766 , n81770 );
xor ( n81772 , n81712 , n81716 );
xor ( n81773 , n81772 , n81721 );
and ( n81774 , n81770 , n81773 );
and ( n81775 , n81766 , n81773 );
or ( n81776 , n81771 , n81774 , n81775 );
and ( n81777 , n80999 , n80376 );
and ( n81778 , n80929 , n80374 );
nor ( n81779 , n81777 , n81778 );
xnor ( n81780 , n81779 , n80338 );
and ( n81781 , n81776 , n81780 );
and ( n81782 , n81129 , n80303 );
and ( n81783 , n81134 , n80301 );
nor ( n81784 , n81782 , n81783 );
xnor ( n81785 , n81784 , n80263 );
and ( n81786 , n81780 , n81785 );
and ( n81787 , n81776 , n81785 );
or ( n81788 , n81781 , n81786 , n81787 );
and ( n81789 , n80526 , n80806 );
and ( n81790 , n80472 , n80804 );
nor ( n81791 , n81789 , n81790 );
xnor ( n81792 , n81791 , n80684 );
and ( n81793 , n81788 , n81792 );
xor ( n81794 , n81646 , n81650 );
xor ( n81795 , n81794 , n81653 );
and ( n81796 , n81792 , n81795 );
and ( n81797 , n81788 , n81795 );
or ( n81798 , n81793 , n81796 , n81797 );
and ( n81799 , n80348 , n81011 );
and ( n81800 , n80353 , n81008 );
nor ( n81801 , n81799 , n81800 );
xnor ( n81802 , n81801 , n80681 );
and ( n81803 , n81798 , n81802 );
xor ( n81804 , n81668 , n81672 );
xor ( n81805 , n81804 , n81675 );
and ( n81806 , n81802 , n81805 );
and ( n81807 , n81798 , n81805 );
or ( n81808 , n81803 , n81806 , n81807 );
xor ( n81809 , n81664 , n81678 );
xor ( n81810 , n81809 , n81683 );
and ( n81811 , n81808 , n81810 );
xor ( n81812 , n81754 , n81756 );
xor ( n81813 , n81812 , n81759 );
and ( n81814 , n81810 , n81813 );
and ( n81815 , n81808 , n81813 );
or ( n81816 , n81811 , n81814 , n81815 );
and ( n81817 , n81762 , n81816 );
xor ( n81818 , n81686 , n81688 );
xor ( n81819 , n81818 , n81691 );
and ( n81820 , n81816 , n81819 );
and ( n81821 , n81762 , n81819 );
or ( n81822 , n81817 , n81820 , n81821 );
and ( n81823 , n81694 , n81822 );
xor ( n81824 , n81587 , n81589 );
xor ( n81825 , n81824 , n81592 );
and ( n81826 , n81822 , n81825 );
and ( n81827 , n81694 , n81825 );
or ( n81828 , n81823 , n81826 , n81827 );
and ( n81829 , n81613 , n81828 );
xor ( n81830 , n81613 , n81828 );
xor ( n81831 , n81694 , n81822 );
xor ( n81832 , n81831 , n81825 );
xor ( n81833 , n81762 , n81816 );
xor ( n81834 , n81833 , n81819 );
and ( n81835 , n80383 , n81011 );
and ( n81836 , n80348 , n81008 );
nor ( n81837 , n81835 , n81836 );
xnor ( n81838 , n81837 , n80681 );
and ( n81839 , n80618 , n80705 );
and ( n81840 , n80587 , n80703 );
nor ( n81841 , n81839 , n81840 );
xnor ( n81842 , n81841 , n80577 );
and ( n81843 , n81838 , n81842 );
xor ( n81844 , n81732 , n81736 );
xor ( n81845 , n81844 , n81741 );
and ( n81846 , n81842 , n81845 );
and ( n81847 , n81838 , n81845 );
or ( n81848 , n81843 , n81846 , n81847 );
xor ( n81849 , n81744 , n81748 );
xor ( n81850 , n81849 , n81751 );
and ( n81851 , n81848 , n81850 );
xor ( n81852 , n81798 , n81802 );
xor ( n81853 , n81852 , n81805 );
and ( n81854 , n81850 , n81853 );
and ( n81855 , n81848 , n81853 );
or ( n81856 , n81851 , n81854 , n81855 );
and ( n81857 , n80587 , n80806 );
and ( n81858 , n80526 , n80804 );
nor ( n81859 , n81857 , n81858 );
xnor ( n81860 , n81859 , n80684 );
and ( n81861 , n80826 , n80503 );
and ( n81862 , n80774 , n80501 );
nor ( n81863 , n81861 , n81862 );
xnor ( n81864 , n81863 , n80462 );
and ( n81865 , n81860 , n81864 );
xor ( n81866 , n81695 , n81724 );
xor ( n81867 , n81866 , n81729 );
and ( n81868 , n81864 , n81867 );
and ( n81869 , n81860 , n81867 );
or ( n81870 , n81865 , n81868 , n81869 );
xor ( n81871 , n81699 , n81711 );
and ( n81872 , n81626 , n80237 );
and ( n81873 , n81497 , n80235 );
nor ( n81874 , n81872 , n81873 );
xnor ( n81875 , n81874 , n80215 );
and ( n81876 , n81708 , n80170 );
and ( n81877 , n81641 , n80168 );
nor ( n81878 , n81876 , n81877 );
xnor ( n81879 , n81878 , n80175 );
and ( n81880 , n81875 , n81879 );
xor ( n81881 , n80003 , n80005 );
buf ( n81882 , n81881 );
buf ( n81883 , n81882 );
buf ( n81884 , n81883 );
and ( n81885 , n81884 , n80155 );
and ( n81886 , n81703 , n80153 );
nor ( n81887 , n81885 , n81886 );
not ( n81888 , n81887 );
and ( n81889 , n81879 , n81888 );
and ( n81890 , n81875 , n81888 );
or ( n81891 , n81880 , n81889 , n81890 );
and ( n81892 , n81871 , n81891 );
and ( n81893 , n81497 , n80237 );
and ( n81894 , n81364 , n80235 );
nor ( n81895 , n81893 , n81894 );
xnor ( n81896 , n81895 , n80215 );
and ( n81897 , n81891 , n81896 );
and ( n81898 , n81871 , n81896 );
or ( n81899 , n81892 , n81897 , n81898 );
and ( n81900 , n80929 , n80503 );
and ( n81901 , n80826 , n80501 );
nor ( n81902 , n81900 , n81901 );
xnor ( n81903 , n81902 , n80462 );
and ( n81904 , n81899 , n81903 );
and ( n81905 , n81134 , n80376 );
and ( n81906 , n80999 , n80374 );
nor ( n81907 , n81905 , n81906 );
xnor ( n81908 , n81907 , n80338 );
and ( n81909 , n81903 , n81908 );
and ( n81910 , n81899 , n81908 );
or ( n81911 , n81904 , n81909 , n81910 );
and ( n81912 , n80694 , n80705 );
and ( n81913 , n80618 , n80703 );
nor ( n81914 , n81912 , n81913 );
xnor ( n81915 , n81914 , n80577 );
and ( n81916 , n81911 , n81915 );
xor ( n81917 , n81776 , n81780 );
xor ( n81918 , n81917 , n81785 );
and ( n81919 , n81915 , n81918 );
and ( n81920 , n81911 , n81918 );
or ( n81921 , n81916 , n81919 , n81920 );
and ( n81922 , n81870 , n81921 );
xor ( n81923 , n81788 , n81792 );
xor ( n81924 , n81923 , n81795 );
and ( n81925 , n81921 , n81924 );
and ( n81926 , n81870 , n81924 );
or ( n81927 , n81922 , n81925 , n81926 );
and ( n81928 , n81129 , n80376 );
and ( n81929 , n81134 , n80374 );
nor ( n81930 , n81928 , n81929 );
xnor ( n81931 , n81930 , n80338 );
and ( n81932 , n81275 , n80303 );
and ( n81933 , n81280 , n80301 );
nor ( n81934 , n81932 , n81933 );
xnor ( n81935 , n81934 , n80263 );
and ( n81936 , n81931 , n81935 );
xor ( n81937 , n81871 , n81891 );
xor ( n81938 , n81937 , n81896 );
and ( n81939 , n81935 , n81938 );
and ( n81940 , n81931 , n81938 );
or ( n81941 , n81936 , n81939 , n81940 );
and ( n81942 , n80774 , n80705 );
and ( n81943 , n80694 , n80703 );
nor ( n81944 , n81942 , n81943 );
xnor ( n81945 , n81944 , n80577 );
and ( n81946 , n81941 , n81945 );
xor ( n81947 , n81766 , n81770 );
xor ( n81948 , n81947 , n81773 );
and ( n81949 , n81945 , n81948 );
and ( n81950 , n81941 , n81948 );
or ( n81951 , n81946 , n81949 , n81950 );
and ( n81952 , n80472 , n81011 );
and ( n81953 , n80383 , n81008 );
nor ( n81954 , n81952 , n81953 );
xnor ( n81955 , n81954 , n80681 );
and ( n81956 , n81951 , n81955 );
xor ( n81957 , n81860 , n81864 );
xor ( n81958 , n81957 , n81867 );
and ( n81959 , n81955 , n81958 );
and ( n81960 , n81951 , n81958 );
or ( n81961 , n81956 , n81959 , n81960 );
xor ( n81962 , n81838 , n81842 );
xor ( n81963 , n81962 , n81845 );
and ( n81964 , n81961 , n81963 );
xor ( n81965 , n81870 , n81921 );
xor ( n81966 , n81965 , n81924 );
and ( n81967 , n81963 , n81966 );
and ( n81968 , n81961 , n81966 );
or ( n81969 , n81964 , n81967 , n81968 );
and ( n81970 , n81927 , n81969 );
xor ( n81971 , n81848 , n81850 );
xor ( n81972 , n81971 , n81853 );
and ( n81973 , n81969 , n81972 );
and ( n81974 , n81927 , n81972 );
or ( n81975 , n81970 , n81973 , n81974 );
and ( n81976 , n81856 , n81975 );
xor ( n81977 , n81808 , n81810 );
xor ( n81978 , n81977 , n81813 );
and ( n81979 , n81975 , n81978 );
and ( n81980 , n81856 , n81978 );
or ( n81981 , n81976 , n81979 , n81980 );
and ( n81982 , n81834 , n81981 );
xor ( n81983 , n81834 , n81981 );
xor ( n81984 , n81856 , n81975 );
xor ( n81985 , n81984 , n81978 );
xor ( n81986 , n81927 , n81969 );
xor ( n81987 , n81986 , n81972 );
and ( n81988 , n80526 , n81011 );
and ( n81989 , n80472 , n81008 );
nor ( n81990 , n81988 , n81989 );
xnor ( n81991 , n81990 , n80681 );
and ( n81992 , n80618 , n80806 );
and ( n81993 , n80587 , n80804 );
nor ( n81994 , n81992 , n81993 );
xnor ( n81995 , n81994 , n80684 );
and ( n81996 , n81991 , n81995 );
xor ( n81997 , n81899 , n81903 );
xor ( n81998 , n81997 , n81908 );
and ( n81999 , n81995 , n81998 );
and ( n82000 , n81991 , n81998 );
or ( n82001 , n81996 , n81999 , n82000 );
and ( n82002 , n81641 , n80237 );
and ( n82003 , n81626 , n80235 );
nor ( n82004 , n82002 , n82003 );
xnor ( n82005 , n82004 , n80215 );
and ( n82006 , n81703 , n80170 );
and ( n82007 , n81708 , n80168 );
nor ( n82008 , n82006 , n82007 );
xnor ( n82009 , n82008 , n80175 );
xor ( n82010 , n82005 , n82009 );
and ( n82011 , n81497 , n80303 );
and ( n82012 , n81364 , n80301 );
nor ( n82013 , n82011 , n82012 );
xnor ( n82014 , n82013 , n80263 );
and ( n82015 , n82010 , n82014 );
xor ( n82016 , n79997 , n79998 );
xor ( n82017 , n82016 , n80000 );
buf ( n82018 , n82017 );
buf ( n82019 , n82018 );
buf ( n82020 , n82019 );
and ( n82021 , n82020 , n80155 );
and ( n82022 , n81884 , n80153 );
nor ( n82023 , n82021 , n82022 );
not ( n82024 , n82023 );
and ( n82025 , n82014 , n82024 );
and ( n82026 , n82010 , n82024 );
or ( n82027 , n82015 , n82025 , n82026 );
and ( n82028 , n81134 , n80503 );
and ( n82029 , n80999 , n80501 );
nor ( n82030 , n82028 , n82029 );
xnor ( n82031 , n82030 , n80462 );
and ( n82032 , n82027 , n82031 );
and ( n82033 , n81280 , n80376 );
and ( n82034 , n81129 , n80374 );
nor ( n82035 , n82033 , n82034 );
xnor ( n82036 , n82035 , n80338 );
and ( n82037 , n82031 , n82036 );
and ( n82038 , n82027 , n82036 );
or ( n82039 , n82032 , n82037 , n82038 );
and ( n82040 , n82005 , n82009 );
and ( n82041 , n81364 , n80303 );
and ( n82042 , n81275 , n80301 );
nor ( n82043 , n82041 , n82042 );
xnor ( n82044 , n82043 , n80263 );
and ( n82045 , n82040 , n82044 );
xor ( n82046 , n81875 , n81879 );
xor ( n82047 , n82046 , n81888 );
and ( n82048 , n82044 , n82047 );
and ( n82049 , n82040 , n82047 );
or ( n82050 , n82045 , n82048 , n82049 );
and ( n82051 , n82039 , n82050 );
and ( n82052 , n80999 , n80503 );
and ( n82053 , n80929 , n80501 );
nor ( n82054 , n82052 , n82053 );
xnor ( n82055 , n82054 , n80462 );
and ( n82056 , n82050 , n82055 );
and ( n82057 , n82039 , n82055 );
or ( n82058 , n82051 , n82056 , n82057 );
and ( n82059 , n80587 , n81011 );
and ( n82060 , n80526 , n81008 );
nor ( n82061 , n82059 , n82060 );
xnor ( n82062 , n82061 , n80681 );
and ( n82063 , n80826 , n80705 );
and ( n82064 , n80774 , n80703 );
nor ( n82065 , n82063 , n82064 );
xnor ( n82066 , n82065 , n80577 );
and ( n82067 , n82062 , n82066 );
xor ( n82068 , n81931 , n81935 );
xor ( n82069 , n82068 , n81938 );
and ( n82070 , n82066 , n82069 );
and ( n82071 , n82062 , n82069 );
or ( n82072 , n82067 , n82070 , n82071 );
and ( n82073 , n82058 , n82072 );
xor ( n82074 , n81941 , n81945 );
xor ( n82075 , n82074 , n81948 );
and ( n82076 , n82072 , n82075 );
and ( n82077 , n82058 , n82075 );
or ( n82078 , n82073 , n82076 , n82077 );
and ( n82079 , n82001 , n82078 );
xor ( n82080 , n81911 , n81915 );
xor ( n82081 , n82080 , n81918 );
and ( n82082 , n82078 , n82081 );
and ( n82083 , n82001 , n82081 );
or ( n82084 , n82079 , n82082 , n82083 );
and ( n82085 , n81708 , n80237 );
and ( n82086 , n81641 , n80235 );
nor ( n82087 , n82085 , n82086 );
xnor ( n82088 , n82087 , n80215 );
and ( n82089 , n81884 , n80170 );
and ( n82090 , n81703 , n80168 );
nor ( n82091 , n82089 , n82090 );
xnor ( n82092 , n82091 , n80175 );
and ( n82093 , n82088 , n82092 );
and ( n82094 , n82020 , n80153 );
and ( n82095 , n82092 , n82094 );
and ( n82096 , n82088 , n82094 );
or ( n82097 , n82093 , n82095 , n82096 );
and ( n82098 , n81129 , n80503 );
and ( n82099 , n81134 , n80501 );
nor ( n82100 , n82098 , n82099 );
xnor ( n82101 , n82100 , n80462 );
and ( n82102 , n82097 , n82101 );
and ( n82103 , n81275 , n80376 );
and ( n82104 , n81280 , n80374 );
nor ( n82105 , n82103 , n82104 );
xnor ( n82106 , n82105 , n80338 );
and ( n82107 , n82101 , n82106 );
and ( n82108 , n82097 , n82106 );
or ( n82109 , n82102 , n82107 , n82108 );
and ( n82110 , n80929 , n80705 );
and ( n82111 , n80826 , n80703 );
nor ( n82112 , n82110 , n82111 );
xnor ( n82113 , n82112 , n80577 );
and ( n82114 , n82109 , n82113 );
xor ( n82115 , n82040 , n82044 );
xor ( n82116 , n82115 , n82047 );
and ( n82117 , n82113 , n82116 );
and ( n82118 , n82109 , n82116 );
or ( n82119 , n82114 , n82117 , n82118 );
and ( n82120 , n80694 , n80806 );
and ( n82121 , n80618 , n80804 );
nor ( n82122 , n82120 , n82121 );
xnor ( n82123 , n82122 , n80684 );
and ( n82124 , n82119 , n82123 );
xor ( n82125 , n82039 , n82050 );
xor ( n82126 , n82125 , n82055 );
and ( n82127 , n82123 , n82126 );
and ( n82128 , n82119 , n82126 );
or ( n82129 , n82124 , n82127 , n82128 );
xor ( n82130 , n81991 , n81995 );
xor ( n82131 , n82130 , n81998 );
and ( n82132 , n82129 , n82131 );
xor ( n82133 , n82058 , n82072 );
xor ( n82134 , n82133 , n82075 );
and ( n82135 , n82131 , n82134 );
and ( n82136 , n82129 , n82134 );
or ( n82137 , n82132 , n82135 , n82136 );
xor ( n82138 , n81951 , n81955 );
xor ( n82139 , n82138 , n81958 );
and ( n82140 , n82137 , n82139 );
xor ( n82141 , n82001 , n82078 );
xor ( n82142 , n82141 , n82081 );
and ( n82143 , n82139 , n82142 );
and ( n82144 , n82137 , n82142 );
or ( n82145 , n82140 , n82143 , n82144 );
and ( n82146 , n82084 , n82145 );
xor ( n82147 , n81961 , n81963 );
xor ( n82148 , n82147 , n81966 );
and ( n82149 , n82145 , n82148 );
and ( n82150 , n82084 , n82148 );
or ( n82151 , n82146 , n82149 , n82150 );
and ( n82152 , n81987 , n82151 );
xor ( n82153 , n81987 , n82151 );
xor ( n82154 , n82084 , n82145 );
xor ( n82155 , n82154 , n82148 );
xor ( n82156 , n82137 , n82139 );
xor ( n82157 , n82156 , n82142 );
and ( n82158 , n80618 , n81011 );
and ( n82159 , n80587 , n81008 );
nor ( n82160 , n82158 , n82159 );
xnor ( n82161 , n82160 , n80681 );
and ( n82162 , n80774 , n80806 );
and ( n82163 , n80694 , n80804 );
nor ( n82164 , n82162 , n82163 );
xnor ( n82165 , n82164 , n80684 );
and ( n82166 , n82161 , n82165 );
xor ( n82167 , n82027 , n82031 );
xor ( n82168 , n82167 , n82036 );
and ( n82169 , n82165 , n82168 );
and ( n82170 , n82161 , n82168 );
or ( n82171 , n82166 , n82169 , n82170 );
and ( n82172 , n80826 , n80806 );
and ( n82173 , n80774 , n80804 );
nor ( n82174 , n82172 , n82173 );
xnor ( n82175 , n82174 , n80684 );
and ( n82176 , n80999 , n80705 );
and ( n82177 , n80929 , n80703 );
nor ( n82178 , n82176 , n82177 );
xnor ( n82179 , n82178 , n80577 );
and ( n82180 , n82175 , n82179 );
xor ( n82181 , n82097 , n82101 );
xor ( n82182 , n82181 , n82106 );
and ( n82183 , n82179 , n82182 );
and ( n82184 , n82175 , n82182 );
or ( n82185 , n82180 , n82183 , n82184 );
and ( n82186 , n81641 , n80303 );
and ( n82187 , n81626 , n80301 );
nor ( n82188 , n82186 , n82187 );
xnor ( n82189 , n82188 , n80263 );
buf ( n82190 , n78840 );
buf ( n82191 , n82190 );
buf ( n82192 , n82191 );
buf ( n82193 , n82192 );
and ( n82194 , n82193 , n80155 );
and ( n82195 , n82189 , n82194 );
and ( n82196 , n81364 , n80376 );
and ( n82197 , n81275 , n80374 );
nor ( n82198 , n82196 , n82197 );
xnor ( n82199 , n82198 , n80338 );
and ( n82200 , n82195 , n82199 );
and ( n82201 , n81626 , n80303 );
and ( n82202 , n81497 , n80301 );
nor ( n82203 , n82201 , n82202 );
xnor ( n82204 , n82203 , n80263 );
and ( n82205 , n82199 , n82204 );
and ( n82206 , n82195 , n82204 );
or ( n82207 , n82200 , n82205 , n82206 );
and ( n82208 , n81708 , n80303 );
and ( n82209 , n81641 , n80301 );
nor ( n82210 , n82208 , n82209 );
xnor ( n82211 , n82210 , n80263 );
and ( n82212 , n82193 , n80153 );
and ( n82213 , n82211 , n82212 );
and ( n82214 , n81703 , n80237 );
and ( n82215 , n81708 , n80235 );
nor ( n82216 , n82214 , n82215 );
xnor ( n82217 , n82216 , n80215 );
and ( n82218 , n82213 , n82217 );
and ( n82219 , n82020 , n80170 );
and ( n82220 , n81884 , n80168 );
nor ( n82221 , n82219 , n82220 );
xnor ( n82222 , n82221 , n80175 );
and ( n82223 , n82217 , n82222 );
and ( n82224 , n82213 , n82222 );
or ( n82225 , n82218 , n82223 , n82224 );
and ( n82226 , n81280 , n80503 );
and ( n82227 , n81129 , n80501 );
nor ( n82228 , n82226 , n82227 );
xnor ( n82229 , n82228 , n80462 );
and ( n82230 , n82225 , n82229 );
xor ( n82231 , n82088 , n82092 );
xor ( n82232 , n82231 , n82094 );
and ( n82233 , n82229 , n82232 );
and ( n82234 , n82225 , n82232 );
or ( n82235 , n82230 , n82233 , n82234 );
and ( n82236 , n82207 , n82235 );
xor ( n82237 , n82010 , n82014 );
xor ( n82238 , n82237 , n82024 );
and ( n82239 , n82235 , n82238 );
and ( n82240 , n82207 , n82238 );
or ( n82241 , n82236 , n82239 , n82240 );
and ( n82242 , n82185 , n82241 );
xor ( n82243 , n82109 , n82113 );
xor ( n82244 , n82243 , n82116 );
and ( n82245 , n82241 , n82244 );
and ( n82246 , n82185 , n82244 );
or ( n82247 , n82242 , n82245 , n82246 );
and ( n82248 , n82171 , n82247 );
xor ( n82249 , n82062 , n82066 );
xor ( n82250 , n82249 , n82069 );
and ( n82251 , n82247 , n82250 );
and ( n82252 , n82171 , n82250 );
or ( n82253 , n82248 , n82251 , n82252 );
xor ( n82254 , n82189 , n82194 );
and ( n82255 , n81626 , n80376 );
and ( n82256 , n81497 , n80374 );
nor ( n82257 , n82255 , n82256 );
xnor ( n82258 , n82257 , n80338 );
and ( n82259 , n81884 , n80237 );
and ( n82260 , n81703 , n80235 );
nor ( n82261 , n82259 , n82260 );
xnor ( n82262 , n82261 , n80215 );
and ( n82263 , n82258 , n82262 );
and ( n82264 , n82020 , n80168 );
not ( n82265 , n82264 );
xnor ( n82266 , n82265 , n80175 );
and ( n82267 , n82262 , n82266 );
and ( n82268 , n82258 , n82266 );
or ( n82269 , n82263 , n82267 , n82268 );
and ( n82270 , n82254 , n82269 );
and ( n82271 , n81497 , n80376 );
and ( n82272 , n81364 , n80374 );
nor ( n82273 , n82271 , n82272 );
xnor ( n82274 , n82273 , n80338 );
and ( n82275 , n82269 , n82274 );
and ( n82276 , n82254 , n82274 );
or ( n82277 , n82270 , n82275 , n82276 );
and ( n82278 , n81134 , n80705 );
and ( n82279 , n80999 , n80703 );
nor ( n82280 , n82278 , n82279 );
xnor ( n82281 , n82280 , n80577 );
and ( n82282 , n82277 , n82281 );
xor ( n82283 , n82195 , n82199 );
xor ( n82284 , n82283 , n82204 );
and ( n82285 , n82281 , n82284 );
and ( n82286 , n82277 , n82284 );
or ( n82287 , n82282 , n82285 , n82286 );
and ( n82288 , n80694 , n81011 );
and ( n82289 , n80618 , n81008 );
nor ( n82290 , n82288 , n82289 );
xnor ( n82291 , n82290 , n80681 );
and ( n82292 , n82287 , n82291 );
xor ( n82293 , n82207 , n82235 );
xor ( n82294 , n82293 , n82238 );
and ( n82295 , n82291 , n82294 );
and ( n82296 , n82287 , n82294 );
or ( n82297 , n82292 , n82295 , n82296 );
xor ( n82298 , n82161 , n82165 );
xor ( n82299 , n82298 , n82168 );
and ( n82300 , n82297 , n82299 );
xor ( n82301 , n82185 , n82241 );
xor ( n82302 , n82301 , n82244 );
and ( n82303 , n82299 , n82302 );
and ( n82304 , n82297 , n82302 );
or ( n82305 , n82300 , n82303 , n82304 );
xor ( n82306 , n82119 , n82123 );
xor ( n82307 , n82306 , n82126 );
and ( n82308 , n82305 , n82307 );
xor ( n82309 , n82171 , n82247 );
xor ( n82310 , n82309 , n82250 );
and ( n82311 , n82307 , n82310 );
and ( n82312 , n82305 , n82310 );
or ( n82313 , n82308 , n82311 , n82312 );
and ( n82314 , n82253 , n82313 );
xor ( n82315 , n82129 , n82131 );
xor ( n82316 , n82315 , n82134 );
and ( n82317 , n82313 , n82316 );
and ( n82318 , n82253 , n82316 );
or ( n82319 , n82314 , n82317 , n82318 );
and ( n82320 , n82157 , n82319 );
xor ( n82321 , n82157 , n82319 );
xor ( n82322 , n82253 , n82313 );
xor ( n82323 , n82322 , n82316 );
xor ( n82324 , n82305 , n82307 );
xor ( n82325 , n82324 , n82310 );
and ( n82326 , n81129 , n80705 );
and ( n82327 , n81134 , n80703 );
nor ( n82328 , n82326 , n82327 );
xnor ( n82329 , n82328 , n80577 );
and ( n82330 , n81275 , n80503 );
and ( n82331 , n81280 , n80501 );
nor ( n82332 , n82330 , n82331 );
xnor ( n82333 , n82332 , n80462 );
and ( n82334 , n82329 , n82333 );
xor ( n82335 , n82213 , n82217 );
xor ( n82336 , n82335 , n82222 );
and ( n82337 , n82333 , n82336 );
and ( n82338 , n82329 , n82336 );
or ( n82339 , n82334 , n82337 , n82338 );
and ( n82340 , n80929 , n80806 );
and ( n82341 , n80826 , n80804 );
nor ( n82342 , n82340 , n82341 );
xnor ( n82343 , n82342 , n80684 );
and ( n82344 , n82339 , n82343 );
xor ( n82345 , n82225 , n82229 );
xor ( n82346 , n82345 , n82232 );
and ( n82347 , n82343 , n82346 );
and ( n82348 , n82339 , n82346 );
or ( n82349 , n82344 , n82347 , n82348 );
xor ( n82350 , n82211 , n82212 );
and ( n82351 , n81641 , n80376 );
and ( n82352 , n81626 , n80374 );
nor ( n82353 , n82351 , n82352 );
xnor ( n82354 , n82353 , n80338 );
and ( n82355 , n81703 , n80303 );
and ( n82356 , n81708 , n80301 );
nor ( n82357 , n82355 , n82356 );
xnor ( n82358 , n82357 , n80263 );
and ( n82359 , n82354 , n82358 );
and ( n82360 , n82193 , n80168 );
not ( n82361 , n82360 );
and ( n82362 , n82361 , n80175 );
and ( n82363 , n82358 , n82362 );
and ( n82364 , n82354 , n82362 );
or ( n82365 , n82359 , n82363 , n82364 );
and ( n82366 , n82350 , n82365 );
and ( n82367 , n81364 , n80503 );
and ( n82368 , n81275 , n80501 );
nor ( n82369 , n82367 , n82368 );
xnor ( n82370 , n82369 , n80462 );
and ( n82371 , n82365 , n82370 );
and ( n82372 , n82350 , n82370 );
or ( n82373 , n82366 , n82371 , n82372 );
and ( n82374 , n80999 , n80806 );
and ( n82375 , n80929 , n80804 );
nor ( n82376 , n82374 , n82375 );
xnor ( n82377 , n82376 , n80684 );
and ( n82378 , n82373 , n82377 );
xor ( n82379 , n82254 , n82269 );
xor ( n82380 , n82379 , n82274 );
and ( n82381 , n82377 , n82380 );
and ( n82382 , n82373 , n82380 );
or ( n82383 , n82378 , n82381 , n82382 );
and ( n82384 , n80774 , n81011 );
and ( n82385 , n80694 , n81008 );
nor ( n82386 , n82384 , n82385 );
xnor ( n82387 , n82386 , n80681 );
and ( n82388 , n82383 , n82387 );
xor ( n82389 , n82277 , n82281 );
xor ( n82390 , n82389 , n82284 );
and ( n82391 , n82387 , n82390 );
and ( n82392 , n82383 , n82390 );
or ( n82393 , n82388 , n82391 , n82392 );
and ( n82394 , n82349 , n82393 );
xor ( n82395 , n82175 , n82179 );
xor ( n82396 , n82395 , n82182 );
and ( n82397 , n82393 , n82396 );
and ( n82398 , n82349 , n82396 );
or ( n82399 , n82394 , n82397 , n82398 );
and ( n82400 , n81708 , n80376 );
and ( n82401 , n81641 , n80374 );
nor ( n82402 , n82400 , n82401 );
xnor ( n82403 , n82402 , n80338 );
and ( n82404 , n82403 , n82360 );
and ( n82405 , n82020 , n80237 );
and ( n82406 , n81884 , n80235 );
nor ( n82407 , n82405 , n82406 );
xnor ( n82408 , n82407 , n80215 );
and ( n82409 , n82404 , n82408 );
and ( n82410 , n82193 , n80170 );
not ( n82411 , n82410 );
xnor ( n82412 , n82411 , n80175 );
and ( n82413 , n82408 , n82412 );
and ( n82414 , n82404 , n82412 );
or ( n82415 , n82409 , n82413 , n82414 );
and ( n82416 , n81280 , n80705 );
and ( n82417 , n81129 , n80703 );
nor ( n82418 , n82416 , n82417 );
xnor ( n82419 , n82418 , n80577 );
and ( n82420 , n82415 , n82419 );
xor ( n82421 , n82258 , n82262 );
xor ( n82422 , n82421 , n82266 );
and ( n82423 , n82419 , n82422 );
and ( n82424 , n82415 , n82422 );
or ( n82425 , n82420 , n82423 , n82424 );
and ( n82426 , n80826 , n81011 );
and ( n82427 , n80774 , n81008 );
nor ( n82428 , n82426 , n82427 );
xnor ( n82429 , n82428 , n80681 );
and ( n82430 , n82425 , n82429 );
xor ( n82431 , n82329 , n82333 );
xor ( n82432 , n82431 , n82336 );
and ( n82433 , n82429 , n82432 );
and ( n82434 , n82425 , n82432 );
or ( n82435 , n82430 , n82433 , n82434 );
xor ( n82436 , n82339 , n82343 );
xor ( n82437 , n82436 , n82346 );
and ( n82438 , n82435 , n82437 );
xor ( n82439 , n82383 , n82387 );
xor ( n82440 , n82439 , n82390 );
and ( n82441 , n82437 , n82440 );
and ( n82442 , n82435 , n82440 );
or ( n82443 , n82438 , n82441 , n82442 );
xor ( n82444 , n82287 , n82291 );
xor ( n82445 , n82444 , n82294 );
and ( n82446 , n82443 , n82445 );
xor ( n82447 , n82349 , n82393 );
xor ( n82448 , n82447 , n82396 );
and ( n82449 , n82445 , n82448 );
and ( n82450 , n82443 , n82448 );
or ( n82451 , n82446 , n82449 , n82450 );
and ( n82452 , n82399 , n82451 );
xor ( n82453 , n82297 , n82299 );
xor ( n82454 , n82453 , n82302 );
and ( n82455 , n82451 , n82454 );
and ( n82456 , n82399 , n82454 );
or ( n82457 , n82452 , n82455 , n82456 );
and ( n82458 , n82325 , n82457 );
xor ( n82459 , n82325 , n82457 );
xor ( n82460 , n82399 , n82451 );
xor ( n82461 , n82460 , n82454 );
xor ( n82462 , n82443 , n82445 );
xor ( n82463 , n82462 , n82448 );
and ( n82464 , n81626 , n80503 );
and ( n82465 , n81497 , n80501 );
nor ( n82466 , n82464 , n82465 );
xnor ( n82467 , n82466 , n80462 );
and ( n82468 , n81884 , n80303 );
and ( n82469 , n81703 , n80301 );
nor ( n82470 , n82468 , n82469 );
xnor ( n82471 , n82470 , n80263 );
and ( n82472 , n82467 , n82471 );
and ( n82473 , n82020 , n80235 );
not ( n82474 , n82473 );
xnor ( n82475 , n82474 , n80215 );
and ( n82476 , n82471 , n82475 );
and ( n82477 , n82467 , n82475 );
or ( n82478 , n82472 , n82476 , n82477 );
and ( n82479 , n81497 , n80503 );
and ( n82480 , n81364 , n80501 );
nor ( n82481 , n82479 , n82480 );
xnor ( n82482 , n82481 , n80462 );
and ( n82483 , n82478 , n82482 );
xor ( n82484 , n82354 , n82358 );
xor ( n82485 , n82484 , n82362 );
and ( n82486 , n82482 , n82485 );
and ( n82487 , n82478 , n82485 );
or ( n82488 , n82483 , n82486 , n82487 );
and ( n82489 , n81134 , n80806 );
and ( n82490 , n80999 , n80804 );
nor ( n82491 , n82489 , n82490 );
xnor ( n82492 , n82491 , n80684 );
and ( n82493 , n82488 , n82492 );
xor ( n82494 , n82350 , n82365 );
xor ( n82495 , n82494 , n82370 );
and ( n82496 , n82492 , n82495 );
and ( n82497 , n82488 , n82495 );
or ( n82498 , n82493 , n82496 , n82497 );
and ( n82499 , n81129 , n80806 );
and ( n82500 , n81134 , n80804 );
nor ( n82501 , n82499 , n82500 );
xnor ( n82502 , n82501 , n80684 );
and ( n82503 , n81275 , n80705 );
and ( n82504 , n81280 , n80703 );
nor ( n82505 , n82503 , n82504 );
xnor ( n82506 , n82505 , n80577 );
and ( n82507 , n82502 , n82506 );
xor ( n82508 , n82404 , n82408 );
xor ( n82509 , n82508 , n82412 );
and ( n82510 , n82506 , n82509 );
and ( n82511 , n82502 , n82509 );
or ( n82512 , n82507 , n82510 , n82511 );
and ( n82513 , n80929 , n81011 );
and ( n82514 , n80826 , n81008 );
nor ( n82515 , n82513 , n82514 );
xnor ( n82516 , n82515 , n80681 );
and ( n82517 , n82512 , n82516 );
xor ( n82518 , n82415 , n82419 );
xor ( n82519 , n82518 , n82422 );
and ( n82520 , n82516 , n82519 );
and ( n82521 , n82512 , n82519 );
or ( n82522 , n82517 , n82520 , n82521 );
and ( n82523 , n82498 , n82522 );
xor ( n82524 , n82373 , n82377 );
xor ( n82525 , n82524 , n82380 );
and ( n82526 , n82522 , n82525 );
and ( n82527 , n82498 , n82525 );
or ( n82528 , n82523 , n82526 , n82527 );
xor ( n82529 , n82403 , n82360 );
and ( n82530 , n81641 , n80503 );
and ( n82531 , n81626 , n80501 );
nor ( n82532 , n82530 , n82531 );
xnor ( n82533 , n82532 , n80462 );
and ( n82534 , n82020 , n80303 );
and ( n82535 , n81884 , n80301 );
nor ( n82536 , n82534 , n82535 );
xnor ( n82537 , n82536 , n80263 );
and ( n82538 , n82533 , n82537 );
and ( n82539 , n82193 , n80235 );
not ( n82540 , n82539 );
and ( n82541 , n82540 , n80215 );
and ( n82542 , n82537 , n82541 );
and ( n82543 , n82533 , n82541 );
or ( n82544 , n82538 , n82542 , n82543 );
and ( n82545 , n82529 , n82544 );
and ( n82546 , n81364 , n80705 );
and ( n82547 , n81275 , n80703 );
nor ( n82548 , n82546 , n82547 );
xnor ( n82549 , n82548 , n80577 );
and ( n82550 , n82544 , n82549 );
and ( n82551 , n82529 , n82549 );
or ( n82552 , n82545 , n82550 , n82551 );
and ( n82553 , n80999 , n81011 );
and ( n82554 , n80929 , n81008 );
nor ( n82555 , n82553 , n82554 );
xnor ( n82556 , n82555 , n80681 );
and ( n82557 , n82552 , n82556 );
xor ( n82558 , n82478 , n82482 );
xor ( n82559 , n82558 , n82485 );
and ( n82560 , n82556 , n82559 );
and ( n82561 , n82552 , n82559 );
or ( n82562 , n82557 , n82560 , n82561 );
xor ( n82563 , n82488 , n82492 );
xor ( n82564 , n82563 , n82495 );
and ( n82565 , n82562 , n82564 );
xor ( n82566 , n82512 , n82516 );
xor ( n82567 , n82566 , n82519 );
and ( n82568 , n82564 , n82567 );
and ( n82569 , n82562 , n82567 );
or ( n82570 , n82565 , n82568 , n82569 );
xor ( n82571 , n82425 , n82429 );
xor ( n82572 , n82571 , n82432 );
and ( n82573 , n82570 , n82572 );
xor ( n82574 , n82498 , n82522 );
xor ( n82575 , n82574 , n82525 );
and ( n82576 , n82572 , n82575 );
and ( n82577 , n82570 , n82575 );
or ( n82578 , n82573 , n82576 , n82577 );
and ( n82579 , n82528 , n82578 );
xor ( n82580 , n82435 , n82437 );
xor ( n82581 , n82580 , n82440 );
and ( n82582 , n82578 , n82581 );
and ( n82583 , n82528 , n82581 );
or ( n82584 , n82579 , n82582 , n82583 );
and ( n82585 , n82463 , n82584 );
xor ( n82586 , n82463 , n82584 );
xor ( n82587 , n82528 , n82578 );
xor ( n82588 , n82587 , n82581 );
xor ( n82589 , n82570 , n82572 );
xor ( n82590 , n82589 , n82575 );
and ( n82591 , n81708 , n80503 );
and ( n82592 , n81641 , n80501 );
nor ( n82593 , n82591 , n82592 );
xnor ( n82594 , n82593 , n80462 );
and ( n82595 , n82594 , n82539 );
and ( n82596 , n81703 , n80376 );
and ( n82597 , n81708 , n80374 );
nor ( n82598 , n82596 , n82597 );
xnor ( n82599 , n82598 , n80338 );
and ( n82600 , n82595 , n82599 );
and ( n82601 , n82193 , n80237 );
not ( n82602 , n82601 );
xnor ( n82603 , n82602 , n80215 );
and ( n82604 , n82599 , n82603 );
and ( n82605 , n82595 , n82603 );
or ( n82606 , n82600 , n82604 , n82605 );
and ( n82607 , n81280 , n80806 );
and ( n82608 , n81129 , n80804 );
nor ( n82609 , n82607 , n82608 );
xnor ( n82610 , n82609 , n80684 );
and ( n82611 , n82606 , n82610 );
xor ( n82612 , n82467 , n82471 );
xor ( n82613 , n82612 , n82475 );
and ( n82614 , n82610 , n82613 );
and ( n82615 , n82606 , n82613 );
or ( n82616 , n82611 , n82614 , n82615 );
and ( n82617 , n81626 , n80705 );
and ( n82618 , n81497 , n80703 );
nor ( n82619 , n82617 , n82618 );
xnor ( n82620 , n82619 , n80577 );
and ( n82621 , n81884 , n80376 );
and ( n82622 , n81703 , n80374 );
nor ( n82623 , n82621 , n82622 );
xnor ( n82624 , n82623 , n80338 );
and ( n82625 , n82620 , n82624 );
and ( n82626 , n82020 , n80301 );
not ( n82627 , n82626 );
xnor ( n82628 , n82627 , n80263 );
and ( n82629 , n82624 , n82628 );
and ( n82630 , n82620 , n82628 );
or ( n82631 , n82625 , n82629 , n82630 );
and ( n82632 , n81497 , n80705 );
and ( n82633 , n81364 , n80703 );
nor ( n82634 , n82632 , n82633 );
xnor ( n82635 , n82634 , n80577 );
and ( n82636 , n82631 , n82635 );
xor ( n82637 , n82533 , n82537 );
xor ( n82638 , n82637 , n82541 );
and ( n82639 , n82635 , n82638 );
and ( n82640 , n82631 , n82638 );
or ( n82641 , n82636 , n82639 , n82640 );
and ( n82642 , n81134 , n81011 );
and ( n82643 , n80999 , n81008 );
nor ( n82644 , n82642 , n82643 );
xnor ( n82645 , n82644 , n80681 );
and ( n82646 , n82641 , n82645 );
xor ( n82647 , n82529 , n82544 );
xor ( n82648 , n82647 , n82549 );
and ( n82649 , n82645 , n82648 );
and ( n82650 , n82641 , n82648 );
or ( n82651 , n82646 , n82649 , n82650 );
and ( n82652 , n82616 , n82651 );
xor ( n82653 , n82502 , n82506 );
xor ( n82654 , n82653 , n82509 );
and ( n82655 , n82651 , n82654 );
and ( n82656 , n82616 , n82654 );
or ( n82657 , n82652 , n82655 , n82656 );
and ( n82658 , n81129 , n81011 );
and ( n82659 , n81134 , n81008 );
nor ( n82660 , n82658 , n82659 );
xnor ( n82661 , n82660 , n80681 );
and ( n82662 , n81275 , n80806 );
and ( n82663 , n81280 , n80804 );
nor ( n82664 , n82662 , n82663 );
xnor ( n82665 , n82664 , n80684 );
and ( n82666 , n82661 , n82665 );
xor ( n82667 , n82595 , n82599 );
xor ( n82668 , n82667 , n82603 );
and ( n82669 , n82665 , n82668 );
and ( n82670 , n82661 , n82668 );
or ( n82671 , n82666 , n82669 , n82670 );
xor ( n82672 , n82606 , n82610 );
xor ( n82673 , n82672 , n82613 );
and ( n82674 , n82671 , n82673 );
xor ( n82675 , n82641 , n82645 );
xor ( n82676 , n82675 , n82648 );
and ( n82677 , n82673 , n82676 );
and ( n82678 , n82671 , n82676 );
or ( n82679 , n82674 , n82677 , n82678 );
xor ( n82680 , n82552 , n82556 );
xor ( n82681 , n82680 , n82559 );
and ( n82682 , n82679 , n82681 );
xor ( n82683 , n82616 , n82651 );
xor ( n82684 , n82683 , n82654 );
and ( n82685 , n82681 , n82684 );
and ( n82686 , n82679 , n82684 );
or ( n82687 , n82682 , n82685 , n82686 );
and ( n82688 , n82657 , n82687 );
xor ( n82689 , n82562 , n82564 );
xor ( n82690 , n82689 , n82567 );
and ( n82691 , n82687 , n82690 );
and ( n82692 , n82657 , n82690 );
or ( n82693 , n82688 , n82691 , n82692 );
and ( n82694 , n82590 , n82693 );
xor ( n82695 , n82590 , n82693 );
xor ( n82696 , n82657 , n82687 );
xor ( n82697 , n82696 , n82690 );
xor ( n82698 , n82679 , n82681 );
xor ( n82699 , n82698 , n82684 );
xor ( n82700 , n82594 , n82539 );
and ( n82701 , n81703 , n80503 );
and ( n82702 , n81708 , n80501 );
nor ( n82703 , n82701 , n82702 );
xnor ( n82704 , n82703 , n80462 );
and ( n82705 , n82020 , n80376 );
and ( n82706 , n81884 , n80374 );
nor ( n82707 , n82705 , n82706 );
xnor ( n82708 , n82707 , n80338 );
and ( n82709 , n82704 , n82708 );
and ( n82710 , n82193 , n80301 );
not ( n82711 , n82710 );
and ( n82712 , n82711 , n80263 );
and ( n82713 , n82708 , n82712 );
and ( n82714 , n82704 , n82712 );
or ( n82715 , n82709 , n82713 , n82714 );
and ( n82716 , n82700 , n82715 );
and ( n82717 , n81364 , n80806 );
and ( n82718 , n81275 , n80804 );
nor ( n82719 , n82717 , n82718 );
xnor ( n82720 , n82719 , n80684 );
and ( n82721 , n82715 , n82720 );
and ( n82722 , n82700 , n82720 );
or ( n82723 , n82716 , n82721 , n82722 );
and ( n82724 , n81884 , n80503 );
and ( n82725 , n81703 , n80501 );
nor ( n82726 , n82724 , n82725 );
xnor ( n82727 , n82726 , n80462 );
and ( n82728 , n82727 , n82710 );
and ( n82729 , n81641 , n80705 );
and ( n82730 , n81626 , n80703 );
nor ( n82731 , n82729 , n82730 );
xnor ( n82732 , n82731 , n80577 );
and ( n82733 , n82728 , n82732 );
and ( n82734 , n82193 , n80303 );
not ( n82735 , n82734 );
xnor ( n82736 , n82735 , n80263 );
and ( n82737 , n82732 , n82736 );
and ( n82738 , n82728 , n82736 );
or ( n82739 , n82733 , n82737 , n82738 );
and ( n82740 , n81280 , n81011 );
and ( n82741 , n81129 , n81008 );
nor ( n82742 , n82740 , n82741 );
xnor ( n82743 , n82742 , n80681 );
and ( n82744 , n82739 , n82743 );
xor ( n82745 , n82620 , n82624 );
xor ( n82746 , n82745 , n82628 );
and ( n82747 , n82743 , n82746 );
and ( n82748 , n82739 , n82746 );
or ( n82749 , n82744 , n82747 , n82748 );
and ( n82750 , n82723 , n82749 );
xor ( n82751 , n82631 , n82635 );
xor ( n82752 , n82751 , n82638 );
and ( n82753 , n82749 , n82752 );
and ( n82754 , n82723 , n82752 );
or ( n82755 , n82750 , n82753 , n82754 );
and ( n82756 , n81626 , n80806 );
and ( n82757 , n81497 , n80804 );
nor ( n82758 , n82756 , n82757 );
xnor ( n82759 , n82758 , n80684 );
and ( n82760 , n81708 , n80705 );
and ( n82761 , n81641 , n80703 );
nor ( n82762 , n82760 , n82761 );
xnor ( n82763 , n82762 , n80577 );
and ( n82764 , n82759 , n82763 );
and ( n82765 , n82020 , n80374 );
not ( n82766 , n82765 );
xnor ( n82767 , n82766 , n80338 );
and ( n82768 , n82763 , n82767 );
and ( n82769 , n82759 , n82767 );
or ( n82770 , n82764 , n82768 , n82769 );
and ( n82771 , n81497 , n80806 );
and ( n82772 , n81364 , n80804 );
nor ( n82773 , n82771 , n82772 );
xnor ( n82774 , n82773 , n80684 );
and ( n82775 , n82770 , n82774 );
xor ( n82776 , n82704 , n82708 );
xor ( n82777 , n82776 , n82712 );
and ( n82778 , n82774 , n82777 );
and ( n82779 , n82770 , n82777 );
or ( n82780 , n82775 , n82778 , n82779 );
xor ( n82781 , n82700 , n82715 );
xor ( n82782 , n82781 , n82720 );
and ( n82783 , n82780 , n82782 );
xor ( n82784 , n82739 , n82743 );
xor ( n82785 , n82784 , n82746 );
and ( n82786 , n82782 , n82785 );
and ( n82787 , n82780 , n82785 );
or ( n82788 , n82783 , n82786 , n82787 );
xor ( n82789 , n82661 , n82665 );
xor ( n82790 , n82789 , n82668 );
and ( n82791 , n82788 , n82790 );
xor ( n82792 , n82723 , n82749 );
xor ( n82793 , n82792 , n82752 );
and ( n82794 , n82790 , n82793 );
and ( n82795 , n82788 , n82793 );
or ( n82796 , n82791 , n82794 , n82795 );
and ( n82797 , n82755 , n82796 );
xor ( n82798 , n82671 , n82673 );
xor ( n82799 , n82798 , n82676 );
and ( n82800 , n82796 , n82799 );
and ( n82801 , n82755 , n82799 );
or ( n82802 , n82797 , n82800 , n82801 );
and ( n82803 , n82699 , n82802 );
xor ( n82804 , n82699 , n82802 );
xor ( n82805 , n82755 , n82796 );
xor ( n82806 , n82805 , n82799 );
xor ( n82807 , n82788 , n82790 );
xor ( n82808 , n82807 , n82793 );
xor ( n82809 , n82727 , n82710 );
and ( n82810 , n81703 , n80705 );
and ( n82811 , n81708 , n80703 );
nor ( n82812 , n82810 , n82811 );
xnor ( n82813 , n82812 , n80577 );
and ( n82814 , n82020 , n80503 );
and ( n82815 , n81884 , n80501 );
nor ( n82816 , n82814 , n82815 );
xnor ( n82817 , n82816 , n80462 );
and ( n82818 , n82813 , n82817 );
and ( n82819 , n82193 , n80374 );
not ( n82820 , n82819 );
and ( n82821 , n82820 , n80338 );
and ( n82822 , n82817 , n82821 );
and ( n82823 , n82813 , n82821 );
or ( n82824 , n82818 , n82822 , n82823 );
and ( n82825 , n82809 , n82824 );
and ( n82826 , n81708 , n80806 );
and ( n82827 , n81641 , n80804 );
nor ( n82828 , n82826 , n82827 );
xnor ( n82829 , n82828 , n80684 );
and ( n82830 , n82829 , n82819 );
and ( n82831 , n81641 , n80806 );
and ( n82832 , n81626 , n80804 );
nor ( n82833 , n82831 , n82832 );
xnor ( n82834 , n82833 , n80684 );
and ( n82835 , n82830 , n82834 );
and ( n82836 , n82193 , n80376 );
not ( n82837 , n82836 );
xnor ( n82838 , n82837 , n80338 );
and ( n82839 , n82834 , n82838 );
and ( n82840 , n82830 , n82838 );
or ( n82841 , n82835 , n82839 , n82840 );
and ( n82842 , n82824 , n82841 );
and ( n82843 , n82809 , n82841 );
or ( n82844 , n82825 , n82842 , n82843 );
and ( n82845 , n81275 , n81011 );
and ( n82846 , n81280 , n81008 );
nor ( n82847 , n82845 , n82846 );
xnor ( n82848 , n82847 , n80681 );
and ( n82849 , n82844 , n82848 );
xor ( n82850 , n82728 , n82732 );
xor ( n82851 , n82850 , n82736 );
and ( n82852 , n82848 , n82851 );
and ( n82853 , n82844 , n82851 );
or ( n82854 , n82849 , n82852 , n82853 );
xor ( n82855 , n82829 , n82819 );
and ( n82856 , n81884 , n80705 );
and ( n82857 , n81703 , n80703 );
nor ( n82858 , n82856 , n82857 );
xnor ( n82859 , n82858 , n80577 );
and ( n82860 , n82855 , n82859 );
and ( n82861 , n82020 , n80501 );
not ( n82862 , n82861 );
xnor ( n82863 , n82862 , n80462 );
and ( n82864 , n82859 , n82863 );
and ( n82865 , n82855 , n82863 );
or ( n82866 , n82860 , n82864 , n82865 );
and ( n82867 , n81497 , n81011 );
and ( n82868 , n81364 , n81008 );
nor ( n82869 , n82867 , n82868 );
xnor ( n82870 , n82869 , n80681 );
and ( n82871 , n82866 , n82870 );
xor ( n82872 , n82813 , n82817 );
xor ( n82873 , n82872 , n82821 );
and ( n82874 , n82870 , n82873 );
and ( n82875 , n82866 , n82873 );
or ( n82876 , n82871 , n82874 , n82875 );
and ( n82877 , n81364 , n81011 );
and ( n82878 , n81275 , n81008 );
nor ( n82879 , n82877 , n82878 );
xnor ( n82880 , n82879 , n80681 );
and ( n82881 , n82876 , n82880 );
xor ( n82882 , n82759 , n82763 );
xor ( n82883 , n82882 , n82767 );
and ( n82884 , n82880 , n82883 );
and ( n82885 , n82876 , n82883 );
or ( n82886 , n82881 , n82884 , n82885 );
xor ( n82887 , n82770 , n82774 );
xor ( n82888 , n82887 , n82777 );
and ( n82889 , n82886 , n82888 );
xor ( n82890 , n82844 , n82848 );
xor ( n82891 , n82890 , n82851 );
and ( n82892 , n82888 , n82891 );
and ( n82893 , n82886 , n82891 );
or ( n82894 , n82889 , n82892 , n82893 );
and ( n82895 , n82854 , n82894 );
xor ( n82896 , n82780 , n82782 );
xor ( n82897 , n82896 , n82785 );
and ( n82898 , n82894 , n82897 );
and ( n82899 , n82854 , n82897 );
or ( n82900 , n82895 , n82898 , n82899 );
and ( n82901 , n82808 , n82900 );
xor ( n82902 , n82808 , n82900 );
xor ( n82903 , n82854 , n82894 );
xor ( n82904 , n82903 , n82897 );
xor ( n82905 , n82886 , n82888 );
xor ( n82906 , n82905 , n82891 );
and ( n82907 , n81884 , n80806 );
and ( n82908 , n81703 , n80804 );
nor ( n82909 , n82907 , n82908 );
xnor ( n82910 , n82909 , n80684 );
and ( n82911 , n82193 , n80501 );
and ( n82912 , n82910 , n82911 );
and ( n82913 , n81703 , n80806 );
and ( n82914 , n81708 , n80804 );
nor ( n82915 , n82913 , n82914 );
xnor ( n82916 , n82915 , n80684 );
and ( n82917 , n82912 , n82916 );
not ( n82918 , n82911 );
and ( n82919 , n82918 , n80462 );
and ( n82920 , n82916 , n82919 );
and ( n82921 , n82912 , n82919 );
or ( n82922 , n82917 , n82920 , n82921 );
and ( n82923 , n81626 , n81011 );
and ( n82924 , n81497 , n81008 );
nor ( n82925 , n82923 , n82924 );
xnor ( n82926 , n82925 , n80681 );
and ( n82927 , n82922 , n82926 );
xor ( n82928 , n82855 , n82859 );
xor ( n82929 , n82928 , n82863 );
and ( n82930 , n82926 , n82929 );
and ( n82931 , n82922 , n82929 );
or ( n82932 , n82927 , n82930 , n82931 );
xor ( n82933 , n82830 , n82834 );
xor ( n82934 , n82933 , n82838 );
and ( n82935 , n82932 , n82934 );
xor ( n82936 , n82866 , n82870 );
xor ( n82937 , n82936 , n82873 );
and ( n82938 , n82934 , n82937 );
and ( n82939 , n82932 , n82937 );
or ( n82940 , n82935 , n82938 , n82939 );
xor ( n82941 , n82809 , n82824 );
xor ( n82942 , n82941 , n82841 );
and ( n82943 , n82940 , n82942 );
xor ( n82944 , n82876 , n82880 );
xor ( n82945 , n82944 , n82883 );
and ( n82946 , n82942 , n82945 );
and ( n82947 , n82940 , n82945 );
or ( n82948 , n82943 , n82946 , n82947 );
and ( n82949 , n82906 , n82948 );
xor ( n82950 , n82906 , n82948 );
xor ( n82951 , n82940 , n82942 );
xor ( n82952 , n82951 , n82945 );
xor ( n82953 , n82932 , n82934 );
xor ( n82954 , n82953 , n82937 );
and ( n82955 , n81641 , n81011 );
and ( n82956 , n81626 , n81008 );
nor ( n82957 , n82955 , n82956 );
xnor ( n82958 , n82957 , n80681 );
and ( n82959 , n82020 , n80705 );
and ( n82960 , n81884 , n80703 );
nor ( n82961 , n82959 , n82960 );
xnor ( n82962 , n82961 , n80577 );
and ( n82963 , n82958 , n82962 );
and ( n82964 , n82193 , n80503 );
not ( n82965 , n82964 );
xnor ( n82966 , n82965 , n80462 );
and ( n82967 , n82962 , n82966 );
and ( n82968 , n82958 , n82966 );
or ( n82969 , n82963 , n82967 , n82968 );
xor ( n82970 , n82910 , n82911 );
and ( n82971 , n81708 , n81011 );
and ( n82972 , n81641 , n81008 );
nor ( n82973 , n82971 , n82972 );
xnor ( n82974 , n82973 , n80681 );
and ( n82975 , n82970 , n82974 );
and ( n82976 , n82020 , n80703 );
not ( n82977 , n82976 );
xnor ( n82978 , n82977 , n80577 );
and ( n82979 , n82974 , n82978 );
and ( n82980 , n82970 , n82978 );
or ( n82981 , n82975 , n82979 , n82980 );
xor ( n82982 , n82958 , n82962 );
xor ( n82983 , n82982 , n82966 );
and ( n82984 , n82981 , n82983 );
xor ( n82985 , n82912 , n82916 );
xor ( n82986 , n82985 , n82919 );
and ( n82987 , n82983 , n82986 );
and ( n82988 , n82981 , n82986 );
or ( n82989 , n82984 , n82987 , n82988 );
and ( n82990 , n82969 , n82989 );
xor ( n82991 , n82922 , n82926 );
xor ( n82992 , n82991 , n82929 );
and ( n82993 , n82989 , n82992 );
and ( n82994 , n82969 , n82992 );
or ( n82995 , n82990 , n82993 , n82994 );
and ( n82996 , n82954 , n82995 );
xor ( n82997 , n82954 , n82995 );
xor ( n82998 , n82969 , n82989 );
xor ( n82999 , n82998 , n82992 );
xor ( n83000 , n82981 , n82983 );
xor ( n83001 , n83000 , n82986 );
and ( n83002 , n81703 , n81011 );
and ( n83003 , n81708 , n81008 );
nor ( n83004 , n83002 , n83003 );
xnor ( n83005 , n83004 , n80681 );
and ( n83006 , n82020 , n80806 );
and ( n83007 , n81884 , n80804 );
nor ( n83008 , n83006 , n83007 );
xnor ( n83009 , n83008 , n80684 );
and ( n83010 , n83005 , n83009 );
and ( n83011 , n82193 , n80703 );
not ( n83012 , n83011 );
and ( n83013 , n83012 , n80577 );
and ( n83014 , n83009 , n83013 );
and ( n83015 , n83005 , n83013 );
or ( n83016 , n83010 , n83014 , n83015 );
and ( n83017 , n82020 , n80804 );
not ( n83018 , n83017 );
xnor ( n83019 , n83018 , n80684 );
and ( n83020 , n83019 , n83011 );
and ( n83021 , n82193 , n80705 );
not ( n83022 , n83021 );
xnor ( n83023 , n83022 , n80577 );
and ( n83024 , n83020 , n83023 );
xor ( n83025 , n83005 , n83009 );
xor ( n83026 , n83025 , n83013 );
and ( n83027 , n83023 , n83026 );
and ( n83028 , n83020 , n83026 );
or ( n83029 , n83024 , n83027 , n83028 );
and ( n83030 , n83016 , n83029 );
xor ( n83031 , n82970 , n82974 );
xor ( n83032 , n83031 , n82978 );
and ( n83033 , n83029 , n83032 );
and ( n83034 , n83016 , n83032 );
or ( n83035 , n83030 , n83033 , n83034 );
and ( n83036 , n83001 , n83035 );
xor ( n83037 , n83001 , n83035 );
xor ( n83038 , n83016 , n83029 );
xor ( n83039 , n83038 , n83032 );
xor ( n83040 , n83020 , n83023 );
xor ( n83041 , n83040 , n83026 );
xor ( n83042 , n83019 , n83011 );
and ( n83043 , n82020 , n81011 );
and ( n83044 , n81884 , n81008 );
nor ( n83045 , n83043 , n83044 );
xnor ( n83046 , n83045 , n80681 );
and ( n83047 , n82193 , n80804 );
not ( n83048 , n83047 );
and ( n83049 , n83048 , n80684 );
and ( n83050 , n83046 , n83049 );
and ( n83051 , n82193 , n80806 );
not ( n83052 , n83051 );
xnor ( n83053 , n83052 , n80684 );
and ( n83054 , n83049 , n83053 );
and ( n83055 , n83046 , n83053 );
or ( n83056 , n83050 , n83054 , n83055 );
and ( n83057 , n83042 , n83056 );
and ( n83058 , n81884 , n81011 );
and ( n83059 , n81703 , n81008 );
nor ( n83060 , n83058 , n83059 );
xnor ( n83061 , n83060 , n80681 );
and ( n83062 , n83056 , n83061 );
and ( n83063 , n83042 , n83061 );
or ( n83064 , n83057 , n83062 , n83063 );
and ( n83065 , n83041 , n83064 );
xor ( n83066 , n83041 , n83064 );
xor ( n83067 , n83042 , n83056 );
xor ( n83068 , n83067 , n83061 );
xor ( n83069 , n83046 , n83049 );
xor ( n83070 , n83069 , n83053 );
and ( n83071 , n82020 , n81008 );
not ( n83072 , n83071 );
xnor ( n83073 , n83072 , n80681 );
and ( n83074 , n83073 , n83047 );
xor ( n83075 , n83073 , n83047 );
and ( n83076 , n82193 , n81011 );
not ( n83077 , n83076 );
xnor ( n83078 , n83077 , n80681 );
and ( n83079 , n82193 , n81008 );
not ( n83080 , n83079 );
and ( n83081 , n83080 , n80681 );
and ( n83082 , n83078 , n83081 );
and ( n83083 , n83075 , n83082 );
or ( n83084 , n83074 , n83083 );
and ( n83085 , n83070 , n83084 );
and ( n83086 , n83068 , n83085 );
and ( n83087 , n83066 , n83086 );
or ( n83088 , n83065 , n83087 );
and ( n83089 , n83039 , n83088 );
and ( n83090 , n83037 , n83089 );
or ( n83091 , n83036 , n83090 );
and ( n83092 , n82999 , n83091 );
and ( n83093 , n82997 , n83092 );
or ( n83094 , n82996 , n83093 );
and ( n83095 , n82952 , n83094 );
and ( n83096 , n82950 , n83095 );
or ( n83097 , n82949 , n83096 );
and ( n83098 , n82904 , n83097 );
and ( n83099 , n82902 , n83098 );
or ( n83100 , n82901 , n83099 );
and ( n83101 , n82806 , n83100 );
and ( n83102 , n82804 , n83101 );
or ( n83103 , n82803 , n83102 );
and ( n83104 , n82697 , n83103 );
and ( n83105 , n82695 , n83104 );
or ( n83106 , n82694 , n83105 );
and ( n83107 , n82588 , n83106 );
and ( n83108 , n82586 , n83107 );
or ( n83109 , n82585 , n83108 );
and ( n83110 , n82461 , n83109 );
and ( n83111 , n82459 , n83110 );
or ( n83112 , n82458 , n83111 );
and ( n83113 , n82323 , n83112 );
and ( n83114 , n82321 , n83113 );
or ( n83115 , n82320 , n83114 );
and ( n83116 , n82155 , n83115 );
and ( n83117 , n82153 , n83116 );
or ( n83118 , n82152 , n83117 );
and ( n83119 , n81985 , n83118 );
and ( n83120 , n81983 , n83119 );
or ( n83121 , n81982 , n83120 );
and ( n83122 , n81832 , n83121 );
and ( n83123 , n81830 , n83122 );
or ( n83124 , n81829 , n83123 );
and ( n83125 , n81611 , n83124 );
and ( n83126 , n81609 , n83125 );
or ( n83127 , n81608 , n83126 );
and ( n83128 , n81453 , n83127 );
and ( n83129 , n81451 , n83128 );
or ( n83130 , n81450 , n83129 );
and ( n83131 , n81265 , n83130 );
and ( n83132 , n81263 , n83131 );
or ( n83133 , n81262 , n83132 );
and ( n83134 , n81091 , n83133 );
and ( n83135 , n81089 , n83134 );
or ( n83136 , n81088 , n83135 );
and ( n83137 , n80914 , n83136 );
and ( n83138 , n80912 , n83137 );
or ( n83139 , n80911 , n83138 );
and ( n83140 , n80746 , n83139 );
and ( n83141 , n80744 , n83140 );
or ( n83142 , n80743 , n83141 );
and ( n83143 , n80561 , n83142 );
and ( n83144 , n80559 , n83143 );
or ( n83145 , n80558 , n83144 );
and ( n83146 , n80422 , n83145 );
and ( n83147 , n80420 , n83146 );
or ( n83148 , n80419 , n83147 );
and ( n83149 , n80297 , n83148 );
and ( n83150 , n80295 , n83149 );
or ( n83151 , n80294 , n83150 );
xor ( n83152 , n80199 , n83151 );
buf ( n83153 , n83152 );
buf ( n83154 , n83153 );
xor ( n83155 , n80295 , n83149 );
buf ( n83156 , n83155 );
buf ( n83157 , n83156 );
xor ( n83158 , n80297 , n83148 );
buf ( n83159 , n83158 );
buf ( n83160 , n83159 );
xor ( n83161 , n80420 , n83146 );
buf ( n83162 , n83161 );
buf ( n83163 , n83162 );
xor ( n83164 , n80422 , n83145 );
buf ( n83165 , n83164 );
buf ( n83166 , n83165 );
xor ( n83167 , n80559 , n83143 );
buf ( n83168 , n83167 );
buf ( n83169 , n83168 );
xor ( n83170 , n80561 , n83142 );
buf ( n83171 , n83170 );
buf ( n83172 , n83171 );
xor ( n83173 , n80744 , n83140 );
buf ( n83174 , n83173 );
buf ( n83175 , n83174 );
xor ( n83176 , n80746 , n83139 );
buf ( n83177 , n83176 );
buf ( n83178 , n83177 );
xor ( n83179 , n80912 , n83137 );
buf ( n83180 , n83179 );
buf ( n83181 , n83180 );
xor ( n83182 , n80914 , n83136 );
buf ( n83183 , n83182 );
buf ( n83184 , n83183 );
xor ( n83185 , n81089 , n83134 );
buf ( n83186 , n83185 );
buf ( n83187 , n83186 );
xor ( n83188 , n81091 , n83133 );
buf ( n83189 , n83188 );
buf ( n83190 , n83189 );
xor ( n83191 , n81263 , n83131 );
buf ( n83192 , n83191 );
buf ( n83193 , n83192 );
xor ( n83194 , n81265 , n83130 );
buf ( n83195 , n83194 );
buf ( n83196 , n83195 );
xor ( n83197 , n81451 , n83128 );
buf ( n83198 , n83197 );
buf ( n83199 , n83198 );
xor ( n83200 , n81453 , n83127 );
buf ( n83201 , n83200 );
buf ( n83202 , n83201 );
xor ( n83203 , n81609 , n83125 );
buf ( n83204 , n83203 );
buf ( n83205 , n83204 );
xor ( n83206 , n81611 , n83124 );
buf ( n83207 , n83206 );
buf ( n83208 , n83207 );
xor ( n83209 , n81830 , n83122 );
buf ( n83210 , n83209 );
buf ( n83211 , n83210 );
xor ( n83212 , n81832 , n83121 );
buf ( n83213 , n83212 );
buf ( n83214 , n83213 );
xor ( n83215 , n81983 , n83119 );
buf ( n83216 , n83215 );
buf ( n83217 , n83216 );
xor ( n83218 , n81985 , n83118 );
buf ( n83219 , n83218 );
buf ( n83220 , n83219 );
xor ( n83221 , n82153 , n83116 );
buf ( n83222 , n83221 );
buf ( n83223 , n83222 );
xor ( n83224 , n82155 , n83115 );
buf ( n83225 , n83224 );
buf ( n83226 , n83225 );
xor ( n83227 , n82321 , n83113 );
buf ( n83228 , n83227 );
buf ( n83229 , n83228 );
xor ( n83230 , n82323 , n83112 );
buf ( n83231 , n83230 );
buf ( n83232 , n83231 );
xor ( n83233 , n82459 , n83110 );
buf ( n83234 , n83233 );
buf ( n83235 , n83234 );
xor ( n83236 , n82461 , n83109 );
buf ( n83237 , n83236 );
buf ( n83238 , n83237 );
xor ( n83239 , n82586 , n83107 );
buf ( n83240 , n83239 );
buf ( n83241 , n83240 );
xor ( n83242 , n82588 , n83106 );
buf ( n83243 , n83242 );
buf ( n83244 , n83243 );
xor ( n83245 , n82695 , n83104 );
buf ( n83246 , n83245 );
buf ( n83247 , n83246 );
xor ( n83248 , n82697 , n83103 );
buf ( n83249 , n83248 );
buf ( n83250 , n83249 );
xor ( n83251 , n82804 , n83101 );
buf ( n83252 , n83251 );
buf ( n83253 , n83252 );
xor ( n83254 , n82806 , n83100 );
buf ( n83255 , n83254 );
buf ( n83256 , n83255 );
xor ( n83257 , n82902 , n83098 );
buf ( n83258 , n83257 );
buf ( n83259 , n83258 );
xor ( n83260 , n82904 , n83097 );
buf ( n83261 , n83260 );
buf ( n83262 , n83261 );
xor ( n83263 , n82950 , n83095 );
buf ( n83264 , n83263 );
buf ( n83265 , n83264 );
xor ( n83266 , n82952 , n83094 );
buf ( n83267 , n83266 );
buf ( n83268 , n83267 );
xor ( n83269 , n82997 , n83092 );
buf ( n83270 , n83269 );
buf ( n83271 , n83270 );
xor ( n83272 , n82999 , n83091 );
buf ( n83273 , n83272 );
buf ( n83274 , n83273 );
xor ( n83275 , n83037 , n83089 );
buf ( n83276 , n83275 );
buf ( n83277 , n83276 );
xor ( n83278 , n83039 , n83088 );
buf ( n83279 , n83278 );
buf ( n83280 , n83279 );
xor ( n83281 , n83066 , n83086 );
buf ( n83282 , n83281 );
buf ( n83283 , n83282 );
xor ( n83284 , n83068 , n83085 );
buf ( n83285 , n83284 );
buf ( n83286 , n83285 );
xor ( n83287 , n83070 , n83084 );
buf ( n83288 , n83287 );
buf ( n83289 , n83288 );
xor ( n83290 , n83075 , n83082 );
buf ( n83291 , n83290 );
buf ( n83292 , n83291 );
xor ( n83293 , n83078 , n83081 );
buf ( n83294 , n83293 );
buf ( n83295 , n83294 );
buf ( n83296 , n83079 );
buf ( n83297 , n83296 );
buf ( n83298 , n83297 );
and ( n83299 , n77811 , n83154 );
and ( n83300 , n77816 , n83157 );
and ( n83301 , n77821 , n83160 );
and ( n83302 , n77826 , n83163 );
and ( n83303 , n77831 , n83166 );
and ( n83304 , n77836 , n83169 );
and ( n83305 , n77841 , n83172 );
and ( n83306 , n77846 , n83175 );
and ( n83307 , n77851 , n83178 );
and ( n83308 , n77856 , n83181 );
and ( n83309 , n77861 , n83184 );
and ( n83310 , n77866 , n83187 );
and ( n83311 , n77871 , n83190 );
and ( n83312 , n77876 , n83193 );
and ( n83313 , n77881 , n83196 );
and ( n83314 , n77886 , n83199 );
and ( n83315 , n77891 , n83202 );
and ( n83316 , n77896 , n83205 );
and ( n83317 , n77901 , n83208 );
and ( n83318 , n77906 , n83211 );
and ( n83319 , n77911 , n83214 );
and ( n83320 , n77916 , n83217 );
and ( n83321 , n77921 , n83220 );
and ( n83322 , n77926 , n83223 );
and ( n83323 , n77931 , n83226 );
and ( n83324 , n77936 , n83229 );
and ( n83325 , n77941 , n83232 );
and ( n83326 , n77946 , n83235 );
and ( n83327 , n77951 , n83238 );
and ( n83328 , n77956 , n83241 );
and ( n83329 , n77961 , n83244 );
and ( n83330 , n77966 , n83247 );
and ( n83331 , n77971 , n83250 );
and ( n83332 , n77976 , n83253 );
and ( n83333 , n77981 , n83256 );
and ( n83334 , n77986 , n83259 );
and ( n83335 , n77991 , n83262 );
and ( n83336 , n77996 , n83265 );
and ( n83337 , n78001 , n83268 );
and ( n83338 , n78006 , n83271 );
and ( n83339 , n78011 , n83274 );
and ( n83340 , n78016 , n83277 );
and ( n83341 , n78021 , n83280 );
and ( n83342 , n78026 , n83283 );
and ( n83343 , n78031 , n83286 );
and ( n83344 , n78036 , n83289 );
and ( n83345 , n78041 , n83292 );
and ( n83346 , n78045 , n83295 );
buf ( n83347 , n83346 );
and ( n83348 , n83292 , n83347 );
and ( n83349 , n78041 , n83347 );
or ( n83350 , n83345 , n83348 , n83349 );
and ( n83351 , n83289 , n83350 );
and ( n83352 , n78036 , n83350 );
or ( n83353 , n83344 , n83351 , n83352 );
and ( n83354 , n83286 , n83353 );
and ( n83355 , n78031 , n83353 );
or ( n83356 , n83343 , n83354 , n83355 );
and ( n83357 , n83283 , n83356 );
and ( n83358 , n78026 , n83356 );
or ( n83359 , n83342 , n83357 , n83358 );
and ( n83360 , n83280 , n83359 );
and ( n83361 , n78021 , n83359 );
or ( n83362 , n83341 , n83360 , n83361 );
and ( n83363 , n83277 , n83362 );
and ( n83364 , n78016 , n83362 );
or ( n83365 , n83340 , n83363 , n83364 );
and ( n83366 , n83274 , n83365 );
and ( n83367 , n78011 , n83365 );
or ( n83368 , n83339 , n83366 , n83367 );
and ( n83369 , n83271 , n83368 );
and ( n83370 , n78006 , n83368 );
or ( n83371 , n83338 , n83369 , n83370 );
and ( n83372 , n83268 , n83371 );
and ( n83373 , n78001 , n83371 );
or ( n83374 , n83337 , n83372 , n83373 );
and ( n83375 , n83265 , n83374 );
and ( n83376 , n77996 , n83374 );
or ( n83377 , n83336 , n83375 , n83376 );
and ( n83378 , n83262 , n83377 );
and ( n83379 , n77991 , n83377 );
or ( n83380 , n83335 , n83378 , n83379 );
and ( n83381 , n83259 , n83380 );
and ( n83382 , n77986 , n83380 );
or ( n83383 , n83334 , n83381 , n83382 );
and ( n83384 , n83256 , n83383 );
and ( n83385 , n77981 , n83383 );
or ( n83386 , n83333 , n83384 , n83385 );
and ( n83387 , n83253 , n83386 );
and ( n83388 , n77976 , n83386 );
or ( n83389 , n83332 , n83387 , n83388 );
and ( n83390 , n83250 , n83389 );
and ( n83391 , n77971 , n83389 );
or ( n83392 , n83331 , n83390 , n83391 );
and ( n83393 , n83247 , n83392 );
and ( n83394 , n77966 , n83392 );
or ( n83395 , n83330 , n83393 , n83394 );
and ( n83396 , n83244 , n83395 );
and ( n83397 , n77961 , n83395 );
or ( n83398 , n83329 , n83396 , n83397 );
and ( n83399 , n83241 , n83398 );
and ( n83400 , n77956 , n83398 );
or ( n83401 , n83328 , n83399 , n83400 );
and ( n83402 , n83238 , n83401 );
and ( n83403 , n77951 , n83401 );
or ( n83404 , n83327 , n83402 , n83403 );
and ( n83405 , n83235 , n83404 );
and ( n83406 , n77946 , n83404 );
or ( n83407 , n83326 , n83405 , n83406 );
and ( n83408 , n83232 , n83407 );
and ( n83409 , n77941 , n83407 );
or ( n83410 , n83325 , n83408 , n83409 );
and ( n83411 , n83229 , n83410 );
and ( n83412 , n77936 , n83410 );
or ( n83413 , n83324 , n83411 , n83412 );
and ( n83414 , n83226 , n83413 );
and ( n83415 , n77931 , n83413 );
or ( n83416 , n83323 , n83414 , n83415 );
and ( n83417 , n83223 , n83416 );
and ( n83418 , n77926 , n83416 );
or ( n83419 , n83322 , n83417 , n83418 );
and ( n83420 , n83220 , n83419 );
and ( n83421 , n77921 , n83419 );
or ( n83422 , n83321 , n83420 , n83421 );
and ( n83423 , n83217 , n83422 );
and ( n83424 , n77916 , n83422 );
or ( n83425 , n83320 , n83423 , n83424 );
and ( n83426 , n83214 , n83425 );
and ( n83427 , n77911 , n83425 );
or ( n83428 , n83319 , n83426 , n83427 );
and ( n83429 , n83211 , n83428 );
and ( n83430 , n77906 , n83428 );
or ( n83431 , n83318 , n83429 , n83430 );
and ( n83432 , n83208 , n83431 );
and ( n83433 , n77901 , n83431 );
or ( n83434 , n83317 , n83432 , n83433 );
and ( n83435 , n83205 , n83434 );
and ( n83436 , n77896 , n83434 );
or ( n83437 , n83316 , n83435 , n83436 );
and ( n83438 , n83202 , n83437 );
and ( n83439 , n77891 , n83437 );
or ( n83440 , n83315 , n83438 , n83439 );
and ( n83441 , n83199 , n83440 );
and ( n83442 , n77886 , n83440 );
or ( n83443 , n83314 , n83441 , n83442 );
and ( n83444 , n83196 , n83443 );
and ( n83445 , n77881 , n83443 );
or ( n83446 , n83313 , n83444 , n83445 );
and ( n83447 , n83193 , n83446 );
and ( n83448 , n77876 , n83446 );
or ( n83449 , n83312 , n83447 , n83448 );
and ( n83450 , n83190 , n83449 );
and ( n83451 , n77871 , n83449 );
or ( n83452 , n83311 , n83450 , n83451 );
and ( n83453 , n83187 , n83452 );
and ( n83454 , n77866 , n83452 );
or ( n83455 , n83310 , n83453 , n83454 );
and ( n83456 , n83184 , n83455 );
and ( n83457 , n77861 , n83455 );
or ( n83458 , n83309 , n83456 , n83457 );
and ( n83459 , n83181 , n83458 );
and ( n83460 , n77856 , n83458 );
or ( n83461 , n83308 , n83459 , n83460 );
and ( n83462 , n83178 , n83461 );
and ( n83463 , n77851 , n83461 );
or ( n83464 , n83307 , n83462 , n83463 );
and ( n83465 , n83175 , n83464 );
and ( n83466 , n77846 , n83464 );
or ( n83467 , n83306 , n83465 , n83466 );
and ( n83468 , n83172 , n83467 );
and ( n83469 , n77841 , n83467 );
or ( n83470 , n83305 , n83468 , n83469 );
and ( n83471 , n83169 , n83470 );
and ( n83472 , n77836 , n83470 );
or ( n83473 , n83304 , n83471 , n83472 );
and ( n83474 , n83166 , n83473 );
and ( n83475 , n77831 , n83473 );
or ( n83476 , n83303 , n83474 , n83475 );
and ( n83477 , n83163 , n83476 );
and ( n83478 , n77826 , n83476 );
or ( n83479 , n83302 , n83477 , n83478 );
and ( n83480 , n83160 , n83479 );
and ( n83481 , n77821 , n83479 );
or ( n83482 , n83301 , n83480 , n83481 );
and ( n83483 , n83157 , n83482 );
and ( n83484 , n77816 , n83482 );
or ( n83485 , n83300 , n83483 , n83484 );
and ( n83486 , n83154 , n83485 );
and ( n83487 , n77811 , n83485 );
or ( n83488 , n83299 , n83486 , n83487 );
and ( n83489 , n77806 , n83488 );
and ( n83490 , n77801 , n83489 );
and ( n83491 , n77796 , n83490 );
and ( n83492 , n77791 , n83491 );
and ( n83493 , n77786 , n83492 );
and ( n83494 , n77781 , n83493 );
and ( n83495 , n77776 , n83494 );
and ( n83496 , n77771 , n83495 );
and ( n83497 , n77766 , n83496 );
and ( n83498 , n77761 , n83497 );
and ( n83499 , n77756 , n83498 );
and ( n83500 , n77751 , n83499 );
and ( n83501 , n77746 , n83500 );
and ( n83502 , n77741 , n83501 );
and ( n83503 , n77736 , n83502 );
and ( n83504 , n77731 , n83503 );
and ( n83505 , n77726 , n83504 );
and ( n83506 , n77721 , n83505 );
and ( n83507 , n77716 , n83506 );
and ( n83508 , n77711 , n83507 );
and ( n83509 , n77706 , n83508 );
and ( n83510 , n77701 , n83509 );
and ( n83511 , n77696 , n83510 );
and ( n83512 , n77691 , n83511 );
and ( n83513 , n77686 , n83512 );
and ( n83514 , n77681 , n83513 );
and ( n83515 , n77676 , n83514 );
and ( n83516 , n77671 , n83515 );
and ( n83517 , n77666 , n83516 );
and ( n83518 , n77661 , n83517 );
and ( n83519 , n77656 , n83518 );
and ( n83520 , n77651 , n83519 );
and ( n83521 , n77646 , n83520 );
and ( n83522 , n77641 , n83521 );
and ( n83523 , n77636 , n83522 );
and ( n83524 , n77631 , n83523 );
and ( n83525 , n77626 , n83524 );
and ( n83526 , n77621 , n83525 );
and ( n83527 , n77616 , n83526 );
and ( n83528 , n77611 , n83527 );
and ( n83529 , n77606 , n83528 );
and ( n83530 , n77601 , n83529 );
and ( n83531 , n77596 , n83530 );
and ( n83532 , n77591 , n83531 );
and ( n83533 , n77586 , n83532 );
and ( n83534 , n77581 , n83533 );
and ( n83535 , n77576 , n83534 );
and ( n83536 , n77571 , n83535 );
and ( n83537 , n77566 , n83536 );
and ( n83538 , n77561 , n83537 );
and ( n83539 , n77556 , n83538 );
and ( n83540 , n77551 , n83539 );
and ( n83541 , n77546 , n83540 );
and ( n83542 , n77541 , n83541 );
and ( n83543 , n77536 , n83542 );
and ( n83544 , n77531 , n83543 );
and ( n83545 , n77526 , n83544 );
and ( n83546 , n77521 , n83545 );
and ( n83547 , n77516 , n83546 );
and ( n83548 , n77511 , n83547 );
and ( n83549 , n77506 , n83548 );
and ( n83550 , n77501 , n83549 );
and ( n83551 , n77496 , n83550 );
and ( n83552 , n77491 , n83551 );
and ( n83553 , n77486 , n83552 );
and ( n83554 , n77481 , n83553 );
and ( n83555 , n77476 , n83554 );
and ( n83556 , n77471 , n83555 );
and ( n83557 , n77466 , n83556 );
and ( n83558 , n77461 , n83557 );
and ( n83559 , n77456 , n83558 );
and ( n83560 , n77451 , n83559 );
and ( n83561 , n77446 , n83560 );
and ( n83562 , n77441 , n83561 );
and ( n83563 , n77436 , n83562 );
and ( n83564 , n77431 , n83563 );
and ( n83565 , n77426 , n83564 );
and ( n83566 , n77421 , n83565 );
xor ( n83567 , n77416 , n83566 );
buf ( n83568 , n83567 );
xor ( n83569 , n77421 , n83565 );
buf ( n83570 , n83569 );
xor ( n83571 , n77426 , n83564 );
buf ( n83572 , n83571 );
xor ( n83573 , n77431 , n83563 );
buf ( n83574 , n83573 );
xor ( n83575 , n77436 , n83562 );
buf ( n83576 , n83575 );
xor ( n83577 , n77441 , n83561 );
buf ( n83578 , n83577 );
xor ( n83579 , n77446 , n83560 );
buf ( n83580 , n83579 );
xor ( n83581 , n77451 , n83559 );
buf ( n83582 , n83581 );
xor ( n83583 , n77456 , n83558 );
buf ( n83584 , n83583 );
xor ( n83585 , n77461 , n83557 );
buf ( n83586 , n83585 );
xor ( n83587 , n77466 , n83556 );
buf ( n83588 , n83587 );
xor ( n83589 , n77471 , n83555 );
buf ( n83590 , n83589 );
xor ( n83591 , n77476 , n83554 );
buf ( n83592 , n83591 );
xor ( n83593 , n77481 , n83553 );
buf ( n83594 , n83593 );
xor ( n83595 , n77486 , n83552 );
buf ( n83596 , n83595 );
xor ( n83597 , n77491 , n83551 );
buf ( n83598 , n83597 );
xor ( n83599 , n77496 , n83550 );
buf ( n83600 , n83599 );
xor ( n83601 , n77501 , n83549 );
buf ( n83602 , n83601 );
xor ( n83603 , n77506 , n83548 );
buf ( n83604 , n83603 );
xor ( n83605 , n77511 , n83547 );
buf ( n83606 , n83605 );
xor ( n83607 , n77516 , n83546 );
buf ( n83608 , n83607 );
xor ( n83609 , n77521 , n83545 );
buf ( n83610 , n83609 );
xor ( n83611 , n77526 , n83544 );
buf ( n83612 , n83611 );
xor ( n83613 , n77531 , n83543 );
buf ( n83614 , n83613 );
xor ( n83615 , n77536 , n83542 );
buf ( n83616 , n83615 );
xor ( n83617 , n77541 , n83541 );
buf ( n83618 , n83617 );
xor ( n83619 , n77546 , n83540 );
buf ( n83620 , n83619 );
xor ( n83621 , n77551 , n83539 );
buf ( n83622 , n83621 );
xor ( n83623 , n77556 , n83538 );
buf ( n83624 , n83623 );
xor ( n83625 , n77561 , n83537 );
buf ( n83626 , n83625 );
xor ( n83627 , n77566 , n83536 );
buf ( n83628 , n83627 );
xor ( n83629 , n77571 , n83535 );
buf ( n83630 , n83629 );
xor ( n83631 , n77576 , n83534 );
buf ( n83632 , n83631 );
xor ( n83633 , n77581 , n83533 );
buf ( n83634 , n83633 );
xor ( n83635 , n77586 , n83532 );
buf ( n83636 , n83635 );
xor ( n83637 , n77591 , n83531 );
buf ( n83638 , n83637 );
xor ( n83639 , n77596 , n83530 );
buf ( n83640 , n83639 );
xor ( n83641 , n77601 , n83529 );
buf ( n83642 , n83641 );
xor ( n83643 , n77606 , n83528 );
buf ( n83644 , n83643 );
xor ( n83645 , n77611 , n83527 );
buf ( n83646 , n83645 );
xor ( n83647 , n77616 , n83526 );
buf ( n83648 , n83647 );
xor ( n83649 , n77621 , n83525 );
buf ( n83650 , n83649 );
xor ( n83651 , n77626 , n83524 );
buf ( n83652 , n83651 );
xor ( n83653 , n77631 , n83523 );
buf ( n83654 , n83653 );
xor ( n83655 , n77636 , n83522 );
buf ( n83656 , n83655 );
xor ( n83657 , n77641 , n83521 );
buf ( n83658 , n83657 );
xor ( n83659 , n77646 , n83520 );
buf ( n83660 , n83659 );
xor ( n83661 , n77651 , n83519 );
buf ( n83662 , n83661 );
xor ( n83663 , n77656 , n83518 );
buf ( n83664 , n83663 );
xor ( n83665 , n77661 , n83517 );
buf ( n83666 , n83665 );
xor ( n83667 , n77666 , n83516 );
buf ( n83668 , n83667 );
xor ( n83669 , n77671 , n83515 );
buf ( n83670 , n83669 );
xor ( n83671 , n77676 , n83514 );
buf ( n83672 , n83671 );
xor ( n83673 , n77681 , n83513 );
buf ( n83674 , n83673 );
xor ( n83675 , n77686 , n83512 );
buf ( n83676 , n83675 );
xor ( n83677 , n77691 , n83511 );
buf ( n83678 , n83677 );
xor ( n83679 , n77696 , n83510 );
buf ( n83680 , n83679 );
xor ( n83681 , n77701 , n83509 );
buf ( n83682 , n83681 );
xor ( n83683 , n77706 , n83508 );
buf ( n83684 , n83683 );
xor ( n83685 , n77711 , n83507 );
buf ( n83686 , n83685 );
xor ( n83687 , n77716 , n83506 );
buf ( n83688 , n83687 );
xor ( n83689 , n77721 , n83505 );
buf ( n83690 , n83689 );
xor ( n83691 , n77726 , n83504 );
buf ( n83692 , n83691 );
xor ( n83693 , n77731 , n83503 );
buf ( n83694 , n83693 );
xor ( n83695 , n77736 , n83502 );
buf ( n83696 , n83695 );
xor ( n83697 , n77741 , n83501 );
buf ( n83698 , n83697 );
xor ( n83699 , n77746 , n83500 );
buf ( n83700 , n83699 );
xor ( n83701 , n77751 , n83499 );
buf ( n83702 , n83701 );
xor ( n83703 , n77756 , n83498 );
buf ( n83704 , n83703 );
xor ( n83705 , n77761 , n83497 );
buf ( n83706 , n83705 );
xor ( n83707 , n77766 , n83496 );
buf ( n83708 , n83707 );
xor ( n83709 , n77771 , n83495 );
buf ( n83710 , n83709 );
xor ( n83711 , n77776 , n83494 );
buf ( n83712 , n83711 );
xor ( n83713 , n77781 , n83493 );
buf ( n83714 , n83713 );
xor ( n83715 , n77786 , n83492 );
buf ( n83716 , n83715 );
xor ( n83717 , n77791 , n83491 );
buf ( n83718 , n83717 );
xor ( n83719 , n77796 , n83490 );
buf ( n83720 , n83719 );
xor ( n83721 , n77801 , n83489 );
buf ( n83722 , n83721 );
xor ( n83723 , n77806 , n83488 );
buf ( n83724 , n83723 );
xor ( n83725 , n77811 , n83154 );
xor ( n83726 , n83725 , n83485 );
buf ( n83727 , n83726 );
xor ( n83728 , n77816 , n83157 );
xor ( n83729 , n83728 , n83482 );
buf ( n83730 , n83729 );
xor ( n83731 , n77821 , n83160 );
xor ( n83732 , n83731 , n83479 );
buf ( n83733 , n83732 );
xor ( n83734 , n77826 , n83163 );
xor ( n83735 , n83734 , n83476 );
buf ( n83736 , n83735 );
xor ( n83737 , n77831 , n83166 );
xor ( n83738 , n83737 , n83473 );
buf ( n83739 , n83738 );
xor ( n83740 , n77836 , n83169 );
xor ( n83741 , n83740 , n83470 );
buf ( n83742 , n83741 );
xor ( n83743 , n77841 , n83172 );
xor ( n83744 , n83743 , n83467 );
buf ( n83745 , n83744 );
xor ( n83746 , n77846 , n83175 );
xor ( n83747 , n83746 , n83464 );
buf ( n83748 , n83747 );
xor ( n83749 , n77851 , n83178 );
xor ( n83750 , n83749 , n83461 );
buf ( n83751 , n83750 );
xor ( n83752 , n77856 , n83181 );
xor ( n83753 , n83752 , n83458 );
buf ( n83754 , n83753 );
xor ( n83755 , n77861 , n83184 );
xor ( n83756 , n83755 , n83455 );
buf ( n83757 , n83756 );
xor ( n83758 , n77866 , n83187 );
xor ( n83759 , n83758 , n83452 );
buf ( n83760 , n83759 );
xor ( n83761 , n77871 , n83190 );
xor ( n83762 , n83761 , n83449 );
buf ( n83763 , n83762 );
xor ( n83764 , n77876 , n83193 );
xor ( n83765 , n83764 , n83446 );
buf ( n83766 , n83765 );
xor ( n83767 , n77881 , n83196 );
xor ( n83768 , n83767 , n83443 );
buf ( n83769 , n83768 );
xor ( n83770 , n77886 , n83199 );
xor ( n83771 , n83770 , n83440 );
buf ( n83772 , n83771 );
xor ( n83773 , n77891 , n83202 );
xor ( n83774 , n83773 , n83437 );
buf ( n83775 , n83774 );
xor ( n83776 , n77896 , n83205 );
xor ( n83777 , n83776 , n83434 );
buf ( n83778 , n83777 );
xor ( n83779 , n77901 , n83208 );
xor ( n83780 , n83779 , n83431 );
buf ( n83781 , n83780 );
xor ( n83782 , n77906 , n83211 );
xor ( n83783 , n83782 , n83428 );
buf ( n83784 , n83783 );
xor ( n83785 , n77911 , n83214 );
xor ( n83786 , n83785 , n83425 );
buf ( n83787 , n83786 );
xor ( n83788 , n77916 , n83217 );
xor ( n83789 , n83788 , n83422 );
buf ( n83790 , n83789 );
xor ( n83791 , n77921 , n83220 );
xor ( n83792 , n83791 , n83419 );
buf ( n83793 , n83792 );
xor ( n83794 , n77926 , n83223 );
xor ( n83795 , n83794 , n83416 );
buf ( n83796 , n83795 );
xor ( n83797 , n77931 , n83226 );
xor ( n83798 , n83797 , n83413 );
buf ( n83799 , n83798 );
xor ( n83800 , n77936 , n83229 );
xor ( n83801 , n83800 , n83410 );
buf ( n83802 , n83801 );
xor ( n83803 , n77941 , n83232 );
xor ( n83804 , n83803 , n83407 );
buf ( n83805 , n83804 );
xor ( n83806 , n77946 , n83235 );
xor ( n83807 , n83806 , n83404 );
buf ( n83808 , n83807 );
xor ( n83809 , n77951 , n83238 );
xor ( n83810 , n83809 , n83401 );
buf ( n83811 , n83810 );
xor ( n83812 , n77956 , n83241 );
xor ( n83813 , n83812 , n83398 );
buf ( n83814 , n83813 );
xor ( n83815 , n77961 , n83244 );
xor ( n83816 , n83815 , n83395 );
buf ( n83817 , n83816 );
xor ( n83818 , n77966 , n83247 );
xor ( n83819 , n83818 , n83392 );
buf ( n83820 , n83819 );
xor ( n83821 , n77971 , n83250 );
xor ( n83822 , n83821 , n83389 );
buf ( n83823 , n83822 );
xor ( n83824 , n77976 , n83253 );
xor ( n83825 , n83824 , n83386 );
buf ( n83826 , n83825 );
xor ( n83827 , n77981 , n83256 );
xor ( n83828 , n83827 , n83383 );
buf ( n83829 , n83828 );
xor ( n83830 , n77986 , n83259 );
xor ( n83831 , n83830 , n83380 );
buf ( n83832 , n83831 );
xor ( n83833 , n77991 , n83262 );
xor ( n83834 , n83833 , n83377 );
buf ( n83835 , n83834 );
xor ( n83836 , n77996 , n83265 );
xor ( n83837 , n83836 , n83374 );
buf ( n83838 , n83837 );
xor ( n83839 , n78001 , n83268 );
xor ( n83840 , n83839 , n83371 );
buf ( n83841 , n83840 );
xor ( n83842 , n78006 , n83271 );
xor ( n83843 , n83842 , n83368 );
buf ( n83844 , n83843 );
xor ( n83845 , n78011 , n83274 );
xor ( n83846 , n83845 , n83365 );
buf ( n83847 , n83846 );
xor ( n83848 , n78016 , n83277 );
xor ( n83849 , n83848 , n83362 );
buf ( n83850 , n83849 );
xor ( n83851 , n78021 , n83280 );
xor ( n83852 , n83851 , n83359 );
buf ( n83853 , n83852 );
xor ( n83854 , n78026 , n83283 );
xor ( n83855 , n83854 , n83356 );
buf ( n83856 , n83855 );
xor ( n83857 , n78031 , n83286 );
xor ( n83858 , n83857 , n83353 );
buf ( n83859 , n83858 );
xor ( n83860 , n78036 , n83289 );
xor ( n83861 , n83860 , n83350 );
buf ( n83862 , n83861 );
xor ( n83863 , n78041 , n83292 );
xor ( n83864 , n83863 , n83347 );
buf ( n83865 , n83864 );
xor ( n83866 , n78045 , n83295 );
buf ( n83867 , n83866 );
buf ( n83868 , n83867 );
buf ( n83869 , n83298 );
buf ( n83870 , n83869 );
buf ( n83871 , n18044 );
buf ( n83872 , n18046 );
buf ( n83873 , n18048 );
buf ( n83874 , n18050 );
buf ( n83875 , n18052 );
buf ( n83876 , n18054 );
buf ( n83877 , n18056 );
buf ( n83878 , n18058 );
buf ( n83879 , n18060 );
buf ( n83880 , n18062 );
buf ( n83881 , n18064 );
buf ( n83882 , n18066 );
buf ( n83883 , n18068 );
buf ( n83884 , n18070 );
buf ( n83885 , n18072 );
buf ( n83886 , n18074 );
buf ( n83887 , n18076 );
buf ( n83888 , n18078 );
buf ( n83889 , n18080 );
buf ( n83890 , n18082 );
buf ( n83891 , n18084 );
buf ( n83892 , n18086 );
buf ( n83893 , n18088 );
buf ( n83894 , n18090 );
buf ( n83895 , n18092 );
buf ( n83896 , n18094 );
buf ( n83897 , n18096 );
buf ( n83898 , n578 );
buf ( n83899 , n83898 );
buf ( n83900 , n579 );
buf ( n83901 , n83900 );
buf ( n83902 , n580 );
buf ( n83903 , n83902 );
and ( n83904 , n83901 , n83903 );
not ( n83905 , n83904 );
and ( n83906 , n83899 , n83905 );
not ( n83907 , n83906 );
buf ( n83908 , n545 );
buf ( n83909 , n83908 );
buf ( n83910 , n576 );
buf ( n83911 , n83910 );
buf ( n83912 , n577 );
buf ( n83913 , n83912 );
xor ( n83914 , n83911 , n83913 );
xor ( n83915 , n83913 , n83899 );
not ( n83916 , n83915 );
and ( n83917 , n83914 , n83916 );
and ( n83918 , n83909 , n83917 );
buf ( n83919 , n544 );
buf ( n83920 , n83919 );
and ( n83921 , n83920 , n83915 );
nor ( n83922 , n83918 , n83921 );
and ( n83923 , n83913 , n83899 );
not ( n83924 , n83923 );
and ( n83925 , n83911 , n83924 );
xnor ( n83926 , n83922 , n83925 );
and ( n83927 , n83907 , n83926 );
buf ( n83928 , n546 );
buf ( n83929 , n83928 );
and ( n83930 , n83929 , n83911 );
and ( n83931 , n83926 , n83930 );
and ( n83932 , n83907 , n83930 );
or ( n83933 , n83927 , n83931 , n83932 );
and ( n83934 , n83920 , n83917 );
not ( n83935 , n83934 );
xnor ( n83936 , n83935 , n83925 );
and ( n83937 , n83933 , n83936 );
and ( n83938 , n83909 , n83911 );
not ( n83939 , n83938 );
and ( n83940 , n83936 , n83939 );
and ( n83941 , n83933 , n83939 );
or ( n83942 , n83937 , n83940 , n83941 );
xor ( n83943 , n83899 , n83901 );
xor ( n83944 , n83901 , n83903 );
not ( n83945 , n83944 );
and ( n83946 , n83943 , n83945 );
and ( n83947 , n83920 , n83946 );
not ( n83948 , n83947 );
xnor ( n83949 , n83948 , n83906 );
not ( n83950 , n83949 );
and ( n83951 , n83929 , n83917 );
and ( n83952 , n83909 , n83915 );
nor ( n83953 , n83951 , n83952 );
xnor ( n83954 , n83953 , n83925 );
and ( n83955 , n83950 , n83954 );
buf ( n83956 , n547 );
buf ( n83957 , n83956 );
and ( n83958 , n83957 , n83911 );
and ( n83959 , n83954 , n83958 );
and ( n83960 , n83950 , n83958 );
or ( n83961 , n83955 , n83959 , n83960 );
buf ( n83962 , n83949 );
and ( n83963 , n83961 , n83962 );
xor ( n83964 , n83907 , n83926 );
xor ( n83965 , n83964 , n83930 );
and ( n83966 , n83962 , n83965 );
and ( n83967 , n83961 , n83965 );
or ( n83968 , n83963 , n83966 , n83967 );
buf ( n83969 , n83871 );
and ( n83970 , n83968 , n83969 );
xor ( n83971 , n83933 , n83936 );
xor ( n83972 , n83971 , n83939 );
and ( n83973 , n83969 , n83972 );
and ( n83974 , n83968 , n83972 );
or ( n83975 , n83970 , n83973 , n83974 );
xor ( n83976 , n83942 , n83975 );
buf ( n83977 , n83938 );
not ( n83978 , n83925 );
xor ( n83979 , n83977 , n83978 );
and ( n83980 , n83920 , n83911 );
xor ( n83981 , n83979 , n83980 );
xor ( n83982 , n83976 , n83981 );
xor ( n83983 , n83968 , n83969 );
xor ( n83984 , n83983 , n83972 );
buf ( n83985 , n581 );
buf ( n83986 , n83985 );
buf ( n83987 , n582 );
buf ( n83988 , n83987 );
and ( n83989 , n83986 , n83988 );
not ( n83990 , n83989 );
and ( n83991 , n83903 , n83990 );
not ( n83992 , n83991 );
and ( n83993 , n83909 , n83946 );
and ( n83994 , n83920 , n83944 );
nor ( n83995 , n83993 , n83994 );
xnor ( n83996 , n83995 , n83906 );
and ( n83997 , n83992 , n83996 );
buf ( n83998 , n548 );
buf ( n83999 , n83998 );
and ( n84000 , n83999 , n83911 );
and ( n84001 , n83996 , n84000 );
and ( n84002 , n83992 , n84000 );
or ( n84003 , n83997 , n84001 , n84002 );
and ( n84004 , n83929 , n83946 );
and ( n84005 , n83909 , n83944 );
nor ( n84006 , n84004 , n84005 );
xnor ( n84007 , n84006 , n83906 );
and ( n84008 , n83999 , n83917 );
and ( n84009 , n83957 , n83915 );
nor ( n84010 , n84008 , n84009 );
xnor ( n84011 , n84010 , n83925 );
and ( n84012 , n84007 , n84011 );
buf ( n84013 , n549 );
buf ( n84014 , n84013 );
and ( n84015 , n84014 , n83911 );
and ( n84016 , n84011 , n84015 );
and ( n84017 , n84007 , n84015 );
or ( n84018 , n84012 , n84016 , n84017 );
xor ( n84019 , n83903 , n83986 );
xor ( n84020 , n83986 , n83988 );
not ( n84021 , n84020 );
and ( n84022 , n84019 , n84021 );
and ( n84023 , n83920 , n84022 );
not ( n84024 , n84023 );
xnor ( n84025 , n84024 , n83991 );
buf ( n84026 , n84025 );
and ( n84027 , n84018 , n84026 );
and ( n84028 , n83957 , n83917 );
and ( n84029 , n83929 , n83915 );
nor ( n84030 , n84028 , n84029 );
xnor ( n84031 , n84030 , n83925 );
and ( n84032 , n84026 , n84031 );
and ( n84033 , n84018 , n84031 );
or ( n84034 , n84027 , n84032 , n84033 );
and ( n84035 , n84003 , n84034 );
xor ( n84036 , n83950 , n83954 );
xor ( n84037 , n84036 , n83958 );
and ( n84038 , n84034 , n84037 );
and ( n84039 , n84003 , n84037 );
or ( n84040 , n84035 , n84038 , n84039 );
buf ( n84041 , n83872 );
and ( n84042 , n84040 , n84041 );
xor ( n84043 , n83961 , n83962 );
xor ( n84044 , n84043 , n83965 );
and ( n84045 , n84041 , n84044 );
and ( n84046 , n84040 , n84044 );
or ( n84047 , n84042 , n84045 , n84046 );
and ( n84048 , n83984 , n84047 );
xor ( n84049 , n83984 , n84047 );
xor ( n84050 , n84040 , n84041 );
xor ( n84051 , n84050 , n84044 );
buf ( n84052 , n583 );
buf ( n84053 , n84052 );
buf ( n84054 , n584 );
buf ( n84055 , n84054 );
and ( n84056 , n84053 , n84055 );
not ( n84057 , n84056 );
and ( n84058 , n83988 , n84057 );
not ( n84059 , n84058 );
and ( n84060 , n83909 , n84022 );
and ( n84061 , n83920 , n84020 );
nor ( n84062 , n84060 , n84061 );
xnor ( n84063 , n84062 , n83991 );
and ( n84064 , n84059 , n84063 );
and ( n84065 , n84014 , n83917 );
and ( n84066 , n83999 , n83915 );
nor ( n84067 , n84065 , n84066 );
xnor ( n84068 , n84067 , n83925 );
and ( n84069 , n84063 , n84068 );
and ( n84070 , n84059 , n84068 );
or ( n84071 , n84064 , n84069 , n84070 );
not ( n84072 , n84025 );
and ( n84073 , n84071 , n84072 );
xor ( n84074 , n84007 , n84011 );
xor ( n84075 , n84074 , n84015 );
and ( n84076 , n84072 , n84075 );
and ( n84077 , n84071 , n84075 );
or ( n84078 , n84073 , n84076 , n84077 );
xor ( n84079 , n83992 , n83996 );
xor ( n84080 , n84079 , n84000 );
and ( n84081 , n84078 , n84080 );
xor ( n84082 , n84018 , n84026 );
xor ( n84083 , n84082 , n84031 );
and ( n84084 , n84080 , n84083 );
and ( n84085 , n84078 , n84083 );
or ( n84086 , n84081 , n84084 , n84085 );
buf ( n84087 , n83873 );
and ( n84088 , n84086 , n84087 );
xor ( n84089 , n84003 , n84034 );
xor ( n84090 , n84089 , n84037 );
and ( n84091 , n84087 , n84090 );
and ( n84092 , n84086 , n84090 );
or ( n84093 , n84088 , n84091 , n84092 );
and ( n84094 , n84051 , n84093 );
xor ( n84095 , n84051 , n84093 );
xor ( n84096 , n84086 , n84087 );
xor ( n84097 , n84096 , n84090 );
and ( n84098 , n83929 , n84022 );
and ( n84099 , n83909 , n84020 );
nor ( n84100 , n84098 , n84099 );
xnor ( n84101 , n84100 , n83991 );
buf ( n84102 , n84101 );
and ( n84103 , n83957 , n83946 );
and ( n84104 , n83929 , n83944 );
nor ( n84105 , n84103 , n84104 );
xnor ( n84106 , n84105 , n83906 );
and ( n84107 , n84102 , n84106 );
buf ( n84108 , n550 );
buf ( n84109 , n84108 );
and ( n84110 , n84109 , n83911 );
and ( n84111 , n84106 , n84110 );
and ( n84112 , n84102 , n84110 );
or ( n84113 , n84107 , n84111 , n84112 );
xor ( n84114 , n83988 , n84053 );
xor ( n84115 , n84053 , n84055 );
not ( n84116 , n84115 );
and ( n84117 , n84114 , n84116 );
and ( n84118 , n83920 , n84117 );
not ( n84119 , n84118 );
xnor ( n84120 , n84119 , n84058 );
and ( n84121 , n84109 , n83917 );
and ( n84122 , n84014 , n83915 );
nor ( n84123 , n84121 , n84122 );
xnor ( n84124 , n84123 , n83925 );
and ( n84125 , n84120 , n84124 );
buf ( n84126 , n551 );
buf ( n84127 , n84126 );
and ( n84128 , n84127 , n83911 );
and ( n84129 , n84124 , n84128 );
and ( n84130 , n84120 , n84128 );
or ( n84131 , n84125 , n84129 , n84130 );
xor ( n84132 , n84059 , n84063 );
xor ( n84133 , n84132 , n84068 );
and ( n84134 , n84131 , n84133 );
xor ( n84135 , n84102 , n84106 );
xor ( n84136 , n84135 , n84110 );
and ( n84137 , n84133 , n84136 );
and ( n84138 , n84131 , n84136 );
or ( n84139 , n84134 , n84137 , n84138 );
and ( n84140 , n84113 , n84139 );
xor ( n84141 , n84071 , n84072 );
xor ( n84142 , n84141 , n84075 );
and ( n84143 , n84139 , n84142 );
and ( n84144 , n84113 , n84142 );
or ( n84145 , n84140 , n84143 , n84144 );
buf ( n84146 , n83874 );
and ( n84147 , n84145 , n84146 );
xor ( n84148 , n84078 , n84080 );
xor ( n84149 , n84148 , n84083 );
and ( n84150 , n84146 , n84149 );
and ( n84151 , n84145 , n84149 );
or ( n84152 , n84147 , n84150 , n84151 );
and ( n84153 , n84097 , n84152 );
xor ( n84154 , n84097 , n84152 );
xor ( n84155 , n84145 , n84146 );
xor ( n84156 , n84155 , n84149 );
and ( n84157 , n83957 , n84022 );
and ( n84158 , n83929 , n84020 );
nor ( n84159 , n84157 , n84158 );
xnor ( n84160 , n84159 , n83991 );
and ( n84161 , n84127 , n83917 );
and ( n84162 , n84109 , n83915 );
nor ( n84163 , n84161 , n84162 );
xnor ( n84164 , n84163 , n83925 );
and ( n84165 , n84160 , n84164 );
buf ( n84166 , n552 );
buf ( n84167 , n84166 );
and ( n84168 , n84167 , n83911 );
and ( n84169 , n84164 , n84168 );
and ( n84170 , n84160 , n84168 );
or ( n84171 , n84165 , n84169 , n84170 );
not ( n84172 , n84101 );
and ( n84173 , n84171 , n84172 );
and ( n84174 , n83999 , n83946 );
and ( n84175 , n83957 , n83944 );
nor ( n84176 , n84174 , n84175 );
xnor ( n84177 , n84176 , n83906 );
and ( n84178 , n84172 , n84177 );
and ( n84179 , n84171 , n84177 );
or ( n84180 , n84173 , n84178 , n84179 );
buf ( n84181 , n585 );
buf ( n84182 , n84181 );
buf ( n84183 , n586 );
buf ( n84184 , n84183 );
and ( n84185 , n84182 , n84184 );
not ( n84186 , n84185 );
and ( n84187 , n84055 , n84186 );
not ( n84188 , n84187 );
and ( n84189 , n83909 , n84117 );
and ( n84190 , n83920 , n84115 );
nor ( n84191 , n84189 , n84190 );
xnor ( n84192 , n84191 , n84058 );
and ( n84193 , n84188 , n84192 );
and ( n84194 , n84014 , n83946 );
and ( n84195 , n83999 , n83944 );
nor ( n84196 , n84194 , n84195 );
xnor ( n84197 , n84196 , n83906 );
and ( n84198 , n84192 , n84197 );
and ( n84199 , n84188 , n84197 );
or ( n84200 , n84193 , n84198 , n84199 );
xor ( n84201 , n84120 , n84124 );
xor ( n84202 , n84201 , n84128 );
and ( n84203 , n84200 , n84202 );
xor ( n84204 , n84171 , n84172 );
xor ( n84205 , n84204 , n84177 );
and ( n84206 , n84202 , n84205 );
and ( n84207 , n84200 , n84205 );
or ( n84208 , n84203 , n84206 , n84207 );
and ( n84209 , n84180 , n84208 );
xor ( n84210 , n84131 , n84133 );
xor ( n84211 , n84210 , n84136 );
and ( n84212 , n84208 , n84211 );
and ( n84213 , n84180 , n84211 );
or ( n84214 , n84209 , n84212 , n84213 );
buf ( n84215 , n83875 );
and ( n84216 , n84214 , n84215 );
xor ( n84217 , n84113 , n84139 );
xor ( n84218 , n84217 , n84142 );
and ( n84219 , n84215 , n84218 );
and ( n84220 , n84214 , n84218 );
or ( n84221 , n84216 , n84219 , n84220 );
and ( n84222 , n84156 , n84221 );
xor ( n84223 , n84156 , n84221 );
xor ( n84224 , n84214 , n84215 );
xor ( n84225 , n84224 , n84218 );
xor ( n84226 , n84055 , n84182 );
xor ( n84227 , n84182 , n84184 );
not ( n84228 , n84227 );
and ( n84229 , n84226 , n84228 );
and ( n84230 , n83920 , n84229 );
not ( n84231 , n84230 );
xnor ( n84232 , n84231 , n84187 );
and ( n84233 , n84109 , n83946 );
and ( n84234 , n84014 , n83944 );
nor ( n84235 , n84233 , n84234 );
xnor ( n84236 , n84235 , n83906 );
and ( n84237 , n84232 , n84236 );
and ( n84238 , n84167 , n83917 );
and ( n84239 , n84127 , n83915 );
nor ( n84240 , n84238 , n84239 );
xnor ( n84241 , n84240 , n83925 );
and ( n84242 , n84236 , n84241 );
and ( n84243 , n84232 , n84241 );
or ( n84244 , n84237 , n84242 , n84243 );
and ( n84245 , n83929 , n84117 );
and ( n84246 , n83909 , n84115 );
nor ( n84247 , n84245 , n84246 );
xnor ( n84248 , n84247 , n84058 );
buf ( n84249 , n84248 );
and ( n84250 , n84244 , n84249 );
xor ( n84251 , n84160 , n84164 );
xor ( n84252 , n84251 , n84168 );
and ( n84253 , n84249 , n84252 );
and ( n84254 , n84244 , n84252 );
or ( n84255 , n84250 , n84253 , n84254 );
not ( n84256 , n84248 );
and ( n84257 , n83999 , n84022 );
and ( n84258 , n83957 , n84020 );
nor ( n84259 , n84257 , n84258 );
xnor ( n84260 , n84259 , n83991 );
and ( n84261 , n84256 , n84260 );
buf ( n84262 , n553 );
buf ( n84263 , n84262 );
and ( n84264 , n84263 , n83911 );
and ( n84265 , n84260 , n84264 );
and ( n84266 , n84256 , n84264 );
or ( n84267 , n84261 , n84265 , n84266 );
xor ( n84268 , n84188 , n84192 );
xor ( n84269 , n84268 , n84197 );
and ( n84270 , n84267 , n84269 );
xor ( n84271 , n84244 , n84249 );
xor ( n84272 , n84271 , n84252 );
and ( n84273 , n84269 , n84272 );
and ( n84274 , n84267 , n84272 );
or ( n84275 , n84270 , n84273 , n84274 );
and ( n84276 , n84255 , n84275 );
xor ( n84277 , n84200 , n84202 );
xor ( n84278 , n84277 , n84205 );
and ( n84279 , n84275 , n84278 );
and ( n84280 , n84255 , n84278 );
or ( n84281 , n84276 , n84279 , n84280 );
buf ( n84282 , n83876 );
and ( n84283 , n84281 , n84282 );
xor ( n84284 , n84180 , n84208 );
xor ( n84285 , n84284 , n84211 );
and ( n84286 , n84282 , n84285 );
and ( n84287 , n84281 , n84285 );
or ( n84288 , n84283 , n84286 , n84287 );
and ( n84289 , n84225 , n84288 );
xor ( n84290 , n84225 , n84288 );
xor ( n84291 , n84281 , n84282 );
xor ( n84292 , n84291 , n84285 );
buf ( n84293 , n587 );
buf ( n84294 , n84293 );
buf ( n84295 , n588 );
buf ( n84296 , n84295 );
and ( n84297 , n84294 , n84296 );
not ( n84298 , n84297 );
and ( n84299 , n84184 , n84298 );
not ( n84300 , n84299 );
and ( n84301 , n83909 , n84229 );
and ( n84302 , n83920 , n84227 );
nor ( n84303 , n84301 , n84302 );
xnor ( n84304 , n84303 , n84187 );
and ( n84305 , n84300 , n84304 );
and ( n84306 , n84014 , n84022 );
and ( n84307 , n83999 , n84020 );
nor ( n84308 , n84306 , n84307 );
xnor ( n84309 , n84308 , n83991 );
and ( n84310 , n84304 , n84309 );
and ( n84311 , n84300 , n84309 );
or ( n84312 , n84305 , n84310 , n84311 );
and ( n84313 , n83957 , n84117 );
and ( n84314 , n83929 , n84115 );
nor ( n84315 , n84313 , n84314 );
xnor ( n84316 , n84315 , n84058 );
and ( n84317 , n84127 , n83946 );
and ( n84318 , n84109 , n83944 );
nor ( n84319 , n84317 , n84318 );
xnor ( n84320 , n84319 , n83906 );
and ( n84321 , n84316 , n84320 );
and ( n84322 , n84263 , n83917 );
and ( n84323 , n84167 , n83915 );
nor ( n84324 , n84322 , n84323 );
xnor ( n84325 , n84324 , n83925 );
and ( n84326 , n84320 , n84325 );
and ( n84327 , n84316 , n84325 );
or ( n84328 , n84321 , n84326 , n84327 );
and ( n84329 , n84312 , n84328 );
xor ( n84330 , n84232 , n84236 );
xor ( n84331 , n84330 , n84241 );
and ( n84332 , n84328 , n84331 );
and ( n84333 , n84312 , n84331 );
or ( n84334 , n84329 , n84332 , n84333 );
and ( n84335 , n83929 , n84229 );
and ( n84336 , n83909 , n84227 );
nor ( n84337 , n84335 , n84336 );
xnor ( n84338 , n84337 , n84187 );
and ( n84339 , n84109 , n84022 );
and ( n84340 , n84014 , n84020 );
nor ( n84341 , n84339 , n84340 );
xnor ( n84342 , n84341 , n83991 );
and ( n84343 , n84338 , n84342 );
and ( n84344 , n84167 , n83946 );
and ( n84345 , n84127 , n83944 );
nor ( n84346 , n84344 , n84345 );
xnor ( n84347 , n84346 , n83906 );
and ( n84348 , n84342 , n84347 );
and ( n84349 , n84338 , n84347 );
or ( n84350 , n84343 , n84348 , n84349 );
xor ( n84351 , n84184 , n84294 );
xor ( n84352 , n84294 , n84296 );
not ( n84353 , n84352 );
and ( n84354 , n84351 , n84353 );
and ( n84355 , n83920 , n84354 );
not ( n84356 , n84355 );
xnor ( n84357 , n84356 , n84299 );
buf ( n84358 , n84357 );
and ( n84359 , n84350 , n84358 );
buf ( n84360 , n554 );
buf ( n84361 , n84360 );
and ( n84362 , n84361 , n83911 );
and ( n84363 , n84358 , n84362 );
and ( n84364 , n84350 , n84362 );
or ( n84365 , n84359 , n84363 , n84364 );
and ( n84366 , n83999 , n84117 );
and ( n84367 , n83957 , n84115 );
nor ( n84368 , n84366 , n84367 );
xnor ( n84369 , n84368 , n84058 );
and ( n84370 , n84361 , n83917 );
and ( n84371 , n84263 , n83915 );
nor ( n84372 , n84370 , n84371 );
xnor ( n84373 , n84372 , n83925 );
and ( n84374 , n84369 , n84373 );
buf ( n84375 , n555 );
buf ( n84376 , n84375 );
and ( n84377 , n84376 , n83911 );
and ( n84378 , n84373 , n84377 );
and ( n84379 , n84369 , n84377 );
or ( n84380 , n84374 , n84378 , n84379 );
xor ( n84381 , n84300 , n84304 );
xor ( n84382 , n84381 , n84309 );
and ( n84383 , n84380 , n84382 );
xor ( n84384 , n84316 , n84320 );
xor ( n84385 , n84384 , n84325 );
and ( n84386 , n84382 , n84385 );
and ( n84387 , n84380 , n84385 );
or ( n84388 , n84383 , n84386 , n84387 );
and ( n84389 , n84365 , n84388 );
xor ( n84390 , n84256 , n84260 );
xor ( n84391 , n84390 , n84264 );
and ( n84392 , n84388 , n84391 );
and ( n84393 , n84365 , n84391 );
or ( n84394 , n84389 , n84392 , n84393 );
and ( n84395 , n84334 , n84394 );
xor ( n84396 , n84267 , n84269 );
xor ( n84397 , n84396 , n84272 );
and ( n84398 , n84394 , n84397 );
and ( n84399 , n84334 , n84397 );
or ( n84400 , n84395 , n84398 , n84399 );
buf ( n84401 , n83877 );
and ( n84402 , n84400 , n84401 );
xor ( n84403 , n84255 , n84275 );
xor ( n84404 , n84403 , n84278 );
and ( n84405 , n84401 , n84404 );
and ( n84406 , n84400 , n84404 );
or ( n84407 , n84402 , n84405 , n84406 );
and ( n84408 , n84292 , n84407 );
xor ( n84409 , n84292 , n84407 );
xor ( n84410 , n84400 , n84401 );
xor ( n84411 , n84410 , n84404 );
and ( n84412 , n83957 , n84229 );
and ( n84413 , n83929 , n84227 );
nor ( n84414 , n84412 , n84413 );
xnor ( n84415 , n84414 , n84187 );
and ( n84416 , n84127 , n84022 );
and ( n84417 , n84109 , n84020 );
nor ( n84418 , n84416 , n84417 );
xnor ( n84419 , n84418 , n83991 );
and ( n84420 , n84415 , n84419 );
buf ( n84421 , n556 );
buf ( n84422 , n84421 );
and ( n84423 , n84422 , n83911 );
and ( n84424 , n84419 , n84423 );
and ( n84425 , n84415 , n84423 );
or ( n84426 , n84420 , n84424 , n84425 );
buf ( n84427 , n589 );
buf ( n84428 , n84427 );
buf ( n84429 , n590 );
buf ( n84430 , n84429 );
and ( n84431 , n84428 , n84430 );
not ( n84432 , n84431 );
and ( n84433 , n84296 , n84432 );
not ( n84434 , n84433 );
and ( n84435 , n83909 , n84354 );
and ( n84436 , n83920 , n84352 );
nor ( n84437 , n84435 , n84436 );
xnor ( n84438 , n84437 , n84299 );
and ( n84439 , n84434 , n84438 );
and ( n84440 , n84014 , n84117 );
and ( n84441 , n83999 , n84115 );
nor ( n84442 , n84440 , n84441 );
xnor ( n84443 , n84442 , n84058 );
and ( n84444 , n84438 , n84443 );
and ( n84445 , n84434 , n84443 );
or ( n84446 , n84439 , n84444 , n84445 );
and ( n84447 , n84426 , n84446 );
not ( n84448 , n84357 );
and ( n84449 , n84446 , n84448 );
and ( n84450 , n84426 , n84448 );
or ( n84451 , n84447 , n84449 , n84450 );
xor ( n84452 , n84296 , n84428 );
xor ( n84453 , n84428 , n84430 );
not ( n84454 , n84453 );
and ( n84455 , n84452 , n84454 );
and ( n84456 , n83920 , n84455 );
not ( n84457 , n84456 );
xnor ( n84458 , n84457 , n84433 );
buf ( n84459 , n84458 );
and ( n84460 , n84263 , n83946 );
and ( n84461 , n84167 , n83944 );
nor ( n84462 , n84460 , n84461 );
xnor ( n84463 , n84462 , n83906 );
and ( n84464 , n84459 , n84463 );
and ( n84465 , n84376 , n83917 );
and ( n84466 , n84361 , n83915 );
nor ( n84467 , n84465 , n84466 );
xnor ( n84468 , n84467 , n83925 );
and ( n84469 , n84463 , n84468 );
and ( n84470 , n84459 , n84468 );
or ( n84471 , n84464 , n84469 , n84470 );
xor ( n84472 , n84369 , n84373 );
xor ( n84473 , n84472 , n84377 );
and ( n84474 , n84471 , n84473 );
xor ( n84475 , n84338 , n84342 );
xor ( n84476 , n84475 , n84347 );
and ( n84477 , n84473 , n84476 );
and ( n84478 , n84471 , n84476 );
or ( n84479 , n84474 , n84477 , n84478 );
and ( n84480 , n84451 , n84479 );
xor ( n84481 , n84350 , n84358 );
xor ( n84482 , n84481 , n84362 );
and ( n84483 , n84479 , n84482 );
and ( n84484 , n84451 , n84482 );
or ( n84485 , n84480 , n84483 , n84484 );
xor ( n84486 , n84312 , n84328 );
xor ( n84487 , n84486 , n84331 );
and ( n84488 , n84485 , n84487 );
xor ( n84489 , n84365 , n84388 );
xor ( n84490 , n84489 , n84391 );
and ( n84491 , n84487 , n84490 );
and ( n84492 , n84485 , n84490 );
or ( n84493 , n84488 , n84491 , n84492 );
buf ( n84494 , n83878 );
and ( n84495 , n84493 , n84494 );
xor ( n84496 , n84334 , n84394 );
xor ( n84497 , n84496 , n84397 );
and ( n84498 , n84494 , n84497 );
and ( n84499 , n84493 , n84497 );
or ( n84500 , n84495 , n84498 , n84499 );
and ( n84501 , n84411 , n84500 );
xor ( n84502 , n84411 , n84500 );
xor ( n84503 , n84493 , n84494 );
xor ( n84504 , n84503 , n84497 );
and ( n84505 , n83929 , n84354 );
and ( n84506 , n83909 , n84352 );
nor ( n84507 , n84505 , n84506 );
xnor ( n84508 , n84507 , n84299 );
and ( n84509 , n84109 , n84117 );
and ( n84510 , n84014 , n84115 );
nor ( n84511 , n84509 , n84510 );
xnor ( n84512 , n84511 , n84058 );
and ( n84513 , n84508 , n84512 );
buf ( n84514 , n557 );
buf ( n84515 , n84514 );
and ( n84516 , n84515 , n83911 );
and ( n84517 , n84512 , n84516 );
and ( n84518 , n84508 , n84516 );
or ( n84519 , n84513 , n84517 , n84518 );
and ( n84520 , n83999 , n84229 );
and ( n84521 , n83957 , n84227 );
nor ( n84522 , n84520 , n84521 );
xnor ( n84523 , n84522 , n84187 );
and ( n84524 , n84167 , n84022 );
and ( n84525 , n84127 , n84020 );
nor ( n84526 , n84524 , n84525 );
xnor ( n84527 , n84526 , n83991 );
and ( n84528 , n84523 , n84527 );
and ( n84529 , n84361 , n83946 );
and ( n84530 , n84263 , n83944 );
nor ( n84531 , n84529 , n84530 );
xnor ( n84532 , n84531 , n83906 );
and ( n84533 , n84527 , n84532 );
and ( n84534 , n84523 , n84532 );
or ( n84535 , n84528 , n84533 , n84534 );
and ( n84536 , n84519 , n84535 );
xor ( n84537 , n84434 , n84438 );
xor ( n84538 , n84537 , n84443 );
and ( n84539 , n84535 , n84538 );
and ( n84540 , n84519 , n84538 );
or ( n84541 , n84536 , n84539 , n84540 );
xor ( n84542 , n84426 , n84446 );
xor ( n84543 , n84542 , n84448 );
and ( n84544 , n84541 , n84543 );
xor ( n84545 , n84471 , n84473 );
xor ( n84546 , n84545 , n84476 );
and ( n84547 , n84543 , n84546 );
and ( n84548 , n84541 , n84546 );
or ( n84549 , n84544 , n84547 , n84548 );
xor ( n84550 , n84380 , n84382 );
xor ( n84551 , n84550 , n84385 );
and ( n84552 , n84549 , n84551 );
xor ( n84553 , n84451 , n84479 );
xor ( n84554 , n84553 , n84482 );
and ( n84555 , n84551 , n84554 );
and ( n84556 , n84549 , n84554 );
or ( n84557 , n84552 , n84555 , n84556 );
buf ( n84558 , n83879 );
and ( n84559 , n84557 , n84558 );
xor ( n84560 , n84485 , n84487 );
xor ( n84561 , n84560 , n84490 );
and ( n84562 , n84558 , n84561 );
and ( n84563 , n84557 , n84561 );
or ( n84564 , n84559 , n84562 , n84563 );
and ( n84565 , n84504 , n84564 );
xor ( n84566 , n84504 , n84564 );
xor ( n84567 , n84557 , n84558 );
xor ( n84568 , n84567 , n84561 );
and ( n84569 , n84014 , n84229 );
and ( n84570 , n83999 , n84227 );
nor ( n84571 , n84569 , n84570 );
xnor ( n84572 , n84571 , n84187 );
buf ( n84573 , n84572 );
not ( n84574 , n84458 );
and ( n84575 , n84573 , n84574 );
and ( n84576 , n84422 , n83917 );
and ( n84577 , n84376 , n83915 );
nor ( n84578 , n84576 , n84577 );
xnor ( n84579 , n84578 , n83925 );
and ( n84580 , n84574 , n84579 );
and ( n84581 , n84573 , n84579 );
or ( n84582 , n84575 , n84580 , n84581 );
xor ( n84583 , n84415 , n84419 );
xor ( n84584 , n84583 , n84423 );
and ( n84585 , n84582 , n84584 );
xor ( n84586 , n84459 , n84463 );
xor ( n84587 , n84586 , n84468 );
and ( n84588 , n84584 , n84587 );
and ( n84589 , n84582 , n84587 );
or ( n84590 , n84585 , n84588 , n84589 );
not ( n84591 , n84430 );
and ( n84592 , n84515 , n83917 );
and ( n84593 , n84422 , n83915 );
nor ( n84594 , n84592 , n84593 );
xnor ( n84595 , n84594 , n83925 );
and ( n84596 , n84591 , n84595 );
buf ( n84597 , n558 );
buf ( n84598 , n84597 );
and ( n84599 , n84598 , n83911 );
and ( n84600 , n84595 , n84599 );
and ( n84601 , n84591 , n84599 );
or ( n84602 , n84596 , n84600 , n84601 );
and ( n84603 , n83909 , n84455 );
and ( n84604 , n83920 , n84453 );
nor ( n84605 , n84603 , n84604 );
xnor ( n84606 , n84605 , n84433 );
and ( n84607 , n83957 , n84354 );
and ( n84608 , n83929 , n84352 );
nor ( n84609 , n84607 , n84608 );
xnor ( n84610 , n84609 , n84299 );
and ( n84611 , n84606 , n84610 );
and ( n84612 , n84127 , n84117 );
and ( n84613 , n84109 , n84115 );
nor ( n84614 , n84612 , n84613 );
xnor ( n84615 , n84614 , n84058 );
and ( n84616 , n84610 , n84615 );
and ( n84617 , n84606 , n84615 );
or ( n84618 , n84611 , n84616 , n84617 );
and ( n84619 , n84602 , n84618 );
xor ( n84620 , n84523 , n84527 );
xor ( n84621 , n84620 , n84532 );
and ( n84622 , n84618 , n84621 );
and ( n84623 , n84602 , n84621 );
or ( n84624 , n84619 , n84622 , n84623 );
and ( n84625 , n83999 , n84354 );
and ( n84626 , n83957 , n84352 );
nor ( n84627 , n84625 , n84626 );
xnor ( n84628 , n84627 , n84299 );
and ( n84629 , n84361 , n84022 );
and ( n84630 , n84263 , n84020 );
nor ( n84631 , n84629 , n84630 );
xnor ( n84632 , n84631 , n83991 );
and ( n84633 , n84628 , n84632 );
and ( n84634 , n84422 , n83946 );
and ( n84635 , n84376 , n83944 );
nor ( n84636 , n84634 , n84635 );
xnor ( n84637 , n84636 , n83906 );
and ( n84638 , n84632 , n84637 );
and ( n84639 , n84628 , n84637 );
or ( n84640 , n84633 , n84638 , n84639 );
buf ( n84641 , n591 );
buf ( n84642 , n84641 );
xor ( n84643 , n84430 , n84642 );
not ( n84644 , n84642 );
and ( n84645 , n84643 , n84644 );
and ( n84646 , n83920 , n84645 );
not ( n84647 , n84646 );
xnor ( n84648 , n84647 , n84430 );
and ( n84649 , n83929 , n84455 );
and ( n84650 , n83909 , n84453 );
nor ( n84651 , n84649 , n84650 );
xnor ( n84652 , n84651 , n84433 );
and ( n84653 , n84648 , n84652 );
buf ( n84654 , n559 );
buf ( n84655 , n84654 );
and ( n84656 , n84655 , n83911 );
and ( n84657 , n84652 , n84656 );
and ( n84658 , n84648 , n84656 );
or ( n84659 , n84653 , n84657 , n84658 );
and ( n84660 , n84640 , n84659 );
and ( n84661 , n84109 , n84229 );
and ( n84662 , n84014 , n84227 );
nor ( n84663 , n84661 , n84662 );
xnor ( n84664 , n84663 , n84187 );
and ( n84665 , n84167 , n84117 );
and ( n84666 , n84127 , n84115 );
nor ( n84667 , n84665 , n84666 );
xnor ( n84668 , n84667 , n84058 );
and ( n84669 , n84664 , n84668 );
and ( n84670 , n84598 , n83917 );
and ( n84671 , n84515 , n83915 );
nor ( n84672 , n84670 , n84671 );
xnor ( n84673 , n84672 , n83925 );
and ( n84674 , n84668 , n84673 );
and ( n84675 , n84664 , n84673 );
or ( n84676 , n84669 , n84674 , n84675 );
and ( n84677 , n84659 , n84676 );
and ( n84678 , n84640 , n84676 );
or ( n84679 , n84660 , n84677 , n84678 );
xor ( n84680 , n84508 , n84512 );
xor ( n84681 , n84680 , n84516 );
and ( n84682 , n84679 , n84681 );
xor ( n84683 , n84573 , n84574 );
xor ( n84684 , n84683 , n84579 );
and ( n84685 , n84681 , n84684 );
and ( n84686 , n84679 , n84684 );
or ( n84687 , n84682 , n84685 , n84686 );
and ( n84688 , n84624 , n84687 );
xor ( n84689 , n84519 , n84535 );
xor ( n84690 , n84689 , n84538 );
and ( n84691 , n84687 , n84690 );
and ( n84692 , n84624 , n84690 );
or ( n84693 , n84688 , n84691 , n84692 );
and ( n84694 , n84590 , n84693 );
xor ( n84695 , n84541 , n84543 );
xor ( n84696 , n84695 , n84546 );
and ( n84697 , n84693 , n84696 );
and ( n84698 , n84590 , n84696 );
or ( n84699 , n84694 , n84697 , n84698 );
buf ( n84700 , n83880 );
and ( n84701 , n84699 , n84700 );
xor ( n84702 , n84549 , n84551 );
xor ( n84703 , n84702 , n84554 );
and ( n84704 , n84700 , n84703 );
and ( n84705 , n84699 , n84703 );
or ( n84706 , n84701 , n84704 , n84705 );
and ( n84707 , n84568 , n84706 );
xor ( n84708 , n84568 , n84706 );
xor ( n84709 , n84699 , n84700 );
xor ( n84710 , n84709 , n84703 );
not ( n84711 , n84572 );
and ( n84712 , n84263 , n84022 );
and ( n84713 , n84167 , n84020 );
nor ( n84714 , n84712 , n84713 );
xnor ( n84715 , n84714 , n83991 );
and ( n84716 , n84711 , n84715 );
and ( n84717 , n84376 , n83946 );
and ( n84718 , n84361 , n83944 );
nor ( n84719 , n84717 , n84718 );
xnor ( n84720 , n84719 , n83906 );
and ( n84721 , n84715 , n84720 );
and ( n84722 , n84711 , n84720 );
or ( n84723 , n84716 , n84721 , n84722 );
and ( n84724 , n84014 , n84354 );
and ( n84725 , n83999 , n84352 );
nor ( n84726 , n84724 , n84725 );
xnor ( n84727 , n84726 , n84299 );
and ( n84728 , n84263 , n84117 );
and ( n84729 , n84167 , n84115 );
nor ( n84730 , n84728 , n84729 );
xnor ( n84731 , n84730 , n84058 );
and ( n84732 , n84727 , n84731 );
and ( n84733 , n84376 , n84022 );
and ( n84734 , n84361 , n84020 );
nor ( n84735 , n84733 , n84734 );
xnor ( n84736 , n84735 , n83991 );
and ( n84737 , n84731 , n84736 );
and ( n84738 , n84727 , n84736 );
or ( n84739 , n84732 , n84737 , n84738 );
and ( n84740 , n83957 , n84455 );
and ( n84741 , n83929 , n84453 );
nor ( n84742 , n84740 , n84741 );
xnor ( n84743 , n84742 , n84433 );
and ( n84744 , n84127 , n84229 );
and ( n84745 , n84109 , n84227 );
nor ( n84746 , n84744 , n84745 );
xnor ( n84747 , n84746 , n84187 );
and ( n84748 , n84743 , n84747 );
and ( n84749 , n84655 , n83917 );
and ( n84750 , n84598 , n83915 );
nor ( n84751 , n84749 , n84750 );
xnor ( n84752 , n84751 , n83925 );
and ( n84753 , n84747 , n84752 );
and ( n84754 , n84743 , n84752 );
or ( n84755 , n84748 , n84753 , n84754 );
and ( n84756 , n84739 , n84755 );
and ( n84757 , n83909 , n84645 );
and ( n84758 , n83920 , n84642 );
nor ( n84759 , n84757 , n84758 );
xnor ( n84760 , n84759 , n84430 );
and ( n84761 , n84655 , n83915 );
not ( n84762 , n84761 );
and ( n84763 , n84762 , n83925 );
and ( n84764 , n84760 , n84763 );
and ( n84765 , n84755 , n84764 );
and ( n84766 , n84739 , n84764 );
or ( n84767 , n84756 , n84765 , n84766 );
xor ( n84768 , n84591 , n84595 );
xor ( n84769 , n84768 , n84599 );
and ( n84770 , n84767 , n84769 );
xor ( n84771 , n84606 , n84610 );
xor ( n84772 , n84771 , n84615 );
and ( n84773 , n84769 , n84772 );
and ( n84774 , n84767 , n84772 );
or ( n84775 , n84770 , n84773 , n84774 );
and ( n84776 , n84723 , n84775 );
xor ( n84777 , n84602 , n84618 );
xor ( n84778 , n84777 , n84621 );
and ( n84779 , n84775 , n84778 );
and ( n84780 , n84723 , n84778 );
or ( n84781 , n84776 , n84779 , n84780 );
xor ( n84782 , n84582 , n84584 );
xor ( n84783 , n84782 , n84587 );
and ( n84784 , n84781 , n84783 );
xor ( n84785 , n84624 , n84687 );
xor ( n84786 , n84785 , n84690 );
and ( n84787 , n84783 , n84786 );
and ( n84788 , n84781 , n84786 );
or ( n84789 , n84784 , n84787 , n84788 );
buf ( n84790 , n83881 );
and ( n84791 , n84789 , n84790 );
xor ( n84792 , n84590 , n84693 );
xor ( n84793 , n84792 , n84696 );
and ( n84794 , n84790 , n84793 );
and ( n84795 , n84789 , n84793 );
or ( n84796 , n84791 , n84794 , n84795 );
and ( n84797 , n84710 , n84796 );
xor ( n84798 , n84710 , n84796 );
xor ( n84799 , n84628 , n84632 );
xor ( n84800 , n84799 , n84637 );
xor ( n84801 , n84648 , n84652 );
xor ( n84802 , n84801 , n84656 );
and ( n84803 , n84800 , n84802 );
xor ( n84804 , n84664 , n84668 );
xor ( n84805 , n84804 , n84673 );
and ( n84806 , n84802 , n84805 );
and ( n84807 , n84800 , n84805 );
or ( n84808 , n84803 , n84806 , n84807 );
xor ( n84809 , n84640 , n84659 );
xor ( n84810 , n84809 , n84676 );
and ( n84811 , n84808 , n84810 );
xor ( n84812 , n84711 , n84715 );
xor ( n84813 , n84812 , n84720 );
and ( n84814 , n84810 , n84813 );
and ( n84815 , n84808 , n84813 );
or ( n84816 , n84811 , n84814 , n84815 );
xor ( n84817 , n84679 , n84681 );
xor ( n84818 , n84817 , n84684 );
and ( n84819 , n84816 , n84818 );
xor ( n84820 , n84723 , n84775 );
xor ( n84821 , n84820 , n84778 );
and ( n84822 , n84818 , n84821 );
and ( n84823 , n84816 , n84821 );
or ( n84824 , n84819 , n84822 , n84823 );
buf ( n84825 , n83882 );
and ( n84826 , n84824 , n84825 );
xor ( n84827 , n84781 , n84783 );
xor ( n84828 , n84827 , n84786 );
and ( n84829 , n84825 , n84828 );
and ( n84830 , n84824 , n84828 );
or ( n84831 , n84826 , n84829 , n84830 );
xor ( n84832 , n84789 , n84790 );
xor ( n84833 , n84832 , n84793 );
and ( n84834 , n84831 , n84833 );
xor ( n84835 , n84831 , n84833 );
xor ( n84836 , n84824 , n84825 );
xor ( n84837 , n84836 , n84828 );
xor ( n84838 , n84760 , n84763 );
and ( n84839 , n83929 , n84645 );
and ( n84840 , n83909 , n84642 );
nor ( n84841 , n84839 , n84840 );
xnor ( n84842 , n84841 , n84430 );
and ( n84843 , n83999 , n84455 );
and ( n84844 , n83957 , n84453 );
nor ( n84845 , n84843 , n84844 );
xnor ( n84846 , n84845 , n84433 );
and ( n84847 , n84842 , n84846 );
and ( n84848 , n84846 , n84761 );
and ( n84849 , n84842 , n84761 );
or ( n84850 , n84847 , n84848 , n84849 );
and ( n84851 , n84838 , n84850 );
and ( n84852 , n84515 , n83946 );
and ( n84853 , n84422 , n83944 );
nor ( n84854 , n84852 , n84853 );
xnor ( n84855 , n84854 , n83906 );
and ( n84856 , n84850 , n84855 );
and ( n84857 , n84838 , n84855 );
or ( n84858 , n84851 , n84856 , n84857 );
and ( n84859 , n84109 , n84354 );
and ( n84860 , n84014 , n84352 );
nor ( n84861 , n84859 , n84860 );
xnor ( n84862 , n84861 , n84299 );
and ( n84863 , n84167 , n84229 );
and ( n84864 , n84127 , n84227 );
nor ( n84865 , n84863 , n84864 );
xnor ( n84866 , n84865 , n84187 );
and ( n84867 , n84862 , n84866 );
and ( n84868 , n84361 , n84117 );
and ( n84869 , n84263 , n84115 );
nor ( n84870 , n84868 , n84869 );
xnor ( n84871 , n84870 , n84058 );
and ( n84872 , n84866 , n84871 );
and ( n84873 , n84862 , n84871 );
or ( n84874 , n84867 , n84872 , n84873 );
xor ( n84875 , n84727 , n84731 );
xor ( n84876 , n84875 , n84736 );
and ( n84877 , n84874 , n84876 );
xor ( n84878 , n84743 , n84747 );
xor ( n84879 , n84878 , n84752 );
and ( n84880 , n84876 , n84879 );
and ( n84881 , n84874 , n84879 );
or ( n84882 , n84877 , n84880 , n84881 );
and ( n84883 , n84858 , n84882 );
xor ( n84884 , n84739 , n84755 );
xor ( n84885 , n84884 , n84764 );
and ( n84886 , n84882 , n84885 );
and ( n84887 , n84858 , n84885 );
or ( n84888 , n84883 , n84886 , n84887 );
xor ( n84889 , n84767 , n84769 );
xor ( n84890 , n84889 , n84772 );
and ( n84891 , n84888 , n84890 );
xor ( n84892 , n84808 , n84810 );
xor ( n84893 , n84892 , n84813 );
and ( n84894 , n84890 , n84893 );
and ( n84895 , n84888 , n84893 );
or ( n84896 , n84891 , n84894 , n84895 );
buf ( n84897 , n83883 );
and ( n84898 , n84896 , n84897 );
xor ( n84899 , n84816 , n84818 );
xor ( n84900 , n84899 , n84821 );
and ( n84901 , n84897 , n84900 );
and ( n84902 , n84896 , n84900 );
or ( n84903 , n84898 , n84901 , n84902 );
and ( n84904 , n84837 , n84903 );
xor ( n84905 , n84837 , n84903 );
and ( n84906 , n83957 , n84645 );
and ( n84907 , n83929 , n84642 );
nor ( n84908 , n84906 , n84907 );
xnor ( n84909 , n84908 , n84430 );
and ( n84910 , n84655 , n83944 );
not ( n84911 , n84910 );
and ( n84912 , n84911 , n83906 );
and ( n84913 , n84909 , n84912 );
and ( n84914 , n84422 , n84022 );
and ( n84915 , n84376 , n84020 );
nor ( n84916 , n84914 , n84915 );
xnor ( n84917 , n84916 , n83991 );
and ( n84918 , n84913 , n84917 );
and ( n84919 , n84598 , n83946 );
and ( n84920 , n84515 , n83944 );
nor ( n84921 , n84919 , n84920 );
xnor ( n84922 , n84921 , n83906 );
and ( n84923 , n84917 , n84922 );
and ( n84924 , n84913 , n84922 );
or ( n84925 , n84918 , n84923 , n84924 );
and ( n84926 , n84014 , n84455 );
and ( n84927 , n83999 , n84453 );
nor ( n84928 , n84926 , n84927 );
xnor ( n84929 , n84928 , n84433 );
and ( n84930 , n84263 , n84229 );
and ( n84931 , n84167 , n84227 );
nor ( n84932 , n84930 , n84931 );
xnor ( n84933 , n84932 , n84187 );
and ( n84934 , n84929 , n84933 );
and ( n84935 , n84376 , n84117 );
and ( n84936 , n84361 , n84115 );
nor ( n84937 , n84935 , n84936 );
xnor ( n84938 , n84937 , n84058 );
and ( n84939 , n84933 , n84938 );
and ( n84940 , n84929 , n84938 );
or ( n84941 , n84934 , n84939 , n84940 );
and ( n84942 , n84127 , n84354 );
and ( n84943 , n84109 , n84352 );
nor ( n84944 , n84942 , n84943 );
xnor ( n84945 , n84944 , n84299 );
and ( n84946 , n84515 , n84022 );
and ( n84947 , n84422 , n84020 );
nor ( n84948 , n84946 , n84947 );
xnor ( n84949 , n84948 , n83991 );
and ( n84950 , n84945 , n84949 );
and ( n84951 , n84655 , n83946 );
and ( n84952 , n84598 , n83944 );
nor ( n84953 , n84951 , n84952 );
xnor ( n84954 , n84953 , n83906 );
and ( n84955 , n84949 , n84954 );
and ( n84956 , n84945 , n84954 );
or ( n84957 , n84950 , n84955 , n84956 );
and ( n84958 , n84941 , n84957 );
xor ( n84959 , n84842 , n84846 );
xor ( n84960 , n84959 , n84761 );
and ( n84961 , n84957 , n84960 );
and ( n84962 , n84941 , n84960 );
or ( n84963 , n84958 , n84961 , n84962 );
and ( n84964 , n84925 , n84963 );
xor ( n84965 , n84838 , n84850 );
xor ( n84966 , n84965 , n84855 );
and ( n84967 , n84963 , n84966 );
and ( n84968 , n84925 , n84966 );
or ( n84969 , n84964 , n84967 , n84968 );
xor ( n84970 , n84800 , n84802 );
xor ( n84971 , n84970 , n84805 );
and ( n84972 , n84969 , n84971 );
xor ( n84973 , n84858 , n84882 );
xor ( n84974 , n84973 , n84885 );
and ( n84975 , n84971 , n84974 );
and ( n84976 , n84969 , n84974 );
or ( n84977 , n84972 , n84975 , n84976 );
buf ( n84978 , n83884 );
and ( n84979 , n84977 , n84978 );
xor ( n84980 , n84888 , n84890 );
xor ( n84981 , n84980 , n84893 );
and ( n84982 , n84978 , n84981 );
and ( n84983 , n84977 , n84981 );
or ( n84984 , n84979 , n84982 , n84983 );
xor ( n84985 , n84896 , n84897 );
xor ( n84986 , n84985 , n84900 );
and ( n84987 , n84984 , n84986 );
xor ( n84988 , n84984 , n84986 );
xor ( n84989 , n84977 , n84978 );
xor ( n84990 , n84989 , n84981 );
xor ( n84991 , n84909 , n84912 );
and ( n84992 , n84109 , n84455 );
and ( n84993 , n84014 , n84453 );
nor ( n84994 , n84992 , n84993 );
xnor ( n84995 , n84994 , n84433 );
and ( n84996 , n84361 , n84229 );
and ( n84997 , n84263 , n84227 );
nor ( n84998 , n84996 , n84997 );
xnor ( n84999 , n84998 , n84187 );
and ( n85000 , n84995 , n84999 );
and ( n85001 , n84999 , n84910 );
and ( n85002 , n84995 , n84910 );
or ( n85003 , n85000 , n85001 , n85002 );
and ( n85004 , n84991 , n85003 );
and ( n85005 , n83999 , n84645 );
and ( n85006 , n83957 , n84642 );
nor ( n85007 , n85005 , n85006 );
xnor ( n85008 , n85007 , n84430 );
and ( n85009 , n84422 , n84117 );
and ( n85010 , n84376 , n84115 );
nor ( n85011 , n85009 , n85010 );
xnor ( n85012 , n85011 , n84058 );
and ( n85013 , n85008 , n85012 );
and ( n85014 , n84598 , n84022 );
and ( n85015 , n84515 , n84020 );
nor ( n85016 , n85014 , n85015 );
xnor ( n85017 , n85016 , n83991 );
and ( n85018 , n85012 , n85017 );
and ( n85019 , n85008 , n85017 );
or ( n85020 , n85013 , n85018 , n85019 );
and ( n85021 , n85003 , n85020 );
and ( n85022 , n84991 , n85020 );
or ( n85023 , n85004 , n85021 , n85022 );
xor ( n85024 , n84862 , n84866 );
xor ( n85025 , n85024 , n84871 );
and ( n85026 , n85023 , n85025 );
xor ( n85027 , n84913 , n84917 );
xor ( n85028 , n85027 , n84922 );
and ( n85029 , n85025 , n85028 );
and ( n85030 , n85023 , n85028 );
or ( n85031 , n85026 , n85029 , n85030 );
xor ( n85032 , n84874 , n84876 );
xor ( n85033 , n85032 , n84879 );
and ( n85034 , n85031 , n85033 );
xor ( n85035 , n84925 , n84963 );
xor ( n85036 , n85035 , n84966 );
and ( n85037 , n85033 , n85036 );
and ( n85038 , n85031 , n85036 );
or ( n85039 , n85034 , n85037 , n85038 );
buf ( n85040 , n83885 );
and ( n85041 , n85039 , n85040 );
xor ( n85042 , n84969 , n84971 );
xor ( n85043 , n85042 , n84974 );
and ( n85044 , n85040 , n85043 );
and ( n85045 , n85039 , n85043 );
or ( n85046 , n85041 , n85044 , n85045 );
and ( n85047 , n84990 , n85046 );
xor ( n85048 , n84990 , n85046 );
xor ( n85049 , n85039 , n85040 );
xor ( n85050 , n85049 , n85043 );
and ( n85051 , n84014 , n84645 );
and ( n85052 , n83999 , n84642 );
nor ( n85053 , n85051 , n85052 );
xnor ( n85054 , n85053 , n84430 );
and ( n85055 , n84376 , n84229 );
and ( n85056 , n84361 , n84227 );
nor ( n85057 , n85055 , n85056 );
xnor ( n85058 , n85057 , n84187 );
and ( n85059 , n85054 , n85058 );
and ( n85060 , n84515 , n84117 );
and ( n85061 , n84422 , n84115 );
nor ( n85062 , n85060 , n85061 );
xnor ( n85063 , n85062 , n84058 );
and ( n85064 , n85058 , n85063 );
and ( n85065 , n85054 , n85063 );
or ( n85066 , n85059 , n85064 , n85065 );
and ( n85067 , n84127 , n84455 );
and ( n85068 , n84109 , n84453 );
nor ( n85069 , n85067 , n85068 );
xnor ( n85070 , n85069 , n84433 );
and ( n85071 , n84655 , n84020 );
not ( n85072 , n85071 );
and ( n85073 , n85072 , n83991 );
and ( n85074 , n85070 , n85073 );
and ( n85075 , n85066 , n85074 );
and ( n85076 , n84167 , n84354 );
and ( n85077 , n84127 , n84352 );
nor ( n85078 , n85076 , n85077 );
xnor ( n85079 , n85078 , n84299 );
and ( n85080 , n85074 , n85079 );
and ( n85081 , n85066 , n85079 );
or ( n85082 , n85075 , n85080 , n85081 );
xor ( n85083 , n84929 , n84933 );
xor ( n85084 , n85083 , n84938 );
and ( n85085 , n85082 , n85084 );
xor ( n85086 , n84945 , n84949 );
xor ( n85087 , n85086 , n84954 );
and ( n85088 , n85084 , n85087 );
and ( n85089 , n85082 , n85087 );
or ( n85090 , n85085 , n85088 , n85089 );
xor ( n85091 , n84941 , n84957 );
xor ( n85092 , n85091 , n84960 );
and ( n85093 , n85090 , n85092 );
xor ( n85094 , n85023 , n85025 );
xor ( n85095 , n85094 , n85028 );
and ( n85096 , n85092 , n85095 );
and ( n85097 , n85090 , n85095 );
or ( n85098 , n85093 , n85096 , n85097 );
buf ( n85099 , n83886 );
and ( n85100 , n85098 , n85099 );
xor ( n85101 , n85031 , n85033 );
xor ( n85102 , n85101 , n85036 );
and ( n85103 , n85099 , n85102 );
and ( n85104 , n85098 , n85102 );
or ( n85105 , n85100 , n85103 , n85104 );
and ( n85106 , n85050 , n85105 );
xor ( n85107 , n85050 , n85105 );
xor ( n85108 , n85098 , n85099 );
xor ( n85109 , n85108 , n85102 );
xor ( n85110 , n85070 , n85073 );
and ( n85111 , n84263 , n84354 );
and ( n85112 , n84167 , n84352 );
nor ( n85113 , n85111 , n85112 );
xnor ( n85114 , n85113 , n84299 );
and ( n85115 , n85110 , n85114 );
and ( n85116 , n84655 , n84022 );
and ( n85117 , n84598 , n84020 );
nor ( n85118 , n85116 , n85117 );
xnor ( n85119 , n85118 , n83991 );
and ( n85120 , n85114 , n85119 );
and ( n85121 , n85110 , n85119 );
or ( n85122 , n85115 , n85120 , n85121 );
xor ( n85123 , n84995 , n84999 );
xor ( n85124 , n85123 , n84910 );
and ( n85125 , n85122 , n85124 );
xor ( n85126 , n85008 , n85012 );
xor ( n85127 , n85126 , n85017 );
and ( n85128 , n85124 , n85127 );
and ( n85129 , n85122 , n85127 );
or ( n85130 , n85125 , n85128 , n85129 );
xor ( n85131 , n84991 , n85003 );
xor ( n85132 , n85131 , n85020 );
and ( n85133 , n85130 , n85132 );
xor ( n85134 , n85082 , n85084 );
xor ( n85135 , n85134 , n85087 );
and ( n85136 , n85132 , n85135 );
and ( n85137 , n85130 , n85135 );
or ( n85138 , n85133 , n85136 , n85137 );
buf ( n85139 , n83887 );
and ( n85140 , n85138 , n85139 );
xor ( n85141 , n85090 , n85092 );
xor ( n85142 , n85141 , n85095 );
and ( n85143 , n85139 , n85142 );
and ( n85144 , n85138 , n85142 );
or ( n85145 , n85140 , n85143 , n85144 );
and ( n85146 , n85109 , n85145 );
xor ( n85147 , n85109 , n85145 );
xor ( n85148 , n85138 , n85139 );
xor ( n85149 , n85148 , n85142 );
and ( n85150 , n84109 , n84645 );
and ( n85151 , n84014 , n84642 );
nor ( n85152 , n85150 , n85151 );
xnor ( n85153 , n85152 , n84430 );
and ( n85154 , n84361 , n84354 );
and ( n85155 , n84263 , n84352 );
nor ( n85156 , n85154 , n85155 );
xnor ( n85157 , n85156 , n84299 );
and ( n85158 , n85153 , n85157 );
and ( n85159 , n84598 , n84117 );
and ( n85160 , n84515 , n84115 );
nor ( n85161 , n85159 , n85160 );
xnor ( n85162 , n85161 , n84058 );
and ( n85163 , n85157 , n85162 );
and ( n85164 , n85153 , n85162 );
or ( n85165 , n85158 , n85163 , n85164 );
and ( n85166 , n84167 , n84455 );
and ( n85167 , n84127 , n84453 );
nor ( n85168 , n85166 , n85167 );
xnor ( n85169 , n85168 , n84433 );
and ( n85170 , n84422 , n84229 );
and ( n85171 , n84376 , n84227 );
nor ( n85172 , n85170 , n85171 );
xnor ( n85173 , n85172 , n84187 );
and ( n85174 , n85169 , n85173 );
and ( n85175 , n85173 , n85071 );
and ( n85176 , n85169 , n85071 );
or ( n85177 , n85174 , n85175 , n85176 );
and ( n85178 , n85165 , n85177 );
xor ( n85179 , n85054 , n85058 );
xor ( n85180 , n85179 , n85063 );
and ( n85181 , n85177 , n85180 );
and ( n85182 , n85165 , n85180 );
or ( n85183 , n85178 , n85181 , n85182 );
xor ( n85184 , n85066 , n85074 );
xor ( n85185 , n85184 , n85079 );
and ( n85186 , n85183 , n85185 );
xor ( n85187 , n85122 , n85124 );
xor ( n85188 , n85187 , n85127 );
and ( n85189 , n85185 , n85188 );
and ( n85190 , n85183 , n85188 );
or ( n85191 , n85186 , n85189 , n85190 );
buf ( n85192 , n83888 );
and ( n85193 , n85191 , n85192 );
xor ( n85194 , n85130 , n85132 );
xor ( n85195 , n85194 , n85135 );
and ( n85196 , n85192 , n85195 );
and ( n85197 , n85191 , n85195 );
or ( n85198 , n85193 , n85196 , n85197 );
and ( n85199 , n85149 , n85198 );
xor ( n85200 , n85149 , n85198 );
xor ( n85201 , n85191 , n85192 );
xor ( n85202 , n85201 , n85195 );
and ( n85203 , n84127 , n84645 );
and ( n85204 , n84109 , n84642 );
nor ( n85205 , n85203 , n85204 );
xnor ( n85206 , n85205 , n84430 );
and ( n85207 , n84515 , n84229 );
and ( n85208 , n84422 , n84227 );
nor ( n85209 , n85207 , n85208 );
xnor ( n85210 , n85209 , n84187 );
and ( n85211 , n85206 , n85210 );
and ( n85212 , n84655 , n84117 );
and ( n85213 , n84598 , n84115 );
nor ( n85214 , n85212 , n85213 );
xnor ( n85215 , n85214 , n84058 );
and ( n85216 , n85210 , n85215 );
and ( n85217 , n85206 , n85215 );
or ( n85218 , n85211 , n85216 , n85217 );
and ( n85219 , n84263 , n84455 );
and ( n85220 , n84167 , n84453 );
nor ( n85221 , n85219 , n85220 );
xnor ( n85222 , n85221 , n84433 );
and ( n85223 , n84655 , n84115 );
not ( n85224 , n85223 );
and ( n85225 , n85224 , n84058 );
and ( n85226 , n85222 , n85225 );
and ( n85227 , n85218 , n85226 );
xor ( n85228 , n85169 , n85173 );
xor ( n85229 , n85228 , n85071 );
and ( n85230 , n85226 , n85229 );
and ( n85231 , n85218 , n85229 );
or ( n85232 , n85227 , n85230 , n85231 );
xor ( n85233 , n85110 , n85114 );
xor ( n85234 , n85233 , n85119 );
and ( n85235 , n85232 , n85234 );
xor ( n85236 , n85165 , n85177 );
xor ( n85237 , n85236 , n85180 );
and ( n85238 , n85234 , n85237 );
and ( n85239 , n85232 , n85237 );
or ( n85240 , n85235 , n85238 , n85239 );
buf ( n85241 , n83889 );
and ( n85242 , n85240 , n85241 );
xor ( n85243 , n85183 , n85185 );
xor ( n85244 , n85243 , n85188 );
and ( n85245 , n85241 , n85244 );
and ( n85246 , n85240 , n85244 );
or ( n85247 , n85242 , n85245 , n85246 );
and ( n85248 , n85202 , n85247 );
xor ( n85249 , n85202 , n85247 );
xor ( n85250 , n85222 , n85225 );
and ( n85251 , n84167 , n84645 );
and ( n85252 , n84127 , n84642 );
nor ( n85253 , n85251 , n85252 );
xnor ( n85254 , n85253 , n84430 );
and ( n85255 , n84598 , n84229 );
and ( n85256 , n84515 , n84227 );
nor ( n85257 , n85255 , n85256 );
xnor ( n85258 , n85257 , n84187 );
and ( n85259 , n85254 , n85258 );
and ( n85260 , n85258 , n85223 );
and ( n85261 , n85254 , n85223 );
or ( n85262 , n85259 , n85260 , n85261 );
and ( n85263 , n85250 , n85262 );
and ( n85264 , n84376 , n84354 );
and ( n85265 , n84361 , n84352 );
nor ( n85266 , n85264 , n85265 );
xnor ( n85267 , n85266 , n84299 );
and ( n85268 , n85262 , n85267 );
and ( n85269 , n85250 , n85267 );
or ( n85270 , n85263 , n85268 , n85269 );
xor ( n85271 , n85153 , n85157 );
xor ( n85272 , n85271 , n85162 );
and ( n85273 , n85270 , n85272 );
xor ( n85274 , n85218 , n85226 );
xor ( n85275 , n85274 , n85229 );
and ( n85276 , n85272 , n85275 );
and ( n85277 , n85270 , n85275 );
or ( n85278 , n85273 , n85276 , n85277 );
buf ( n85279 , n83890 );
and ( n85280 , n85278 , n85279 );
xor ( n85281 , n85232 , n85234 );
xor ( n85282 , n85281 , n85237 );
and ( n85283 , n85279 , n85282 );
and ( n85284 , n85278 , n85282 );
or ( n85285 , n85280 , n85283 , n85284 );
xor ( n85286 , n85240 , n85241 );
xor ( n85287 , n85286 , n85244 );
and ( n85288 , n85285 , n85287 );
xor ( n85289 , n85285 , n85287 );
xor ( n85290 , n85278 , n85279 );
xor ( n85291 , n85290 , n85282 );
and ( n85292 , n84263 , n84645 );
and ( n85293 , n84167 , n84642 );
nor ( n85294 , n85292 , n85293 );
xnor ( n85295 , n85294 , n84430 );
and ( n85296 , n84655 , n84227 );
not ( n85297 , n85296 );
and ( n85298 , n85297 , n84187 );
and ( n85299 , n85295 , n85298 );
and ( n85300 , n84361 , n84455 );
and ( n85301 , n84263 , n84453 );
nor ( n85302 , n85300 , n85301 );
xnor ( n85303 , n85302 , n84433 );
and ( n85304 , n85299 , n85303 );
and ( n85305 , n84422 , n84354 );
and ( n85306 , n84376 , n84352 );
nor ( n85307 , n85305 , n85306 );
xnor ( n85308 , n85307 , n84299 );
and ( n85309 , n85303 , n85308 );
and ( n85310 , n85299 , n85308 );
or ( n85311 , n85304 , n85309 , n85310 );
xor ( n85312 , n85206 , n85210 );
xor ( n85313 , n85312 , n85215 );
and ( n85314 , n85311 , n85313 );
xor ( n85315 , n85250 , n85262 );
xor ( n85316 , n85315 , n85267 );
and ( n85317 , n85313 , n85316 );
and ( n85318 , n85311 , n85316 );
or ( n85319 , n85314 , n85317 , n85318 );
buf ( n85320 , n83891 );
and ( n85321 , n85319 , n85320 );
xor ( n85322 , n85270 , n85272 );
xor ( n85323 , n85322 , n85275 );
and ( n85324 , n85320 , n85323 );
and ( n85325 , n85319 , n85323 );
or ( n85326 , n85321 , n85324 , n85325 );
and ( n85327 , n85291 , n85326 );
xor ( n85328 , n85291 , n85326 );
xor ( n85329 , n85319 , n85320 );
xor ( n85330 , n85329 , n85323 );
and ( n85331 , n84376 , n84455 );
and ( n85332 , n84361 , n84453 );
nor ( n85333 , n85331 , n85332 );
xnor ( n85334 , n85333 , n84433 );
and ( n85335 , n84515 , n84354 );
and ( n85336 , n84422 , n84352 );
nor ( n85337 , n85335 , n85336 );
xnor ( n85338 , n85337 , n84299 );
and ( n85339 , n85334 , n85338 );
and ( n85340 , n84655 , n84229 );
and ( n85341 , n84598 , n84227 );
nor ( n85342 , n85340 , n85341 );
xnor ( n85343 , n85342 , n84187 );
and ( n85344 , n85338 , n85343 );
and ( n85345 , n85334 , n85343 );
or ( n85346 , n85339 , n85344 , n85345 );
xor ( n85347 , n85254 , n85258 );
xor ( n85348 , n85347 , n85223 );
and ( n85349 , n85346 , n85348 );
xor ( n85350 , n85299 , n85303 );
xor ( n85351 , n85350 , n85308 );
and ( n85352 , n85348 , n85351 );
and ( n85353 , n85346 , n85351 );
or ( n85354 , n85349 , n85352 , n85353 );
buf ( n85355 , n83892 );
and ( n85356 , n85354 , n85355 );
xor ( n85357 , n85311 , n85313 );
xor ( n85358 , n85357 , n85316 );
and ( n85359 , n85355 , n85358 );
and ( n85360 , n85354 , n85358 );
or ( n85361 , n85356 , n85359 , n85360 );
and ( n85362 , n85330 , n85361 );
xor ( n85363 , n85330 , n85361 );
xor ( n85364 , n85354 , n85355 );
xor ( n85365 , n85364 , n85358 );
xor ( n85366 , n85295 , n85298 );
and ( n85367 , n84361 , n84645 );
and ( n85368 , n84263 , n84642 );
nor ( n85369 , n85367 , n85368 );
xnor ( n85370 , n85369 , n84430 );
and ( n85371 , n84422 , n84455 );
and ( n85372 , n84376 , n84453 );
nor ( n85373 , n85371 , n85372 );
xnor ( n85374 , n85373 , n84433 );
and ( n85375 , n85370 , n85374 );
and ( n85376 , n85374 , n85296 );
and ( n85377 , n85370 , n85296 );
or ( n85378 , n85375 , n85376 , n85377 );
and ( n85379 , n85366 , n85378 );
xor ( n85380 , n85334 , n85338 );
xor ( n85381 , n85380 , n85343 );
and ( n85382 , n85378 , n85381 );
and ( n85383 , n85366 , n85381 );
or ( n85384 , n85379 , n85382 , n85383 );
buf ( n85385 , n83893 );
and ( n85386 , n85384 , n85385 );
xor ( n85387 , n85346 , n85348 );
xor ( n85388 , n85387 , n85351 );
and ( n85389 , n85385 , n85388 );
and ( n85390 , n85384 , n85388 );
or ( n85391 , n85386 , n85389 , n85390 );
and ( n85392 , n85365 , n85391 );
xor ( n85393 , n85365 , n85391 );
and ( n85394 , n84376 , n84645 );
and ( n85395 , n84361 , n84642 );
nor ( n85396 , n85394 , n85395 );
xnor ( n85397 , n85396 , n84430 );
and ( n85398 , n84655 , n84352 );
not ( n85399 , n85398 );
and ( n85400 , n85399 , n84299 );
and ( n85401 , n85397 , n85400 );
and ( n85402 , n84598 , n84354 );
and ( n85403 , n84515 , n84352 );
nor ( n85404 , n85402 , n85403 );
xnor ( n85405 , n85404 , n84299 );
and ( n85406 , n85401 , n85405 );
xor ( n85407 , n85370 , n85374 );
xor ( n85408 , n85407 , n85296 );
and ( n85409 , n85405 , n85408 );
and ( n85410 , n85401 , n85408 );
or ( n85411 , n85406 , n85409 , n85410 );
buf ( n85412 , n83894 );
and ( n85413 , n85411 , n85412 );
xor ( n85414 , n85366 , n85378 );
xor ( n85415 , n85414 , n85381 );
and ( n85416 , n85412 , n85415 );
and ( n85417 , n85411 , n85415 );
or ( n85418 , n85413 , n85416 , n85417 );
xor ( n85419 , n85384 , n85385 );
xor ( n85420 , n85419 , n85388 );
and ( n85421 , n85418 , n85420 );
xor ( n85422 , n85418 , n85420 );
xor ( n85423 , n85411 , n85412 );
xor ( n85424 , n85423 , n85415 );
xor ( n85425 , n85397 , n85400 );
and ( n85426 , n84515 , n84455 );
and ( n85427 , n84422 , n84453 );
nor ( n85428 , n85426 , n85427 );
xnor ( n85429 , n85428 , n84433 );
and ( n85430 , n85425 , n85429 );
and ( n85431 , n84655 , n84354 );
and ( n85432 , n84598 , n84352 );
nor ( n85433 , n85431 , n85432 );
xnor ( n85434 , n85433 , n84299 );
and ( n85435 , n85429 , n85434 );
and ( n85436 , n85425 , n85434 );
or ( n85437 , n85430 , n85435 , n85436 );
buf ( n85438 , n83895 );
and ( n85439 , n85437 , n85438 );
xor ( n85440 , n85401 , n85405 );
xor ( n85441 , n85440 , n85408 );
and ( n85442 , n85438 , n85441 );
and ( n85443 , n85437 , n85441 );
or ( n85444 , n85439 , n85442 , n85443 );
and ( n85445 , n85424 , n85444 );
xor ( n85446 , n85424 , n85444 );
xor ( n85447 , n85437 , n85438 );
xor ( n85448 , n85447 , n85441 );
and ( n85449 , n84422 , n84645 );
and ( n85450 , n84376 , n84642 );
nor ( n85451 , n85449 , n85450 );
xnor ( n85452 , n85451 , n84430 );
and ( n85453 , n84598 , n84455 );
and ( n85454 , n84515 , n84453 );
nor ( n85455 , n85453 , n85454 );
xnor ( n85456 , n85455 , n84433 );
and ( n85457 , n85452 , n85456 );
and ( n85458 , n85456 , n85398 );
and ( n85459 , n85452 , n85398 );
or ( n85460 , n85457 , n85458 , n85459 );
buf ( n85461 , n83896 );
and ( n85462 , n85460 , n85461 );
xor ( n85463 , n85425 , n85429 );
xor ( n85464 , n85463 , n85434 );
and ( n85465 , n85461 , n85464 );
and ( n85466 , n85460 , n85464 );
or ( n85467 , n85462 , n85465 , n85466 );
and ( n85468 , n85448 , n85467 );
xor ( n85469 , n85448 , n85467 );
and ( n85470 , n84515 , n84645 );
and ( n85471 , n84422 , n84642 );
nor ( n85472 , n85470 , n85471 );
xnor ( n85473 , n85472 , n84430 );
and ( n85474 , n84655 , n84453 );
not ( n85475 , n85474 );
and ( n85476 , n85475 , n84433 );
and ( n85477 , n85473 , n85476 );
buf ( n85478 , n83897 );
and ( n85479 , n85477 , n85478 );
xor ( n85480 , n85452 , n85456 );
xor ( n85481 , n85480 , n85398 );
and ( n85482 , n85478 , n85481 );
and ( n85483 , n85477 , n85481 );
or ( n85484 , n85479 , n85482 , n85483 );
xor ( n85485 , n85460 , n85461 );
xor ( n85486 , n85485 , n85464 );
and ( n85487 , n85484 , n85486 );
xor ( n85488 , n85484 , n85486 );
xor ( n85489 , n85477 , n85478 );
xor ( n85490 , n85489 , n85481 );
and ( n85491 , n84655 , n84455 );
and ( n85492 , n84598 , n84453 );
nor ( n85493 , n85491 , n85492 );
xnor ( n85494 , n85493 , n84433 );
xor ( n85495 , n85473 , n85476 );
and ( n85496 , n85494 , n85495 );
and ( n85497 , n85490 , n85496 );
xor ( n85498 , n85490 , n85496 );
and ( n85499 , n84598 , n84645 );
and ( n85500 , n84515 , n84642 );
nor ( n85501 , n85499 , n85500 );
xnor ( n85502 , n85501 , n84430 );
or ( n85503 , n85502 , n85474 );
xor ( n85504 , n85494 , n85495 );
and ( n85505 , n85503 , n85504 );
xor ( n85506 , n85503 , n85504 );
and ( n85507 , n84655 , n84645 );
and ( n85508 , n84598 , n84642 );
nor ( n85509 , n85507 , n85508 );
xnor ( n85510 , n85509 , n84430 );
and ( n85511 , n84655 , n84642 );
not ( n85512 , n85511 );
and ( n85513 , n85512 , n84430 );
and ( n85514 , n85510 , n85513 );
xnor ( n85515 , n85502 , n85474 );
and ( n85516 , n85514 , n85515 );
xor ( n85517 , n85514 , n85515 );
xor ( n85518 , n85510 , n85513 );
and ( n85519 , n85518 , n85511 );
and ( n85520 , n85517 , n85519 );
or ( n85521 , n85516 , n85520 );
and ( n85522 , n85506 , n85521 );
or ( n85523 , n85505 , n85522 );
and ( n85524 , n85498 , n85523 );
or ( n85525 , n85497 , n85524 );
and ( n85526 , n85488 , n85525 );
or ( n85527 , n85487 , n85526 );
and ( n85528 , n85469 , n85527 );
or ( n85529 , n85468 , n85528 );
and ( n85530 , n85446 , n85529 );
or ( n85531 , n85445 , n85530 );
and ( n85532 , n85422 , n85531 );
or ( n85533 , n85421 , n85532 );
and ( n85534 , n85393 , n85533 );
or ( n85535 , n85392 , n85534 );
and ( n85536 , n85363 , n85535 );
or ( n85537 , n85362 , n85536 );
and ( n85538 , n85328 , n85537 );
or ( n85539 , n85327 , n85538 );
and ( n85540 , n85289 , n85539 );
or ( n85541 , n85288 , n85540 );
and ( n85542 , n85249 , n85541 );
or ( n85543 , n85248 , n85542 );
and ( n85544 , n85200 , n85543 );
or ( n85545 , n85199 , n85544 );
and ( n85546 , n85147 , n85545 );
or ( n85547 , n85146 , n85546 );
and ( n85548 , n85107 , n85547 );
or ( n85549 , n85106 , n85548 );
and ( n85550 , n85048 , n85549 );
or ( n85551 , n85047 , n85550 );
and ( n85552 , n84988 , n85551 );
or ( n85553 , n84987 , n85552 );
and ( n85554 , n84905 , n85553 );
or ( n85555 , n84904 , n85554 );
and ( n85556 , n84835 , n85555 );
or ( n85557 , n84834 , n85556 );
and ( n85558 , n84798 , n85557 );
or ( n85559 , n84797 , n85558 );
and ( n85560 , n84708 , n85559 );
or ( n85561 , n84707 , n85560 );
and ( n85562 , n84566 , n85561 );
or ( n85563 , n84565 , n85562 );
and ( n85564 , n84502 , n85563 );
or ( n85565 , n84501 , n85564 );
and ( n85566 , n84409 , n85565 );
or ( n85567 , n84408 , n85566 );
and ( n85568 , n84290 , n85567 );
or ( n85569 , n84289 , n85568 );
and ( n85570 , n84223 , n85569 );
or ( n85571 , n84222 , n85570 );
and ( n85572 , n84154 , n85571 );
or ( n85573 , n84153 , n85572 );
and ( n85574 , n84095 , n85573 );
or ( n85575 , n84094 , n85574 );
and ( n85576 , n84049 , n85575 );
or ( n85577 , n84048 , n85576 );
xor ( n85578 , n83982 , n85577 );
buf ( n85579 , n85578 );
xor ( n85580 , n84049 , n85575 );
buf ( n85581 , n85580 );
xor ( n85582 , n84095 , n85573 );
buf ( n85583 , n85582 );
xor ( n85584 , n84154 , n85571 );
buf ( n85585 , n85584 );
xor ( n85586 , n84223 , n85569 );
buf ( n85587 , n85586 );
xor ( n85588 , n84290 , n85567 );
buf ( n85589 , n85588 );
xor ( n85590 , n84409 , n85565 );
buf ( n85591 , n85590 );
xor ( n85592 , n84502 , n85563 );
buf ( n85593 , n85592 );
xor ( n85594 , n84566 , n85561 );
buf ( n85595 , n85594 );
xor ( n85596 , n84708 , n85559 );
buf ( n85597 , n85596 );
xor ( n85598 , n84798 , n85557 );
buf ( n85599 , n85598 );
xor ( n85600 , n84835 , n85555 );
buf ( n85601 , n85600 );
xor ( n85602 , n84905 , n85553 );
buf ( n85603 , n85602 );
xor ( n85604 , n84988 , n85551 );
buf ( n85605 , n85604 );
xor ( n85606 , n85048 , n85549 );
buf ( n85607 , n85606 );
xor ( n85608 , n85107 , n85547 );
buf ( n85609 , n85608 );
xor ( n85610 , n85147 , n85545 );
buf ( n85611 , n85610 );
xor ( n85612 , n85200 , n85543 );
buf ( n85613 , n85612 );
xor ( n85614 , n85249 , n85541 );
buf ( n85615 , n85614 );
xor ( n85616 , n85289 , n85539 );
buf ( n85617 , n85616 );
xor ( n85618 , n85328 , n85537 );
buf ( n85619 , n85618 );
xor ( n85620 , n85363 , n85535 );
buf ( n85621 , n85620 );
xor ( n85622 , n85393 , n85533 );
buf ( n85623 , n85622 );
xor ( n85624 , n85422 , n85531 );
buf ( n85625 , n85624 );
xor ( n85626 , n85446 , n85529 );
buf ( n85627 , n85626 );
xor ( n85628 , n85469 , n85527 );
buf ( n85629 , n85628 );
xor ( n85630 , n85488 , n85525 );
buf ( n85631 , n85630 );
xor ( n85632 , n85498 , n85523 );
buf ( n85633 , n85632 );
xor ( n85634 , n85506 , n85521 );
buf ( n85635 , n85634 );
xor ( n85636 , n85517 , n85519 );
buf ( n85637 , n85636 );
xor ( n85638 , n85518 , n85511 );
buf ( n85639 , n85638 );
buf ( n85640 , n85512 );
buf ( n85641 , n85640 );
buf ( n85642 , n29719 );
buf ( n85643 , n29721 );
buf ( n85644 , n29723 );
buf ( n85645 , n29725 );
buf ( n85646 , n29727 );
buf ( n85647 , n29729 );
buf ( n85648 , n29731 );
buf ( n85649 , n29733 );
buf ( n85650 , n29735 );
buf ( n85651 , n29737 );
buf ( n85652 , n29739 );
buf ( n85653 , n29741 );
buf ( n85654 , n29743 );
buf ( n85655 , n29745 );
buf ( n85656 , n29747 );
buf ( n85657 , n29749 );
buf ( n85658 , n29751 );
buf ( n85659 , n29753 );
buf ( n85660 , n29755 );
buf ( n85661 , n29757 );
buf ( n85662 , n29759 );
buf ( n85663 , n29761 );
buf ( n85664 , n29763 );
buf ( n85665 , n29765 );
buf ( n85666 , n29767 );
buf ( n85667 , n29769 );
buf ( n85668 , n29771 );
buf ( n85669 , n544 );
buf ( n85670 , n85669 );
buf ( n85671 , n562 );
buf ( n85672 , n85671 );
buf ( n85673 , n563 );
buf ( n85674 , n85673 );
xor ( n85675 , n85672 , n85674 );
buf ( n85676 , n564 );
buf ( n85677 , n85676 );
xor ( n85678 , n85674 , n85677 );
not ( n85679 , n85678 );
and ( n85680 , n85675 , n85679 );
and ( n85681 , n85670 , n85680 );
not ( n85682 , n85681 );
and ( n85683 , n85674 , n85677 );
not ( n85684 , n85683 );
and ( n85685 , n85672 , n85684 );
xnor ( n85686 , n85682 , n85685 );
not ( n85687 , n85686 );
buf ( n85688 , n546 );
buf ( n85689 , n85688 );
buf ( n85690 , n560 );
buf ( n85691 , n85690 );
buf ( n85692 , n561 );
buf ( n85693 , n85692 );
xor ( n85694 , n85691 , n85693 );
xor ( n85695 , n85693 , n85672 );
not ( n85696 , n85695 );
and ( n85697 , n85694 , n85696 );
and ( n85698 , n85689 , n85697 );
buf ( n85699 , n545 );
buf ( n85700 , n85699 );
and ( n85701 , n85700 , n85695 );
nor ( n85702 , n85698 , n85701 );
and ( n85703 , n85693 , n85672 );
not ( n85704 , n85703 );
and ( n85705 , n85691 , n85704 );
xnor ( n85706 , n85702 , n85705 );
and ( n85707 , n85687 , n85706 );
buf ( n85708 , n547 );
buf ( n85709 , n85708 );
and ( n85710 , n85709 , n85691 );
and ( n85711 , n85706 , n85710 );
and ( n85712 , n85687 , n85710 );
or ( n85713 , n85707 , n85711 , n85712 );
buf ( n85714 , n85686 );
and ( n85715 , n85713 , n85714 );
not ( n85716 , n85685 );
and ( n85717 , n85700 , n85697 );
and ( n85718 , n85670 , n85695 );
nor ( n85719 , n85717 , n85718 );
xnor ( n85720 , n85719 , n85705 );
xor ( n85721 , n85716 , n85720 );
and ( n85722 , n85689 , n85691 );
xor ( n85723 , n85721 , n85722 );
and ( n85724 , n85714 , n85723 );
and ( n85725 , n85713 , n85723 );
or ( n85726 , n85715 , n85724 , n85725 );
and ( n85727 , n85716 , n85720 );
and ( n85728 , n85720 , n85722 );
and ( n85729 , n85716 , n85722 );
or ( n85730 , n85727 , n85728 , n85729 );
and ( n85731 , n85670 , n85697 );
not ( n85732 , n85731 );
xnor ( n85733 , n85732 , n85705 );
xor ( n85734 , n85730 , n85733 );
and ( n85735 , n85700 , n85691 );
not ( n85736 , n85735 );
xor ( n85737 , n85734 , n85736 );
and ( n85738 , n85726 , n85737 );
and ( n85739 , n85730 , n85733 );
and ( n85740 , n85733 , n85736 );
and ( n85741 , n85730 , n85736 );
or ( n85742 , n85739 , n85740 , n85741 );
buf ( n85743 , n85735 );
not ( n85744 , n85705 );
xor ( n85745 , n85743 , n85744 );
and ( n85746 , n85670 , n85691 );
xor ( n85747 , n85745 , n85746 );
xor ( n85748 , n85742 , n85747 );
xor ( n85749 , n85738 , n85748 );
buf ( n85750 , n85642 );
xor ( n85751 , n85726 , n85737 );
and ( n85752 , n85750 , n85751 );
buf ( n85753 , n565 );
buf ( n85754 , n85753 );
buf ( n85755 , n566 );
buf ( n85756 , n85755 );
and ( n85757 , n85754 , n85756 );
not ( n85758 , n85757 );
and ( n85759 , n85677 , n85758 );
not ( n85760 , n85759 );
and ( n85761 , n85700 , n85680 );
and ( n85762 , n85670 , n85678 );
nor ( n85763 , n85761 , n85762 );
xnor ( n85764 , n85763 , n85685 );
and ( n85765 , n85760 , n85764 );
buf ( n85766 , n548 );
buf ( n85767 , n85766 );
and ( n85768 , n85767 , n85691 );
and ( n85769 , n85764 , n85768 );
and ( n85770 , n85760 , n85768 );
or ( n85771 , n85765 , n85769 , n85770 );
and ( n85772 , n85689 , n85680 );
and ( n85773 , n85700 , n85678 );
nor ( n85774 , n85772 , n85773 );
xnor ( n85775 , n85774 , n85685 );
and ( n85776 , n85767 , n85697 );
and ( n85777 , n85709 , n85695 );
nor ( n85778 , n85776 , n85777 );
xnor ( n85779 , n85778 , n85705 );
and ( n85780 , n85775 , n85779 );
buf ( n85781 , n549 );
buf ( n85782 , n85781 );
and ( n85783 , n85782 , n85691 );
and ( n85784 , n85779 , n85783 );
and ( n85785 , n85775 , n85783 );
or ( n85786 , n85780 , n85784 , n85785 );
xor ( n85787 , n85677 , n85754 );
xor ( n85788 , n85754 , n85756 );
not ( n85789 , n85788 );
and ( n85790 , n85787 , n85789 );
and ( n85791 , n85670 , n85790 );
not ( n85792 , n85791 );
xnor ( n85793 , n85792 , n85759 );
buf ( n85794 , n85793 );
and ( n85795 , n85786 , n85794 );
and ( n85796 , n85709 , n85697 );
and ( n85797 , n85689 , n85695 );
nor ( n85798 , n85796 , n85797 );
xnor ( n85799 , n85798 , n85705 );
and ( n85800 , n85794 , n85799 );
and ( n85801 , n85786 , n85799 );
or ( n85802 , n85795 , n85800 , n85801 );
and ( n85803 , n85771 , n85802 );
xor ( n85804 , n85687 , n85706 );
xor ( n85805 , n85804 , n85710 );
and ( n85806 , n85802 , n85805 );
and ( n85807 , n85771 , n85805 );
or ( n85808 , n85803 , n85806 , n85807 );
xor ( n85809 , n85713 , n85714 );
xor ( n85810 , n85809 , n85723 );
and ( n85811 , n85808 , n85810 );
and ( n85812 , n85751 , n85811 );
and ( n85813 , n85750 , n85811 );
or ( n85814 , n85752 , n85812 , n85813 );
xor ( n85815 , n85749 , n85814 );
buf ( n85816 , n85643 );
xor ( n85817 , n85808 , n85810 );
and ( n85818 , n85816 , n85817 );
buf ( n85819 , n567 );
buf ( n85820 , n85819 );
buf ( n85821 , n568 );
buf ( n85822 , n85821 );
and ( n85823 , n85820 , n85822 );
not ( n85824 , n85823 );
and ( n85825 , n85756 , n85824 );
not ( n85826 , n85825 );
and ( n85827 , n85700 , n85790 );
and ( n85828 , n85670 , n85788 );
nor ( n85829 , n85827 , n85828 );
xnor ( n85830 , n85829 , n85759 );
and ( n85831 , n85826 , n85830 );
and ( n85832 , n85782 , n85697 );
and ( n85833 , n85767 , n85695 );
nor ( n85834 , n85832 , n85833 );
xnor ( n85835 , n85834 , n85705 );
and ( n85836 , n85830 , n85835 );
and ( n85837 , n85826 , n85835 );
or ( n85838 , n85831 , n85836 , n85837 );
not ( n85839 , n85793 );
and ( n85840 , n85838 , n85839 );
xor ( n85841 , n85775 , n85779 );
xor ( n85842 , n85841 , n85783 );
and ( n85843 , n85839 , n85842 );
and ( n85844 , n85838 , n85842 );
or ( n85845 , n85840 , n85843 , n85844 );
xor ( n85846 , n85760 , n85764 );
xor ( n85847 , n85846 , n85768 );
and ( n85848 , n85845 , n85847 );
xor ( n85849 , n85786 , n85794 );
xor ( n85850 , n85849 , n85799 );
and ( n85851 , n85847 , n85850 );
and ( n85852 , n85845 , n85850 );
or ( n85853 , n85848 , n85851 , n85852 );
xor ( n85854 , n85771 , n85802 );
xor ( n85855 , n85854 , n85805 );
and ( n85856 , n85853 , n85855 );
and ( n85857 , n85817 , n85856 );
and ( n85858 , n85816 , n85856 );
or ( n85859 , n85818 , n85857 , n85858 );
xor ( n85860 , n85750 , n85751 );
xor ( n85861 , n85860 , n85811 );
and ( n85862 , n85859 , n85861 );
xor ( n85863 , n85816 , n85817 );
xor ( n85864 , n85863 , n85856 );
buf ( n85865 , n85644 );
xor ( n85866 , n85853 , n85855 );
and ( n85867 , n85865 , n85866 );
and ( n85868 , n85689 , n85790 );
and ( n85869 , n85700 , n85788 );
nor ( n85870 , n85868 , n85869 );
xnor ( n85871 , n85870 , n85759 );
buf ( n85872 , n85871 );
and ( n85873 , n85709 , n85680 );
and ( n85874 , n85689 , n85678 );
nor ( n85875 , n85873 , n85874 );
xnor ( n85876 , n85875 , n85685 );
and ( n85877 , n85872 , n85876 );
buf ( n85878 , n550 );
buf ( n85879 , n85878 );
and ( n85880 , n85879 , n85691 );
and ( n85881 , n85876 , n85880 );
and ( n85882 , n85872 , n85880 );
or ( n85883 , n85877 , n85881 , n85882 );
xor ( n85884 , n85756 , n85820 );
xor ( n85885 , n85820 , n85822 );
not ( n85886 , n85885 );
and ( n85887 , n85884 , n85886 );
and ( n85888 , n85670 , n85887 );
not ( n85889 , n85888 );
xnor ( n85890 , n85889 , n85825 );
and ( n85891 , n85879 , n85697 );
and ( n85892 , n85782 , n85695 );
nor ( n85893 , n85891 , n85892 );
xnor ( n85894 , n85893 , n85705 );
and ( n85895 , n85890 , n85894 );
buf ( n85896 , n551 );
buf ( n85897 , n85896 );
and ( n85898 , n85897 , n85691 );
and ( n85899 , n85894 , n85898 );
and ( n85900 , n85890 , n85898 );
or ( n85901 , n85895 , n85899 , n85900 );
xor ( n85902 , n85826 , n85830 );
xor ( n85903 , n85902 , n85835 );
and ( n85904 , n85901 , n85903 );
xor ( n85905 , n85872 , n85876 );
xor ( n85906 , n85905 , n85880 );
and ( n85907 , n85903 , n85906 );
and ( n85908 , n85901 , n85906 );
or ( n85909 , n85904 , n85907 , n85908 );
and ( n85910 , n85883 , n85909 );
xor ( n85911 , n85838 , n85839 );
xor ( n85912 , n85911 , n85842 );
and ( n85913 , n85909 , n85912 );
and ( n85914 , n85883 , n85912 );
or ( n85915 , n85910 , n85913 , n85914 );
xor ( n85916 , n85845 , n85847 );
xor ( n85917 , n85916 , n85850 );
and ( n85918 , n85915 , n85917 );
and ( n85919 , n85866 , n85918 );
and ( n85920 , n85865 , n85918 );
or ( n85921 , n85867 , n85919 , n85920 );
and ( n85922 , n85864 , n85921 );
buf ( n85923 , n85645 );
xor ( n85924 , n85915 , n85917 );
and ( n85925 , n85923 , n85924 );
and ( n85926 , n85709 , n85790 );
and ( n85927 , n85689 , n85788 );
nor ( n85928 , n85926 , n85927 );
xnor ( n85929 , n85928 , n85759 );
and ( n85930 , n85897 , n85697 );
and ( n85931 , n85879 , n85695 );
nor ( n85932 , n85930 , n85931 );
xnor ( n85933 , n85932 , n85705 );
and ( n85934 , n85929 , n85933 );
buf ( n85935 , n552 );
buf ( n85936 , n85935 );
and ( n85937 , n85936 , n85691 );
and ( n85938 , n85933 , n85937 );
and ( n85939 , n85929 , n85937 );
or ( n85940 , n85934 , n85938 , n85939 );
not ( n85941 , n85871 );
and ( n85942 , n85940 , n85941 );
and ( n85943 , n85767 , n85680 );
and ( n85944 , n85709 , n85678 );
nor ( n85945 , n85943 , n85944 );
xnor ( n85946 , n85945 , n85685 );
and ( n85947 , n85941 , n85946 );
and ( n85948 , n85940 , n85946 );
or ( n85949 , n85942 , n85947 , n85948 );
buf ( n85950 , n569 );
buf ( n85951 , n85950 );
buf ( n85952 , n570 );
buf ( n85953 , n85952 );
and ( n85954 , n85951 , n85953 );
not ( n85955 , n85954 );
and ( n85956 , n85822 , n85955 );
not ( n85957 , n85956 );
and ( n85958 , n85700 , n85887 );
and ( n85959 , n85670 , n85885 );
nor ( n85960 , n85958 , n85959 );
xnor ( n85961 , n85960 , n85825 );
and ( n85962 , n85957 , n85961 );
and ( n85963 , n85782 , n85680 );
and ( n85964 , n85767 , n85678 );
nor ( n85965 , n85963 , n85964 );
xnor ( n85966 , n85965 , n85685 );
and ( n85967 , n85961 , n85966 );
and ( n85968 , n85957 , n85966 );
or ( n85969 , n85962 , n85967 , n85968 );
xor ( n85970 , n85890 , n85894 );
xor ( n85971 , n85970 , n85898 );
and ( n85972 , n85969 , n85971 );
xor ( n85973 , n85940 , n85941 );
xor ( n85974 , n85973 , n85946 );
and ( n85975 , n85971 , n85974 );
and ( n85976 , n85969 , n85974 );
or ( n85977 , n85972 , n85975 , n85976 );
and ( n85978 , n85949 , n85977 );
xor ( n85979 , n85901 , n85903 );
xor ( n85980 , n85979 , n85906 );
and ( n85981 , n85977 , n85980 );
and ( n85982 , n85949 , n85980 );
or ( n85983 , n85978 , n85981 , n85982 );
xor ( n85984 , n85883 , n85909 );
xor ( n85985 , n85984 , n85912 );
and ( n85986 , n85983 , n85985 );
and ( n85987 , n85924 , n85986 );
and ( n85988 , n85923 , n85986 );
or ( n85989 , n85925 , n85987 , n85988 );
xor ( n85990 , n85865 , n85866 );
xor ( n85991 , n85990 , n85918 );
and ( n85992 , n85989 , n85991 );
buf ( n85993 , n85646 );
xor ( n85994 , n85983 , n85985 );
and ( n85995 , n85993 , n85994 );
xor ( n85996 , n85822 , n85951 );
xor ( n85997 , n85951 , n85953 );
not ( n85998 , n85997 );
and ( n85999 , n85996 , n85998 );
and ( n86000 , n85670 , n85999 );
not ( n86001 , n86000 );
xnor ( n86002 , n86001 , n85956 );
and ( n86003 , n85879 , n85680 );
and ( n86004 , n85782 , n85678 );
nor ( n86005 , n86003 , n86004 );
xnor ( n86006 , n86005 , n85685 );
and ( n86007 , n86002 , n86006 );
and ( n86008 , n85936 , n85697 );
and ( n86009 , n85897 , n85695 );
nor ( n86010 , n86008 , n86009 );
xnor ( n86011 , n86010 , n85705 );
and ( n86012 , n86006 , n86011 );
and ( n86013 , n86002 , n86011 );
or ( n86014 , n86007 , n86012 , n86013 );
and ( n86015 , n85689 , n85887 );
and ( n86016 , n85700 , n85885 );
nor ( n86017 , n86015 , n86016 );
xnor ( n86018 , n86017 , n85825 );
buf ( n86019 , n86018 );
and ( n86020 , n86014 , n86019 );
xor ( n86021 , n85929 , n85933 );
xor ( n86022 , n86021 , n85937 );
and ( n86023 , n86019 , n86022 );
and ( n86024 , n86014 , n86022 );
or ( n86025 , n86020 , n86023 , n86024 );
not ( n86026 , n86018 );
and ( n86027 , n85767 , n85790 );
and ( n86028 , n85709 , n85788 );
nor ( n86029 , n86027 , n86028 );
xnor ( n86030 , n86029 , n85759 );
and ( n86031 , n86026 , n86030 );
buf ( n86032 , n553 );
buf ( n86033 , n86032 );
and ( n86034 , n86033 , n85691 );
and ( n86035 , n86030 , n86034 );
and ( n86036 , n86026 , n86034 );
or ( n86037 , n86031 , n86035 , n86036 );
xor ( n86038 , n85957 , n85961 );
xor ( n86039 , n86038 , n85966 );
and ( n86040 , n86037 , n86039 );
xor ( n86041 , n86014 , n86019 );
xor ( n86042 , n86041 , n86022 );
and ( n86043 , n86039 , n86042 );
and ( n86044 , n86037 , n86042 );
or ( n86045 , n86040 , n86043 , n86044 );
and ( n86046 , n86025 , n86045 );
xor ( n86047 , n85969 , n85971 );
xor ( n86048 , n86047 , n85974 );
and ( n86049 , n86045 , n86048 );
and ( n86050 , n86025 , n86048 );
or ( n86051 , n86046 , n86049 , n86050 );
xor ( n86052 , n85949 , n85977 );
xor ( n86053 , n86052 , n85980 );
and ( n86054 , n86051 , n86053 );
and ( n86055 , n85994 , n86054 );
and ( n86056 , n85993 , n86054 );
or ( n86057 , n85995 , n86055 , n86056 );
xor ( n86058 , n85923 , n85924 );
xor ( n86059 , n86058 , n85986 );
and ( n86060 , n86057 , n86059 );
buf ( n86061 , n85647 );
xor ( n86062 , n86051 , n86053 );
and ( n86063 , n86061 , n86062 );
buf ( n86064 , n571 );
buf ( n86065 , n86064 );
buf ( n86066 , n572 );
buf ( n86067 , n86066 );
and ( n86068 , n86065 , n86067 );
not ( n86069 , n86068 );
and ( n86070 , n85953 , n86069 );
not ( n86071 , n86070 );
and ( n86072 , n85700 , n85999 );
and ( n86073 , n85670 , n85997 );
nor ( n86074 , n86072 , n86073 );
xnor ( n86075 , n86074 , n85956 );
and ( n86076 , n86071 , n86075 );
and ( n86077 , n85782 , n85790 );
and ( n86078 , n85767 , n85788 );
nor ( n86079 , n86077 , n86078 );
xnor ( n86080 , n86079 , n85759 );
and ( n86081 , n86075 , n86080 );
and ( n86082 , n86071 , n86080 );
or ( n86083 , n86076 , n86081 , n86082 );
and ( n86084 , n85709 , n85887 );
and ( n86085 , n85689 , n85885 );
nor ( n86086 , n86084 , n86085 );
xnor ( n86087 , n86086 , n85825 );
and ( n86088 , n85897 , n85680 );
and ( n86089 , n85879 , n85678 );
nor ( n86090 , n86088 , n86089 );
xnor ( n86091 , n86090 , n85685 );
and ( n86092 , n86087 , n86091 );
and ( n86093 , n86033 , n85697 );
and ( n86094 , n85936 , n85695 );
nor ( n86095 , n86093 , n86094 );
xnor ( n86096 , n86095 , n85705 );
and ( n86097 , n86091 , n86096 );
and ( n86098 , n86087 , n86096 );
or ( n86099 , n86092 , n86097 , n86098 );
and ( n86100 , n86083 , n86099 );
xor ( n86101 , n86002 , n86006 );
xor ( n86102 , n86101 , n86011 );
and ( n86103 , n86099 , n86102 );
and ( n86104 , n86083 , n86102 );
or ( n86105 , n86100 , n86103 , n86104 );
and ( n86106 , n85689 , n85999 );
and ( n86107 , n85700 , n85997 );
nor ( n86108 , n86106 , n86107 );
xnor ( n86109 , n86108 , n85956 );
and ( n86110 , n85879 , n85790 );
and ( n86111 , n85782 , n85788 );
nor ( n86112 , n86110 , n86111 );
xnor ( n86113 , n86112 , n85759 );
and ( n86114 , n86109 , n86113 );
and ( n86115 , n85936 , n85680 );
and ( n86116 , n85897 , n85678 );
nor ( n86117 , n86115 , n86116 );
xnor ( n86118 , n86117 , n85685 );
and ( n86119 , n86113 , n86118 );
and ( n86120 , n86109 , n86118 );
or ( n86121 , n86114 , n86119 , n86120 );
xor ( n86122 , n85953 , n86065 );
xor ( n86123 , n86065 , n86067 );
not ( n86124 , n86123 );
and ( n86125 , n86122 , n86124 );
and ( n86126 , n85670 , n86125 );
not ( n86127 , n86126 );
xnor ( n86128 , n86127 , n86070 );
buf ( n86129 , n86128 );
and ( n86130 , n86121 , n86129 );
buf ( n86131 , n554 );
buf ( n86132 , n86131 );
and ( n86133 , n86132 , n85691 );
and ( n86134 , n86129 , n86133 );
and ( n86135 , n86121 , n86133 );
or ( n86136 , n86130 , n86134 , n86135 );
and ( n86137 , n85767 , n85887 );
and ( n86138 , n85709 , n85885 );
nor ( n86139 , n86137 , n86138 );
xnor ( n86140 , n86139 , n85825 );
and ( n86141 , n86132 , n85697 );
and ( n86142 , n86033 , n85695 );
nor ( n86143 , n86141 , n86142 );
xnor ( n86144 , n86143 , n85705 );
and ( n86145 , n86140 , n86144 );
buf ( n86146 , n555 );
buf ( n86147 , n86146 );
and ( n86148 , n86147 , n85691 );
and ( n86149 , n86144 , n86148 );
and ( n86150 , n86140 , n86148 );
or ( n86151 , n86145 , n86149 , n86150 );
xor ( n86152 , n86071 , n86075 );
xor ( n86153 , n86152 , n86080 );
and ( n86154 , n86151 , n86153 );
xor ( n86155 , n86087 , n86091 );
xor ( n86156 , n86155 , n86096 );
and ( n86157 , n86153 , n86156 );
and ( n86158 , n86151 , n86156 );
or ( n86159 , n86154 , n86157 , n86158 );
and ( n86160 , n86136 , n86159 );
xor ( n86161 , n86026 , n86030 );
xor ( n86162 , n86161 , n86034 );
and ( n86163 , n86159 , n86162 );
and ( n86164 , n86136 , n86162 );
or ( n86165 , n86160 , n86163 , n86164 );
and ( n86166 , n86105 , n86165 );
xor ( n86167 , n86037 , n86039 );
xor ( n86168 , n86167 , n86042 );
and ( n86169 , n86165 , n86168 );
and ( n86170 , n86105 , n86168 );
or ( n86171 , n86166 , n86169 , n86170 );
xor ( n86172 , n86025 , n86045 );
xor ( n86173 , n86172 , n86048 );
and ( n86174 , n86171 , n86173 );
and ( n86175 , n86062 , n86174 );
and ( n86176 , n86061 , n86174 );
or ( n86177 , n86063 , n86175 , n86176 );
xor ( n86178 , n85993 , n85994 );
xor ( n86179 , n86178 , n86054 );
and ( n86180 , n86177 , n86179 );
xor ( n86181 , n86061 , n86062 );
xor ( n86182 , n86181 , n86174 );
buf ( n86183 , n85648 );
xor ( n86184 , n86171 , n86173 );
and ( n86185 , n86183 , n86184 );
and ( n86186 , n85709 , n85999 );
and ( n86187 , n85689 , n85997 );
nor ( n86188 , n86186 , n86187 );
xnor ( n86189 , n86188 , n85956 );
and ( n86190 , n85897 , n85790 );
and ( n86191 , n85879 , n85788 );
nor ( n86192 , n86190 , n86191 );
xnor ( n86193 , n86192 , n85759 );
and ( n86194 , n86189 , n86193 );
buf ( n86195 , n556 );
buf ( n86196 , n86195 );
and ( n86197 , n86196 , n85691 );
and ( n86198 , n86193 , n86197 );
and ( n86199 , n86189 , n86197 );
or ( n86200 , n86194 , n86198 , n86199 );
buf ( n86201 , n573 );
buf ( n86202 , n86201 );
buf ( n86203 , n574 );
buf ( n86204 , n86203 );
and ( n86205 , n86202 , n86204 );
not ( n86206 , n86205 );
and ( n86207 , n86067 , n86206 );
not ( n86208 , n86207 );
and ( n86209 , n85700 , n86125 );
and ( n86210 , n85670 , n86123 );
nor ( n86211 , n86209 , n86210 );
xnor ( n86212 , n86211 , n86070 );
and ( n86213 , n86208 , n86212 );
and ( n86214 , n85782 , n85887 );
and ( n86215 , n85767 , n85885 );
nor ( n86216 , n86214 , n86215 );
xnor ( n86217 , n86216 , n85825 );
and ( n86218 , n86212 , n86217 );
and ( n86219 , n86208 , n86217 );
or ( n86220 , n86213 , n86218 , n86219 );
and ( n86221 , n86200 , n86220 );
not ( n86222 , n86128 );
and ( n86223 , n86220 , n86222 );
and ( n86224 , n86200 , n86222 );
or ( n86225 , n86221 , n86223 , n86224 );
xor ( n86226 , n86067 , n86202 );
xor ( n86227 , n86202 , n86204 );
not ( n86228 , n86227 );
and ( n86229 , n86226 , n86228 );
and ( n86230 , n85670 , n86229 );
not ( n86231 , n86230 );
xnor ( n86232 , n86231 , n86207 );
buf ( n86233 , n86232 );
and ( n86234 , n86033 , n85680 );
and ( n86235 , n85936 , n85678 );
nor ( n86236 , n86234 , n86235 );
xnor ( n86237 , n86236 , n85685 );
and ( n86238 , n86233 , n86237 );
and ( n86239 , n86147 , n85697 );
and ( n86240 , n86132 , n85695 );
nor ( n86241 , n86239 , n86240 );
xnor ( n86242 , n86241 , n85705 );
and ( n86243 , n86237 , n86242 );
and ( n86244 , n86233 , n86242 );
or ( n86245 , n86238 , n86243 , n86244 );
xor ( n86246 , n86140 , n86144 );
xor ( n86247 , n86246 , n86148 );
and ( n86248 , n86245 , n86247 );
xor ( n86249 , n86109 , n86113 );
xor ( n86250 , n86249 , n86118 );
and ( n86251 , n86247 , n86250 );
and ( n86252 , n86245 , n86250 );
or ( n86253 , n86248 , n86251 , n86252 );
and ( n86254 , n86225 , n86253 );
xor ( n86255 , n86121 , n86129 );
xor ( n86256 , n86255 , n86133 );
and ( n86257 , n86253 , n86256 );
and ( n86258 , n86225 , n86256 );
or ( n86259 , n86254 , n86257 , n86258 );
xor ( n86260 , n86083 , n86099 );
xor ( n86261 , n86260 , n86102 );
and ( n86262 , n86259 , n86261 );
xor ( n86263 , n86136 , n86159 );
xor ( n86264 , n86263 , n86162 );
and ( n86265 , n86261 , n86264 );
and ( n86266 , n86259 , n86264 );
or ( n86267 , n86262 , n86265 , n86266 );
xor ( n86268 , n86105 , n86165 );
xor ( n86269 , n86268 , n86168 );
and ( n86270 , n86267 , n86269 );
and ( n86271 , n86184 , n86270 );
and ( n86272 , n86183 , n86270 );
or ( n86273 , n86185 , n86271 , n86272 );
and ( n86274 , n86182 , n86273 );
buf ( n86275 , n85649 );
xor ( n86276 , n86267 , n86269 );
and ( n86277 , n86275 , n86276 );
and ( n86278 , n85689 , n86125 );
and ( n86279 , n85700 , n86123 );
nor ( n86280 , n86278 , n86279 );
xnor ( n86281 , n86280 , n86070 );
and ( n86282 , n85879 , n85887 );
and ( n86283 , n85782 , n85885 );
nor ( n86284 , n86282 , n86283 );
xnor ( n86285 , n86284 , n85825 );
and ( n86286 , n86281 , n86285 );
buf ( n86287 , n557 );
buf ( n86288 , n86287 );
and ( n86289 , n86288 , n85691 );
and ( n86290 , n86285 , n86289 );
and ( n86291 , n86281 , n86289 );
or ( n86292 , n86286 , n86290 , n86291 );
and ( n86293 , n85767 , n85999 );
and ( n86294 , n85709 , n85997 );
nor ( n86295 , n86293 , n86294 );
xnor ( n86296 , n86295 , n85956 );
and ( n86297 , n85936 , n85790 );
and ( n86298 , n85897 , n85788 );
nor ( n86299 , n86297 , n86298 );
xnor ( n86300 , n86299 , n85759 );
and ( n86301 , n86296 , n86300 );
and ( n86302 , n86132 , n85680 );
and ( n86303 , n86033 , n85678 );
nor ( n86304 , n86302 , n86303 );
xnor ( n86305 , n86304 , n85685 );
and ( n86306 , n86300 , n86305 );
and ( n86307 , n86296 , n86305 );
or ( n86308 , n86301 , n86306 , n86307 );
and ( n86309 , n86292 , n86308 );
xor ( n86310 , n86208 , n86212 );
xor ( n86311 , n86310 , n86217 );
and ( n86312 , n86308 , n86311 );
and ( n86313 , n86292 , n86311 );
or ( n86314 , n86309 , n86312 , n86313 );
xor ( n86315 , n86200 , n86220 );
xor ( n86316 , n86315 , n86222 );
and ( n86317 , n86314 , n86316 );
xor ( n86318 , n86245 , n86247 );
xor ( n86319 , n86318 , n86250 );
and ( n86320 , n86316 , n86319 );
and ( n86321 , n86314 , n86319 );
or ( n86322 , n86317 , n86320 , n86321 );
xor ( n86323 , n86151 , n86153 );
xor ( n86324 , n86323 , n86156 );
and ( n86325 , n86322 , n86324 );
xor ( n86326 , n86225 , n86253 );
xor ( n86327 , n86326 , n86256 );
and ( n86328 , n86324 , n86327 );
and ( n86329 , n86322 , n86327 );
or ( n86330 , n86325 , n86328 , n86329 );
xor ( n86331 , n86259 , n86261 );
xor ( n86332 , n86331 , n86264 );
and ( n86333 , n86330 , n86332 );
and ( n86334 , n86276 , n86333 );
and ( n86335 , n86275 , n86333 );
or ( n86336 , n86277 , n86334 , n86335 );
xor ( n86337 , n86183 , n86184 );
xor ( n86338 , n86337 , n86270 );
and ( n86339 , n86336 , n86338 );
buf ( n86340 , n85650 );
xor ( n86341 , n86330 , n86332 );
and ( n86342 , n86340 , n86341 );
and ( n86343 , n85782 , n85999 );
and ( n86344 , n85767 , n85997 );
nor ( n86345 , n86343 , n86344 );
xnor ( n86346 , n86345 , n85956 );
buf ( n86347 , n86346 );
not ( n86348 , n86232 );
and ( n86349 , n86347 , n86348 );
and ( n86350 , n86196 , n85697 );
and ( n86351 , n86147 , n85695 );
nor ( n86352 , n86350 , n86351 );
xnor ( n86353 , n86352 , n85705 );
and ( n86354 , n86348 , n86353 );
and ( n86355 , n86347 , n86353 );
or ( n86356 , n86349 , n86354 , n86355 );
xor ( n86357 , n86189 , n86193 );
xor ( n86358 , n86357 , n86197 );
and ( n86359 , n86356 , n86358 );
xor ( n86360 , n86233 , n86237 );
xor ( n86361 , n86360 , n86242 );
and ( n86362 , n86358 , n86361 );
and ( n86363 , n86356 , n86361 );
or ( n86364 , n86359 , n86362 , n86363 );
not ( n86365 , n86204 );
and ( n86366 , n86288 , n85697 );
and ( n86367 , n86196 , n85695 );
nor ( n86368 , n86366 , n86367 );
xnor ( n86369 , n86368 , n85705 );
and ( n86370 , n86365 , n86369 );
buf ( n86371 , n558 );
buf ( n86372 , n86371 );
and ( n86373 , n86372 , n85691 );
and ( n86374 , n86369 , n86373 );
and ( n86375 , n86365 , n86373 );
or ( n86376 , n86370 , n86374 , n86375 );
and ( n86377 , n85700 , n86229 );
and ( n86378 , n85670 , n86227 );
nor ( n86379 , n86377 , n86378 );
xnor ( n86380 , n86379 , n86207 );
and ( n86381 , n85709 , n86125 );
and ( n86382 , n85689 , n86123 );
nor ( n86383 , n86381 , n86382 );
xnor ( n86384 , n86383 , n86070 );
and ( n86385 , n86380 , n86384 );
and ( n86386 , n85897 , n85887 );
and ( n86387 , n85879 , n85885 );
nor ( n86388 , n86386 , n86387 );
xnor ( n86389 , n86388 , n85825 );
and ( n86390 , n86384 , n86389 );
and ( n86391 , n86380 , n86389 );
or ( n86392 , n86385 , n86390 , n86391 );
and ( n86393 , n86376 , n86392 );
xor ( n86394 , n86296 , n86300 );
xor ( n86395 , n86394 , n86305 );
and ( n86396 , n86392 , n86395 );
and ( n86397 , n86376 , n86395 );
or ( n86398 , n86393 , n86396 , n86397 );
buf ( n86399 , n575 );
buf ( n86400 , n86399 );
xor ( n86401 , n86204 , n86400 );
not ( n86402 , n86400 );
and ( n86403 , n86401 , n86402 );
and ( n86404 , n85670 , n86403 );
not ( n86405 , n86404 );
xnor ( n86406 , n86405 , n86204 );
and ( n86407 , n85689 , n86229 );
and ( n86408 , n85700 , n86227 );
nor ( n86409 , n86407 , n86408 );
xnor ( n86410 , n86409 , n86207 );
and ( n86411 , n86406 , n86410 );
buf ( n86412 , n559 );
buf ( n86413 , n86412 );
and ( n86414 , n86413 , n85691 );
and ( n86415 , n86410 , n86414 );
and ( n86416 , n86406 , n86414 );
or ( n86417 , n86411 , n86415 , n86416 );
and ( n86418 , n85767 , n86125 );
and ( n86419 , n85709 , n86123 );
nor ( n86420 , n86418 , n86419 );
xnor ( n86421 , n86420 , n86070 );
and ( n86422 , n86132 , n85790 );
and ( n86423 , n86033 , n85788 );
nor ( n86424 , n86422 , n86423 );
xnor ( n86425 , n86424 , n85759 );
and ( n86426 , n86421 , n86425 );
and ( n86427 , n86196 , n85680 );
and ( n86428 , n86147 , n85678 );
nor ( n86429 , n86427 , n86428 );
xnor ( n86430 , n86429 , n85685 );
and ( n86431 , n86425 , n86430 );
and ( n86432 , n86421 , n86430 );
or ( n86433 , n86426 , n86431 , n86432 );
and ( n86434 , n86417 , n86433 );
and ( n86435 , n85879 , n85999 );
and ( n86436 , n85782 , n85997 );
nor ( n86437 , n86435 , n86436 );
xnor ( n86438 , n86437 , n85956 );
and ( n86439 , n85936 , n85887 );
and ( n86440 , n85897 , n85885 );
nor ( n86441 , n86439 , n86440 );
xnor ( n86442 , n86441 , n85825 );
and ( n86443 , n86438 , n86442 );
and ( n86444 , n86372 , n85697 );
and ( n86445 , n86288 , n85695 );
nor ( n86446 , n86444 , n86445 );
xnor ( n86447 , n86446 , n85705 );
and ( n86448 , n86442 , n86447 );
and ( n86449 , n86438 , n86447 );
or ( n86450 , n86443 , n86448 , n86449 );
and ( n86451 , n86433 , n86450 );
and ( n86452 , n86417 , n86450 );
or ( n86453 , n86434 , n86451 , n86452 );
xor ( n86454 , n86281 , n86285 );
xor ( n86455 , n86454 , n86289 );
and ( n86456 , n86453 , n86455 );
xor ( n86457 , n86347 , n86348 );
xor ( n86458 , n86457 , n86353 );
and ( n86459 , n86455 , n86458 );
and ( n86460 , n86453 , n86458 );
or ( n86461 , n86456 , n86459 , n86460 );
and ( n86462 , n86398 , n86461 );
xor ( n86463 , n86292 , n86308 );
xor ( n86464 , n86463 , n86311 );
and ( n86465 , n86461 , n86464 );
and ( n86466 , n86398 , n86464 );
or ( n86467 , n86462 , n86465 , n86466 );
and ( n86468 , n86364 , n86467 );
xor ( n86469 , n86314 , n86316 );
xor ( n86470 , n86469 , n86319 );
and ( n86471 , n86467 , n86470 );
and ( n86472 , n86364 , n86470 );
or ( n86473 , n86468 , n86471 , n86472 );
xor ( n86474 , n86322 , n86324 );
xor ( n86475 , n86474 , n86327 );
and ( n86476 , n86473 , n86475 );
and ( n86477 , n86341 , n86476 );
and ( n86478 , n86340 , n86476 );
or ( n86479 , n86342 , n86477 , n86478 );
xor ( n86480 , n86275 , n86276 );
xor ( n86481 , n86480 , n86333 );
and ( n86482 , n86479 , n86481 );
buf ( n86483 , n85651 );
xor ( n86484 , n86473 , n86475 );
and ( n86485 , n86483 , n86484 );
not ( n86486 , n86346 );
and ( n86487 , n86033 , n85790 );
and ( n86488 , n85936 , n85788 );
nor ( n86489 , n86487 , n86488 );
xnor ( n86490 , n86489 , n85759 );
and ( n86491 , n86486 , n86490 );
and ( n86492 , n86147 , n85680 );
and ( n86493 , n86132 , n85678 );
nor ( n86494 , n86492 , n86493 );
xnor ( n86495 , n86494 , n85685 );
and ( n86496 , n86490 , n86495 );
and ( n86497 , n86486 , n86495 );
or ( n86498 , n86491 , n86496 , n86497 );
and ( n86499 , n85782 , n86125 );
and ( n86500 , n85767 , n86123 );
nor ( n86501 , n86499 , n86500 );
xnor ( n86502 , n86501 , n86070 );
and ( n86503 , n86033 , n85887 );
and ( n86504 , n85936 , n85885 );
nor ( n86505 , n86503 , n86504 );
xnor ( n86506 , n86505 , n85825 );
and ( n86507 , n86502 , n86506 );
and ( n86508 , n86147 , n85790 );
and ( n86509 , n86132 , n85788 );
nor ( n86510 , n86508 , n86509 );
xnor ( n86511 , n86510 , n85759 );
and ( n86512 , n86506 , n86511 );
and ( n86513 , n86502 , n86511 );
or ( n86514 , n86507 , n86512 , n86513 );
and ( n86515 , n85709 , n86229 );
and ( n86516 , n85689 , n86227 );
nor ( n86517 , n86515 , n86516 );
xnor ( n86518 , n86517 , n86207 );
and ( n86519 , n85897 , n85999 );
and ( n86520 , n85879 , n85997 );
nor ( n86521 , n86519 , n86520 );
xnor ( n86522 , n86521 , n85956 );
and ( n86523 , n86518 , n86522 );
and ( n86524 , n86413 , n85697 );
and ( n86525 , n86372 , n85695 );
nor ( n86526 , n86524 , n86525 );
xnor ( n86527 , n86526 , n85705 );
and ( n86528 , n86522 , n86527 );
and ( n86529 , n86518 , n86527 );
or ( n86530 , n86523 , n86528 , n86529 );
and ( n86531 , n86514 , n86530 );
and ( n86532 , n85700 , n86403 );
and ( n86533 , n85670 , n86400 );
nor ( n86534 , n86532 , n86533 );
xnor ( n86535 , n86534 , n86204 );
and ( n86536 , n86413 , n85695 );
not ( n86537 , n86536 );
and ( n86538 , n86537 , n85705 );
and ( n86539 , n86535 , n86538 );
and ( n86540 , n86530 , n86539 );
and ( n86541 , n86514 , n86539 );
or ( n86542 , n86531 , n86540 , n86541 );
xor ( n86543 , n86365 , n86369 );
xor ( n86544 , n86543 , n86373 );
and ( n86545 , n86542 , n86544 );
xor ( n86546 , n86380 , n86384 );
xor ( n86547 , n86546 , n86389 );
and ( n86548 , n86544 , n86547 );
and ( n86549 , n86542 , n86547 );
or ( n86550 , n86545 , n86548 , n86549 );
and ( n86551 , n86498 , n86550 );
xor ( n86552 , n86376 , n86392 );
xor ( n86553 , n86552 , n86395 );
and ( n86554 , n86550 , n86553 );
and ( n86555 , n86498 , n86553 );
or ( n86556 , n86551 , n86554 , n86555 );
xor ( n86557 , n86356 , n86358 );
xor ( n86558 , n86557 , n86361 );
and ( n86559 , n86556 , n86558 );
xor ( n86560 , n86398 , n86461 );
xor ( n86561 , n86560 , n86464 );
and ( n86562 , n86558 , n86561 );
and ( n86563 , n86556 , n86561 );
or ( n86564 , n86559 , n86562 , n86563 );
xor ( n86565 , n86364 , n86467 );
xor ( n86566 , n86565 , n86470 );
and ( n86567 , n86564 , n86566 );
and ( n86568 , n86484 , n86567 );
and ( n86569 , n86483 , n86567 );
or ( n86570 , n86485 , n86568 , n86569 );
xor ( n86571 , n86340 , n86341 );
xor ( n86572 , n86571 , n86476 );
and ( n86573 , n86570 , n86572 );
buf ( n86574 , n85652 );
xor ( n86575 , n86406 , n86410 );
xor ( n86576 , n86575 , n86414 );
xor ( n86577 , n86421 , n86425 );
xor ( n86578 , n86577 , n86430 );
and ( n86579 , n86576 , n86578 );
xor ( n86580 , n86438 , n86442 );
xor ( n86581 , n86580 , n86447 );
and ( n86582 , n86578 , n86581 );
and ( n86583 , n86576 , n86581 );
or ( n86584 , n86579 , n86582 , n86583 );
xor ( n86585 , n86417 , n86433 );
xor ( n86586 , n86585 , n86450 );
and ( n86587 , n86584 , n86586 );
xor ( n86588 , n86486 , n86490 );
xor ( n86589 , n86588 , n86495 );
and ( n86590 , n86586 , n86589 );
and ( n86591 , n86584 , n86589 );
or ( n86592 , n86587 , n86590 , n86591 );
xor ( n86593 , n86453 , n86455 );
xor ( n86594 , n86593 , n86458 );
and ( n86595 , n86592 , n86594 );
xor ( n86596 , n86498 , n86550 );
xor ( n86597 , n86596 , n86553 );
and ( n86598 , n86594 , n86597 );
and ( n86599 , n86592 , n86597 );
or ( n86600 , n86595 , n86598 , n86599 );
xor ( n86601 , n86556 , n86558 );
xor ( n86602 , n86601 , n86561 );
and ( n86603 , n86600 , n86602 );
and ( n86604 , n86574 , n86603 );
xor ( n86605 , n86564 , n86566 );
and ( n86606 , n86603 , n86605 );
and ( n86607 , n86574 , n86605 );
or ( n86608 , n86604 , n86606 , n86607 );
xor ( n86609 , n86483 , n86484 );
xor ( n86610 , n86609 , n86567 );
and ( n86611 , n86608 , n86610 );
buf ( n86612 , n85653 );
xor ( n86613 , n86600 , n86602 );
and ( n86614 , n86612 , n86613 );
xor ( n86615 , n86535 , n86538 );
and ( n86616 , n85689 , n86403 );
and ( n86617 , n85700 , n86400 );
nor ( n86618 , n86616 , n86617 );
xnor ( n86619 , n86618 , n86204 );
and ( n86620 , n85767 , n86229 );
and ( n86621 , n85709 , n86227 );
nor ( n86622 , n86620 , n86621 );
xnor ( n86623 , n86622 , n86207 );
and ( n86624 , n86619 , n86623 );
and ( n86625 , n86623 , n86536 );
and ( n86626 , n86619 , n86536 );
or ( n86627 , n86624 , n86625 , n86626 );
and ( n86628 , n86615 , n86627 );
and ( n86629 , n86288 , n85680 );
and ( n86630 , n86196 , n85678 );
nor ( n86631 , n86629 , n86630 );
xnor ( n86632 , n86631 , n85685 );
and ( n86633 , n86627 , n86632 );
and ( n86634 , n86615 , n86632 );
or ( n86635 , n86628 , n86633 , n86634 );
and ( n86636 , n85879 , n86125 );
and ( n86637 , n85782 , n86123 );
nor ( n86638 , n86636 , n86637 );
xnor ( n86639 , n86638 , n86070 );
and ( n86640 , n85936 , n85999 );
and ( n86641 , n85897 , n85997 );
nor ( n86642 , n86640 , n86641 );
xnor ( n86643 , n86642 , n85956 );
and ( n86644 , n86639 , n86643 );
and ( n86645 , n86132 , n85887 );
and ( n86646 , n86033 , n85885 );
nor ( n86647 , n86645 , n86646 );
xnor ( n86648 , n86647 , n85825 );
and ( n86649 , n86643 , n86648 );
and ( n86650 , n86639 , n86648 );
or ( n86651 , n86644 , n86649 , n86650 );
xor ( n86652 , n86502 , n86506 );
xor ( n86653 , n86652 , n86511 );
and ( n86654 , n86651 , n86653 );
xor ( n86655 , n86518 , n86522 );
xor ( n86656 , n86655 , n86527 );
and ( n86657 , n86653 , n86656 );
and ( n86658 , n86651 , n86656 );
or ( n86659 , n86654 , n86657 , n86658 );
and ( n86660 , n86635 , n86659 );
xor ( n86661 , n86514 , n86530 );
xor ( n86662 , n86661 , n86539 );
and ( n86663 , n86659 , n86662 );
and ( n86664 , n86635 , n86662 );
or ( n86665 , n86660 , n86663 , n86664 );
xor ( n86666 , n86542 , n86544 );
xor ( n86667 , n86666 , n86547 );
and ( n86668 , n86665 , n86667 );
xor ( n86669 , n86584 , n86586 );
xor ( n86670 , n86669 , n86589 );
and ( n86671 , n86667 , n86670 );
and ( n86672 , n86665 , n86670 );
or ( n86673 , n86668 , n86671 , n86672 );
xor ( n86674 , n86592 , n86594 );
xor ( n86675 , n86674 , n86597 );
and ( n86676 , n86673 , n86675 );
and ( n86677 , n86613 , n86676 );
and ( n86678 , n86612 , n86676 );
or ( n86679 , n86614 , n86677 , n86678 );
xor ( n86680 , n86574 , n86603 );
xor ( n86681 , n86680 , n86605 );
and ( n86682 , n86679 , n86681 );
buf ( n86683 , n85654 );
and ( n86684 , n85709 , n86403 );
and ( n86685 , n85689 , n86400 );
nor ( n86686 , n86684 , n86685 );
xnor ( n86687 , n86686 , n86204 );
and ( n86688 , n86413 , n85678 );
not ( n86689 , n86688 );
and ( n86690 , n86689 , n85685 );
and ( n86691 , n86687 , n86690 );
and ( n86692 , n86196 , n85790 );
and ( n86693 , n86147 , n85788 );
nor ( n86694 , n86692 , n86693 );
xnor ( n86695 , n86694 , n85759 );
and ( n86696 , n86691 , n86695 );
and ( n86697 , n86372 , n85680 );
and ( n86698 , n86288 , n85678 );
nor ( n86699 , n86697 , n86698 );
xnor ( n86700 , n86699 , n85685 );
and ( n86701 , n86695 , n86700 );
and ( n86702 , n86691 , n86700 );
or ( n86703 , n86696 , n86701 , n86702 );
and ( n86704 , n85897 , n86125 );
and ( n86705 , n85879 , n86123 );
nor ( n86706 , n86704 , n86705 );
xnor ( n86707 , n86706 , n86070 );
and ( n86708 , n86288 , n85790 );
and ( n86709 , n86196 , n85788 );
nor ( n86710 , n86708 , n86709 );
xnor ( n86711 , n86710 , n85759 );
and ( n86712 , n86707 , n86711 );
and ( n86713 , n86413 , n85680 );
and ( n86714 , n86372 , n85678 );
nor ( n86715 , n86713 , n86714 );
xnor ( n86716 , n86715 , n85685 );
and ( n86717 , n86711 , n86716 );
and ( n86718 , n86707 , n86716 );
or ( n86719 , n86712 , n86717 , n86718 );
and ( n86720 , n85782 , n86229 );
and ( n86721 , n85767 , n86227 );
nor ( n86722 , n86720 , n86721 );
xnor ( n86723 , n86722 , n86207 );
and ( n86724 , n86033 , n85999 );
and ( n86725 , n85936 , n85997 );
nor ( n86726 , n86724 , n86725 );
xnor ( n86727 , n86726 , n85956 );
and ( n86728 , n86723 , n86727 );
and ( n86729 , n86147 , n85887 );
and ( n86730 , n86132 , n85885 );
nor ( n86731 , n86729 , n86730 );
xnor ( n86732 , n86731 , n85825 );
and ( n86733 , n86727 , n86732 );
and ( n86734 , n86723 , n86732 );
or ( n86735 , n86728 , n86733 , n86734 );
and ( n86736 , n86719 , n86735 );
xor ( n86737 , n86619 , n86623 );
xor ( n86738 , n86737 , n86536 );
and ( n86739 , n86735 , n86738 );
and ( n86740 , n86719 , n86738 );
or ( n86741 , n86736 , n86739 , n86740 );
and ( n86742 , n86703 , n86741 );
xor ( n86743 , n86615 , n86627 );
xor ( n86744 , n86743 , n86632 );
and ( n86745 , n86741 , n86744 );
and ( n86746 , n86703 , n86744 );
or ( n86747 , n86742 , n86745 , n86746 );
xor ( n86748 , n86576 , n86578 );
xor ( n86749 , n86748 , n86581 );
and ( n86750 , n86747 , n86749 );
xor ( n86751 , n86635 , n86659 );
xor ( n86752 , n86751 , n86662 );
and ( n86753 , n86749 , n86752 );
and ( n86754 , n86747 , n86752 );
or ( n86755 , n86750 , n86753 , n86754 );
xor ( n86756 , n86665 , n86667 );
xor ( n86757 , n86756 , n86670 );
and ( n86758 , n86755 , n86757 );
and ( n86759 , n86683 , n86758 );
xor ( n86760 , n86673 , n86675 );
and ( n86761 , n86758 , n86760 );
and ( n86762 , n86683 , n86760 );
or ( n86763 , n86759 , n86761 , n86762 );
xor ( n86764 , n86612 , n86613 );
xor ( n86765 , n86764 , n86676 );
and ( n86766 , n86763 , n86765 );
buf ( n86767 , n85655 );
xor ( n86768 , n86755 , n86757 );
and ( n86769 , n86767 , n86768 );
xor ( n86770 , n86687 , n86690 );
and ( n86771 , n85767 , n86403 );
and ( n86772 , n85709 , n86400 );
nor ( n86773 , n86771 , n86772 );
xnor ( n86774 , n86773 , n86204 );
and ( n86775 , n86196 , n85887 );
and ( n86776 , n86147 , n85885 );
nor ( n86777 , n86775 , n86776 );
xnor ( n86778 , n86777 , n85825 );
and ( n86779 , n86774 , n86778 );
and ( n86780 , n86372 , n85790 );
and ( n86781 , n86288 , n85788 );
nor ( n86782 , n86780 , n86781 );
xnor ( n86783 , n86782 , n85759 );
and ( n86784 , n86778 , n86783 );
and ( n86785 , n86774 , n86783 );
or ( n86786 , n86779 , n86784 , n86785 );
and ( n86787 , n86770 , n86786 );
and ( n86788 , n85879 , n86229 );
and ( n86789 , n85782 , n86227 );
nor ( n86790 , n86788 , n86789 );
xnor ( n86791 , n86790 , n86207 );
and ( n86792 , n86132 , n85999 );
and ( n86793 , n86033 , n85997 );
nor ( n86794 , n86792 , n86793 );
xnor ( n86795 , n86794 , n85956 );
and ( n86796 , n86791 , n86795 );
and ( n86797 , n86795 , n86688 );
and ( n86798 , n86791 , n86688 );
or ( n86799 , n86796 , n86797 , n86798 );
and ( n86800 , n86786 , n86799 );
and ( n86801 , n86770 , n86799 );
or ( n86802 , n86787 , n86800 , n86801 );
xor ( n86803 , n86639 , n86643 );
xor ( n86804 , n86803 , n86648 );
and ( n86805 , n86802 , n86804 );
xor ( n86806 , n86691 , n86695 );
xor ( n86807 , n86806 , n86700 );
and ( n86808 , n86804 , n86807 );
and ( n86809 , n86802 , n86807 );
or ( n86810 , n86805 , n86808 , n86809 );
xor ( n86811 , n86651 , n86653 );
xor ( n86812 , n86811 , n86656 );
and ( n86813 , n86810 , n86812 );
xor ( n86814 , n86703 , n86741 );
xor ( n86815 , n86814 , n86744 );
and ( n86816 , n86812 , n86815 );
and ( n86817 , n86810 , n86815 );
or ( n86818 , n86813 , n86816 , n86817 );
xor ( n86819 , n86747 , n86749 );
xor ( n86820 , n86819 , n86752 );
and ( n86821 , n86818 , n86820 );
and ( n86822 , n86768 , n86821 );
and ( n86823 , n86767 , n86821 );
or ( n86824 , n86769 , n86822 , n86823 );
xor ( n86825 , n86683 , n86758 );
xor ( n86826 , n86825 , n86760 );
and ( n86827 , n86824 , n86826 );
buf ( n86828 , n85656 );
xor ( n86829 , n86818 , n86820 );
and ( n86830 , n86828 , n86829 );
and ( n86831 , n85782 , n86403 );
and ( n86832 , n85767 , n86400 );
nor ( n86833 , n86831 , n86832 );
xnor ( n86834 , n86833 , n86204 );
and ( n86835 , n86147 , n85999 );
and ( n86836 , n86132 , n85997 );
nor ( n86837 , n86835 , n86836 );
xnor ( n86838 , n86837 , n85956 );
and ( n86839 , n86834 , n86838 );
and ( n86840 , n86288 , n85887 );
and ( n86841 , n86196 , n85885 );
nor ( n86842 , n86840 , n86841 );
xnor ( n86843 , n86842 , n85825 );
and ( n86844 , n86838 , n86843 );
and ( n86845 , n86834 , n86843 );
or ( n86846 , n86839 , n86844 , n86845 );
and ( n86847 , n85897 , n86229 );
and ( n86848 , n85879 , n86227 );
nor ( n86849 , n86847 , n86848 );
xnor ( n86850 , n86849 , n86207 );
and ( n86851 , n86413 , n85788 );
not ( n86852 , n86851 );
and ( n86853 , n86852 , n85759 );
and ( n86854 , n86850 , n86853 );
and ( n86855 , n86846 , n86854 );
and ( n86856 , n85936 , n86125 );
and ( n86857 , n85897 , n86123 );
nor ( n86858 , n86856 , n86857 );
xnor ( n86859 , n86858 , n86070 );
and ( n86860 , n86854 , n86859 );
and ( n86861 , n86846 , n86859 );
or ( n86862 , n86855 , n86860 , n86861 );
xor ( n86863 , n86707 , n86711 );
xor ( n86864 , n86863 , n86716 );
and ( n86865 , n86862 , n86864 );
xor ( n86866 , n86723 , n86727 );
xor ( n86867 , n86866 , n86732 );
and ( n86868 , n86864 , n86867 );
and ( n86869 , n86862 , n86867 );
or ( n86870 , n86865 , n86868 , n86869 );
xor ( n86871 , n86719 , n86735 );
xor ( n86872 , n86871 , n86738 );
and ( n86873 , n86870 , n86872 );
xor ( n86874 , n86802 , n86804 );
xor ( n86875 , n86874 , n86807 );
and ( n86876 , n86872 , n86875 );
and ( n86877 , n86870 , n86875 );
or ( n86878 , n86873 , n86876 , n86877 );
xor ( n86879 , n86810 , n86812 );
xor ( n86880 , n86879 , n86815 );
and ( n86881 , n86878 , n86880 );
and ( n86882 , n86829 , n86881 );
and ( n86883 , n86828 , n86881 );
or ( n86884 , n86830 , n86882 , n86883 );
xor ( n86885 , n86767 , n86768 );
xor ( n86886 , n86885 , n86821 );
and ( n86887 , n86884 , n86886 );
buf ( n86888 , n85657 );
xor ( n86889 , n86878 , n86880 );
and ( n86890 , n86888 , n86889 );
xor ( n86891 , n86850 , n86853 );
and ( n86892 , n86033 , n86125 );
and ( n86893 , n85936 , n86123 );
nor ( n86894 , n86892 , n86893 );
xnor ( n86895 , n86894 , n86070 );
and ( n86896 , n86891 , n86895 );
and ( n86897 , n86413 , n85790 );
and ( n86898 , n86372 , n85788 );
nor ( n86899 , n86897 , n86898 );
xnor ( n86900 , n86899 , n85759 );
and ( n86901 , n86895 , n86900 );
and ( n86902 , n86891 , n86900 );
or ( n86903 , n86896 , n86901 , n86902 );
xor ( n86904 , n86774 , n86778 );
xor ( n86905 , n86904 , n86783 );
and ( n86906 , n86903 , n86905 );
xor ( n86907 , n86791 , n86795 );
xor ( n86908 , n86907 , n86688 );
and ( n86909 , n86905 , n86908 );
and ( n86910 , n86903 , n86908 );
or ( n86911 , n86906 , n86909 , n86910 );
xor ( n86912 , n86770 , n86786 );
xor ( n86913 , n86912 , n86799 );
and ( n86914 , n86911 , n86913 );
xor ( n86915 , n86862 , n86864 );
xor ( n86916 , n86915 , n86867 );
and ( n86917 , n86913 , n86916 );
and ( n86918 , n86911 , n86916 );
or ( n86919 , n86914 , n86917 , n86918 );
xor ( n86920 , n86870 , n86872 );
xor ( n86921 , n86920 , n86875 );
and ( n86922 , n86919 , n86921 );
and ( n86923 , n86889 , n86922 );
and ( n86924 , n86888 , n86922 );
or ( n86925 , n86890 , n86923 , n86924 );
xor ( n86926 , n86828 , n86829 );
xor ( n86927 , n86926 , n86881 );
and ( n86928 , n86925 , n86927 );
buf ( n86929 , n85658 );
xor ( n86930 , n86919 , n86921 );
and ( n86931 , n86929 , n86930 );
and ( n86932 , n85879 , n86403 );
and ( n86933 , n85782 , n86400 );
nor ( n86934 , n86932 , n86933 );
xnor ( n86935 , n86934 , n86204 );
and ( n86936 , n86132 , n86125 );
and ( n86937 , n86033 , n86123 );
nor ( n86938 , n86936 , n86937 );
xnor ( n86939 , n86938 , n86070 );
and ( n86940 , n86935 , n86939 );
and ( n86941 , n86372 , n85887 );
and ( n86942 , n86288 , n85885 );
nor ( n86943 , n86941 , n86942 );
xnor ( n86944 , n86943 , n85825 );
and ( n86945 , n86939 , n86944 );
and ( n86946 , n86935 , n86944 );
or ( n86947 , n86940 , n86945 , n86946 );
and ( n86948 , n85936 , n86229 );
and ( n86949 , n85897 , n86227 );
nor ( n86950 , n86948 , n86949 );
xnor ( n86951 , n86950 , n86207 );
and ( n86952 , n86196 , n85999 );
and ( n86953 , n86147 , n85997 );
nor ( n86954 , n86952 , n86953 );
xnor ( n86955 , n86954 , n85956 );
and ( n86956 , n86951 , n86955 );
and ( n86957 , n86955 , n86851 );
and ( n86958 , n86951 , n86851 );
or ( n86959 , n86956 , n86957 , n86958 );
and ( n86960 , n86947 , n86959 );
xor ( n86961 , n86834 , n86838 );
xor ( n86962 , n86961 , n86843 );
and ( n86963 , n86959 , n86962 );
and ( n86964 , n86947 , n86962 );
or ( n86965 , n86960 , n86963 , n86964 );
xor ( n86966 , n86846 , n86854 );
xor ( n86967 , n86966 , n86859 );
and ( n86968 , n86965 , n86967 );
xor ( n86969 , n86903 , n86905 );
xor ( n86970 , n86969 , n86908 );
and ( n86971 , n86967 , n86970 );
and ( n86972 , n86965 , n86970 );
or ( n86973 , n86968 , n86971 , n86972 );
xor ( n86974 , n86911 , n86913 );
xor ( n86975 , n86974 , n86916 );
and ( n86976 , n86973 , n86975 );
and ( n86977 , n86930 , n86976 );
and ( n86978 , n86929 , n86976 );
or ( n86979 , n86931 , n86977 , n86978 );
xor ( n86980 , n86888 , n86889 );
xor ( n86981 , n86980 , n86922 );
and ( n86982 , n86979 , n86981 );
buf ( n86983 , n85659 );
xor ( n86984 , n86973 , n86975 );
and ( n86985 , n86983 , n86984 );
and ( n86986 , n85897 , n86403 );
and ( n86987 , n85879 , n86400 );
nor ( n86988 , n86986 , n86987 );
xnor ( n86989 , n86988 , n86204 );
and ( n86990 , n86288 , n85999 );
and ( n86991 , n86196 , n85997 );
nor ( n86992 , n86990 , n86991 );
xnor ( n86993 , n86992 , n85956 );
and ( n86994 , n86989 , n86993 );
and ( n86995 , n86413 , n85887 );
and ( n86996 , n86372 , n85885 );
nor ( n86997 , n86995 , n86996 );
xnor ( n86998 , n86997 , n85825 );
and ( n86999 , n86993 , n86998 );
and ( n87000 , n86989 , n86998 );
or ( n87001 , n86994 , n86999 , n87000 );
and ( n87002 , n86033 , n86229 );
and ( n87003 , n85936 , n86227 );
nor ( n87004 , n87002 , n87003 );
xnor ( n87005 , n87004 , n86207 );
and ( n87006 , n86413 , n85885 );
not ( n87007 , n87006 );
and ( n87008 , n87007 , n85825 );
and ( n87009 , n87005 , n87008 );
and ( n87010 , n87001 , n87009 );
xor ( n87011 , n86951 , n86955 );
xor ( n87012 , n87011 , n86851 );
and ( n87013 , n87009 , n87012 );
and ( n87014 , n87001 , n87012 );
or ( n87015 , n87010 , n87013 , n87014 );
xor ( n87016 , n86891 , n86895 );
xor ( n87017 , n87016 , n86900 );
and ( n87018 , n87015 , n87017 );
xor ( n87019 , n86947 , n86959 );
xor ( n87020 , n87019 , n86962 );
and ( n87021 , n87017 , n87020 );
and ( n87022 , n87015 , n87020 );
or ( n87023 , n87018 , n87021 , n87022 );
xor ( n87024 , n86965 , n86967 );
xor ( n87025 , n87024 , n86970 );
and ( n87026 , n87023 , n87025 );
and ( n87027 , n86984 , n87026 );
and ( n87028 , n86983 , n87026 );
or ( n87029 , n86985 , n87027 , n87028 );
xor ( n87030 , n86929 , n86930 );
xor ( n87031 , n87030 , n86976 );
and ( n87032 , n87029 , n87031 );
buf ( n87033 , n85660 );
xor ( n87034 , n87005 , n87008 );
and ( n87035 , n85936 , n86403 );
and ( n87036 , n85897 , n86400 );
nor ( n87037 , n87035 , n87036 );
xnor ( n87038 , n87037 , n86204 );
and ( n87039 , n86372 , n85999 );
and ( n87040 , n86288 , n85997 );
nor ( n87041 , n87039 , n87040 );
xnor ( n87042 , n87041 , n85956 );
and ( n87043 , n87038 , n87042 );
and ( n87044 , n87042 , n87006 );
and ( n87045 , n87038 , n87006 );
or ( n87046 , n87043 , n87044 , n87045 );
and ( n87047 , n87034 , n87046 );
and ( n87048 , n86147 , n86125 );
and ( n87049 , n86132 , n86123 );
nor ( n87050 , n87048 , n87049 );
xnor ( n87051 , n87050 , n86070 );
and ( n87052 , n87046 , n87051 );
and ( n87053 , n87034 , n87051 );
or ( n87054 , n87047 , n87052 , n87053 );
xor ( n87055 , n86935 , n86939 );
xor ( n87056 , n87055 , n86944 );
and ( n87057 , n87054 , n87056 );
xor ( n87058 , n87001 , n87009 );
xor ( n87059 , n87058 , n87012 );
and ( n87060 , n87056 , n87059 );
and ( n87061 , n87054 , n87059 );
or ( n87062 , n87057 , n87060 , n87061 );
xor ( n87063 , n87015 , n87017 );
xor ( n87064 , n87063 , n87020 );
and ( n87065 , n87062 , n87064 );
and ( n87066 , n87033 , n87065 );
xor ( n87067 , n87023 , n87025 );
and ( n87068 , n87065 , n87067 );
and ( n87069 , n87033 , n87067 );
or ( n87070 , n87066 , n87068 , n87069 );
xor ( n87071 , n86983 , n86984 );
xor ( n87072 , n87071 , n87026 );
and ( n87073 , n87070 , n87072 );
buf ( n87074 , n85661 );
xor ( n87075 , n87062 , n87064 );
and ( n87076 , n87074 , n87075 );
and ( n87077 , n86033 , n86403 );
and ( n87078 , n85936 , n86400 );
nor ( n87079 , n87077 , n87078 );
xnor ( n87080 , n87079 , n86204 );
and ( n87081 , n86413 , n85997 );
not ( n87082 , n87081 );
and ( n87083 , n87082 , n85956 );
and ( n87084 , n87080 , n87083 );
and ( n87085 , n86132 , n86229 );
and ( n87086 , n86033 , n86227 );
nor ( n87087 , n87085 , n87086 );
xnor ( n87088 , n87087 , n86207 );
and ( n87089 , n87084 , n87088 );
and ( n87090 , n86196 , n86125 );
and ( n87091 , n86147 , n86123 );
nor ( n87092 , n87090 , n87091 );
xnor ( n87093 , n87092 , n86070 );
and ( n87094 , n87088 , n87093 );
and ( n87095 , n87084 , n87093 );
or ( n87096 , n87089 , n87094 , n87095 );
xor ( n87097 , n86989 , n86993 );
xor ( n87098 , n87097 , n86998 );
and ( n87099 , n87096 , n87098 );
xor ( n87100 , n87034 , n87046 );
xor ( n87101 , n87100 , n87051 );
and ( n87102 , n87098 , n87101 );
and ( n87103 , n87096 , n87101 );
or ( n87104 , n87099 , n87102 , n87103 );
xor ( n87105 , n87054 , n87056 );
xor ( n87106 , n87105 , n87059 );
and ( n87107 , n87104 , n87106 );
and ( n87108 , n87075 , n87107 );
and ( n87109 , n87074 , n87107 );
or ( n87110 , n87076 , n87108 , n87109 );
xor ( n87111 , n87033 , n87065 );
xor ( n87112 , n87111 , n87067 );
and ( n87113 , n87110 , n87112 );
buf ( n87114 , n85662 );
xor ( n87115 , n87104 , n87106 );
and ( n87116 , n87114 , n87115 );
and ( n87117 , n86147 , n86229 );
and ( n87118 , n86132 , n86227 );
nor ( n87119 , n87117 , n87118 );
xnor ( n87120 , n87119 , n86207 );
and ( n87121 , n86288 , n86125 );
and ( n87122 , n86196 , n86123 );
nor ( n87123 , n87121 , n87122 );
xnor ( n87124 , n87123 , n86070 );
and ( n87125 , n87120 , n87124 );
and ( n87126 , n86413 , n85999 );
and ( n87127 , n86372 , n85997 );
nor ( n87128 , n87126 , n87127 );
xnor ( n87129 , n87128 , n85956 );
and ( n87130 , n87124 , n87129 );
and ( n87131 , n87120 , n87129 );
or ( n87132 , n87125 , n87130 , n87131 );
xor ( n87133 , n87038 , n87042 );
xor ( n87134 , n87133 , n87006 );
and ( n87135 , n87132 , n87134 );
xor ( n87136 , n87084 , n87088 );
xor ( n87137 , n87136 , n87093 );
and ( n87138 , n87134 , n87137 );
and ( n87139 , n87132 , n87137 );
or ( n87140 , n87135 , n87138 , n87139 );
xor ( n87141 , n87096 , n87098 );
xor ( n87142 , n87141 , n87101 );
and ( n87143 , n87140 , n87142 );
and ( n87144 , n87115 , n87143 );
and ( n87145 , n87114 , n87143 );
or ( n87146 , n87116 , n87144 , n87145 );
xor ( n87147 , n87074 , n87075 );
xor ( n87148 , n87147 , n87107 );
and ( n87149 , n87146 , n87148 );
buf ( n87150 , n85663 );
xor ( n87151 , n87140 , n87142 );
and ( n87152 , n87150 , n87151 );
xor ( n87153 , n87080 , n87083 );
and ( n87154 , n86132 , n86403 );
and ( n87155 , n86033 , n86400 );
nor ( n87156 , n87154 , n87155 );
xnor ( n87157 , n87156 , n86204 );
and ( n87158 , n86196 , n86229 );
and ( n87159 , n86147 , n86227 );
nor ( n87160 , n87158 , n87159 );
xnor ( n87161 , n87160 , n86207 );
and ( n87162 , n87157 , n87161 );
and ( n87163 , n87161 , n87081 );
and ( n87164 , n87157 , n87081 );
or ( n87165 , n87162 , n87163 , n87164 );
and ( n87166 , n87153 , n87165 );
xor ( n87167 , n87120 , n87124 );
xor ( n87168 , n87167 , n87129 );
and ( n87169 , n87165 , n87168 );
and ( n87170 , n87153 , n87168 );
or ( n87171 , n87166 , n87169 , n87170 );
xor ( n87172 , n87132 , n87134 );
xor ( n87173 , n87172 , n87137 );
and ( n87174 , n87171 , n87173 );
and ( n87175 , n87151 , n87174 );
and ( n87176 , n87150 , n87174 );
or ( n87177 , n87152 , n87175 , n87176 );
xor ( n87178 , n87114 , n87115 );
xor ( n87179 , n87178 , n87143 );
and ( n87180 , n87177 , n87179 );
buf ( n87181 , n85664 );
and ( n87182 , n86147 , n86403 );
and ( n87183 , n86132 , n86400 );
nor ( n87184 , n87182 , n87183 );
xnor ( n87185 , n87184 , n86204 );
and ( n87186 , n86413 , n86123 );
not ( n87187 , n87186 );
and ( n87188 , n87187 , n86070 );
and ( n87189 , n87185 , n87188 );
and ( n87190 , n86372 , n86125 );
and ( n87191 , n86288 , n86123 );
nor ( n87192 , n87190 , n87191 );
xnor ( n87193 , n87192 , n86070 );
and ( n87194 , n87189 , n87193 );
xor ( n87195 , n87157 , n87161 );
xor ( n87196 , n87195 , n87081 );
and ( n87197 , n87193 , n87196 );
and ( n87198 , n87189 , n87196 );
or ( n87199 , n87194 , n87197 , n87198 );
xor ( n87200 , n87153 , n87165 );
xor ( n87201 , n87200 , n87168 );
and ( n87202 , n87199 , n87201 );
and ( n87203 , n87181 , n87202 );
xor ( n87204 , n87171 , n87173 );
and ( n87205 , n87202 , n87204 );
and ( n87206 , n87181 , n87204 );
or ( n87207 , n87203 , n87205 , n87206 );
xor ( n87208 , n87150 , n87151 );
xor ( n87209 , n87208 , n87174 );
and ( n87210 , n87207 , n87209 );
buf ( n87211 , n85665 );
xor ( n87212 , n87199 , n87201 );
and ( n87213 , n87211 , n87212 );
xor ( n87214 , n87185 , n87188 );
and ( n87215 , n86288 , n86229 );
and ( n87216 , n86196 , n86227 );
nor ( n87217 , n87215 , n87216 );
xnor ( n87218 , n87217 , n86207 );
and ( n87219 , n87214 , n87218 );
and ( n87220 , n86413 , n86125 );
and ( n87221 , n86372 , n86123 );
nor ( n87222 , n87220 , n87221 );
xnor ( n87223 , n87222 , n86070 );
and ( n87224 , n87218 , n87223 );
and ( n87225 , n87214 , n87223 );
or ( n87226 , n87219 , n87224 , n87225 );
xor ( n87227 , n87189 , n87193 );
xor ( n87228 , n87227 , n87196 );
and ( n87229 , n87226 , n87228 );
and ( n87230 , n87212 , n87229 );
and ( n87231 , n87211 , n87229 );
or ( n87232 , n87213 , n87230 , n87231 );
xor ( n87233 , n87181 , n87202 );
xor ( n87234 , n87233 , n87204 );
and ( n87235 , n87232 , n87234 );
buf ( n87236 , n85666 );
xor ( n87237 , n87226 , n87228 );
and ( n87238 , n87236 , n87237 );
and ( n87239 , n86196 , n86403 );
and ( n87240 , n86147 , n86400 );
nor ( n87241 , n87239 , n87240 );
xnor ( n87242 , n87241 , n86204 );
and ( n87243 , n86372 , n86229 );
and ( n87244 , n86288 , n86227 );
nor ( n87245 , n87243 , n87244 );
xnor ( n87246 , n87245 , n86207 );
and ( n87247 , n87242 , n87246 );
and ( n87248 , n87246 , n87186 );
and ( n87249 , n87242 , n87186 );
or ( n87250 , n87247 , n87248 , n87249 );
xor ( n87251 , n87214 , n87218 );
xor ( n87252 , n87251 , n87223 );
and ( n87253 , n87250 , n87252 );
and ( n87254 , n87237 , n87253 );
and ( n87255 , n87236 , n87253 );
or ( n87256 , n87238 , n87254 , n87255 );
xor ( n87257 , n87211 , n87212 );
xor ( n87258 , n87257 , n87229 );
and ( n87259 , n87256 , n87258 );
buf ( n87260 , n85667 );
buf ( n87261 , n85668 );
xor ( n87262 , n87242 , n87246 );
xor ( n87263 , n87262 , n87186 );
and ( n87264 , n87261 , n87263 );
and ( n87265 , n86288 , n86403 );
and ( n87266 , n86196 , n86400 );
nor ( n87267 , n87265 , n87266 );
xnor ( n87268 , n87267 , n86204 );
and ( n87269 , n86413 , n86227 );
not ( n87270 , n87269 );
and ( n87271 , n87270 , n86207 );
or ( n87272 , n87268 , n87271 );
and ( n87273 , n87263 , n87272 );
and ( n87274 , n87261 , n87272 );
or ( n87275 , n87264 , n87273 , n87274 );
and ( n87276 , n87260 , n87275 );
xor ( n87277 , n87250 , n87252 );
and ( n87278 , n87275 , n87277 );
and ( n87279 , n87260 , n87277 );
or ( n87280 , n87276 , n87278 , n87279 );
xor ( n87281 , n87236 , n87237 );
xor ( n87282 , n87281 , n87253 );
and ( n87283 , n87280 , n87282 );
and ( n87284 , n86413 , n86229 );
and ( n87285 , n86372 , n86227 );
nor ( n87286 , n87284 , n87285 );
xnor ( n87287 , n87286 , n86207 );
xnor ( n87288 , n87268 , n87271 );
or ( n87289 , n87287 , n87288 );
xor ( n87290 , n87261 , n87263 );
xor ( n87291 , n87290 , n87272 );
and ( n87292 , n87289 , n87291 );
and ( n87293 , n86372 , n86403 );
and ( n87294 , n86288 , n86400 );
nor ( n87295 , n87293 , n87294 );
xnor ( n87296 , n87295 , n86204 );
and ( n87297 , n87296 , n87269 );
xnor ( n87298 , n87287 , n87288 );
or ( n87299 , n87297 , n87298 );
and ( n87300 , n87291 , n87299 );
and ( n87301 , n87289 , n87299 );
or ( n87302 , n87292 , n87300 , n87301 );
xor ( n87303 , n87260 , n87275 );
xor ( n87304 , n87303 , n87277 );
or ( n87305 , n87302 , n87304 );
and ( n87306 , n87282 , n87305 );
and ( n87307 , n87280 , n87305 );
or ( n87308 , n87283 , n87306 , n87307 );
and ( n87309 , n87258 , n87308 );
and ( n87310 , n87256 , n87308 );
or ( n87311 , n87259 , n87309 , n87310 );
and ( n87312 , n87234 , n87311 );
and ( n87313 , n87232 , n87311 );
or ( n87314 , n87235 , n87312 , n87313 );
and ( n87315 , n87209 , n87314 );
and ( n87316 , n87207 , n87314 );
or ( n87317 , n87210 , n87315 , n87316 );
and ( n87318 , n87179 , n87317 );
and ( n87319 , n87177 , n87317 );
or ( n87320 , n87180 , n87318 , n87319 );
and ( n87321 , n87148 , n87320 );
and ( n87322 , n87146 , n87320 );
or ( n87323 , n87149 , n87321 , n87322 );
and ( n87324 , n87112 , n87323 );
and ( n87325 , n87110 , n87323 );
or ( n87326 , n87113 , n87324 , n87325 );
and ( n87327 , n87072 , n87326 );
and ( n87328 , n87070 , n87326 );
or ( n87329 , n87073 , n87327 , n87328 );
and ( n87330 , n87031 , n87329 );
and ( n87331 , n87029 , n87329 );
or ( n87332 , n87032 , n87330 , n87331 );
and ( n87333 , n86981 , n87332 );
and ( n87334 , n86979 , n87332 );
or ( n87335 , n86982 , n87333 , n87334 );
and ( n87336 , n86927 , n87335 );
and ( n87337 , n86925 , n87335 );
or ( n87338 , n86928 , n87336 , n87337 );
and ( n87339 , n86886 , n87338 );
and ( n87340 , n86884 , n87338 );
or ( n87341 , n86887 , n87339 , n87340 );
and ( n87342 , n86826 , n87341 );
and ( n87343 , n86824 , n87341 );
or ( n87344 , n86827 , n87342 , n87343 );
and ( n87345 , n86765 , n87344 );
and ( n87346 , n86763 , n87344 );
or ( n87347 , n86766 , n87345 , n87346 );
and ( n87348 , n86681 , n87347 );
and ( n87349 , n86679 , n87347 );
or ( n87350 , n86682 , n87348 , n87349 );
and ( n87351 , n86610 , n87350 );
and ( n87352 , n86608 , n87350 );
or ( n87353 , n86611 , n87351 , n87352 );
and ( n87354 , n86572 , n87353 );
and ( n87355 , n86570 , n87353 );
or ( n87356 , n86573 , n87354 , n87355 );
and ( n87357 , n86481 , n87356 );
and ( n87358 , n86479 , n87356 );
or ( n87359 , n86482 , n87357 , n87358 );
and ( n87360 , n86338 , n87359 );
and ( n87361 , n86336 , n87359 );
or ( n87362 , n86339 , n87360 , n87361 );
and ( n87363 , n86273 , n87362 );
and ( n87364 , n86182 , n87362 );
or ( n87365 , n86274 , n87363 , n87364 );
and ( n87366 , n86179 , n87365 );
and ( n87367 , n86177 , n87365 );
or ( n87368 , n86180 , n87366 , n87367 );
and ( n87369 , n86059 , n87368 );
and ( n87370 , n86057 , n87368 );
or ( n87371 , n86060 , n87369 , n87370 );
and ( n87372 , n85991 , n87371 );
and ( n87373 , n85989 , n87371 );
or ( n87374 , n85992 , n87372 , n87373 );
and ( n87375 , n85921 , n87374 );
and ( n87376 , n85864 , n87374 );
or ( n87377 , n85922 , n87375 , n87376 );
and ( n87378 , n85861 , n87377 );
and ( n87379 , n85859 , n87377 );
or ( n87380 , n85862 , n87378 , n87379 );
xor ( n87381 , n85815 , n87380 );
not ( n87382 , n87381 );
xor ( n87383 , n85859 , n85861 );
xor ( n87384 , n87383 , n87377 );
not ( n87385 , n87384 );
xor ( n87386 , n85864 , n85921 );
xor ( n87387 , n87386 , n87374 );
not ( n87388 , n87387 );
xor ( n87389 , n85989 , n85991 );
xor ( n87390 , n87389 , n87371 );
not ( n87391 , n87390 );
xor ( n87392 , n86057 , n86059 );
xor ( n87393 , n87392 , n87368 );
not ( n87394 , n87393 );
xor ( n87395 , n86177 , n86179 );
xor ( n87396 , n87395 , n87365 );
not ( n87397 , n87396 );
xor ( n87398 , n86182 , n86273 );
xor ( n87399 , n87398 , n87362 );
not ( n87400 , n87399 );
xor ( n87401 , n86336 , n86338 );
xor ( n87402 , n87401 , n87359 );
not ( n87403 , n87402 );
xor ( n87404 , n86479 , n86481 );
xor ( n87405 , n87404 , n87356 );
not ( n87406 , n87405 );
xor ( n87407 , n86570 , n86572 );
xor ( n87408 , n87407 , n87353 );
not ( n87409 , n87408 );
xor ( n87410 , n86608 , n86610 );
xor ( n87411 , n87410 , n87350 );
not ( n87412 , n87411 );
xor ( n87413 , n86679 , n86681 );
xor ( n87414 , n87413 , n87347 );
not ( n87415 , n87414 );
xor ( n87416 , n86763 , n86765 );
xor ( n87417 , n87416 , n87344 );
not ( n87418 , n87417 );
xor ( n87419 , n86824 , n86826 );
xor ( n87420 , n87419 , n87341 );
not ( n87421 , n87420 );
xor ( n87422 , n86884 , n86886 );
xor ( n87423 , n87422 , n87338 );
not ( n87424 , n87423 );
xor ( n87425 , n86925 , n86927 );
xor ( n87426 , n87425 , n87335 );
not ( n87427 , n87426 );
xor ( n87428 , n86979 , n86981 );
xor ( n87429 , n87428 , n87332 );
not ( n87430 , n87429 );
xor ( n87431 , n87029 , n87031 );
xor ( n87432 , n87431 , n87329 );
not ( n87433 , n87432 );
xor ( n87434 , n87070 , n87072 );
xor ( n87435 , n87434 , n87326 );
not ( n87436 , n87435 );
xor ( n87437 , n87110 , n87112 );
xor ( n87438 , n87437 , n87323 );
not ( n87439 , n87438 );
xor ( n87440 , n87146 , n87148 );
xor ( n87441 , n87440 , n87320 );
not ( n87442 , n87441 );
xor ( n87443 , n87177 , n87179 );
xor ( n87444 , n87443 , n87317 );
not ( n87445 , n87444 );
xor ( n87446 , n87207 , n87209 );
xor ( n87447 , n87446 , n87314 );
not ( n87448 , n87447 );
xor ( n87449 , n87232 , n87234 );
xor ( n87450 , n87449 , n87311 );
not ( n87451 , n87450 );
xor ( n87452 , n87256 , n87258 );
xor ( n87453 , n87452 , n87308 );
not ( n87454 , n87453 );
xor ( n87455 , n87280 , n87282 );
xor ( n87456 , n87455 , n87305 );
not ( n87457 , n87456 );
xnor ( n87458 , n87302 , n87304 );
xor ( n87459 , n87289 , n87291 );
xor ( n87460 , n87459 , n87299 );
not ( n87461 , n87460 );
xnor ( n87462 , n87297 , n87298 );
and ( n87463 , n86413 , n86403 );
and ( n87464 , n86372 , n86400 );
nor ( n87465 , n87463 , n87464 );
xnor ( n87466 , n87465 , n86204 );
and ( n87467 , n86413 , n86400 );
not ( n87468 , n87467 );
and ( n87469 , n87468 , n86204 );
or ( n87470 , n87466 , n87469 );
xor ( n87471 , n87296 , n87269 );
and ( n87472 , n87470 , n87471 );
and ( n87473 , n87462 , n87472 );
and ( n87474 , n87461 , n87473 );
or ( n87475 , n87460 , n87474 );
and ( n87476 , n87458 , n87475 );
and ( n87477 , n87457 , n87476 );
or ( n87478 , n87456 , n87477 );
and ( n87479 , n87454 , n87478 );
or ( n87480 , n87453 , n87479 );
and ( n87481 , n87451 , n87480 );
or ( n87482 , n87450 , n87481 );
and ( n87483 , n87448 , n87482 );
or ( n87484 , n87447 , n87483 );
and ( n87485 , n87445 , n87484 );
or ( n87486 , n87444 , n87485 );
and ( n87487 , n87442 , n87486 );
or ( n87488 , n87441 , n87487 );
and ( n87489 , n87439 , n87488 );
or ( n87490 , n87438 , n87489 );
and ( n87491 , n87436 , n87490 );
or ( n87492 , n87435 , n87491 );
and ( n87493 , n87433 , n87492 );
or ( n87494 , n87432 , n87493 );
and ( n87495 , n87430 , n87494 );
or ( n87496 , n87429 , n87495 );
and ( n87497 , n87427 , n87496 );
or ( n87498 , n87426 , n87497 );
and ( n87499 , n87424 , n87498 );
or ( n87500 , n87423 , n87499 );
and ( n87501 , n87421 , n87500 );
or ( n87502 , n87420 , n87501 );
and ( n87503 , n87418 , n87502 );
or ( n87504 , n87417 , n87503 );
and ( n87505 , n87415 , n87504 );
or ( n87506 , n87414 , n87505 );
and ( n87507 , n87412 , n87506 );
or ( n87508 , n87411 , n87507 );
and ( n87509 , n87409 , n87508 );
or ( n87510 , n87408 , n87509 );
and ( n87511 , n87406 , n87510 );
or ( n87512 , n87405 , n87511 );
and ( n87513 , n87403 , n87512 );
or ( n87514 , n87402 , n87513 );
and ( n87515 , n87400 , n87514 );
or ( n87516 , n87399 , n87515 );
and ( n87517 , n87397 , n87516 );
or ( n87518 , n87396 , n87517 );
and ( n87519 , n87394 , n87518 );
or ( n87520 , n87393 , n87519 );
and ( n87521 , n87391 , n87520 );
or ( n87522 , n87390 , n87521 );
and ( n87523 , n87388 , n87522 );
or ( n87524 , n87387 , n87523 );
and ( n87525 , n87385 , n87524 );
or ( n87526 , n87384 , n87525 );
xor ( n87527 , n87382 , n87526 );
buf ( n87528 , n87527 );
xor ( n87529 , n87385 , n87524 );
buf ( n87530 , n87529 );
xor ( n87531 , n87388 , n87522 );
buf ( n87532 , n87531 );
xor ( n87533 , n87391 , n87520 );
buf ( n87534 , n87533 );
xor ( n87535 , n87394 , n87518 );
buf ( n87536 , n87535 );
xor ( n87537 , n87397 , n87516 );
buf ( n87538 , n87537 );
xor ( n87539 , n87400 , n87514 );
buf ( n87540 , n87539 );
xor ( n87541 , n87403 , n87512 );
buf ( n87542 , n87541 );
xor ( n87543 , n87406 , n87510 );
buf ( n87544 , n87543 );
xor ( n87545 , n87409 , n87508 );
buf ( n87546 , n87545 );
xor ( n87547 , n87412 , n87506 );
buf ( n87548 , n87547 );
xor ( n87549 , n87415 , n87504 );
buf ( n87550 , n87549 );
xor ( n87551 , n87418 , n87502 );
buf ( n87552 , n87551 );
xor ( n87553 , n87421 , n87500 );
buf ( n87554 , n87553 );
xor ( n87555 , n87424 , n87498 );
buf ( n87556 , n87555 );
xor ( n87557 , n87427 , n87496 );
buf ( n87558 , n87557 );
xor ( n87559 , n87430 , n87494 );
buf ( n87560 , n87559 );
xor ( n87561 , n87433 , n87492 );
buf ( n87562 , n87561 );
xor ( n87563 , n87436 , n87490 );
buf ( n87564 , n87563 );
xor ( n87565 , n87439 , n87488 );
buf ( n87566 , n87565 );
xor ( n87567 , n87442 , n87486 );
buf ( n87568 , n87567 );
xor ( n87569 , n87445 , n87484 );
buf ( n87570 , n87569 );
xor ( n87571 , n87448 , n87482 );
buf ( n87572 , n87571 );
xor ( n87573 , n87451 , n87480 );
buf ( n87574 , n87573 );
xor ( n87575 , n87454 , n87478 );
buf ( n87576 , n87575 );
xor ( n87577 , n87457 , n87476 );
buf ( n87578 , n87577 );
xor ( n87579 , n87458 , n87475 );
buf ( n87580 , n87579 );
xor ( n87581 , n87461 , n87473 );
buf ( n87582 , n87581 );
xor ( n87583 , n87462 , n87472 );
buf ( n87584 , n87583 );
xor ( n87585 , n87470 , n87471 );
buf ( n87586 , n87585 );
xnor ( n87587 , n87466 , n87469 );
buf ( n87588 , n87587 );
buf ( n87589 , n87467 );
buf ( n87590 , n87589 );
endmodule
