module DMDbuf (I, O);

input [15:0] I;
output [15:0] O;

assign O = I;
endmodule
