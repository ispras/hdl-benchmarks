//NOTE: no-implementation module stub

module REG14L (
    input wire DSPCLK,
    input wire RST,
    input wire CLKI4enb,
    input wire ldI,
    input wire [13:0] Iin,
    output wire [13:0] I4,
    input wire SCAN_TEST
);

endmodule
