// IWLS benchmark module "vda" printed on Wed May 29 17:30:25 2002
module vda(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q;
output
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  a1,
  b0,
  b1,
  c0,
  c1,
  d0,
  d1,
  e0,
  f0,
  g0,
  h0,
  i0,
  j0,
  k0,
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0,
  t0,
  u0,
  v0,
  w0,
  x0,
  y0,
  z0;
wire
  \[15] ,
  \[16] ,
  \[17] ,
  \[18] ,
  \[19] ,
  \[0] ,
  \[1] ,
  \[20] ,
  \[2] ,
  \[21] ,
  \[3] ,
  \[22] ,
  \[4] ,
  \[23] ,
  \[5] ,
  \[24] ,
  \[6] ,
  \[25] ,
  \[7] ,
  \[26] ,
  \[8] ,
  \[27] ,
  \[9] ,
  \[28] ,
  \[29] ,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  a5,
  a6,
  a7,
  \[35] ,
  b5,
  b6,
  b7,
  \[36] ,
  c5,
  c6,
  c7,
  \[37] ,
  d5,
  d6,
  d7,
  \[38] ,
  e4,
  e5,
  e6,
  e7,
  f4,
  f5,
  f6,
  f7,
  g4,
  g5,
  g6,
  g7,
  h4,
  h5,
  h6,
  h7,
  i4,
  i5,
  i6,
  i7,
  j4,
  j5,
  j6,
  j7,
  k4,
  k5,
  k6,
  l4,
  l5,
  l6,
  m4,
  m5,
  m6,
  n4,
  n5,
  n6,
  o4,
  o5,
  o6,
  p4,
  p5,
  p6,
  q4,
  q5,
  q6,
  r4,
  r5,
  r6,
  s4,
  s5,
  s6,
  t4,
  t5,
  t6,
  u4,
  u5,
  u6,
  v4,
  v5,
  v6,
  w4,
  w5,
  w6,
  x4,
  x5,
  x6,
  y4,
  y5,
  y6,
  z4,
  z5,
  z6,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[14] ;
assign
  \[15]  = p5 | (q5 | (r5 | (t5 | (u5 | (v5 | (n4 | (a6 | (c6 | (d6 | (g6 | (k6 | (m6 | (n6 | (s6 | (\[35]  | (e6 | (l4 | (f4 | (g4 | (i4 | (j4 | (k4 | (o5 | (m4 | (p4 | (r4 | (s4 | (t4 | (u4 | (w4 | (y4 | (a5 | (c5 | (e5 | (f5 | (g5 | (h5 | (m5 | (b7 | (l5 | (q6 | (j7 | (g7 | (f7 | (d7 | (x6 | (e7 | (v6 | (e4 | z6))))))))))))))))))))))))))))))))))))))))))))))))),
  \[16]  = (q & (p & (o & (n & (~l & (~i & (~g & ~c))))))) | (p5 | (r5 | (s5 | (t5 | (v5 | (w5 | (n4 | (d6 | (j5 | (h6 | (k6 | (l6 | (m6 | (n6 | (\[11]  | (y5 | (s6 | (t6 | (\[38]  | (w6 | (e6 | (l4 | (f4 | (g4 | (h4 | (i4 | (p4 | (q4 | (r4 | (w4 | (x4 | (\[34]  | (y4 | (z4 | (h7 | (\[36]  | (x6 | (e7 | (v6 | (p6 | (a7 | z6))))))))))))))))))))))))))))))))))))))))),
  \[17]  = (~p & (~o & (~n & (~m & (~l & ~c))))) | (p5 | (r5 | (s5 | (u5 | (v5 | (w5 | (n4 | (z5 | (c6 | (d6 | (j5 | (g6 | (h6 | (j6 | (l6 | (y5 | (t6 | (u6 | (w6 | (i4 | (j4 | (m4 | (p4 | (r4 | (v4 | (w4 | (b5 | (d5 | (i5 | (i7 | (c7 | (y6 | (p6 | (a7 | o6)))))))))))))))))))))))))))))))))),
  \[18]  = k4 | (u4 | (d5 | (h5 | (b7 | (g7 | (f7 | (d7 | e4))))))),
  \[19]  = p5 | (q5 | (r5 | (s5 | (t5 | (u5 | (v5 | (w5 | (x5 | (z5 | (a6 | (b6 | (o4 | (f6 | (g6 | (i6 | (n5 | (s6 | (\[38]  | (k4 | (q4 | (u4 | (d5 | (h5 | (b7 | (\[36]  | (g7 | (f7 | (d7 | e4)))))))))))))))))))))))))))),
  r = \[0] ,
  s = \[1] ,
  t = \[2] ,
  u = \[3] ,
  v = \[4] ,
  w = \[5] ,
  \x  = \[6] ,
  y = \[7] ,
  z = \[8] ,
  \[0]  = p5 | (q5 | (r5 | (s5 | (t5 | (u5 | (v5 | (w5 | (x5 | (n4 | (z5 | (a6 | (b6 | (c6 | (d6 | (o4 | (f6 | (g6 | (h6 | (i6 | (j6 | (l6 | (m6 | (n6 | (n5 | (t6 | (h4 | (s4 | (t4 | (a5 | (i7 | (c7 | y6))))))))))))))))))))))))))))))),
  \[1]  = \[35]  | (k4 | (d5 | (h5 | (b7 | (j7 | (g7 | (f7 | (d7 | e4)))))))),
  \[20]  = p5 | (q5 | (r5 | (s5 | (t5 | (u5 | (v5 | (x5 | (n4 | (z5 | (a6 | (b6 | (c6 | (d6 | (f6 | (i6 | (j6 | (l6 | (n6 | (\[11]  | (t6 | (\[35]  | (\[38]  | (h4 | (\[10]  | (\[34]  | \[36] ))))))))))))))))))))))))),
  \[2]  = p5 | (q5 | (r5 | (s5 | (t5 | (u5 | (v5 | (w5 | (x5 | (n4 | (z5 | (a6 | (b6 | (c6 | (d6 | (o4 | (g6 | (h6 | (l6 | (m6 | (h4 | (s4 | (t4 | (a5 | (i7 | (c7 | y6))))))))))))))))))))))))),
  \[21]  = p5 | (r5 | (t5 | (v5 | (w5 | (z5 | (b6 | (c6 | (d6 | (o4 | (g6 | (l6 | (m6 | (n5 | (s6 | (h4 | (q4 | (s4 | (t4 | a5)))))))))))))))))),
  \[3]  = j5 | (k6 | (\[11]  | (k5 | (r6 | u6)))),
  \[22]  = p5 | (q5 | (r5 | (s5 | (t5 | (u5 | (v5 | (w5 | (x5 | (n4 | (z5 | (a6 | (b6 | (o4 | (f6 | (g6 | (i6 | (j6 | (n6 | (\[11]  | (n5 | (s6 | (t6 | (\[35]  | (\[38]  | (\[10]  | (q4 | (\[34]  | \[36] ))))))))))))))))))))))))))),
  \[4]  = j5 | (f6 | (i6 | (j6 | (k6 | (\[11]  | (k5 | (n5 | (r6 | (u6 | (e6 | (l4 | (f4 | (g4 | (\[10]  | m4)))))))))))))),
  \[23]  = q5 | (x5 | (n4 | (a6 | (c6 | (f6 | (i6 | (j6 | (h4 | (\[10]  | (k4 | (s4 | (t4 | (u4 | (\[34]  | (a5 | (d5 | (h5 | (b7 | (\[36]  | (g7 | (f7 | (d7 | (i7 | (c7 | (y6 | e4))))))))))))))))))))))))),
  \[5]  = p5 | (q5 | (r5 | (s5 | (t5 | (u5 | (v5 | (w5 | (x5 | (n4 | (z5 | (a6 | (b6 | (c6 | (d6 | (o4 | (g6 | (h6 | (l6 | (m6 | (h4 | (s4 | (t4 | (a5 | (i7 | (c7 | y6))))))))))))))))))))))))),
  \[24]  = p5 | (q5 | (r5 | (s5 | (t5 | (u5 | (v5 | (w5 | (x5 | (z5 | (a6 | (b6 | (o4 | (j5 | (f6 | (g6 | (i6 | (k5 | (n5 | (r6 | (u6 | (e6 | (l4 | (f4 | (g4 | m4)))))))))))))))))))))))),
  \[6]  = p5 | (q5 | (r5 | (s5 | (t5 | (u5 | (v5 | (w5 | (x5 | (n4 | (z5 | (a6 | (b6 | (c6 | (d6 | (o4 | (g6 | (h6 | (l6 | (m6 | (h4 | (s4 | (t4 | (a5 | (i7 | (c7 | y6))))))))))))))))))))))))),
  \[25]  = p5 | (q5 | (r5 | (s5 | (t5 | (u5 | (v5 | (x5 | (z5 | (a6 | (b6 | (c6 | (d6 | (j5 | (f6 | (g6 | (h6 | (i6 | (j6 | (k6 | (n6 | (\[11]  | (k5 | (t6 | (u6 | (e6 | (l4 | (f4 | (g4 | (\[10]  | (m4 | (i7 | (c7 | y6)))))))))))))))))))))))))))))))),
  \[7]  = j5 | (f6 | (i6 | (k6 | (\[11]  | (k5 | (n5 | (r6 | (u6 | (e6 | (l4 | (f4 | (g4 | (\[10]  | m4))))))))))))),
  \[26]  = p5 | (r5 | (v5 | (w5 | (x5 | (b6 | (c6 | (d6 | (o4 | (j6 | (k6 | (m6 | (n6 | (\[11]  | (k5 | (n5 | (r6 | (t6 | (u6 | (\[10]  | (m4 | (s4 | (t4 | a5)))))))))))))))))))))),
  \[8]  = c6 | d6,
  \[27]  = p5 | (q5 | (r5 | (s5 | (t5 | (u5 | (v5 | (w5 | (x5 | (z5 | (a6 | (b6 | (o4 | (j5 | (f6 | (g6 | (h6 | (i6 | (k5 | (n5 | (r6 | (u6 | (e6 | (l4 | (f4 | (g4 | (m4 | (i7 | (c7 | y6)))))))))))))))))))))))))))),
  \[9]  = f6 | (i6 | (\[11]  | \[10] )),
  \[28]  = q5 | (t5 | (n4 | (z5 | (a6 | (c6 | (j5 | (f6 | (i6 | (j6 | (k6 | (e6 | (l4 | (f4 | (g4 | (h4 | (\[10]  | (s4 | (t4 | (a5 | (i7 | (c7 | y6))))))))))))))))))))),
  \[29]  = p5 | (q5 | (r5 | (s5 | (t5 | (u5 | (v5 | (w5 | (x5 | (n4 | (z5 | (a6 | (b6 | (o4 | (f6 | (g6 | (h6 | (i6 | (l6 | (n5 | (r6 | (h4 | (i7 | (c7 | y6))))))))))))))))))))))),
  \[30]  = r5 | (s5 | (t5 | (u5 | (v5 | (w5 | (c6 | (d6 | (o4 | (j5 | (f6 | (g6 | (i6 | (k6 | (k5 | (u6 | (e6 | (l4 | (f4 | (g4 | m4))))))))))))))))))),
  \[31]  = p5 | (q5 | (a6 | (b6 | (k6 | (m6 | (s4 | (t4 | a5))))))),
  \[32]  = p5 | (q5 | (a6 | (b6 | (j5 | (m6 | (k5 | (r6 | (u6 | (e6 | (l4 | (f4 | (g4 | (m4 | (s4 | (t4 | a5))))))))))))))),
  \[33]  = p5 | (q5 | (s5 | (u5 | (w5 | (a6 | (b6 | (c6 | (o4 | (j5 | (g6 | (n6 | (\[11]  | (k5 | (t6 | (u6 | (e6 | (l4 | (f4 | (g4 | (m4 | (s4 | (t4 | a5)))))))))))))))))))))),
  \[34]  = q & (~p & (~o & (~n & (~m & l)))),
  a0 = \[9] ,
  a1 = \[35] ,
  a5 = ~q & (~p & (o & (~n & (~m & (l & (e & a)))))),
  a6 = q & (p & (~o & (n & (~m & (~l & i))))),
  a7 = q & (p & (~o & (~n & (~m & (~l & (f & (~e & b))))))),
  \[35]  = q & (p & (~o & (~n & (~m & l)))),
  b0 = \[10] ,
  b1 = \[36] ,
  b5 = ~q & (~p & (~o & (n & (m & ~l)))),
  b6 = ~q & (~p & (o & (n & (~m & ~l)))),
  b7 = ~q & (o & (n & (m & (~l & (~i & ~h))))),
  \[36]  = ~q & (~p & (o & (n & (m & (~l & (j & h)))))),
  c0 = \[11] ,
  c1 = \[37] ,
  c5 = ~q & (p & (~o & (n & (m & ~l)))),
  c6 = ~q & (~p & (o & (~n & (~m & ~l)))),
  c7 = ~q & (p & (o & (n & (m & (~l & (j & (~i & (h & (e & ~c))))))))),
  \[37]  = s6 | q4,
  d0 = \[12] ,
  d1 = \[38] ,
  d5 = ~q & (~p & (~o & (~n & (~m & ~l)))),
  d6 = ~q & (p & (o & (~n & (~m & ~l)))),
  d7 = ~q & (p & (o & (n & (m & (~l & (~i & (~e & b))))))),
  \[38]  = q & (~p & (~o & (n & (m & l)))),
  e0 = \[13] ,
  e4 = ~q & (~p & (o & (~n & (~m & (l & (~f & (~e & a))))))),
  e5 = q & (p & (o & (n & (~l & ~g)))),
  e6 = ~q & (p & (o & (~n & (m & (~l & (g & c)))))),
  e7 = p & (o & (n & (m & (~l & (~j & (h & (e & ~c))))))),
  f0 = \[14] ,
  f4 = ~q & (p & (o & (~n & (m & (~l & (k & g)))))),
  f5 = q & (p & (n & (m & (~l & g)))),
  f6 = q & (p & (o & (n & (~m & (~l & g))))),
  f7 = ~q & (p & (o & (n & (m & (~l & (~i & (~e & ~c))))))),
  g0 = \[15] ,
  g4 = q & (p & (~o & (n & (~m & (~l & (~i & d)))))),
  g5 = q & (~p & (n & (~m & l))),
  g6 = q & (p & (~o & (~n & (~m & (~l & (f & ~b)))))),
  g7 = ~q & (p & (o & (n & (m & (~l & (~i & (~f & ~e))))))),
  h0 = \[16] ,
  h4 = q & (~p & (~o & (~n & (~m & (~l & c))))),
  h5 = ~q & (~p & (o & (n & (m & (~l & ~h))))),
  h6 = ~q & (p & (~o & (~n & (~m & l)))),
  h7 = q & (p & (o & (~n & (~m & (~l & k))))),
  i0 = \[17] ,
  i4 = p & (o & (~n & (m & l))),
  i5 = ~q & (~p & (~o & (n & (~m & l)))),
  i6 = ~q & (~p & (o & (~n & (m & (~l & g))))),
  i7 = ~q & (p & (o & (n & (m & (~l & (j & (~i & (h & (~f & e))))))))),
  j0 = \[18] ,
  j4 = q & (p & (~o & (~n & (m & ~l)))),
  j5 = ~q & (p & (~o & (~n & (m & ~l)))),
  j6 = ~q & (~p & (~o & (n & (~m & ~l)))),
  j7 = q & (p & (~o & (~n & (~m & (~f & ~e))))),
  k0 = \[19] ,
  k4 = ~q & (p & (o & (n & (~m & l)))),
  k5 = q & (~p & (~o & (n & (m & ~l)))),
  k6 = q & (~p & (o & (~n & (m & l)))),
  l0 = \[20] ,
  l4 = ~q & (p & (o & (~n & (m & (~l & (i & g)))))),
  l5 = ~q & (~p & (o & (n & (m & (~l & h))))),
  l6 = ~q & (p & (~o & (~n & (~m & ~l)))),
  m0 = \[21] ,
  m4 = q & (p & (~o & (n & (~m & (~l & (~i & ~d)))))),
  m5 = ~p & (o & (~n & (l & ~a))),
  m6 = q & (~p & (o & (~n & (~m & ~l)))),
  n0 = \[22] ,
  n4 = ~q & (p & (o & (~n & (~m & l)))),
  n5 = q & (p & (o & (~n & (~m & (l & g))))),
  n6 = ~q & (p & (~o & (n & (~m & (~l & ~f))))),
  o0 = \[23] ,
  o4 = q & (p & (o & (~n & (~m & (l & ~g))))),
  o5 = ~q & (p & (~n & (m & l))),
  o6 = ~q & (p & (o & (n & (m & (~l & (~i & (h & (f & (c & ~b))))))))),
  p0 = \[24] ,
  p4 = q & (p & (~o & (n & (~m & l)))),
  p5 = ~q & (~p & (o & (~n & (m & l)))),
  p6 = ~q & (o & (~n & (~m & (l & (f & (~e & a)))))),
  q0 = \[25] ,
  q4 = q & (p & (o & (n & (m & ~l)))),
  q5 = q & (p & (~o & (~n & (m & l)))),
  q6 = ~q & (~p & (o & (~n & (m & (~l & ~g))))),
  r0 = \[26] ,
  r4 = ~q & (p & (o & (n & (m & (~l & i))))),
  r5 = ~q & (p & (o & (~n & (m & (~l & ~g))))),
  r6 = q & (p & (o & (n & (~m & l)))),
  s0 = \[27] ,
  s4 = q & (p & (~o & (~n & (~m & (~l & (~f & e)))))),
  s5 = ~q & (~p & (~o & (n & (m & l)))),
  s6 = ~q & (~p & (~o & (~n & (~m & l)))),
  t0 = \[28] ,
  t4 = q & (p & (~o & (~n & (~m & (~l & (e & b)))))),
  t5 = q & (~p & (o & (~n & (~m & l)))),
  t6 = ~q & (p & (~o & (n & (~m & (~l & f))))),
  u0 = \[29] ,
  u4 = ~q & (~p & (o & (n & (m & l)))),
  u5 = q & (p & (~o & (n & (m & l)))),
  u6 = q & (~p & (~o & (n & (~m & l)))),
  v0 = \[30] ,
  v4 = ~q & (~o & (~n & (m & l))),
  v5 = q & (p & (~o & (n & (m & (~l & ~g))))),
  v6 = p & (o & (n & (m & (~l & (~j & (h & (e & b))))))),
  w0 = \[31] ,
  w4 = q & (~p & (~o & (~n & (m & l)))),
  w5 = q & (~p & (o & (n & (~m & ~l)))),
  w6 = ~q & (~p & (o & (n & ~m))),
  x0 = \[32] ,
  x4 = q & (~p & (o & (~n & (m & ~l)))),
  x5 = q & (p & (o & (~n & (m & ~l)))),
  x6 = p & (o & (n & (m & (~l & (~j & (h & (~f & e))))))),
  y0 = \[33] ,
  y4 = ~q & (p & (~o & (n & (~m & l)))),
  y5 = ~q & (o & (n & (~m & ~l))),
  y6 = ~q & (p & (o & (n & (m & (~l & (j & (~i & (h & (e & b))))))))),
  z0 = \[34] ,
  z4 = q & (~p & (~o & (m & ~l))),
  z5 = ~q & (~p & (~o & (~n & (m & ~l)))),
  z6 = ~q & (p & (o & (~n & (m & (~l & (~k & (~i & (g & ~c)))))))),
  \[10]  = q & (p & (o & (~n & (~m & (~l & ~k))))),
  \[11]  = q & (~p & (~o & (n & (~m & ~l)))),
  \[12]  = (~q & (p & (~o & (n & m)))) | (p5 | (q5 | (s5 | (t5 | (n4 | (o4 | (g6 | (h6 | (k6 | (n5 | (y5 | (r6 | (s6 | (\[35]  | (\[38]  | (j4 | (k4 | (o5 | (u4 | (v4 | (w4 | (x4 | (\[34]  | (h5 | (i5 | (m5 | (b7 | (h7 | (j7 | (g7 | (f7 | (d7 | (i7 | (c7 | (y6 | (e4 | o6)))))))))))))))))))))))))))))))))))),
  \[13]  = q5 | (r5 | (s5 | (v5 | (x5 | (z5 | (o4 | (j5 | (f6 | (i6 | (k6 | (n6 | (r6 | (\[35]  | (\[38]  | (w6 | (o5 | (m4 | (r4 | (v4 | (y4 | (z4 | (b5 | (e5 | (f5 | (g5 | (l5 | (q6 | (h7 | (x6 | (e7 | (v6 | (z6 | o6)))))))))))))))))))))))))))))))),
  \[14]  = p5 | (u5 | (w5 | (x5 | (n4 | (a6 | (o4 | (j6 | (n6 | (\[11]  | (k5 | (n5 | (y5 | (s6 | (t6 | (\[35]  | (\[38]  | (w6 | (e6 | (l4 | (f4 | (g4 | (j4 | (\[10]  | (p4 | (r4 | (x4 | (b5 | (c5 | (e5 | (f5 | (i5 | (l5 | (q6 | (x6 | (e7 | (v6 | (p6 | (a7 | (z6 | o6)))))))))))))))))))))))))))))))))))))));
endmodule

