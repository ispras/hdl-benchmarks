//NOTE: no-implementation module stub

module BTBmem (
    input DSPCLK,
    input [4:0] BTB_wa,
    input BTB_web,
    input PWRDn,
    input [25:0] BTB_wd,
    input [4:0] BTB_ra,
    output [25:0] BTB_rd
);

endmodule
