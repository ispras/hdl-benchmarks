// IWLS benchmark module "i9" printed on Wed May 29 17:27:06 2002
module i9(\V9(3) , \V9(1) , \V9(2) , \V9(10) , \V9(0) , \V9(5) , \V9(6) , \V9(7) , \V9(8) , \V56(31) , \V56(30) , \V56(29) , \V56(28) , \V56(27) , \V56(26) , \V56(25) , \V56(24) , \V56(23) , \V56(22) , \V56(21) , \V56(20) , \V56(19) , \V56(18) , \V56(17) , \V56(16) , \V56(15) , \V56(14) , \V56(13) , \V56(12) , \V56(11) , \V56(10) , \V56(9) , \V56(8) , \V56(7) , \V56(6) , \V56(5) , \V56(4) , \V56(3) , \V56(2) , \V56(1) , \V56(0) , \V88(11) , \V88(10) , \V88(9) , \V88(8) , \V88(7) , \V88(6) , \V88(5) , \V88(4) , \V88(3) , \V88(2) , \V88(1) , \V24(14) , \V24(13) , \V24(12) , \V24(11) , \V24(10) , \V24(9) , \V24(8) , \V24(7) , \V24(6) , \V24(5) , \V24(4) , \V24(3) , \V24(2) , \V24(1) , \V24(0) , \V88(31) , \V88(30) , \V88(29) , \V88(28) , \V88(27) , \V88(26) , \V88(25) , \V88(24) , \V88(23) , \V88(22) , \V88(21) , \V88(20) , \V88(19) , \V88(18) , \V88(17) , \V88(16) , \V88(15) , \V88(14) , \V88(13) , \V88(12) , \V88(0) , \V119(30) , \V119(29) , \V119(28) , \V119(27) , \V119(26) , \V119(25) , \V119(24) , \V119(23) , \V119(22) , \V119(21) , \V119(20) , \V119(19) , \V119(18) , \V119(17) , \V119(16) , \V119(15) , \V119(14) , \V119(13) , \V119(12) , \V119(11) , \V119(10) , \V119(9) , \V119(8) , \V119(7) , \V119(6) , \V119(5) , \V119(4) , \V119(3) , \V119(2) , \V119(1) , \V119(0) , \V151(15) , \V151(14) , \V151(13) , \V151(12) , \V151(11) , \V151(10) , \V151(9) , \V151(8) , \V151(7) , \V151(6) , \V151(5) , \V151(4) , \V151(3) , \V151(2) , \V151(1) , \V151(0) , \V151(31) , \V151(30) , \V151(29) , \V151(28) , \V151(27) , \V151(26) , \V151(25) , \V151(24) , \V151(23) , \V151(22) , \V151(21) , \V151(20) , \V151(19) , \V151(18) , \V151(17) , \V151(16) );
input
  \V9(10) ,
  \V56(0) ,
  \V56(1) ,
  \V56(2) ,
  \V56(3) ,
  \V56(4) ,
  \V56(5) ,
  \V56(6) ,
  \V56(7) ,
  \V56(8) ,
  \V56(9) ,
  \V24(13) ,
  \V24(12) ,
  \V24(14) ,
  \V24(11) ,
  \V24(10) ,
  \V9(0) ,
  \V9(1) ,
  \V9(2) ,
  \V9(3) ,
  \V9(5) ,
  \V9(6) ,
  \V9(7) ,
  \V9(8) ,
  \V88(13) ,
  \V88(12) ,
  \V88(15) ,
  \V88(14) ,
  \V88(11) ,
  \V88(10) ,
  \V88(0) ,
  \V88(1) ,
  \V88(2) ,
  \V88(3) ,
  \V88(17) ,
  \V88(4) ,
  \V88(16) ,
  \V88(5) ,
  \V88(19) ,
  \V88(6) ,
  \V88(18) ,
  \V88(7) ,
  \V88(23) ,
  \V88(8) ,
  \V88(22) ,
  \V88(9) ,
  \V88(25) ,
  \V88(24) ,
  \V88(21) ,
  \V88(20) ,
  \V88(27) ,
  \V88(26) ,
  \V88(29) ,
  \V88(28) ,
  \V88(31) ,
  \V88(30) ,
  \V56(13) ,
  \V56(12) ,
  \V56(15) ,
  \V56(14) ,
  \V24(0) ,
  \V56(11) ,
  \V24(1) ,
  \V56(10) ,
  \V24(2) ,
  \V24(3) ,
  \V24(4) ,
  \V24(5) ,
  \V24(6) ,
  \V56(17) ,
  \V24(7) ,
  \V56(16) ,
  \V24(8) ,
  \V56(19) ,
  \V24(9) ,
  \V56(18) ,
  \V56(23) ,
  \V56(22) ,
  \V56(25) ,
  \V56(24) ,
  \V56(21) ,
  \V56(20) ,
  \V56(27) ,
  \V56(26) ,
  \V56(29) ,
  \V56(28) ,
  \V56(31) ,
  \V56(30) ;
output
  \V151(27) ,
  \V151(26) ,
  \V151(29) ,
  \V151(28) ,
  \V151(21) ,
  \V151(20) ,
  \V151(23) ,
  \V151(22) ,
  \V119(27) ,
  \V151(25) ,
  \V119(26) ,
  \V151(24) ,
  \V119(29) ,
  \V151(17) ,
  \V119(28) ,
  \V151(16) ,
  \V151(19) ,
  \V151(18) ,
  \V119(21) ,
  \V119(20) ,
  \V119(23) ,
  \V151(11) ,
  \V119(22) ,
  \V151(10) ,
  \V119(25) ,
  \V151(3) ,
  \V151(13) ,
  \V119(24) ,
  \V151(2) ,
  \V151(12) ,
  \V119(17) ,
  \V151(5) ,
  \V151(15) ,
  \V119(16) ,
  \V151(4) ,
  \V151(14) ,
  \V119(19) ,
  \V119(18) ,
  \V151(1) ,
  \V151(0) ,
  \V119(11) ,
  \V151(7) ,
  \V119(10) ,
  \V151(6) ,
  \V119(13) ,
  \V151(9) ,
  \V119(12) ,
  \V151(8) ,
  \V119(15) ,
  \V119(14) ,
  \V151(31) ,
  \V151(30) ,
  \V119(30) ,
  \V119(3) ,
  \V119(2) ,
  \V119(5) ,
  \V119(4) ,
  \V119(1) ,
  \V119(0) ,
  \V119(7) ,
  \V119(6) ,
  \V119(9) ,
  \V119(8) ;
wire
  \[0] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \[5] ,
  \[6] ,
  \[7] ,
  \[8] ,
  \[9] ,
  V152,
  V153,
  V154,
  V155,
  V156,
  V157,
  V158,
  V159,
  V160,
  V161,
  V162,
  V163,
  V164,
  V165,
  V166,
  V167,
  V168,
  V169,
  V170,
  V171,
  V175,
  V176,
  V177,
  V178,
  V179,
  V180,
  V181,
  V182,
  V183,
  V184,
  V185,
  V186,
  V187,
  V188,
  V189,
  V190,
  V191,
  V192,
  V193,
  V194,
  V195,
  V196,
  V197,
  V198,
  V199,
  V200,
  V201,
  V202,
  V203,
  V204,
  V205,
  V206,
  V207,
  V208,
  V209,
  V210,
  V211,
  V212,
  V213,
  V214,
  V215,
  V216,
  V217,
  V218,
  V219,
  V220,
  V221,
  V222,
  V223,
  V224,
  V225,
  V226,
  V227,
  V228,
  V229,
  V230,
  V231,
  V232,
  V233,
  V234,
  V235,
  V236,
  V237,
  V238,
  V239,
  V240,
  V241,
  V242,
  V243,
  V244,
  V245,
  V246,
  V247,
  V248,
  V249,
  V250,
  V251,
  V252,
  V253,
  V254,
  V255,
  V256,
  V257,
  V258,
  V259,
  V260,
  V261,
  V262,
  V263,
  V264,
  V265,
  V266,
  V267,
  V268,
  V269,
  V270,
  V271,
  V272,
  V273,
  V274,
  V275,
  V276,
  V277,
  V278,
  V279,
  V280,
  V281,
  V282,
  V283,
  V284,
  V285,
  V286,
  V287,
  V288,
  V289,
  V290,
  V291,
  V292,
  V293,
  V294,
  V295,
  V296,
  V297,
  V298,
  V299,
  V300,
  V301,
  V302,
  V303,
  V304,
  V305,
  V306,
  V307,
  V308,
  V309,
  V310,
  V311,
  V312,
  V313,
  V314,
  V315,
  V316,
  V317,
  V318,
  V319,
  V320,
  V321,
  V322,
  V323,
  V324,
  V325,
  V326,
  V327,
  V328,
  V329,
  V330,
  V331,
  V332,
  V333,
  V334,
  V335,
  V336,
  V337,
  V338,
  V339,
  V340,
  V341,
  V342,
  V343,
  V344,
  V345,
  V346,
  V347,
  V348,
  V349,
  V350,
  V351,
  V352,
  V353,
  V354,
  V355,
  V356,
  V357,
  V358,
  V359,
  V360,
  V361,
  V362,
  V363,
  V364,
  V365,
  V366,
  V367,
  V368,
  V369,
  V370,
  V371,
  V372,
  V373,
  V374,
  V375,
  V376,
  V377,
  V378,
  V379,
  V380,
  V381,
  V382,
  V383,
  V384,
  V385,
  V386,
  V387,
  V388,
  V389,
  V390,
  V391,
  V392,
  V393,
  V394,
  V395,
  V396,
  V397,
  V398,
  V399,
  V400,
  V401,
  V402,
  V403,
  V404,
  V405,
  V406,
  V407,
  V408,
  V409,
  V410,
  V411,
  V412,
  V413,
  V414,
  V415,
  V416,
  V417,
  V418,
  V419,
  V420,
  V421,
  V422,
  V423,
  V424,
  V425,
  V426,
  V427,
  V428,
  V429,
  V430,
  V431,
  V432,
  V433,
  V434,
  V435,
  V436,
  V437,
  V438,
  V439,
  V440,
  V441,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[14] ,
  \[15] ,
  \[16] ,
  \[17] ,
  \[18] ,
  \[19] ,
  \[20] ,
  \[21] ,
  \[22] ,
  \[23] ,
  \[24] ,
  \[25] ,
  \[26] ,
  \[27] ,
  \[28] ,
  \[29] ,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \V174(2) ,
  \[34] ,
  \[35] ,
  \[36] ,
  \[37] ,
  \[38] ,
  \V174(1) ,
  \[39] ,
  \V174(0) ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ,
  \[59] ,
  \[60] ,
  \[61] ,
  \[62] ;
assign
  \V151(27)  = \[51] ,
  \V151(26)  = \[52] ,
  \V151(29)  = \[49] ,
  \V151(28)  = \[50] ,
  \V151(21)  = \[57] ,
  \V151(20)  = \[58] ,
  \V151(23)  = \[55] ,
  \V151(22)  = \[56] ,
  \V119(27)  = \[3] ,
  \V151(25)  = \[53] ,
  \V119(26)  = \[4] ,
  \V151(24)  = \[54] ,
  \V119(29)  = \[1] ,
  \V151(17)  = \[61] ,
  \V119(28)  = \[2] ,
  \V151(16)  = \[62] ,
  \V151(19)  = \[59] ,
  \V151(18)  = \[60] ,
  \V119(21)  = \[9] ,
  \V119(20)  = \[10] ,
  \V119(23)  = \[7] ,
  \V151(11)  = \[35] ,
  \V119(22)  = \[8] ,
  \V151(10)  = \[36] ,
  \V119(25)  = \[5] ,
  \V151(3)  = \[43] ,
  \V151(13)  = \[33] ,
  \V119(24)  = \[6] ,
  \V151(2)  = \[44] ,
  \V151(12)  = \[34] ,
  \V119(17)  = \[13] ,
  \V151(5)  = \[41] ,
  \V151(15)  = \[31] ,
  \V119(16)  = \[14] ,
  \V151(4)  = \[42] ,
  \V151(14)  = \[32] ,
  \V119(19)  = \[11] ,
  \V119(18)  = \[12] ,
  \V151(1)  = \[45] ,
  \V151(0)  = \[46] ,
  \[0]  = V263 | (V232 | (V208 | (V176 | V175))),
  \V119(11)  = \[19] ,
  \[1]  = V264 | (V233 | (V209 | (V177 | V175))),
  \V151(7)  = \[39] ,
  \V119(10)  = \[20] ,
  \[2]  = V265 | (V234 | (V210 | (V178 | V175))),
  \V151(6)  = \[40] ,
  \V119(13)  = \[17] ,
  \[3]  = V266 | (V235 | (V211 | (V179 | V175))),
  \V151(9)  = \[37] ,
  \V119(12)  = \[18] ,
  \[4]  = V267 | (V236 | (V212 | (V180 | V175))),
  \V151(8)  = \[38] ,
  \V119(15)  = \[15] ,
  \[5]  = V268 | (V237 | (V213 | (V181 | V175))),
  \V119(14)  = \[16] ,
  \[6]  = V269 | (V238 | (V214 | (V182 | V175))),
  \[7]  = V270 | (V239 | (V215 | (V183 | V175))),
  \[8]  = V271 | (V240 | (V216 | (V184 | V175))),
  \[9]  = V272 | (V241 | (V217 | (V185 | V175))),
  \V151(31)  = \[47] ,
  \V151(30)  = \[48] ,
  \V119(30)  = \[0] ,
  V152 = \V9(2)  & (\V9(1)  & \V9(3) ),
  V153 = \V9(1)  & \V9(10) ,
  V154 = \V9(2)  & \V9(10) ,
  V155 = ~\V9(0) ,
  V156 = ~\V9(5) ,
  V157 = ~\V9(10) ,
  V158 = V156 & (V155 & V157),
  V159 = ~\V9(2) ,
  V160 = ~\V9(6) ,
  V161 = V160 & (V159 & (\V9(1)  & (V156 & V157))),
  V162 = \V9(7)  & (V155 & V157),
  V163 = \V9(8)  & (\V9(1)  & V157),
  V164 = ~\V9(3) ,
  V165 = V164 & (\V9(1)  & (\V9(2)  & V157)),
  V166 = ~\V9(1) ,
  V167 = V160 & (\V9(2)  & (\V9(0)  & (V166 & (V156 & V157)))),
  V168 = \V9(8)  & (V166 & (\V9(2)  & V157)),
  V169 = V156 & (V166 & (V159 & V160)),
  V170 = V159 & (V166 & \V9(7) ),
  V171 = V159 & (V166 & \V9(10) ),
  V175 = ~\V174(0) ,
  V176 = \V174(0)  & (V426 & (V427 & \V56(31) )),
  V177 = \V174(0)  & (V426 & (V427 & \V56(30) )),
  V178 = \V174(0)  & (V426 & (V427 & \V56(29) )),
  V179 = \V174(0)  & (V426 & (V427 & \V56(28) )),
  V180 = \V174(0)  & (V426 & (V427 & \V56(27) )),
  V181 = \V174(0)  & (V426 & (V427 & \V56(26) )),
  V182 = \V174(0)  & (V426 & (V427 & \V56(25) )),
  V183 = \V174(0)  & (V426 & (V427 & \V56(24) )),
  V184 = \V174(0)  & (V426 & (V427 & \V56(23) )),
  V185 = \V174(0)  & (V426 & (V427 & \V56(22) )),
  V186 = \V174(0)  & (V426 & (V427 & \V56(21) )),
  V187 = \V174(0)  & (V426 & (V427 & \V56(20) )),
  V188 = \V174(0)  & (V426 & (V427 & \V56(19) )),
  V189 = \V174(0)  & (V426 & (V427 & \V56(18) )),
  V190 = \V174(0)  & (V426 & (V427 & \V56(17) )),
  V191 = \V174(0)  & (V426 & (V427 & \V56(16) )),
  V192 = \V174(0)  & (V426 & (V427 & \V56(15) )),
  V193 = \V174(0)  & (V426 & (V427 & \V56(14) )),
  V194 = \V174(0)  & (V426 & (V427 & \V56(13) )),
  V195 = \V174(0)  & (V426 & (V427 & \V56(12) )),
  V196 = \V174(0)  & (V426 & (V427 & \V56(11) )),
  V197 = \V174(0)  & (V426 & (V427 & \V56(10) )),
  V198 = \V174(0)  & (V426 & (V427 & \V56(9) )),
  V199 = \V174(0)  & (V426 & (V427 & \V56(8) )),
  V200 = \V174(0)  & (V426 & (V427 & \V56(7) )),
  V201 = \V174(0)  & (V426 & (V427 & \V56(6) )),
  V202 = \V174(0)  & (V426 & (V427 & \V56(5) )),
  V203 = \V174(0)  & (V426 & (V427 & \V56(4) )),
  V204 = \V174(0)  & (V426 & (V427 & \V56(3) )),
  V205 = \V174(0)  & (V426 & (V427 & \V56(2) )),
  V206 = \V174(0)  & (V426 & (V427 & \V56(1) )),
  V207 = \V174(2)  & (V428 & \V174(0) ),
  V208 = \V56(23)  & V207,
  V209 = \V56(22)  & V207,
  V210 = \V56(21)  & V207,
  V211 = \V56(20)  & V207,
  V212 = \V56(19)  & V207,
  V213 = \V56(18)  & V207,
  V214 = \V56(17)  & V207,
  V215 = \V56(16)  & V207,
  V216 = \V56(15)  & V207,
  V217 = \V56(14)  & V207,
  V218 = \V56(13)  & V207,
  V219 = \V56(12)  & V207,
  V220 = \V56(11)  & V207,
  V221 = \V56(10)  & V207,
  V222 = \V56(9)  & V207,
  V223 = \V56(8)  & V207,
  V224 = \V56(7)  & V207,
  V225 = \V56(6)  & V207,
  V226 = \V56(5)  & V207,
  V227 = \V56(4)  & V207,
  V228 = \V56(3)  & V207,
  V229 = \V56(2)  & V207,
  V230 = \V56(1)  & V207,
  V231 = \V56(0)  & V207,
  V232 = \V174(0)  & (\V174(1)  & (V429 & \V56(20) )),
  V233 = \V174(0)  & (\V174(1)  & (V429 & \V56(19) )),
  V234 = \V174(0)  & (\V174(1)  & (V429 & \V56(18) )),
  V235 = \V174(0)  & (\V174(1)  & (V429 & \V56(17) )),
  V236 = \V174(0)  & (\V174(1)  & (V429 & \V56(16) )),
  V237 = \V174(0)  & (\V174(1)  & (V429 & \V56(15) )),
  V238 = \V174(0)  & (\V174(1)  & (V429 & \V56(14) )),
  V239 = \V174(0)  & (\V174(1)  & (V429 & \V56(13) )),
  V240 = \V174(0)  & (\V174(1)  & (V429 & \V56(12) )),
  V241 = \V174(0)  & (\V174(1)  & (V429 & \V56(11) )),
  V242 = \V174(0)  & (\V174(1)  & (V429 & \V56(10) )),
  V243 = \V174(0)  & (\V174(1)  & (V429 & \V56(9) )),
  V244 = \V174(0)  & (\V174(1)  & (V429 & \V56(8) )),
  V245 = \V174(0)  & (\V174(1)  & (V429 & \V56(7) )),
  V246 = \V174(0)  & (\V174(1)  & (V429 & \V56(6) )),
  V247 = \V174(0)  & (\V174(1)  & (V429 & \V56(5) )),
  V248 = \V174(0)  & (\V174(1)  & (V429 & \V56(4) )),
  V249 = \V174(0)  & (\V174(1)  & (V429 & \V56(3) )),
  V250 = \V174(0)  & (\V174(1)  & (V429 & \V56(2) )),
  V251 = \V174(0)  & (\V174(1)  & (V429 & \V56(1) )),
  V252 = \V174(0)  & (\V174(1)  & (V429 & \V88(11) )),
  V253 = \V174(0)  & (\V174(1)  & (V429 & \V88(10) )),
  V254 = \V174(0)  & (\V174(1)  & (V429 & \V88(9) )),
  V255 = \V174(0)  & (\V174(1)  & (V429 & \V88(8) )),
  V256 = \V174(0)  & (\V174(1)  & (V429 & \V88(7) )),
  V257 = \V174(0)  & (\V174(1)  & (V429 & \V88(6) )),
  V258 = \V174(0)  & (\V174(1)  & (V429 & \V88(5) )),
  V259 = \V174(0)  & (\V174(1)  & (V429 & \V88(4) )),
  V260 = \V174(0)  & (\V174(1)  & (V429 & \V88(3) )),
  V261 = \V174(0)  & (\V174(1)  & (V429 & \V88(2) )),
  V262 = \V174(0)  & (\V174(1)  & (V429 & \V88(1) )),
  V263 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(16) )),
  V264 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(15) )),
  V265 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(14) )),
  V266 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(13) )),
  V267 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(12) )),
  V268 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(11) )),
  V269 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(10) )),
  V270 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(9) )),
  V271 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(8) )),
  V272 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(7) )),
  V273 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(6) )),
  V274 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(5) )),
  V275 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(4) )),
  V276 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(3) )),
  V277 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(2) )),
  V278 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(1) )),
  V279 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V24(14) )),
  V280 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V24(13) )),
  V281 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V24(12) )),
  V282 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V24(11) )),
  V283 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V24(10) )),
  V284 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V24(9) )),
  V285 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V24(8) )),
  V286 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V24(7) )),
  V287 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V24(6) )),
  V288 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V24(5) )),
  V289 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V24(4) )),
  V290 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V24(3) )),
  V291 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V24(2) )),
  V292 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V24(1) )),
  V293 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V24(0) )),
  V294 = V432 & (V431 & V430),
  V295 = \V174(2)  & (V434 & V433),
  V296 = V436 & (\V174(1)  & V435),
  V297 = \V174(2)  & (\V174(1)  & V437),
  V298 = \V174(0)  & (V438 & (V439 & \V88(31) )),
  V299 = \V174(0)  & (V438 & (V439 & \V88(30) )),
  V300 = \V174(0)  & (V438 & (V439 & \V88(29) )),
  V301 = \V174(0)  & (V438 & (V439 & \V88(28) )),
  V302 = \V174(0)  & (V438 & (V439 & \V88(27) )),
  V303 = \V174(0)  & (V438 & (V439 & \V88(26) )),
  V304 = \V174(0)  & (V438 & (V439 & \V88(25) )),
  V305 = \V174(0)  & (V438 & (V439 & \V88(24) )),
  V306 = \V174(0)  & (V438 & (V439 & \V88(23) )),
  V307 = \V174(0)  & (V438 & (V439 & \V88(22) )),
  V308 = \V174(0)  & (V438 & (V439 & \V88(21) )),
  V309 = \V174(0)  & (V438 & (V439 & \V88(20) )),
  V310 = \V174(0)  & (V438 & (V439 & \V88(19) )),
  V311 = \V174(0)  & (V438 & (V439 & \V88(18) )),
  V312 = \V174(0)  & (V438 & (V439 & \V88(17) )),
  V313 = \V174(0)  & (V438 & (V439 & \V88(16) )),
  V314 = \V174(0)  & (V438 & (V439 & \V88(15) )),
  V315 = \V174(0)  & (V438 & (V439 & \V88(14) )),
  V316 = \V174(0)  & (V438 & (V439 & \V88(13) )),
  V317 = \V174(0)  & (V438 & (V439 & \V88(12) )),
  V318 = \V174(0)  & (V438 & (V439 & \V88(11) )),
  V319 = \V174(0)  & (V438 & (V439 & \V88(10) )),
  V320 = \V174(0)  & (V438 & (V439 & \V88(9) )),
  V321 = \V174(0)  & (V438 & (V439 & \V88(8) )),
  V322 = \V174(0)  & (V438 & (V439 & \V88(7) )),
  V323 = \V174(0)  & (V438 & (V439 & \V88(6) )),
  V324 = \V174(0)  & (V438 & (V439 & \V88(5) )),
  V325 = \V174(0)  & (V438 & (V439 & \V88(4) )),
  V326 = \V174(0)  & (V438 & (V439 & \V88(3) )),
  V327 = \V174(0)  & (V438 & (V439 & \V88(2) )),
  V328 = \V174(0)  & (V438 & (V439 & \V88(1) )),
  V329 = \V174(0)  & (V438 & (V439 & \V88(0) )),
  V330 = \V174(0)  & (V440 & (\V174(2)  & \V88(23) )),
  V331 = \V174(0)  & (V440 & (\V174(2)  & \V88(22) )),
  V332 = \V174(0)  & (V440 & (\V174(2)  & \V88(21) )),
  V333 = \V174(0)  & (V440 & (\V174(2)  & \V88(20) )),
  V334 = \V174(0)  & (V440 & (\V174(2)  & \V88(19) )),
  V335 = \V174(0)  & (V440 & (\V174(2)  & \V88(18) )),
  V336 = \V174(0)  & (V440 & (\V174(2)  & \V88(17) )),
  V337 = \V174(0)  & (V440 & (\V174(2)  & \V88(16) )),
  V338 = \V174(0)  & (V440 & (\V174(2)  & \V88(15) )),
  V339 = \V174(0)  & (V440 & (\V174(2)  & \V88(14) )),
  V340 = \V174(0)  & (V440 & (\V174(2)  & \V88(13) )),
  V341 = \V174(0)  & (V440 & (\V174(2)  & \V88(12) )),
  V342 = \V174(0)  & (V440 & (\V174(2)  & \V88(11) )),
  V343 = \V174(0)  & (V440 & (\V174(2)  & \V88(10) )),
  V344 = \V174(0)  & (V440 & (\V174(2)  & \V88(9) )),
  V345 = \V174(0)  & (V440 & (\V174(2)  & \V88(8) )),
  V346 = \V174(0)  & (V440 & (\V174(2)  & \V88(7) )),
  V347 = \V174(0)  & (V440 & (\V174(2)  & \V88(6) )),
  V348 = \V174(0)  & (V440 & (\V174(2)  & \V88(5) )),
  V349 = \V174(0)  & (V440 & (\V174(2)  & \V88(4) )),
  V350 = \V174(0)  & (V440 & (\V174(2)  & \V88(3) )),
  V351 = \V174(0)  & (V440 & (\V174(2)  & \V88(2) )),
  V352 = \V174(0)  & (V440 & (\V174(2)  & \V88(1) )),
  V353 = \V174(0)  & (V440 & (\V174(2)  & \V88(0) )),
  V354 = \V174(0)  & (V440 & (\V174(2)  & \V56(31) )),
  V355 = \V174(0)  & (V440 & (\V174(2)  & \V56(30) )),
  V356 = \V174(0)  & (V440 & (\V174(2)  & \V56(29) )),
  V357 = \V174(0)  & (V440 & (\V174(2)  & \V56(28) )),
  V358 = \V174(0)  & (V440 & (\V174(2)  & \V56(27) )),
  V359 = \V174(0)  & (V440 & (\V174(2)  & \V56(26) )),
  V360 = \V174(0)  & (V440 & (\V174(2)  & \V56(25) )),
  V361 = \V174(0)  & (V440 & (\V174(2)  & \V56(24) )),
  V362 = \V174(0)  & (\V174(1)  & (V441 & \V88(20) )),
  V363 = \V174(0)  & (\V174(1)  & (V441 & \V88(19) )),
  V364 = \V174(0)  & (\V174(1)  & (V441 & \V88(18) )),
  V365 = \V174(0)  & (\V174(1)  & (V441 & \V88(17) )),
  V366 = \V174(0)  & (\V174(1)  & (V441 & \V88(16) )),
  V367 = \V174(0)  & (\V174(1)  & (V441 & \V88(15) )),
  V368 = \V174(0)  & (\V174(1)  & (V441 & \V88(14) )),
  V369 = \V174(0)  & (\V174(1)  & (V441 & \V88(13) )),
  V370 = \V174(0)  & (\V174(1)  & (V441 & \V88(12) )),
  V371 = \V174(0)  & (\V174(1)  & (V441 & \V88(11) )),
  V372 = \V174(0)  & (\V174(1)  & (V441 & \V88(10) )),
  V373 = \V174(0)  & (\V174(1)  & (V441 & \V88(9) )),
  V374 = \V174(0)  & (\V174(1)  & (V441 & \V88(8) )),
  V375 = \V174(0)  & (\V174(1)  & (V441 & \V88(7) )),
  V376 = \V174(0)  & (\V174(1)  & (V441 & \V88(6) )),
  V377 = \V174(0)  & (\V174(1)  & (V441 & \V88(5) )),
  V378 = \V174(0)  & (\V174(1)  & (V441 & \V88(4) )),
  V379 = \V174(0)  & (\V174(1)  & (V441 & \V88(3) )),
  V380 = \V174(0)  & (\V174(1)  & (V441 & \V88(2) )),
  V381 = \V174(0)  & (\V174(1)  & (V441 & \V88(1) )),
  V382 = \V174(0)  & (\V174(1)  & (V441 & \V88(0) )),
  V383 = \V174(0)  & (\V174(1)  & (V441 & \V56(31) )),
  V384 = \V174(0)  & (\V174(1)  & (V441 & \V56(30) )),
  V385 = \V174(0)  & (\V174(1)  & (V441 & \V56(29) )),
  V386 = \V174(0)  & (\V174(1)  & (V441 & \V56(28) )),
  V387 = \V174(0)  & (\V174(1)  & (V441 & \V56(27) )),
  V388 = \V174(0)  & (\V174(1)  & (V441 & \V56(26) )),
  V389 = \V174(0)  & (\V174(1)  & (V441 & \V56(25) )),
  V390 = \V174(0)  & (\V174(1)  & (V441 & \V56(24) )),
  V391 = \V174(0)  & (\V174(1)  & (V441 & \V56(23) )),
  V392 = \V174(0)  & (\V174(1)  & (V441 & \V56(22) )),
  V393 = \V174(0)  & (\V174(1)  & (V441 & \V56(21) )),
  V394 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(16) )),
  V395 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(15) )),
  V396 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(14) )),
  V397 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(13) )),
  V398 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(12) )),
  V399 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(11) )),
  V400 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(10) )),
  V401 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(9) )),
  V402 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(8) )),
  V403 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(7) )),
  V404 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(6) )),
  V405 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(5) )),
  V406 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(4) )),
  V407 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(3) )),
  V408 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(2) )),
  V409 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(1) )),
  V410 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V88(0) )),
  V411 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(31) )),
  V412 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(30) )),
  V413 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(29) )),
  V414 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(28) )),
  V415 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(27) )),
  V416 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(26) )),
  V417 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(25) )),
  V418 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(24) )),
  V419 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(23) )),
  V420 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(22) )),
  V421 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(21) )),
  V422 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(20) )),
  V423 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(19) )),
  V424 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(18) )),
  V425 = \V174(0)  & (\V174(1)  & (\V174(2)  & \V56(17) )),
  V426 = ~\V174(1) ,
  V427 = ~\V174(2) ,
  V428 = ~\V174(1) ,
  V429 = ~\V174(2) ,
  V430 = ~\V174(0) ,
  V431 = ~\V174(1) ,
  V432 = ~\V174(2) ,
  V433 = ~\V174(0) ,
  V434 = ~\V174(1) ,
  V435 = ~\V174(0) ,
  V436 = ~\V174(2) ,
  V437 = ~\V174(0) ,
  V438 = ~\V174(1) ,
  V439 = ~\V174(2) ,
  V440 = ~\V174(1) ,
  V441 = ~\V174(2) ,
  \V119(3)  = \[27] ,
  \V119(2)  = \[28] ,
  \V119(5)  = \[25] ,
  \V119(4)  = \[26] ,
  \[10]  = V273 | (V242 | (V218 | (V186 | V175))),
  \[11]  = V274 | (V243 | (V219 | (V187 | V175))),
  \V119(1)  = \[29] ,
  \[12]  = V275 | (V244 | (V220 | (V188 | V175))),
  \V119(0)  = \[30] ,
  \[13]  = V276 | (V245 | (V221 | (V189 | V175))),
  \[14]  = V277 | (V246 | (V222 | (V190 | V175))),
  \[15]  = V278 | (V247 | (V223 | (V191 | V175))),
  \[16]  = V279 | (V248 | (V224 | (V192 | V175))),
  \[17]  = V280 | (V249 | (V225 | (V193 | V175))),
  \V119(7)  = \[23] ,
  \[18]  = V281 | (V250 | (V226 | (V194 | V175))),
  \V119(6)  = \[24] ,
  \[19]  = V282 | (V251 | (V227 | (V195 | V175))),
  \V119(9)  = \[21] ,
  \V119(8)  = \[22] ,
  \[20]  = V283 | (V252 | (V228 | (V196 | V175))),
  \[21]  = V284 | (V253 | (V229 | (V197 | V175))),
  \[22]  = V285 | (V254 | (V230 | (V198 | V175))),
  \[23]  = V286 | (V255 | (V231 | (V199 | V175))),
  \[24]  = V287 | (V256 | (V207 | (V200 | V175))),
  \[25]  = V288 | (V257 | (V207 | (V201 | V175))),
  \[26]  = V289 | (V258 | (V207 | (V202 | V175))),
  \[27]  = V290 | (V259 | (V207 | (V203 | V175))),
  \[28]  = V291 | (V260 | (V207 | (V204 | V175))),
  \[29]  = V292 | (V261 | (V207 | (V205 | V175))),
  \[30]  = V293 | (V262 | (V207 | (V206 | V175))),
  \[31]  = V410 | (V378 | (V346 | (V314 | (V297 | (V296 | (V295 | V294)))))),
  \[32]  = V411 | (V379 | (V347 | (V315 | (V297 | (V296 | (V295 | V294)))))),
  \[33]  = V412 | (V380 | (V348 | (V316 | (V297 | (V296 | (V295 | V294)))))),
  \V174(2)  = V171 | (V169 | (V170 | (V161 | (V158 | (V162 | V163))))),
  \[34]  = V413 | (V381 | (V349 | (V317 | (V297 | (V296 | (V295 | V294)))))),
  \[35]  = V414 | (V382 | (V350 | (V318 | (V297 | (V296 | (V295 | V294)))))),
  \[36]  = V415 | (V383 | (V351 | (V319 | (V297 | (V296 | (V295 | V294)))))),
  \[37]  = V416 | (V384 | (V352 | (V320 | (V297 | (V296 | (V295 | V294)))))),
  \[38]  = V417 | (V385 | (V353 | (V321 | (V297 | (V296 | (V295 | V294)))))),
  \V174(1)  = V171 | (V169 | (V170 | (V165 | (V167 | V168)))),
  \[39]  = V418 | (V386 | (V354 | (V322 | (V297 | (V296 | (V295 | V294)))))),
  \V174(0)  = V168 | (V167 | (V165 | (V163 | (V161 | (V158 | (V162 | (V152 | (V153 | (V154 | (V169 | (V170 | V171))))))))))),
  \[40]  = V419 | (V387 | (V355 | (V323 | (V297 | (V296 | (V295 | V294)))))),
  \[41]  = V420 | (V388 | (V356 | (V324 | (V297 | (V296 | (V295 | V294)))))),
  \[42]  = V421 | (V389 | (V357 | (V325 | (V297 | (V296 | (V295 | V294)))))),
  \[43]  = V422 | (V390 | (V358 | (V326 | (V297 | (V296 | (V295 | V294)))))),
  \[44]  = V423 | (V391 | (V359 | (V327 | (V297 | (V296 | (V295 | V294)))))),
  \[45]  = V424 | (V392 | (V360 | (V328 | (V297 | (V296 | (V295 | V294)))))),
  \[46]  = V425 | (V393 | (V361 | (V329 | (V297 | (V296 | (V295 | V294)))))),
  \[47]  = V394 | (V362 | (V330 | (V298 | (V297 | (V296 | (V295 | V294)))))),
  \[48]  = V395 | (V363 | (V331 | (V299 | (V297 | (V296 | (V295 | V294)))))),
  \[49]  = V396 | (V364 | (V332 | (V300 | (V297 | (V296 | (V295 | V294)))))),
  \[50]  = V397 | (V365 | (V333 | (V301 | (V297 | (V296 | (V295 | V294)))))),
  \[51]  = V398 | (V366 | (V334 | (V302 | (V297 | (V296 | (V295 | V294)))))),
  \[52]  = V399 | (V367 | (V335 | (V303 | (V297 | (V296 | (V295 | V294)))))),
  \[53]  = V400 | (V368 | (V336 | (V304 | (V297 | (V296 | (V295 | V294)))))),
  \[54]  = V401 | (V369 | (V337 | (V305 | (V297 | (V296 | (V295 | V294)))))),
  \[55]  = V402 | (V370 | (V338 | (V306 | (V297 | (V296 | (V295 | V294)))))),
  \[56]  = V403 | (V371 | (V339 | (V307 | (V297 | (V296 | (V295 | V294)))))),
  \[57]  = V404 | (V372 | (V340 | (V308 | (V297 | (V296 | (V295 | V294)))))),
  \[58]  = V405 | (V373 | (V341 | (V309 | (V297 | (V296 | (V295 | V294)))))),
  \[59]  = V406 | (V374 | (V342 | (V310 | (V297 | (V296 | (V295 | V294)))))),
  \[60]  = V407 | (V375 | (V343 | (V311 | (V297 | (V296 | (V295 | V294)))))),
  \[61]  = V408 | (V376 | (V344 | (V312 | (V297 | (V296 | (V295 | V294)))))),
  \[62]  = V409 | (V377 | (V345 | (V313 | (V297 | (V296 | (V295 | V294))))));
endmodule

