//NOTE: no-implementation module stub

module lmi_dram (
    input wire CLK,
    input wire TMODE,
    input wire RESET_D1_R_N,
    input wire DISABLEC,
    input wire CFG_DWDISW,
    input wire EXT_DWREQRAM_R,
    input wire DW_GNTRAM_R,
    input wire DATAIN,
    output wire DW_DATAOUT,
    output wire DW_DATAOE,
    input wire NEXTADDR,
    input wire NEXTRDOP,
    input wire NEXTWROP,
    input wire NEXTBE,
    input wire NEXTSX,
    output wire EXCP,
    output wire DW_VAL,
    output wire DW_ACK,
    output wire X_HALT_R,
    output wire DC_RPQUIETIFNBA,
    output wire DC_RPQUIETIFB,
    output wire DC_RPALGNIFNBNA,
    output wire DC_RPALGNIFB,
    output wire DW_HALT_W_R,
    input wire DW_DATAINDEX,
    input wire DWR_DATARD,
    input wire DW_DATAWR,
    input wire DW_DATAWE,
    input wire DW_DATAWEN,
    input wire DW_DATARE,
    input wire DW_DATAREN,
    input wire DW_DATACS,
    input wire DW_DATACSN,
    input wire CONFIGBASE,
    input wire CONFIGTOP
);

endmodule
