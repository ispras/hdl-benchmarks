`timescale 1 ps / 1 ps

module carry (goofy_bach, ceres_elian_outwire);
  input goofy_bach;
  output ceres_elian_outwire;
endmodule
