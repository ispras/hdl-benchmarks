module s953_bench(
  blif_clk_net,
  blif_reset_net,
  Rdy1RtHS1,
  Rdy2RtHS1,
  Rdy1BmHS1,
  Rdy2BmHS1,
  IInDoneHS1,
  RtTSHS1,
  TpArrayHS1,
  OutputHS1,
  WantBmHS1,
  WantRtHS1,
  OutAvHS1,
  FullOHS1,
  FullIIHS1,
  Prog_2,
  Prog_1,
  Prog_0,
  ReWhBufHS1,
  TgWhBufHS1,
  SeOutAvHS1,
  LdProgHS1,
  Mode2HS1,
  ReRtTSHS1,
  ShftIIRHS1,
  NewTrHS1,
  Mode1HS1,
  ShftORHS1,
  ActRtHS1,
  Mode0HS1,
  TxHIInHS1,
  LxHIInHS1,
  NewLineHS1,
  ActBmHS1,
  GoBmHS1,
  LoadOHHS1,
  DumpIIHS1,
  SeFullOHS1,
  GoRtHS1,
  LoadIIHHS1,
  SeFullIIHS1);
input blif_clk_net;
input blif_reset_net;
input Rdy1RtHS1;
input Rdy2RtHS1;
input Rdy1BmHS1;
input Rdy2BmHS1;
input IInDoneHS1;
input RtTSHS1;
input TpArrayHS1;
input OutputHS1;
input WantBmHS1;
input WantRtHS1;
input OutAvHS1;
input FullOHS1;
input FullIIHS1;
input Prog_2;
input Prog_1;
input Prog_0;
output ReWhBufHS1;
output TgWhBufHS1;
output SeOutAvHS1;
output LdProgHS1;
output Mode2HS1;
output ReRtTSHS1;
output ShftIIRHS1;
output NewTrHS1;
output Mode1HS1;
output ShftORHS1;
output ActRtHS1;
output Mode0HS1;
output TxHIInHS1;
output LxHIInHS1;
output NewLineHS1;
output ActBmHS1;
output GoBmHS1;
output LoadOHHS1;
output DumpIIHS1;
output SeFullOHS1;
output GoRtHS1;
output LoadIIHHS1;
output SeFullIIHS1;
reg State_5;
reg State_4;
reg State_3;
reg State_2;
reg State_1;
reg State_0;
reg _8383_;
reg _8388_;
reg _8393_;
reg _8389_;
reg _8380_;
reg _8378_;
reg _8384_;
reg _8381_;
reg _8377_;
reg _8387_;
reg _8382_;
reg _8379_;
reg _8386_;
reg _8385_;
reg _8390_;
reg _8394_;
reg _8375_;
reg _8392_;
reg _8395_;
reg _8374_;
reg _8373_;
reg _8376_;
reg _8391_;
wire II372;
wire II425;
wire II699;
wire II789_1;
wire II351;
wire II1154_1;
wire II263;
wire II1166_2;
wire II1031_1;
wire II504;
wire II663;
wire II476;
wire II599;
wire II810_1;
wire II861_1;
wire II339;
wire II407;
wire II725;
wire II715;
wire II595;
wire II587;
wire II517;
wire II531;
wire II682;
wire II796_1;
wire II523;
wire II731;
wire II9;
wire II585;
wire II1160_1;
wire II1077_1;
wire II447;
wire II497;
wire II1047_1;
wire II1028_1;
wire II1196_1;
wire II418;
wire II1125_1;
wire II659;
wire II1207_1;
wire II779;
wire II571;
wire II686;
wire II577;
wire II363;
wire II283;
wire II689;
wire II1163_1;
wire II509;
wire II469;
wire II15;
wire II266;
wire II1103_2;
wire II474;
wire II4;
wire II366;
wire II343;
wire II278;
wire II440;
wire II513;
wire II481;
wire II25;
wire II466;
wire II704;
wire II514;
wire II348;
wire II1143_1;
wire II768;
wire II362;
wire II415;
wire II8;
wire II487;
wire II1083_1;
wire II609;
wire II422;
wire II750;
wire II1044_1;
wire II556;
wire II503;
wire II840_1;
wire II892_2;
wire II532;
wire II511;
wire II437;
wire II493;
wire II297;
wire II771;
wire II1157_1;
wire II379;
wire II521;
wire II671;
wire II382;
wire II18;
wire II1080_1;
wire II439;
wire II29;
wire II543;
wire II695;
wire II431;
wire II300;
wire II1173_1;
wire II336;
wire II355;
wire II555;
wire II1136_1;
wire II498;
wire II399;
wire II347;
wire II328;
wire II279;
wire II508;
wire II829_1;
wire II1184_2;
wire II1140_1;
wire II315;
wire II1040_1;
wire II655;
wire II333;
wire II746;
wire II318;
wire II735;
wire II568;
wire II479;
wire II21;
wire II551;
wire II624;
wire II458;
wire II1037_1;
wire II489;
wire II16;
wire II446;
wire II338;
wire II770;
wire II1176_2;
wire II596;
wire II575;
wire II1151_1;
wire II485;
wire II548;
wire II390;
wire II12;
wire II614;
wire II691;
wire II1199_1;
wire II398;
wire II404;
wire II386;
wire II1193_1;
wire II376;
wire II5;
wire II274;
wire II364;
wire II545;
wire II562;
wire II282;
wire II475;
wire II534;
wire II1132_2;
wire II1213_1;
wire II329;
wire II311;
wire II1216_1;
wire II1210_1;
wire II1113_1;
wire II410;
wire II13;
wire II450;
wire II423;
wire II697;
wire II405;
wire II275;
wire II580;
wire II537;
wire II1091_1;
wire II465;
wire II559;
wire II449;
wire II30;
wire II1107_1;
wire II24;
wire II740;
wire II711;
wire II359;
wire II512;
wire II442;
wire II680;
wire II367;
wire II554;
wire II416;
wire II1188_1;
wire II519;
wire II370;
wire II294;
wire II457;
wire II1188_2;
wire II414;
wire II723;
wire II567;
wire II264;
wire II335;
wire II673;
wire II354;
wire II1148_1;
wire II267;
wire II434;
wire II393;
wire II1118_1;
wire II461;
wire II910_1;
wire II17;
wire II660;
wire II342;
wire II357;
wire II665;
wire II539;
wire II27;
wire II20;
wire II702;
wire II1199_2;
wire II593;
wire II377;
wire II661;
wire II494;
wire II394;
wire II269;
wire II657;
wire II547;
wire II840_2;
wire II535;
wire II326;
wire II397;
wire II1184_1;
wire II565;
wire II693;
wire II625;
wire II896_1;
wire II676;
wire II767;
wire II495;
wire II963_1;
wire II7;
wire II733;
wire II271;
wire II1110_1;
wire II1034_1;
wire II322;
wire II451;
wire II1121_1;
wire II850_2;
wire II6;
wire II486;
wire II506;
wire II525;
wire II411;
wire II526;
wire II10;
wire II353;
wire II445;
wire II281;
wire II1203_1;
wire II325;
wire II1103_1;
wire II966_1;
wire II23;
wire II561;
wire II14;
wire II430;
wire II690;
wire II491;
wire II396;
wire II1056_1;
wire II529;
wire II276;
wire II1180_2;
wire II403;
wire II706;
wire II684;
wire II380;
wire II873_1;
wire II295;
wire II814_1;
wire II424;
wire II553;
wire II1166_1;
wire II738;
wire II468;
wire II717;
wire II287;
wire II360;
wire II341;
wire II350;
wire II881_2;
wire II330;
wire II345;
wire II374;
wire II1180_1;
wire II505;
wire II435;
wire II1094_1;
wire II284;
wire II1121_2;
wire II881_1;
wire II861_2;
wire II470;
wire II573;
wire II857_1;
wire II1100_1;
wire II331;
wire II1047_2;
wire II500;
wire II744;
wire II1087_1;
wire II610;
wire II667;
wire II11;
wire II1025_1;
wire II371;
wire II675;
wire II729;
wire II303;
wire II384;
wire II327;
wire II552;
wire II381;
wire II358;
wire II388;
wire II320;
wire II721;
wire II850_1;
wire II1132_1;
wire II477;
wire II1203_2;
wire II408;
wire II323;
wire II452;
wire II566;
wire II1216_2;
wire II272;
wire II277;
wire II421;
wire II540;
wire II634;
wire II600;
wire II2;
wire II441;
wire II429;
wire II778;
wire II317;
wire II708;
wire II590;
wire II412;
wire II570;
wire II612;
wire II737;
wire II1170_1;
wire II834_1;
wire II719;
wire II459;
wire II1128_1;
wire II455;
wire II19;
wire II467;
wire II579;
wire II428;
wire II1176_1;
wire II713;
wire II582;
wire II391;
wire II26;
wire II1097_1;
wire II340;
wire II669;
wire II280;
wire II662;
wire II463;
wire II453;
wire II742;
wire II769;
wire II589;
wire II700;
wire II777;
wire II432;
wire II344;
wire II265;
wire II22;
wire II482;
wire II678;
wire II28;
wire II436;
wire II473;
wire II3;
wire II892_1;
wire II1143_2;
wire II444;
wire II378;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    State_5 <= 0;
  else
    State_5 <= II2;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    State_4 <= 0;
  else
    State_4 <= II3;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    State_3 <= 0;
  else
    State_3 <= II4;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    State_2 <= 0;
  else
    State_2 <= II5;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    State_1 <= 0;
  else
    State_1 <= II6;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    State_0 <= 0;
  else
    State_0 <= II7;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8383_ <= 0;
  else
    _8383_ <= II8;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8388_ <= 0;
  else
    _8388_ <= II9;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8393_ <= 0;
  else
    _8393_ <= II10;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8389_ <= 0;
  else
    _8389_ <= II11;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8380_ <= 0;
  else
    _8380_ <= II12;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8378_ <= 0;
  else
    _8378_ <= II13;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8384_ <= 0;
  else
    _8384_ <= II14;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8381_ <= 0;
  else
    _8381_ <= II15;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8377_ <= 0;
  else
    _8377_ <= II16;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8387_ <= 0;
  else
    _8387_ <= II17;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8382_ <= 0;
  else
    _8382_ <= II18;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8379_ <= 0;
  else
    _8379_ <= II19;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8386_ <= 0;
  else
    _8386_ <= II20;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8385_ <= 0;
  else
    _8385_ <= II21;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8390_ <= 0;
  else
    _8390_ <= II22;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8394_ <= 0;
  else
    _8394_ <= II23;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8375_ <= 0;
  else
    _8375_ <= II24;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8392_ <= 0;
  else
    _8392_ <= II25;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8395_ <= 0;
  else
    _8395_ <= II26;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8374_ <= 0;
  else
    _8374_ <= II27;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8373_ <= 0;
  else
    _8373_ <= II28;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8376_ <= 0;
  else
    _8376_ <= II29;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    _8391_ <= 0;
  else
    _8391_ <= II30;
assign II372 = ((~II892_1))|((~II892_2));
assign II699 = ((~II1143_1)&(~II1143_2));
assign II425 = ((~State_2))|((~II281))|((~II508));
assign II789_1 = (II278&II580);
assign II351 = ((~II350));
assign II1154_1 = (II267)|(II371);
assign II263 = ((~Rdy1RtHS1));
assign II1166_2 = (Prog_2&II452);
assign II1031_1 = (II317&II398);
assign II504 = ((~II505));
assign II663 = ((~II662));
assign II476 = ((~II519)&(~II545));
assign II599 = ((~II275))|((~II354));
assign II810_1 = (II364&II562);
assign II861_1 = (II263)|(II455);
assign II339 = ((~II338));
assign II725 = ((~II1184_1)&(~II1184_2));
assign II407 = ((~II412))|((~II532));
assign II715 = ((~II1166_1)&(~II1166_2));
assign II595 = ((~Rdy2BmHS1))|((~II274));
assign II517 = ((~II264))|((~II358));
assign II682 = ((~II1118_1))|((~II323));
assign II587 = ((~Prog_0))|((~II317));
assign II796_1 = (II283)|(II323);
assign II531 = ((~II429))|((~II491));
assign II523 = ((~II274))|((~Prog_2));
assign II731 = ((~II540)&(~II474));
assign II9 = ((~II377))|((~II661))|((~II659));
assign II585 = ((~II353))|((~II422));
assign II1160_1 = (II281&II412);
assign II1077_1 = (II458&II512);
assign II447 = ((~Rdy2RtHS1))|((~II362));
assign II497 = ((~II455))|((~II457));
assign II1047_1 = (II264)|(II284);
assign II1028_1 = (II367)|(II493);
assign II1196_1 = (II345&II418);
assign II418 = ((~II279)&(~II485));
assign II659 = ((~II322)&(~II1083_1));
assign II1125_1 = (Rdy2RtHS1)|(II561);
assign II1207_1 = (II519)|(II579);
assign II779 = ((~II778));
assign II571 = ((~II570));
assign II686 = ((~II1125_1))|((~II441));
assign II577 = ((~State_0))|((~II318))|((~II436));
assign II363 = ((~II362));
assign II283 = ((~Prog_1));
assign II689 = ((~II440)&(~II1128_1));
assign II1163_1 = (II345&II531);
assign II469 = ((~II468));
assign II509 = ((~II276))|((~II277));
assign II15 = ((~II796_1))|((~II675));
assign II266 = ((~Rdy2BmHS1));
assign II1103_2 = (Prog_0&II322);
assign II474 = ((~II493)&(~II577));
assign II4 = ((~II725))|((~II381))|((~II551));
assign II366 = ((~State_0)&(~II335)&(~II399));
assign II343 = ((~II276))|((~II394))|((~II482));
assign II278 = ((~State_3));
assign II481 = ((~II372))|((~II486));
assign II25 = ((~II814_1))|((~II767));
assign II513 = ((~II512));
assign II440 = ((~II495)&(~II509));
assign II466 = ((~Rdy1BmHS1)&(~II503));
assign II704 = ((~II1151_1))|((~II329));
assign II514 = ((~II263)&(~Rdy2RtHS1));
assign II348 = ((~II315)&(~II363));
assign II1143_1 = (II353&II404);
assign II768 = ((~II719))|((~II717));
assign II362 = ((~State_0)&(~II407));
assign II415 = ((~II414));
assign II8 = ((~II655))|((~II657));
assign II487 = ((~State_3))|((~II508));
assign II1083_1 = (II458&II506);
assign II609 = ((~II265))|((~II434));
assign II422 = ((~II431)&(~II525));
assign II750 = ((~II665))|((~II663));
assign II1044_1 = (II497&II570);
assign II556 = ((~II1028_1))|((~II355));
assign II503 = ((~II277))|((~II504));
assign II840_1 = (II283&II284);
assign II532 = ((~State_4)&(~II327));
assign II511 = ((~State_1))|((~State_0));
assign II892_2 = (II269)|(II625);
assign II437 = ((~II436));
assign II493 = ((~Rdy1BmHS1))|((~II266));
assign II297 = ((~II376)&(~II686)&(~II684));
assign II771 = ((~II770));
assign II1157_1 = (II274)|(II599);
assign II521 = ((~RtTSHS1))|((~II278));
assign II379 = ((~II378));
assign II671 = ((~II1103_1)&(~II1103_2));
assign II382 = ((~II276)&(~Prog_2)&(~II485));
assign II18 = ((~II295));
assign II1080_1 = (Prog_0&II382);
assign II439 = ((~Prog_0))|((~II514));
assign II29 = ((~II278)&(~State_2)&(~II441));
assign II543 = ((~II265))|((~Rdy2BmHS1));
assign II695 = ((~II408)&(~II328));
assign II431 = ((~II430));
assign II300 = ((~II700)&(~II810_1));
assign II1173_1 = (II263&II466);
assign II336 = ((~II473))|((~II357));
assign II355 = ((~II354));
assign II555 = ((~II330)&(~II1025_1));
assign II1136_1 = (II282&II590);
assign II498 = ((~II271)&(~II473));
assign II399 = ((~II284))|((~II436));
assign II347 = ((~State_3)&(~II394));
assign II328 = ((~II609)&(~II511)&(~II539));
assign II279 = ((~State_2));
assign II829_1 = (II547)|(II575);
assign II508 = ((~II509));
assign II1184_2 = (II269&II376);
assign II315 = ((~II272)&(~II514));
assign II655 = ((~II322)&(~II1077_1));
assign II1140_1 = (II271&II573);
assign II1040_1 = (OutputHS1&II322);
assign II333 = ((~II850_1)&(~II850_2));
assign II746 = ((~II1216_1))|((~II1216_2));
assign II318 = ((~II834_1))|((~II277));
assign II735 = ((~II552)&(~II1196_1));
assign II568 = ((~II1047_1))|((~II1047_2));
assign II479 = ((~II279))|((~II486));
assign II551 = ((~II279))|((~II442));
assign II21 = ((~II689))|((~II693))|((~II691));
assign II624 = ((~State_2)&(~II511));
assign II458 = ((~II279)&(~II571));
assign II1037_1 = (Prog_0)|(II336);
assign II489 = ((~II506))|((~II570));
assign II16 = ((~II323));
assign II446 = ((~II447));
assign II338 = ((~II857_1))|((~II439));
assign II770 = ((~II715))|((~II713));
assign II575 = ((~II271))|((~II284));
assign II1176_2 = (Prog_0&II600);
assign II596 = ((~II336)&(~II367));
assign II1151_1 = (II405)|(II537);
assign II485 = ((~II277))|((~II548));
assign II548 = ((~State_3)&(~II513));
assign II390 = ((~II391));
assign II12 = ((~II377))|((~II469));
assign II614 = ((~II523)&(~II575));
assign II691 = ((~II690));
assign II1199_1 = (II338&II364);
assign II398 = ((~II399));
assign II386 = ((~State_2)&(~II280));
assign II404 = ((~II284)&(~II421));
assign II1193_1 = (II424&II521);
assign II5 = ((~II733))|((~II729))|((~II731))|((~II397));
assign II376 = ((~II281)&(~II479));
assign II274 = ((~FullOHS1));
assign II545 = ((~II272))|((~II362));
assign II364 = ((~II274)&(~II379)&(~II525));
assign II562 = ((~II1037_1))|((~II439));
assign II282 = ((~Prog_2));
assign II475 = ((~II474));
assign II534 = ((~State_4)&(~II571));
assign II1132_2 = (II281)|(II467);
assign II1213_1 = (II498)|(II547);
assign II311 = ((~II742)&(~II746)&(~II744));
assign II329 = ((~II328));
assign II1216_1 = (II449)|(II537);
assign II1210_1 = (II339)|(II421);
assign II1113_1 = (II282)|(II415);
assign II410 = ((~II411));
assign II13 = ((~II415));
assign II450 = ((~State_0)&(~II505));
assign II697 = ((~II384)&(~II1140_1));
assign II423 = ((~II422));
assign II405 = ((~II404));
assign II275 = ((~FullIIHS1));
assign II580 = ((~II345)&(~II397));
assign II537 = ((~II263))|((~Rdy2RtHS1));
assign II1091_1 = (II585)|(II587);
assign II465 = ((~II390)&(~II966_1));
assign II559 = ((~II412)&(~II1031_1));
assign II449 = ((~State_1))|((~II318))|((~II450));
assign II30 = ((~II829_1))|((~II351));
assign II1107_1 = (II284&II382);
assign II24 = ((~OutAvHS1)&(~II326));
assign II740 = ((~II1207_1))|((~II477));
assign II711 = ((~II388)&(~II1160_1));
assign II359 = ((~Rdy1RtHS1))|((~II432))|((~II532));
assign II512 = ((~II280)&(~State_0));
assign II680 = ((~II445))|((~II381));
assign II442 = ((~State_1)&(~II347)&(~II509));
assign II554 = ((~II555));
assign II367 = ((~II366));
assign II416 = ((~II461)&(~II535));
assign II519 = ((~Rdy2BmHS1))|((~WantBmHS1));
assign II1188_1 = (State_1&II376);
assign II294 = ((~II408)&(~II678)&(~II676));
assign II370 = ((~II371));
assign II457 = ((~II266))|((~II506));
assign II723 = ((~II1180_1)&(~II1180_2));
assign II1188_2 = (II267&II388);
assign II414 = ((~State_1)&(~II425)&(~II521));
assign II264 = ((~Rdy2RtHS1));
assign II567 = ((~II388)&(~II1044_1));
assign II335 = ((~II277))|((~II282));
assign II673 = ((~II410)&(~II1107_1));
assign II354 = ((~II367)&(~II543));
assign II1148_1 = (II267)|(II565);
assign II267 = ((~IInDoneHS1));
assign II434 = ((~FullIIHS1)&(~II503));
assign II393 = ((~II282))|((~II283));
assign II1118_1 = (State_1)|(II479);
assign II461 = ((~II282))|((~II506));
assign II910_1 = (II277&II360);
assign II17 = ((~II294));
assign II660 = ((~II1087_1))|((~II469));
assign II342 = ((~II343));
assign II357 = ((~Rdy1BmHS1))|((~Rdy2BmHS1));
assign II665 = ((~II540)&(~II1094_1));
assign II539 = ((~II263))|((~II274));
assign II27 = ((~OutAvHS1)&(~II275));
assign II20 = ((~II297));
assign II702 = ((~II1148_1))|((~II481));
assign II1199_2 = (II267&II380);
assign II593 = ((~II284))|((~II430));
assign II377 = ((~II376));
assign II661 = ((~II660));
assign II394 = ((~State_0)&(~II327)&(~II357));
assign II494 = ((~II495));
assign II269 = ((~TpArrayHS1));
assign II657 = ((~II410)&(~II1080_1));
assign II547 = ((~WantRtHS1))|((~II446));
assign II535 = ((~II534));
assign II840_2 = (Prog_1&Prog_0);
assign II326 = ((~FullOHS1)&(~FullIIHS1));
assign II397 = ((~II396));
assign II1184_1 = (II486&II506);
assign II693 = ((~II376)&(~II1136_1));
assign II565 = ((~II444)&(~II1040_1));
assign II625 = ((~II624));
assign II896_1 = (II279)|(II320);
assign II676 = ((~II1113_1))|((~II343));
assign II767 = ((~II704)&(~II702));
assign II495 = ((~II280))|((~II281));
assign II733 = ((~II342)&(~II1193_1));
assign II7 = ((~II311));
assign II963_1 = (II335&II345);
assign II271 = ((~WantBmHS1));
assign II1110_1 = (II277&II388);
assign II322 = ((~II323));
assign II1034_1 = (II317&II428);
assign II451 = ((~II450));
assign II1121_1 = (State_0)|(II589);
assign II6 = ((~II377))|((~II779))|((~II777));
assign II486 = ((~II487));
assign II850_2 = (WantRtHS1&II614);
assign II525 = ((~II277))|((~II280));
assign II506 = ((~State_1)&(~II281));
assign II411 = ((~II279))|((~Prog_0))|((~II416));
assign II526 = ((~II370)&(~II416));
assign II10 = ((~II287));
assign II353 = ((~II344)&(~II873_1));
assign II445 = ((~II374))|((~II534));
assign II281 = ((~State_0));
assign II1203_1 = (II463)|(II491);
assign II325 = ((~II840_1)&(~II840_2));
assign II1103_1 = (State_5&II418);
assign II966_1 = (II335&II357);
assign II23 = ((~II300));
assign II561 = ((~II432)&(~II1034_1));
assign II14 = ((~II671))|((~II673));
assign II430 = ((~Prog_2)&(~II451));
assign II690 = ((~II1132_1))|((~II1132_2));
assign II491 = ((~State_5))|((~II548));
assign II396 = ((~II280)&(~II425));
assign II276 = ((~State_5));
assign II529 = ((~II399))|((~II489));
assign II1056_1 = (II280&II358);
assign II1180_2 = (II348&II554);
assign II403 = ((~II634))|((~II434))|((~II494));
assign II706 = ((~II1154_1))|((~II403));
assign II684 = ((~II1121_1))|((~II1121_2));
assign II380 = ((~II381));
assign II873_1 = (II263&II264);
assign II814_1 = (FullOHS1)|(II355);
assign II424 = ((~II425));
assign II295 = ((~II376)&(~II682)&(~II680));
assign II553 = ((~State_1))|((~II500));
assign II1166_1 = (II357&II529);
assign II738 = ((~II1203_1))|((~II1203_2));
assign II468 = ((~State_0)&(~II386)&(~II487));
assign II717 = ((~II322)&(~II1170_1));
assign II287 = ((~II750)&(~II789_1));
assign II341 = ((~II340));
assign II360 = ((~II881_1))|((~II881_2));
assign II350 = ((~II325)&(~II477));
assign II881_2 = (II282)|(II326);
assign II330 = ((~WantBmHS1))|((~II493));
assign II345 = ((~Rdy1RtHS1))|((~Rdy2RtHS1));
assign II374 = ((~II896_1))|((~II461));
assign II1180_1 = (II267&II322);
assign II505 = ((~II279))|((~II570));
assign II435 = ((~II434));
assign II1094_1 = (WantRtHS1&II582);
assign II284 = ((~Prog_0));
assign II1121_2 = (Rdy2BmHS1)|(II559);
assign II861_2 = (II265)|(II457);
assign II881_1 = (IInDoneHS1)|(Prog_2);
assign II470 = ((~II320)&(~II335)&(~II571));
assign II573 = ((~II517))|((~II545));
assign II857_1 = (Prog_0)|(II493);
assign II1100_1 = (WantBmHS1&II384);
assign II331 = ((~II330));
assign II500 = ((~II281)&(~II453));
assign II1047_2 = (Rdy1BmHS1)|(Prog_0);
assign II744 = ((~II1213_1))|((~II553));
assign II1087_1 = (Prog_0)|(II526);
assign II667 = ((~II328)&(~II1097_1));
assign II11 = ((~II475))|((~II669))|((~II667));
assign II610 = ((~Prog_2)&(~II284));
assign II1025_1 = (Rdy2BmHS1&II325);
assign II729 = ((~II1188_1)&(~II1188_2));
assign II675 = ((~II470)&(~II1110_1));
assign II371 = ((~II279))|((~II382));
assign II303 = ((~II706)&(~II708));
assign II552 = ((~II553));
assign II327 = ((~II326));
assign II384 = ((~II315)&(~II407)&(~II493));
assign II358 = ((~II359));
assign II381 = ((~State_3))|((~II396));
assign II388 = ((~II320)&(~II459));
assign II320 = ((~II495))|((~II511));
assign II721 = ((~II1176_1)&(~II1176_2));
assign II1132_1 = (II593)|(II595);
assign II850_1 = (II610&II612);
assign II477 = ((~II476));
assign II1203_2 = (II543)|(II577);
assign II408 = ((~II341)&(~II435)&(~II523));
assign II323 = ((~State_4))|((~II281))|((~II436));
assign II452 = ((~II453));
assign II566 = ((~II567));
assign II1216_2 = (II465)|(II489);
assign II272 = ((~WantRtHS1));
assign II277 = ((~State_4));
assign II421 = ((~II274))|((~II422));
assign II540 = ((~Rdy2RtHS1)&(~II263)&(~II449));
assign II634 = ((~II264)&(~II333));
assign II600 = ((~II331)&(~II447));
assign II441 = ((~II440));
assign II2 = ((~II711))|((~II771))|((~II769));
assign II429 = ((~Prog_0))|((~II450));
assign II778 = ((~II737))|((~II735));
assign II708 = ((~II1157_1))|((~II351));
assign II317 = ((~FullOHS1))|((~FullIIHS1));
assign II590 = ((~II429)&(~II539));
assign II570 = ((~II276)&(~State_3));
assign II412 = ((~II282)&(~II437));
assign II612 = ((~Rdy1RtHS1)&(~II274));
assign II737 = ((~II1199_1)&(~II1199_2));
assign II1170_1 = (II393&II414);
assign II834_1 = (FullIIHS1)|(II523);
assign II719 = ((~II500)&(~II1173_1));
assign II459 = ((~II458));
assign II1128_1 = (II378&II568);
assign II455 = ((~II264))|((~II512));
assign II19 = ((~II371))|((~II323));
assign II467 = ((~II466));
assign II579 = ((~II446)&(~II1056_1));
assign II428 = ((~II429));
assign II1176_1 = (State_4&II566);
assign II713 = ((~II470)&(~II1163_1));
assign II391 = ((~State_2)&(~II910_1));
assign II582 = ((~II331)&(~II517));
assign II26 = ((~II303));
assign II340 = ((~II861_1))|((~II861_2));
assign II1097_1 = (II317&II556);
assign II669 = ((~II342)&(~II1100_1));
assign II280 = ((~State_1));
assign II662 = ((~II1091_1))|((~II329));
assign II463 = ((~II390)&(~II963_1));
assign II453 = ((~II277))|((~II327))|((~II504));
assign II742 = ((~II1210_1))|((~II551));
assign II769 = ((~II768));
assign II777 = ((~II740)&(~II738));
assign II700 = ((~II403))|((~II351));
assign II432 = ((~II282)&(~II451));
assign II589 = ((~Prog_2))|((~II482));
assign II344 = ((~II345));
assign II265 = ((~Rdy1BmHS1));
assign II482 = ((~State_3)&(~State_2)&(~II525));
assign II22 = ((~II699))|((~II695))|((~II697))|((~II481));
assign II678 = ((~II329))|((~II423));
assign II28 = ((~OutAvHS1)&(~FullIIHS1));
assign II436 = ((~State_1)&(~II505));
assign II473 = ((~II265))|((~II266));
assign II3 = ((~II721))|((~II723));
assign II444 = ((~II445));
assign II1143_2 = (II274&II596);
assign II892_1 = (II279)|(II495);
assign II378 = ((~FullIIHS1)&(~II431));
endmodule
