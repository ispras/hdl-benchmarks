//NOTE: no-implementation module stub

module REG16L (
    input wire DSPCLK,
    input wire CLKMX0renb,
    input wire GO_C,
    input wire [15:0] Xin,
    output reg [15:0] MX0r
);

endmodule
