//NOTE: no-implementation module stub

module REG12LC (
    input wire DSPCLK,
    input wire MMR_web,
    input wire PMASK_we,
    input wire [15:0] DMD,
    output reg [11:0] PMASK,
    input wire T_RST
);

endmodule
