module OptKuznechikDecoder(
  input wire clk,
  input wire [127:0] encoded,
  input wire [255:0] key,
  output wire [127:0] out
);
  wire [7:0] literal_2043896[256] = '{8'hfc, 8'hee, 8'hdd, 8'h11, 8'hcf, 8'h6e, 8'h31, 8'h16, 8'hfb, 8'hc4, 8'hfa, 8'hda, 8'h23, 8'hc5, 8'h04, 8'h4d, 8'he9, 8'h77, 8'hf0, 8'hdb, 8'h93, 8'h2e, 8'h99, 8'hba, 8'h17, 8'h36, 8'hf1, 8'hbb, 8'h14, 8'hcd, 8'h5f, 8'hc1, 8'hf9, 8'h18, 8'h65, 8'h5a, 8'he2, 8'h5c, 8'hef, 8'h21, 8'h81, 8'h1c, 8'h3c, 8'h42, 8'h8b, 8'h01, 8'h8e, 8'h4f, 8'h05, 8'h84, 8'h02, 8'hae, 8'he3, 8'h6a, 8'h8f, 8'ha0, 8'h06, 8'h0b, 8'hed, 8'h98, 8'h7f, 8'hd4, 8'hd3, 8'h1f, 8'heb, 8'h34, 8'h2c, 8'h51, 8'hea, 8'hc8, 8'h48, 8'hab, 8'hf2, 8'h2a, 8'h68, 8'ha2, 8'hfd, 8'h3a, 8'hce, 8'hcc, 8'hb5, 8'h70, 8'h0e, 8'h56, 8'h08, 8'h0c, 8'h76, 8'h12, 8'hbf, 8'h72, 8'h13, 8'h47, 8'h9c, 8'hb7, 8'h5d, 8'h87, 8'h15, 8'ha1, 8'h96, 8'h29, 8'h10, 8'h7b, 8'h9a, 8'hc7, 8'hf3, 8'h91, 8'h78, 8'h6f, 8'h9d, 8'h9e, 8'hb2, 8'hb1, 8'h32, 8'h75, 8'h19, 8'h3d, 8'hff, 8'h35, 8'h8a, 8'h7e, 8'h6d, 8'h54, 8'hc6, 8'h80, 8'hc3, 8'hbd, 8'h0d, 8'h57, 8'hdf, 8'hf5, 8'h24, 8'ha9, 8'h3e, 8'ha8, 8'h43, 8'hc9, 8'hd7, 8'h79, 8'hd6, 8'hf6, 8'h7c, 8'h22, 8'hb9, 8'h03, 8'he0, 8'h0f, 8'hec, 8'hde, 8'h7a, 8'h94, 8'hb0, 8'hbc, 8'hdc, 8'he8, 8'h28, 8'h50, 8'h4e, 8'h33, 8'h0a, 8'h4a, 8'ha7, 8'h97, 8'h60, 8'h73, 8'h1e, 8'h00, 8'h62, 8'h44, 8'h1a, 8'hb8, 8'h38, 8'h82, 8'h64, 8'h9f, 8'h26, 8'h41, 8'had, 8'h45, 8'h46, 8'h92, 8'h27, 8'h5e, 8'h55, 8'h2f, 8'h8c, 8'ha3, 8'ha5, 8'h7d, 8'h69, 8'hd5, 8'h95, 8'h3b, 8'h07, 8'h58, 8'hb3, 8'h40, 8'h86, 8'hac, 8'h1d, 8'hf7, 8'h30, 8'h37, 8'h6b, 8'he4, 8'h88, 8'hd9, 8'he7, 8'h89, 8'he1, 8'h1b, 8'h83, 8'h49, 8'h4c, 8'h3f, 8'hf8, 8'hfe, 8'h8d, 8'h53, 8'haa, 8'h90, 8'hca, 8'hd8, 8'h85, 8'h61, 8'h20, 8'h71, 8'h67, 8'ha4, 8'h2d, 8'h2b, 8'h09, 8'h5b, 8'hcb, 8'h9b, 8'h25, 8'hd0, 8'hbe, 8'he5, 8'h6c, 8'h52, 8'h59, 8'ha6, 8'h74, 8'hd2, 8'he6, 8'hf4, 8'hb4, 8'hc0, 8'hd1, 8'h66, 8'haf, 8'hc2, 8'h39, 8'h4b, 8'h63, 8'hb6};
  wire [7:0] literal_2043910[256] = '{8'h00, 8'h94, 8'heb, 8'h7f, 8'h15, 8'h81, 8'hfe, 8'h6a, 8'h2a, 8'hbe, 8'hc1, 8'h55, 8'h3f, 8'hab, 8'hd4, 8'h40, 8'h54, 8'hc0, 8'hbf, 8'h2b, 8'h41, 8'hd5, 8'haa, 8'h3e, 8'h7e, 8'hea, 8'h95, 8'h01, 8'h6b, 8'hff, 8'h80, 8'h14, 8'ha8, 8'h3c, 8'h43, 8'hd7, 8'hbd, 8'h29, 8'h56, 8'hc2, 8'h82, 8'h16, 8'h69, 8'hfd, 8'h97, 8'h03, 8'h7c, 8'he8, 8'hfc, 8'h68, 8'h17, 8'h83, 8'he9, 8'h7d, 8'h02, 8'h96, 8'hd6, 8'h42, 8'h3d, 8'ha9, 8'hc3, 8'h57, 8'h28, 8'hbc, 8'h93, 8'h07, 8'h78, 8'hec, 8'h86, 8'h12, 8'h6d, 8'hf9, 8'hb9, 8'h2d, 8'h52, 8'hc6, 8'hac, 8'h38, 8'h47, 8'hd3, 8'hc7, 8'h53, 8'h2c, 8'hb8, 8'hd2, 8'h46, 8'h39, 8'had, 8'hed, 8'h79, 8'h06, 8'h92, 8'hf8, 8'h6c, 8'h13, 8'h87, 8'h3b, 8'haf, 8'hd0, 8'h44, 8'h2e, 8'hba, 8'hc5, 8'h51, 8'h11, 8'h85, 8'hfa, 8'h6e, 8'h04, 8'h90, 8'hef, 8'h7b, 8'h6f, 8'hfb, 8'h84, 8'h10, 8'h7a, 8'hee, 8'h91, 8'h05, 8'h45, 8'hd1, 8'hae, 8'h3a, 8'h50, 8'hc4, 8'hbb, 8'h2f, 8'he5, 8'h71, 8'h0e, 8'h9a, 8'hf0, 8'h64, 8'h1b, 8'h8f, 8'hcf, 8'h5b, 8'h24, 8'hb0, 8'hda, 8'h4e, 8'h31, 8'ha5, 8'hb1, 8'h25, 8'h5a, 8'hce, 8'ha4, 8'h30, 8'h4f, 8'hdb, 8'h9b, 8'h0f, 8'h70, 8'he4, 8'h8e, 8'h1a, 8'h65, 8'hf1, 8'h4d, 8'hd9, 8'ha6, 8'h32, 8'h58, 8'hcc, 8'hb3, 8'h27, 8'h67, 8'hf3, 8'h8c, 8'h18, 8'h72, 8'he6, 8'h99, 8'h0d, 8'h19, 8'h8d, 8'hf2, 8'h66, 8'h0c, 8'h98, 8'he7, 8'h73, 8'h33, 8'ha7, 8'hd8, 8'h4c, 8'h26, 8'hb2, 8'hcd, 8'h59, 8'h76, 8'he2, 8'h9d, 8'h09, 8'h63, 8'hf7, 8'h88, 8'h1c, 8'h5c, 8'hc8, 8'hb7, 8'h23, 8'h49, 8'hdd, 8'ha2, 8'h36, 8'h22, 8'hb6, 8'hc9, 8'h5d, 8'h37, 8'ha3, 8'hdc, 8'h48, 8'h08, 8'h9c, 8'he3, 8'h77, 8'h1d, 8'h89, 8'hf6, 8'h62, 8'hde, 8'h4a, 8'h35, 8'ha1, 8'hcb, 8'h5f, 8'h20, 8'hb4, 8'hf4, 8'h60, 8'h1f, 8'h8b, 8'he1, 8'h75, 8'h0a, 8'h9e, 8'h8a, 8'h1e, 8'h61, 8'hf5, 8'h9f, 8'h0b, 8'h74, 8'he0, 8'ha0, 8'h34, 8'h4b, 8'hdf, 8'hb5, 8'h21, 8'h5e, 8'hca};
  wire [7:0] literal_2043912[256] = '{8'h00, 8'h20, 8'h40, 8'h60, 8'h80, 8'ha0, 8'hc0, 8'he0, 8'hc3, 8'he3, 8'h83, 8'ha3, 8'h43, 8'h63, 8'h03, 8'h23, 8'h45, 8'h65, 8'h05, 8'h25, 8'hc5, 8'he5, 8'h85, 8'ha5, 8'h86, 8'ha6, 8'hc6, 8'he6, 8'h06, 8'h26, 8'h46, 8'h66, 8'h8a, 8'haa, 8'hca, 8'hea, 8'h0a, 8'h2a, 8'h4a, 8'h6a, 8'h49, 8'h69, 8'h09, 8'h29, 8'hc9, 8'he9, 8'h89, 8'ha9, 8'hcf, 8'hef, 8'h8f, 8'haf, 8'h4f, 8'h6f, 8'h0f, 8'h2f, 8'h0c, 8'h2c, 8'h4c, 8'h6c, 8'h8c, 8'hac, 8'hcc, 8'hec, 8'hd7, 8'hf7, 8'h97, 8'hb7, 8'h57, 8'h77, 8'h17, 8'h37, 8'h14, 8'h34, 8'h54, 8'h74, 8'h94, 8'hb4, 8'hd4, 8'hf4, 8'h92, 8'hb2, 8'hd2, 8'hf2, 8'h12, 8'h32, 8'h52, 8'h72, 8'h51, 8'h71, 8'h11, 8'h31, 8'hd1, 8'hf1, 8'h91, 8'hb1, 8'h5d, 8'h7d, 8'h1d, 8'h3d, 8'hdd, 8'hfd, 8'h9d, 8'hbd, 8'h9e, 8'hbe, 8'hde, 8'hfe, 8'h1e, 8'h3e, 8'h5e, 8'h7e, 8'h18, 8'h38, 8'h58, 8'h78, 8'h98, 8'hb8, 8'hd8, 8'hf8, 8'hdb, 8'hfb, 8'h9b, 8'hbb, 8'h5b, 8'h7b, 8'h1b, 8'h3b, 8'h6d, 8'h4d, 8'h2d, 8'h0d, 8'hed, 8'hcd, 8'had, 8'h8d, 8'hae, 8'h8e, 8'hee, 8'hce, 8'h2e, 8'h0e, 8'h6e, 8'h4e, 8'h28, 8'h08, 8'h68, 8'h48, 8'ha8, 8'h88, 8'he8, 8'hc8, 8'heb, 8'hcb, 8'hab, 8'h8b, 8'h6b, 8'h4b, 8'h2b, 8'h0b, 8'he7, 8'hc7, 8'ha7, 8'h87, 8'h67, 8'h47, 8'h27, 8'h07, 8'h24, 8'h04, 8'h64, 8'h44, 8'ha4, 8'h84, 8'he4, 8'hc4, 8'ha2, 8'h82, 8'he2, 8'hc2, 8'h22, 8'h02, 8'h62, 8'h42, 8'h61, 8'h41, 8'h21, 8'h01, 8'he1, 8'hc1, 8'ha1, 8'h81, 8'hba, 8'h9a, 8'hfa, 8'hda, 8'h3a, 8'h1a, 8'h7a, 8'h5a, 8'h79, 8'h59, 8'h39, 8'h19, 8'hf9, 8'hd9, 8'hb9, 8'h99, 8'hff, 8'hdf, 8'hbf, 8'h9f, 8'h7f, 8'h5f, 8'h3f, 8'h1f, 8'h3c, 8'h1c, 8'h7c, 8'h5c, 8'hbc, 8'h9c, 8'hfc, 8'hdc, 8'h30, 8'h10, 8'h70, 8'h50, 8'hb0, 8'h90, 8'hf0, 8'hd0, 8'hf3, 8'hd3, 8'hb3, 8'h93, 8'h73, 8'h53, 8'h33, 8'h13, 8'h75, 8'h55, 8'h35, 8'h15, 8'hf5, 8'hd5, 8'hb5, 8'h95, 8'hb6, 8'h96, 8'hf6, 8'hd6, 8'h36, 8'h16, 8'h76, 8'h56};
  wire [7:0] literal_2043914[256] = '{8'h00, 8'h85, 8'hc9, 8'h4c, 8'h51, 8'hd4, 8'h98, 8'h1d, 8'ha2, 8'h27, 8'h6b, 8'hee, 8'hf3, 8'h76, 8'h3a, 8'hbf, 8'h87, 8'h02, 8'h4e, 8'hcb, 8'hd6, 8'h53, 8'h1f, 8'h9a, 8'h25, 8'ha0, 8'hec, 8'h69, 8'h74, 8'hf1, 8'hbd, 8'h38, 8'hcd, 8'h48, 8'h04, 8'h81, 8'h9c, 8'h19, 8'h55, 8'hd0, 8'h6f, 8'hea, 8'ha6, 8'h23, 8'h3e, 8'hbb, 8'hf7, 8'h72, 8'h4a, 8'hcf, 8'h83, 8'h06, 8'h1b, 8'h9e, 8'hd2, 8'h57, 8'he8, 8'h6d, 8'h21, 8'ha4, 8'hb9, 8'h3c, 8'h70, 8'hf5, 8'h59, 8'hdc, 8'h90, 8'h15, 8'h08, 8'h8d, 8'hc1, 8'h44, 8'hfb, 8'h7e, 8'h32, 8'hb7, 8'haa, 8'h2f, 8'h63, 8'he6, 8'hde, 8'h5b, 8'h17, 8'h92, 8'h8f, 8'h0a, 8'h46, 8'hc3, 8'h7c, 8'hf9, 8'hb5, 8'h30, 8'h2d, 8'ha8, 8'he4, 8'h61, 8'h94, 8'h11, 8'h5d, 8'hd8, 8'hc5, 8'h40, 8'h0c, 8'h89, 8'h36, 8'hb3, 8'hff, 8'h7a, 8'h67, 8'he2, 8'hae, 8'h2b, 8'h13, 8'h96, 8'hda, 8'h5f, 8'h42, 8'hc7, 8'h8b, 8'h0e, 8'hb1, 8'h34, 8'h78, 8'hfd, 8'he0, 8'h65, 8'h29, 8'hac, 8'hb2, 8'h37, 8'h7b, 8'hfe, 8'he3, 8'h66, 8'h2a, 8'haf, 8'h10, 8'h95, 8'hd9, 8'h5c, 8'h41, 8'hc4, 8'h88, 8'h0d, 8'h35, 8'hb0, 8'hfc, 8'h79, 8'h64, 8'he1, 8'had, 8'h28, 8'h97, 8'h12, 8'h5e, 8'hdb, 8'hc6, 8'h43, 8'h0f, 8'h8a, 8'h7f, 8'hfa, 8'hb6, 8'h33, 8'h2e, 8'hab, 8'he7, 8'h62, 8'hdd, 8'h58, 8'h14, 8'h91, 8'h8c, 8'h09, 8'h45, 8'hc0, 8'hf8, 8'h7d, 8'h31, 8'hb4, 8'ha9, 8'h2c, 8'h60, 8'he5, 8'h5a, 8'hdf, 8'h93, 8'h16, 8'h0b, 8'h8e, 8'hc2, 8'h47, 8'heb, 8'h6e, 8'h22, 8'ha7, 8'hba, 8'h3f, 8'h73, 8'hf6, 8'h49, 8'hcc, 8'h80, 8'h05, 8'h18, 8'h9d, 8'hd1, 8'h54, 8'h6c, 8'he9, 8'ha5, 8'h20, 8'h3d, 8'hb8, 8'hf4, 8'h71, 8'hce, 8'h4b, 8'h07, 8'h82, 8'h9f, 8'h1a, 8'h56, 8'hd3, 8'h26, 8'ha3, 8'hef, 8'h6a, 8'h77, 8'hf2, 8'hbe, 8'h3b, 8'h84, 8'h01, 8'h4d, 8'hc8, 8'hd5, 8'h50, 8'h1c, 8'h99, 8'ha1, 8'h24, 8'h68, 8'hed, 8'hf0, 8'h75, 8'h39, 8'hbc, 8'h03, 8'h86, 8'hca, 8'h4f, 8'h52, 8'hd7, 8'h9b, 8'h1e};
  wire [7:0] literal_2043916[256] = '{8'h00, 8'h10, 8'h20, 8'h30, 8'h40, 8'h50, 8'h60, 8'h70, 8'h80, 8'h90, 8'ha0, 8'hb0, 8'hc0, 8'hd0, 8'he0, 8'hf0, 8'hc3, 8'hd3, 8'he3, 8'hf3, 8'h83, 8'h93, 8'ha3, 8'hb3, 8'h43, 8'h53, 8'h63, 8'h73, 8'h03, 8'h13, 8'h23, 8'h33, 8'h45, 8'h55, 8'h65, 8'h75, 8'h05, 8'h15, 8'h25, 8'h35, 8'hc5, 8'hd5, 8'he5, 8'hf5, 8'h85, 8'h95, 8'ha5, 8'hb5, 8'h86, 8'h96, 8'ha6, 8'hb6, 8'hc6, 8'hd6, 8'he6, 8'hf6, 8'h06, 8'h16, 8'h26, 8'h36, 8'h46, 8'h56, 8'h66, 8'h76, 8'h8a, 8'h9a, 8'haa, 8'hba, 8'hca, 8'hda, 8'hea, 8'hfa, 8'h0a, 8'h1a, 8'h2a, 8'h3a, 8'h4a, 8'h5a, 8'h6a, 8'h7a, 8'h49, 8'h59, 8'h69, 8'h79, 8'h09, 8'h19, 8'h29, 8'h39, 8'hc9, 8'hd9, 8'he9, 8'hf9, 8'h89, 8'h99, 8'ha9, 8'hb9, 8'hcf, 8'hdf, 8'hef, 8'hff, 8'h8f, 8'h9f, 8'haf, 8'hbf, 8'h4f, 8'h5f, 8'h6f, 8'h7f, 8'h0f, 8'h1f, 8'h2f, 8'h3f, 8'h0c, 8'h1c, 8'h2c, 8'h3c, 8'h4c, 8'h5c, 8'h6c, 8'h7c, 8'h8c, 8'h9c, 8'hac, 8'hbc, 8'hcc, 8'hdc, 8'hec, 8'hfc, 8'hd7, 8'hc7, 8'hf7, 8'he7, 8'h97, 8'h87, 8'hb7, 8'ha7, 8'h57, 8'h47, 8'h77, 8'h67, 8'h17, 8'h07, 8'h37, 8'h27, 8'h14, 8'h04, 8'h34, 8'h24, 8'h54, 8'h44, 8'h74, 8'h64, 8'h94, 8'h84, 8'hb4, 8'ha4, 8'hd4, 8'hc4, 8'hf4, 8'he4, 8'h92, 8'h82, 8'hb2, 8'ha2, 8'hd2, 8'hc2, 8'hf2, 8'he2, 8'h12, 8'h02, 8'h32, 8'h22, 8'h52, 8'h42, 8'h72, 8'h62, 8'h51, 8'h41, 8'h71, 8'h61, 8'h11, 8'h01, 8'h31, 8'h21, 8'hd1, 8'hc1, 8'hf1, 8'he1, 8'h91, 8'h81, 8'hb1, 8'ha1, 8'h5d, 8'h4d, 8'h7d, 8'h6d, 8'h1d, 8'h0d, 8'h3d, 8'h2d, 8'hdd, 8'hcd, 8'hfd, 8'hed, 8'h9d, 8'h8d, 8'hbd, 8'had, 8'h9e, 8'h8e, 8'hbe, 8'hae, 8'hde, 8'hce, 8'hfe, 8'hee, 8'h1e, 8'h0e, 8'h3e, 8'h2e, 8'h5e, 8'h4e, 8'h7e, 8'h6e, 8'h18, 8'h08, 8'h38, 8'h28, 8'h58, 8'h48, 8'h78, 8'h68, 8'h98, 8'h88, 8'hb8, 8'ha8, 8'hd8, 8'hc8, 8'hf8, 8'he8, 8'hdb, 8'hcb, 8'hfb, 8'heb, 8'h9b, 8'h8b, 8'hbb, 8'hab, 8'h5b, 8'h4b, 8'h7b, 8'h6b, 8'h1b, 8'h0b, 8'h3b, 8'h2b};
  wire [7:0] literal_2043918[256] = '{8'h00, 8'hc2, 8'h47, 8'h85, 8'h8e, 8'h4c, 8'hc9, 8'h0b, 8'hdf, 8'h1d, 8'h98, 8'h5a, 8'h51, 8'h93, 8'h16, 8'hd4, 8'h7d, 8'hbf, 8'h3a, 8'hf8, 8'hf3, 8'h31, 8'hb4, 8'h76, 8'ha2, 8'h60, 8'he5, 8'h27, 8'h2c, 8'hee, 8'h6b, 8'ha9, 8'hfa, 8'h38, 8'hbd, 8'h7f, 8'h74, 8'hb6, 8'h33, 8'hf1, 8'h25, 8'he7, 8'h62, 8'ha0, 8'hab, 8'h69, 8'hec, 8'h2e, 8'h87, 8'h45, 8'hc0, 8'h02, 8'h09, 8'hcb, 8'h4e, 8'h8c, 8'h58, 8'h9a, 8'h1f, 8'hdd, 8'hd6, 8'h14, 8'h91, 8'h53, 8'h37, 8'hf5, 8'h70, 8'hb2, 8'hb9, 8'h7b, 8'hfe, 8'h3c, 8'he8, 8'h2a, 8'haf, 8'h6d, 8'h66, 8'ha4, 8'h21, 8'he3, 8'h4a, 8'h88, 8'h0d, 8'hcf, 8'hc4, 8'h06, 8'h83, 8'h41, 8'h95, 8'h57, 8'hd2, 8'h10, 8'h1b, 8'hd9, 8'h5c, 8'h9e, 8'hcd, 8'h0f, 8'h8a, 8'h48, 8'h43, 8'h81, 8'h04, 8'hc6, 8'h12, 8'hd0, 8'h55, 8'h97, 8'h9c, 8'h5e, 8'hdb, 8'h19, 8'hb0, 8'h72, 8'hf7, 8'h35, 8'h3e, 8'hfc, 8'h79, 8'hbb, 8'h6f, 8'had, 8'h28, 8'hea, 8'he1, 8'h23, 8'ha6, 8'h64, 8'h6e, 8'hac, 8'h29, 8'heb, 8'he0, 8'h22, 8'ha7, 8'h65, 8'hb1, 8'h73, 8'hf6, 8'h34, 8'h3f, 8'hfd, 8'h78, 8'hba, 8'h13, 8'hd1, 8'h54, 8'h96, 8'h9d, 8'h5f, 8'hda, 8'h18, 8'hcc, 8'h0e, 8'h8b, 8'h49, 8'h42, 8'h80, 8'h05, 8'hc7, 8'h94, 8'h56, 8'hd3, 8'h11, 8'h1a, 8'hd8, 8'h5d, 8'h9f, 8'h4b, 8'h89, 8'h0c, 8'hce, 8'hc5, 8'h07, 8'h82, 8'h40, 8'he9, 8'h2b, 8'hae, 8'h6c, 8'h67, 8'ha5, 8'h20, 8'he2, 8'h36, 8'hf4, 8'h71, 8'hb3, 8'hb8, 8'h7a, 8'hff, 8'h3d, 8'h59, 8'h9b, 8'h1e, 8'hdc, 8'hd7, 8'h15, 8'h90, 8'h52, 8'h86, 8'h44, 8'hc1, 8'h03, 8'h08, 8'hca, 8'h4f, 8'h8d, 8'h24, 8'he6, 8'h63, 8'ha1, 8'haa, 8'h68, 8'hed, 8'h2f, 8'hfb, 8'h39, 8'hbc, 8'h7e, 8'h75, 8'hb7, 8'h32, 8'hf0, 8'ha3, 8'h61, 8'he4, 8'h26, 8'h2d, 8'hef, 8'h6a, 8'ha8, 8'h7c, 8'hbe, 8'h3b, 8'hf9, 8'hf2, 8'h30, 8'hb5, 8'h77, 8'hde, 8'h1c, 8'h99, 8'h5b, 8'h50, 8'h92, 8'h17, 8'hd5, 8'h01, 8'hc3, 8'h46, 8'h84, 8'h8f, 8'h4d, 8'hc8, 8'h0a};
  wire [7:0] literal_2043920[256] = '{8'h00, 8'hc0, 8'h43, 8'h83, 8'h86, 8'h46, 8'hc5, 8'h05, 8'hcf, 8'h0f, 8'h8c, 8'h4c, 8'h49, 8'h89, 8'h0a, 8'hca, 8'h5d, 8'h9d, 8'h1e, 8'hde, 8'hdb, 8'h1b, 8'h98, 8'h58, 8'h92, 8'h52, 8'hd1, 8'h11, 8'h14, 8'hd4, 8'h57, 8'h97, 8'hba, 8'h7a, 8'hf9, 8'h39, 8'h3c, 8'hfc, 8'h7f, 8'hbf, 8'h75, 8'hb5, 8'h36, 8'hf6, 8'hf3, 8'h33, 8'hb0, 8'h70, 8'he7, 8'h27, 8'ha4, 8'h64, 8'h61, 8'ha1, 8'h22, 8'he2, 8'h28, 8'he8, 8'h6b, 8'hab, 8'hae, 8'h6e, 8'hed, 8'h2d, 8'hb7, 8'h77, 8'hf4, 8'h34, 8'h31, 8'hf1, 8'h72, 8'hb2, 8'h78, 8'hb8, 8'h3b, 8'hfb, 8'hfe, 8'h3e, 8'hbd, 8'h7d, 8'hea, 8'h2a, 8'ha9, 8'h69, 8'h6c, 8'hac, 8'h2f, 8'hef, 8'h25, 8'he5, 8'h66, 8'ha6, 8'ha3, 8'h63, 8'he0, 8'h20, 8'h0d, 8'hcd, 8'h4e, 8'h8e, 8'h8b, 8'h4b, 8'hc8, 8'h08, 8'hc2, 8'h02, 8'h81, 8'h41, 8'h44, 8'h84, 8'h07, 8'hc7, 8'h50, 8'h90, 8'h13, 8'hd3, 8'hd6, 8'h16, 8'h95, 8'h55, 8'h9f, 8'h5f, 8'hdc, 8'h1c, 8'h19, 8'hd9, 8'h5a, 8'h9a, 8'had, 8'h6d, 8'hee, 8'h2e, 8'h2b, 8'heb, 8'h68, 8'ha8, 8'h62, 8'ha2, 8'h21, 8'he1, 8'he4, 8'h24, 8'ha7, 8'h67, 8'hf0, 8'h30, 8'hb3, 8'h73, 8'h76, 8'hb6, 8'h35, 8'hf5, 8'h3f, 8'hff, 8'h7c, 8'hbc, 8'hb9, 8'h79, 8'hfa, 8'h3a, 8'h17, 8'hd7, 8'h54, 8'h94, 8'h91, 8'h51, 8'hd2, 8'h12, 8'hd8, 8'h18, 8'h9b, 8'h5b, 8'h5e, 8'h9e, 8'h1d, 8'hdd, 8'h4a, 8'h8a, 8'h09, 8'hc9, 8'hcc, 8'h0c, 8'h8f, 8'h4f, 8'h85, 8'h45, 8'hc6, 8'h06, 8'h03, 8'hc3, 8'h40, 8'h80, 8'h1a, 8'hda, 8'h59, 8'h99, 8'h9c, 8'h5c, 8'hdf, 8'h1f, 8'hd5, 8'h15, 8'h96, 8'h56, 8'h53, 8'h93, 8'h10, 8'hd0, 8'h47, 8'h87, 8'h04, 8'hc4, 8'hc1, 8'h01, 8'h82, 8'h42, 8'h88, 8'h48, 8'hcb, 8'h0b, 8'h0e, 8'hce, 8'h4d, 8'h8d, 8'ha0, 8'h60, 8'he3, 8'h23, 8'h26, 8'he6, 8'h65, 8'ha5, 8'h6f, 8'haf, 8'h2c, 8'hec, 8'he9, 8'h29, 8'haa, 8'h6a, 8'hfd, 8'h3d, 8'hbe, 8'h7e, 8'h7b, 8'hbb, 8'h38, 8'hf8, 8'h32, 8'hf2, 8'h71, 8'hb1, 8'hb4, 8'h74, 8'hf7, 8'h37};
  wire [7:0] literal_2043923[256] = '{8'h00, 8'hfb, 8'h35, 8'hce, 8'h6a, 8'h91, 8'h5f, 8'ha4, 8'hd4, 8'h2f, 8'he1, 8'h1a, 8'hbe, 8'h45, 8'h8b, 8'h70, 8'h6b, 8'h90, 8'h5e, 8'ha5, 8'h01, 8'hfa, 8'h34, 8'hcf, 8'hbf, 8'h44, 8'h8a, 8'h71, 8'hd5, 8'h2e, 8'he0, 8'h1b, 8'hd6, 8'h2d, 8'he3, 8'h18, 8'hbc, 8'h47, 8'h89, 8'h72, 8'h02, 8'hf9, 8'h37, 8'hcc, 8'h68, 8'h93, 8'h5d, 8'ha6, 8'hbd, 8'h46, 8'h88, 8'h73, 8'hd7, 8'h2c, 8'he2, 8'h19, 8'h69, 8'h92, 8'h5c, 8'ha7, 8'h03, 8'hf8, 8'h36, 8'hcd, 8'h6f, 8'h94, 8'h5a, 8'ha1, 8'h05, 8'hfe, 8'h30, 8'hcb, 8'hbb, 8'h40, 8'h8e, 8'h75, 8'hd1, 8'h2a, 8'he4, 8'h1f, 8'h04, 8'hff, 8'h31, 8'hca, 8'h6e, 8'h95, 8'h5b, 8'ha0, 8'hd0, 8'h2b, 8'he5, 8'h1e, 8'hba, 8'h41, 8'h8f, 8'h74, 8'hb9, 8'h42, 8'h8c, 8'h77, 8'hd3, 8'h28, 8'he6, 8'h1d, 8'h6d, 8'h96, 8'h58, 8'ha3, 8'h07, 8'hfc, 8'h32, 8'hc9, 8'hd2, 8'h29, 8'he7, 8'h1c, 8'hb8, 8'h43, 8'h8d, 8'h76, 8'h06, 8'hfd, 8'h33, 8'hc8, 8'h6c, 8'h97, 8'h59, 8'ha2, 8'hde, 8'h25, 8'heb, 8'h10, 8'hb4, 8'h4f, 8'h81, 8'h7a, 8'h0a, 8'hf1, 8'h3f, 8'hc4, 8'h60, 8'h9b, 8'h55, 8'hae, 8'hb5, 8'h4e, 8'h80, 8'h7b, 8'hdf, 8'h24, 8'hea, 8'h11, 8'h61, 8'h9a, 8'h54, 8'haf, 8'h0b, 8'hf0, 8'h3e, 8'hc5, 8'h08, 8'hf3, 8'h3d, 8'hc6, 8'h62, 8'h99, 8'h57, 8'hac, 8'hdc, 8'h27, 8'he9, 8'h12, 8'hb6, 8'h4d, 8'h83, 8'h78, 8'h63, 8'h98, 8'h56, 8'had, 8'h09, 8'hf2, 8'h3c, 8'hc7, 8'hb7, 8'h4c, 8'h82, 8'h79, 8'hdd, 8'h26, 8'he8, 8'h13, 8'hb1, 8'h4a, 8'h84, 8'h7f, 8'hdb, 8'h20, 8'hee, 8'h15, 8'h65, 8'h9e, 8'h50, 8'hab, 8'h0f, 8'hf4, 8'h3a, 8'hc1, 8'hda, 8'h21, 8'hef, 8'h14, 8'hb0, 8'h4b, 8'h85, 8'h7e, 8'h0e, 8'hf5, 8'h3b, 8'hc0, 8'h64, 8'h9f, 8'h51, 8'haa, 8'h67, 8'h9c, 8'h52, 8'ha9, 8'h0d, 8'hf6, 8'h38, 8'hc3, 8'hb3, 8'h48, 8'h86, 8'h7d, 8'hd9, 8'h22, 8'hec, 8'h17, 8'h0c, 8'hf7, 8'h39, 8'hc2, 8'h66, 8'h9d, 8'h53, 8'ha8, 8'hd8, 8'h23, 8'hed, 8'h16, 8'hb2, 8'h49, 8'h87, 8'h7c};
  wire [7:0] literal_2058836[256] = '{8'ha5, 8'h2d, 8'h32, 8'h8f, 8'h0e, 8'h30, 8'h38, 8'hc0, 8'h54, 8'he6, 8'h9e, 8'h39, 8'h55, 8'h7e, 8'h52, 8'h91, 8'h64, 8'h03, 8'h57, 8'h5a, 8'h1c, 8'h60, 8'h07, 8'h18, 8'h21, 8'h72, 8'ha8, 8'hd1, 8'h29, 8'hc6, 8'ha4, 8'h3f, 8'he0, 8'h27, 8'h8d, 8'h0c, 8'h82, 8'hea, 8'hae, 8'hb4, 8'h9a, 8'h63, 8'h49, 8'he5, 8'h42, 8'he4, 8'h15, 8'hb7, 8'hc8, 8'h06, 8'h70, 8'h9d, 8'h41, 8'h75, 8'h19, 8'hc9, 8'haa, 8'hfc, 8'h4d, 8'hbf, 8'h2a, 8'h73, 8'h84, 8'hd5, 8'hc3, 8'haf, 8'h2b, 8'h86, 8'ha7, 8'hb1, 8'hb2, 8'h5b, 8'h46, 8'hd3, 8'h9f, 8'hfd, 8'hd4, 8'h0f, 8'h9c, 8'h2f, 8'h9b, 8'h43, 8'hef, 8'hd9, 8'h79, 8'hb6, 8'h53, 8'h7f, 8'hc1, 8'hf0, 8'h23, 8'he7, 8'h25, 8'h5e, 8'hb5, 8'h1e, 8'ha2, 8'hdf, 8'ha6, 8'hfe, 8'hac, 8'h22, 8'hf9, 8'he2, 8'h4a, 8'hbc, 8'h35, 8'hca, 8'hee, 8'h78, 8'h05, 8'h6b, 8'h51, 8'he1, 8'h59, 8'ha3, 8'hf2, 8'h71, 8'h56, 8'h11, 8'h6a, 8'h89, 8'h94, 8'h65, 8'h8c, 8'hbb, 8'h77, 8'h3c, 8'h7b, 8'h28, 8'hab, 8'hd2, 8'h31, 8'hde, 8'hc4, 8'h5f, 8'hcc, 8'hcf, 8'h76, 8'h2c, 8'hb8, 8'hd8, 8'h2e, 8'h36, 8'hdb, 8'h69, 8'hb3, 8'h14, 8'h95, 8'hbe, 8'h62, 8'ha1, 8'h3b, 8'h16, 8'h66, 8'he9, 8'h5c, 8'h6c, 8'h6d, 8'had, 8'h37, 8'h61, 8'h4b, 8'hb9, 8'he3, 8'hba, 8'hf1, 8'ha0, 8'h85, 8'h83, 8'hda, 8'h47, 8'hc5, 8'hb0, 8'h33, 8'hfa, 8'h96, 8'h6f, 8'h6e, 8'hc2, 8'hf6, 8'h50, 8'hff, 8'h5d, 8'ha9, 8'h8e, 8'h17, 8'h1b, 8'h97, 8'h7d, 8'hec, 8'h58, 8'hf7, 8'h1f, 8'hfb, 8'h7c, 8'h09, 8'h0d, 8'h7a, 8'h67, 8'h45, 8'h87, 8'hdc, 8'he8, 8'h4f, 8'h1d, 8'h4e, 8'h04, 8'heb, 8'hf8, 8'hf3, 8'h3e, 8'h3d, 8'hbd, 8'h8a, 8'h88, 8'hdd, 8'hcd, 8'h0b, 8'h13, 8'h98, 8'h02, 8'h93, 8'h80, 8'h90, 8'hd0, 8'h24, 8'h34, 8'hcb, 8'hed, 8'hf4, 8'hce, 8'h99, 8'h10, 8'h44, 8'h40, 8'h92, 8'h3a, 8'h01, 8'h26, 8'h12, 8'h1a, 8'h48, 8'h68, 8'hf5, 8'h81, 8'h8b, 8'hc7, 8'hd6, 8'h20, 8'h0a, 8'h08, 8'h00, 8'h4c, 8'hd7, 8'h74};

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [127:0] p0_encoded;
  reg [255:0] p0_key;
  reg [7:0] p1_literal_2043896[256];
  reg [7:0] p1_literal_2043910[256];
  reg [7:0] p1_literal_2043912[256];
  reg [7:0] p1_literal_2043914[256];
  reg [7:0] p1_literal_2043916[256];
  reg [7:0] p1_literal_2043918[256];
  reg [7:0] p1_literal_2043920[256];
  reg [7:0] p1_literal_2043923[256];
  reg [7:0] p78_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p0_encoded <= encoded;
    p0_key <= key;
    p1_literal_2043896 <= literal_2043896;
    p1_literal_2043910 <= literal_2043910;
    p1_literal_2043912 <= literal_2043912;
    p1_literal_2043914 <= literal_2043914;
    p1_literal_2043916 <= literal_2043916;
    p1_literal_2043918 <= literal_2043918;
    p1_literal_2043920 <= literal_2043920;
    p1_literal_2043923 <= literal_2043923;
    p78_literal_2058836 <= literal_2058836;
  end

  // ===== Pipe stage 1:
  wire [127:0] p1_bit_slice_2043893_comb;
  wire [127:0] p1_addedKey__32_comb;
  wire [7:0] p1_array_index_2043911_comb;
  wire [7:0] p1_array_index_2043913_comb;
  wire [7:0] p1_array_index_2043915_comb;
  wire [7:0] p1_array_index_2043917_comb;
  wire [7:0] p1_array_index_2043919_comb;
  wire [7:0] p1_array_index_2043921_comb;
  wire [7:0] p1_array_index_2043924_comb;
  wire [7:0] p1_array_index_2043926_comb;
  wire [7:0] p1_array_index_2043927_comb;
  wire [7:0] p1_array_index_2043928_comb;
  wire [7:0] p1_array_index_2043929_comb;
  wire [7:0] p1_array_index_2043930_comb;
  wire [7:0] p1_array_index_2043931_comb;
  wire [7:0] p1_array_index_2043933_comb;
  wire [7:0] p1_array_index_2043934_comb;
  wire [7:0] p1_array_index_2043935_comb;
  wire [7:0] p1_array_index_2043936_comb;
  wire [7:0] p1_array_index_2043937_comb;
  wire [7:0] p1_array_index_2043938_comb;
  wire [7:0] p1_array_index_2043939_comb;
  wire [7:0] p1_array_index_2043941_comb;
  wire [7:0] p1_res7_comb;
  wire [7:0] p1_array_index_2043950_comb;
  wire [7:0] p1_array_index_2043951_comb;
  wire [7:0] p1_array_index_2043952_comb;
  wire [7:0] p1_array_index_2043953_comb;
  wire [7:0] p1_array_index_2043954_comb;
  wire [7:0] p1_array_index_2043955_comb;
  wire [7:0] p1_res7__2_comb;
  wire [7:0] p1_array_index_2043965_comb;
  wire [7:0] p1_array_index_2043966_comb;
  wire [7:0] p1_array_index_2043967_comb;
  wire [7:0] p1_array_index_2043968_comb;
  wire [7:0] p1_array_index_2043969_comb;
  wire [7:0] p1_res7__4_comb;
  wire [7:0] p1_array_index_2043979_comb;
  wire [7:0] p1_array_index_2043980_comb;
  wire [7:0] p1_array_index_2043981_comb;
  wire [7:0] p1_array_index_2043982_comb;
  wire [7:0] p1_array_index_2043983_comb;
  wire [7:0] p1_res7__6_comb;
  wire [7:0] p1_array_index_2043994_comb;
  wire [7:0] p1_array_index_2043995_comb;
  wire [7:0] p1_array_index_2043996_comb;
  wire [7:0] p1_array_index_2043997_comb;
  wire [7:0] p1_res7__8_comb;
  wire [7:0] p1_array_index_2044007_comb;
  wire [7:0] p1_array_index_2044008_comb;
  wire [7:0] p1_array_index_2044009_comb;
  wire [7:0] p1_array_index_2044010_comb;
  wire [7:0] p1_res7__10_comb;
  wire [127:0] p1_bit_slice_2044018_comb;
  assign p1_bit_slice_2043893_comb = p0_key[255:128];
  assign p1_addedKey__32_comb = p1_bit_slice_2043893_comb ^ 128'h6ea2_7672_6c48_7ab8_5d27_bd10_dd84_9401;
  assign p1_array_index_2043911_comb = literal_2043896[p1_addedKey__32_comb[127:120]];
  assign p1_array_index_2043913_comb = literal_2043896[p1_addedKey__32_comb[119:112]];
  assign p1_array_index_2043915_comb = literal_2043896[p1_addedKey__32_comb[111:104]];
  assign p1_array_index_2043917_comb = literal_2043896[p1_addedKey__32_comb[103:96]];
  assign p1_array_index_2043919_comb = literal_2043896[p1_addedKey__32_comb[95:88]];
  assign p1_array_index_2043921_comb = literal_2043896[p1_addedKey__32_comb[87:80]];
  assign p1_array_index_2043924_comb = literal_2043896[p1_addedKey__32_comb[71:64]];
  assign p1_array_index_2043926_comb = literal_2043896[p1_addedKey__32_comb[55:48]];
  assign p1_array_index_2043927_comb = literal_2043896[p1_addedKey__32_comb[47:40]];
  assign p1_array_index_2043928_comb = literal_2043896[p1_addedKey__32_comb[39:32]];
  assign p1_array_index_2043929_comb = literal_2043896[p1_addedKey__32_comb[31:24]];
  assign p1_array_index_2043930_comb = literal_2043896[p1_addedKey__32_comb[23:16]];
  assign p1_array_index_2043931_comb = literal_2043896[p1_addedKey__32_comb[15:8]];
  assign p1_array_index_2043933_comb = literal_2043910[p1_array_index_2043911_comb];
  assign p1_array_index_2043934_comb = literal_2043912[p1_array_index_2043913_comb];
  assign p1_array_index_2043935_comb = literal_2043914[p1_array_index_2043915_comb];
  assign p1_array_index_2043936_comb = literal_2043916[p1_array_index_2043917_comb];
  assign p1_array_index_2043937_comb = literal_2043918[p1_array_index_2043919_comb];
  assign p1_array_index_2043938_comb = literal_2043920[p1_array_index_2043921_comb];
  assign p1_array_index_2043939_comb = literal_2043896[p1_addedKey__32_comb[79:72]];
  assign p1_array_index_2043941_comb = literal_2043896[p1_addedKey__32_comb[63:56]];
  assign p1_res7_comb = p1_array_index_2043933_comb ^ p1_array_index_2043934_comb ^ p1_array_index_2043935_comb ^ p1_array_index_2043936_comb ^ p1_array_index_2043937_comb ^ p1_array_index_2043938_comb ^ p1_array_index_2043939_comb ^ literal_2043923[p1_array_index_2043924_comb] ^ p1_array_index_2043941_comb ^ literal_2043920[p1_array_index_2043926_comb] ^ literal_2043918[p1_array_index_2043927_comb] ^ literal_2043916[p1_array_index_2043928_comb] ^ literal_2043914[p1_array_index_2043929_comb] ^ literal_2043912[p1_array_index_2043930_comb] ^ literal_2043910[p1_array_index_2043931_comb] ^ literal_2043896[p1_addedKey__32_comb[7:0]];
  assign p1_array_index_2043950_comb = literal_2043910[p1_res7_comb];
  assign p1_array_index_2043951_comb = literal_2043912[p1_array_index_2043911_comb];
  assign p1_array_index_2043952_comb = literal_2043914[p1_array_index_2043913_comb];
  assign p1_array_index_2043953_comb = literal_2043916[p1_array_index_2043915_comb];
  assign p1_array_index_2043954_comb = literal_2043918[p1_array_index_2043917_comb];
  assign p1_array_index_2043955_comb = literal_2043920[p1_array_index_2043919_comb];
  assign p1_res7__2_comb = p1_array_index_2043950_comb ^ p1_array_index_2043951_comb ^ p1_array_index_2043952_comb ^ p1_array_index_2043953_comb ^ p1_array_index_2043954_comb ^ p1_array_index_2043955_comb ^ p1_array_index_2043921_comb ^ literal_2043923[p1_array_index_2043939_comb] ^ p1_array_index_2043924_comb ^ literal_2043920[p1_array_index_2043941_comb] ^ literal_2043918[p1_array_index_2043926_comb] ^ literal_2043916[p1_array_index_2043927_comb] ^ literal_2043914[p1_array_index_2043928_comb] ^ literal_2043912[p1_array_index_2043929_comb] ^ literal_2043910[p1_array_index_2043930_comb] ^ p1_array_index_2043931_comb;
  assign p1_array_index_2043965_comb = literal_2043912[p1_res7_comb];
  assign p1_array_index_2043966_comb = literal_2043914[p1_array_index_2043911_comb];
  assign p1_array_index_2043967_comb = literal_2043916[p1_array_index_2043913_comb];
  assign p1_array_index_2043968_comb = literal_2043918[p1_array_index_2043915_comb];
  assign p1_array_index_2043969_comb = literal_2043920[p1_array_index_2043917_comb];
  assign p1_res7__4_comb = literal_2043910[p1_res7__2_comb] ^ p1_array_index_2043965_comb ^ p1_array_index_2043966_comb ^ p1_array_index_2043967_comb ^ p1_array_index_2043968_comb ^ p1_array_index_2043969_comb ^ p1_array_index_2043919_comb ^ literal_2043923[p1_array_index_2043921_comb] ^ p1_array_index_2043939_comb ^ literal_2043920[p1_array_index_2043924_comb] ^ literal_2043918[p1_array_index_2043941_comb] ^ literal_2043916[p1_array_index_2043926_comb] ^ literal_2043914[p1_array_index_2043927_comb] ^ literal_2043912[p1_array_index_2043928_comb] ^ literal_2043910[p1_array_index_2043929_comb] ^ p1_array_index_2043930_comb;
  assign p1_array_index_2043979_comb = literal_2043912[p1_res7__2_comb];
  assign p1_array_index_2043980_comb = literal_2043914[p1_res7_comb];
  assign p1_array_index_2043981_comb = literal_2043916[p1_array_index_2043911_comb];
  assign p1_array_index_2043982_comb = literal_2043918[p1_array_index_2043913_comb];
  assign p1_array_index_2043983_comb = literal_2043920[p1_array_index_2043915_comb];
  assign p1_res7__6_comb = literal_2043910[p1_res7__4_comb] ^ p1_array_index_2043979_comb ^ p1_array_index_2043980_comb ^ p1_array_index_2043981_comb ^ p1_array_index_2043982_comb ^ p1_array_index_2043983_comb ^ p1_array_index_2043917_comb ^ literal_2043923[p1_array_index_2043919_comb] ^ p1_array_index_2043921_comb ^ literal_2043920[p1_array_index_2043939_comb] ^ literal_2043918[p1_array_index_2043924_comb] ^ literal_2043916[p1_array_index_2043941_comb] ^ literal_2043914[p1_array_index_2043926_comb] ^ literal_2043912[p1_array_index_2043927_comb] ^ literal_2043910[p1_array_index_2043928_comb] ^ p1_array_index_2043929_comb;
  assign p1_array_index_2043994_comb = literal_2043914[p1_res7__2_comb];
  assign p1_array_index_2043995_comb = literal_2043916[p1_res7_comb];
  assign p1_array_index_2043996_comb = literal_2043918[p1_array_index_2043911_comb];
  assign p1_array_index_2043997_comb = literal_2043920[p1_array_index_2043913_comb];
  assign p1_res7__8_comb = literal_2043910[p1_res7__6_comb] ^ literal_2043912[p1_res7__4_comb] ^ p1_array_index_2043994_comb ^ p1_array_index_2043995_comb ^ p1_array_index_2043996_comb ^ p1_array_index_2043997_comb ^ p1_array_index_2043915_comb ^ literal_2043923[p1_array_index_2043917_comb] ^ p1_array_index_2043919_comb ^ p1_array_index_2043938_comb ^ literal_2043918[p1_array_index_2043939_comb] ^ literal_2043916[p1_array_index_2043924_comb] ^ literal_2043914[p1_array_index_2043941_comb] ^ literal_2043912[p1_array_index_2043926_comb] ^ literal_2043910[p1_array_index_2043927_comb] ^ p1_array_index_2043928_comb;
  assign p1_array_index_2044007_comb = literal_2043914[p1_res7__4_comb];
  assign p1_array_index_2044008_comb = literal_2043916[p1_res7__2_comb];
  assign p1_array_index_2044009_comb = literal_2043918[p1_res7_comb];
  assign p1_array_index_2044010_comb = literal_2043920[p1_array_index_2043911_comb];
  assign p1_res7__10_comb = literal_2043910[p1_res7__8_comb] ^ literal_2043912[p1_res7__6_comb] ^ p1_array_index_2044007_comb ^ p1_array_index_2044008_comb ^ p1_array_index_2044009_comb ^ p1_array_index_2044010_comb ^ p1_array_index_2043913_comb ^ literal_2043923[p1_array_index_2043915_comb] ^ p1_array_index_2043917_comb ^ p1_array_index_2043955_comb ^ literal_2043918[p1_array_index_2043921_comb] ^ literal_2043916[p1_array_index_2043939_comb] ^ literal_2043914[p1_array_index_2043924_comb] ^ literal_2043912[p1_array_index_2043941_comb] ^ literal_2043910[p1_array_index_2043926_comb] ^ p1_array_index_2043927_comb;
  assign p1_bit_slice_2044018_comb = p0_key[127:0];

  // Registers for pipe stage 1:
  reg [127:0] p1_encoded;
  reg [127:0] p1_bit_slice_2043893;
  reg [7:0] p1_array_index_2043911;
  reg [7:0] p1_array_index_2043913;
  reg [7:0] p1_array_index_2043915;
  reg [7:0] p1_array_index_2043917;
  reg [7:0] p1_array_index_2043919;
  reg [7:0] p1_array_index_2043921;
  reg [7:0] p1_array_index_2043924;
  reg [7:0] p1_array_index_2043926;
  reg [7:0] p1_array_index_2043933;
  reg [7:0] p1_array_index_2043934;
  reg [7:0] p1_array_index_2043935;
  reg [7:0] p1_array_index_2043936;
  reg [7:0] p1_array_index_2043937;
  reg [7:0] p1_array_index_2043939;
  reg [7:0] p1_array_index_2043941;
  reg [7:0] p1_res7;
  reg [7:0] p1_array_index_2043950;
  reg [7:0] p1_array_index_2043951;
  reg [7:0] p1_array_index_2043952;
  reg [7:0] p1_array_index_2043953;
  reg [7:0] p1_array_index_2043954;
  reg [7:0] p1_res7__2;
  reg [7:0] p1_array_index_2043965;
  reg [7:0] p1_array_index_2043966;
  reg [7:0] p1_array_index_2043967;
  reg [7:0] p1_array_index_2043968;
  reg [7:0] p1_array_index_2043969;
  reg [7:0] p1_res7__4;
  reg [7:0] p1_array_index_2043979;
  reg [7:0] p1_array_index_2043980;
  reg [7:0] p1_array_index_2043981;
  reg [7:0] p1_array_index_2043982;
  reg [7:0] p1_array_index_2043983;
  reg [7:0] p1_res7__6;
  reg [7:0] p1_array_index_2043994;
  reg [7:0] p1_array_index_2043995;
  reg [7:0] p1_array_index_2043996;
  reg [7:0] p1_array_index_2043997;
  reg [7:0] p1_res7__8;
  reg [7:0] p1_array_index_2044007;
  reg [7:0] p1_array_index_2044008;
  reg [7:0] p1_array_index_2044009;
  reg [7:0] p1_array_index_2044010;
  reg [7:0] p1_res7__10;
  reg [127:0] p1_bit_slice_2044018;
  reg [7:0] p2_literal_2043896[256];
  reg [7:0] p2_literal_2043910[256];
  reg [7:0] p2_literal_2043912[256];
  reg [7:0] p2_literal_2043914[256];
  reg [7:0] p2_literal_2043916[256];
  reg [7:0] p2_literal_2043918[256];
  reg [7:0] p2_literal_2043920[256];
  reg [7:0] p2_literal_2043923[256];
  reg [7:0] p79_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p1_encoded <= p0_encoded;
    p1_bit_slice_2043893 <= p1_bit_slice_2043893_comb;
    p1_array_index_2043911 <= p1_array_index_2043911_comb;
    p1_array_index_2043913 <= p1_array_index_2043913_comb;
    p1_array_index_2043915 <= p1_array_index_2043915_comb;
    p1_array_index_2043917 <= p1_array_index_2043917_comb;
    p1_array_index_2043919 <= p1_array_index_2043919_comb;
    p1_array_index_2043921 <= p1_array_index_2043921_comb;
    p1_array_index_2043924 <= p1_array_index_2043924_comb;
    p1_array_index_2043926 <= p1_array_index_2043926_comb;
    p1_array_index_2043933 <= p1_array_index_2043933_comb;
    p1_array_index_2043934 <= p1_array_index_2043934_comb;
    p1_array_index_2043935 <= p1_array_index_2043935_comb;
    p1_array_index_2043936 <= p1_array_index_2043936_comb;
    p1_array_index_2043937 <= p1_array_index_2043937_comb;
    p1_array_index_2043939 <= p1_array_index_2043939_comb;
    p1_array_index_2043941 <= p1_array_index_2043941_comb;
    p1_res7 <= p1_res7_comb;
    p1_array_index_2043950 <= p1_array_index_2043950_comb;
    p1_array_index_2043951 <= p1_array_index_2043951_comb;
    p1_array_index_2043952 <= p1_array_index_2043952_comb;
    p1_array_index_2043953 <= p1_array_index_2043953_comb;
    p1_array_index_2043954 <= p1_array_index_2043954_comb;
    p1_res7__2 <= p1_res7__2_comb;
    p1_array_index_2043965 <= p1_array_index_2043965_comb;
    p1_array_index_2043966 <= p1_array_index_2043966_comb;
    p1_array_index_2043967 <= p1_array_index_2043967_comb;
    p1_array_index_2043968 <= p1_array_index_2043968_comb;
    p1_array_index_2043969 <= p1_array_index_2043969_comb;
    p1_res7__4 <= p1_res7__4_comb;
    p1_array_index_2043979 <= p1_array_index_2043979_comb;
    p1_array_index_2043980 <= p1_array_index_2043980_comb;
    p1_array_index_2043981 <= p1_array_index_2043981_comb;
    p1_array_index_2043982 <= p1_array_index_2043982_comb;
    p1_array_index_2043983 <= p1_array_index_2043983_comb;
    p1_res7__6 <= p1_res7__6_comb;
    p1_array_index_2043994 <= p1_array_index_2043994_comb;
    p1_array_index_2043995 <= p1_array_index_2043995_comb;
    p1_array_index_2043996 <= p1_array_index_2043996_comb;
    p1_array_index_2043997 <= p1_array_index_2043997_comb;
    p1_res7__8 <= p1_res7__8_comb;
    p1_array_index_2044007 <= p1_array_index_2044007_comb;
    p1_array_index_2044008 <= p1_array_index_2044008_comb;
    p1_array_index_2044009 <= p1_array_index_2044009_comb;
    p1_array_index_2044010 <= p1_array_index_2044010_comb;
    p1_res7__10 <= p1_res7__10_comb;
    p1_bit_slice_2044018 <= p1_bit_slice_2044018_comb;
    p2_literal_2043896 <= p1_literal_2043896;
    p2_literal_2043910 <= p1_literal_2043910;
    p2_literal_2043912 <= p1_literal_2043912;
    p2_literal_2043914 <= p1_literal_2043914;
    p2_literal_2043916 <= p1_literal_2043916;
    p2_literal_2043918 <= p1_literal_2043918;
    p2_literal_2043920 <= p1_literal_2043920;
    p2_literal_2043923 <= p1_literal_2043923;
    p79_literal_2058836 <= p78_literal_2058836;
  end

  // ===== Pipe stage 2:
  wire [7:0] p2_array_index_2044132_comb;
  wire [7:0] p2_array_index_2044133_comb;
  wire [7:0] p2_array_index_2044134_comb;
  wire [7:0] p2_res7__12_comb;
  wire [7:0] p2_array_index_2044144_comb;
  wire [7:0] p2_array_index_2044145_comb;
  wire [7:0] p2_array_index_2044146_comb;
  wire [7:0] p2_res7__14_comb;
  wire [7:0] p2_array_index_2044157_comb;
  wire [7:0] p2_array_index_2044158_comb;
  wire [7:0] p2_res7__16_comb;
  wire [7:0] p2_array_index_2044168_comb;
  wire [7:0] p2_array_index_2044169_comb;
  wire [7:0] p2_res7__18_comb;
  wire [7:0] p2_array_index_2044180_comb;
  wire [7:0] p2_res7__20_comb;
  wire [7:0] p2_array_index_2044190_comb;
  wire [7:0] p2_res7__22_comb;
  wire [7:0] p2_res7__24_comb;
  assign p2_array_index_2044132_comb = p1_literal_2043916[p1_res7__4];
  assign p2_array_index_2044133_comb = p1_literal_2043918[p1_res7__2];
  assign p2_array_index_2044134_comb = p1_literal_2043920[p1_res7];
  assign p2_res7__12_comb = p1_literal_2043910[p1_res7__10] ^ p1_literal_2043912[p1_res7__8] ^ p1_literal_2043914[p1_res7__6] ^ p2_array_index_2044132_comb ^ p2_array_index_2044133_comb ^ p2_array_index_2044134_comb ^ p1_array_index_2043911 ^ p1_literal_2043923[p1_array_index_2043913] ^ p1_array_index_2043915 ^ p1_array_index_2043969 ^ p1_array_index_2043937 ^ p1_literal_2043916[p1_array_index_2043921] ^ p1_literal_2043914[p1_array_index_2043939] ^ p1_literal_2043912[p1_array_index_2043924] ^ p1_literal_2043910[p1_array_index_2043941] ^ p1_array_index_2043926;
  assign p2_array_index_2044144_comb = p1_literal_2043916[p1_res7__6];
  assign p2_array_index_2044145_comb = p1_literal_2043918[p1_res7__4];
  assign p2_array_index_2044146_comb = p1_literal_2043920[p1_res7__2];
  assign p2_res7__14_comb = p1_literal_2043910[p2_res7__12_comb] ^ p1_literal_2043912[p1_res7__10] ^ p1_literal_2043914[p1_res7__8] ^ p2_array_index_2044144_comb ^ p2_array_index_2044145_comb ^ p2_array_index_2044146_comb ^ p1_res7 ^ p1_literal_2043923[p1_array_index_2043911] ^ p1_array_index_2043913 ^ p1_array_index_2043983 ^ p1_array_index_2043954 ^ p1_literal_2043916[p1_array_index_2043919] ^ p1_literal_2043914[p1_array_index_2043921] ^ p1_literal_2043912[p1_array_index_2043939] ^ p1_literal_2043910[p1_array_index_2043924] ^ p1_array_index_2043941;
  assign p2_array_index_2044157_comb = p1_literal_2043918[p1_res7__6];
  assign p2_array_index_2044158_comb = p1_literal_2043920[p1_res7__4];
  assign p2_res7__16_comb = p1_literal_2043910[p2_res7__14_comb] ^ p1_literal_2043912[p2_res7__12_comb] ^ p1_literal_2043914[p1_res7__10] ^ p1_literal_2043916[p1_res7__8] ^ p2_array_index_2044157_comb ^ p2_array_index_2044158_comb ^ p1_res7__2 ^ p1_literal_2043923[p1_res7] ^ p1_array_index_2043911 ^ p1_array_index_2043997 ^ p1_array_index_2043968 ^ p1_array_index_2043936 ^ p1_literal_2043914[p1_array_index_2043919] ^ p1_literal_2043912[p1_array_index_2043921] ^ p1_literal_2043910[p1_array_index_2043939] ^ p1_array_index_2043924;
  assign p2_array_index_2044168_comb = p1_literal_2043918[p1_res7__8];
  assign p2_array_index_2044169_comb = p1_literal_2043920[p1_res7__6];
  assign p2_res7__18_comb = p1_literal_2043910[p2_res7__16_comb] ^ p1_literal_2043912[p2_res7__14_comb] ^ p1_literal_2043914[p2_res7__12_comb] ^ p1_literal_2043916[p1_res7__10] ^ p2_array_index_2044168_comb ^ p2_array_index_2044169_comb ^ p1_res7__4 ^ p1_literal_2043923[p1_res7__2] ^ p1_res7 ^ p1_array_index_2044010 ^ p1_array_index_2043982 ^ p1_array_index_2043953 ^ p1_literal_2043914[p1_array_index_2043917] ^ p1_literal_2043912[p1_array_index_2043919] ^ p1_literal_2043910[p1_array_index_2043921] ^ p1_array_index_2043939;
  assign p2_array_index_2044180_comb = p1_literal_2043920[p1_res7__8];
  assign p2_res7__20_comb = p1_literal_2043910[p2_res7__18_comb] ^ p1_literal_2043912[p2_res7__16_comb] ^ p1_literal_2043914[p2_res7__14_comb] ^ p1_literal_2043916[p2_res7__12_comb] ^ p1_literal_2043918[p1_res7__10] ^ p2_array_index_2044180_comb ^ p1_res7__6 ^ p1_literal_2043923[p1_res7__4] ^ p1_res7__2 ^ p2_array_index_2044134_comb ^ p1_array_index_2043996 ^ p1_array_index_2043967 ^ p1_array_index_2043935 ^ p1_literal_2043912[p1_array_index_2043917] ^ p1_literal_2043910[p1_array_index_2043919] ^ p1_array_index_2043921;
  assign p2_array_index_2044190_comb = p1_literal_2043920[p1_res7__10];
  assign p2_res7__22_comb = p1_literal_2043910[p2_res7__20_comb] ^ p1_literal_2043912[p2_res7__18_comb] ^ p1_literal_2043914[p2_res7__16_comb] ^ p1_literal_2043916[p2_res7__14_comb] ^ p1_literal_2043918[p2_res7__12_comb] ^ p2_array_index_2044190_comb ^ p1_res7__8 ^ p1_literal_2043923[p1_res7__6] ^ p1_res7__4 ^ p2_array_index_2044146_comb ^ p1_array_index_2044009 ^ p1_array_index_2043981 ^ p1_array_index_2043952 ^ p1_literal_2043912[p1_array_index_2043915] ^ p1_literal_2043910[p1_array_index_2043917] ^ p1_array_index_2043919;
  assign p2_res7__24_comb = p1_literal_2043910[p2_res7__22_comb] ^ p1_literal_2043912[p2_res7__20_comb] ^ p1_literal_2043914[p2_res7__18_comb] ^ p1_literal_2043916[p2_res7__16_comb] ^ p1_literal_2043918[p2_res7__14_comb] ^ p1_literal_2043920[p2_res7__12_comb] ^ p1_res7__10 ^ p1_literal_2043923[p1_res7__8] ^ p1_res7__6 ^ p2_array_index_2044158_comb ^ p2_array_index_2044133_comb ^ p1_array_index_2043995 ^ p1_array_index_2043966 ^ p1_array_index_2043934 ^ p1_literal_2043910[p1_array_index_2043915] ^ p1_array_index_2043917;

  // Registers for pipe stage 2:
  reg [127:0] p2_encoded;
  reg [127:0] p2_bit_slice_2043893;
  reg [7:0] p2_array_index_2043911;
  reg [7:0] p2_array_index_2043913;
  reg [7:0] p2_array_index_2043915;
  reg [7:0] p2_array_index_2043933;
  reg [7:0] p2_res7;
  reg [7:0] p2_array_index_2043950;
  reg [7:0] p2_array_index_2043951;
  reg [7:0] p2_res7__2;
  reg [7:0] p2_array_index_2043965;
  reg [7:0] p2_res7__4;
  reg [7:0] p2_array_index_2043979;
  reg [7:0] p2_array_index_2043980;
  reg [7:0] p2_res7__6;
  reg [7:0] p2_array_index_2043994;
  reg [7:0] p2_res7__8;
  reg [7:0] p2_array_index_2044007;
  reg [7:0] p2_array_index_2044008;
  reg [7:0] p2_res7__10;
  reg [7:0] p2_array_index_2044132;
  reg [7:0] p2_res7__12;
  reg [7:0] p2_array_index_2044144;
  reg [7:0] p2_array_index_2044145;
  reg [7:0] p2_res7__14;
  reg [7:0] p2_array_index_2044157;
  reg [7:0] p2_res7__16;
  reg [7:0] p2_array_index_2044168;
  reg [7:0] p2_array_index_2044169;
  reg [7:0] p2_res7__18;
  reg [7:0] p2_array_index_2044180;
  reg [7:0] p2_res7__20;
  reg [7:0] p2_array_index_2044190;
  reg [7:0] p2_res7__22;
  reg [7:0] p2_res7__24;
  reg [127:0] p2_bit_slice_2044018;
  reg [7:0] p3_literal_2043896[256];
  reg [7:0] p3_literal_2043910[256];
  reg [7:0] p3_literal_2043912[256];
  reg [7:0] p3_literal_2043914[256];
  reg [7:0] p3_literal_2043916[256];
  reg [7:0] p3_literal_2043918[256];
  reg [7:0] p3_literal_2043920[256];
  reg [7:0] p3_literal_2043923[256];
  reg [7:0] p80_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p2_encoded <= p1_encoded;
    p2_bit_slice_2043893 <= p1_bit_slice_2043893;
    p2_array_index_2043911 <= p1_array_index_2043911;
    p2_array_index_2043913 <= p1_array_index_2043913;
    p2_array_index_2043915 <= p1_array_index_2043915;
    p2_array_index_2043933 <= p1_array_index_2043933;
    p2_res7 <= p1_res7;
    p2_array_index_2043950 <= p1_array_index_2043950;
    p2_array_index_2043951 <= p1_array_index_2043951;
    p2_res7__2 <= p1_res7__2;
    p2_array_index_2043965 <= p1_array_index_2043965;
    p2_res7__4 <= p1_res7__4;
    p2_array_index_2043979 <= p1_array_index_2043979;
    p2_array_index_2043980 <= p1_array_index_2043980;
    p2_res7__6 <= p1_res7__6;
    p2_array_index_2043994 <= p1_array_index_2043994;
    p2_res7__8 <= p1_res7__8;
    p2_array_index_2044007 <= p1_array_index_2044007;
    p2_array_index_2044008 <= p1_array_index_2044008;
    p2_res7__10 <= p1_res7__10;
    p2_array_index_2044132 <= p2_array_index_2044132_comb;
    p2_res7__12 <= p2_res7__12_comb;
    p2_array_index_2044144 <= p2_array_index_2044144_comb;
    p2_array_index_2044145 <= p2_array_index_2044145_comb;
    p2_res7__14 <= p2_res7__14_comb;
    p2_array_index_2044157 <= p2_array_index_2044157_comb;
    p2_res7__16 <= p2_res7__16_comb;
    p2_array_index_2044168 <= p2_array_index_2044168_comb;
    p2_array_index_2044169 <= p2_array_index_2044169_comb;
    p2_res7__18 <= p2_res7__18_comb;
    p2_array_index_2044180 <= p2_array_index_2044180_comb;
    p2_res7__20 <= p2_res7__20_comb;
    p2_array_index_2044190 <= p2_array_index_2044190_comb;
    p2_res7__22 <= p2_res7__22_comb;
    p2_res7__24 <= p2_res7__24_comb;
    p2_bit_slice_2044018 <= p1_bit_slice_2044018;
    p3_literal_2043896 <= p2_literal_2043896;
    p3_literal_2043910 <= p2_literal_2043910;
    p3_literal_2043912 <= p2_literal_2043912;
    p3_literal_2043914 <= p2_literal_2043914;
    p3_literal_2043916 <= p2_literal_2043916;
    p3_literal_2043918 <= p2_literal_2043918;
    p3_literal_2043920 <= p2_literal_2043920;
    p3_literal_2043923 <= p2_literal_2043923;
    p80_literal_2058836 <= p79_literal_2058836;
  end

  // ===== Pipe stage 3:
  wire [7:0] p3_res7__26_comb;
  wire [7:0] p3_res7__28_comb;
  wire [7:0] p3_res7__30_comb;
  wire [127:0] p3_res_comb;
  wire [127:0] p3_xor_2044318_comb;
  wire [127:0] p3_addedKey__33_comb;
  wire [7:0] p3_array_index_2044334_comb;
  wire [7:0] p3_array_index_2044335_comb;
  wire [7:0] p3_array_index_2044336_comb;
  wire [7:0] p3_array_index_2044337_comb;
  wire [7:0] p3_array_index_2044338_comb;
  wire [7:0] p3_array_index_2044339_comb;
  wire [7:0] p3_array_index_2044341_comb;
  wire [7:0] p3_array_index_2044343_comb;
  wire [7:0] p3_array_index_2044344_comb;
  wire [7:0] p3_array_index_2044345_comb;
  wire [7:0] p3_array_index_2044346_comb;
  wire [7:0] p3_array_index_2044347_comb;
  wire [7:0] p3_array_index_2044348_comb;
  wire [7:0] p3_array_index_2044350_comb;
  wire [7:0] p3_array_index_2044351_comb;
  wire [7:0] p3_array_index_2044352_comb;
  wire [7:0] p3_array_index_2044353_comb;
  wire [7:0] p3_array_index_2044354_comb;
  wire [7:0] p3_array_index_2044355_comb;
  wire [7:0] p3_array_index_2044356_comb;
  wire [7:0] p3_array_index_2044358_comb;
  wire [7:0] p3_res7__32_comb;
  wire [7:0] p3_array_index_2044367_comb;
  wire [7:0] p3_array_index_2044368_comb;
  wire [7:0] p3_array_index_2044369_comb;
  wire [7:0] p3_array_index_2044370_comb;
  wire [7:0] p3_array_index_2044371_comb;
  wire [7:0] p3_array_index_2044372_comb;
  wire [7:0] p3_res7__34_comb;
  wire [7:0] p3_array_index_2044382_comb;
  wire [7:0] p3_array_index_2044383_comb;
  wire [7:0] p3_array_index_2044384_comb;
  wire [7:0] p3_array_index_2044385_comb;
  wire [7:0] p3_array_index_2044386_comb;
  wire [7:0] p3_res7__36_comb;
  assign p3_res7__26_comb = p2_literal_2043910[p2_res7__24] ^ p2_literal_2043912[p2_res7__22] ^ p2_literal_2043914[p2_res7__20] ^ p2_literal_2043916[p2_res7__18] ^ p2_literal_2043918[p2_res7__16] ^ p2_literal_2043920[p2_res7__14] ^ p2_res7__12 ^ p2_literal_2043923[p2_res7__10] ^ p2_res7__8 ^ p2_array_index_2044169 ^ p2_array_index_2044145 ^ p2_array_index_2044008 ^ p2_array_index_2043980 ^ p2_array_index_2043951 ^ p2_literal_2043910[p2_array_index_2043913] ^ p2_array_index_2043915;
  assign p3_res7__28_comb = p2_literal_2043910[p3_res7__26_comb] ^ p2_literal_2043912[p2_res7__24] ^ p2_literal_2043914[p2_res7__22] ^ p2_literal_2043916[p2_res7__20] ^ p2_literal_2043918[p2_res7__18] ^ p2_literal_2043920[p2_res7__16] ^ p2_res7__14 ^ p2_literal_2043923[p2_res7__12] ^ p2_res7__10 ^ p2_array_index_2044180 ^ p2_array_index_2044157 ^ p2_array_index_2044132 ^ p2_array_index_2043994 ^ p2_array_index_2043965 ^ p2_array_index_2043933 ^ p2_array_index_2043913;
  assign p3_res7__30_comb = p2_literal_2043910[p3_res7__28_comb] ^ p2_literal_2043912[p3_res7__26_comb] ^ p2_literal_2043914[p2_res7__24] ^ p2_literal_2043916[p2_res7__22] ^ p2_literal_2043918[p2_res7__20] ^ p2_literal_2043920[p2_res7__18] ^ p2_res7__16 ^ p2_literal_2043923[p2_res7__14] ^ p2_res7__12 ^ p2_array_index_2044190 ^ p2_array_index_2044168 ^ p2_array_index_2044144 ^ p2_array_index_2044007 ^ p2_array_index_2043979 ^ p2_array_index_2043950 ^ p2_array_index_2043911;
  assign p3_res_comb = {p3_res7__30_comb, p3_res7__28_comb, p3_res7__26_comb, p2_res7__24, p2_res7__22, p2_res7__20, p2_res7__18, p2_res7__16, p2_res7__14, p2_res7__12, p2_res7__10, p2_res7__8, p2_res7__6, p2_res7__4, p2_res7__2, p2_res7};
  assign p3_xor_2044318_comb = p3_res_comb ^ p2_bit_slice_2044018;
  assign p3_addedKey__33_comb = p3_xor_2044318_comb ^ 128'hdc87_ece4_d890_f4b3_ba4e_b920_79cb_eb02;
  assign p3_array_index_2044334_comb = p2_literal_2043896[p3_addedKey__33_comb[127:120]];
  assign p3_array_index_2044335_comb = p2_literal_2043896[p3_addedKey__33_comb[119:112]];
  assign p3_array_index_2044336_comb = p2_literal_2043896[p3_addedKey__33_comb[111:104]];
  assign p3_array_index_2044337_comb = p2_literal_2043896[p3_addedKey__33_comb[103:96]];
  assign p3_array_index_2044338_comb = p2_literal_2043896[p3_addedKey__33_comb[95:88]];
  assign p3_array_index_2044339_comb = p2_literal_2043896[p3_addedKey__33_comb[87:80]];
  assign p3_array_index_2044341_comb = p2_literal_2043896[p3_addedKey__33_comb[71:64]];
  assign p3_array_index_2044343_comb = p2_literal_2043896[p3_addedKey__33_comb[55:48]];
  assign p3_array_index_2044344_comb = p2_literal_2043896[p3_addedKey__33_comb[47:40]];
  assign p3_array_index_2044345_comb = p2_literal_2043896[p3_addedKey__33_comb[39:32]];
  assign p3_array_index_2044346_comb = p2_literal_2043896[p3_addedKey__33_comb[31:24]];
  assign p3_array_index_2044347_comb = p2_literal_2043896[p3_addedKey__33_comb[23:16]];
  assign p3_array_index_2044348_comb = p2_literal_2043896[p3_addedKey__33_comb[15:8]];
  assign p3_array_index_2044350_comb = p2_literal_2043910[p3_array_index_2044334_comb];
  assign p3_array_index_2044351_comb = p2_literal_2043912[p3_array_index_2044335_comb];
  assign p3_array_index_2044352_comb = p2_literal_2043914[p3_array_index_2044336_comb];
  assign p3_array_index_2044353_comb = p2_literal_2043916[p3_array_index_2044337_comb];
  assign p3_array_index_2044354_comb = p2_literal_2043918[p3_array_index_2044338_comb];
  assign p3_array_index_2044355_comb = p2_literal_2043920[p3_array_index_2044339_comb];
  assign p3_array_index_2044356_comb = p2_literal_2043896[p3_addedKey__33_comb[79:72]];
  assign p3_array_index_2044358_comb = p2_literal_2043896[p3_addedKey__33_comb[63:56]];
  assign p3_res7__32_comb = p3_array_index_2044350_comb ^ p3_array_index_2044351_comb ^ p3_array_index_2044352_comb ^ p3_array_index_2044353_comb ^ p3_array_index_2044354_comb ^ p3_array_index_2044355_comb ^ p3_array_index_2044356_comb ^ p2_literal_2043923[p3_array_index_2044341_comb] ^ p3_array_index_2044358_comb ^ p2_literal_2043920[p3_array_index_2044343_comb] ^ p2_literal_2043918[p3_array_index_2044344_comb] ^ p2_literal_2043916[p3_array_index_2044345_comb] ^ p2_literal_2043914[p3_array_index_2044346_comb] ^ p2_literal_2043912[p3_array_index_2044347_comb] ^ p2_literal_2043910[p3_array_index_2044348_comb] ^ p2_literal_2043896[p3_addedKey__33_comb[7:0]];
  assign p3_array_index_2044367_comb = p2_literal_2043910[p3_res7__32_comb];
  assign p3_array_index_2044368_comb = p2_literal_2043912[p3_array_index_2044334_comb];
  assign p3_array_index_2044369_comb = p2_literal_2043914[p3_array_index_2044335_comb];
  assign p3_array_index_2044370_comb = p2_literal_2043916[p3_array_index_2044336_comb];
  assign p3_array_index_2044371_comb = p2_literal_2043918[p3_array_index_2044337_comb];
  assign p3_array_index_2044372_comb = p2_literal_2043920[p3_array_index_2044338_comb];
  assign p3_res7__34_comb = p3_array_index_2044367_comb ^ p3_array_index_2044368_comb ^ p3_array_index_2044369_comb ^ p3_array_index_2044370_comb ^ p3_array_index_2044371_comb ^ p3_array_index_2044372_comb ^ p3_array_index_2044339_comb ^ p2_literal_2043923[p3_array_index_2044356_comb] ^ p3_array_index_2044341_comb ^ p2_literal_2043920[p3_array_index_2044358_comb] ^ p2_literal_2043918[p3_array_index_2044343_comb] ^ p2_literal_2043916[p3_array_index_2044344_comb] ^ p2_literal_2043914[p3_array_index_2044345_comb] ^ p2_literal_2043912[p3_array_index_2044346_comb] ^ p2_literal_2043910[p3_array_index_2044347_comb] ^ p3_array_index_2044348_comb;
  assign p3_array_index_2044382_comb = p2_literal_2043912[p3_res7__32_comb];
  assign p3_array_index_2044383_comb = p2_literal_2043914[p3_array_index_2044334_comb];
  assign p3_array_index_2044384_comb = p2_literal_2043916[p3_array_index_2044335_comb];
  assign p3_array_index_2044385_comb = p2_literal_2043918[p3_array_index_2044336_comb];
  assign p3_array_index_2044386_comb = p2_literal_2043920[p3_array_index_2044337_comb];
  assign p3_res7__36_comb = p2_literal_2043910[p3_res7__34_comb] ^ p3_array_index_2044382_comb ^ p3_array_index_2044383_comb ^ p3_array_index_2044384_comb ^ p3_array_index_2044385_comb ^ p3_array_index_2044386_comb ^ p3_array_index_2044338_comb ^ p2_literal_2043923[p3_array_index_2044339_comb] ^ p3_array_index_2044356_comb ^ p2_literal_2043920[p3_array_index_2044341_comb] ^ p2_literal_2043918[p3_array_index_2044358_comb] ^ p2_literal_2043916[p3_array_index_2044343_comb] ^ p2_literal_2043914[p3_array_index_2044344_comb] ^ p2_literal_2043912[p3_array_index_2044345_comb] ^ p2_literal_2043910[p3_array_index_2044346_comb] ^ p3_array_index_2044347_comb;

  // Registers for pipe stage 3:
  reg [127:0] p3_encoded;
  reg [127:0] p3_bit_slice_2043893;
  reg [127:0] p3_bit_slice_2044018;
  reg [127:0] p3_xor_2044318;
  reg [7:0] p3_array_index_2044334;
  reg [7:0] p3_array_index_2044335;
  reg [7:0] p3_array_index_2044336;
  reg [7:0] p3_array_index_2044337;
  reg [7:0] p3_array_index_2044338;
  reg [7:0] p3_array_index_2044339;
  reg [7:0] p3_array_index_2044341;
  reg [7:0] p3_array_index_2044343;
  reg [7:0] p3_array_index_2044344;
  reg [7:0] p3_array_index_2044345;
  reg [7:0] p3_array_index_2044346;
  reg [7:0] p3_array_index_2044350;
  reg [7:0] p3_array_index_2044351;
  reg [7:0] p3_array_index_2044352;
  reg [7:0] p3_array_index_2044353;
  reg [7:0] p3_array_index_2044354;
  reg [7:0] p3_array_index_2044355;
  reg [7:0] p3_array_index_2044356;
  reg [7:0] p3_array_index_2044358;
  reg [7:0] p3_res7__32;
  reg [7:0] p3_array_index_2044367;
  reg [7:0] p3_array_index_2044368;
  reg [7:0] p3_array_index_2044369;
  reg [7:0] p3_array_index_2044370;
  reg [7:0] p3_array_index_2044371;
  reg [7:0] p3_array_index_2044372;
  reg [7:0] p3_res7__34;
  reg [7:0] p3_array_index_2044382;
  reg [7:0] p3_array_index_2044383;
  reg [7:0] p3_array_index_2044384;
  reg [7:0] p3_array_index_2044385;
  reg [7:0] p3_array_index_2044386;
  reg [7:0] p3_res7__36;
  reg [7:0] p4_literal_2043896[256];
  reg [7:0] p4_literal_2043910[256];
  reg [7:0] p4_literal_2043912[256];
  reg [7:0] p4_literal_2043914[256];
  reg [7:0] p4_literal_2043916[256];
  reg [7:0] p4_literal_2043918[256];
  reg [7:0] p4_literal_2043920[256];
  reg [7:0] p4_literal_2043923[256];
  reg [7:0] p81_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p3_encoded <= p2_encoded;
    p3_bit_slice_2043893 <= p2_bit_slice_2043893;
    p3_bit_slice_2044018 <= p2_bit_slice_2044018;
    p3_xor_2044318 <= p3_xor_2044318_comb;
    p3_array_index_2044334 <= p3_array_index_2044334_comb;
    p3_array_index_2044335 <= p3_array_index_2044335_comb;
    p3_array_index_2044336 <= p3_array_index_2044336_comb;
    p3_array_index_2044337 <= p3_array_index_2044337_comb;
    p3_array_index_2044338 <= p3_array_index_2044338_comb;
    p3_array_index_2044339 <= p3_array_index_2044339_comb;
    p3_array_index_2044341 <= p3_array_index_2044341_comb;
    p3_array_index_2044343 <= p3_array_index_2044343_comb;
    p3_array_index_2044344 <= p3_array_index_2044344_comb;
    p3_array_index_2044345 <= p3_array_index_2044345_comb;
    p3_array_index_2044346 <= p3_array_index_2044346_comb;
    p3_array_index_2044350 <= p3_array_index_2044350_comb;
    p3_array_index_2044351 <= p3_array_index_2044351_comb;
    p3_array_index_2044352 <= p3_array_index_2044352_comb;
    p3_array_index_2044353 <= p3_array_index_2044353_comb;
    p3_array_index_2044354 <= p3_array_index_2044354_comb;
    p3_array_index_2044355 <= p3_array_index_2044355_comb;
    p3_array_index_2044356 <= p3_array_index_2044356_comb;
    p3_array_index_2044358 <= p3_array_index_2044358_comb;
    p3_res7__32 <= p3_res7__32_comb;
    p3_array_index_2044367 <= p3_array_index_2044367_comb;
    p3_array_index_2044368 <= p3_array_index_2044368_comb;
    p3_array_index_2044369 <= p3_array_index_2044369_comb;
    p3_array_index_2044370 <= p3_array_index_2044370_comb;
    p3_array_index_2044371 <= p3_array_index_2044371_comb;
    p3_array_index_2044372 <= p3_array_index_2044372_comb;
    p3_res7__34 <= p3_res7__34_comb;
    p3_array_index_2044382 <= p3_array_index_2044382_comb;
    p3_array_index_2044383 <= p3_array_index_2044383_comb;
    p3_array_index_2044384 <= p3_array_index_2044384_comb;
    p3_array_index_2044385 <= p3_array_index_2044385_comb;
    p3_array_index_2044386 <= p3_array_index_2044386_comb;
    p3_res7__36 <= p3_res7__36_comb;
    p4_literal_2043896 <= p3_literal_2043896;
    p4_literal_2043910 <= p3_literal_2043910;
    p4_literal_2043912 <= p3_literal_2043912;
    p4_literal_2043914 <= p3_literal_2043914;
    p4_literal_2043916 <= p3_literal_2043916;
    p4_literal_2043918 <= p3_literal_2043918;
    p4_literal_2043920 <= p3_literal_2043920;
    p4_literal_2043923 <= p3_literal_2043923;
    p81_literal_2058836 <= p80_literal_2058836;
  end

  // ===== Pipe stage 4:
  wire [7:0] p4_array_index_2044486_comb;
  wire [7:0] p4_array_index_2044487_comb;
  wire [7:0] p4_array_index_2044488_comb;
  wire [7:0] p4_array_index_2044489_comb;
  wire [7:0] p4_array_index_2044490_comb;
  wire [7:0] p4_res7__38_comb;
  wire [7:0] p4_array_index_2044501_comb;
  wire [7:0] p4_array_index_2044502_comb;
  wire [7:0] p4_array_index_2044503_comb;
  wire [7:0] p4_array_index_2044504_comb;
  wire [7:0] p4_res7__40_comb;
  wire [7:0] p4_array_index_2044514_comb;
  wire [7:0] p4_array_index_2044515_comb;
  wire [7:0] p4_array_index_2044516_comb;
  wire [7:0] p4_array_index_2044517_comb;
  wire [7:0] p4_res7__42_comb;
  wire [7:0] p4_array_index_2044528_comb;
  wire [7:0] p4_array_index_2044529_comb;
  wire [7:0] p4_array_index_2044530_comb;
  wire [7:0] p4_res7__44_comb;
  wire [7:0] p4_array_index_2044540_comb;
  wire [7:0] p4_array_index_2044541_comb;
  wire [7:0] p4_array_index_2044542_comb;
  wire [7:0] p4_res7__46_comb;
  wire [7:0] p4_array_index_2044553_comb;
  wire [7:0] p4_array_index_2044554_comb;
  wire [7:0] p4_res7__48_comb;
  wire [7:0] p4_array_index_2044564_comb;
  wire [7:0] p4_array_index_2044565_comb;
  wire [7:0] p4_res7__50_comb;
  assign p4_array_index_2044486_comb = p3_literal_2043912[p3_res7__34];
  assign p4_array_index_2044487_comb = p3_literal_2043914[p3_res7__32];
  assign p4_array_index_2044488_comb = p3_literal_2043916[p3_array_index_2044334];
  assign p4_array_index_2044489_comb = p3_literal_2043918[p3_array_index_2044335];
  assign p4_array_index_2044490_comb = p3_literal_2043920[p3_array_index_2044336];
  assign p4_res7__38_comb = p3_literal_2043910[p3_res7__36] ^ p4_array_index_2044486_comb ^ p4_array_index_2044487_comb ^ p4_array_index_2044488_comb ^ p4_array_index_2044489_comb ^ p4_array_index_2044490_comb ^ p3_array_index_2044337 ^ p3_literal_2043923[p3_array_index_2044338] ^ p3_array_index_2044339 ^ p3_literal_2043920[p3_array_index_2044356] ^ p3_literal_2043918[p3_array_index_2044341] ^ p3_literal_2043916[p3_array_index_2044358] ^ p3_literal_2043914[p3_array_index_2044343] ^ p3_literal_2043912[p3_array_index_2044344] ^ p3_literal_2043910[p3_array_index_2044345] ^ p3_array_index_2044346;
  assign p4_array_index_2044501_comb = p3_literal_2043914[p3_res7__34];
  assign p4_array_index_2044502_comb = p3_literal_2043916[p3_res7__32];
  assign p4_array_index_2044503_comb = p3_literal_2043918[p3_array_index_2044334];
  assign p4_array_index_2044504_comb = p3_literal_2043920[p3_array_index_2044335];
  assign p4_res7__40_comb = p3_literal_2043910[p4_res7__38_comb] ^ p3_literal_2043912[p3_res7__36] ^ p4_array_index_2044501_comb ^ p4_array_index_2044502_comb ^ p4_array_index_2044503_comb ^ p4_array_index_2044504_comb ^ p3_array_index_2044336 ^ p3_literal_2043923[p3_array_index_2044337] ^ p3_array_index_2044338 ^ p3_array_index_2044355 ^ p3_literal_2043918[p3_array_index_2044356] ^ p3_literal_2043916[p3_array_index_2044341] ^ p3_literal_2043914[p3_array_index_2044358] ^ p3_literal_2043912[p3_array_index_2044343] ^ p3_literal_2043910[p3_array_index_2044344] ^ p3_array_index_2044345;
  assign p4_array_index_2044514_comb = p3_literal_2043914[p3_res7__36];
  assign p4_array_index_2044515_comb = p3_literal_2043916[p3_res7__34];
  assign p4_array_index_2044516_comb = p3_literal_2043918[p3_res7__32];
  assign p4_array_index_2044517_comb = p3_literal_2043920[p3_array_index_2044334];
  assign p4_res7__42_comb = p3_literal_2043910[p4_res7__40_comb] ^ p3_literal_2043912[p4_res7__38_comb] ^ p4_array_index_2044514_comb ^ p4_array_index_2044515_comb ^ p4_array_index_2044516_comb ^ p4_array_index_2044517_comb ^ p3_array_index_2044335 ^ p3_literal_2043923[p3_array_index_2044336] ^ p3_array_index_2044337 ^ p3_array_index_2044372 ^ p3_literal_2043918[p3_array_index_2044339] ^ p3_literal_2043916[p3_array_index_2044356] ^ p3_literal_2043914[p3_array_index_2044341] ^ p3_literal_2043912[p3_array_index_2044358] ^ p3_literal_2043910[p3_array_index_2044343] ^ p3_array_index_2044344;
  assign p4_array_index_2044528_comb = p3_literal_2043916[p3_res7__36];
  assign p4_array_index_2044529_comb = p3_literal_2043918[p3_res7__34];
  assign p4_array_index_2044530_comb = p3_literal_2043920[p3_res7__32];
  assign p4_res7__44_comb = p3_literal_2043910[p4_res7__42_comb] ^ p3_literal_2043912[p4_res7__40_comb] ^ p3_literal_2043914[p4_res7__38_comb] ^ p4_array_index_2044528_comb ^ p4_array_index_2044529_comb ^ p4_array_index_2044530_comb ^ p3_array_index_2044334 ^ p3_literal_2043923[p3_array_index_2044335] ^ p3_array_index_2044336 ^ p3_array_index_2044386 ^ p3_array_index_2044354 ^ p3_literal_2043916[p3_array_index_2044339] ^ p3_literal_2043914[p3_array_index_2044356] ^ p3_literal_2043912[p3_array_index_2044341] ^ p3_literal_2043910[p3_array_index_2044358] ^ p3_array_index_2044343;
  assign p4_array_index_2044540_comb = p3_literal_2043916[p4_res7__38_comb];
  assign p4_array_index_2044541_comb = p3_literal_2043918[p3_res7__36];
  assign p4_array_index_2044542_comb = p3_literal_2043920[p3_res7__34];
  assign p4_res7__46_comb = p3_literal_2043910[p4_res7__44_comb] ^ p3_literal_2043912[p4_res7__42_comb] ^ p3_literal_2043914[p4_res7__40_comb] ^ p4_array_index_2044540_comb ^ p4_array_index_2044541_comb ^ p4_array_index_2044542_comb ^ p3_res7__32 ^ p3_literal_2043923[p3_array_index_2044334] ^ p3_array_index_2044335 ^ p4_array_index_2044490_comb ^ p3_array_index_2044371 ^ p3_literal_2043916[p3_array_index_2044338] ^ p3_literal_2043914[p3_array_index_2044339] ^ p3_literal_2043912[p3_array_index_2044356] ^ p3_literal_2043910[p3_array_index_2044341] ^ p3_array_index_2044358;
  assign p4_array_index_2044553_comb = p3_literal_2043918[p4_res7__38_comb];
  assign p4_array_index_2044554_comb = p3_literal_2043920[p3_res7__36];
  assign p4_res7__48_comb = p3_literal_2043910[p4_res7__46_comb] ^ p3_literal_2043912[p4_res7__44_comb] ^ p3_literal_2043914[p4_res7__42_comb] ^ p3_literal_2043916[p4_res7__40_comb] ^ p4_array_index_2044553_comb ^ p4_array_index_2044554_comb ^ p3_res7__34 ^ p3_literal_2043923[p3_res7__32] ^ p3_array_index_2044334 ^ p4_array_index_2044504_comb ^ p3_array_index_2044385 ^ p3_array_index_2044353 ^ p3_literal_2043914[p3_array_index_2044338] ^ p3_literal_2043912[p3_array_index_2044339] ^ p3_literal_2043910[p3_array_index_2044356] ^ p3_array_index_2044341;
  assign p4_array_index_2044564_comb = p3_literal_2043918[p4_res7__40_comb];
  assign p4_array_index_2044565_comb = p3_literal_2043920[p4_res7__38_comb];
  assign p4_res7__50_comb = p3_literal_2043910[p4_res7__48_comb] ^ p3_literal_2043912[p4_res7__46_comb] ^ p3_literal_2043914[p4_res7__44_comb] ^ p3_literal_2043916[p4_res7__42_comb] ^ p4_array_index_2044564_comb ^ p4_array_index_2044565_comb ^ p3_res7__36 ^ p3_literal_2043923[p3_res7__34] ^ p3_res7__32 ^ p4_array_index_2044517_comb ^ p4_array_index_2044489_comb ^ p3_array_index_2044370 ^ p3_literal_2043914[p3_array_index_2044337] ^ p3_literal_2043912[p3_array_index_2044338] ^ p3_literal_2043910[p3_array_index_2044339] ^ p3_array_index_2044356;

  // Registers for pipe stage 4:
  reg [127:0] p4_encoded;
  reg [127:0] p4_bit_slice_2043893;
  reg [127:0] p4_bit_slice_2044018;
  reg [127:0] p4_xor_2044318;
  reg [7:0] p4_array_index_2044334;
  reg [7:0] p4_array_index_2044335;
  reg [7:0] p4_array_index_2044336;
  reg [7:0] p4_array_index_2044337;
  reg [7:0] p4_array_index_2044338;
  reg [7:0] p4_array_index_2044339;
  reg [7:0] p4_array_index_2044350;
  reg [7:0] p4_array_index_2044351;
  reg [7:0] p4_array_index_2044352;
  reg [7:0] p4_res7__32;
  reg [7:0] p4_array_index_2044367;
  reg [7:0] p4_array_index_2044368;
  reg [7:0] p4_array_index_2044369;
  reg [7:0] p4_res7__34;
  reg [7:0] p4_array_index_2044382;
  reg [7:0] p4_array_index_2044383;
  reg [7:0] p4_array_index_2044384;
  reg [7:0] p4_res7__36;
  reg [7:0] p4_array_index_2044486;
  reg [7:0] p4_array_index_2044487;
  reg [7:0] p4_array_index_2044488;
  reg [7:0] p4_res7__38;
  reg [7:0] p4_array_index_2044501;
  reg [7:0] p4_array_index_2044502;
  reg [7:0] p4_array_index_2044503;
  reg [7:0] p4_res7__40;
  reg [7:0] p4_array_index_2044514;
  reg [7:0] p4_array_index_2044515;
  reg [7:0] p4_array_index_2044516;
  reg [7:0] p4_res7__42;
  reg [7:0] p4_array_index_2044528;
  reg [7:0] p4_array_index_2044529;
  reg [7:0] p4_array_index_2044530;
  reg [7:0] p4_res7__44;
  reg [7:0] p4_array_index_2044540;
  reg [7:0] p4_array_index_2044541;
  reg [7:0] p4_array_index_2044542;
  reg [7:0] p4_res7__46;
  reg [7:0] p4_array_index_2044553;
  reg [7:0] p4_array_index_2044554;
  reg [7:0] p4_res7__48;
  reg [7:0] p4_array_index_2044564;
  reg [7:0] p4_array_index_2044565;
  reg [7:0] p4_res7__50;
  reg [7:0] p5_literal_2043896[256];
  reg [7:0] p5_literal_2043910[256];
  reg [7:0] p5_literal_2043912[256];
  reg [7:0] p5_literal_2043914[256];
  reg [7:0] p5_literal_2043916[256];
  reg [7:0] p5_literal_2043918[256];
  reg [7:0] p5_literal_2043920[256];
  reg [7:0] p5_literal_2043923[256];
  reg [7:0] p82_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p4_encoded <= p3_encoded;
    p4_bit_slice_2043893 <= p3_bit_slice_2043893;
    p4_bit_slice_2044018 <= p3_bit_slice_2044018;
    p4_xor_2044318 <= p3_xor_2044318;
    p4_array_index_2044334 <= p3_array_index_2044334;
    p4_array_index_2044335 <= p3_array_index_2044335;
    p4_array_index_2044336 <= p3_array_index_2044336;
    p4_array_index_2044337 <= p3_array_index_2044337;
    p4_array_index_2044338 <= p3_array_index_2044338;
    p4_array_index_2044339 <= p3_array_index_2044339;
    p4_array_index_2044350 <= p3_array_index_2044350;
    p4_array_index_2044351 <= p3_array_index_2044351;
    p4_array_index_2044352 <= p3_array_index_2044352;
    p4_res7__32 <= p3_res7__32;
    p4_array_index_2044367 <= p3_array_index_2044367;
    p4_array_index_2044368 <= p3_array_index_2044368;
    p4_array_index_2044369 <= p3_array_index_2044369;
    p4_res7__34 <= p3_res7__34;
    p4_array_index_2044382 <= p3_array_index_2044382;
    p4_array_index_2044383 <= p3_array_index_2044383;
    p4_array_index_2044384 <= p3_array_index_2044384;
    p4_res7__36 <= p3_res7__36;
    p4_array_index_2044486 <= p4_array_index_2044486_comb;
    p4_array_index_2044487 <= p4_array_index_2044487_comb;
    p4_array_index_2044488 <= p4_array_index_2044488_comb;
    p4_res7__38 <= p4_res7__38_comb;
    p4_array_index_2044501 <= p4_array_index_2044501_comb;
    p4_array_index_2044502 <= p4_array_index_2044502_comb;
    p4_array_index_2044503 <= p4_array_index_2044503_comb;
    p4_res7__40 <= p4_res7__40_comb;
    p4_array_index_2044514 <= p4_array_index_2044514_comb;
    p4_array_index_2044515 <= p4_array_index_2044515_comb;
    p4_array_index_2044516 <= p4_array_index_2044516_comb;
    p4_res7__42 <= p4_res7__42_comb;
    p4_array_index_2044528 <= p4_array_index_2044528_comb;
    p4_array_index_2044529 <= p4_array_index_2044529_comb;
    p4_array_index_2044530 <= p4_array_index_2044530_comb;
    p4_res7__44 <= p4_res7__44_comb;
    p4_array_index_2044540 <= p4_array_index_2044540_comb;
    p4_array_index_2044541 <= p4_array_index_2044541_comb;
    p4_array_index_2044542 <= p4_array_index_2044542_comb;
    p4_res7__46 <= p4_res7__46_comb;
    p4_array_index_2044553 <= p4_array_index_2044553_comb;
    p4_array_index_2044554 <= p4_array_index_2044554_comb;
    p4_res7__48 <= p4_res7__48_comb;
    p4_array_index_2044564 <= p4_array_index_2044564_comb;
    p4_array_index_2044565 <= p4_array_index_2044565_comb;
    p4_res7__50 <= p4_res7__50_comb;
    p5_literal_2043896 <= p4_literal_2043896;
    p5_literal_2043910 <= p4_literal_2043910;
    p5_literal_2043912 <= p4_literal_2043912;
    p5_literal_2043914 <= p4_literal_2043914;
    p5_literal_2043916 <= p4_literal_2043916;
    p5_literal_2043918 <= p4_literal_2043918;
    p5_literal_2043920 <= p4_literal_2043920;
    p5_literal_2043923 <= p4_literal_2043923;
    p82_literal_2058836 <= p81_literal_2058836;
  end

  // ===== Pipe stage 5:
  wire [7:0] p5_array_index_2044688_comb;
  wire [7:0] p5_res7__52_comb;
  wire [7:0] p5_array_index_2044698_comb;
  wire [7:0] p5_res7__54_comb;
  wire [7:0] p5_res7__56_comb;
  wire [7:0] p5_res7__58_comb;
  wire [7:0] p5_res7__60_comb;
  wire [7:0] p5_res7__62_comb;
  wire [127:0] p5_res__1_comb;
  wire [127:0] p5_xor_2044738_comb;
  wire [127:0] p5_addedKey__34_comb;
  wire [7:0] p5_array_index_2044754_comb;
  wire [7:0] p5_array_index_2044755_comb;
  wire [7:0] p5_array_index_2044756_comb;
  wire [7:0] p5_array_index_2044757_comb;
  wire [7:0] p5_array_index_2044758_comb;
  wire [7:0] p5_array_index_2044759_comb;
  wire [7:0] p5_array_index_2044761_comb;
  wire [7:0] p5_array_index_2044763_comb;
  wire [7:0] p5_array_index_2044764_comb;
  wire [7:0] p5_array_index_2044765_comb;
  wire [7:0] p5_array_index_2044766_comb;
  wire [7:0] p5_array_index_2044767_comb;
  wire [7:0] p5_array_index_2044768_comb;
  wire [7:0] p5_array_index_2044770_comb;
  wire [7:0] p5_array_index_2044771_comb;
  wire [7:0] p5_array_index_2044772_comb;
  assign p5_array_index_2044688_comb = p4_literal_2043920[p4_res7__40];
  assign p5_res7__52_comb = p4_literal_2043910[p4_res7__50] ^ p4_literal_2043912[p4_res7__48] ^ p4_literal_2043914[p4_res7__46] ^ p4_literal_2043916[p4_res7__44] ^ p4_literal_2043918[p4_res7__42] ^ p5_array_index_2044688_comb ^ p4_res7__38 ^ p4_literal_2043923[p4_res7__36] ^ p4_res7__34 ^ p4_array_index_2044530 ^ p4_array_index_2044503 ^ p4_array_index_2044384 ^ p4_array_index_2044352 ^ p4_literal_2043912[p4_array_index_2044337] ^ p4_literal_2043910[p4_array_index_2044338] ^ p4_array_index_2044339;
  assign p5_array_index_2044698_comb = p4_literal_2043920[p4_res7__42];
  assign p5_res7__54_comb = p4_literal_2043910[p5_res7__52_comb] ^ p4_literal_2043912[p4_res7__50] ^ p4_literal_2043914[p4_res7__48] ^ p4_literal_2043916[p4_res7__46] ^ p4_literal_2043918[p4_res7__44] ^ p5_array_index_2044698_comb ^ p4_res7__40 ^ p4_literal_2043923[p4_res7__38] ^ p4_res7__36 ^ p4_array_index_2044542 ^ p4_array_index_2044516 ^ p4_array_index_2044488 ^ p4_array_index_2044369 ^ p4_literal_2043912[p4_array_index_2044336] ^ p4_literal_2043910[p4_array_index_2044337] ^ p4_array_index_2044338;
  assign p5_res7__56_comb = p4_literal_2043910[p5_res7__54_comb] ^ p4_literal_2043912[p5_res7__52_comb] ^ p4_literal_2043914[p4_res7__50] ^ p4_literal_2043916[p4_res7__48] ^ p4_literal_2043918[p4_res7__46] ^ p4_literal_2043920[p4_res7__44] ^ p4_res7__42 ^ p4_literal_2043923[p4_res7__40] ^ p4_res7__38 ^ p4_array_index_2044554 ^ p4_array_index_2044529 ^ p4_array_index_2044502 ^ p4_array_index_2044383 ^ p4_array_index_2044351 ^ p4_literal_2043910[p4_array_index_2044336] ^ p4_array_index_2044337;
  assign p5_res7__58_comb = p4_literal_2043910[p5_res7__56_comb] ^ p4_literal_2043912[p5_res7__54_comb] ^ p4_literal_2043914[p5_res7__52_comb] ^ p4_literal_2043916[p4_res7__50] ^ p4_literal_2043918[p4_res7__48] ^ p4_literal_2043920[p4_res7__46] ^ p4_res7__44 ^ p4_literal_2043923[p4_res7__42] ^ p4_res7__40 ^ p4_array_index_2044565 ^ p4_array_index_2044541 ^ p4_array_index_2044515 ^ p4_array_index_2044487 ^ p4_array_index_2044368 ^ p4_literal_2043910[p4_array_index_2044335] ^ p4_array_index_2044336;
  assign p5_res7__60_comb = p4_literal_2043910[p5_res7__58_comb] ^ p4_literal_2043912[p5_res7__56_comb] ^ p4_literal_2043914[p5_res7__54_comb] ^ p4_literal_2043916[p5_res7__52_comb] ^ p4_literal_2043918[p4_res7__50] ^ p4_literal_2043920[p4_res7__48] ^ p4_res7__46 ^ p4_literal_2043923[p4_res7__44] ^ p4_res7__42 ^ p5_array_index_2044688_comb ^ p4_array_index_2044553 ^ p4_array_index_2044528 ^ p4_array_index_2044501 ^ p4_array_index_2044382 ^ p4_array_index_2044350 ^ p4_array_index_2044335;
  assign p5_res7__62_comb = p4_literal_2043910[p5_res7__60_comb] ^ p4_literal_2043912[p5_res7__58_comb] ^ p4_literal_2043914[p5_res7__56_comb] ^ p4_literal_2043916[p5_res7__54_comb] ^ p4_literal_2043918[p5_res7__52_comb] ^ p4_literal_2043920[p4_res7__50] ^ p4_res7__48 ^ p4_literal_2043923[p4_res7__46] ^ p4_res7__44 ^ p5_array_index_2044698_comb ^ p4_array_index_2044564 ^ p4_array_index_2044540 ^ p4_array_index_2044514 ^ p4_array_index_2044486 ^ p4_array_index_2044367 ^ p4_array_index_2044334;
  assign p5_res__1_comb = {p5_res7__62_comb, p5_res7__60_comb, p5_res7__58_comb, p5_res7__56_comb, p5_res7__54_comb, p5_res7__52_comb, p4_res7__50, p4_res7__48, p4_res7__46, p4_res7__44, p4_res7__42, p4_res7__40, p4_res7__38, p4_res7__36, p4_res7__34, p4_res7__32};
  assign p5_xor_2044738_comb = p5_res__1_comb ^ p4_bit_slice_2043893;
  assign p5_addedKey__34_comb = p5_xor_2044738_comb ^ 128'hb225_9a96_b4d8_8e0b_e769_0430_a44f_7f03;
  assign p5_array_index_2044754_comb = p4_literal_2043896[p5_addedKey__34_comb[127:120]];
  assign p5_array_index_2044755_comb = p4_literal_2043896[p5_addedKey__34_comb[119:112]];
  assign p5_array_index_2044756_comb = p4_literal_2043896[p5_addedKey__34_comb[111:104]];
  assign p5_array_index_2044757_comb = p4_literal_2043896[p5_addedKey__34_comb[103:96]];
  assign p5_array_index_2044758_comb = p4_literal_2043896[p5_addedKey__34_comb[95:88]];
  assign p5_array_index_2044759_comb = p4_literal_2043896[p5_addedKey__34_comb[87:80]];
  assign p5_array_index_2044761_comb = p4_literal_2043896[p5_addedKey__34_comb[71:64]];
  assign p5_array_index_2044763_comb = p4_literal_2043896[p5_addedKey__34_comb[55:48]];
  assign p5_array_index_2044764_comb = p4_literal_2043896[p5_addedKey__34_comb[47:40]];
  assign p5_array_index_2044765_comb = p4_literal_2043896[p5_addedKey__34_comb[39:32]];
  assign p5_array_index_2044766_comb = p4_literal_2043896[p5_addedKey__34_comb[31:24]];
  assign p5_array_index_2044767_comb = p4_literal_2043896[p5_addedKey__34_comb[23:16]];
  assign p5_array_index_2044768_comb = p4_literal_2043896[p5_addedKey__34_comb[15:8]];
  assign p5_array_index_2044770_comb = p4_literal_2043896[p5_addedKey__34_comb[79:72]];
  assign p5_array_index_2044771_comb = p4_literal_2043896[p5_addedKey__34_comb[63:56]];
  assign p5_array_index_2044772_comb = p4_literal_2043896[p5_addedKey__34_comb[7:0]];

  // Registers for pipe stage 5:
  reg [127:0] p5_encoded;
  reg [127:0] p5_bit_slice_2043893;
  reg [127:0] p5_bit_slice_2044018;
  reg [127:0] p5_xor_2044318;
  reg [127:0] p5_xor_2044738;
  reg [7:0] p5_array_index_2044754;
  reg [7:0] p5_array_index_2044755;
  reg [7:0] p5_array_index_2044756;
  reg [7:0] p5_array_index_2044757;
  reg [7:0] p5_array_index_2044758;
  reg [7:0] p5_array_index_2044759;
  reg [7:0] p5_array_index_2044761;
  reg [7:0] p5_array_index_2044763;
  reg [7:0] p5_array_index_2044764;
  reg [7:0] p5_array_index_2044765;
  reg [7:0] p5_array_index_2044766;
  reg [7:0] p5_array_index_2044767;
  reg [7:0] p5_array_index_2044768;
  reg [7:0] p5_array_index_2044770;
  reg [7:0] p5_array_index_2044771;
  reg [7:0] p5_array_index_2044772;
  reg [7:0] p6_literal_2043896[256];
  reg [7:0] p6_literal_2043910[256];
  reg [7:0] p6_literal_2043912[256];
  reg [7:0] p6_literal_2043914[256];
  reg [7:0] p6_literal_2043916[256];
  reg [7:0] p6_literal_2043918[256];
  reg [7:0] p6_literal_2043920[256];
  reg [7:0] p6_literal_2043923[256];
  reg [7:0] p83_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p5_encoded <= p4_encoded;
    p5_bit_slice_2043893 <= p4_bit_slice_2043893;
    p5_bit_slice_2044018 <= p4_bit_slice_2044018;
    p5_xor_2044318 <= p4_xor_2044318;
    p5_xor_2044738 <= p5_xor_2044738_comb;
    p5_array_index_2044754 <= p5_array_index_2044754_comb;
    p5_array_index_2044755 <= p5_array_index_2044755_comb;
    p5_array_index_2044756 <= p5_array_index_2044756_comb;
    p5_array_index_2044757 <= p5_array_index_2044757_comb;
    p5_array_index_2044758 <= p5_array_index_2044758_comb;
    p5_array_index_2044759 <= p5_array_index_2044759_comb;
    p5_array_index_2044761 <= p5_array_index_2044761_comb;
    p5_array_index_2044763 <= p5_array_index_2044763_comb;
    p5_array_index_2044764 <= p5_array_index_2044764_comb;
    p5_array_index_2044765 <= p5_array_index_2044765_comb;
    p5_array_index_2044766 <= p5_array_index_2044766_comb;
    p5_array_index_2044767 <= p5_array_index_2044767_comb;
    p5_array_index_2044768 <= p5_array_index_2044768_comb;
    p5_array_index_2044770 <= p5_array_index_2044770_comb;
    p5_array_index_2044771 <= p5_array_index_2044771_comb;
    p5_array_index_2044772 <= p5_array_index_2044772_comb;
    p6_literal_2043896 <= p5_literal_2043896;
    p6_literal_2043910 <= p5_literal_2043910;
    p6_literal_2043912 <= p5_literal_2043912;
    p6_literal_2043914 <= p5_literal_2043914;
    p6_literal_2043916 <= p5_literal_2043916;
    p6_literal_2043918 <= p5_literal_2043918;
    p6_literal_2043920 <= p5_literal_2043920;
    p6_literal_2043923 <= p5_literal_2043923;
    p83_literal_2058836 <= p82_literal_2058836;
  end

  // ===== Pipe stage 6:
  wire [7:0] p6_array_index_2044831_comb;
  wire [7:0] p6_array_index_2044832_comb;
  wire [7:0] p6_array_index_2044833_comb;
  wire [7:0] p6_array_index_2044834_comb;
  wire [7:0] p6_array_index_2044835_comb;
  wire [7:0] p6_array_index_2044836_comb;
  wire [7:0] p6_res7__64_comb;
  wire [7:0] p6_array_index_2044845_comb;
  wire [7:0] p6_array_index_2044846_comb;
  wire [7:0] p6_array_index_2044847_comb;
  wire [7:0] p6_array_index_2044848_comb;
  wire [7:0] p6_array_index_2044849_comb;
  wire [7:0] p6_array_index_2044850_comb;
  wire [7:0] p6_res7__66_comb;
  wire [7:0] p6_array_index_2044860_comb;
  wire [7:0] p6_array_index_2044861_comb;
  wire [7:0] p6_array_index_2044862_comb;
  wire [7:0] p6_array_index_2044863_comb;
  wire [7:0] p6_array_index_2044864_comb;
  wire [7:0] p6_res7__68_comb;
  wire [7:0] p6_array_index_2044874_comb;
  wire [7:0] p6_array_index_2044875_comb;
  wire [7:0] p6_array_index_2044876_comb;
  wire [7:0] p6_array_index_2044877_comb;
  wire [7:0] p6_array_index_2044878_comb;
  wire [7:0] p6_res7__70_comb;
  wire [7:0] p6_array_index_2044889_comb;
  wire [7:0] p6_array_index_2044890_comb;
  wire [7:0] p6_array_index_2044891_comb;
  wire [7:0] p6_array_index_2044892_comb;
  wire [7:0] p6_res7__72_comb;
  wire [7:0] p6_array_index_2044902_comb;
  wire [7:0] p6_array_index_2044903_comb;
  wire [7:0] p6_array_index_2044904_comb;
  wire [7:0] p6_array_index_2044905_comb;
  wire [7:0] p6_res7__74_comb;
  wire [7:0] p6_array_index_2044916_comb;
  wire [7:0] p6_array_index_2044917_comb;
  wire [7:0] p6_array_index_2044918_comb;
  wire [7:0] p6_res7__76_comb;
  assign p6_array_index_2044831_comb = p5_literal_2043910[p5_array_index_2044754];
  assign p6_array_index_2044832_comb = p5_literal_2043912[p5_array_index_2044755];
  assign p6_array_index_2044833_comb = p5_literal_2043914[p5_array_index_2044756];
  assign p6_array_index_2044834_comb = p5_literal_2043916[p5_array_index_2044757];
  assign p6_array_index_2044835_comb = p5_literal_2043918[p5_array_index_2044758];
  assign p6_array_index_2044836_comb = p5_literal_2043920[p5_array_index_2044759];
  assign p6_res7__64_comb = p6_array_index_2044831_comb ^ p6_array_index_2044832_comb ^ p6_array_index_2044833_comb ^ p6_array_index_2044834_comb ^ p6_array_index_2044835_comb ^ p6_array_index_2044836_comb ^ p5_array_index_2044770 ^ p5_literal_2043923[p5_array_index_2044761] ^ p5_array_index_2044771 ^ p5_literal_2043920[p5_array_index_2044763] ^ p5_literal_2043918[p5_array_index_2044764] ^ p5_literal_2043916[p5_array_index_2044765] ^ p5_literal_2043914[p5_array_index_2044766] ^ p5_literal_2043912[p5_array_index_2044767] ^ p5_literal_2043910[p5_array_index_2044768] ^ p5_array_index_2044772;
  assign p6_array_index_2044845_comb = p5_literal_2043910[p6_res7__64_comb];
  assign p6_array_index_2044846_comb = p5_literal_2043912[p5_array_index_2044754];
  assign p6_array_index_2044847_comb = p5_literal_2043914[p5_array_index_2044755];
  assign p6_array_index_2044848_comb = p5_literal_2043916[p5_array_index_2044756];
  assign p6_array_index_2044849_comb = p5_literal_2043918[p5_array_index_2044757];
  assign p6_array_index_2044850_comb = p5_literal_2043920[p5_array_index_2044758];
  assign p6_res7__66_comb = p6_array_index_2044845_comb ^ p6_array_index_2044846_comb ^ p6_array_index_2044847_comb ^ p6_array_index_2044848_comb ^ p6_array_index_2044849_comb ^ p6_array_index_2044850_comb ^ p5_array_index_2044759 ^ p5_literal_2043923[p5_array_index_2044770] ^ p5_array_index_2044761 ^ p5_literal_2043920[p5_array_index_2044771] ^ p5_literal_2043918[p5_array_index_2044763] ^ p5_literal_2043916[p5_array_index_2044764] ^ p5_literal_2043914[p5_array_index_2044765] ^ p5_literal_2043912[p5_array_index_2044766] ^ p5_literal_2043910[p5_array_index_2044767] ^ p5_array_index_2044768;
  assign p6_array_index_2044860_comb = p5_literal_2043912[p6_res7__64_comb];
  assign p6_array_index_2044861_comb = p5_literal_2043914[p5_array_index_2044754];
  assign p6_array_index_2044862_comb = p5_literal_2043916[p5_array_index_2044755];
  assign p6_array_index_2044863_comb = p5_literal_2043918[p5_array_index_2044756];
  assign p6_array_index_2044864_comb = p5_literal_2043920[p5_array_index_2044757];
  assign p6_res7__68_comb = p5_literal_2043910[p6_res7__66_comb] ^ p6_array_index_2044860_comb ^ p6_array_index_2044861_comb ^ p6_array_index_2044862_comb ^ p6_array_index_2044863_comb ^ p6_array_index_2044864_comb ^ p5_array_index_2044758 ^ p5_literal_2043923[p5_array_index_2044759] ^ p5_array_index_2044770 ^ p5_literal_2043920[p5_array_index_2044761] ^ p5_literal_2043918[p5_array_index_2044771] ^ p5_literal_2043916[p5_array_index_2044763] ^ p5_literal_2043914[p5_array_index_2044764] ^ p5_literal_2043912[p5_array_index_2044765] ^ p5_literal_2043910[p5_array_index_2044766] ^ p5_array_index_2044767;
  assign p6_array_index_2044874_comb = p5_literal_2043912[p6_res7__66_comb];
  assign p6_array_index_2044875_comb = p5_literal_2043914[p6_res7__64_comb];
  assign p6_array_index_2044876_comb = p5_literal_2043916[p5_array_index_2044754];
  assign p6_array_index_2044877_comb = p5_literal_2043918[p5_array_index_2044755];
  assign p6_array_index_2044878_comb = p5_literal_2043920[p5_array_index_2044756];
  assign p6_res7__70_comb = p5_literal_2043910[p6_res7__68_comb] ^ p6_array_index_2044874_comb ^ p6_array_index_2044875_comb ^ p6_array_index_2044876_comb ^ p6_array_index_2044877_comb ^ p6_array_index_2044878_comb ^ p5_array_index_2044757 ^ p5_literal_2043923[p5_array_index_2044758] ^ p5_array_index_2044759 ^ p5_literal_2043920[p5_array_index_2044770] ^ p5_literal_2043918[p5_array_index_2044761] ^ p5_literal_2043916[p5_array_index_2044771] ^ p5_literal_2043914[p5_array_index_2044763] ^ p5_literal_2043912[p5_array_index_2044764] ^ p5_literal_2043910[p5_array_index_2044765] ^ p5_array_index_2044766;
  assign p6_array_index_2044889_comb = p5_literal_2043914[p6_res7__66_comb];
  assign p6_array_index_2044890_comb = p5_literal_2043916[p6_res7__64_comb];
  assign p6_array_index_2044891_comb = p5_literal_2043918[p5_array_index_2044754];
  assign p6_array_index_2044892_comb = p5_literal_2043920[p5_array_index_2044755];
  assign p6_res7__72_comb = p5_literal_2043910[p6_res7__70_comb] ^ p5_literal_2043912[p6_res7__68_comb] ^ p6_array_index_2044889_comb ^ p6_array_index_2044890_comb ^ p6_array_index_2044891_comb ^ p6_array_index_2044892_comb ^ p5_array_index_2044756 ^ p5_literal_2043923[p5_array_index_2044757] ^ p5_array_index_2044758 ^ p6_array_index_2044836_comb ^ p5_literal_2043918[p5_array_index_2044770] ^ p5_literal_2043916[p5_array_index_2044761] ^ p5_literal_2043914[p5_array_index_2044771] ^ p5_literal_2043912[p5_array_index_2044763] ^ p5_literal_2043910[p5_array_index_2044764] ^ p5_array_index_2044765;
  assign p6_array_index_2044902_comb = p5_literal_2043914[p6_res7__68_comb];
  assign p6_array_index_2044903_comb = p5_literal_2043916[p6_res7__66_comb];
  assign p6_array_index_2044904_comb = p5_literal_2043918[p6_res7__64_comb];
  assign p6_array_index_2044905_comb = p5_literal_2043920[p5_array_index_2044754];
  assign p6_res7__74_comb = p5_literal_2043910[p6_res7__72_comb] ^ p5_literal_2043912[p6_res7__70_comb] ^ p6_array_index_2044902_comb ^ p6_array_index_2044903_comb ^ p6_array_index_2044904_comb ^ p6_array_index_2044905_comb ^ p5_array_index_2044755 ^ p5_literal_2043923[p5_array_index_2044756] ^ p5_array_index_2044757 ^ p6_array_index_2044850_comb ^ p5_literal_2043918[p5_array_index_2044759] ^ p5_literal_2043916[p5_array_index_2044770] ^ p5_literal_2043914[p5_array_index_2044761] ^ p5_literal_2043912[p5_array_index_2044771] ^ p5_literal_2043910[p5_array_index_2044763] ^ p5_array_index_2044764;
  assign p6_array_index_2044916_comb = p5_literal_2043916[p6_res7__68_comb];
  assign p6_array_index_2044917_comb = p5_literal_2043918[p6_res7__66_comb];
  assign p6_array_index_2044918_comb = p5_literal_2043920[p6_res7__64_comb];
  assign p6_res7__76_comb = p5_literal_2043910[p6_res7__74_comb] ^ p5_literal_2043912[p6_res7__72_comb] ^ p5_literal_2043914[p6_res7__70_comb] ^ p6_array_index_2044916_comb ^ p6_array_index_2044917_comb ^ p6_array_index_2044918_comb ^ p5_array_index_2044754 ^ p5_literal_2043923[p5_array_index_2044755] ^ p5_array_index_2044756 ^ p6_array_index_2044864_comb ^ p6_array_index_2044835_comb ^ p5_literal_2043916[p5_array_index_2044759] ^ p5_literal_2043914[p5_array_index_2044770] ^ p5_literal_2043912[p5_array_index_2044761] ^ p5_literal_2043910[p5_array_index_2044771] ^ p5_array_index_2044763;

  // Registers for pipe stage 6:
  reg [127:0] p6_encoded;
  reg [127:0] p6_bit_slice_2043893;
  reg [127:0] p6_bit_slice_2044018;
  reg [127:0] p6_xor_2044318;
  reg [127:0] p6_xor_2044738;
  reg [7:0] p6_array_index_2044754;
  reg [7:0] p6_array_index_2044755;
  reg [7:0] p6_array_index_2044756;
  reg [7:0] p6_array_index_2044757;
  reg [7:0] p6_array_index_2044758;
  reg [7:0] p6_array_index_2044759;
  reg [7:0] p6_array_index_2044761;
  reg [7:0] p6_array_index_2044831;
  reg [7:0] p6_array_index_2044832;
  reg [7:0] p6_array_index_2044833;
  reg [7:0] p6_array_index_2044834;
  reg [7:0] p6_array_index_2044770;
  reg [7:0] p6_array_index_2044771;
  reg [7:0] p6_res7__64;
  reg [7:0] p6_array_index_2044845;
  reg [7:0] p6_array_index_2044846;
  reg [7:0] p6_array_index_2044847;
  reg [7:0] p6_array_index_2044848;
  reg [7:0] p6_array_index_2044849;
  reg [7:0] p6_res7__66;
  reg [7:0] p6_array_index_2044860;
  reg [7:0] p6_array_index_2044861;
  reg [7:0] p6_array_index_2044862;
  reg [7:0] p6_array_index_2044863;
  reg [7:0] p6_res7__68;
  reg [7:0] p6_array_index_2044874;
  reg [7:0] p6_array_index_2044875;
  reg [7:0] p6_array_index_2044876;
  reg [7:0] p6_array_index_2044877;
  reg [7:0] p6_array_index_2044878;
  reg [7:0] p6_res7__70;
  reg [7:0] p6_array_index_2044889;
  reg [7:0] p6_array_index_2044890;
  reg [7:0] p6_array_index_2044891;
  reg [7:0] p6_array_index_2044892;
  reg [7:0] p6_res7__72;
  reg [7:0] p6_array_index_2044902;
  reg [7:0] p6_array_index_2044903;
  reg [7:0] p6_array_index_2044904;
  reg [7:0] p6_array_index_2044905;
  reg [7:0] p6_res7__74;
  reg [7:0] p6_array_index_2044916;
  reg [7:0] p6_array_index_2044917;
  reg [7:0] p6_array_index_2044918;
  reg [7:0] p6_res7__76;
  reg [7:0] p7_literal_2043896[256];
  reg [7:0] p7_literal_2043910[256];
  reg [7:0] p7_literal_2043912[256];
  reg [7:0] p7_literal_2043914[256];
  reg [7:0] p7_literal_2043916[256];
  reg [7:0] p7_literal_2043918[256];
  reg [7:0] p7_literal_2043920[256];
  reg [7:0] p7_literal_2043923[256];
  reg [7:0] p84_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p6_encoded <= p5_encoded;
    p6_bit_slice_2043893 <= p5_bit_slice_2043893;
    p6_bit_slice_2044018 <= p5_bit_slice_2044018;
    p6_xor_2044318 <= p5_xor_2044318;
    p6_xor_2044738 <= p5_xor_2044738;
    p6_array_index_2044754 <= p5_array_index_2044754;
    p6_array_index_2044755 <= p5_array_index_2044755;
    p6_array_index_2044756 <= p5_array_index_2044756;
    p6_array_index_2044757 <= p5_array_index_2044757;
    p6_array_index_2044758 <= p5_array_index_2044758;
    p6_array_index_2044759 <= p5_array_index_2044759;
    p6_array_index_2044761 <= p5_array_index_2044761;
    p6_array_index_2044831 <= p6_array_index_2044831_comb;
    p6_array_index_2044832 <= p6_array_index_2044832_comb;
    p6_array_index_2044833 <= p6_array_index_2044833_comb;
    p6_array_index_2044834 <= p6_array_index_2044834_comb;
    p6_array_index_2044770 <= p5_array_index_2044770;
    p6_array_index_2044771 <= p5_array_index_2044771;
    p6_res7__64 <= p6_res7__64_comb;
    p6_array_index_2044845 <= p6_array_index_2044845_comb;
    p6_array_index_2044846 <= p6_array_index_2044846_comb;
    p6_array_index_2044847 <= p6_array_index_2044847_comb;
    p6_array_index_2044848 <= p6_array_index_2044848_comb;
    p6_array_index_2044849 <= p6_array_index_2044849_comb;
    p6_res7__66 <= p6_res7__66_comb;
    p6_array_index_2044860 <= p6_array_index_2044860_comb;
    p6_array_index_2044861 <= p6_array_index_2044861_comb;
    p6_array_index_2044862 <= p6_array_index_2044862_comb;
    p6_array_index_2044863 <= p6_array_index_2044863_comb;
    p6_res7__68 <= p6_res7__68_comb;
    p6_array_index_2044874 <= p6_array_index_2044874_comb;
    p6_array_index_2044875 <= p6_array_index_2044875_comb;
    p6_array_index_2044876 <= p6_array_index_2044876_comb;
    p6_array_index_2044877 <= p6_array_index_2044877_comb;
    p6_array_index_2044878 <= p6_array_index_2044878_comb;
    p6_res7__70 <= p6_res7__70_comb;
    p6_array_index_2044889 <= p6_array_index_2044889_comb;
    p6_array_index_2044890 <= p6_array_index_2044890_comb;
    p6_array_index_2044891 <= p6_array_index_2044891_comb;
    p6_array_index_2044892 <= p6_array_index_2044892_comb;
    p6_res7__72 <= p6_res7__72_comb;
    p6_array_index_2044902 <= p6_array_index_2044902_comb;
    p6_array_index_2044903 <= p6_array_index_2044903_comb;
    p6_array_index_2044904 <= p6_array_index_2044904_comb;
    p6_array_index_2044905 <= p6_array_index_2044905_comb;
    p6_res7__74 <= p6_res7__74_comb;
    p6_array_index_2044916 <= p6_array_index_2044916_comb;
    p6_array_index_2044917 <= p6_array_index_2044917_comb;
    p6_array_index_2044918 <= p6_array_index_2044918_comb;
    p6_res7__76 <= p6_res7__76_comb;
    p7_literal_2043896 <= p6_literal_2043896;
    p7_literal_2043910 <= p6_literal_2043910;
    p7_literal_2043912 <= p6_literal_2043912;
    p7_literal_2043914 <= p6_literal_2043914;
    p7_literal_2043916 <= p6_literal_2043916;
    p7_literal_2043918 <= p6_literal_2043918;
    p7_literal_2043920 <= p6_literal_2043920;
    p7_literal_2043923 <= p6_literal_2043923;
    p84_literal_2058836 <= p83_literal_2058836;
  end

  // ===== Pipe stage 7:
  wire [7:0] p7_array_index_2045044_comb;
  wire [7:0] p7_array_index_2045045_comb;
  wire [7:0] p7_array_index_2045046_comb;
  wire [7:0] p7_res7__78_comb;
  wire [7:0] p7_array_index_2045057_comb;
  wire [7:0] p7_array_index_2045058_comb;
  wire [7:0] p7_res7__80_comb;
  wire [7:0] p7_array_index_2045068_comb;
  wire [7:0] p7_array_index_2045069_comb;
  wire [7:0] p7_res7__82_comb;
  wire [7:0] p7_array_index_2045080_comb;
  wire [7:0] p7_res7__84_comb;
  wire [7:0] p7_array_index_2045090_comb;
  wire [7:0] p7_res7__86_comb;
  wire [7:0] p7_res7__88_comb;
  wire [7:0] p7_res7__90_comb;
  assign p7_array_index_2045044_comb = p6_literal_2043916[p6_res7__70];
  assign p7_array_index_2045045_comb = p6_literal_2043918[p6_res7__68];
  assign p7_array_index_2045046_comb = p6_literal_2043920[p6_res7__66];
  assign p7_res7__78_comb = p6_literal_2043910[p6_res7__76] ^ p6_literal_2043912[p6_res7__74] ^ p6_literal_2043914[p6_res7__72] ^ p7_array_index_2045044_comb ^ p7_array_index_2045045_comb ^ p7_array_index_2045046_comb ^ p6_res7__64 ^ p6_literal_2043923[p6_array_index_2044754] ^ p6_array_index_2044755 ^ p6_array_index_2044878 ^ p6_array_index_2044849 ^ p6_literal_2043916[p6_array_index_2044758] ^ p6_literal_2043914[p6_array_index_2044759] ^ p6_literal_2043912[p6_array_index_2044770] ^ p6_literal_2043910[p6_array_index_2044761] ^ p6_array_index_2044771;
  assign p7_array_index_2045057_comb = p6_literal_2043918[p6_res7__70];
  assign p7_array_index_2045058_comb = p6_literal_2043920[p6_res7__68];
  assign p7_res7__80_comb = p6_literal_2043910[p7_res7__78_comb] ^ p6_literal_2043912[p6_res7__76] ^ p6_literal_2043914[p6_res7__74] ^ p6_literal_2043916[p6_res7__72] ^ p7_array_index_2045057_comb ^ p7_array_index_2045058_comb ^ p6_res7__66 ^ p6_literal_2043923[p6_res7__64] ^ p6_array_index_2044754 ^ p6_array_index_2044892 ^ p6_array_index_2044863 ^ p6_array_index_2044834 ^ p6_literal_2043914[p6_array_index_2044758] ^ p6_literal_2043912[p6_array_index_2044759] ^ p6_literal_2043910[p6_array_index_2044770] ^ p6_array_index_2044761;
  assign p7_array_index_2045068_comb = p6_literal_2043918[p6_res7__72];
  assign p7_array_index_2045069_comb = p6_literal_2043920[p6_res7__70];
  assign p7_res7__82_comb = p6_literal_2043910[p7_res7__80_comb] ^ p6_literal_2043912[p7_res7__78_comb] ^ p6_literal_2043914[p6_res7__76] ^ p6_literal_2043916[p6_res7__74] ^ p7_array_index_2045068_comb ^ p7_array_index_2045069_comb ^ p6_res7__68 ^ p6_literal_2043923[p6_res7__66] ^ p6_res7__64 ^ p6_array_index_2044905 ^ p6_array_index_2044877 ^ p6_array_index_2044848 ^ p6_literal_2043914[p6_array_index_2044757] ^ p6_literal_2043912[p6_array_index_2044758] ^ p6_literal_2043910[p6_array_index_2044759] ^ p6_array_index_2044770;
  assign p7_array_index_2045080_comb = p6_literal_2043920[p6_res7__72];
  assign p7_res7__84_comb = p6_literal_2043910[p7_res7__82_comb] ^ p6_literal_2043912[p7_res7__80_comb] ^ p6_literal_2043914[p7_res7__78_comb] ^ p6_literal_2043916[p6_res7__76] ^ p6_literal_2043918[p6_res7__74] ^ p7_array_index_2045080_comb ^ p6_res7__70 ^ p6_literal_2043923[p6_res7__68] ^ p6_res7__66 ^ p6_array_index_2044918 ^ p6_array_index_2044891 ^ p6_array_index_2044862 ^ p6_array_index_2044833 ^ p6_literal_2043912[p6_array_index_2044757] ^ p6_literal_2043910[p6_array_index_2044758] ^ p6_array_index_2044759;
  assign p7_array_index_2045090_comb = p6_literal_2043920[p6_res7__74];
  assign p7_res7__86_comb = p6_literal_2043910[p7_res7__84_comb] ^ p6_literal_2043912[p7_res7__82_comb] ^ p6_literal_2043914[p7_res7__80_comb] ^ p6_literal_2043916[p7_res7__78_comb] ^ p6_literal_2043918[p6_res7__76] ^ p7_array_index_2045090_comb ^ p6_res7__72 ^ p6_literal_2043923[p6_res7__70] ^ p6_res7__68 ^ p7_array_index_2045046_comb ^ p6_array_index_2044904 ^ p6_array_index_2044876 ^ p6_array_index_2044847 ^ p6_literal_2043912[p6_array_index_2044756] ^ p6_literal_2043910[p6_array_index_2044757] ^ p6_array_index_2044758;
  assign p7_res7__88_comb = p6_literal_2043910[p7_res7__86_comb] ^ p6_literal_2043912[p7_res7__84_comb] ^ p6_literal_2043914[p7_res7__82_comb] ^ p6_literal_2043916[p7_res7__80_comb] ^ p6_literal_2043918[p7_res7__78_comb] ^ p6_literal_2043920[p6_res7__76] ^ p6_res7__74 ^ p6_literal_2043923[p6_res7__72] ^ p6_res7__70 ^ p7_array_index_2045058_comb ^ p6_array_index_2044917 ^ p6_array_index_2044890 ^ p6_array_index_2044861 ^ p6_array_index_2044832 ^ p6_literal_2043910[p6_array_index_2044756] ^ p6_array_index_2044757;
  assign p7_res7__90_comb = p6_literal_2043910[p7_res7__88_comb] ^ p6_literal_2043912[p7_res7__86_comb] ^ p6_literal_2043914[p7_res7__84_comb] ^ p6_literal_2043916[p7_res7__82_comb] ^ p6_literal_2043918[p7_res7__80_comb] ^ p6_literal_2043920[p7_res7__78_comb] ^ p6_res7__76 ^ p6_literal_2043923[p6_res7__74] ^ p6_res7__72 ^ p7_array_index_2045069_comb ^ p7_array_index_2045045_comb ^ p6_array_index_2044903 ^ p6_array_index_2044875 ^ p6_array_index_2044846 ^ p6_literal_2043910[p6_array_index_2044755] ^ p6_array_index_2044756;

  // Registers for pipe stage 7:
  reg [127:0] p7_encoded;
  reg [127:0] p7_bit_slice_2043893;
  reg [127:0] p7_bit_slice_2044018;
  reg [127:0] p7_xor_2044318;
  reg [127:0] p7_xor_2044738;
  reg [7:0] p7_array_index_2044754;
  reg [7:0] p7_array_index_2044755;
  reg [7:0] p7_array_index_2044831;
  reg [7:0] p7_res7__64;
  reg [7:0] p7_array_index_2044845;
  reg [7:0] p7_res7__66;
  reg [7:0] p7_array_index_2044860;
  reg [7:0] p7_res7__68;
  reg [7:0] p7_array_index_2044874;
  reg [7:0] p7_res7__70;
  reg [7:0] p7_array_index_2044889;
  reg [7:0] p7_res7__72;
  reg [7:0] p7_array_index_2044902;
  reg [7:0] p7_res7__74;
  reg [7:0] p7_array_index_2044916;
  reg [7:0] p7_res7__76;
  reg [7:0] p7_array_index_2045044;
  reg [7:0] p7_res7__78;
  reg [7:0] p7_array_index_2045057;
  reg [7:0] p7_res7__80;
  reg [7:0] p7_array_index_2045068;
  reg [7:0] p7_res7__82;
  reg [7:0] p7_array_index_2045080;
  reg [7:0] p7_res7__84;
  reg [7:0] p7_array_index_2045090;
  reg [7:0] p7_res7__86;
  reg [7:0] p7_res7__88;
  reg [7:0] p7_res7__90;
  reg [7:0] p8_literal_2043896[256];
  reg [7:0] p8_literal_2043910[256];
  reg [7:0] p8_literal_2043912[256];
  reg [7:0] p8_literal_2043914[256];
  reg [7:0] p8_literal_2043916[256];
  reg [7:0] p8_literal_2043918[256];
  reg [7:0] p8_literal_2043920[256];
  reg [7:0] p8_literal_2043923[256];
  reg [7:0] p85_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p7_encoded <= p6_encoded;
    p7_bit_slice_2043893 <= p6_bit_slice_2043893;
    p7_bit_slice_2044018 <= p6_bit_slice_2044018;
    p7_xor_2044318 <= p6_xor_2044318;
    p7_xor_2044738 <= p6_xor_2044738;
    p7_array_index_2044754 <= p6_array_index_2044754;
    p7_array_index_2044755 <= p6_array_index_2044755;
    p7_array_index_2044831 <= p6_array_index_2044831;
    p7_res7__64 <= p6_res7__64;
    p7_array_index_2044845 <= p6_array_index_2044845;
    p7_res7__66 <= p6_res7__66;
    p7_array_index_2044860 <= p6_array_index_2044860;
    p7_res7__68 <= p6_res7__68;
    p7_array_index_2044874 <= p6_array_index_2044874;
    p7_res7__70 <= p6_res7__70;
    p7_array_index_2044889 <= p6_array_index_2044889;
    p7_res7__72 <= p6_res7__72;
    p7_array_index_2044902 <= p6_array_index_2044902;
    p7_res7__74 <= p6_res7__74;
    p7_array_index_2044916 <= p6_array_index_2044916;
    p7_res7__76 <= p6_res7__76;
    p7_array_index_2045044 <= p7_array_index_2045044_comb;
    p7_res7__78 <= p7_res7__78_comb;
    p7_array_index_2045057 <= p7_array_index_2045057_comb;
    p7_res7__80 <= p7_res7__80_comb;
    p7_array_index_2045068 <= p7_array_index_2045068_comb;
    p7_res7__82 <= p7_res7__82_comb;
    p7_array_index_2045080 <= p7_array_index_2045080_comb;
    p7_res7__84 <= p7_res7__84_comb;
    p7_array_index_2045090 <= p7_array_index_2045090_comb;
    p7_res7__86 <= p7_res7__86_comb;
    p7_res7__88 <= p7_res7__88_comb;
    p7_res7__90 <= p7_res7__90_comb;
    p8_literal_2043896 <= p7_literal_2043896;
    p8_literal_2043910 <= p7_literal_2043910;
    p8_literal_2043912 <= p7_literal_2043912;
    p8_literal_2043914 <= p7_literal_2043914;
    p8_literal_2043916 <= p7_literal_2043916;
    p8_literal_2043918 <= p7_literal_2043918;
    p8_literal_2043920 <= p7_literal_2043920;
    p8_literal_2043923 <= p7_literal_2043923;
    p85_literal_2058836 <= p84_literal_2058836;
  end

  // ===== Pipe stage 8:
  wire [7:0] p8_res7__92_comb;
  wire [7:0] p8_res7__94_comb;
  wire [127:0] p8_res__2_comb;
  wire [127:0] p8_xor_2045212_comb;
  wire [127:0] p8_addedKey__35_comb;
  wire [7:0] p8_array_index_2045228_comb;
  wire [7:0] p8_array_index_2045229_comb;
  wire [7:0] p8_array_index_2045230_comb;
  wire [7:0] p8_array_index_2045231_comb;
  wire [7:0] p8_array_index_2045232_comb;
  wire [7:0] p8_array_index_2045233_comb;
  wire [7:0] p8_array_index_2045235_comb;
  wire [7:0] p8_array_index_2045237_comb;
  wire [7:0] p8_array_index_2045238_comb;
  wire [7:0] p8_array_index_2045239_comb;
  wire [7:0] p8_array_index_2045240_comb;
  wire [7:0] p8_array_index_2045241_comb;
  wire [7:0] p8_array_index_2045242_comb;
  wire [7:0] p8_array_index_2045244_comb;
  wire [7:0] p8_array_index_2045245_comb;
  wire [7:0] p8_array_index_2045246_comb;
  wire [7:0] p8_array_index_2045247_comb;
  wire [7:0] p8_array_index_2045248_comb;
  wire [7:0] p8_array_index_2045249_comb;
  wire [7:0] p8_array_index_2045250_comb;
  wire [7:0] p8_array_index_2045252_comb;
  wire [7:0] p8_res7__96_comb;
  wire [7:0] p8_array_index_2045261_comb;
  wire [7:0] p8_array_index_2045262_comb;
  wire [7:0] p8_array_index_2045263_comb;
  wire [7:0] p8_array_index_2045264_comb;
  wire [7:0] p8_array_index_2045265_comb;
  wire [7:0] p8_array_index_2045266_comb;
  wire [7:0] p8_res7__98_comb;
  wire [7:0] p8_array_index_2045276_comb;
  wire [7:0] p8_array_index_2045277_comb;
  wire [7:0] p8_array_index_2045278_comb;
  wire [7:0] p8_array_index_2045279_comb;
  wire [7:0] p8_array_index_2045280_comb;
  wire [7:0] p8_res7__100_comb;
  wire [7:0] p8_array_index_2045290_comb;
  wire [7:0] p8_array_index_2045291_comb;
  wire [7:0] p8_array_index_2045292_comb;
  wire [7:0] p8_array_index_2045293_comb;
  wire [7:0] p8_array_index_2045294_comb;
  wire [7:0] p8_res7__102_comb;
  assign p8_res7__92_comb = p7_literal_2043910[p7_res7__90] ^ p7_literal_2043912[p7_res7__88] ^ p7_literal_2043914[p7_res7__86] ^ p7_literal_2043916[p7_res7__84] ^ p7_literal_2043918[p7_res7__82] ^ p7_literal_2043920[p7_res7__80] ^ p7_res7__78 ^ p7_literal_2043923[p7_res7__76] ^ p7_res7__74 ^ p7_array_index_2045080 ^ p7_array_index_2045057 ^ p7_array_index_2044916 ^ p7_array_index_2044889 ^ p7_array_index_2044860 ^ p7_array_index_2044831 ^ p7_array_index_2044755;
  assign p8_res7__94_comb = p7_literal_2043910[p8_res7__92_comb] ^ p7_literal_2043912[p7_res7__90] ^ p7_literal_2043914[p7_res7__88] ^ p7_literal_2043916[p7_res7__86] ^ p7_literal_2043918[p7_res7__84] ^ p7_literal_2043920[p7_res7__82] ^ p7_res7__80 ^ p7_literal_2043923[p7_res7__78] ^ p7_res7__76 ^ p7_array_index_2045090 ^ p7_array_index_2045068 ^ p7_array_index_2045044 ^ p7_array_index_2044902 ^ p7_array_index_2044874 ^ p7_array_index_2044845 ^ p7_array_index_2044754;
  assign p8_res__2_comb = {p8_res7__94_comb, p8_res7__92_comb, p7_res7__90, p7_res7__88, p7_res7__86, p7_res7__84, p7_res7__82, p7_res7__80, p7_res7__78, p7_res7__76, p7_res7__74, p7_res7__72, p7_res7__70, p7_res7__68, p7_res7__66, p7_res7__64};
  assign p8_xor_2045212_comb = p8_res__2_comb ^ p7_xor_2044318;
  assign p8_addedKey__35_comb = p8_xor_2045212_comb ^ 128'h7bcd_1b0b_73e3_2ba5_b79c_b140_f255_1504;
  assign p8_array_index_2045228_comb = p7_literal_2043896[p8_addedKey__35_comb[127:120]];
  assign p8_array_index_2045229_comb = p7_literal_2043896[p8_addedKey__35_comb[119:112]];
  assign p8_array_index_2045230_comb = p7_literal_2043896[p8_addedKey__35_comb[111:104]];
  assign p8_array_index_2045231_comb = p7_literal_2043896[p8_addedKey__35_comb[103:96]];
  assign p8_array_index_2045232_comb = p7_literal_2043896[p8_addedKey__35_comb[95:88]];
  assign p8_array_index_2045233_comb = p7_literal_2043896[p8_addedKey__35_comb[87:80]];
  assign p8_array_index_2045235_comb = p7_literal_2043896[p8_addedKey__35_comb[71:64]];
  assign p8_array_index_2045237_comb = p7_literal_2043896[p8_addedKey__35_comb[55:48]];
  assign p8_array_index_2045238_comb = p7_literal_2043896[p8_addedKey__35_comb[47:40]];
  assign p8_array_index_2045239_comb = p7_literal_2043896[p8_addedKey__35_comb[39:32]];
  assign p8_array_index_2045240_comb = p7_literal_2043896[p8_addedKey__35_comb[31:24]];
  assign p8_array_index_2045241_comb = p7_literal_2043896[p8_addedKey__35_comb[23:16]];
  assign p8_array_index_2045242_comb = p7_literal_2043896[p8_addedKey__35_comb[15:8]];
  assign p8_array_index_2045244_comb = p7_literal_2043910[p8_array_index_2045228_comb];
  assign p8_array_index_2045245_comb = p7_literal_2043912[p8_array_index_2045229_comb];
  assign p8_array_index_2045246_comb = p7_literal_2043914[p8_array_index_2045230_comb];
  assign p8_array_index_2045247_comb = p7_literal_2043916[p8_array_index_2045231_comb];
  assign p8_array_index_2045248_comb = p7_literal_2043918[p8_array_index_2045232_comb];
  assign p8_array_index_2045249_comb = p7_literal_2043920[p8_array_index_2045233_comb];
  assign p8_array_index_2045250_comb = p7_literal_2043896[p8_addedKey__35_comb[79:72]];
  assign p8_array_index_2045252_comb = p7_literal_2043896[p8_addedKey__35_comb[63:56]];
  assign p8_res7__96_comb = p8_array_index_2045244_comb ^ p8_array_index_2045245_comb ^ p8_array_index_2045246_comb ^ p8_array_index_2045247_comb ^ p8_array_index_2045248_comb ^ p8_array_index_2045249_comb ^ p8_array_index_2045250_comb ^ p7_literal_2043923[p8_array_index_2045235_comb] ^ p8_array_index_2045252_comb ^ p7_literal_2043920[p8_array_index_2045237_comb] ^ p7_literal_2043918[p8_array_index_2045238_comb] ^ p7_literal_2043916[p8_array_index_2045239_comb] ^ p7_literal_2043914[p8_array_index_2045240_comb] ^ p7_literal_2043912[p8_array_index_2045241_comb] ^ p7_literal_2043910[p8_array_index_2045242_comb] ^ p7_literal_2043896[p8_addedKey__35_comb[7:0]];
  assign p8_array_index_2045261_comb = p7_literal_2043910[p8_res7__96_comb];
  assign p8_array_index_2045262_comb = p7_literal_2043912[p8_array_index_2045228_comb];
  assign p8_array_index_2045263_comb = p7_literal_2043914[p8_array_index_2045229_comb];
  assign p8_array_index_2045264_comb = p7_literal_2043916[p8_array_index_2045230_comb];
  assign p8_array_index_2045265_comb = p7_literal_2043918[p8_array_index_2045231_comb];
  assign p8_array_index_2045266_comb = p7_literal_2043920[p8_array_index_2045232_comb];
  assign p8_res7__98_comb = p8_array_index_2045261_comb ^ p8_array_index_2045262_comb ^ p8_array_index_2045263_comb ^ p8_array_index_2045264_comb ^ p8_array_index_2045265_comb ^ p8_array_index_2045266_comb ^ p8_array_index_2045233_comb ^ p7_literal_2043923[p8_array_index_2045250_comb] ^ p8_array_index_2045235_comb ^ p7_literal_2043920[p8_array_index_2045252_comb] ^ p7_literal_2043918[p8_array_index_2045237_comb] ^ p7_literal_2043916[p8_array_index_2045238_comb] ^ p7_literal_2043914[p8_array_index_2045239_comb] ^ p7_literal_2043912[p8_array_index_2045240_comb] ^ p7_literal_2043910[p8_array_index_2045241_comb] ^ p8_array_index_2045242_comb;
  assign p8_array_index_2045276_comb = p7_literal_2043912[p8_res7__96_comb];
  assign p8_array_index_2045277_comb = p7_literal_2043914[p8_array_index_2045228_comb];
  assign p8_array_index_2045278_comb = p7_literal_2043916[p8_array_index_2045229_comb];
  assign p8_array_index_2045279_comb = p7_literal_2043918[p8_array_index_2045230_comb];
  assign p8_array_index_2045280_comb = p7_literal_2043920[p8_array_index_2045231_comb];
  assign p8_res7__100_comb = p7_literal_2043910[p8_res7__98_comb] ^ p8_array_index_2045276_comb ^ p8_array_index_2045277_comb ^ p8_array_index_2045278_comb ^ p8_array_index_2045279_comb ^ p8_array_index_2045280_comb ^ p8_array_index_2045232_comb ^ p7_literal_2043923[p8_array_index_2045233_comb] ^ p8_array_index_2045250_comb ^ p7_literal_2043920[p8_array_index_2045235_comb] ^ p7_literal_2043918[p8_array_index_2045252_comb] ^ p7_literal_2043916[p8_array_index_2045237_comb] ^ p7_literal_2043914[p8_array_index_2045238_comb] ^ p7_literal_2043912[p8_array_index_2045239_comb] ^ p7_literal_2043910[p8_array_index_2045240_comb] ^ p8_array_index_2045241_comb;
  assign p8_array_index_2045290_comb = p7_literal_2043912[p8_res7__98_comb];
  assign p8_array_index_2045291_comb = p7_literal_2043914[p8_res7__96_comb];
  assign p8_array_index_2045292_comb = p7_literal_2043916[p8_array_index_2045228_comb];
  assign p8_array_index_2045293_comb = p7_literal_2043918[p8_array_index_2045229_comb];
  assign p8_array_index_2045294_comb = p7_literal_2043920[p8_array_index_2045230_comb];
  assign p8_res7__102_comb = p7_literal_2043910[p8_res7__100_comb] ^ p8_array_index_2045290_comb ^ p8_array_index_2045291_comb ^ p8_array_index_2045292_comb ^ p8_array_index_2045293_comb ^ p8_array_index_2045294_comb ^ p8_array_index_2045231_comb ^ p7_literal_2043923[p8_array_index_2045232_comb] ^ p8_array_index_2045233_comb ^ p7_literal_2043920[p8_array_index_2045250_comb] ^ p7_literal_2043918[p8_array_index_2045235_comb] ^ p7_literal_2043916[p8_array_index_2045252_comb] ^ p7_literal_2043914[p8_array_index_2045237_comb] ^ p7_literal_2043912[p8_array_index_2045238_comb] ^ p7_literal_2043910[p8_array_index_2045239_comb] ^ p8_array_index_2045240_comb;

  // Registers for pipe stage 8:
  reg [127:0] p8_encoded;
  reg [127:0] p8_bit_slice_2043893;
  reg [127:0] p8_bit_slice_2044018;
  reg [127:0] p8_xor_2044738;
  reg [127:0] p8_xor_2045212;
  reg [7:0] p8_array_index_2045228;
  reg [7:0] p8_array_index_2045229;
  reg [7:0] p8_array_index_2045230;
  reg [7:0] p8_array_index_2045231;
  reg [7:0] p8_array_index_2045232;
  reg [7:0] p8_array_index_2045233;
  reg [7:0] p8_array_index_2045235;
  reg [7:0] p8_array_index_2045237;
  reg [7:0] p8_array_index_2045238;
  reg [7:0] p8_array_index_2045239;
  reg [7:0] p8_array_index_2045244;
  reg [7:0] p8_array_index_2045245;
  reg [7:0] p8_array_index_2045246;
  reg [7:0] p8_array_index_2045247;
  reg [7:0] p8_array_index_2045248;
  reg [7:0] p8_array_index_2045249;
  reg [7:0] p8_array_index_2045250;
  reg [7:0] p8_array_index_2045252;
  reg [7:0] p8_res7__96;
  reg [7:0] p8_array_index_2045261;
  reg [7:0] p8_array_index_2045262;
  reg [7:0] p8_array_index_2045263;
  reg [7:0] p8_array_index_2045264;
  reg [7:0] p8_array_index_2045265;
  reg [7:0] p8_array_index_2045266;
  reg [7:0] p8_res7__98;
  reg [7:0] p8_array_index_2045276;
  reg [7:0] p8_array_index_2045277;
  reg [7:0] p8_array_index_2045278;
  reg [7:0] p8_array_index_2045279;
  reg [7:0] p8_array_index_2045280;
  reg [7:0] p8_res7__100;
  reg [7:0] p8_array_index_2045290;
  reg [7:0] p8_array_index_2045291;
  reg [7:0] p8_array_index_2045292;
  reg [7:0] p8_array_index_2045293;
  reg [7:0] p8_array_index_2045294;
  reg [7:0] p8_res7__102;
  reg [7:0] p9_literal_2043896[256];
  reg [7:0] p9_literal_2043910[256];
  reg [7:0] p9_literal_2043912[256];
  reg [7:0] p9_literal_2043914[256];
  reg [7:0] p9_literal_2043916[256];
  reg [7:0] p9_literal_2043918[256];
  reg [7:0] p9_literal_2043920[256];
  reg [7:0] p9_literal_2043923[256];
  reg [7:0] p86_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p8_encoded <= p7_encoded;
    p8_bit_slice_2043893 <= p7_bit_slice_2043893;
    p8_bit_slice_2044018 <= p7_bit_slice_2044018;
    p8_xor_2044738 <= p7_xor_2044738;
    p8_xor_2045212 <= p8_xor_2045212_comb;
    p8_array_index_2045228 <= p8_array_index_2045228_comb;
    p8_array_index_2045229 <= p8_array_index_2045229_comb;
    p8_array_index_2045230 <= p8_array_index_2045230_comb;
    p8_array_index_2045231 <= p8_array_index_2045231_comb;
    p8_array_index_2045232 <= p8_array_index_2045232_comb;
    p8_array_index_2045233 <= p8_array_index_2045233_comb;
    p8_array_index_2045235 <= p8_array_index_2045235_comb;
    p8_array_index_2045237 <= p8_array_index_2045237_comb;
    p8_array_index_2045238 <= p8_array_index_2045238_comb;
    p8_array_index_2045239 <= p8_array_index_2045239_comb;
    p8_array_index_2045244 <= p8_array_index_2045244_comb;
    p8_array_index_2045245 <= p8_array_index_2045245_comb;
    p8_array_index_2045246 <= p8_array_index_2045246_comb;
    p8_array_index_2045247 <= p8_array_index_2045247_comb;
    p8_array_index_2045248 <= p8_array_index_2045248_comb;
    p8_array_index_2045249 <= p8_array_index_2045249_comb;
    p8_array_index_2045250 <= p8_array_index_2045250_comb;
    p8_array_index_2045252 <= p8_array_index_2045252_comb;
    p8_res7__96 <= p8_res7__96_comb;
    p8_array_index_2045261 <= p8_array_index_2045261_comb;
    p8_array_index_2045262 <= p8_array_index_2045262_comb;
    p8_array_index_2045263 <= p8_array_index_2045263_comb;
    p8_array_index_2045264 <= p8_array_index_2045264_comb;
    p8_array_index_2045265 <= p8_array_index_2045265_comb;
    p8_array_index_2045266 <= p8_array_index_2045266_comb;
    p8_res7__98 <= p8_res7__98_comb;
    p8_array_index_2045276 <= p8_array_index_2045276_comb;
    p8_array_index_2045277 <= p8_array_index_2045277_comb;
    p8_array_index_2045278 <= p8_array_index_2045278_comb;
    p8_array_index_2045279 <= p8_array_index_2045279_comb;
    p8_array_index_2045280 <= p8_array_index_2045280_comb;
    p8_res7__100 <= p8_res7__100_comb;
    p8_array_index_2045290 <= p8_array_index_2045290_comb;
    p8_array_index_2045291 <= p8_array_index_2045291_comb;
    p8_array_index_2045292 <= p8_array_index_2045292_comb;
    p8_array_index_2045293 <= p8_array_index_2045293_comb;
    p8_array_index_2045294 <= p8_array_index_2045294_comb;
    p8_res7__102 <= p8_res7__102_comb;
    p9_literal_2043896 <= p8_literal_2043896;
    p9_literal_2043910 <= p8_literal_2043910;
    p9_literal_2043912 <= p8_literal_2043912;
    p9_literal_2043914 <= p8_literal_2043914;
    p9_literal_2043916 <= p8_literal_2043916;
    p9_literal_2043918 <= p8_literal_2043918;
    p9_literal_2043920 <= p8_literal_2043920;
    p9_literal_2043923 <= p8_literal_2043923;
    p86_literal_2058836 <= p85_literal_2058836;
  end

  // ===== Pipe stage 9:
  wire [7:0] p9_array_index_2045407_comb;
  wire [7:0] p9_array_index_2045408_comb;
  wire [7:0] p9_array_index_2045409_comb;
  wire [7:0] p9_array_index_2045410_comb;
  wire [7:0] p9_res7__104_comb;
  wire [7:0] p9_array_index_2045420_comb;
  wire [7:0] p9_array_index_2045421_comb;
  wire [7:0] p9_array_index_2045422_comb;
  wire [7:0] p9_array_index_2045423_comb;
  wire [7:0] p9_res7__106_comb;
  wire [7:0] p9_array_index_2045434_comb;
  wire [7:0] p9_array_index_2045435_comb;
  wire [7:0] p9_array_index_2045436_comb;
  wire [7:0] p9_res7__108_comb;
  wire [7:0] p9_array_index_2045446_comb;
  wire [7:0] p9_array_index_2045447_comb;
  wire [7:0] p9_array_index_2045448_comb;
  wire [7:0] p9_res7__110_comb;
  wire [7:0] p9_array_index_2045459_comb;
  wire [7:0] p9_array_index_2045460_comb;
  wire [7:0] p9_res7__112_comb;
  wire [7:0] p9_array_index_2045470_comb;
  wire [7:0] p9_array_index_2045471_comb;
  wire [7:0] p9_res7__114_comb;
  wire [7:0] p9_array_index_2045482_comb;
  wire [7:0] p9_res7__116_comb;
  assign p9_array_index_2045407_comb = p8_literal_2043914[p8_res7__98];
  assign p9_array_index_2045408_comb = p8_literal_2043916[p8_res7__96];
  assign p9_array_index_2045409_comb = p8_literal_2043918[p8_array_index_2045228];
  assign p9_array_index_2045410_comb = p8_literal_2043920[p8_array_index_2045229];
  assign p9_res7__104_comb = p8_literal_2043910[p8_res7__102] ^ p8_literal_2043912[p8_res7__100] ^ p9_array_index_2045407_comb ^ p9_array_index_2045408_comb ^ p9_array_index_2045409_comb ^ p9_array_index_2045410_comb ^ p8_array_index_2045230 ^ p8_literal_2043923[p8_array_index_2045231] ^ p8_array_index_2045232 ^ p8_array_index_2045249 ^ p8_literal_2043918[p8_array_index_2045250] ^ p8_literal_2043916[p8_array_index_2045235] ^ p8_literal_2043914[p8_array_index_2045252] ^ p8_literal_2043912[p8_array_index_2045237] ^ p8_literal_2043910[p8_array_index_2045238] ^ p8_array_index_2045239;
  assign p9_array_index_2045420_comb = p8_literal_2043914[p8_res7__100];
  assign p9_array_index_2045421_comb = p8_literal_2043916[p8_res7__98];
  assign p9_array_index_2045422_comb = p8_literal_2043918[p8_res7__96];
  assign p9_array_index_2045423_comb = p8_literal_2043920[p8_array_index_2045228];
  assign p9_res7__106_comb = p8_literal_2043910[p9_res7__104_comb] ^ p8_literal_2043912[p8_res7__102] ^ p9_array_index_2045420_comb ^ p9_array_index_2045421_comb ^ p9_array_index_2045422_comb ^ p9_array_index_2045423_comb ^ p8_array_index_2045229 ^ p8_literal_2043923[p8_array_index_2045230] ^ p8_array_index_2045231 ^ p8_array_index_2045266 ^ p8_literal_2043918[p8_array_index_2045233] ^ p8_literal_2043916[p8_array_index_2045250] ^ p8_literal_2043914[p8_array_index_2045235] ^ p8_literal_2043912[p8_array_index_2045252] ^ p8_literal_2043910[p8_array_index_2045237] ^ p8_array_index_2045238;
  assign p9_array_index_2045434_comb = p8_literal_2043916[p8_res7__100];
  assign p9_array_index_2045435_comb = p8_literal_2043918[p8_res7__98];
  assign p9_array_index_2045436_comb = p8_literal_2043920[p8_res7__96];
  assign p9_res7__108_comb = p8_literal_2043910[p9_res7__106_comb] ^ p8_literal_2043912[p9_res7__104_comb] ^ p8_literal_2043914[p8_res7__102] ^ p9_array_index_2045434_comb ^ p9_array_index_2045435_comb ^ p9_array_index_2045436_comb ^ p8_array_index_2045228 ^ p8_literal_2043923[p8_array_index_2045229] ^ p8_array_index_2045230 ^ p8_array_index_2045280 ^ p8_array_index_2045248 ^ p8_literal_2043916[p8_array_index_2045233] ^ p8_literal_2043914[p8_array_index_2045250] ^ p8_literal_2043912[p8_array_index_2045235] ^ p8_literal_2043910[p8_array_index_2045252] ^ p8_array_index_2045237;
  assign p9_array_index_2045446_comb = p8_literal_2043916[p8_res7__102];
  assign p9_array_index_2045447_comb = p8_literal_2043918[p8_res7__100];
  assign p9_array_index_2045448_comb = p8_literal_2043920[p8_res7__98];
  assign p9_res7__110_comb = p8_literal_2043910[p9_res7__108_comb] ^ p8_literal_2043912[p9_res7__106_comb] ^ p8_literal_2043914[p9_res7__104_comb] ^ p9_array_index_2045446_comb ^ p9_array_index_2045447_comb ^ p9_array_index_2045448_comb ^ p8_res7__96 ^ p8_literal_2043923[p8_array_index_2045228] ^ p8_array_index_2045229 ^ p8_array_index_2045294 ^ p8_array_index_2045265 ^ p8_literal_2043916[p8_array_index_2045232] ^ p8_literal_2043914[p8_array_index_2045233] ^ p8_literal_2043912[p8_array_index_2045250] ^ p8_literal_2043910[p8_array_index_2045235] ^ p8_array_index_2045252;
  assign p9_array_index_2045459_comb = p8_literal_2043918[p8_res7__102];
  assign p9_array_index_2045460_comb = p8_literal_2043920[p8_res7__100];
  assign p9_res7__112_comb = p8_literal_2043910[p9_res7__110_comb] ^ p8_literal_2043912[p9_res7__108_comb] ^ p8_literal_2043914[p9_res7__106_comb] ^ p8_literal_2043916[p9_res7__104_comb] ^ p9_array_index_2045459_comb ^ p9_array_index_2045460_comb ^ p8_res7__98 ^ p8_literal_2043923[p8_res7__96] ^ p8_array_index_2045228 ^ p9_array_index_2045410_comb ^ p8_array_index_2045279 ^ p8_array_index_2045247 ^ p8_literal_2043914[p8_array_index_2045232] ^ p8_literal_2043912[p8_array_index_2045233] ^ p8_literal_2043910[p8_array_index_2045250] ^ p8_array_index_2045235;
  assign p9_array_index_2045470_comb = p8_literal_2043918[p9_res7__104_comb];
  assign p9_array_index_2045471_comb = p8_literal_2043920[p8_res7__102];
  assign p9_res7__114_comb = p8_literal_2043910[p9_res7__112_comb] ^ p8_literal_2043912[p9_res7__110_comb] ^ p8_literal_2043914[p9_res7__108_comb] ^ p8_literal_2043916[p9_res7__106_comb] ^ p9_array_index_2045470_comb ^ p9_array_index_2045471_comb ^ p8_res7__100 ^ p8_literal_2043923[p8_res7__98] ^ p8_res7__96 ^ p9_array_index_2045423_comb ^ p8_array_index_2045293 ^ p8_array_index_2045264 ^ p8_literal_2043914[p8_array_index_2045231] ^ p8_literal_2043912[p8_array_index_2045232] ^ p8_literal_2043910[p8_array_index_2045233] ^ p8_array_index_2045250;
  assign p9_array_index_2045482_comb = p8_literal_2043920[p9_res7__104_comb];
  assign p9_res7__116_comb = p8_literal_2043910[p9_res7__114_comb] ^ p8_literal_2043912[p9_res7__112_comb] ^ p8_literal_2043914[p9_res7__110_comb] ^ p8_literal_2043916[p9_res7__108_comb] ^ p8_literal_2043918[p9_res7__106_comb] ^ p9_array_index_2045482_comb ^ p8_res7__102 ^ p8_literal_2043923[p8_res7__100] ^ p8_res7__98 ^ p9_array_index_2045436_comb ^ p9_array_index_2045409_comb ^ p8_array_index_2045278 ^ p8_array_index_2045246 ^ p8_literal_2043912[p8_array_index_2045231] ^ p8_literal_2043910[p8_array_index_2045232] ^ p8_array_index_2045233;

  // Registers for pipe stage 9:
  reg [127:0] p9_encoded;
  reg [127:0] p9_bit_slice_2043893;
  reg [127:0] p9_bit_slice_2044018;
  reg [127:0] p9_xor_2044738;
  reg [127:0] p9_xor_2045212;
  reg [7:0] p9_array_index_2045228;
  reg [7:0] p9_array_index_2045229;
  reg [7:0] p9_array_index_2045230;
  reg [7:0] p9_array_index_2045231;
  reg [7:0] p9_array_index_2045232;
  reg [7:0] p9_array_index_2045244;
  reg [7:0] p9_array_index_2045245;
  reg [7:0] p9_res7__96;
  reg [7:0] p9_array_index_2045261;
  reg [7:0] p9_array_index_2045262;
  reg [7:0] p9_array_index_2045263;
  reg [7:0] p9_res7__98;
  reg [7:0] p9_array_index_2045276;
  reg [7:0] p9_array_index_2045277;
  reg [7:0] p9_res7__100;
  reg [7:0] p9_array_index_2045290;
  reg [7:0] p9_array_index_2045291;
  reg [7:0] p9_array_index_2045292;
  reg [7:0] p9_res7__102;
  reg [7:0] p9_array_index_2045407;
  reg [7:0] p9_array_index_2045408;
  reg [7:0] p9_res7__104;
  reg [7:0] p9_array_index_2045420;
  reg [7:0] p9_array_index_2045421;
  reg [7:0] p9_array_index_2045422;
  reg [7:0] p9_res7__106;
  reg [7:0] p9_array_index_2045434;
  reg [7:0] p9_array_index_2045435;
  reg [7:0] p9_res7__108;
  reg [7:0] p9_array_index_2045446;
  reg [7:0] p9_array_index_2045447;
  reg [7:0] p9_array_index_2045448;
  reg [7:0] p9_res7__110;
  reg [7:0] p9_array_index_2045459;
  reg [7:0] p9_array_index_2045460;
  reg [7:0] p9_res7__112;
  reg [7:0] p9_array_index_2045470;
  reg [7:0] p9_array_index_2045471;
  reg [7:0] p9_res7__114;
  reg [7:0] p9_array_index_2045482;
  reg [7:0] p9_res7__116;
  reg [7:0] p10_literal_2043896[256];
  reg [7:0] p10_literal_2043910[256];
  reg [7:0] p10_literal_2043912[256];
  reg [7:0] p10_literal_2043914[256];
  reg [7:0] p10_literal_2043916[256];
  reg [7:0] p10_literal_2043918[256];
  reg [7:0] p10_literal_2043920[256];
  reg [7:0] p10_literal_2043923[256];
  reg [7:0] p87_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p9_encoded <= p8_encoded;
    p9_bit_slice_2043893 <= p8_bit_slice_2043893;
    p9_bit_slice_2044018 <= p8_bit_slice_2044018;
    p9_xor_2044738 <= p8_xor_2044738;
    p9_xor_2045212 <= p8_xor_2045212;
    p9_array_index_2045228 <= p8_array_index_2045228;
    p9_array_index_2045229 <= p8_array_index_2045229;
    p9_array_index_2045230 <= p8_array_index_2045230;
    p9_array_index_2045231 <= p8_array_index_2045231;
    p9_array_index_2045232 <= p8_array_index_2045232;
    p9_array_index_2045244 <= p8_array_index_2045244;
    p9_array_index_2045245 <= p8_array_index_2045245;
    p9_res7__96 <= p8_res7__96;
    p9_array_index_2045261 <= p8_array_index_2045261;
    p9_array_index_2045262 <= p8_array_index_2045262;
    p9_array_index_2045263 <= p8_array_index_2045263;
    p9_res7__98 <= p8_res7__98;
    p9_array_index_2045276 <= p8_array_index_2045276;
    p9_array_index_2045277 <= p8_array_index_2045277;
    p9_res7__100 <= p8_res7__100;
    p9_array_index_2045290 <= p8_array_index_2045290;
    p9_array_index_2045291 <= p8_array_index_2045291;
    p9_array_index_2045292 <= p8_array_index_2045292;
    p9_res7__102 <= p8_res7__102;
    p9_array_index_2045407 <= p9_array_index_2045407_comb;
    p9_array_index_2045408 <= p9_array_index_2045408_comb;
    p9_res7__104 <= p9_res7__104_comb;
    p9_array_index_2045420 <= p9_array_index_2045420_comb;
    p9_array_index_2045421 <= p9_array_index_2045421_comb;
    p9_array_index_2045422 <= p9_array_index_2045422_comb;
    p9_res7__106 <= p9_res7__106_comb;
    p9_array_index_2045434 <= p9_array_index_2045434_comb;
    p9_array_index_2045435 <= p9_array_index_2045435_comb;
    p9_res7__108 <= p9_res7__108_comb;
    p9_array_index_2045446 <= p9_array_index_2045446_comb;
    p9_array_index_2045447 <= p9_array_index_2045447_comb;
    p9_array_index_2045448 <= p9_array_index_2045448_comb;
    p9_res7__110 <= p9_res7__110_comb;
    p9_array_index_2045459 <= p9_array_index_2045459_comb;
    p9_array_index_2045460 <= p9_array_index_2045460_comb;
    p9_res7__112 <= p9_res7__112_comb;
    p9_array_index_2045470 <= p9_array_index_2045470_comb;
    p9_array_index_2045471 <= p9_array_index_2045471_comb;
    p9_res7__114 <= p9_res7__114_comb;
    p9_array_index_2045482 <= p9_array_index_2045482_comb;
    p9_res7__116 <= p9_res7__116_comb;
    p10_literal_2043896 <= p9_literal_2043896;
    p10_literal_2043910 <= p9_literal_2043910;
    p10_literal_2043912 <= p9_literal_2043912;
    p10_literal_2043914 <= p9_literal_2043914;
    p10_literal_2043916 <= p9_literal_2043916;
    p10_literal_2043918 <= p9_literal_2043918;
    p10_literal_2043920 <= p9_literal_2043920;
    p10_literal_2043923 <= p9_literal_2043923;
    p87_literal_2058836 <= p86_literal_2058836;
  end

  // ===== Pipe stage 10:
  wire [7:0] p10_array_index_2045600_comb;
  wire [7:0] p10_res7__118_comb;
  wire [7:0] p10_res7__120_comb;
  wire [7:0] p10_res7__122_comb;
  wire [7:0] p10_res7__124_comb;
  wire [7:0] p10_res7__126_comb;
  wire [127:0] p10_res__3_comb;
  wire [127:0] p10_xor_2045640_comb;
  wire [127:0] p10_addedKey__36_comb;
  wire [7:0] p10_array_index_2045656_comb;
  wire [7:0] p10_array_index_2045657_comb;
  wire [7:0] p10_array_index_2045658_comb;
  wire [7:0] p10_array_index_2045659_comb;
  wire [7:0] p10_array_index_2045660_comb;
  wire [7:0] p10_array_index_2045661_comb;
  wire [7:0] p10_array_index_2045663_comb;
  wire [7:0] p10_array_index_2045665_comb;
  wire [7:0] p10_array_index_2045666_comb;
  wire [7:0] p10_array_index_2045667_comb;
  wire [7:0] p10_array_index_2045668_comb;
  wire [7:0] p10_array_index_2045669_comb;
  wire [7:0] p10_array_index_2045670_comb;
  wire [7:0] p10_array_index_2045672_comb;
  wire [7:0] p10_array_index_2045673_comb;
  wire [7:0] p10_array_index_2045674_comb;
  wire [7:0] p10_array_index_2045675_comb;
  wire [7:0] p10_array_index_2045676_comb;
  wire [7:0] p10_array_index_2045677_comb;
  wire [7:0] p10_array_index_2045678_comb;
  wire [7:0] p10_array_index_2045680_comb;
  wire [7:0] p10_res7__128_comb;
  assign p10_array_index_2045600_comb = p9_literal_2043920[p9_res7__106];
  assign p10_res7__118_comb = p9_literal_2043910[p9_res7__116] ^ p9_literal_2043912[p9_res7__114] ^ p9_literal_2043914[p9_res7__112] ^ p9_literal_2043916[p9_res7__110] ^ p9_literal_2043918[p9_res7__108] ^ p10_array_index_2045600_comb ^ p9_res7__104 ^ p9_literal_2043923[p9_res7__102] ^ p9_res7__100 ^ p9_array_index_2045448 ^ p9_array_index_2045422 ^ p9_array_index_2045292 ^ p9_array_index_2045263 ^ p9_literal_2043912[p9_array_index_2045230] ^ p9_literal_2043910[p9_array_index_2045231] ^ p9_array_index_2045232;
  assign p10_res7__120_comb = p9_literal_2043910[p10_res7__118_comb] ^ p9_literal_2043912[p9_res7__116] ^ p9_literal_2043914[p9_res7__114] ^ p9_literal_2043916[p9_res7__112] ^ p9_literal_2043918[p9_res7__110] ^ p9_literal_2043920[p9_res7__108] ^ p9_res7__106 ^ p9_literal_2043923[p9_res7__104] ^ p9_res7__102 ^ p9_array_index_2045460 ^ p9_array_index_2045435 ^ p9_array_index_2045408 ^ p9_array_index_2045277 ^ p9_array_index_2045245 ^ p9_literal_2043910[p9_array_index_2045230] ^ p9_array_index_2045231;
  assign p10_res7__122_comb = p9_literal_2043910[p10_res7__120_comb] ^ p9_literal_2043912[p10_res7__118_comb] ^ p9_literal_2043914[p9_res7__116] ^ p9_literal_2043916[p9_res7__114] ^ p9_literal_2043918[p9_res7__112] ^ p9_literal_2043920[p9_res7__110] ^ p9_res7__108 ^ p9_literal_2043923[p9_res7__106] ^ p9_res7__104 ^ p9_array_index_2045471 ^ p9_array_index_2045447 ^ p9_array_index_2045421 ^ p9_array_index_2045291 ^ p9_array_index_2045262 ^ p9_literal_2043910[p9_array_index_2045229] ^ p9_array_index_2045230;
  assign p10_res7__124_comb = p9_literal_2043910[p10_res7__122_comb] ^ p9_literal_2043912[p10_res7__120_comb] ^ p9_literal_2043914[p10_res7__118_comb] ^ p9_literal_2043916[p9_res7__116] ^ p9_literal_2043918[p9_res7__114] ^ p9_literal_2043920[p9_res7__112] ^ p9_res7__110 ^ p9_literal_2043923[p9_res7__108] ^ p9_res7__106 ^ p9_array_index_2045482 ^ p9_array_index_2045459 ^ p9_array_index_2045434 ^ p9_array_index_2045407 ^ p9_array_index_2045276 ^ p9_array_index_2045244 ^ p9_array_index_2045229;
  assign p10_res7__126_comb = p9_literal_2043910[p10_res7__124_comb] ^ p9_literal_2043912[p10_res7__122_comb] ^ p9_literal_2043914[p10_res7__120_comb] ^ p9_literal_2043916[p10_res7__118_comb] ^ p9_literal_2043918[p9_res7__116] ^ p9_literal_2043920[p9_res7__114] ^ p9_res7__112 ^ p9_literal_2043923[p9_res7__110] ^ p9_res7__108 ^ p10_array_index_2045600_comb ^ p9_array_index_2045470 ^ p9_array_index_2045446 ^ p9_array_index_2045420 ^ p9_array_index_2045290 ^ p9_array_index_2045261 ^ p9_array_index_2045228;
  assign p10_res__3_comb = {p10_res7__126_comb, p10_res7__124_comb, p10_res7__122_comb, p10_res7__120_comb, p10_res7__118_comb, p9_res7__116, p9_res7__114, p9_res7__112, p9_res7__110, p9_res7__108, p9_res7__106, p9_res7__104, p9_res7__102, p9_res7__100, p9_res7__98, p9_res7__96};
  assign p10_xor_2045640_comb = p10_res__3_comb ^ p9_xor_2044738;
  assign p10_addedKey__36_comb = p10_xor_2045640_comb ^ 128'h156f_6d79_1fab_511d_eabb_0c50_2fd1_8105;
  assign p10_array_index_2045656_comb = p9_literal_2043896[p10_addedKey__36_comb[127:120]];
  assign p10_array_index_2045657_comb = p9_literal_2043896[p10_addedKey__36_comb[119:112]];
  assign p10_array_index_2045658_comb = p9_literal_2043896[p10_addedKey__36_comb[111:104]];
  assign p10_array_index_2045659_comb = p9_literal_2043896[p10_addedKey__36_comb[103:96]];
  assign p10_array_index_2045660_comb = p9_literal_2043896[p10_addedKey__36_comb[95:88]];
  assign p10_array_index_2045661_comb = p9_literal_2043896[p10_addedKey__36_comb[87:80]];
  assign p10_array_index_2045663_comb = p9_literal_2043896[p10_addedKey__36_comb[71:64]];
  assign p10_array_index_2045665_comb = p9_literal_2043896[p10_addedKey__36_comb[55:48]];
  assign p10_array_index_2045666_comb = p9_literal_2043896[p10_addedKey__36_comb[47:40]];
  assign p10_array_index_2045667_comb = p9_literal_2043896[p10_addedKey__36_comb[39:32]];
  assign p10_array_index_2045668_comb = p9_literal_2043896[p10_addedKey__36_comb[31:24]];
  assign p10_array_index_2045669_comb = p9_literal_2043896[p10_addedKey__36_comb[23:16]];
  assign p10_array_index_2045670_comb = p9_literal_2043896[p10_addedKey__36_comb[15:8]];
  assign p10_array_index_2045672_comb = p9_literal_2043910[p10_array_index_2045656_comb];
  assign p10_array_index_2045673_comb = p9_literal_2043912[p10_array_index_2045657_comb];
  assign p10_array_index_2045674_comb = p9_literal_2043914[p10_array_index_2045658_comb];
  assign p10_array_index_2045675_comb = p9_literal_2043916[p10_array_index_2045659_comb];
  assign p10_array_index_2045676_comb = p9_literal_2043918[p10_array_index_2045660_comb];
  assign p10_array_index_2045677_comb = p9_literal_2043920[p10_array_index_2045661_comb];
  assign p10_array_index_2045678_comb = p9_literal_2043896[p10_addedKey__36_comb[79:72]];
  assign p10_array_index_2045680_comb = p9_literal_2043896[p10_addedKey__36_comb[63:56]];
  assign p10_res7__128_comb = p10_array_index_2045672_comb ^ p10_array_index_2045673_comb ^ p10_array_index_2045674_comb ^ p10_array_index_2045675_comb ^ p10_array_index_2045676_comb ^ p10_array_index_2045677_comb ^ p10_array_index_2045678_comb ^ p9_literal_2043923[p10_array_index_2045663_comb] ^ p10_array_index_2045680_comb ^ p9_literal_2043920[p10_array_index_2045665_comb] ^ p9_literal_2043918[p10_array_index_2045666_comb] ^ p9_literal_2043916[p10_array_index_2045667_comb] ^ p9_literal_2043914[p10_array_index_2045668_comb] ^ p9_literal_2043912[p10_array_index_2045669_comb] ^ p9_literal_2043910[p10_array_index_2045670_comb] ^ p9_literal_2043896[p10_addedKey__36_comb[7:0]];

  // Registers for pipe stage 10:
  reg [127:0] p10_encoded;
  reg [127:0] p10_bit_slice_2043893;
  reg [127:0] p10_bit_slice_2044018;
  reg [127:0] p10_xor_2045212;
  reg [127:0] p10_xor_2045640;
  reg [7:0] p10_array_index_2045656;
  reg [7:0] p10_array_index_2045657;
  reg [7:0] p10_array_index_2045658;
  reg [7:0] p10_array_index_2045659;
  reg [7:0] p10_array_index_2045660;
  reg [7:0] p10_array_index_2045661;
  reg [7:0] p10_array_index_2045663;
  reg [7:0] p10_array_index_2045665;
  reg [7:0] p10_array_index_2045666;
  reg [7:0] p10_array_index_2045667;
  reg [7:0] p10_array_index_2045668;
  reg [7:0] p10_array_index_2045669;
  reg [7:0] p10_array_index_2045670;
  reg [7:0] p10_array_index_2045672;
  reg [7:0] p10_array_index_2045673;
  reg [7:0] p10_array_index_2045674;
  reg [7:0] p10_array_index_2045675;
  reg [7:0] p10_array_index_2045676;
  reg [7:0] p10_array_index_2045677;
  reg [7:0] p10_array_index_2045678;
  reg [7:0] p10_array_index_2045680;
  reg [7:0] p10_res7__128;
  reg [7:0] p11_literal_2043896[256];
  reg [7:0] p11_literal_2043910[256];
  reg [7:0] p11_literal_2043912[256];
  reg [7:0] p11_literal_2043914[256];
  reg [7:0] p11_literal_2043916[256];
  reg [7:0] p11_literal_2043918[256];
  reg [7:0] p11_literal_2043920[256];
  reg [7:0] p11_literal_2043923[256];
  reg [7:0] p88_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p10_encoded <= p9_encoded;
    p10_bit_slice_2043893 <= p9_bit_slice_2043893;
    p10_bit_slice_2044018 <= p9_bit_slice_2044018;
    p10_xor_2045212 <= p9_xor_2045212;
    p10_xor_2045640 <= p10_xor_2045640_comb;
    p10_array_index_2045656 <= p10_array_index_2045656_comb;
    p10_array_index_2045657 <= p10_array_index_2045657_comb;
    p10_array_index_2045658 <= p10_array_index_2045658_comb;
    p10_array_index_2045659 <= p10_array_index_2045659_comb;
    p10_array_index_2045660 <= p10_array_index_2045660_comb;
    p10_array_index_2045661 <= p10_array_index_2045661_comb;
    p10_array_index_2045663 <= p10_array_index_2045663_comb;
    p10_array_index_2045665 <= p10_array_index_2045665_comb;
    p10_array_index_2045666 <= p10_array_index_2045666_comb;
    p10_array_index_2045667 <= p10_array_index_2045667_comb;
    p10_array_index_2045668 <= p10_array_index_2045668_comb;
    p10_array_index_2045669 <= p10_array_index_2045669_comb;
    p10_array_index_2045670 <= p10_array_index_2045670_comb;
    p10_array_index_2045672 <= p10_array_index_2045672_comb;
    p10_array_index_2045673 <= p10_array_index_2045673_comb;
    p10_array_index_2045674 <= p10_array_index_2045674_comb;
    p10_array_index_2045675 <= p10_array_index_2045675_comb;
    p10_array_index_2045676 <= p10_array_index_2045676_comb;
    p10_array_index_2045677 <= p10_array_index_2045677_comb;
    p10_array_index_2045678 <= p10_array_index_2045678_comb;
    p10_array_index_2045680 <= p10_array_index_2045680_comb;
    p10_res7__128 <= p10_res7__128_comb;
    p11_literal_2043896 <= p10_literal_2043896;
    p11_literal_2043910 <= p10_literal_2043910;
    p11_literal_2043912 <= p10_literal_2043912;
    p11_literal_2043914 <= p10_literal_2043914;
    p11_literal_2043916 <= p10_literal_2043916;
    p11_literal_2043918 <= p10_literal_2043918;
    p11_literal_2043920 <= p10_literal_2043920;
    p11_literal_2043923 <= p10_literal_2043923;
    p88_literal_2058836 <= p87_literal_2058836;
  end

  // ===== Pipe stage 11:
  wire [7:0] p11_array_index_2045759_comb;
  wire [7:0] p11_array_index_2045760_comb;
  wire [7:0] p11_array_index_2045761_comb;
  wire [7:0] p11_array_index_2045762_comb;
  wire [7:0] p11_array_index_2045763_comb;
  wire [7:0] p11_array_index_2045764_comb;
  wire [7:0] p11_res7__130_comb;
  wire [7:0] p11_array_index_2045774_comb;
  wire [7:0] p11_array_index_2045775_comb;
  wire [7:0] p11_array_index_2045776_comb;
  wire [7:0] p11_array_index_2045777_comb;
  wire [7:0] p11_array_index_2045778_comb;
  wire [7:0] p11_res7__132_comb;
  wire [7:0] p11_array_index_2045788_comb;
  wire [7:0] p11_array_index_2045789_comb;
  wire [7:0] p11_array_index_2045790_comb;
  wire [7:0] p11_array_index_2045791_comb;
  wire [7:0] p11_array_index_2045792_comb;
  wire [7:0] p11_res7__134_comb;
  wire [7:0] p11_array_index_2045803_comb;
  wire [7:0] p11_array_index_2045804_comb;
  wire [7:0] p11_array_index_2045805_comb;
  wire [7:0] p11_array_index_2045806_comb;
  wire [7:0] p11_res7__136_comb;
  wire [7:0] p11_array_index_2045816_comb;
  wire [7:0] p11_array_index_2045817_comb;
  wire [7:0] p11_array_index_2045818_comb;
  wire [7:0] p11_array_index_2045819_comb;
  wire [7:0] p11_res7__138_comb;
  wire [7:0] p11_array_index_2045830_comb;
  wire [7:0] p11_array_index_2045831_comb;
  wire [7:0] p11_array_index_2045832_comb;
  wire [7:0] p11_res7__140_comb;
  wire [7:0] p11_array_index_2045842_comb;
  wire [7:0] p11_array_index_2045843_comb;
  wire [7:0] p11_array_index_2045844_comb;
  wire [7:0] p11_res7__142_comb;
  assign p11_array_index_2045759_comb = p10_literal_2043910[p10_res7__128];
  assign p11_array_index_2045760_comb = p10_literal_2043912[p10_array_index_2045656];
  assign p11_array_index_2045761_comb = p10_literal_2043914[p10_array_index_2045657];
  assign p11_array_index_2045762_comb = p10_literal_2043916[p10_array_index_2045658];
  assign p11_array_index_2045763_comb = p10_literal_2043918[p10_array_index_2045659];
  assign p11_array_index_2045764_comb = p10_literal_2043920[p10_array_index_2045660];
  assign p11_res7__130_comb = p11_array_index_2045759_comb ^ p11_array_index_2045760_comb ^ p11_array_index_2045761_comb ^ p11_array_index_2045762_comb ^ p11_array_index_2045763_comb ^ p11_array_index_2045764_comb ^ p10_array_index_2045661 ^ p10_literal_2043923[p10_array_index_2045678] ^ p10_array_index_2045663 ^ p10_literal_2043920[p10_array_index_2045680] ^ p10_literal_2043918[p10_array_index_2045665] ^ p10_literal_2043916[p10_array_index_2045666] ^ p10_literal_2043914[p10_array_index_2045667] ^ p10_literal_2043912[p10_array_index_2045668] ^ p10_literal_2043910[p10_array_index_2045669] ^ p10_array_index_2045670;
  assign p11_array_index_2045774_comb = p10_literal_2043912[p10_res7__128];
  assign p11_array_index_2045775_comb = p10_literal_2043914[p10_array_index_2045656];
  assign p11_array_index_2045776_comb = p10_literal_2043916[p10_array_index_2045657];
  assign p11_array_index_2045777_comb = p10_literal_2043918[p10_array_index_2045658];
  assign p11_array_index_2045778_comb = p10_literal_2043920[p10_array_index_2045659];
  assign p11_res7__132_comb = p10_literal_2043910[p11_res7__130_comb] ^ p11_array_index_2045774_comb ^ p11_array_index_2045775_comb ^ p11_array_index_2045776_comb ^ p11_array_index_2045777_comb ^ p11_array_index_2045778_comb ^ p10_array_index_2045660 ^ p10_literal_2043923[p10_array_index_2045661] ^ p10_array_index_2045678 ^ p10_literal_2043920[p10_array_index_2045663] ^ p10_literal_2043918[p10_array_index_2045680] ^ p10_literal_2043916[p10_array_index_2045665] ^ p10_literal_2043914[p10_array_index_2045666] ^ p10_literal_2043912[p10_array_index_2045667] ^ p10_literal_2043910[p10_array_index_2045668] ^ p10_array_index_2045669;
  assign p11_array_index_2045788_comb = p10_literal_2043912[p11_res7__130_comb];
  assign p11_array_index_2045789_comb = p10_literal_2043914[p10_res7__128];
  assign p11_array_index_2045790_comb = p10_literal_2043916[p10_array_index_2045656];
  assign p11_array_index_2045791_comb = p10_literal_2043918[p10_array_index_2045657];
  assign p11_array_index_2045792_comb = p10_literal_2043920[p10_array_index_2045658];
  assign p11_res7__134_comb = p10_literal_2043910[p11_res7__132_comb] ^ p11_array_index_2045788_comb ^ p11_array_index_2045789_comb ^ p11_array_index_2045790_comb ^ p11_array_index_2045791_comb ^ p11_array_index_2045792_comb ^ p10_array_index_2045659 ^ p10_literal_2043923[p10_array_index_2045660] ^ p10_array_index_2045661 ^ p10_literal_2043920[p10_array_index_2045678] ^ p10_literal_2043918[p10_array_index_2045663] ^ p10_literal_2043916[p10_array_index_2045680] ^ p10_literal_2043914[p10_array_index_2045665] ^ p10_literal_2043912[p10_array_index_2045666] ^ p10_literal_2043910[p10_array_index_2045667] ^ p10_array_index_2045668;
  assign p11_array_index_2045803_comb = p10_literal_2043914[p11_res7__130_comb];
  assign p11_array_index_2045804_comb = p10_literal_2043916[p10_res7__128];
  assign p11_array_index_2045805_comb = p10_literal_2043918[p10_array_index_2045656];
  assign p11_array_index_2045806_comb = p10_literal_2043920[p10_array_index_2045657];
  assign p11_res7__136_comb = p10_literal_2043910[p11_res7__134_comb] ^ p10_literal_2043912[p11_res7__132_comb] ^ p11_array_index_2045803_comb ^ p11_array_index_2045804_comb ^ p11_array_index_2045805_comb ^ p11_array_index_2045806_comb ^ p10_array_index_2045658 ^ p10_literal_2043923[p10_array_index_2045659] ^ p10_array_index_2045660 ^ p10_array_index_2045677 ^ p10_literal_2043918[p10_array_index_2045678] ^ p10_literal_2043916[p10_array_index_2045663] ^ p10_literal_2043914[p10_array_index_2045680] ^ p10_literal_2043912[p10_array_index_2045665] ^ p10_literal_2043910[p10_array_index_2045666] ^ p10_array_index_2045667;
  assign p11_array_index_2045816_comb = p10_literal_2043914[p11_res7__132_comb];
  assign p11_array_index_2045817_comb = p10_literal_2043916[p11_res7__130_comb];
  assign p11_array_index_2045818_comb = p10_literal_2043918[p10_res7__128];
  assign p11_array_index_2045819_comb = p10_literal_2043920[p10_array_index_2045656];
  assign p11_res7__138_comb = p10_literal_2043910[p11_res7__136_comb] ^ p10_literal_2043912[p11_res7__134_comb] ^ p11_array_index_2045816_comb ^ p11_array_index_2045817_comb ^ p11_array_index_2045818_comb ^ p11_array_index_2045819_comb ^ p10_array_index_2045657 ^ p10_literal_2043923[p10_array_index_2045658] ^ p10_array_index_2045659 ^ p11_array_index_2045764_comb ^ p10_literal_2043918[p10_array_index_2045661] ^ p10_literal_2043916[p10_array_index_2045678] ^ p10_literal_2043914[p10_array_index_2045663] ^ p10_literal_2043912[p10_array_index_2045680] ^ p10_literal_2043910[p10_array_index_2045665] ^ p10_array_index_2045666;
  assign p11_array_index_2045830_comb = p10_literal_2043916[p11_res7__132_comb];
  assign p11_array_index_2045831_comb = p10_literal_2043918[p11_res7__130_comb];
  assign p11_array_index_2045832_comb = p10_literal_2043920[p10_res7__128];
  assign p11_res7__140_comb = p10_literal_2043910[p11_res7__138_comb] ^ p10_literal_2043912[p11_res7__136_comb] ^ p10_literal_2043914[p11_res7__134_comb] ^ p11_array_index_2045830_comb ^ p11_array_index_2045831_comb ^ p11_array_index_2045832_comb ^ p10_array_index_2045656 ^ p10_literal_2043923[p10_array_index_2045657] ^ p10_array_index_2045658 ^ p11_array_index_2045778_comb ^ p10_array_index_2045676 ^ p10_literal_2043916[p10_array_index_2045661] ^ p10_literal_2043914[p10_array_index_2045678] ^ p10_literal_2043912[p10_array_index_2045663] ^ p10_literal_2043910[p10_array_index_2045680] ^ p10_array_index_2045665;
  assign p11_array_index_2045842_comb = p10_literal_2043916[p11_res7__134_comb];
  assign p11_array_index_2045843_comb = p10_literal_2043918[p11_res7__132_comb];
  assign p11_array_index_2045844_comb = p10_literal_2043920[p11_res7__130_comb];
  assign p11_res7__142_comb = p10_literal_2043910[p11_res7__140_comb] ^ p10_literal_2043912[p11_res7__138_comb] ^ p10_literal_2043914[p11_res7__136_comb] ^ p11_array_index_2045842_comb ^ p11_array_index_2045843_comb ^ p11_array_index_2045844_comb ^ p10_res7__128 ^ p10_literal_2043923[p10_array_index_2045656] ^ p10_array_index_2045657 ^ p11_array_index_2045792_comb ^ p11_array_index_2045763_comb ^ p10_literal_2043916[p10_array_index_2045660] ^ p10_literal_2043914[p10_array_index_2045661] ^ p10_literal_2043912[p10_array_index_2045678] ^ p10_literal_2043910[p10_array_index_2045663] ^ p10_array_index_2045680;

  // Registers for pipe stage 11:
  reg [127:0] p11_encoded;
  reg [127:0] p11_bit_slice_2043893;
  reg [127:0] p11_bit_slice_2044018;
  reg [127:0] p11_xor_2045212;
  reg [127:0] p11_xor_2045640;
  reg [7:0] p11_array_index_2045656;
  reg [7:0] p11_array_index_2045657;
  reg [7:0] p11_array_index_2045658;
  reg [7:0] p11_array_index_2045659;
  reg [7:0] p11_array_index_2045660;
  reg [7:0] p11_array_index_2045661;
  reg [7:0] p11_array_index_2045663;
  reg [7:0] p11_array_index_2045672;
  reg [7:0] p11_array_index_2045673;
  reg [7:0] p11_array_index_2045674;
  reg [7:0] p11_array_index_2045675;
  reg [7:0] p11_array_index_2045678;
  reg [7:0] p11_res7__128;
  reg [7:0] p11_array_index_2045759;
  reg [7:0] p11_array_index_2045760;
  reg [7:0] p11_array_index_2045761;
  reg [7:0] p11_array_index_2045762;
  reg [7:0] p11_res7__130;
  reg [7:0] p11_array_index_2045774;
  reg [7:0] p11_array_index_2045775;
  reg [7:0] p11_array_index_2045776;
  reg [7:0] p11_array_index_2045777;
  reg [7:0] p11_res7__132;
  reg [7:0] p11_array_index_2045788;
  reg [7:0] p11_array_index_2045789;
  reg [7:0] p11_array_index_2045790;
  reg [7:0] p11_array_index_2045791;
  reg [7:0] p11_res7__134;
  reg [7:0] p11_array_index_2045803;
  reg [7:0] p11_array_index_2045804;
  reg [7:0] p11_array_index_2045805;
  reg [7:0] p11_array_index_2045806;
  reg [7:0] p11_res7__136;
  reg [7:0] p11_array_index_2045816;
  reg [7:0] p11_array_index_2045817;
  reg [7:0] p11_array_index_2045818;
  reg [7:0] p11_array_index_2045819;
  reg [7:0] p11_res7__138;
  reg [7:0] p11_array_index_2045830;
  reg [7:0] p11_array_index_2045831;
  reg [7:0] p11_array_index_2045832;
  reg [7:0] p11_res7__140;
  reg [7:0] p11_array_index_2045842;
  reg [7:0] p11_array_index_2045843;
  reg [7:0] p11_array_index_2045844;
  reg [7:0] p11_res7__142;
  reg [7:0] p12_literal_2043896[256];
  reg [7:0] p12_literal_2043910[256];
  reg [7:0] p12_literal_2043912[256];
  reg [7:0] p12_literal_2043914[256];
  reg [7:0] p12_literal_2043916[256];
  reg [7:0] p12_literal_2043918[256];
  reg [7:0] p12_literal_2043920[256];
  reg [7:0] p12_literal_2043923[256];
  reg [7:0] p89_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p11_encoded <= p10_encoded;
    p11_bit_slice_2043893 <= p10_bit_slice_2043893;
    p11_bit_slice_2044018 <= p10_bit_slice_2044018;
    p11_xor_2045212 <= p10_xor_2045212;
    p11_xor_2045640 <= p10_xor_2045640;
    p11_array_index_2045656 <= p10_array_index_2045656;
    p11_array_index_2045657 <= p10_array_index_2045657;
    p11_array_index_2045658 <= p10_array_index_2045658;
    p11_array_index_2045659 <= p10_array_index_2045659;
    p11_array_index_2045660 <= p10_array_index_2045660;
    p11_array_index_2045661 <= p10_array_index_2045661;
    p11_array_index_2045663 <= p10_array_index_2045663;
    p11_array_index_2045672 <= p10_array_index_2045672;
    p11_array_index_2045673 <= p10_array_index_2045673;
    p11_array_index_2045674 <= p10_array_index_2045674;
    p11_array_index_2045675 <= p10_array_index_2045675;
    p11_array_index_2045678 <= p10_array_index_2045678;
    p11_res7__128 <= p10_res7__128;
    p11_array_index_2045759 <= p11_array_index_2045759_comb;
    p11_array_index_2045760 <= p11_array_index_2045760_comb;
    p11_array_index_2045761 <= p11_array_index_2045761_comb;
    p11_array_index_2045762 <= p11_array_index_2045762_comb;
    p11_res7__130 <= p11_res7__130_comb;
    p11_array_index_2045774 <= p11_array_index_2045774_comb;
    p11_array_index_2045775 <= p11_array_index_2045775_comb;
    p11_array_index_2045776 <= p11_array_index_2045776_comb;
    p11_array_index_2045777 <= p11_array_index_2045777_comb;
    p11_res7__132 <= p11_res7__132_comb;
    p11_array_index_2045788 <= p11_array_index_2045788_comb;
    p11_array_index_2045789 <= p11_array_index_2045789_comb;
    p11_array_index_2045790 <= p11_array_index_2045790_comb;
    p11_array_index_2045791 <= p11_array_index_2045791_comb;
    p11_res7__134 <= p11_res7__134_comb;
    p11_array_index_2045803 <= p11_array_index_2045803_comb;
    p11_array_index_2045804 <= p11_array_index_2045804_comb;
    p11_array_index_2045805 <= p11_array_index_2045805_comb;
    p11_array_index_2045806 <= p11_array_index_2045806_comb;
    p11_res7__136 <= p11_res7__136_comb;
    p11_array_index_2045816 <= p11_array_index_2045816_comb;
    p11_array_index_2045817 <= p11_array_index_2045817_comb;
    p11_array_index_2045818 <= p11_array_index_2045818_comb;
    p11_array_index_2045819 <= p11_array_index_2045819_comb;
    p11_res7__138 <= p11_res7__138_comb;
    p11_array_index_2045830 <= p11_array_index_2045830_comb;
    p11_array_index_2045831 <= p11_array_index_2045831_comb;
    p11_array_index_2045832 <= p11_array_index_2045832_comb;
    p11_res7__140 <= p11_res7__140_comb;
    p11_array_index_2045842 <= p11_array_index_2045842_comb;
    p11_array_index_2045843 <= p11_array_index_2045843_comb;
    p11_array_index_2045844 <= p11_array_index_2045844_comb;
    p11_res7__142 <= p11_res7__142_comb;
    p12_literal_2043896 <= p11_literal_2043896;
    p12_literal_2043910 <= p11_literal_2043910;
    p12_literal_2043912 <= p11_literal_2043912;
    p12_literal_2043914 <= p11_literal_2043914;
    p12_literal_2043916 <= p11_literal_2043916;
    p12_literal_2043918 <= p11_literal_2043918;
    p12_literal_2043920 <= p11_literal_2043920;
    p12_literal_2043923 <= p11_literal_2043923;
    p89_literal_2058836 <= p88_literal_2058836;
  end

  // ===== Pipe stage 12:
  wire [7:0] p12_array_index_2045973_comb;
  wire [7:0] p12_array_index_2045974_comb;
  wire [7:0] p12_res7__144_comb;
  wire [7:0] p12_array_index_2045984_comb;
  wire [7:0] p12_array_index_2045985_comb;
  wire [7:0] p12_res7__146_comb;
  wire [7:0] p12_array_index_2045996_comb;
  wire [7:0] p12_res7__148_comb;
  wire [7:0] p12_array_index_2046006_comb;
  wire [7:0] p12_res7__150_comb;
  wire [7:0] p12_res7__152_comb;
  wire [7:0] p12_res7__154_comb;
  wire [7:0] p12_res7__156_comb;
  assign p12_array_index_2045973_comb = p11_literal_2043918[p11_res7__134];
  assign p12_array_index_2045974_comb = p11_literal_2043920[p11_res7__132];
  assign p12_res7__144_comb = p11_literal_2043910[p11_res7__142] ^ p11_literal_2043912[p11_res7__140] ^ p11_literal_2043914[p11_res7__138] ^ p11_literal_2043916[p11_res7__136] ^ p12_array_index_2045973_comb ^ p12_array_index_2045974_comb ^ p11_res7__130 ^ p11_literal_2043923[p11_res7__128] ^ p11_array_index_2045656 ^ p11_array_index_2045806 ^ p11_array_index_2045777 ^ p11_array_index_2045675 ^ p11_literal_2043914[p11_array_index_2045660] ^ p11_literal_2043912[p11_array_index_2045661] ^ p11_literal_2043910[p11_array_index_2045678] ^ p11_array_index_2045663;
  assign p12_array_index_2045984_comb = p11_literal_2043918[p11_res7__136];
  assign p12_array_index_2045985_comb = p11_literal_2043920[p11_res7__134];
  assign p12_res7__146_comb = p11_literal_2043910[p12_res7__144_comb] ^ p11_literal_2043912[p11_res7__142] ^ p11_literal_2043914[p11_res7__140] ^ p11_literal_2043916[p11_res7__138] ^ p12_array_index_2045984_comb ^ p12_array_index_2045985_comb ^ p11_res7__132 ^ p11_literal_2043923[p11_res7__130] ^ p11_res7__128 ^ p11_array_index_2045819 ^ p11_array_index_2045791 ^ p11_array_index_2045762 ^ p11_literal_2043914[p11_array_index_2045659] ^ p11_literal_2043912[p11_array_index_2045660] ^ p11_literal_2043910[p11_array_index_2045661] ^ p11_array_index_2045678;
  assign p12_array_index_2045996_comb = p11_literal_2043920[p11_res7__136];
  assign p12_res7__148_comb = p11_literal_2043910[p12_res7__146_comb] ^ p11_literal_2043912[p12_res7__144_comb] ^ p11_literal_2043914[p11_res7__142] ^ p11_literal_2043916[p11_res7__140] ^ p11_literal_2043918[p11_res7__138] ^ p12_array_index_2045996_comb ^ p11_res7__134 ^ p11_literal_2043923[p11_res7__132] ^ p11_res7__130 ^ p11_array_index_2045832 ^ p11_array_index_2045805 ^ p11_array_index_2045776 ^ p11_array_index_2045674 ^ p11_literal_2043912[p11_array_index_2045659] ^ p11_literal_2043910[p11_array_index_2045660] ^ p11_array_index_2045661;
  assign p12_array_index_2046006_comb = p11_literal_2043920[p11_res7__138];
  assign p12_res7__150_comb = p11_literal_2043910[p12_res7__148_comb] ^ p11_literal_2043912[p12_res7__146_comb] ^ p11_literal_2043914[p12_res7__144_comb] ^ p11_literal_2043916[p11_res7__142] ^ p11_literal_2043918[p11_res7__140] ^ p12_array_index_2046006_comb ^ p11_res7__136 ^ p11_literal_2043923[p11_res7__134] ^ p11_res7__132 ^ p11_array_index_2045844 ^ p11_array_index_2045818 ^ p11_array_index_2045790 ^ p11_array_index_2045761 ^ p11_literal_2043912[p11_array_index_2045658] ^ p11_literal_2043910[p11_array_index_2045659] ^ p11_array_index_2045660;
  assign p12_res7__152_comb = p11_literal_2043910[p12_res7__150_comb] ^ p11_literal_2043912[p12_res7__148_comb] ^ p11_literal_2043914[p12_res7__146_comb] ^ p11_literal_2043916[p12_res7__144_comb] ^ p11_literal_2043918[p11_res7__142] ^ p11_literal_2043920[p11_res7__140] ^ p11_res7__138 ^ p11_literal_2043923[p11_res7__136] ^ p11_res7__134 ^ p12_array_index_2045974_comb ^ p11_array_index_2045831 ^ p11_array_index_2045804 ^ p11_array_index_2045775 ^ p11_array_index_2045673 ^ p11_literal_2043910[p11_array_index_2045658] ^ p11_array_index_2045659;
  assign p12_res7__154_comb = p11_literal_2043910[p12_res7__152_comb] ^ p11_literal_2043912[p12_res7__150_comb] ^ p11_literal_2043914[p12_res7__148_comb] ^ p11_literal_2043916[p12_res7__146_comb] ^ p11_literal_2043918[p12_res7__144_comb] ^ p11_literal_2043920[p11_res7__142] ^ p11_res7__140 ^ p11_literal_2043923[p11_res7__138] ^ p11_res7__136 ^ p12_array_index_2045985_comb ^ p11_array_index_2045843 ^ p11_array_index_2045817 ^ p11_array_index_2045789 ^ p11_array_index_2045760 ^ p11_literal_2043910[p11_array_index_2045657] ^ p11_array_index_2045658;
  assign p12_res7__156_comb = p11_literal_2043910[p12_res7__154_comb] ^ p11_literal_2043912[p12_res7__152_comb] ^ p11_literal_2043914[p12_res7__150_comb] ^ p11_literal_2043916[p12_res7__148_comb] ^ p11_literal_2043918[p12_res7__146_comb] ^ p11_literal_2043920[p12_res7__144_comb] ^ p11_res7__142 ^ p11_literal_2043923[p11_res7__140] ^ p11_res7__138 ^ p12_array_index_2045996_comb ^ p12_array_index_2045973_comb ^ p11_array_index_2045830 ^ p11_array_index_2045803 ^ p11_array_index_2045774 ^ p11_array_index_2045672 ^ p11_array_index_2045657;

  // Registers for pipe stage 12:
  reg [127:0] p12_encoded;
  reg [127:0] p12_bit_slice_2043893;
  reg [127:0] p12_bit_slice_2044018;
  reg [127:0] p12_xor_2045212;
  reg [127:0] p12_xor_2045640;
  reg [7:0] p12_array_index_2045656;
  reg [7:0] p12_res7__128;
  reg [7:0] p12_array_index_2045759;
  reg [7:0] p12_res7__130;
  reg [7:0] p12_res7__132;
  reg [7:0] p12_array_index_2045788;
  reg [7:0] p12_res7__134;
  reg [7:0] p12_res7__136;
  reg [7:0] p12_array_index_2045816;
  reg [7:0] p12_res7__138;
  reg [7:0] p12_res7__140;
  reg [7:0] p12_array_index_2045842;
  reg [7:0] p12_res7__142;
  reg [7:0] p12_res7__144;
  reg [7:0] p12_array_index_2045984;
  reg [7:0] p12_res7__146;
  reg [7:0] p12_res7__148;
  reg [7:0] p12_array_index_2046006;
  reg [7:0] p12_res7__150;
  reg [7:0] p12_res7__152;
  reg [7:0] p12_res7__154;
  reg [7:0] p12_res7__156;
  reg [7:0] p13_literal_2043896[256];
  reg [7:0] p13_literal_2043910[256];
  reg [7:0] p13_literal_2043912[256];
  reg [7:0] p13_literal_2043914[256];
  reg [7:0] p13_literal_2043916[256];
  reg [7:0] p13_literal_2043918[256];
  reg [7:0] p13_literal_2043920[256];
  reg [7:0] p13_literal_2043923[256];
  reg [7:0] p90_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p12_encoded <= p11_encoded;
    p12_bit_slice_2043893 <= p11_bit_slice_2043893;
    p12_bit_slice_2044018 <= p11_bit_slice_2044018;
    p12_xor_2045212 <= p11_xor_2045212;
    p12_xor_2045640 <= p11_xor_2045640;
    p12_array_index_2045656 <= p11_array_index_2045656;
    p12_res7__128 <= p11_res7__128;
    p12_array_index_2045759 <= p11_array_index_2045759;
    p12_res7__130 <= p11_res7__130;
    p12_res7__132 <= p11_res7__132;
    p12_array_index_2045788 <= p11_array_index_2045788;
    p12_res7__134 <= p11_res7__134;
    p12_res7__136 <= p11_res7__136;
    p12_array_index_2045816 <= p11_array_index_2045816;
    p12_res7__138 <= p11_res7__138;
    p12_res7__140 <= p11_res7__140;
    p12_array_index_2045842 <= p11_array_index_2045842;
    p12_res7__142 <= p11_res7__142;
    p12_res7__144 <= p12_res7__144_comb;
    p12_array_index_2045984 <= p12_array_index_2045984_comb;
    p12_res7__146 <= p12_res7__146_comb;
    p12_res7__148 <= p12_res7__148_comb;
    p12_array_index_2046006 <= p12_array_index_2046006_comb;
    p12_res7__150 <= p12_res7__150_comb;
    p12_res7__152 <= p12_res7__152_comb;
    p12_res7__154 <= p12_res7__154_comb;
    p12_res7__156 <= p12_res7__156_comb;
    p13_literal_2043896 <= p12_literal_2043896;
    p13_literal_2043910 <= p12_literal_2043910;
    p13_literal_2043912 <= p12_literal_2043912;
    p13_literal_2043914 <= p12_literal_2043914;
    p13_literal_2043916 <= p12_literal_2043916;
    p13_literal_2043918 <= p12_literal_2043918;
    p13_literal_2043920 <= p12_literal_2043920;
    p13_literal_2043923 <= p12_literal_2043923;
    p90_literal_2058836 <= p89_literal_2058836;
  end

  // ===== Pipe stage 13:
  wire [7:0] p13_res7__158_comb;
  wire [127:0] p13_res__4_comb;
  wire [127:0] p13_xor_2046116_comb;
  wire [127:0] p13_addedKey__37_comb;
  wire [7:0] p13_array_index_2046132_comb;
  wire [7:0] p13_array_index_2046133_comb;
  wire [7:0] p13_array_index_2046134_comb;
  wire [7:0] p13_array_index_2046135_comb;
  wire [7:0] p13_array_index_2046136_comb;
  wire [7:0] p13_array_index_2046137_comb;
  wire [7:0] p13_array_index_2046139_comb;
  wire [7:0] p13_array_index_2046141_comb;
  wire [7:0] p13_array_index_2046142_comb;
  wire [7:0] p13_array_index_2046143_comb;
  wire [7:0] p13_array_index_2046144_comb;
  wire [7:0] p13_array_index_2046145_comb;
  wire [7:0] p13_array_index_2046146_comb;
  wire [7:0] p13_array_index_2046148_comb;
  wire [7:0] p13_array_index_2046149_comb;
  wire [7:0] p13_array_index_2046150_comb;
  wire [7:0] p13_array_index_2046151_comb;
  wire [7:0] p13_array_index_2046152_comb;
  wire [7:0] p13_array_index_2046153_comb;
  wire [7:0] p13_array_index_2046154_comb;
  wire [7:0] p13_array_index_2046156_comb;
  wire [7:0] p13_res7__160_comb;
  wire [7:0] p13_array_index_2046165_comb;
  wire [7:0] p13_array_index_2046166_comb;
  wire [7:0] p13_array_index_2046167_comb;
  wire [7:0] p13_array_index_2046168_comb;
  wire [7:0] p13_array_index_2046169_comb;
  wire [7:0] p13_array_index_2046170_comb;
  wire [7:0] p13_res7__162_comb;
  wire [7:0] p13_array_index_2046180_comb;
  wire [7:0] p13_array_index_2046181_comb;
  wire [7:0] p13_array_index_2046182_comb;
  wire [7:0] p13_array_index_2046183_comb;
  wire [7:0] p13_array_index_2046184_comb;
  wire [7:0] p13_res7__164_comb;
  wire [7:0] p13_array_index_2046194_comb;
  wire [7:0] p13_array_index_2046195_comb;
  wire [7:0] p13_array_index_2046196_comb;
  wire [7:0] p13_array_index_2046197_comb;
  wire [7:0] p13_array_index_2046198_comb;
  wire [7:0] p13_res7__166_comb;
  wire [7:0] p13_array_index_2046209_comb;
  wire [7:0] p13_array_index_2046210_comb;
  wire [7:0] p13_array_index_2046211_comb;
  wire [7:0] p13_array_index_2046212_comb;
  wire [7:0] p13_res7__168_comb;
  assign p13_res7__158_comb = p12_literal_2043910[p12_res7__156] ^ p12_literal_2043912[p12_res7__154] ^ p12_literal_2043914[p12_res7__152] ^ p12_literal_2043916[p12_res7__150] ^ p12_literal_2043918[p12_res7__148] ^ p12_literal_2043920[p12_res7__146] ^ p12_res7__144 ^ p12_literal_2043923[p12_res7__142] ^ p12_res7__140 ^ p12_array_index_2046006 ^ p12_array_index_2045984 ^ p12_array_index_2045842 ^ p12_array_index_2045816 ^ p12_array_index_2045788 ^ p12_array_index_2045759 ^ p12_array_index_2045656;
  assign p13_res__4_comb = {p13_res7__158_comb, p12_res7__156, p12_res7__154, p12_res7__152, p12_res7__150, p12_res7__148, p12_res7__146, p12_res7__144, p12_res7__142, p12_res7__140, p12_res7__138, p12_res7__136, p12_res7__134, p12_res7__132, p12_res7__130, p12_res7__128};
  assign p13_xor_2046116_comb = p13_res__4_comb ^ p12_xor_2045212;
  assign p13_addedKey__37_comb = p13_xor_2046116_comb ^ 128'ha74a_f7ef_ab73_df16_0dd2_0860_8b9e_fe06;
  assign p13_array_index_2046132_comb = p12_literal_2043896[p13_addedKey__37_comb[127:120]];
  assign p13_array_index_2046133_comb = p12_literal_2043896[p13_addedKey__37_comb[119:112]];
  assign p13_array_index_2046134_comb = p12_literal_2043896[p13_addedKey__37_comb[111:104]];
  assign p13_array_index_2046135_comb = p12_literal_2043896[p13_addedKey__37_comb[103:96]];
  assign p13_array_index_2046136_comb = p12_literal_2043896[p13_addedKey__37_comb[95:88]];
  assign p13_array_index_2046137_comb = p12_literal_2043896[p13_addedKey__37_comb[87:80]];
  assign p13_array_index_2046139_comb = p12_literal_2043896[p13_addedKey__37_comb[71:64]];
  assign p13_array_index_2046141_comb = p12_literal_2043896[p13_addedKey__37_comb[55:48]];
  assign p13_array_index_2046142_comb = p12_literal_2043896[p13_addedKey__37_comb[47:40]];
  assign p13_array_index_2046143_comb = p12_literal_2043896[p13_addedKey__37_comb[39:32]];
  assign p13_array_index_2046144_comb = p12_literal_2043896[p13_addedKey__37_comb[31:24]];
  assign p13_array_index_2046145_comb = p12_literal_2043896[p13_addedKey__37_comb[23:16]];
  assign p13_array_index_2046146_comb = p12_literal_2043896[p13_addedKey__37_comb[15:8]];
  assign p13_array_index_2046148_comb = p12_literal_2043910[p13_array_index_2046132_comb];
  assign p13_array_index_2046149_comb = p12_literal_2043912[p13_array_index_2046133_comb];
  assign p13_array_index_2046150_comb = p12_literal_2043914[p13_array_index_2046134_comb];
  assign p13_array_index_2046151_comb = p12_literal_2043916[p13_array_index_2046135_comb];
  assign p13_array_index_2046152_comb = p12_literal_2043918[p13_array_index_2046136_comb];
  assign p13_array_index_2046153_comb = p12_literal_2043920[p13_array_index_2046137_comb];
  assign p13_array_index_2046154_comb = p12_literal_2043896[p13_addedKey__37_comb[79:72]];
  assign p13_array_index_2046156_comb = p12_literal_2043896[p13_addedKey__37_comb[63:56]];
  assign p13_res7__160_comb = p13_array_index_2046148_comb ^ p13_array_index_2046149_comb ^ p13_array_index_2046150_comb ^ p13_array_index_2046151_comb ^ p13_array_index_2046152_comb ^ p13_array_index_2046153_comb ^ p13_array_index_2046154_comb ^ p12_literal_2043923[p13_array_index_2046139_comb] ^ p13_array_index_2046156_comb ^ p12_literal_2043920[p13_array_index_2046141_comb] ^ p12_literal_2043918[p13_array_index_2046142_comb] ^ p12_literal_2043916[p13_array_index_2046143_comb] ^ p12_literal_2043914[p13_array_index_2046144_comb] ^ p12_literal_2043912[p13_array_index_2046145_comb] ^ p12_literal_2043910[p13_array_index_2046146_comb] ^ p12_literal_2043896[p13_addedKey__37_comb[7:0]];
  assign p13_array_index_2046165_comb = p12_literal_2043910[p13_res7__160_comb];
  assign p13_array_index_2046166_comb = p12_literal_2043912[p13_array_index_2046132_comb];
  assign p13_array_index_2046167_comb = p12_literal_2043914[p13_array_index_2046133_comb];
  assign p13_array_index_2046168_comb = p12_literal_2043916[p13_array_index_2046134_comb];
  assign p13_array_index_2046169_comb = p12_literal_2043918[p13_array_index_2046135_comb];
  assign p13_array_index_2046170_comb = p12_literal_2043920[p13_array_index_2046136_comb];
  assign p13_res7__162_comb = p13_array_index_2046165_comb ^ p13_array_index_2046166_comb ^ p13_array_index_2046167_comb ^ p13_array_index_2046168_comb ^ p13_array_index_2046169_comb ^ p13_array_index_2046170_comb ^ p13_array_index_2046137_comb ^ p12_literal_2043923[p13_array_index_2046154_comb] ^ p13_array_index_2046139_comb ^ p12_literal_2043920[p13_array_index_2046156_comb] ^ p12_literal_2043918[p13_array_index_2046141_comb] ^ p12_literal_2043916[p13_array_index_2046142_comb] ^ p12_literal_2043914[p13_array_index_2046143_comb] ^ p12_literal_2043912[p13_array_index_2046144_comb] ^ p12_literal_2043910[p13_array_index_2046145_comb] ^ p13_array_index_2046146_comb;
  assign p13_array_index_2046180_comb = p12_literal_2043912[p13_res7__160_comb];
  assign p13_array_index_2046181_comb = p12_literal_2043914[p13_array_index_2046132_comb];
  assign p13_array_index_2046182_comb = p12_literal_2043916[p13_array_index_2046133_comb];
  assign p13_array_index_2046183_comb = p12_literal_2043918[p13_array_index_2046134_comb];
  assign p13_array_index_2046184_comb = p12_literal_2043920[p13_array_index_2046135_comb];
  assign p13_res7__164_comb = p12_literal_2043910[p13_res7__162_comb] ^ p13_array_index_2046180_comb ^ p13_array_index_2046181_comb ^ p13_array_index_2046182_comb ^ p13_array_index_2046183_comb ^ p13_array_index_2046184_comb ^ p13_array_index_2046136_comb ^ p12_literal_2043923[p13_array_index_2046137_comb] ^ p13_array_index_2046154_comb ^ p12_literal_2043920[p13_array_index_2046139_comb] ^ p12_literal_2043918[p13_array_index_2046156_comb] ^ p12_literal_2043916[p13_array_index_2046141_comb] ^ p12_literal_2043914[p13_array_index_2046142_comb] ^ p12_literal_2043912[p13_array_index_2046143_comb] ^ p12_literal_2043910[p13_array_index_2046144_comb] ^ p13_array_index_2046145_comb;
  assign p13_array_index_2046194_comb = p12_literal_2043912[p13_res7__162_comb];
  assign p13_array_index_2046195_comb = p12_literal_2043914[p13_res7__160_comb];
  assign p13_array_index_2046196_comb = p12_literal_2043916[p13_array_index_2046132_comb];
  assign p13_array_index_2046197_comb = p12_literal_2043918[p13_array_index_2046133_comb];
  assign p13_array_index_2046198_comb = p12_literal_2043920[p13_array_index_2046134_comb];
  assign p13_res7__166_comb = p12_literal_2043910[p13_res7__164_comb] ^ p13_array_index_2046194_comb ^ p13_array_index_2046195_comb ^ p13_array_index_2046196_comb ^ p13_array_index_2046197_comb ^ p13_array_index_2046198_comb ^ p13_array_index_2046135_comb ^ p12_literal_2043923[p13_array_index_2046136_comb] ^ p13_array_index_2046137_comb ^ p12_literal_2043920[p13_array_index_2046154_comb] ^ p12_literal_2043918[p13_array_index_2046139_comb] ^ p12_literal_2043916[p13_array_index_2046156_comb] ^ p12_literal_2043914[p13_array_index_2046141_comb] ^ p12_literal_2043912[p13_array_index_2046142_comb] ^ p12_literal_2043910[p13_array_index_2046143_comb] ^ p13_array_index_2046144_comb;
  assign p13_array_index_2046209_comb = p12_literal_2043914[p13_res7__162_comb];
  assign p13_array_index_2046210_comb = p12_literal_2043916[p13_res7__160_comb];
  assign p13_array_index_2046211_comb = p12_literal_2043918[p13_array_index_2046132_comb];
  assign p13_array_index_2046212_comb = p12_literal_2043920[p13_array_index_2046133_comb];
  assign p13_res7__168_comb = p12_literal_2043910[p13_res7__166_comb] ^ p12_literal_2043912[p13_res7__164_comb] ^ p13_array_index_2046209_comb ^ p13_array_index_2046210_comb ^ p13_array_index_2046211_comb ^ p13_array_index_2046212_comb ^ p13_array_index_2046134_comb ^ p12_literal_2043923[p13_array_index_2046135_comb] ^ p13_array_index_2046136_comb ^ p13_array_index_2046153_comb ^ p12_literal_2043918[p13_array_index_2046154_comb] ^ p12_literal_2043916[p13_array_index_2046139_comb] ^ p12_literal_2043914[p13_array_index_2046156_comb] ^ p12_literal_2043912[p13_array_index_2046141_comb] ^ p12_literal_2043910[p13_array_index_2046142_comb] ^ p13_array_index_2046143_comb;

  // Registers for pipe stage 13:
  reg [127:0] p13_encoded;
  reg [127:0] p13_bit_slice_2043893;
  reg [127:0] p13_bit_slice_2044018;
  reg [127:0] p13_xor_2045640;
  reg [127:0] p13_xor_2046116;
  reg [7:0] p13_array_index_2046132;
  reg [7:0] p13_array_index_2046133;
  reg [7:0] p13_array_index_2046134;
  reg [7:0] p13_array_index_2046135;
  reg [7:0] p13_array_index_2046136;
  reg [7:0] p13_array_index_2046137;
  reg [7:0] p13_array_index_2046139;
  reg [7:0] p13_array_index_2046141;
  reg [7:0] p13_array_index_2046142;
  reg [7:0] p13_array_index_2046148;
  reg [7:0] p13_array_index_2046149;
  reg [7:0] p13_array_index_2046150;
  reg [7:0] p13_array_index_2046151;
  reg [7:0] p13_array_index_2046152;
  reg [7:0] p13_array_index_2046154;
  reg [7:0] p13_array_index_2046156;
  reg [7:0] p13_res7__160;
  reg [7:0] p13_array_index_2046165;
  reg [7:0] p13_array_index_2046166;
  reg [7:0] p13_array_index_2046167;
  reg [7:0] p13_array_index_2046168;
  reg [7:0] p13_array_index_2046169;
  reg [7:0] p13_array_index_2046170;
  reg [7:0] p13_res7__162;
  reg [7:0] p13_array_index_2046180;
  reg [7:0] p13_array_index_2046181;
  reg [7:0] p13_array_index_2046182;
  reg [7:0] p13_array_index_2046183;
  reg [7:0] p13_array_index_2046184;
  reg [7:0] p13_res7__164;
  reg [7:0] p13_array_index_2046194;
  reg [7:0] p13_array_index_2046195;
  reg [7:0] p13_array_index_2046196;
  reg [7:0] p13_array_index_2046197;
  reg [7:0] p13_array_index_2046198;
  reg [7:0] p13_res7__166;
  reg [7:0] p13_array_index_2046209;
  reg [7:0] p13_array_index_2046210;
  reg [7:0] p13_array_index_2046211;
  reg [7:0] p13_array_index_2046212;
  reg [7:0] p13_res7__168;
  reg [7:0] p14_literal_2043896[256];
  reg [7:0] p14_literal_2043910[256];
  reg [7:0] p14_literal_2043912[256];
  reg [7:0] p14_literal_2043914[256];
  reg [7:0] p14_literal_2043916[256];
  reg [7:0] p14_literal_2043918[256];
  reg [7:0] p14_literal_2043920[256];
  reg [7:0] p14_literal_2043923[256];
  reg [7:0] p91_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p13_encoded <= p12_encoded;
    p13_bit_slice_2043893 <= p12_bit_slice_2043893;
    p13_bit_slice_2044018 <= p12_bit_slice_2044018;
    p13_xor_2045640 <= p12_xor_2045640;
    p13_xor_2046116 <= p13_xor_2046116_comb;
    p13_array_index_2046132 <= p13_array_index_2046132_comb;
    p13_array_index_2046133 <= p13_array_index_2046133_comb;
    p13_array_index_2046134 <= p13_array_index_2046134_comb;
    p13_array_index_2046135 <= p13_array_index_2046135_comb;
    p13_array_index_2046136 <= p13_array_index_2046136_comb;
    p13_array_index_2046137 <= p13_array_index_2046137_comb;
    p13_array_index_2046139 <= p13_array_index_2046139_comb;
    p13_array_index_2046141 <= p13_array_index_2046141_comb;
    p13_array_index_2046142 <= p13_array_index_2046142_comb;
    p13_array_index_2046148 <= p13_array_index_2046148_comb;
    p13_array_index_2046149 <= p13_array_index_2046149_comb;
    p13_array_index_2046150 <= p13_array_index_2046150_comb;
    p13_array_index_2046151 <= p13_array_index_2046151_comb;
    p13_array_index_2046152 <= p13_array_index_2046152_comb;
    p13_array_index_2046154 <= p13_array_index_2046154_comb;
    p13_array_index_2046156 <= p13_array_index_2046156_comb;
    p13_res7__160 <= p13_res7__160_comb;
    p13_array_index_2046165 <= p13_array_index_2046165_comb;
    p13_array_index_2046166 <= p13_array_index_2046166_comb;
    p13_array_index_2046167 <= p13_array_index_2046167_comb;
    p13_array_index_2046168 <= p13_array_index_2046168_comb;
    p13_array_index_2046169 <= p13_array_index_2046169_comb;
    p13_array_index_2046170 <= p13_array_index_2046170_comb;
    p13_res7__162 <= p13_res7__162_comb;
    p13_array_index_2046180 <= p13_array_index_2046180_comb;
    p13_array_index_2046181 <= p13_array_index_2046181_comb;
    p13_array_index_2046182 <= p13_array_index_2046182_comb;
    p13_array_index_2046183 <= p13_array_index_2046183_comb;
    p13_array_index_2046184 <= p13_array_index_2046184_comb;
    p13_res7__164 <= p13_res7__164_comb;
    p13_array_index_2046194 <= p13_array_index_2046194_comb;
    p13_array_index_2046195 <= p13_array_index_2046195_comb;
    p13_array_index_2046196 <= p13_array_index_2046196_comb;
    p13_array_index_2046197 <= p13_array_index_2046197_comb;
    p13_array_index_2046198 <= p13_array_index_2046198_comb;
    p13_res7__166 <= p13_res7__166_comb;
    p13_array_index_2046209 <= p13_array_index_2046209_comb;
    p13_array_index_2046210 <= p13_array_index_2046210_comb;
    p13_array_index_2046211 <= p13_array_index_2046211_comb;
    p13_array_index_2046212 <= p13_array_index_2046212_comb;
    p13_res7__168 <= p13_res7__168_comb;
    p14_literal_2043896 <= p13_literal_2043896;
    p14_literal_2043910 <= p13_literal_2043910;
    p14_literal_2043912 <= p13_literal_2043912;
    p14_literal_2043914 <= p13_literal_2043914;
    p14_literal_2043916 <= p13_literal_2043916;
    p14_literal_2043918 <= p13_literal_2043918;
    p14_literal_2043920 <= p13_literal_2043920;
    p14_literal_2043923 <= p13_literal_2043923;
    p91_literal_2058836 <= p90_literal_2058836;
  end

  // ===== Pipe stage 14:
  wire [7:0] p14_array_index_2046330_comb;
  wire [7:0] p14_array_index_2046331_comb;
  wire [7:0] p14_array_index_2046332_comb;
  wire [7:0] p14_array_index_2046333_comb;
  wire [7:0] p14_res7__170_comb;
  wire [7:0] p14_array_index_2046344_comb;
  wire [7:0] p14_array_index_2046345_comb;
  wire [7:0] p14_array_index_2046346_comb;
  wire [7:0] p14_res7__172_comb;
  wire [7:0] p14_array_index_2046356_comb;
  wire [7:0] p14_array_index_2046357_comb;
  wire [7:0] p14_array_index_2046358_comb;
  wire [7:0] p14_res7__174_comb;
  wire [7:0] p14_array_index_2046369_comb;
  wire [7:0] p14_array_index_2046370_comb;
  wire [7:0] p14_res7__176_comb;
  wire [7:0] p14_array_index_2046380_comb;
  wire [7:0] p14_array_index_2046381_comb;
  wire [7:0] p14_res7__178_comb;
  wire [7:0] p14_array_index_2046392_comb;
  wire [7:0] p14_res7__180_comb;
  wire [7:0] p14_array_index_2046402_comb;
  wire [7:0] p14_res7__182_comb;
  assign p14_array_index_2046330_comb = p13_literal_2043914[p13_res7__164];
  assign p14_array_index_2046331_comb = p13_literal_2043916[p13_res7__162];
  assign p14_array_index_2046332_comb = p13_literal_2043918[p13_res7__160];
  assign p14_array_index_2046333_comb = p13_literal_2043920[p13_array_index_2046132];
  assign p14_res7__170_comb = p13_literal_2043910[p13_res7__168] ^ p13_literal_2043912[p13_res7__166] ^ p14_array_index_2046330_comb ^ p14_array_index_2046331_comb ^ p14_array_index_2046332_comb ^ p14_array_index_2046333_comb ^ p13_array_index_2046133 ^ p13_literal_2043923[p13_array_index_2046134] ^ p13_array_index_2046135 ^ p13_array_index_2046170 ^ p13_literal_2043918[p13_array_index_2046137] ^ p13_literal_2043916[p13_array_index_2046154] ^ p13_literal_2043914[p13_array_index_2046139] ^ p13_literal_2043912[p13_array_index_2046156] ^ p13_literal_2043910[p13_array_index_2046141] ^ p13_array_index_2046142;
  assign p14_array_index_2046344_comb = p13_literal_2043916[p13_res7__164];
  assign p14_array_index_2046345_comb = p13_literal_2043918[p13_res7__162];
  assign p14_array_index_2046346_comb = p13_literal_2043920[p13_res7__160];
  assign p14_res7__172_comb = p13_literal_2043910[p14_res7__170_comb] ^ p13_literal_2043912[p13_res7__168] ^ p13_literal_2043914[p13_res7__166] ^ p14_array_index_2046344_comb ^ p14_array_index_2046345_comb ^ p14_array_index_2046346_comb ^ p13_array_index_2046132 ^ p13_literal_2043923[p13_array_index_2046133] ^ p13_array_index_2046134 ^ p13_array_index_2046184 ^ p13_array_index_2046152 ^ p13_literal_2043916[p13_array_index_2046137] ^ p13_literal_2043914[p13_array_index_2046154] ^ p13_literal_2043912[p13_array_index_2046139] ^ p13_literal_2043910[p13_array_index_2046156] ^ p13_array_index_2046141;
  assign p14_array_index_2046356_comb = p13_literal_2043916[p13_res7__166];
  assign p14_array_index_2046357_comb = p13_literal_2043918[p13_res7__164];
  assign p14_array_index_2046358_comb = p13_literal_2043920[p13_res7__162];
  assign p14_res7__174_comb = p13_literal_2043910[p14_res7__172_comb] ^ p13_literal_2043912[p14_res7__170_comb] ^ p13_literal_2043914[p13_res7__168] ^ p14_array_index_2046356_comb ^ p14_array_index_2046357_comb ^ p14_array_index_2046358_comb ^ p13_res7__160 ^ p13_literal_2043923[p13_array_index_2046132] ^ p13_array_index_2046133 ^ p13_array_index_2046198 ^ p13_array_index_2046169 ^ p13_literal_2043916[p13_array_index_2046136] ^ p13_literal_2043914[p13_array_index_2046137] ^ p13_literal_2043912[p13_array_index_2046154] ^ p13_literal_2043910[p13_array_index_2046139] ^ p13_array_index_2046156;
  assign p14_array_index_2046369_comb = p13_literal_2043918[p13_res7__166];
  assign p14_array_index_2046370_comb = p13_literal_2043920[p13_res7__164];
  assign p14_res7__176_comb = p13_literal_2043910[p14_res7__174_comb] ^ p13_literal_2043912[p14_res7__172_comb] ^ p13_literal_2043914[p14_res7__170_comb] ^ p13_literal_2043916[p13_res7__168] ^ p14_array_index_2046369_comb ^ p14_array_index_2046370_comb ^ p13_res7__162 ^ p13_literal_2043923[p13_res7__160] ^ p13_array_index_2046132 ^ p13_array_index_2046212 ^ p13_array_index_2046183 ^ p13_array_index_2046151 ^ p13_literal_2043914[p13_array_index_2046136] ^ p13_literal_2043912[p13_array_index_2046137] ^ p13_literal_2043910[p13_array_index_2046154] ^ p13_array_index_2046139;
  assign p14_array_index_2046380_comb = p13_literal_2043918[p13_res7__168];
  assign p14_array_index_2046381_comb = p13_literal_2043920[p13_res7__166];
  assign p14_res7__178_comb = p13_literal_2043910[p14_res7__176_comb] ^ p13_literal_2043912[p14_res7__174_comb] ^ p13_literal_2043914[p14_res7__172_comb] ^ p13_literal_2043916[p14_res7__170_comb] ^ p14_array_index_2046380_comb ^ p14_array_index_2046381_comb ^ p13_res7__164 ^ p13_literal_2043923[p13_res7__162] ^ p13_res7__160 ^ p14_array_index_2046333_comb ^ p13_array_index_2046197 ^ p13_array_index_2046168 ^ p13_literal_2043914[p13_array_index_2046135] ^ p13_literal_2043912[p13_array_index_2046136] ^ p13_literal_2043910[p13_array_index_2046137] ^ p13_array_index_2046154;
  assign p14_array_index_2046392_comb = p13_literal_2043920[p13_res7__168];
  assign p14_res7__180_comb = p13_literal_2043910[p14_res7__178_comb] ^ p13_literal_2043912[p14_res7__176_comb] ^ p13_literal_2043914[p14_res7__174_comb] ^ p13_literal_2043916[p14_res7__172_comb] ^ p13_literal_2043918[p14_res7__170_comb] ^ p14_array_index_2046392_comb ^ p13_res7__166 ^ p13_literal_2043923[p13_res7__164] ^ p13_res7__162 ^ p14_array_index_2046346_comb ^ p13_array_index_2046211 ^ p13_array_index_2046182 ^ p13_array_index_2046150 ^ p13_literal_2043912[p13_array_index_2046135] ^ p13_literal_2043910[p13_array_index_2046136] ^ p13_array_index_2046137;
  assign p14_array_index_2046402_comb = p13_literal_2043920[p14_res7__170_comb];
  assign p14_res7__182_comb = p13_literal_2043910[p14_res7__180_comb] ^ p13_literal_2043912[p14_res7__178_comb] ^ p13_literal_2043914[p14_res7__176_comb] ^ p13_literal_2043916[p14_res7__174_comb] ^ p13_literal_2043918[p14_res7__172_comb] ^ p14_array_index_2046402_comb ^ p13_res7__168 ^ p13_literal_2043923[p13_res7__166] ^ p13_res7__164 ^ p14_array_index_2046358_comb ^ p14_array_index_2046332_comb ^ p13_array_index_2046196 ^ p13_array_index_2046167 ^ p13_literal_2043912[p13_array_index_2046134] ^ p13_literal_2043910[p13_array_index_2046135] ^ p13_array_index_2046136;

  // Registers for pipe stage 14:
  reg [127:0] p14_encoded;
  reg [127:0] p14_bit_slice_2043893;
  reg [127:0] p14_bit_slice_2044018;
  reg [127:0] p14_xor_2045640;
  reg [127:0] p14_xor_2046116;
  reg [7:0] p14_array_index_2046132;
  reg [7:0] p14_array_index_2046133;
  reg [7:0] p14_array_index_2046134;
  reg [7:0] p14_array_index_2046135;
  reg [7:0] p14_array_index_2046148;
  reg [7:0] p14_array_index_2046149;
  reg [7:0] p14_res7__160;
  reg [7:0] p14_array_index_2046165;
  reg [7:0] p14_array_index_2046166;
  reg [7:0] p14_res7__162;
  reg [7:0] p14_array_index_2046180;
  reg [7:0] p14_array_index_2046181;
  reg [7:0] p14_res7__164;
  reg [7:0] p14_array_index_2046194;
  reg [7:0] p14_array_index_2046195;
  reg [7:0] p14_res7__166;
  reg [7:0] p14_array_index_2046209;
  reg [7:0] p14_array_index_2046210;
  reg [7:0] p14_res7__168;
  reg [7:0] p14_array_index_2046330;
  reg [7:0] p14_array_index_2046331;
  reg [7:0] p14_res7__170;
  reg [7:0] p14_array_index_2046344;
  reg [7:0] p14_array_index_2046345;
  reg [7:0] p14_res7__172;
  reg [7:0] p14_array_index_2046356;
  reg [7:0] p14_array_index_2046357;
  reg [7:0] p14_res7__174;
  reg [7:0] p14_array_index_2046369;
  reg [7:0] p14_array_index_2046370;
  reg [7:0] p14_res7__176;
  reg [7:0] p14_array_index_2046380;
  reg [7:0] p14_array_index_2046381;
  reg [7:0] p14_res7__178;
  reg [7:0] p14_array_index_2046392;
  reg [7:0] p14_res7__180;
  reg [7:0] p14_array_index_2046402;
  reg [7:0] p14_res7__182;
  reg [7:0] p15_literal_2043896[256];
  reg [7:0] p15_literal_2043910[256];
  reg [7:0] p15_literal_2043912[256];
  reg [7:0] p15_literal_2043914[256];
  reg [7:0] p15_literal_2043916[256];
  reg [7:0] p15_literal_2043918[256];
  reg [7:0] p15_literal_2043920[256];
  reg [7:0] p15_literal_2043923[256];
  reg [7:0] p92_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p14_encoded <= p13_encoded;
    p14_bit_slice_2043893 <= p13_bit_slice_2043893;
    p14_bit_slice_2044018 <= p13_bit_slice_2044018;
    p14_xor_2045640 <= p13_xor_2045640;
    p14_xor_2046116 <= p13_xor_2046116;
    p14_array_index_2046132 <= p13_array_index_2046132;
    p14_array_index_2046133 <= p13_array_index_2046133;
    p14_array_index_2046134 <= p13_array_index_2046134;
    p14_array_index_2046135 <= p13_array_index_2046135;
    p14_array_index_2046148 <= p13_array_index_2046148;
    p14_array_index_2046149 <= p13_array_index_2046149;
    p14_res7__160 <= p13_res7__160;
    p14_array_index_2046165 <= p13_array_index_2046165;
    p14_array_index_2046166 <= p13_array_index_2046166;
    p14_res7__162 <= p13_res7__162;
    p14_array_index_2046180 <= p13_array_index_2046180;
    p14_array_index_2046181 <= p13_array_index_2046181;
    p14_res7__164 <= p13_res7__164;
    p14_array_index_2046194 <= p13_array_index_2046194;
    p14_array_index_2046195 <= p13_array_index_2046195;
    p14_res7__166 <= p13_res7__166;
    p14_array_index_2046209 <= p13_array_index_2046209;
    p14_array_index_2046210 <= p13_array_index_2046210;
    p14_res7__168 <= p13_res7__168;
    p14_array_index_2046330 <= p14_array_index_2046330_comb;
    p14_array_index_2046331 <= p14_array_index_2046331_comb;
    p14_res7__170 <= p14_res7__170_comb;
    p14_array_index_2046344 <= p14_array_index_2046344_comb;
    p14_array_index_2046345 <= p14_array_index_2046345_comb;
    p14_res7__172 <= p14_res7__172_comb;
    p14_array_index_2046356 <= p14_array_index_2046356_comb;
    p14_array_index_2046357 <= p14_array_index_2046357_comb;
    p14_res7__174 <= p14_res7__174_comb;
    p14_array_index_2046369 <= p14_array_index_2046369_comb;
    p14_array_index_2046370 <= p14_array_index_2046370_comb;
    p14_res7__176 <= p14_res7__176_comb;
    p14_array_index_2046380 <= p14_array_index_2046380_comb;
    p14_array_index_2046381 <= p14_array_index_2046381_comb;
    p14_res7__178 <= p14_res7__178_comb;
    p14_array_index_2046392 <= p14_array_index_2046392_comb;
    p14_res7__180 <= p14_res7__180_comb;
    p14_array_index_2046402 <= p14_array_index_2046402_comb;
    p14_res7__182 <= p14_res7__182_comb;
    p15_literal_2043896 <= p14_literal_2043896;
    p15_literal_2043910 <= p14_literal_2043910;
    p15_literal_2043912 <= p14_literal_2043912;
    p15_literal_2043914 <= p14_literal_2043914;
    p15_literal_2043916 <= p14_literal_2043916;
    p15_literal_2043918 <= p14_literal_2043918;
    p15_literal_2043920 <= p14_literal_2043920;
    p15_literal_2043923 <= p14_literal_2043923;
    p92_literal_2058836 <= p91_literal_2058836;
  end

  // ===== Pipe stage 15:
  wire [7:0] p15_res7__184_comb;
  wire [7:0] p15_res7__186_comb;
  wire [7:0] p15_res7__188_comb;
  wire [7:0] p15_res7__190_comb;
  wire [127:0] p15_res__5_comb;
  wire [127:0] p15_xor_2046544_comb;
  wire [127:0] p15_addedKey__38_comb;
  wire [7:0] p15_array_index_2046560_comb;
  wire [7:0] p15_array_index_2046561_comb;
  wire [7:0] p15_array_index_2046562_comb;
  wire [7:0] p15_array_index_2046563_comb;
  wire [7:0] p15_array_index_2046564_comb;
  wire [7:0] p15_array_index_2046565_comb;
  wire [7:0] p15_array_index_2046567_comb;
  wire [7:0] p15_array_index_2046569_comb;
  wire [7:0] p15_array_index_2046570_comb;
  wire [7:0] p15_array_index_2046571_comb;
  wire [7:0] p15_array_index_2046572_comb;
  wire [7:0] p15_array_index_2046573_comb;
  wire [7:0] p15_array_index_2046574_comb;
  wire [7:0] p15_array_index_2046576_comb;
  wire [7:0] p15_array_index_2046577_comb;
  wire [7:0] p15_array_index_2046578_comb;
  wire [7:0] p15_array_index_2046579_comb;
  wire [7:0] p15_array_index_2046580_comb;
  wire [7:0] p15_array_index_2046581_comb;
  wire [7:0] p15_array_index_2046582_comb;
  wire [7:0] p15_array_index_2046584_comb;
  wire [7:0] p15_res7__192_comb;
  wire [7:0] p15_array_index_2046593_comb;
  wire [7:0] p15_array_index_2046594_comb;
  wire [7:0] p15_array_index_2046595_comb;
  wire [7:0] p15_array_index_2046596_comb;
  wire [7:0] p15_array_index_2046597_comb;
  wire [7:0] p15_array_index_2046598_comb;
  wire [7:0] p15_res7__194_comb;
  assign p15_res7__184_comb = p14_literal_2043910[p14_res7__182] ^ p14_literal_2043912[p14_res7__180] ^ p14_literal_2043914[p14_res7__178] ^ p14_literal_2043916[p14_res7__176] ^ p14_literal_2043918[p14_res7__174] ^ p14_literal_2043920[p14_res7__172] ^ p14_res7__170 ^ p14_literal_2043923[p14_res7__168] ^ p14_res7__166 ^ p14_array_index_2046370 ^ p14_array_index_2046345 ^ p14_array_index_2046210 ^ p14_array_index_2046181 ^ p14_array_index_2046149 ^ p14_literal_2043910[p14_array_index_2046134] ^ p14_array_index_2046135;
  assign p15_res7__186_comb = p14_literal_2043910[p15_res7__184_comb] ^ p14_literal_2043912[p14_res7__182] ^ p14_literal_2043914[p14_res7__180] ^ p14_literal_2043916[p14_res7__178] ^ p14_literal_2043918[p14_res7__176] ^ p14_literal_2043920[p14_res7__174] ^ p14_res7__172 ^ p14_literal_2043923[p14_res7__170] ^ p14_res7__168 ^ p14_array_index_2046381 ^ p14_array_index_2046357 ^ p14_array_index_2046331 ^ p14_array_index_2046195 ^ p14_array_index_2046166 ^ p14_literal_2043910[p14_array_index_2046133] ^ p14_array_index_2046134;
  assign p15_res7__188_comb = p14_literal_2043910[p15_res7__186_comb] ^ p14_literal_2043912[p15_res7__184_comb] ^ p14_literal_2043914[p14_res7__182] ^ p14_literal_2043916[p14_res7__180] ^ p14_literal_2043918[p14_res7__178] ^ p14_literal_2043920[p14_res7__176] ^ p14_res7__174 ^ p14_literal_2043923[p14_res7__172] ^ p14_res7__170 ^ p14_array_index_2046392 ^ p14_array_index_2046369 ^ p14_array_index_2046344 ^ p14_array_index_2046209 ^ p14_array_index_2046180 ^ p14_array_index_2046148 ^ p14_array_index_2046133;
  assign p15_res7__190_comb = p14_literal_2043910[p15_res7__188_comb] ^ p14_literal_2043912[p15_res7__186_comb] ^ p14_literal_2043914[p15_res7__184_comb] ^ p14_literal_2043916[p14_res7__182] ^ p14_literal_2043918[p14_res7__180] ^ p14_literal_2043920[p14_res7__178] ^ p14_res7__176 ^ p14_literal_2043923[p14_res7__174] ^ p14_res7__172 ^ p14_array_index_2046402 ^ p14_array_index_2046380 ^ p14_array_index_2046356 ^ p14_array_index_2046330 ^ p14_array_index_2046194 ^ p14_array_index_2046165 ^ p14_array_index_2046132;
  assign p15_res__5_comb = {p15_res7__190_comb, p15_res7__188_comb, p15_res7__186_comb, p15_res7__184_comb, p14_res7__182, p14_res7__180, p14_res7__178, p14_res7__176, p14_res7__174, p14_res7__172, p14_res7__170, p14_res7__168, p14_res7__166, p14_res7__164, p14_res7__162, p14_res7__160};
  assign p15_xor_2046544_comb = p15_res__5_comb ^ p14_xor_2045640;
  assign p15_addedKey__38_comb = p15_xor_2046544_comb ^ 128'hc9e8_819d_c73b_a5ae_50f5_b570_561a_6a07;
  assign p15_array_index_2046560_comb = p14_literal_2043896[p15_addedKey__38_comb[127:120]];
  assign p15_array_index_2046561_comb = p14_literal_2043896[p15_addedKey__38_comb[119:112]];
  assign p15_array_index_2046562_comb = p14_literal_2043896[p15_addedKey__38_comb[111:104]];
  assign p15_array_index_2046563_comb = p14_literal_2043896[p15_addedKey__38_comb[103:96]];
  assign p15_array_index_2046564_comb = p14_literal_2043896[p15_addedKey__38_comb[95:88]];
  assign p15_array_index_2046565_comb = p14_literal_2043896[p15_addedKey__38_comb[87:80]];
  assign p15_array_index_2046567_comb = p14_literal_2043896[p15_addedKey__38_comb[71:64]];
  assign p15_array_index_2046569_comb = p14_literal_2043896[p15_addedKey__38_comb[55:48]];
  assign p15_array_index_2046570_comb = p14_literal_2043896[p15_addedKey__38_comb[47:40]];
  assign p15_array_index_2046571_comb = p14_literal_2043896[p15_addedKey__38_comb[39:32]];
  assign p15_array_index_2046572_comb = p14_literal_2043896[p15_addedKey__38_comb[31:24]];
  assign p15_array_index_2046573_comb = p14_literal_2043896[p15_addedKey__38_comb[23:16]];
  assign p15_array_index_2046574_comb = p14_literal_2043896[p15_addedKey__38_comb[15:8]];
  assign p15_array_index_2046576_comb = p14_literal_2043910[p15_array_index_2046560_comb];
  assign p15_array_index_2046577_comb = p14_literal_2043912[p15_array_index_2046561_comb];
  assign p15_array_index_2046578_comb = p14_literal_2043914[p15_array_index_2046562_comb];
  assign p15_array_index_2046579_comb = p14_literal_2043916[p15_array_index_2046563_comb];
  assign p15_array_index_2046580_comb = p14_literal_2043918[p15_array_index_2046564_comb];
  assign p15_array_index_2046581_comb = p14_literal_2043920[p15_array_index_2046565_comb];
  assign p15_array_index_2046582_comb = p14_literal_2043896[p15_addedKey__38_comb[79:72]];
  assign p15_array_index_2046584_comb = p14_literal_2043896[p15_addedKey__38_comb[63:56]];
  assign p15_res7__192_comb = p15_array_index_2046576_comb ^ p15_array_index_2046577_comb ^ p15_array_index_2046578_comb ^ p15_array_index_2046579_comb ^ p15_array_index_2046580_comb ^ p15_array_index_2046581_comb ^ p15_array_index_2046582_comb ^ p14_literal_2043923[p15_array_index_2046567_comb] ^ p15_array_index_2046584_comb ^ p14_literal_2043920[p15_array_index_2046569_comb] ^ p14_literal_2043918[p15_array_index_2046570_comb] ^ p14_literal_2043916[p15_array_index_2046571_comb] ^ p14_literal_2043914[p15_array_index_2046572_comb] ^ p14_literal_2043912[p15_array_index_2046573_comb] ^ p14_literal_2043910[p15_array_index_2046574_comb] ^ p14_literal_2043896[p15_addedKey__38_comb[7:0]];
  assign p15_array_index_2046593_comb = p14_literal_2043910[p15_res7__192_comb];
  assign p15_array_index_2046594_comb = p14_literal_2043912[p15_array_index_2046560_comb];
  assign p15_array_index_2046595_comb = p14_literal_2043914[p15_array_index_2046561_comb];
  assign p15_array_index_2046596_comb = p14_literal_2043916[p15_array_index_2046562_comb];
  assign p15_array_index_2046597_comb = p14_literal_2043918[p15_array_index_2046563_comb];
  assign p15_array_index_2046598_comb = p14_literal_2043920[p15_array_index_2046564_comb];
  assign p15_res7__194_comb = p15_array_index_2046593_comb ^ p15_array_index_2046594_comb ^ p15_array_index_2046595_comb ^ p15_array_index_2046596_comb ^ p15_array_index_2046597_comb ^ p15_array_index_2046598_comb ^ p15_array_index_2046565_comb ^ p14_literal_2043923[p15_array_index_2046582_comb] ^ p15_array_index_2046567_comb ^ p14_literal_2043920[p15_array_index_2046584_comb] ^ p14_literal_2043918[p15_array_index_2046569_comb] ^ p14_literal_2043916[p15_array_index_2046570_comb] ^ p14_literal_2043914[p15_array_index_2046571_comb] ^ p14_literal_2043912[p15_array_index_2046572_comb] ^ p14_literal_2043910[p15_array_index_2046573_comb] ^ p15_array_index_2046574_comb;

  // Registers for pipe stage 15:
  reg [127:0] p15_encoded;
  reg [127:0] p15_bit_slice_2043893;
  reg [127:0] p15_bit_slice_2044018;
  reg [127:0] p15_xor_2046116;
  reg [127:0] p15_xor_2046544;
  reg [7:0] p15_array_index_2046560;
  reg [7:0] p15_array_index_2046561;
  reg [7:0] p15_array_index_2046562;
  reg [7:0] p15_array_index_2046563;
  reg [7:0] p15_array_index_2046564;
  reg [7:0] p15_array_index_2046565;
  reg [7:0] p15_array_index_2046567;
  reg [7:0] p15_array_index_2046569;
  reg [7:0] p15_array_index_2046570;
  reg [7:0] p15_array_index_2046571;
  reg [7:0] p15_array_index_2046572;
  reg [7:0] p15_array_index_2046573;
  reg [7:0] p15_array_index_2046576;
  reg [7:0] p15_array_index_2046577;
  reg [7:0] p15_array_index_2046578;
  reg [7:0] p15_array_index_2046579;
  reg [7:0] p15_array_index_2046580;
  reg [7:0] p15_array_index_2046581;
  reg [7:0] p15_array_index_2046582;
  reg [7:0] p15_array_index_2046584;
  reg [7:0] p15_res7__192;
  reg [7:0] p15_array_index_2046593;
  reg [7:0] p15_array_index_2046594;
  reg [7:0] p15_array_index_2046595;
  reg [7:0] p15_array_index_2046596;
  reg [7:0] p15_array_index_2046597;
  reg [7:0] p15_array_index_2046598;
  reg [7:0] p15_res7__194;
  reg [7:0] p16_literal_2043896[256];
  reg [7:0] p16_literal_2043910[256];
  reg [7:0] p16_literal_2043912[256];
  reg [7:0] p16_literal_2043914[256];
  reg [7:0] p16_literal_2043916[256];
  reg [7:0] p16_literal_2043918[256];
  reg [7:0] p16_literal_2043920[256];
  reg [7:0] p16_literal_2043923[256];
  reg [7:0] p93_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p15_encoded <= p14_encoded;
    p15_bit_slice_2043893 <= p14_bit_slice_2043893;
    p15_bit_slice_2044018 <= p14_bit_slice_2044018;
    p15_xor_2046116 <= p14_xor_2046116;
    p15_xor_2046544 <= p15_xor_2046544_comb;
    p15_array_index_2046560 <= p15_array_index_2046560_comb;
    p15_array_index_2046561 <= p15_array_index_2046561_comb;
    p15_array_index_2046562 <= p15_array_index_2046562_comb;
    p15_array_index_2046563 <= p15_array_index_2046563_comb;
    p15_array_index_2046564 <= p15_array_index_2046564_comb;
    p15_array_index_2046565 <= p15_array_index_2046565_comb;
    p15_array_index_2046567 <= p15_array_index_2046567_comb;
    p15_array_index_2046569 <= p15_array_index_2046569_comb;
    p15_array_index_2046570 <= p15_array_index_2046570_comb;
    p15_array_index_2046571 <= p15_array_index_2046571_comb;
    p15_array_index_2046572 <= p15_array_index_2046572_comb;
    p15_array_index_2046573 <= p15_array_index_2046573_comb;
    p15_array_index_2046576 <= p15_array_index_2046576_comb;
    p15_array_index_2046577 <= p15_array_index_2046577_comb;
    p15_array_index_2046578 <= p15_array_index_2046578_comb;
    p15_array_index_2046579 <= p15_array_index_2046579_comb;
    p15_array_index_2046580 <= p15_array_index_2046580_comb;
    p15_array_index_2046581 <= p15_array_index_2046581_comb;
    p15_array_index_2046582 <= p15_array_index_2046582_comb;
    p15_array_index_2046584 <= p15_array_index_2046584_comb;
    p15_res7__192 <= p15_res7__192_comb;
    p15_array_index_2046593 <= p15_array_index_2046593_comb;
    p15_array_index_2046594 <= p15_array_index_2046594_comb;
    p15_array_index_2046595 <= p15_array_index_2046595_comb;
    p15_array_index_2046596 <= p15_array_index_2046596_comb;
    p15_array_index_2046597 <= p15_array_index_2046597_comb;
    p15_array_index_2046598 <= p15_array_index_2046598_comb;
    p15_res7__194 <= p15_res7__194_comb;
    p16_literal_2043896 <= p15_literal_2043896;
    p16_literal_2043910 <= p15_literal_2043910;
    p16_literal_2043912 <= p15_literal_2043912;
    p16_literal_2043914 <= p15_literal_2043914;
    p16_literal_2043916 <= p15_literal_2043916;
    p16_literal_2043918 <= p15_literal_2043918;
    p16_literal_2043920 <= p15_literal_2043920;
    p16_literal_2043923 <= p15_literal_2043923;
    p93_literal_2058836 <= p92_literal_2058836;
  end

  // ===== Pipe stage 16:
  wire [7:0] p16_array_index_2046690_comb;
  wire [7:0] p16_array_index_2046691_comb;
  wire [7:0] p16_array_index_2046692_comb;
  wire [7:0] p16_array_index_2046693_comb;
  wire [7:0] p16_array_index_2046694_comb;
  wire [7:0] p16_res7__196_comb;
  wire [7:0] p16_array_index_2046704_comb;
  wire [7:0] p16_array_index_2046705_comb;
  wire [7:0] p16_array_index_2046706_comb;
  wire [7:0] p16_array_index_2046707_comb;
  wire [7:0] p16_array_index_2046708_comb;
  wire [7:0] p16_res7__198_comb;
  wire [7:0] p16_array_index_2046719_comb;
  wire [7:0] p16_array_index_2046720_comb;
  wire [7:0] p16_array_index_2046721_comb;
  wire [7:0] p16_array_index_2046722_comb;
  wire [7:0] p16_res7__200_comb;
  wire [7:0] p16_array_index_2046732_comb;
  wire [7:0] p16_array_index_2046733_comb;
  wire [7:0] p16_array_index_2046734_comb;
  wire [7:0] p16_array_index_2046735_comb;
  wire [7:0] p16_res7__202_comb;
  wire [7:0] p16_array_index_2046746_comb;
  wire [7:0] p16_array_index_2046747_comb;
  wire [7:0] p16_array_index_2046748_comb;
  wire [7:0] p16_res7__204_comb;
  wire [7:0] p16_array_index_2046758_comb;
  wire [7:0] p16_array_index_2046759_comb;
  wire [7:0] p16_array_index_2046760_comb;
  wire [7:0] p16_res7__206_comb;
  wire [7:0] p16_array_index_2046771_comb;
  wire [7:0] p16_array_index_2046772_comb;
  wire [7:0] p16_res7__208_comb;
  assign p16_array_index_2046690_comb = p15_literal_2043912[p15_res7__192];
  assign p16_array_index_2046691_comb = p15_literal_2043914[p15_array_index_2046560];
  assign p16_array_index_2046692_comb = p15_literal_2043916[p15_array_index_2046561];
  assign p16_array_index_2046693_comb = p15_literal_2043918[p15_array_index_2046562];
  assign p16_array_index_2046694_comb = p15_literal_2043920[p15_array_index_2046563];
  assign p16_res7__196_comb = p15_literal_2043910[p15_res7__194] ^ p16_array_index_2046690_comb ^ p16_array_index_2046691_comb ^ p16_array_index_2046692_comb ^ p16_array_index_2046693_comb ^ p16_array_index_2046694_comb ^ p15_array_index_2046564 ^ p15_literal_2043923[p15_array_index_2046565] ^ p15_array_index_2046582 ^ p15_literal_2043920[p15_array_index_2046567] ^ p15_literal_2043918[p15_array_index_2046584] ^ p15_literal_2043916[p15_array_index_2046569] ^ p15_literal_2043914[p15_array_index_2046570] ^ p15_literal_2043912[p15_array_index_2046571] ^ p15_literal_2043910[p15_array_index_2046572] ^ p15_array_index_2046573;
  assign p16_array_index_2046704_comb = p15_literal_2043912[p15_res7__194];
  assign p16_array_index_2046705_comb = p15_literal_2043914[p15_res7__192];
  assign p16_array_index_2046706_comb = p15_literal_2043916[p15_array_index_2046560];
  assign p16_array_index_2046707_comb = p15_literal_2043918[p15_array_index_2046561];
  assign p16_array_index_2046708_comb = p15_literal_2043920[p15_array_index_2046562];
  assign p16_res7__198_comb = p15_literal_2043910[p16_res7__196_comb] ^ p16_array_index_2046704_comb ^ p16_array_index_2046705_comb ^ p16_array_index_2046706_comb ^ p16_array_index_2046707_comb ^ p16_array_index_2046708_comb ^ p15_array_index_2046563 ^ p15_literal_2043923[p15_array_index_2046564] ^ p15_array_index_2046565 ^ p15_literal_2043920[p15_array_index_2046582] ^ p15_literal_2043918[p15_array_index_2046567] ^ p15_literal_2043916[p15_array_index_2046584] ^ p15_literal_2043914[p15_array_index_2046569] ^ p15_literal_2043912[p15_array_index_2046570] ^ p15_literal_2043910[p15_array_index_2046571] ^ p15_array_index_2046572;
  assign p16_array_index_2046719_comb = p15_literal_2043914[p15_res7__194];
  assign p16_array_index_2046720_comb = p15_literal_2043916[p15_res7__192];
  assign p16_array_index_2046721_comb = p15_literal_2043918[p15_array_index_2046560];
  assign p16_array_index_2046722_comb = p15_literal_2043920[p15_array_index_2046561];
  assign p16_res7__200_comb = p15_literal_2043910[p16_res7__198_comb] ^ p15_literal_2043912[p16_res7__196_comb] ^ p16_array_index_2046719_comb ^ p16_array_index_2046720_comb ^ p16_array_index_2046721_comb ^ p16_array_index_2046722_comb ^ p15_array_index_2046562 ^ p15_literal_2043923[p15_array_index_2046563] ^ p15_array_index_2046564 ^ p15_array_index_2046581 ^ p15_literal_2043918[p15_array_index_2046582] ^ p15_literal_2043916[p15_array_index_2046567] ^ p15_literal_2043914[p15_array_index_2046584] ^ p15_literal_2043912[p15_array_index_2046569] ^ p15_literal_2043910[p15_array_index_2046570] ^ p15_array_index_2046571;
  assign p16_array_index_2046732_comb = p15_literal_2043914[p16_res7__196_comb];
  assign p16_array_index_2046733_comb = p15_literal_2043916[p15_res7__194];
  assign p16_array_index_2046734_comb = p15_literal_2043918[p15_res7__192];
  assign p16_array_index_2046735_comb = p15_literal_2043920[p15_array_index_2046560];
  assign p16_res7__202_comb = p15_literal_2043910[p16_res7__200_comb] ^ p15_literal_2043912[p16_res7__198_comb] ^ p16_array_index_2046732_comb ^ p16_array_index_2046733_comb ^ p16_array_index_2046734_comb ^ p16_array_index_2046735_comb ^ p15_array_index_2046561 ^ p15_literal_2043923[p15_array_index_2046562] ^ p15_array_index_2046563 ^ p15_array_index_2046598 ^ p15_literal_2043918[p15_array_index_2046565] ^ p15_literal_2043916[p15_array_index_2046582] ^ p15_literal_2043914[p15_array_index_2046567] ^ p15_literal_2043912[p15_array_index_2046584] ^ p15_literal_2043910[p15_array_index_2046569] ^ p15_array_index_2046570;
  assign p16_array_index_2046746_comb = p15_literal_2043916[p16_res7__196_comb];
  assign p16_array_index_2046747_comb = p15_literal_2043918[p15_res7__194];
  assign p16_array_index_2046748_comb = p15_literal_2043920[p15_res7__192];
  assign p16_res7__204_comb = p15_literal_2043910[p16_res7__202_comb] ^ p15_literal_2043912[p16_res7__200_comb] ^ p15_literal_2043914[p16_res7__198_comb] ^ p16_array_index_2046746_comb ^ p16_array_index_2046747_comb ^ p16_array_index_2046748_comb ^ p15_array_index_2046560 ^ p15_literal_2043923[p15_array_index_2046561] ^ p15_array_index_2046562 ^ p16_array_index_2046694_comb ^ p15_array_index_2046580 ^ p15_literal_2043916[p15_array_index_2046565] ^ p15_literal_2043914[p15_array_index_2046582] ^ p15_literal_2043912[p15_array_index_2046567] ^ p15_literal_2043910[p15_array_index_2046584] ^ p15_array_index_2046569;
  assign p16_array_index_2046758_comb = p15_literal_2043916[p16_res7__198_comb];
  assign p16_array_index_2046759_comb = p15_literal_2043918[p16_res7__196_comb];
  assign p16_array_index_2046760_comb = p15_literal_2043920[p15_res7__194];
  assign p16_res7__206_comb = p15_literal_2043910[p16_res7__204_comb] ^ p15_literal_2043912[p16_res7__202_comb] ^ p15_literal_2043914[p16_res7__200_comb] ^ p16_array_index_2046758_comb ^ p16_array_index_2046759_comb ^ p16_array_index_2046760_comb ^ p15_res7__192 ^ p15_literal_2043923[p15_array_index_2046560] ^ p15_array_index_2046561 ^ p16_array_index_2046708_comb ^ p15_array_index_2046597 ^ p15_literal_2043916[p15_array_index_2046564] ^ p15_literal_2043914[p15_array_index_2046565] ^ p15_literal_2043912[p15_array_index_2046582] ^ p15_literal_2043910[p15_array_index_2046567] ^ p15_array_index_2046584;
  assign p16_array_index_2046771_comb = p15_literal_2043918[p16_res7__198_comb];
  assign p16_array_index_2046772_comb = p15_literal_2043920[p16_res7__196_comb];
  assign p16_res7__208_comb = p15_literal_2043910[p16_res7__206_comb] ^ p15_literal_2043912[p16_res7__204_comb] ^ p15_literal_2043914[p16_res7__202_comb] ^ p15_literal_2043916[p16_res7__200_comb] ^ p16_array_index_2046771_comb ^ p16_array_index_2046772_comb ^ p15_res7__194 ^ p15_literal_2043923[p15_res7__192] ^ p15_array_index_2046560 ^ p16_array_index_2046722_comb ^ p16_array_index_2046693_comb ^ p15_array_index_2046579 ^ p15_literal_2043914[p15_array_index_2046564] ^ p15_literal_2043912[p15_array_index_2046565] ^ p15_literal_2043910[p15_array_index_2046582] ^ p15_array_index_2046567;

  // Registers for pipe stage 16:
  reg [127:0] p16_encoded;
  reg [127:0] p16_bit_slice_2043893;
  reg [127:0] p16_bit_slice_2044018;
  reg [127:0] p16_xor_2046116;
  reg [127:0] p16_xor_2046544;
  reg [7:0] p16_array_index_2046560;
  reg [7:0] p16_array_index_2046561;
  reg [7:0] p16_array_index_2046562;
  reg [7:0] p16_array_index_2046563;
  reg [7:0] p16_array_index_2046564;
  reg [7:0] p16_array_index_2046565;
  reg [7:0] p16_array_index_2046576;
  reg [7:0] p16_array_index_2046577;
  reg [7:0] p16_array_index_2046578;
  reg [7:0] p16_array_index_2046582;
  reg [7:0] p16_res7__192;
  reg [7:0] p16_array_index_2046593;
  reg [7:0] p16_array_index_2046594;
  reg [7:0] p16_array_index_2046595;
  reg [7:0] p16_array_index_2046596;
  reg [7:0] p16_res7__194;
  reg [7:0] p16_array_index_2046690;
  reg [7:0] p16_array_index_2046691;
  reg [7:0] p16_array_index_2046692;
  reg [7:0] p16_res7__196;
  reg [7:0] p16_array_index_2046704;
  reg [7:0] p16_array_index_2046705;
  reg [7:0] p16_array_index_2046706;
  reg [7:0] p16_array_index_2046707;
  reg [7:0] p16_res7__198;
  reg [7:0] p16_array_index_2046719;
  reg [7:0] p16_array_index_2046720;
  reg [7:0] p16_array_index_2046721;
  reg [7:0] p16_res7__200;
  reg [7:0] p16_array_index_2046732;
  reg [7:0] p16_array_index_2046733;
  reg [7:0] p16_array_index_2046734;
  reg [7:0] p16_array_index_2046735;
  reg [7:0] p16_res7__202;
  reg [7:0] p16_array_index_2046746;
  reg [7:0] p16_array_index_2046747;
  reg [7:0] p16_array_index_2046748;
  reg [7:0] p16_res7__204;
  reg [7:0] p16_array_index_2046758;
  reg [7:0] p16_array_index_2046759;
  reg [7:0] p16_array_index_2046760;
  reg [7:0] p16_res7__206;
  reg [7:0] p16_array_index_2046771;
  reg [7:0] p16_array_index_2046772;
  reg [7:0] p16_res7__208;
  reg [7:0] p17_literal_2043896[256];
  reg [7:0] p17_literal_2043910[256];
  reg [7:0] p17_literal_2043912[256];
  reg [7:0] p17_literal_2043914[256];
  reg [7:0] p17_literal_2043916[256];
  reg [7:0] p17_literal_2043918[256];
  reg [7:0] p17_literal_2043920[256];
  reg [7:0] p17_literal_2043923[256];
  reg [7:0] p94_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p16_encoded <= p15_encoded;
    p16_bit_slice_2043893 <= p15_bit_slice_2043893;
    p16_bit_slice_2044018 <= p15_bit_slice_2044018;
    p16_xor_2046116 <= p15_xor_2046116;
    p16_xor_2046544 <= p15_xor_2046544;
    p16_array_index_2046560 <= p15_array_index_2046560;
    p16_array_index_2046561 <= p15_array_index_2046561;
    p16_array_index_2046562 <= p15_array_index_2046562;
    p16_array_index_2046563 <= p15_array_index_2046563;
    p16_array_index_2046564 <= p15_array_index_2046564;
    p16_array_index_2046565 <= p15_array_index_2046565;
    p16_array_index_2046576 <= p15_array_index_2046576;
    p16_array_index_2046577 <= p15_array_index_2046577;
    p16_array_index_2046578 <= p15_array_index_2046578;
    p16_array_index_2046582 <= p15_array_index_2046582;
    p16_res7__192 <= p15_res7__192;
    p16_array_index_2046593 <= p15_array_index_2046593;
    p16_array_index_2046594 <= p15_array_index_2046594;
    p16_array_index_2046595 <= p15_array_index_2046595;
    p16_array_index_2046596 <= p15_array_index_2046596;
    p16_res7__194 <= p15_res7__194;
    p16_array_index_2046690 <= p16_array_index_2046690_comb;
    p16_array_index_2046691 <= p16_array_index_2046691_comb;
    p16_array_index_2046692 <= p16_array_index_2046692_comb;
    p16_res7__196 <= p16_res7__196_comb;
    p16_array_index_2046704 <= p16_array_index_2046704_comb;
    p16_array_index_2046705 <= p16_array_index_2046705_comb;
    p16_array_index_2046706 <= p16_array_index_2046706_comb;
    p16_array_index_2046707 <= p16_array_index_2046707_comb;
    p16_res7__198 <= p16_res7__198_comb;
    p16_array_index_2046719 <= p16_array_index_2046719_comb;
    p16_array_index_2046720 <= p16_array_index_2046720_comb;
    p16_array_index_2046721 <= p16_array_index_2046721_comb;
    p16_res7__200 <= p16_res7__200_comb;
    p16_array_index_2046732 <= p16_array_index_2046732_comb;
    p16_array_index_2046733 <= p16_array_index_2046733_comb;
    p16_array_index_2046734 <= p16_array_index_2046734_comb;
    p16_array_index_2046735 <= p16_array_index_2046735_comb;
    p16_res7__202 <= p16_res7__202_comb;
    p16_array_index_2046746 <= p16_array_index_2046746_comb;
    p16_array_index_2046747 <= p16_array_index_2046747_comb;
    p16_array_index_2046748 <= p16_array_index_2046748_comb;
    p16_res7__204 <= p16_res7__204_comb;
    p16_array_index_2046758 <= p16_array_index_2046758_comb;
    p16_array_index_2046759 <= p16_array_index_2046759_comb;
    p16_array_index_2046760 <= p16_array_index_2046760_comb;
    p16_res7__206 <= p16_res7__206_comb;
    p16_array_index_2046771 <= p16_array_index_2046771_comb;
    p16_array_index_2046772 <= p16_array_index_2046772_comb;
    p16_res7__208 <= p16_res7__208_comb;
    p17_literal_2043896 <= p16_literal_2043896;
    p17_literal_2043910 <= p16_literal_2043910;
    p17_literal_2043912 <= p16_literal_2043912;
    p17_literal_2043914 <= p16_literal_2043914;
    p17_literal_2043916 <= p16_literal_2043916;
    p17_literal_2043918 <= p16_literal_2043918;
    p17_literal_2043920 <= p16_literal_2043920;
    p17_literal_2043923 <= p16_literal_2043923;
    p94_literal_2058836 <= p93_literal_2058836;
  end

  // ===== Pipe stage 17:
  wire [7:0] p17_array_index_2046898_comb;
  wire [7:0] p17_array_index_2046899_comb;
  wire [7:0] p17_res7__210_comb;
  wire [7:0] p17_array_index_2046910_comb;
  wire [7:0] p17_res7__212_comb;
  wire [7:0] p17_array_index_2046920_comb;
  wire [7:0] p17_res7__214_comb;
  wire [7:0] p17_res7__216_comb;
  wire [7:0] p17_res7__218_comb;
  wire [7:0] p17_res7__220_comb;
  wire [7:0] p17_res7__222_comb;
  wire [127:0] p17_res__6_comb;
  assign p17_array_index_2046898_comb = p16_literal_2043918[p16_res7__200];
  assign p17_array_index_2046899_comb = p16_literal_2043920[p16_res7__198];
  assign p17_res7__210_comb = p16_literal_2043910[p16_res7__208] ^ p16_literal_2043912[p16_res7__206] ^ p16_literal_2043914[p16_res7__204] ^ p16_literal_2043916[p16_res7__202] ^ p17_array_index_2046898_comb ^ p17_array_index_2046899_comb ^ p16_res7__196 ^ p16_literal_2043923[p16_res7__194] ^ p16_res7__192 ^ p16_array_index_2046735 ^ p16_array_index_2046707 ^ p16_array_index_2046596 ^ p16_literal_2043914[p16_array_index_2046563] ^ p16_literal_2043912[p16_array_index_2046564] ^ p16_literal_2043910[p16_array_index_2046565] ^ p16_array_index_2046582;
  assign p17_array_index_2046910_comb = p16_literal_2043920[p16_res7__200];
  assign p17_res7__212_comb = p16_literal_2043910[p17_res7__210_comb] ^ p16_literal_2043912[p16_res7__208] ^ p16_literal_2043914[p16_res7__206] ^ p16_literal_2043916[p16_res7__204] ^ p16_literal_2043918[p16_res7__202] ^ p17_array_index_2046910_comb ^ p16_res7__198 ^ p16_literal_2043923[p16_res7__196] ^ p16_res7__194 ^ p16_array_index_2046748 ^ p16_array_index_2046721 ^ p16_array_index_2046692 ^ p16_array_index_2046578 ^ p16_literal_2043912[p16_array_index_2046563] ^ p16_literal_2043910[p16_array_index_2046564] ^ p16_array_index_2046565;
  assign p17_array_index_2046920_comb = p16_literal_2043920[p16_res7__202];
  assign p17_res7__214_comb = p16_literal_2043910[p17_res7__212_comb] ^ p16_literal_2043912[p17_res7__210_comb] ^ p16_literal_2043914[p16_res7__208] ^ p16_literal_2043916[p16_res7__206] ^ p16_literal_2043918[p16_res7__204] ^ p17_array_index_2046920_comb ^ p16_res7__200 ^ p16_literal_2043923[p16_res7__198] ^ p16_res7__196 ^ p16_array_index_2046760 ^ p16_array_index_2046734 ^ p16_array_index_2046706 ^ p16_array_index_2046595 ^ p16_literal_2043912[p16_array_index_2046562] ^ p16_literal_2043910[p16_array_index_2046563] ^ p16_array_index_2046564;
  assign p17_res7__216_comb = p16_literal_2043910[p17_res7__214_comb] ^ p16_literal_2043912[p17_res7__212_comb] ^ p16_literal_2043914[p17_res7__210_comb] ^ p16_literal_2043916[p16_res7__208] ^ p16_literal_2043918[p16_res7__206] ^ p16_literal_2043920[p16_res7__204] ^ p16_res7__202 ^ p16_literal_2043923[p16_res7__200] ^ p16_res7__198 ^ p16_array_index_2046772 ^ p16_array_index_2046747 ^ p16_array_index_2046720 ^ p16_array_index_2046691 ^ p16_array_index_2046577 ^ p16_literal_2043910[p16_array_index_2046562] ^ p16_array_index_2046563;
  assign p17_res7__218_comb = p16_literal_2043910[p17_res7__216_comb] ^ p16_literal_2043912[p17_res7__214_comb] ^ p16_literal_2043914[p17_res7__212_comb] ^ p16_literal_2043916[p17_res7__210_comb] ^ p16_literal_2043918[p16_res7__208] ^ p16_literal_2043920[p16_res7__206] ^ p16_res7__204 ^ p16_literal_2043923[p16_res7__202] ^ p16_res7__200 ^ p17_array_index_2046899_comb ^ p16_array_index_2046759 ^ p16_array_index_2046733 ^ p16_array_index_2046705 ^ p16_array_index_2046594 ^ p16_literal_2043910[p16_array_index_2046561] ^ p16_array_index_2046562;
  assign p17_res7__220_comb = p16_literal_2043910[p17_res7__218_comb] ^ p16_literal_2043912[p17_res7__216_comb] ^ p16_literal_2043914[p17_res7__214_comb] ^ p16_literal_2043916[p17_res7__212_comb] ^ p16_literal_2043918[p17_res7__210_comb] ^ p16_literal_2043920[p16_res7__208] ^ p16_res7__206 ^ p16_literal_2043923[p16_res7__204] ^ p16_res7__202 ^ p17_array_index_2046910_comb ^ p16_array_index_2046771 ^ p16_array_index_2046746 ^ p16_array_index_2046719 ^ p16_array_index_2046690 ^ p16_array_index_2046576 ^ p16_array_index_2046561;
  assign p17_res7__222_comb = p16_literal_2043910[p17_res7__220_comb] ^ p16_literal_2043912[p17_res7__218_comb] ^ p16_literal_2043914[p17_res7__216_comb] ^ p16_literal_2043916[p17_res7__214_comb] ^ p16_literal_2043918[p17_res7__212_comb] ^ p16_literal_2043920[p17_res7__210_comb] ^ p16_res7__208 ^ p16_literal_2043923[p16_res7__206] ^ p16_res7__204 ^ p17_array_index_2046920_comb ^ p17_array_index_2046898_comb ^ p16_array_index_2046758 ^ p16_array_index_2046732 ^ p16_array_index_2046704 ^ p16_array_index_2046593 ^ p16_array_index_2046560;
  assign p17_res__6_comb = {p17_res7__222_comb, p17_res7__220_comb, p17_res7__218_comb, p17_res7__216_comb, p17_res7__214_comb, p17_res7__212_comb, p17_res7__210_comb, p16_res7__208, p16_res7__206, p16_res7__204, p16_res7__202, p16_res7__200, p16_res7__198, p16_res7__196, p16_res7__194, p16_res7__192};

  // Registers for pipe stage 17:
  reg [127:0] p17_encoded;
  reg [127:0] p17_bit_slice_2043893;
  reg [127:0] p17_bit_slice_2044018;
  reg [127:0] p17_xor_2046116;
  reg [127:0] p17_xor_2046544;
  reg [127:0] p17_res__6;
  reg [7:0] p18_literal_2043896[256];
  reg [7:0] p18_literal_2043910[256];
  reg [7:0] p18_literal_2043912[256];
  reg [7:0] p18_literal_2043914[256];
  reg [7:0] p18_literal_2043916[256];
  reg [7:0] p18_literal_2043918[256];
  reg [7:0] p18_literal_2043920[256];
  reg [7:0] p18_literal_2043923[256];
  reg [7:0] p95_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p17_encoded <= p16_encoded;
    p17_bit_slice_2043893 <= p16_bit_slice_2043893;
    p17_bit_slice_2044018 <= p16_bit_slice_2044018;
    p17_xor_2046116 <= p16_xor_2046116;
    p17_xor_2046544 <= p16_xor_2046544;
    p17_res__6 <= p17_res__6_comb;
    p18_literal_2043896 <= p17_literal_2043896;
    p18_literal_2043910 <= p17_literal_2043910;
    p18_literal_2043912 <= p17_literal_2043912;
    p18_literal_2043914 <= p17_literal_2043914;
    p18_literal_2043916 <= p17_literal_2043916;
    p18_literal_2043918 <= p17_literal_2043918;
    p18_literal_2043920 <= p17_literal_2043920;
    p18_literal_2043923 <= p17_literal_2043923;
    p95_literal_2058836 <= p94_literal_2058836;
  end

  // ===== Pipe stage 18:
  wire [127:0] p18_k3_comb;
  wire [127:0] p18_addedKey__39_comb;
  wire [7:0] p18_array_index_2047004_comb;
  wire [7:0] p18_array_index_2047005_comb;
  wire [7:0] p18_array_index_2047006_comb;
  wire [7:0] p18_array_index_2047007_comb;
  wire [7:0] p18_array_index_2047008_comb;
  wire [7:0] p18_array_index_2047009_comb;
  wire [7:0] p18_array_index_2047011_comb;
  wire [7:0] p18_array_index_2047013_comb;
  wire [7:0] p18_array_index_2047014_comb;
  wire [7:0] p18_array_index_2047015_comb;
  wire [7:0] p18_array_index_2047016_comb;
  wire [7:0] p18_array_index_2047017_comb;
  wire [7:0] p18_array_index_2047018_comb;
  wire [7:0] p18_array_index_2047020_comb;
  wire [7:0] p18_array_index_2047021_comb;
  wire [7:0] p18_array_index_2047022_comb;
  wire [7:0] p18_array_index_2047023_comb;
  wire [7:0] p18_array_index_2047024_comb;
  wire [7:0] p18_array_index_2047025_comb;
  wire [7:0] p18_array_index_2047026_comb;
  wire [7:0] p18_array_index_2047028_comb;
  wire [7:0] p18_res7__224_comb;
  wire [7:0] p18_array_index_2047037_comb;
  wire [7:0] p18_array_index_2047038_comb;
  wire [7:0] p18_array_index_2047039_comb;
  wire [7:0] p18_array_index_2047040_comb;
  wire [7:0] p18_array_index_2047041_comb;
  wire [7:0] p18_array_index_2047042_comb;
  wire [7:0] p18_res7__226_comb;
  wire [7:0] p18_array_index_2047052_comb;
  wire [7:0] p18_array_index_2047053_comb;
  wire [7:0] p18_array_index_2047054_comb;
  wire [7:0] p18_array_index_2047055_comb;
  wire [7:0] p18_array_index_2047056_comb;
  wire [7:0] p18_res7__228_comb;
  wire [7:0] p18_array_index_2047066_comb;
  wire [7:0] p18_array_index_2047067_comb;
  wire [7:0] p18_array_index_2047068_comb;
  wire [7:0] p18_array_index_2047069_comb;
  wire [7:0] p18_array_index_2047070_comb;
  wire [7:0] p18_res7__230_comb;
  wire [7:0] p18_array_index_2047081_comb;
  wire [7:0] p18_array_index_2047082_comb;
  wire [7:0] p18_array_index_2047083_comb;
  wire [7:0] p18_array_index_2047084_comb;
  wire [7:0] p18_res7__232_comb;
  wire [7:0] p18_array_index_2047094_comb;
  wire [7:0] p18_array_index_2047095_comb;
  wire [7:0] p18_array_index_2047096_comb;
  wire [7:0] p18_array_index_2047097_comb;
  wire [7:0] p18_res7__234_comb;
  assign p18_k3_comb = p17_res__6 ^ p17_xor_2046116;
  assign p18_addedKey__39_comb = p18_k3_comb ^ 128'hf659_3616_e605_5689_adfb_a180_27aa_2a08;
  assign p18_array_index_2047004_comb = p17_literal_2043896[p18_addedKey__39_comb[127:120]];
  assign p18_array_index_2047005_comb = p17_literal_2043896[p18_addedKey__39_comb[119:112]];
  assign p18_array_index_2047006_comb = p17_literal_2043896[p18_addedKey__39_comb[111:104]];
  assign p18_array_index_2047007_comb = p17_literal_2043896[p18_addedKey__39_comb[103:96]];
  assign p18_array_index_2047008_comb = p17_literal_2043896[p18_addedKey__39_comb[95:88]];
  assign p18_array_index_2047009_comb = p17_literal_2043896[p18_addedKey__39_comb[87:80]];
  assign p18_array_index_2047011_comb = p17_literal_2043896[p18_addedKey__39_comb[71:64]];
  assign p18_array_index_2047013_comb = p17_literal_2043896[p18_addedKey__39_comb[55:48]];
  assign p18_array_index_2047014_comb = p17_literal_2043896[p18_addedKey__39_comb[47:40]];
  assign p18_array_index_2047015_comb = p17_literal_2043896[p18_addedKey__39_comb[39:32]];
  assign p18_array_index_2047016_comb = p17_literal_2043896[p18_addedKey__39_comb[31:24]];
  assign p18_array_index_2047017_comb = p17_literal_2043896[p18_addedKey__39_comb[23:16]];
  assign p18_array_index_2047018_comb = p17_literal_2043896[p18_addedKey__39_comb[15:8]];
  assign p18_array_index_2047020_comb = p17_literal_2043910[p18_array_index_2047004_comb];
  assign p18_array_index_2047021_comb = p17_literal_2043912[p18_array_index_2047005_comb];
  assign p18_array_index_2047022_comb = p17_literal_2043914[p18_array_index_2047006_comb];
  assign p18_array_index_2047023_comb = p17_literal_2043916[p18_array_index_2047007_comb];
  assign p18_array_index_2047024_comb = p17_literal_2043918[p18_array_index_2047008_comb];
  assign p18_array_index_2047025_comb = p17_literal_2043920[p18_array_index_2047009_comb];
  assign p18_array_index_2047026_comb = p17_literal_2043896[p18_addedKey__39_comb[79:72]];
  assign p18_array_index_2047028_comb = p17_literal_2043896[p18_addedKey__39_comb[63:56]];
  assign p18_res7__224_comb = p18_array_index_2047020_comb ^ p18_array_index_2047021_comb ^ p18_array_index_2047022_comb ^ p18_array_index_2047023_comb ^ p18_array_index_2047024_comb ^ p18_array_index_2047025_comb ^ p18_array_index_2047026_comb ^ p17_literal_2043923[p18_array_index_2047011_comb] ^ p18_array_index_2047028_comb ^ p17_literal_2043920[p18_array_index_2047013_comb] ^ p17_literal_2043918[p18_array_index_2047014_comb] ^ p17_literal_2043916[p18_array_index_2047015_comb] ^ p17_literal_2043914[p18_array_index_2047016_comb] ^ p17_literal_2043912[p18_array_index_2047017_comb] ^ p17_literal_2043910[p18_array_index_2047018_comb] ^ p17_literal_2043896[p18_addedKey__39_comb[7:0]];
  assign p18_array_index_2047037_comb = p17_literal_2043910[p18_res7__224_comb];
  assign p18_array_index_2047038_comb = p17_literal_2043912[p18_array_index_2047004_comb];
  assign p18_array_index_2047039_comb = p17_literal_2043914[p18_array_index_2047005_comb];
  assign p18_array_index_2047040_comb = p17_literal_2043916[p18_array_index_2047006_comb];
  assign p18_array_index_2047041_comb = p17_literal_2043918[p18_array_index_2047007_comb];
  assign p18_array_index_2047042_comb = p17_literal_2043920[p18_array_index_2047008_comb];
  assign p18_res7__226_comb = p18_array_index_2047037_comb ^ p18_array_index_2047038_comb ^ p18_array_index_2047039_comb ^ p18_array_index_2047040_comb ^ p18_array_index_2047041_comb ^ p18_array_index_2047042_comb ^ p18_array_index_2047009_comb ^ p17_literal_2043923[p18_array_index_2047026_comb] ^ p18_array_index_2047011_comb ^ p17_literal_2043920[p18_array_index_2047028_comb] ^ p17_literal_2043918[p18_array_index_2047013_comb] ^ p17_literal_2043916[p18_array_index_2047014_comb] ^ p17_literal_2043914[p18_array_index_2047015_comb] ^ p17_literal_2043912[p18_array_index_2047016_comb] ^ p17_literal_2043910[p18_array_index_2047017_comb] ^ p18_array_index_2047018_comb;
  assign p18_array_index_2047052_comb = p17_literal_2043912[p18_res7__224_comb];
  assign p18_array_index_2047053_comb = p17_literal_2043914[p18_array_index_2047004_comb];
  assign p18_array_index_2047054_comb = p17_literal_2043916[p18_array_index_2047005_comb];
  assign p18_array_index_2047055_comb = p17_literal_2043918[p18_array_index_2047006_comb];
  assign p18_array_index_2047056_comb = p17_literal_2043920[p18_array_index_2047007_comb];
  assign p18_res7__228_comb = p17_literal_2043910[p18_res7__226_comb] ^ p18_array_index_2047052_comb ^ p18_array_index_2047053_comb ^ p18_array_index_2047054_comb ^ p18_array_index_2047055_comb ^ p18_array_index_2047056_comb ^ p18_array_index_2047008_comb ^ p17_literal_2043923[p18_array_index_2047009_comb] ^ p18_array_index_2047026_comb ^ p17_literal_2043920[p18_array_index_2047011_comb] ^ p17_literal_2043918[p18_array_index_2047028_comb] ^ p17_literal_2043916[p18_array_index_2047013_comb] ^ p17_literal_2043914[p18_array_index_2047014_comb] ^ p17_literal_2043912[p18_array_index_2047015_comb] ^ p17_literal_2043910[p18_array_index_2047016_comb] ^ p18_array_index_2047017_comb;
  assign p18_array_index_2047066_comb = p17_literal_2043912[p18_res7__226_comb];
  assign p18_array_index_2047067_comb = p17_literal_2043914[p18_res7__224_comb];
  assign p18_array_index_2047068_comb = p17_literal_2043916[p18_array_index_2047004_comb];
  assign p18_array_index_2047069_comb = p17_literal_2043918[p18_array_index_2047005_comb];
  assign p18_array_index_2047070_comb = p17_literal_2043920[p18_array_index_2047006_comb];
  assign p18_res7__230_comb = p17_literal_2043910[p18_res7__228_comb] ^ p18_array_index_2047066_comb ^ p18_array_index_2047067_comb ^ p18_array_index_2047068_comb ^ p18_array_index_2047069_comb ^ p18_array_index_2047070_comb ^ p18_array_index_2047007_comb ^ p17_literal_2043923[p18_array_index_2047008_comb] ^ p18_array_index_2047009_comb ^ p17_literal_2043920[p18_array_index_2047026_comb] ^ p17_literal_2043918[p18_array_index_2047011_comb] ^ p17_literal_2043916[p18_array_index_2047028_comb] ^ p17_literal_2043914[p18_array_index_2047013_comb] ^ p17_literal_2043912[p18_array_index_2047014_comb] ^ p17_literal_2043910[p18_array_index_2047015_comb] ^ p18_array_index_2047016_comb;
  assign p18_array_index_2047081_comb = p17_literal_2043914[p18_res7__226_comb];
  assign p18_array_index_2047082_comb = p17_literal_2043916[p18_res7__224_comb];
  assign p18_array_index_2047083_comb = p17_literal_2043918[p18_array_index_2047004_comb];
  assign p18_array_index_2047084_comb = p17_literal_2043920[p18_array_index_2047005_comb];
  assign p18_res7__232_comb = p17_literal_2043910[p18_res7__230_comb] ^ p17_literal_2043912[p18_res7__228_comb] ^ p18_array_index_2047081_comb ^ p18_array_index_2047082_comb ^ p18_array_index_2047083_comb ^ p18_array_index_2047084_comb ^ p18_array_index_2047006_comb ^ p17_literal_2043923[p18_array_index_2047007_comb] ^ p18_array_index_2047008_comb ^ p18_array_index_2047025_comb ^ p17_literal_2043918[p18_array_index_2047026_comb] ^ p17_literal_2043916[p18_array_index_2047011_comb] ^ p17_literal_2043914[p18_array_index_2047028_comb] ^ p17_literal_2043912[p18_array_index_2047013_comb] ^ p17_literal_2043910[p18_array_index_2047014_comb] ^ p18_array_index_2047015_comb;
  assign p18_array_index_2047094_comb = p17_literal_2043914[p18_res7__228_comb];
  assign p18_array_index_2047095_comb = p17_literal_2043916[p18_res7__226_comb];
  assign p18_array_index_2047096_comb = p17_literal_2043918[p18_res7__224_comb];
  assign p18_array_index_2047097_comb = p17_literal_2043920[p18_array_index_2047004_comb];
  assign p18_res7__234_comb = p17_literal_2043910[p18_res7__232_comb] ^ p17_literal_2043912[p18_res7__230_comb] ^ p18_array_index_2047094_comb ^ p18_array_index_2047095_comb ^ p18_array_index_2047096_comb ^ p18_array_index_2047097_comb ^ p18_array_index_2047005_comb ^ p17_literal_2043923[p18_array_index_2047006_comb] ^ p18_array_index_2047007_comb ^ p18_array_index_2047042_comb ^ p17_literal_2043918[p18_array_index_2047009_comb] ^ p17_literal_2043916[p18_array_index_2047026_comb] ^ p17_literal_2043914[p18_array_index_2047011_comb] ^ p17_literal_2043912[p18_array_index_2047028_comb] ^ p17_literal_2043910[p18_array_index_2047013_comb] ^ p18_array_index_2047014_comb;

  // Registers for pipe stage 18:
  reg [127:0] p18_encoded;
  reg [127:0] p18_bit_slice_2043893;
  reg [127:0] p18_bit_slice_2044018;
  reg [127:0] p18_xor_2046544;
  reg [127:0] p18_k3;
  reg [7:0] p18_array_index_2047004;
  reg [7:0] p18_array_index_2047005;
  reg [7:0] p18_array_index_2047006;
  reg [7:0] p18_array_index_2047007;
  reg [7:0] p18_array_index_2047008;
  reg [7:0] p18_array_index_2047009;
  reg [7:0] p18_array_index_2047011;
  reg [7:0] p18_array_index_2047013;
  reg [7:0] p18_array_index_2047020;
  reg [7:0] p18_array_index_2047021;
  reg [7:0] p18_array_index_2047022;
  reg [7:0] p18_array_index_2047023;
  reg [7:0] p18_array_index_2047024;
  reg [7:0] p18_array_index_2047026;
  reg [7:0] p18_array_index_2047028;
  reg [7:0] p18_res7__224;
  reg [7:0] p18_array_index_2047037;
  reg [7:0] p18_array_index_2047038;
  reg [7:0] p18_array_index_2047039;
  reg [7:0] p18_array_index_2047040;
  reg [7:0] p18_array_index_2047041;
  reg [7:0] p18_res7__226;
  reg [7:0] p18_array_index_2047052;
  reg [7:0] p18_array_index_2047053;
  reg [7:0] p18_array_index_2047054;
  reg [7:0] p18_array_index_2047055;
  reg [7:0] p18_array_index_2047056;
  reg [7:0] p18_res7__228;
  reg [7:0] p18_array_index_2047066;
  reg [7:0] p18_array_index_2047067;
  reg [7:0] p18_array_index_2047068;
  reg [7:0] p18_array_index_2047069;
  reg [7:0] p18_array_index_2047070;
  reg [7:0] p18_res7__230;
  reg [7:0] p18_array_index_2047081;
  reg [7:0] p18_array_index_2047082;
  reg [7:0] p18_array_index_2047083;
  reg [7:0] p18_array_index_2047084;
  reg [7:0] p18_res7__232;
  reg [7:0] p18_array_index_2047094;
  reg [7:0] p18_array_index_2047095;
  reg [7:0] p18_array_index_2047096;
  reg [7:0] p18_array_index_2047097;
  reg [7:0] p18_res7__234;
  reg [7:0] p19_literal_2043896[256];
  reg [7:0] p19_literal_2043910[256];
  reg [7:0] p19_literal_2043912[256];
  reg [7:0] p19_literal_2043914[256];
  reg [7:0] p19_literal_2043916[256];
  reg [7:0] p19_literal_2043918[256];
  reg [7:0] p19_literal_2043920[256];
  reg [7:0] p19_literal_2043923[256];
  reg [7:0] p96_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p18_encoded <= p17_encoded;
    p18_bit_slice_2043893 <= p17_bit_slice_2043893;
    p18_bit_slice_2044018 <= p17_bit_slice_2044018;
    p18_xor_2046544 <= p17_xor_2046544;
    p18_k3 <= p18_k3_comb;
    p18_array_index_2047004 <= p18_array_index_2047004_comb;
    p18_array_index_2047005 <= p18_array_index_2047005_comb;
    p18_array_index_2047006 <= p18_array_index_2047006_comb;
    p18_array_index_2047007 <= p18_array_index_2047007_comb;
    p18_array_index_2047008 <= p18_array_index_2047008_comb;
    p18_array_index_2047009 <= p18_array_index_2047009_comb;
    p18_array_index_2047011 <= p18_array_index_2047011_comb;
    p18_array_index_2047013 <= p18_array_index_2047013_comb;
    p18_array_index_2047020 <= p18_array_index_2047020_comb;
    p18_array_index_2047021 <= p18_array_index_2047021_comb;
    p18_array_index_2047022 <= p18_array_index_2047022_comb;
    p18_array_index_2047023 <= p18_array_index_2047023_comb;
    p18_array_index_2047024 <= p18_array_index_2047024_comb;
    p18_array_index_2047026 <= p18_array_index_2047026_comb;
    p18_array_index_2047028 <= p18_array_index_2047028_comb;
    p18_res7__224 <= p18_res7__224_comb;
    p18_array_index_2047037 <= p18_array_index_2047037_comb;
    p18_array_index_2047038 <= p18_array_index_2047038_comb;
    p18_array_index_2047039 <= p18_array_index_2047039_comb;
    p18_array_index_2047040 <= p18_array_index_2047040_comb;
    p18_array_index_2047041 <= p18_array_index_2047041_comb;
    p18_res7__226 <= p18_res7__226_comb;
    p18_array_index_2047052 <= p18_array_index_2047052_comb;
    p18_array_index_2047053 <= p18_array_index_2047053_comb;
    p18_array_index_2047054 <= p18_array_index_2047054_comb;
    p18_array_index_2047055 <= p18_array_index_2047055_comb;
    p18_array_index_2047056 <= p18_array_index_2047056_comb;
    p18_res7__228 <= p18_res7__228_comb;
    p18_array_index_2047066 <= p18_array_index_2047066_comb;
    p18_array_index_2047067 <= p18_array_index_2047067_comb;
    p18_array_index_2047068 <= p18_array_index_2047068_comb;
    p18_array_index_2047069 <= p18_array_index_2047069_comb;
    p18_array_index_2047070 <= p18_array_index_2047070_comb;
    p18_res7__230 <= p18_res7__230_comb;
    p18_array_index_2047081 <= p18_array_index_2047081_comb;
    p18_array_index_2047082 <= p18_array_index_2047082_comb;
    p18_array_index_2047083 <= p18_array_index_2047083_comb;
    p18_array_index_2047084 <= p18_array_index_2047084_comb;
    p18_res7__232 <= p18_res7__232_comb;
    p18_array_index_2047094 <= p18_array_index_2047094_comb;
    p18_array_index_2047095 <= p18_array_index_2047095_comb;
    p18_array_index_2047096 <= p18_array_index_2047096_comb;
    p18_array_index_2047097 <= p18_array_index_2047097_comb;
    p18_res7__234 <= p18_res7__234_comb;
    p19_literal_2043896 <= p18_literal_2043896;
    p19_literal_2043910 <= p18_literal_2043910;
    p19_literal_2043912 <= p18_literal_2043912;
    p19_literal_2043914 <= p18_literal_2043914;
    p19_literal_2043916 <= p18_literal_2043916;
    p19_literal_2043918 <= p18_literal_2043918;
    p19_literal_2043920 <= p18_literal_2043920;
    p19_literal_2043923 <= p18_literal_2043923;
    p96_literal_2058836 <= p95_literal_2058836;
  end

  // ===== Pipe stage 19:
  wire [7:0] p19_array_index_2047222_comb;
  wire [7:0] p19_array_index_2047223_comb;
  wire [7:0] p19_array_index_2047224_comb;
  wire [7:0] p19_res7__236_comb;
  wire [7:0] p19_array_index_2047234_comb;
  wire [7:0] p19_array_index_2047235_comb;
  wire [7:0] p19_array_index_2047236_comb;
  wire [7:0] p19_res7__238_comb;
  wire [7:0] p19_array_index_2047247_comb;
  wire [7:0] p19_array_index_2047248_comb;
  wire [7:0] p19_res7__240_comb;
  wire [7:0] p19_array_index_2047258_comb;
  wire [7:0] p19_array_index_2047259_comb;
  wire [7:0] p19_res7__242_comb;
  wire [7:0] p19_array_index_2047270_comb;
  wire [7:0] p19_res7__244_comb;
  wire [7:0] p19_array_index_2047280_comb;
  wire [7:0] p19_res7__246_comb;
  wire [7:0] p19_res7__248_comb;
  assign p19_array_index_2047222_comb = p18_literal_2043916[p18_res7__228];
  assign p19_array_index_2047223_comb = p18_literal_2043918[p18_res7__226];
  assign p19_array_index_2047224_comb = p18_literal_2043920[p18_res7__224];
  assign p19_res7__236_comb = p18_literal_2043910[p18_res7__234] ^ p18_literal_2043912[p18_res7__232] ^ p18_literal_2043914[p18_res7__230] ^ p19_array_index_2047222_comb ^ p19_array_index_2047223_comb ^ p19_array_index_2047224_comb ^ p18_array_index_2047004 ^ p18_literal_2043923[p18_array_index_2047005] ^ p18_array_index_2047006 ^ p18_array_index_2047056 ^ p18_array_index_2047024 ^ p18_literal_2043916[p18_array_index_2047009] ^ p18_literal_2043914[p18_array_index_2047026] ^ p18_literal_2043912[p18_array_index_2047011] ^ p18_literal_2043910[p18_array_index_2047028] ^ p18_array_index_2047013;
  assign p19_array_index_2047234_comb = p18_literal_2043916[p18_res7__230];
  assign p19_array_index_2047235_comb = p18_literal_2043918[p18_res7__228];
  assign p19_array_index_2047236_comb = p18_literal_2043920[p18_res7__226];
  assign p19_res7__238_comb = p18_literal_2043910[p19_res7__236_comb] ^ p18_literal_2043912[p18_res7__234] ^ p18_literal_2043914[p18_res7__232] ^ p19_array_index_2047234_comb ^ p19_array_index_2047235_comb ^ p19_array_index_2047236_comb ^ p18_res7__224 ^ p18_literal_2043923[p18_array_index_2047004] ^ p18_array_index_2047005 ^ p18_array_index_2047070 ^ p18_array_index_2047041 ^ p18_literal_2043916[p18_array_index_2047008] ^ p18_literal_2043914[p18_array_index_2047009] ^ p18_literal_2043912[p18_array_index_2047026] ^ p18_literal_2043910[p18_array_index_2047011] ^ p18_array_index_2047028;
  assign p19_array_index_2047247_comb = p18_literal_2043918[p18_res7__230];
  assign p19_array_index_2047248_comb = p18_literal_2043920[p18_res7__228];
  assign p19_res7__240_comb = p18_literal_2043910[p19_res7__238_comb] ^ p18_literal_2043912[p19_res7__236_comb] ^ p18_literal_2043914[p18_res7__234] ^ p18_literal_2043916[p18_res7__232] ^ p19_array_index_2047247_comb ^ p19_array_index_2047248_comb ^ p18_res7__226 ^ p18_literal_2043923[p18_res7__224] ^ p18_array_index_2047004 ^ p18_array_index_2047084 ^ p18_array_index_2047055 ^ p18_array_index_2047023 ^ p18_literal_2043914[p18_array_index_2047008] ^ p18_literal_2043912[p18_array_index_2047009] ^ p18_literal_2043910[p18_array_index_2047026] ^ p18_array_index_2047011;
  assign p19_array_index_2047258_comb = p18_literal_2043918[p18_res7__232];
  assign p19_array_index_2047259_comb = p18_literal_2043920[p18_res7__230];
  assign p19_res7__242_comb = p18_literal_2043910[p19_res7__240_comb] ^ p18_literal_2043912[p19_res7__238_comb] ^ p18_literal_2043914[p19_res7__236_comb] ^ p18_literal_2043916[p18_res7__234] ^ p19_array_index_2047258_comb ^ p19_array_index_2047259_comb ^ p18_res7__228 ^ p18_literal_2043923[p18_res7__226] ^ p18_res7__224 ^ p18_array_index_2047097 ^ p18_array_index_2047069 ^ p18_array_index_2047040 ^ p18_literal_2043914[p18_array_index_2047007] ^ p18_literal_2043912[p18_array_index_2047008] ^ p18_literal_2043910[p18_array_index_2047009] ^ p18_array_index_2047026;
  assign p19_array_index_2047270_comb = p18_literal_2043920[p18_res7__232];
  assign p19_res7__244_comb = p18_literal_2043910[p19_res7__242_comb] ^ p18_literal_2043912[p19_res7__240_comb] ^ p18_literal_2043914[p19_res7__238_comb] ^ p18_literal_2043916[p19_res7__236_comb] ^ p18_literal_2043918[p18_res7__234] ^ p19_array_index_2047270_comb ^ p18_res7__230 ^ p18_literal_2043923[p18_res7__228] ^ p18_res7__226 ^ p19_array_index_2047224_comb ^ p18_array_index_2047083 ^ p18_array_index_2047054 ^ p18_array_index_2047022 ^ p18_literal_2043912[p18_array_index_2047007] ^ p18_literal_2043910[p18_array_index_2047008] ^ p18_array_index_2047009;
  assign p19_array_index_2047280_comb = p18_literal_2043920[p18_res7__234];
  assign p19_res7__246_comb = p18_literal_2043910[p19_res7__244_comb] ^ p18_literal_2043912[p19_res7__242_comb] ^ p18_literal_2043914[p19_res7__240_comb] ^ p18_literal_2043916[p19_res7__238_comb] ^ p18_literal_2043918[p19_res7__236_comb] ^ p19_array_index_2047280_comb ^ p18_res7__232 ^ p18_literal_2043923[p18_res7__230] ^ p18_res7__228 ^ p19_array_index_2047236_comb ^ p18_array_index_2047096 ^ p18_array_index_2047068 ^ p18_array_index_2047039 ^ p18_literal_2043912[p18_array_index_2047006] ^ p18_literal_2043910[p18_array_index_2047007] ^ p18_array_index_2047008;
  assign p19_res7__248_comb = p18_literal_2043910[p19_res7__246_comb] ^ p18_literal_2043912[p19_res7__244_comb] ^ p18_literal_2043914[p19_res7__242_comb] ^ p18_literal_2043916[p19_res7__240_comb] ^ p18_literal_2043918[p19_res7__238_comb] ^ p18_literal_2043920[p19_res7__236_comb] ^ p18_res7__234 ^ p18_literal_2043923[p18_res7__232] ^ p18_res7__230 ^ p19_array_index_2047248_comb ^ p19_array_index_2047223_comb ^ p18_array_index_2047082 ^ p18_array_index_2047053 ^ p18_array_index_2047021 ^ p18_literal_2043910[p18_array_index_2047006] ^ p18_array_index_2047007;

  // Registers for pipe stage 19:
  reg [127:0] p19_encoded;
  reg [127:0] p19_bit_slice_2043893;
  reg [127:0] p19_bit_slice_2044018;
  reg [127:0] p19_xor_2046544;
  reg [127:0] p19_k3;
  reg [7:0] p19_array_index_2047004;
  reg [7:0] p19_array_index_2047005;
  reg [7:0] p19_array_index_2047006;
  reg [7:0] p19_array_index_2047020;
  reg [7:0] p19_res7__224;
  reg [7:0] p19_array_index_2047037;
  reg [7:0] p19_array_index_2047038;
  reg [7:0] p19_res7__226;
  reg [7:0] p19_array_index_2047052;
  reg [7:0] p19_res7__228;
  reg [7:0] p19_array_index_2047066;
  reg [7:0] p19_array_index_2047067;
  reg [7:0] p19_res7__230;
  reg [7:0] p19_array_index_2047081;
  reg [7:0] p19_res7__232;
  reg [7:0] p19_array_index_2047094;
  reg [7:0] p19_array_index_2047095;
  reg [7:0] p19_res7__234;
  reg [7:0] p19_array_index_2047222;
  reg [7:0] p19_res7__236;
  reg [7:0] p19_array_index_2047234;
  reg [7:0] p19_array_index_2047235;
  reg [7:0] p19_res7__238;
  reg [7:0] p19_array_index_2047247;
  reg [7:0] p19_res7__240;
  reg [7:0] p19_array_index_2047258;
  reg [7:0] p19_array_index_2047259;
  reg [7:0] p19_res7__242;
  reg [7:0] p19_array_index_2047270;
  reg [7:0] p19_res7__244;
  reg [7:0] p19_array_index_2047280;
  reg [7:0] p19_res7__246;
  reg [7:0] p19_res7__248;
  reg [7:0] p20_literal_2043896[256];
  reg [7:0] p20_literal_2043910[256];
  reg [7:0] p20_literal_2043912[256];
  reg [7:0] p20_literal_2043914[256];
  reg [7:0] p20_literal_2043916[256];
  reg [7:0] p20_literal_2043918[256];
  reg [7:0] p20_literal_2043920[256];
  reg [7:0] p20_literal_2043923[256];
  reg [7:0] p97_literal_2058836[256];
  always_ff @ (posedge clk) begin
    p19_encoded <= p18_encoded;
    p19_bit_slice_2043893 <= p18_bit_slice_2043893;
    p19_bit_slice_2044018 <= p18_bit_slice_2044018;
    p19_xor_2046544 <= p18_xor_2046544;
    p19_k3 <= p18_k3;
    p19_array_index_2047004 <= p18_array_index_2047004;
    p19_array_index_2047005 <= p18_array_index_2047005;
    p19_array_index_2047006 <= p18_array_index_2047006;
    p19_array_index_2047020 <= p18_array_index_2047020;
    p19_res7__224 <= p18_res7__224;
    p19_array_index_2047037 <= p18_array_index_2047037;
    p19_array_index_2047038 <= p18_array_index_2047038;
    p19_res7__226 <= p18_res7__226;
    p19_array_index_2047052 <= p18_array_index_2047052;
    p19_res7__228 <= p18_res7__228;
    p19_array_index_2047066 <= p18_array_index_2047066;
    p19_array_index_2047067 <= p18_array_index_2047067;
    p19_res7__230 <= p18_res7__230;
    p19_array_index_2047081 <= p18_array_index_2047081;
    p19_res7__232 <= p18_res7__232;
    p19_array_index_2047094 <= p18_array_index_2047094;
    p19_array_index_2047095 <= p18_array_index_2047095;
    p19_res7__234 <= p18_res7__234;
    p19_array_index_2047222 <= p19_array_index_2047222_comb;
    p19_res7__236 <= p19_res7__236_comb;
    p19_array_index_2047234 <= p19_array_index_2047234_comb;
    p19_array_index_2047235 <= p19_array_index_2047235_comb;
    p19_res7__238 <= p19_res7__238_comb;
    p19_array_index_2047247 <= p19_array_index_2047247_comb;
    p19_res7__240 <= p19_res7__240_comb;
    p19_array_index_2047258 <= p19_array_index_2047258_comb;
    p19_array_index_2047259 <= p19_array_index_2047259_comb;
    p19_res7__242 <= p19_res7__242_comb;
    p19_array_index_2047270 <= p19_array_index_2047270_comb;
    p19_res7__244 <= p19_res7__244_comb;
    p19_array_index_2047280 <= p19_array_index_2047280_comb;
    p19_res7__246 <= p19_res7__246_comb;
    p19_res7__248 <= p19_res7__248_comb;
    p20_literal_2043896 <= p19_literal_2043896;
    p20_literal_2043910 <= p19_literal_2043910;
    p20_literal_2043912 <= p19_literal_2043912;
    p20_literal_2043914 <= p19_literal_2043914;
    p20_literal_2043916 <= p19_literal_2043916;
    p20_literal_2043918 <= p19_literal_2043918;
    p20_literal_2043920 <= p19_literal_2043920;
    p20_literal_2043923 <= p19_literal_2043923;
    p97_literal_2058836 <= p96_literal_2058836;
  end

  // ===== Pipe stage 20:
  wire [7:0] p20_res7__250_comb;
  wire [7:0] p20_res7__252_comb;
  wire [7:0] p20_res7__254_comb;
  wire [127:0] p20_res__7_comb;
  wire [127:0] p20_k2_comb;
  wire [127:0] p20_addedKey__40_comb;
  wire [7:0] p20_array_index_2047428_comb;
  wire [7:0] p20_array_index_2047429_comb;
  wire [7:0] p20_array_index_2047430_comb;
  wire [7:0] p20_array_index_2047431_comb;
  wire [7:0] p20_array_index_2047432_comb;
  wire [7:0] p20_array_index_2047433_comb;
  wire [7:0] p20_array_index_2047435_comb;
  wire [7:0] p20_array_index_2047437_comb;
  wire [7:0] p20_array_index_2047438_comb;
  wire [7:0] p20_array_index_2047439_comb;
  wire [7:0] p20_array_index_2047440_comb;
  wire [7:0] p20_array_index_2047441_comb;
  wire [7:0] p20_array_index_2047442_comb;
  wire [7:0] p20_array_index_2047444_comb;
  wire [7:0] p20_array_index_2047445_comb;
  wire [7:0] p20_array_index_2047446_comb;
  wire [7:0] p20_array_index_2047447_comb;
  wire [7:0] p20_array_index_2047448_comb;
  wire [7:0] p20_array_index_2047449_comb;
  wire [7:0] p20_array_index_2047450_comb;
  wire [7:0] p20_array_index_2047452_comb;
  wire [7:0] p20_res7__256_comb;
  wire [7:0] p20_array_index_2047461_comb;
  wire [7:0] p20_array_index_2047462_comb;
  wire [7:0] p20_array_index_2047463_comb;
  wire [7:0] p20_array_index_2047464_comb;
  wire [7:0] p20_array_index_2047465_comb;
  wire [7:0] p20_array_index_2047466_comb;
  wire [7:0] p20_res7__258_comb;
  wire [7:0] p20_array_index_2047476_comb;
  wire [7:0] p20_array_index_2047477_comb;
  wire [7:0] p20_array_index_2047478_comb;
  wire [7:0] p20_array_index_2047479_comb;
  wire [7:0] p20_array_index_2047480_comb;
  wire [7:0] p20_res7__260_comb;
  assign p20_res7__250_comb = p19_literal_2043910[p19_res7__248] ^ p19_literal_2043912[p19_res7__246] ^ p19_literal_2043914[p19_res7__244] ^ p19_literal_2043916[p19_res7__242] ^ p19_literal_2043918[p19_res7__240] ^ p19_literal_2043920[p19_res7__238] ^ p19_res7__236 ^ p19_literal_2043923[p19_res7__234] ^ p19_res7__232 ^ p19_array_index_2047259 ^ p19_array_index_2047235 ^ p19_array_index_2047095 ^ p19_array_index_2047067 ^ p19_array_index_2047038 ^ p19_literal_2043910[p19_array_index_2047005] ^ p19_array_index_2047006;
  assign p20_res7__252_comb = p19_literal_2043910[p20_res7__250_comb] ^ p19_literal_2043912[p19_res7__248] ^ p19_literal_2043914[p19_res7__246] ^ p19_literal_2043916[p19_res7__244] ^ p19_literal_2043918[p19_res7__242] ^ p19_literal_2043920[p19_res7__240] ^ p19_res7__238 ^ p19_literal_2043923[p19_res7__236] ^ p19_res7__234 ^ p19_array_index_2047270 ^ p19_array_index_2047247 ^ p19_array_index_2047222 ^ p19_array_index_2047081 ^ p19_array_index_2047052 ^ p19_array_index_2047020 ^ p19_array_index_2047005;
  assign p20_res7__254_comb = p19_literal_2043910[p20_res7__252_comb] ^ p19_literal_2043912[p20_res7__250_comb] ^ p19_literal_2043914[p19_res7__248] ^ p19_literal_2043916[p19_res7__246] ^ p19_literal_2043918[p19_res7__244] ^ p19_literal_2043920[p19_res7__242] ^ p19_res7__240 ^ p19_literal_2043923[p19_res7__238] ^ p19_res7__236 ^ p19_array_index_2047280 ^ p19_array_index_2047258 ^ p19_array_index_2047234 ^ p19_array_index_2047094 ^ p19_array_index_2047066 ^ p19_array_index_2047037 ^ p19_array_index_2047004;
  assign p20_res__7_comb = {p20_res7__254_comb, p20_res7__252_comb, p20_res7__250_comb, p19_res7__248, p19_res7__246, p19_res7__244, p19_res7__242, p19_res7__240, p19_res7__238, p19_res7__236, p19_res7__234, p19_res7__232, p19_res7__230, p19_res7__228, p19_res7__226, p19_res7__224};
  assign p20_k2_comb = p20_res__7_comb ^ p19_xor_2046544;
  assign p20_addedKey__40_comb = p20_k2_comb ^ 128'h98fb_4064_8a4d_2c31_f0dc_1c90_fa2e_be09;
  assign p20_array_index_2047428_comb = p19_literal_2043896[p20_addedKey__40_comb[127:120]];
  assign p20_array_index_2047429_comb = p19_literal_2043896[p20_addedKey__40_comb[119:112]];
  assign p20_array_index_2047430_comb = p19_literal_2043896[p20_addedKey__40_comb[111:104]];
  assign p20_array_index_2047431_comb = p19_literal_2043896[p20_addedKey__40_comb[103:96]];
  assign p20_array_index_2047432_comb = p19_literal_2043896[p20_addedKey__40_comb[95:88]];
  assign p20_array_index_2047433_comb = p19_literal_2043896[p20_addedKey__40_comb[87:80]];
  assign p20_array_index_2047435_comb = p19_literal_2043896[p20_addedKey__40_comb[71:64]];
  assign p20_array_index_2047437_comb = p19_literal_2043896[p20_addedKey__40_comb[55:48]];
  assign p20_array_index_2047438_comb = p19_literal_2043896[p20_addedKey__40_comb[47:40]];
  assign p20_array_index_2047439_comb = p19_literal_2043896[p20_addedKey__40_comb[39:32]];
  assign p20_array_index_2047440_comb = p19_literal_2043896[p20_addedKey__40_comb[31:24]];
  assign p20_array_index_2047441_comb = p19_literal_2043896[p20_addedKey__40_comb[23:16]];
  assign p20_array_index_2047442_comb = p19_literal_2043896[p20_addedKey__40_comb[15:8]];
  assign p20_array_index_2047444_comb = p19_literal_2043910[p20_array_index_2047428_comb];
  assign p20_array_index_2047445_comb = p19_literal_2043912[p20_array_index_2047429_comb];
  assign p20_array_index_2047446_comb = p19_literal_2043914[p20_array_index_2047430_comb];
  assign p20_array_index_2047447_comb = p19_literal_2043916[p20_array_index_2047431_comb];
  assign p20_array_index_2047448_comb = p19_literal_2043918[p20_array_index_2047432_comb];
  assign p20_array_index_2047449_comb = p19_literal_2043920[p20_array_index_2047433_comb];
  assign p20_array_index_2047450_comb = p19_literal_2043896[p20_addedKey__40_comb[79:72]];
  assign p20_array_index_2047452_comb = p19_literal_2043896[p20_addedKey__40_comb[63:56]];
  assign p20_res7__256_comb = p20_array_index_2047444_comb ^ p20_array_index_2047445_comb ^ p20_array_index_2047446_comb ^ p20_array_index_2047447_comb ^ p20_array_index_2047448_comb ^ p20_array_index_2047449_comb ^ p20_array_index_2047450_comb ^ p19_literal_2043923[p20_array_index_2047435_comb] ^ p20_array_index_2047452_comb ^ p19_literal_2043920[p20_array_index_2047437_comb] ^ p19_literal_2043918[p20_array_index_2047438_comb] ^ p19_literal_2043916[p20_array_index_2047439_comb] ^ p19_literal_2043914[p20_array_index_2047440_comb] ^ p19_literal_2043912[p20_array_index_2047441_comb] ^ p19_literal_2043910[p20_array_index_2047442_comb] ^ p19_literal_2043896[p20_addedKey__40_comb[7:0]];
  assign p20_array_index_2047461_comb = p19_literal_2043910[p20_res7__256_comb];
  assign p20_array_index_2047462_comb = p19_literal_2043912[p20_array_index_2047428_comb];
  assign p20_array_index_2047463_comb = p19_literal_2043914[p20_array_index_2047429_comb];
  assign p20_array_index_2047464_comb = p19_literal_2043916[p20_array_index_2047430_comb];
  assign p20_array_index_2047465_comb = p19_literal_2043918[p20_array_index_2047431_comb];
  assign p20_array_index_2047466_comb = p19_literal_2043920[p20_array_index_2047432_comb];
  assign p20_res7__258_comb = p20_array_index_2047461_comb ^ p20_array_index_2047462_comb ^ p20_array_index_2047463_comb ^ p20_array_index_2047464_comb ^ p20_array_index_2047465_comb ^ p20_array_index_2047466_comb ^ p20_array_index_2047433_comb ^ p19_literal_2043923[p20_array_index_2047450_comb] ^ p20_array_index_2047435_comb ^ p19_literal_2043920[p20_array_index_2047452_comb] ^ p19_literal_2043918[p20_array_index_2047437_comb] ^ p19_literal_2043916[p20_array_index_2047438_comb] ^ p19_literal_2043914[p20_array_index_2047439_comb] ^ p19_literal_2043912[p20_array_index_2047440_comb] ^ p19_literal_2043910[p20_array_index_2047441_comb] ^ p20_array_index_2047442_comb;
  assign p20_array_index_2047476_comb = p19_literal_2043912[p20_res7__256_comb];
  assign p20_array_index_2047477_comb = p19_literal_2043914[p20_array_index_2047428_comb];
  assign p20_array_index_2047478_comb = p19_literal_2043916[p20_array_index_2047429_comb];
  assign p20_array_index_2047479_comb = p19_literal_2043918[p20_array_index_2047430_comb];
  assign p20_array_index_2047480_comb = p19_literal_2043920[p20_array_index_2047431_comb];
  assign p20_res7__260_comb = p19_literal_2043910[p20_res7__258_comb] ^ p20_array_index_2047476_comb ^ p20_array_index_2047477_comb ^ p20_array_index_2047478_comb ^ p20_array_index_2047479_comb ^ p20_array_index_2047480_comb ^ p20_array_index_2047432_comb ^ p19_literal_2043923[p20_array_index_2047433_comb] ^ p20_array_index_2047450_comb ^ p19_literal_2043920[p20_array_index_2047435_comb] ^ p19_literal_2043918[p20_array_index_2047452_comb] ^ p19_literal_2043916[p20_array_index_2047437_comb] ^ p19_literal_2043914[p20_array_index_2047438_comb] ^ p19_literal_2043912[p20_array_index_2047439_comb] ^ p19_literal_2043910[p20_array_index_2047440_comb] ^ p20_array_index_2047441_comb;

  // Registers for pipe stage 20:
  reg [127:0] p20_encoded;
  reg [127:0] p20_bit_slice_2043893;
  reg [127:0] p20_bit_slice_2044018;
  reg [127:0] p20_k3;
  reg [127:0] p20_k2;
  reg [7:0] p20_array_index_2047428;
  reg [7:0] p20_array_index_2047429;
  reg [7:0] p20_array_index_2047430;
  reg [7:0] p20_array_index_2047431;
  reg [7:0] p20_array_index_2047432;
  reg [7:0] p20_array_index_2047433;
  reg [7:0] p20_array_index_2047435;
  reg [7:0] p20_array_index_2047437;
  reg [7:0] p20_array_index_2047438;
  reg [7:0] p20_array_index_2047439;
  reg [7:0] p20_array_index_2047440;
  reg [7:0] p20_array_index_2047444;
  reg [7:0] p20_array_index_2047445;
  reg [7:0] p20_array_index_2047446;
  reg [7:0] p20_array_index_2047447;
  reg [7:0] p20_array_index_2047448;
  reg [7:0] p20_array_index_2047449;
  reg [7:0] p20_array_index_2047450;
  reg [7:0] p20_array_index_2047452;
  reg [7:0] p20_res7__256;
  reg [7:0] p20_array_index_2047461;
  reg [7:0] p20_array_index_2047462;
  reg [7:0] p20_array_index_2047463;
  reg [7:0] p20_array_index_2047464;
  reg [7:0] p20_array_index_2047465;
  reg [7:0] p20_array_index_2047466;
  reg [7:0] p20_res7__258;
  reg [7:0] p20_array_index_2047476;
  reg [7:0] p20_array_index_2047477;
  reg [7:0] p20_array_index_2047478;
  reg [7:0] p20_array_index_2047479;
  reg [7:0] p20_array_index_2047480;
  reg [7:0] p20_res7__260;
  reg [7:0] p21_literal_2043896[256];
  reg [7:0] p21_literal_2043910[256];
  reg [7:0] p21_literal_2043912[256];
  reg [7:0] p21_literal_2043914[256];
  reg [7:0] p21_literal_2043916[256];
  reg [7:0] p21_literal_2043918[256];
  reg [7:0] p21_literal_2043920[256];
  reg [7:0] p21_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p20_encoded <= p19_encoded;
    p20_bit_slice_2043893 <= p19_bit_slice_2043893;
    p20_bit_slice_2044018 <= p19_bit_slice_2044018;
    p20_k3 <= p19_k3;
    p20_k2 <= p20_k2_comb;
    p20_array_index_2047428 <= p20_array_index_2047428_comb;
    p20_array_index_2047429 <= p20_array_index_2047429_comb;
    p20_array_index_2047430 <= p20_array_index_2047430_comb;
    p20_array_index_2047431 <= p20_array_index_2047431_comb;
    p20_array_index_2047432 <= p20_array_index_2047432_comb;
    p20_array_index_2047433 <= p20_array_index_2047433_comb;
    p20_array_index_2047435 <= p20_array_index_2047435_comb;
    p20_array_index_2047437 <= p20_array_index_2047437_comb;
    p20_array_index_2047438 <= p20_array_index_2047438_comb;
    p20_array_index_2047439 <= p20_array_index_2047439_comb;
    p20_array_index_2047440 <= p20_array_index_2047440_comb;
    p20_array_index_2047444 <= p20_array_index_2047444_comb;
    p20_array_index_2047445 <= p20_array_index_2047445_comb;
    p20_array_index_2047446 <= p20_array_index_2047446_comb;
    p20_array_index_2047447 <= p20_array_index_2047447_comb;
    p20_array_index_2047448 <= p20_array_index_2047448_comb;
    p20_array_index_2047449 <= p20_array_index_2047449_comb;
    p20_array_index_2047450 <= p20_array_index_2047450_comb;
    p20_array_index_2047452 <= p20_array_index_2047452_comb;
    p20_res7__256 <= p20_res7__256_comb;
    p20_array_index_2047461 <= p20_array_index_2047461_comb;
    p20_array_index_2047462 <= p20_array_index_2047462_comb;
    p20_array_index_2047463 <= p20_array_index_2047463_comb;
    p20_array_index_2047464 <= p20_array_index_2047464_comb;
    p20_array_index_2047465 <= p20_array_index_2047465_comb;
    p20_array_index_2047466 <= p20_array_index_2047466_comb;
    p20_res7__258 <= p20_res7__258_comb;
    p20_array_index_2047476 <= p20_array_index_2047476_comb;
    p20_array_index_2047477 <= p20_array_index_2047477_comb;
    p20_array_index_2047478 <= p20_array_index_2047478_comb;
    p20_array_index_2047479 <= p20_array_index_2047479_comb;
    p20_array_index_2047480 <= p20_array_index_2047480_comb;
    p20_res7__260 <= p20_res7__260_comb;
    p21_literal_2043896 <= p20_literal_2043896;
    p21_literal_2043910 <= p20_literal_2043910;
    p21_literal_2043912 <= p20_literal_2043912;
    p21_literal_2043914 <= p20_literal_2043914;
    p21_literal_2043916 <= p20_literal_2043916;
    p21_literal_2043918 <= p20_literal_2043918;
    p21_literal_2043920 <= p20_literal_2043920;
    p21_literal_2043923 <= p20_literal_2043923;
  end

  // ===== Pipe stage 21:
  wire [7:0] p21_array_index_2047582_comb;
  wire [7:0] p21_array_index_2047583_comb;
  wire [7:0] p21_array_index_2047584_comb;
  wire [7:0] p21_array_index_2047585_comb;
  wire [7:0] p21_array_index_2047586_comb;
  wire [7:0] p21_res7__262_comb;
  wire [7:0] p21_array_index_2047597_comb;
  wire [7:0] p21_array_index_2047598_comb;
  wire [7:0] p21_array_index_2047599_comb;
  wire [7:0] p21_array_index_2047600_comb;
  wire [7:0] p21_res7__264_comb;
  wire [7:0] p21_array_index_2047610_comb;
  wire [7:0] p21_array_index_2047611_comb;
  wire [7:0] p21_array_index_2047612_comb;
  wire [7:0] p21_array_index_2047613_comb;
  wire [7:0] p21_res7__266_comb;
  wire [7:0] p21_array_index_2047624_comb;
  wire [7:0] p21_array_index_2047625_comb;
  wire [7:0] p21_array_index_2047626_comb;
  wire [7:0] p21_res7__268_comb;
  wire [7:0] p21_array_index_2047636_comb;
  wire [7:0] p21_array_index_2047637_comb;
  wire [7:0] p21_array_index_2047638_comb;
  wire [7:0] p21_res7__270_comb;
  wire [7:0] p21_array_index_2047649_comb;
  wire [7:0] p21_array_index_2047650_comb;
  wire [7:0] p21_res7__272_comb;
  wire [7:0] p21_array_index_2047660_comb;
  wire [7:0] p21_array_index_2047661_comb;
  wire [7:0] p21_res7__274_comb;
  assign p21_array_index_2047582_comb = p20_literal_2043912[p20_res7__258];
  assign p21_array_index_2047583_comb = p20_literal_2043914[p20_res7__256];
  assign p21_array_index_2047584_comb = p20_literal_2043916[p20_array_index_2047428];
  assign p21_array_index_2047585_comb = p20_literal_2043918[p20_array_index_2047429];
  assign p21_array_index_2047586_comb = p20_literal_2043920[p20_array_index_2047430];
  assign p21_res7__262_comb = p20_literal_2043910[p20_res7__260] ^ p21_array_index_2047582_comb ^ p21_array_index_2047583_comb ^ p21_array_index_2047584_comb ^ p21_array_index_2047585_comb ^ p21_array_index_2047586_comb ^ p20_array_index_2047431 ^ p20_literal_2043923[p20_array_index_2047432] ^ p20_array_index_2047433 ^ p20_literal_2043920[p20_array_index_2047450] ^ p20_literal_2043918[p20_array_index_2047435] ^ p20_literal_2043916[p20_array_index_2047452] ^ p20_literal_2043914[p20_array_index_2047437] ^ p20_literal_2043912[p20_array_index_2047438] ^ p20_literal_2043910[p20_array_index_2047439] ^ p20_array_index_2047440;
  assign p21_array_index_2047597_comb = p20_literal_2043914[p20_res7__258];
  assign p21_array_index_2047598_comb = p20_literal_2043916[p20_res7__256];
  assign p21_array_index_2047599_comb = p20_literal_2043918[p20_array_index_2047428];
  assign p21_array_index_2047600_comb = p20_literal_2043920[p20_array_index_2047429];
  assign p21_res7__264_comb = p20_literal_2043910[p21_res7__262_comb] ^ p20_literal_2043912[p20_res7__260] ^ p21_array_index_2047597_comb ^ p21_array_index_2047598_comb ^ p21_array_index_2047599_comb ^ p21_array_index_2047600_comb ^ p20_array_index_2047430 ^ p20_literal_2043923[p20_array_index_2047431] ^ p20_array_index_2047432 ^ p20_array_index_2047449 ^ p20_literal_2043918[p20_array_index_2047450] ^ p20_literal_2043916[p20_array_index_2047435] ^ p20_literal_2043914[p20_array_index_2047452] ^ p20_literal_2043912[p20_array_index_2047437] ^ p20_literal_2043910[p20_array_index_2047438] ^ p20_array_index_2047439;
  assign p21_array_index_2047610_comb = p20_literal_2043914[p20_res7__260];
  assign p21_array_index_2047611_comb = p20_literal_2043916[p20_res7__258];
  assign p21_array_index_2047612_comb = p20_literal_2043918[p20_res7__256];
  assign p21_array_index_2047613_comb = p20_literal_2043920[p20_array_index_2047428];
  assign p21_res7__266_comb = p20_literal_2043910[p21_res7__264_comb] ^ p20_literal_2043912[p21_res7__262_comb] ^ p21_array_index_2047610_comb ^ p21_array_index_2047611_comb ^ p21_array_index_2047612_comb ^ p21_array_index_2047613_comb ^ p20_array_index_2047429 ^ p20_literal_2043923[p20_array_index_2047430] ^ p20_array_index_2047431 ^ p20_array_index_2047466 ^ p20_literal_2043918[p20_array_index_2047433] ^ p20_literal_2043916[p20_array_index_2047450] ^ p20_literal_2043914[p20_array_index_2047435] ^ p20_literal_2043912[p20_array_index_2047452] ^ p20_literal_2043910[p20_array_index_2047437] ^ p20_array_index_2047438;
  assign p21_array_index_2047624_comb = p20_literal_2043916[p20_res7__260];
  assign p21_array_index_2047625_comb = p20_literal_2043918[p20_res7__258];
  assign p21_array_index_2047626_comb = p20_literal_2043920[p20_res7__256];
  assign p21_res7__268_comb = p20_literal_2043910[p21_res7__266_comb] ^ p20_literal_2043912[p21_res7__264_comb] ^ p20_literal_2043914[p21_res7__262_comb] ^ p21_array_index_2047624_comb ^ p21_array_index_2047625_comb ^ p21_array_index_2047626_comb ^ p20_array_index_2047428 ^ p20_literal_2043923[p20_array_index_2047429] ^ p20_array_index_2047430 ^ p20_array_index_2047480 ^ p20_array_index_2047448 ^ p20_literal_2043916[p20_array_index_2047433] ^ p20_literal_2043914[p20_array_index_2047450] ^ p20_literal_2043912[p20_array_index_2047435] ^ p20_literal_2043910[p20_array_index_2047452] ^ p20_array_index_2047437;
  assign p21_array_index_2047636_comb = p20_literal_2043916[p21_res7__262_comb];
  assign p21_array_index_2047637_comb = p20_literal_2043918[p20_res7__260];
  assign p21_array_index_2047638_comb = p20_literal_2043920[p20_res7__258];
  assign p21_res7__270_comb = p20_literal_2043910[p21_res7__268_comb] ^ p20_literal_2043912[p21_res7__266_comb] ^ p20_literal_2043914[p21_res7__264_comb] ^ p21_array_index_2047636_comb ^ p21_array_index_2047637_comb ^ p21_array_index_2047638_comb ^ p20_res7__256 ^ p20_literal_2043923[p20_array_index_2047428] ^ p20_array_index_2047429 ^ p21_array_index_2047586_comb ^ p20_array_index_2047465 ^ p20_literal_2043916[p20_array_index_2047432] ^ p20_literal_2043914[p20_array_index_2047433] ^ p20_literal_2043912[p20_array_index_2047450] ^ p20_literal_2043910[p20_array_index_2047435] ^ p20_array_index_2047452;
  assign p21_array_index_2047649_comb = p20_literal_2043918[p21_res7__262_comb];
  assign p21_array_index_2047650_comb = p20_literal_2043920[p20_res7__260];
  assign p21_res7__272_comb = p20_literal_2043910[p21_res7__270_comb] ^ p20_literal_2043912[p21_res7__268_comb] ^ p20_literal_2043914[p21_res7__266_comb] ^ p20_literal_2043916[p21_res7__264_comb] ^ p21_array_index_2047649_comb ^ p21_array_index_2047650_comb ^ p20_res7__258 ^ p20_literal_2043923[p20_res7__256] ^ p20_array_index_2047428 ^ p21_array_index_2047600_comb ^ p20_array_index_2047479 ^ p20_array_index_2047447 ^ p20_literal_2043914[p20_array_index_2047432] ^ p20_literal_2043912[p20_array_index_2047433] ^ p20_literal_2043910[p20_array_index_2047450] ^ p20_array_index_2047435;
  assign p21_array_index_2047660_comb = p20_literal_2043918[p21_res7__264_comb];
  assign p21_array_index_2047661_comb = p20_literal_2043920[p21_res7__262_comb];
  assign p21_res7__274_comb = p20_literal_2043910[p21_res7__272_comb] ^ p20_literal_2043912[p21_res7__270_comb] ^ p20_literal_2043914[p21_res7__268_comb] ^ p20_literal_2043916[p21_res7__266_comb] ^ p21_array_index_2047660_comb ^ p21_array_index_2047661_comb ^ p20_res7__260 ^ p20_literal_2043923[p20_res7__258] ^ p20_res7__256 ^ p21_array_index_2047613_comb ^ p21_array_index_2047585_comb ^ p20_array_index_2047464 ^ p20_literal_2043914[p20_array_index_2047431] ^ p20_literal_2043912[p20_array_index_2047432] ^ p20_literal_2043910[p20_array_index_2047433] ^ p20_array_index_2047450;

  // Registers for pipe stage 21:
  reg [127:0] p21_encoded;
  reg [127:0] p21_bit_slice_2043893;
  reg [127:0] p21_bit_slice_2044018;
  reg [127:0] p21_k3;
  reg [127:0] p21_k2;
  reg [7:0] p21_array_index_2047428;
  reg [7:0] p21_array_index_2047429;
  reg [7:0] p21_array_index_2047430;
  reg [7:0] p21_array_index_2047431;
  reg [7:0] p21_array_index_2047432;
  reg [7:0] p21_array_index_2047433;
  reg [7:0] p21_array_index_2047444;
  reg [7:0] p21_array_index_2047445;
  reg [7:0] p21_array_index_2047446;
  reg [7:0] p21_res7__256;
  reg [7:0] p21_array_index_2047461;
  reg [7:0] p21_array_index_2047462;
  reg [7:0] p21_array_index_2047463;
  reg [7:0] p21_res7__258;
  reg [7:0] p21_array_index_2047476;
  reg [7:0] p21_array_index_2047477;
  reg [7:0] p21_array_index_2047478;
  reg [7:0] p21_res7__260;
  reg [7:0] p21_array_index_2047582;
  reg [7:0] p21_array_index_2047583;
  reg [7:0] p21_array_index_2047584;
  reg [7:0] p21_res7__262;
  reg [7:0] p21_array_index_2047597;
  reg [7:0] p21_array_index_2047598;
  reg [7:0] p21_array_index_2047599;
  reg [7:0] p21_res7__264;
  reg [7:0] p21_array_index_2047610;
  reg [7:0] p21_array_index_2047611;
  reg [7:0] p21_array_index_2047612;
  reg [7:0] p21_res7__266;
  reg [7:0] p21_array_index_2047624;
  reg [7:0] p21_array_index_2047625;
  reg [7:0] p21_array_index_2047626;
  reg [7:0] p21_res7__268;
  reg [7:0] p21_array_index_2047636;
  reg [7:0] p21_array_index_2047637;
  reg [7:0] p21_array_index_2047638;
  reg [7:0] p21_res7__270;
  reg [7:0] p21_array_index_2047649;
  reg [7:0] p21_array_index_2047650;
  reg [7:0] p21_res7__272;
  reg [7:0] p21_array_index_2047660;
  reg [7:0] p21_array_index_2047661;
  reg [7:0] p21_res7__274;
  reg [7:0] p22_literal_2043896[256];
  reg [7:0] p22_literal_2043910[256];
  reg [7:0] p22_literal_2043912[256];
  reg [7:0] p22_literal_2043914[256];
  reg [7:0] p22_literal_2043916[256];
  reg [7:0] p22_literal_2043918[256];
  reg [7:0] p22_literal_2043920[256];
  reg [7:0] p22_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p21_encoded <= p20_encoded;
    p21_bit_slice_2043893 <= p20_bit_slice_2043893;
    p21_bit_slice_2044018 <= p20_bit_slice_2044018;
    p21_k3 <= p20_k3;
    p21_k2 <= p20_k2;
    p21_array_index_2047428 <= p20_array_index_2047428;
    p21_array_index_2047429 <= p20_array_index_2047429;
    p21_array_index_2047430 <= p20_array_index_2047430;
    p21_array_index_2047431 <= p20_array_index_2047431;
    p21_array_index_2047432 <= p20_array_index_2047432;
    p21_array_index_2047433 <= p20_array_index_2047433;
    p21_array_index_2047444 <= p20_array_index_2047444;
    p21_array_index_2047445 <= p20_array_index_2047445;
    p21_array_index_2047446 <= p20_array_index_2047446;
    p21_res7__256 <= p20_res7__256;
    p21_array_index_2047461 <= p20_array_index_2047461;
    p21_array_index_2047462 <= p20_array_index_2047462;
    p21_array_index_2047463 <= p20_array_index_2047463;
    p21_res7__258 <= p20_res7__258;
    p21_array_index_2047476 <= p20_array_index_2047476;
    p21_array_index_2047477 <= p20_array_index_2047477;
    p21_array_index_2047478 <= p20_array_index_2047478;
    p21_res7__260 <= p20_res7__260;
    p21_array_index_2047582 <= p21_array_index_2047582_comb;
    p21_array_index_2047583 <= p21_array_index_2047583_comb;
    p21_array_index_2047584 <= p21_array_index_2047584_comb;
    p21_res7__262 <= p21_res7__262_comb;
    p21_array_index_2047597 <= p21_array_index_2047597_comb;
    p21_array_index_2047598 <= p21_array_index_2047598_comb;
    p21_array_index_2047599 <= p21_array_index_2047599_comb;
    p21_res7__264 <= p21_res7__264_comb;
    p21_array_index_2047610 <= p21_array_index_2047610_comb;
    p21_array_index_2047611 <= p21_array_index_2047611_comb;
    p21_array_index_2047612 <= p21_array_index_2047612_comb;
    p21_res7__266 <= p21_res7__266_comb;
    p21_array_index_2047624 <= p21_array_index_2047624_comb;
    p21_array_index_2047625 <= p21_array_index_2047625_comb;
    p21_array_index_2047626 <= p21_array_index_2047626_comb;
    p21_res7__268 <= p21_res7__268_comb;
    p21_array_index_2047636 <= p21_array_index_2047636_comb;
    p21_array_index_2047637 <= p21_array_index_2047637_comb;
    p21_array_index_2047638 <= p21_array_index_2047638_comb;
    p21_res7__270 <= p21_res7__270_comb;
    p21_array_index_2047649 <= p21_array_index_2047649_comb;
    p21_array_index_2047650 <= p21_array_index_2047650_comb;
    p21_res7__272 <= p21_res7__272_comb;
    p21_array_index_2047660 <= p21_array_index_2047660_comb;
    p21_array_index_2047661 <= p21_array_index_2047661_comb;
    p21_res7__274 <= p21_res7__274_comb;
    p22_literal_2043896 <= p21_literal_2043896;
    p22_literal_2043910 <= p21_literal_2043910;
    p22_literal_2043912 <= p21_literal_2043912;
    p22_literal_2043914 <= p21_literal_2043914;
    p22_literal_2043916 <= p21_literal_2043916;
    p22_literal_2043918 <= p21_literal_2043918;
    p22_literal_2043920 <= p21_literal_2043920;
    p22_literal_2043923 <= p21_literal_2043923;
  end

  // ===== Pipe stage 22:
  wire [7:0] p22_array_index_2047786_comb;
  wire [7:0] p22_res7__276_comb;
  wire [7:0] p22_array_index_2047796_comb;
  wire [7:0] p22_res7__278_comb;
  wire [7:0] p22_res7__280_comb;
  wire [7:0] p22_res7__282_comb;
  wire [7:0] p22_res7__284_comb;
  wire [7:0] p22_res7__286_comb;
  wire [127:0] p22_res__8_comb;
  wire [127:0] p22_xor_2047836_comb;
  wire [127:0] p22_addedKey__41_comb;
  wire [7:0] p22_array_index_2047852_comb;
  wire [7:0] p22_array_index_2047853_comb;
  wire [7:0] p22_array_index_2047854_comb;
  wire [7:0] p22_array_index_2047855_comb;
  wire [7:0] p22_array_index_2047856_comb;
  wire [7:0] p22_array_index_2047857_comb;
  wire [7:0] p22_array_index_2047859_comb;
  wire [7:0] p22_array_index_2047861_comb;
  wire [7:0] p22_array_index_2047862_comb;
  wire [7:0] p22_array_index_2047863_comb;
  wire [7:0] p22_array_index_2047864_comb;
  wire [7:0] p22_array_index_2047865_comb;
  wire [7:0] p22_array_index_2047866_comb;
  wire [7:0] p22_array_index_2047868_comb;
  wire [7:0] p22_array_index_2047869_comb;
  wire [7:0] p22_array_index_2047870_comb;
  assign p22_array_index_2047786_comb = p21_literal_2043920[p21_res7__264];
  assign p22_res7__276_comb = p21_literal_2043910[p21_res7__274] ^ p21_literal_2043912[p21_res7__272] ^ p21_literal_2043914[p21_res7__270] ^ p21_literal_2043916[p21_res7__268] ^ p21_literal_2043918[p21_res7__266] ^ p22_array_index_2047786_comb ^ p21_res7__262 ^ p21_literal_2043923[p21_res7__260] ^ p21_res7__258 ^ p21_array_index_2047626 ^ p21_array_index_2047599 ^ p21_array_index_2047478 ^ p21_array_index_2047446 ^ p21_literal_2043912[p21_array_index_2047431] ^ p21_literal_2043910[p21_array_index_2047432] ^ p21_array_index_2047433;
  assign p22_array_index_2047796_comb = p21_literal_2043920[p21_res7__266];
  assign p22_res7__278_comb = p21_literal_2043910[p22_res7__276_comb] ^ p21_literal_2043912[p21_res7__274] ^ p21_literal_2043914[p21_res7__272] ^ p21_literal_2043916[p21_res7__270] ^ p21_literal_2043918[p21_res7__268] ^ p22_array_index_2047796_comb ^ p21_res7__264 ^ p21_literal_2043923[p21_res7__262] ^ p21_res7__260 ^ p21_array_index_2047638 ^ p21_array_index_2047612 ^ p21_array_index_2047584 ^ p21_array_index_2047463 ^ p21_literal_2043912[p21_array_index_2047430] ^ p21_literal_2043910[p21_array_index_2047431] ^ p21_array_index_2047432;
  assign p22_res7__280_comb = p21_literal_2043910[p22_res7__278_comb] ^ p21_literal_2043912[p22_res7__276_comb] ^ p21_literal_2043914[p21_res7__274] ^ p21_literal_2043916[p21_res7__272] ^ p21_literal_2043918[p21_res7__270] ^ p21_literal_2043920[p21_res7__268] ^ p21_res7__266 ^ p21_literal_2043923[p21_res7__264] ^ p21_res7__262 ^ p21_array_index_2047650 ^ p21_array_index_2047625 ^ p21_array_index_2047598 ^ p21_array_index_2047477 ^ p21_array_index_2047445 ^ p21_literal_2043910[p21_array_index_2047430] ^ p21_array_index_2047431;
  assign p22_res7__282_comb = p21_literal_2043910[p22_res7__280_comb] ^ p21_literal_2043912[p22_res7__278_comb] ^ p21_literal_2043914[p22_res7__276_comb] ^ p21_literal_2043916[p21_res7__274] ^ p21_literal_2043918[p21_res7__272] ^ p21_literal_2043920[p21_res7__270] ^ p21_res7__268 ^ p21_literal_2043923[p21_res7__266] ^ p21_res7__264 ^ p21_array_index_2047661 ^ p21_array_index_2047637 ^ p21_array_index_2047611 ^ p21_array_index_2047583 ^ p21_array_index_2047462 ^ p21_literal_2043910[p21_array_index_2047429] ^ p21_array_index_2047430;
  assign p22_res7__284_comb = p21_literal_2043910[p22_res7__282_comb] ^ p21_literal_2043912[p22_res7__280_comb] ^ p21_literal_2043914[p22_res7__278_comb] ^ p21_literal_2043916[p22_res7__276_comb] ^ p21_literal_2043918[p21_res7__274] ^ p21_literal_2043920[p21_res7__272] ^ p21_res7__270 ^ p21_literal_2043923[p21_res7__268] ^ p21_res7__266 ^ p22_array_index_2047786_comb ^ p21_array_index_2047649 ^ p21_array_index_2047624 ^ p21_array_index_2047597 ^ p21_array_index_2047476 ^ p21_array_index_2047444 ^ p21_array_index_2047429;
  assign p22_res7__286_comb = p21_literal_2043910[p22_res7__284_comb] ^ p21_literal_2043912[p22_res7__282_comb] ^ p21_literal_2043914[p22_res7__280_comb] ^ p21_literal_2043916[p22_res7__278_comb] ^ p21_literal_2043918[p22_res7__276_comb] ^ p21_literal_2043920[p21_res7__274] ^ p21_res7__272 ^ p21_literal_2043923[p21_res7__270] ^ p21_res7__268 ^ p22_array_index_2047796_comb ^ p21_array_index_2047660 ^ p21_array_index_2047636 ^ p21_array_index_2047610 ^ p21_array_index_2047582 ^ p21_array_index_2047461 ^ p21_array_index_2047428;
  assign p22_res__8_comb = {p22_res7__286_comb, p22_res7__284_comb, p22_res7__282_comb, p22_res7__280_comb, p22_res7__278_comb, p22_res7__276_comb, p21_res7__274, p21_res7__272, p21_res7__270, p21_res7__268, p21_res7__266, p21_res7__264, p21_res7__262, p21_res7__260, p21_res7__258, p21_res7__256};
  assign p22_xor_2047836_comb = p22_res__8_comb ^ p21_k3;
  assign p22_addedKey__41_comb = p22_xor_2047836_comb ^ 128'h2ade_daf2_3e95_a23a_17b5_18a0_5e61_c10a;
  assign p22_array_index_2047852_comb = p21_literal_2043896[p22_addedKey__41_comb[127:120]];
  assign p22_array_index_2047853_comb = p21_literal_2043896[p22_addedKey__41_comb[119:112]];
  assign p22_array_index_2047854_comb = p21_literal_2043896[p22_addedKey__41_comb[111:104]];
  assign p22_array_index_2047855_comb = p21_literal_2043896[p22_addedKey__41_comb[103:96]];
  assign p22_array_index_2047856_comb = p21_literal_2043896[p22_addedKey__41_comb[95:88]];
  assign p22_array_index_2047857_comb = p21_literal_2043896[p22_addedKey__41_comb[87:80]];
  assign p22_array_index_2047859_comb = p21_literal_2043896[p22_addedKey__41_comb[71:64]];
  assign p22_array_index_2047861_comb = p21_literal_2043896[p22_addedKey__41_comb[55:48]];
  assign p22_array_index_2047862_comb = p21_literal_2043896[p22_addedKey__41_comb[47:40]];
  assign p22_array_index_2047863_comb = p21_literal_2043896[p22_addedKey__41_comb[39:32]];
  assign p22_array_index_2047864_comb = p21_literal_2043896[p22_addedKey__41_comb[31:24]];
  assign p22_array_index_2047865_comb = p21_literal_2043896[p22_addedKey__41_comb[23:16]];
  assign p22_array_index_2047866_comb = p21_literal_2043896[p22_addedKey__41_comb[15:8]];
  assign p22_array_index_2047868_comb = p21_literal_2043896[p22_addedKey__41_comb[79:72]];
  assign p22_array_index_2047869_comb = p21_literal_2043896[p22_addedKey__41_comb[63:56]];
  assign p22_array_index_2047870_comb = p21_literal_2043896[p22_addedKey__41_comb[7:0]];

  // Registers for pipe stage 22:
  reg [127:0] p22_encoded;
  reg [127:0] p22_bit_slice_2043893;
  reg [127:0] p22_bit_slice_2044018;
  reg [127:0] p22_k3;
  reg [127:0] p22_k2;
  reg [127:0] p22_xor_2047836;
  reg [7:0] p22_array_index_2047852;
  reg [7:0] p22_array_index_2047853;
  reg [7:0] p22_array_index_2047854;
  reg [7:0] p22_array_index_2047855;
  reg [7:0] p22_array_index_2047856;
  reg [7:0] p22_array_index_2047857;
  reg [7:0] p22_array_index_2047859;
  reg [7:0] p22_array_index_2047861;
  reg [7:0] p22_array_index_2047862;
  reg [7:0] p22_array_index_2047863;
  reg [7:0] p22_array_index_2047864;
  reg [7:0] p22_array_index_2047865;
  reg [7:0] p22_array_index_2047866;
  reg [7:0] p22_array_index_2047868;
  reg [7:0] p22_array_index_2047869;
  reg [7:0] p22_array_index_2047870;
  reg [7:0] p23_literal_2043896[256];
  reg [7:0] p23_literal_2043910[256];
  reg [7:0] p23_literal_2043912[256];
  reg [7:0] p23_literal_2043914[256];
  reg [7:0] p23_literal_2043916[256];
  reg [7:0] p23_literal_2043918[256];
  reg [7:0] p23_literal_2043920[256];
  reg [7:0] p23_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p22_encoded <= p21_encoded;
    p22_bit_slice_2043893 <= p21_bit_slice_2043893;
    p22_bit_slice_2044018 <= p21_bit_slice_2044018;
    p22_k3 <= p21_k3;
    p22_k2 <= p21_k2;
    p22_xor_2047836 <= p22_xor_2047836_comb;
    p22_array_index_2047852 <= p22_array_index_2047852_comb;
    p22_array_index_2047853 <= p22_array_index_2047853_comb;
    p22_array_index_2047854 <= p22_array_index_2047854_comb;
    p22_array_index_2047855 <= p22_array_index_2047855_comb;
    p22_array_index_2047856 <= p22_array_index_2047856_comb;
    p22_array_index_2047857 <= p22_array_index_2047857_comb;
    p22_array_index_2047859 <= p22_array_index_2047859_comb;
    p22_array_index_2047861 <= p22_array_index_2047861_comb;
    p22_array_index_2047862 <= p22_array_index_2047862_comb;
    p22_array_index_2047863 <= p22_array_index_2047863_comb;
    p22_array_index_2047864 <= p22_array_index_2047864_comb;
    p22_array_index_2047865 <= p22_array_index_2047865_comb;
    p22_array_index_2047866 <= p22_array_index_2047866_comb;
    p22_array_index_2047868 <= p22_array_index_2047868_comb;
    p22_array_index_2047869 <= p22_array_index_2047869_comb;
    p22_array_index_2047870 <= p22_array_index_2047870_comb;
    p23_literal_2043896 <= p22_literal_2043896;
    p23_literal_2043910 <= p22_literal_2043910;
    p23_literal_2043912 <= p22_literal_2043912;
    p23_literal_2043914 <= p22_literal_2043914;
    p23_literal_2043916 <= p22_literal_2043916;
    p23_literal_2043918 <= p22_literal_2043918;
    p23_literal_2043920 <= p22_literal_2043920;
    p23_literal_2043923 <= p22_literal_2043923;
  end

  // ===== Pipe stage 23:
  wire [7:0] p23_array_index_2047931_comb;
  wire [7:0] p23_array_index_2047932_comb;
  wire [7:0] p23_array_index_2047933_comb;
  wire [7:0] p23_array_index_2047934_comb;
  wire [7:0] p23_array_index_2047935_comb;
  wire [7:0] p23_array_index_2047936_comb;
  wire [7:0] p23_res7__288_comb;
  wire [7:0] p23_array_index_2047945_comb;
  wire [7:0] p23_array_index_2047946_comb;
  wire [7:0] p23_array_index_2047947_comb;
  wire [7:0] p23_array_index_2047948_comb;
  wire [7:0] p23_array_index_2047949_comb;
  wire [7:0] p23_array_index_2047950_comb;
  wire [7:0] p23_res7__290_comb;
  wire [7:0] p23_array_index_2047960_comb;
  wire [7:0] p23_array_index_2047961_comb;
  wire [7:0] p23_array_index_2047962_comb;
  wire [7:0] p23_array_index_2047963_comb;
  wire [7:0] p23_array_index_2047964_comb;
  wire [7:0] p23_res7__292_comb;
  wire [7:0] p23_array_index_2047974_comb;
  wire [7:0] p23_array_index_2047975_comb;
  wire [7:0] p23_array_index_2047976_comb;
  wire [7:0] p23_array_index_2047977_comb;
  wire [7:0] p23_array_index_2047978_comb;
  wire [7:0] p23_res7__294_comb;
  wire [7:0] p23_array_index_2047989_comb;
  wire [7:0] p23_array_index_2047990_comb;
  wire [7:0] p23_array_index_2047991_comb;
  wire [7:0] p23_array_index_2047992_comb;
  wire [7:0] p23_res7__296_comb;
  wire [7:0] p23_array_index_2048002_comb;
  wire [7:0] p23_array_index_2048003_comb;
  wire [7:0] p23_array_index_2048004_comb;
  wire [7:0] p23_array_index_2048005_comb;
  wire [7:0] p23_res7__298_comb;
  wire [7:0] p23_array_index_2048016_comb;
  wire [7:0] p23_array_index_2048017_comb;
  wire [7:0] p23_array_index_2048018_comb;
  wire [7:0] p23_res7__300_comb;
  assign p23_array_index_2047931_comb = p22_literal_2043910[p22_array_index_2047852];
  assign p23_array_index_2047932_comb = p22_literal_2043912[p22_array_index_2047853];
  assign p23_array_index_2047933_comb = p22_literal_2043914[p22_array_index_2047854];
  assign p23_array_index_2047934_comb = p22_literal_2043916[p22_array_index_2047855];
  assign p23_array_index_2047935_comb = p22_literal_2043918[p22_array_index_2047856];
  assign p23_array_index_2047936_comb = p22_literal_2043920[p22_array_index_2047857];
  assign p23_res7__288_comb = p23_array_index_2047931_comb ^ p23_array_index_2047932_comb ^ p23_array_index_2047933_comb ^ p23_array_index_2047934_comb ^ p23_array_index_2047935_comb ^ p23_array_index_2047936_comb ^ p22_array_index_2047868 ^ p22_literal_2043923[p22_array_index_2047859] ^ p22_array_index_2047869 ^ p22_literal_2043920[p22_array_index_2047861] ^ p22_literal_2043918[p22_array_index_2047862] ^ p22_literal_2043916[p22_array_index_2047863] ^ p22_literal_2043914[p22_array_index_2047864] ^ p22_literal_2043912[p22_array_index_2047865] ^ p22_literal_2043910[p22_array_index_2047866] ^ p22_array_index_2047870;
  assign p23_array_index_2047945_comb = p22_literal_2043910[p23_res7__288_comb];
  assign p23_array_index_2047946_comb = p22_literal_2043912[p22_array_index_2047852];
  assign p23_array_index_2047947_comb = p22_literal_2043914[p22_array_index_2047853];
  assign p23_array_index_2047948_comb = p22_literal_2043916[p22_array_index_2047854];
  assign p23_array_index_2047949_comb = p22_literal_2043918[p22_array_index_2047855];
  assign p23_array_index_2047950_comb = p22_literal_2043920[p22_array_index_2047856];
  assign p23_res7__290_comb = p23_array_index_2047945_comb ^ p23_array_index_2047946_comb ^ p23_array_index_2047947_comb ^ p23_array_index_2047948_comb ^ p23_array_index_2047949_comb ^ p23_array_index_2047950_comb ^ p22_array_index_2047857 ^ p22_literal_2043923[p22_array_index_2047868] ^ p22_array_index_2047859 ^ p22_literal_2043920[p22_array_index_2047869] ^ p22_literal_2043918[p22_array_index_2047861] ^ p22_literal_2043916[p22_array_index_2047862] ^ p22_literal_2043914[p22_array_index_2047863] ^ p22_literal_2043912[p22_array_index_2047864] ^ p22_literal_2043910[p22_array_index_2047865] ^ p22_array_index_2047866;
  assign p23_array_index_2047960_comb = p22_literal_2043912[p23_res7__288_comb];
  assign p23_array_index_2047961_comb = p22_literal_2043914[p22_array_index_2047852];
  assign p23_array_index_2047962_comb = p22_literal_2043916[p22_array_index_2047853];
  assign p23_array_index_2047963_comb = p22_literal_2043918[p22_array_index_2047854];
  assign p23_array_index_2047964_comb = p22_literal_2043920[p22_array_index_2047855];
  assign p23_res7__292_comb = p22_literal_2043910[p23_res7__290_comb] ^ p23_array_index_2047960_comb ^ p23_array_index_2047961_comb ^ p23_array_index_2047962_comb ^ p23_array_index_2047963_comb ^ p23_array_index_2047964_comb ^ p22_array_index_2047856 ^ p22_literal_2043923[p22_array_index_2047857] ^ p22_array_index_2047868 ^ p22_literal_2043920[p22_array_index_2047859] ^ p22_literal_2043918[p22_array_index_2047869] ^ p22_literal_2043916[p22_array_index_2047861] ^ p22_literal_2043914[p22_array_index_2047862] ^ p22_literal_2043912[p22_array_index_2047863] ^ p22_literal_2043910[p22_array_index_2047864] ^ p22_array_index_2047865;
  assign p23_array_index_2047974_comb = p22_literal_2043912[p23_res7__290_comb];
  assign p23_array_index_2047975_comb = p22_literal_2043914[p23_res7__288_comb];
  assign p23_array_index_2047976_comb = p22_literal_2043916[p22_array_index_2047852];
  assign p23_array_index_2047977_comb = p22_literal_2043918[p22_array_index_2047853];
  assign p23_array_index_2047978_comb = p22_literal_2043920[p22_array_index_2047854];
  assign p23_res7__294_comb = p22_literal_2043910[p23_res7__292_comb] ^ p23_array_index_2047974_comb ^ p23_array_index_2047975_comb ^ p23_array_index_2047976_comb ^ p23_array_index_2047977_comb ^ p23_array_index_2047978_comb ^ p22_array_index_2047855 ^ p22_literal_2043923[p22_array_index_2047856] ^ p22_array_index_2047857 ^ p22_literal_2043920[p22_array_index_2047868] ^ p22_literal_2043918[p22_array_index_2047859] ^ p22_literal_2043916[p22_array_index_2047869] ^ p22_literal_2043914[p22_array_index_2047861] ^ p22_literal_2043912[p22_array_index_2047862] ^ p22_literal_2043910[p22_array_index_2047863] ^ p22_array_index_2047864;
  assign p23_array_index_2047989_comb = p22_literal_2043914[p23_res7__290_comb];
  assign p23_array_index_2047990_comb = p22_literal_2043916[p23_res7__288_comb];
  assign p23_array_index_2047991_comb = p22_literal_2043918[p22_array_index_2047852];
  assign p23_array_index_2047992_comb = p22_literal_2043920[p22_array_index_2047853];
  assign p23_res7__296_comb = p22_literal_2043910[p23_res7__294_comb] ^ p22_literal_2043912[p23_res7__292_comb] ^ p23_array_index_2047989_comb ^ p23_array_index_2047990_comb ^ p23_array_index_2047991_comb ^ p23_array_index_2047992_comb ^ p22_array_index_2047854 ^ p22_literal_2043923[p22_array_index_2047855] ^ p22_array_index_2047856 ^ p23_array_index_2047936_comb ^ p22_literal_2043918[p22_array_index_2047868] ^ p22_literal_2043916[p22_array_index_2047859] ^ p22_literal_2043914[p22_array_index_2047869] ^ p22_literal_2043912[p22_array_index_2047861] ^ p22_literal_2043910[p22_array_index_2047862] ^ p22_array_index_2047863;
  assign p23_array_index_2048002_comb = p22_literal_2043914[p23_res7__292_comb];
  assign p23_array_index_2048003_comb = p22_literal_2043916[p23_res7__290_comb];
  assign p23_array_index_2048004_comb = p22_literal_2043918[p23_res7__288_comb];
  assign p23_array_index_2048005_comb = p22_literal_2043920[p22_array_index_2047852];
  assign p23_res7__298_comb = p22_literal_2043910[p23_res7__296_comb] ^ p22_literal_2043912[p23_res7__294_comb] ^ p23_array_index_2048002_comb ^ p23_array_index_2048003_comb ^ p23_array_index_2048004_comb ^ p23_array_index_2048005_comb ^ p22_array_index_2047853 ^ p22_literal_2043923[p22_array_index_2047854] ^ p22_array_index_2047855 ^ p23_array_index_2047950_comb ^ p22_literal_2043918[p22_array_index_2047857] ^ p22_literal_2043916[p22_array_index_2047868] ^ p22_literal_2043914[p22_array_index_2047859] ^ p22_literal_2043912[p22_array_index_2047869] ^ p22_literal_2043910[p22_array_index_2047861] ^ p22_array_index_2047862;
  assign p23_array_index_2048016_comb = p22_literal_2043916[p23_res7__292_comb];
  assign p23_array_index_2048017_comb = p22_literal_2043918[p23_res7__290_comb];
  assign p23_array_index_2048018_comb = p22_literal_2043920[p23_res7__288_comb];
  assign p23_res7__300_comb = p22_literal_2043910[p23_res7__298_comb] ^ p22_literal_2043912[p23_res7__296_comb] ^ p22_literal_2043914[p23_res7__294_comb] ^ p23_array_index_2048016_comb ^ p23_array_index_2048017_comb ^ p23_array_index_2048018_comb ^ p22_array_index_2047852 ^ p22_literal_2043923[p22_array_index_2047853] ^ p22_array_index_2047854 ^ p23_array_index_2047964_comb ^ p23_array_index_2047935_comb ^ p22_literal_2043916[p22_array_index_2047857] ^ p22_literal_2043914[p22_array_index_2047868] ^ p22_literal_2043912[p22_array_index_2047859] ^ p22_literal_2043910[p22_array_index_2047869] ^ p22_array_index_2047861;

  // Registers for pipe stage 23:
  reg [127:0] p23_encoded;
  reg [127:0] p23_bit_slice_2043893;
  reg [127:0] p23_bit_slice_2044018;
  reg [127:0] p23_k3;
  reg [127:0] p23_k2;
  reg [127:0] p23_xor_2047836;
  reg [7:0] p23_array_index_2047852;
  reg [7:0] p23_array_index_2047853;
  reg [7:0] p23_array_index_2047854;
  reg [7:0] p23_array_index_2047855;
  reg [7:0] p23_array_index_2047856;
  reg [7:0] p23_array_index_2047857;
  reg [7:0] p23_array_index_2047859;
  reg [7:0] p23_array_index_2047931;
  reg [7:0] p23_array_index_2047932;
  reg [7:0] p23_array_index_2047933;
  reg [7:0] p23_array_index_2047934;
  reg [7:0] p23_array_index_2047868;
  reg [7:0] p23_array_index_2047869;
  reg [7:0] p23_res7__288;
  reg [7:0] p23_array_index_2047945;
  reg [7:0] p23_array_index_2047946;
  reg [7:0] p23_array_index_2047947;
  reg [7:0] p23_array_index_2047948;
  reg [7:0] p23_array_index_2047949;
  reg [7:0] p23_res7__290;
  reg [7:0] p23_array_index_2047960;
  reg [7:0] p23_array_index_2047961;
  reg [7:0] p23_array_index_2047962;
  reg [7:0] p23_array_index_2047963;
  reg [7:0] p23_res7__292;
  reg [7:0] p23_array_index_2047974;
  reg [7:0] p23_array_index_2047975;
  reg [7:0] p23_array_index_2047976;
  reg [7:0] p23_array_index_2047977;
  reg [7:0] p23_array_index_2047978;
  reg [7:0] p23_res7__294;
  reg [7:0] p23_array_index_2047989;
  reg [7:0] p23_array_index_2047990;
  reg [7:0] p23_array_index_2047991;
  reg [7:0] p23_array_index_2047992;
  reg [7:0] p23_res7__296;
  reg [7:0] p23_array_index_2048002;
  reg [7:0] p23_array_index_2048003;
  reg [7:0] p23_array_index_2048004;
  reg [7:0] p23_array_index_2048005;
  reg [7:0] p23_res7__298;
  reg [7:0] p23_array_index_2048016;
  reg [7:0] p23_array_index_2048017;
  reg [7:0] p23_array_index_2048018;
  reg [7:0] p23_res7__300;
  reg [7:0] p24_literal_2043896[256];
  reg [7:0] p24_literal_2043910[256];
  reg [7:0] p24_literal_2043912[256];
  reg [7:0] p24_literal_2043914[256];
  reg [7:0] p24_literal_2043916[256];
  reg [7:0] p24_literal_2043918[256];
  reg [7:0] p24_literal_2043920[256];
  reg [7:0] p24_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p23_encoded <= p22_encoded;
    p23_bit_slice_2043893 <= p22_bit_slice_2043893;
    p23_bit_slice_2044018 <= p22_bit_slice_2044018;
    p23_k3 <= p22_k3;
    p23_k2 <= p22_k2;
    p23_xor_2047836 <= p22_xor_2047836;
    p23_array_index_2047852 <= p22_array_index_2047852;
    p23_array_index_2047853 <= p22_array_index_2047853;
    p23_array_index_2047854 <= p22_array_index_2047854;
    p23_array_index_2047855 <= p22_array_index_2047855;
    p23_array_index_2047856 <= p22_array_index_2047856;
    p23_array_index_2047857 <= p22_array_index_2047857;
    p23_array_index_2047859 <= p22_array_index_2047859;
    p23_array_index_2047931 <= p23_array_index_2047931_comb;
    p23_array_index_2047932 <= p23_array_index_2047932_comb;
    p23_array_index_2047933 <= p23_array_index_2047933_comb;
    p23_array_index_2047934 <= p23_array_index_2047934_comb;
    p23_array_index_2047868 <= p22_array_index_2047868;
    p23_array_index_2047869 <= p22_array_index_2047869;
    p23_res7__288 <= p23_res7__288_comb;
    p23_array_index_2047945 <= p23_array_index_2047945_comb;
    p23_array_index_2047946 <= p23_array_index_2047946_comb;
    p23_array_index_2047947 <= p23_array_index_2047947_comb;
    p23_array_index_2047948 <= p23_array_index_2047948_comb;
    p23_array_index_2047949 <= p23_array_index_2047949_comb;
    p23_res7__290 <= p23_res7__290_comb;
    p23_array_index_2047960 <= p23_array_index_2047960_comb;
    p23_array_index_2047961 <= p23_array_index_2047961_comb;
    p23_array_index_2047962 <= p23_array_index_2047962_comb;
    p23_array_index_2047963 <= p23_array_index_2047963_comb;
    p23_res7__292 <= p23_res7__292_comb;
    p23_array_index_2047974 <= p23_array_index_2047974_comb;
    p23_array_index_2047975 <= p23_array_index_2047975_comb;
    p23_array_index_2047976 <= p23_array_index_2047976_comb;
    p23_array_index_2047977 <= p23_array_index_2047977_comb;
    p23_array_index_2047978 <= p23_array_index_2047978_comb;
    p23_res7__294 <= p23_res7__294_comb;
    p23_array_index_2047989 <= p23_array_index_2047989_comb;
    p23_array_index_2047990 <= p23_array_index_2047990_comb;
    p23_array_index_2047991 <= p23_array_index_2047991_comb;
    p23_array_index_2047992 <= p23_array_index_2047992_comb;
    p23_res7__296 <= p23_res7__296_comb;
    p23_array_index_2048002 <= p23_array_index_2048002_comb;
    p23_array_index_2048003 <= p23_array_index_2048003_comb;
    p23_array_index_2048004 <= p23_array_index_2048004_comb;
    p23_array_index_2048005 <= p23_array_index_2048005_comb;
    p23_res7__298 <= p23_res7__298_comb;
    p23_array_index_2048016 <= p23_array_index_2048016_comb;
    p23_array_index_2048017 <= p23_array_index_2048017_comb;
    p23_array_index_2048018 <= p23_array_index_2048018_comb;
    p23_res7__300 <= p23_res7__300_comb;
    p24_literal_2043896 <= p23_literal_2043896;
    p24_literal_2043910 <= p23_literal_2043910;
    p24_literal_2043912 <= p23_literal_2043912;
    p24_literal_2043914 <= p23_literal_2043914;
    p24_literal_2043916 <= p23_literal_2043916;
    p24_literal_2043918 <= p23_literal_2043918;
    p24_literal_2043920 <= p23_literal_2043920;
    p24_literal_2043923 <= p23_literal_2043923;
  end

  // ===== Pipe stage 24:
  wire [7:0] p24_array_index_2048146_comb;
  wire [7:0] p24_array_index_2048147_comb;
  wire [7:0] p24_array_index_2048148_comb;
  wire [7:0] p24_res7__302_comb;
  wire [7:0] p24_array_index_2048159_comb;
  wire [7:0] p24_array_index_2048160_comb;
  wire [7:0] p24_res7__304_comb;
  wire [7:0] p24_array_index_2048170_comb;
  wire [7:0] p24_array_index_2048171_comb;
  wire [7:0] p24_res7__306_comb;
  wire [7:0] p24_array_index_2048182_comb;
  wire [7:0] p24_res7__308_comb;
  wire [7:0] p24_array_index_2048192_comb;
  wire [7:0] p24_res7__310_comb;
  wire [7:0] p24_res7__312_comb;
  wire [7:0] p24_res7__314_comb;
  assign p24_array_index_2048146_comb = p23_literal_2043916[p23_res7__294];
  assign p24_array_index_2048147_comb = p23_literal_2043918[p23_res7__292];
  assign p24_array_index_2048148_comb = p23_literal_2043920[p23_res7__290];
  assign p24_res7__302_comb = p23_literal_2043910[p23_res7__300] ^ p23_literal_2043912[p23_res7__298] ^ p23_literal_2043914[p23_res7__296] ^ p24_array_index_2048146_comb ^ p24_array_index_2048147_comb ^ p24_array_index_2048148_comb ^ p23_res7__288 ^ p23_literal_2043923[p23_array_index_2047852] ^ p23_array_index_2047853 ^ p23_array_index_2047978 ^ p23_array_index_2047949 ^ p23_literal_2043916[p23_array_index_2047856] ^ p23_literal_2043914[p23_array_index_2047857] ^ p23_literal_2043912[p23_array_index_2047868] ^ p23_literal_2043910[p23_array_index_2047859] ^ p23_array_index_2047869;
  assign p24_array_index_2048159_comb = p23_literal_2043918[p23_res7__294];
  assign p24_array_index_2048160_comb = p23_literal_2043920[p23_res7__292];
  assign p24_res7__304_comb = p23_literal_2043910[p24_res7__302_comb] ^ p23_literal_2043912[p23_res7__300] ^ p23_literal_2043914[p23_res7__298] ^ p23_literal_2043916[p23_res7__296] ^ p24_array_index_2048159_comb ^ p24_array_index_2048160_comb ^ p23_res7__290 ^ p23_literal_2043923[p23_res7__288] ^ p23_array_index_2047852 ^ p23_array_index_2047992 ^ p23_array_index_2047963 ^ p23_array_index_2047934 ^ p23_literal_2043914[p23_array_index_2047856] ^ p23_literal_2043912[p23_array_index_2047857] ^ p23_literal_2043910[p23_array_index_2047868] ^ p23_array_index_2047859;
  assign p24_array_index_2048170_comb = p23_literal_2043918[p23_res7__296];
  assign p24_array_index_2048171_comb = p23_literal_2043920[p23_res7__294];
  assign p24_res7__306_comb = p23_literal_2043910[p24_res7__304_comb] ^ p23_literal_2043912[p24_res7__302_comb] ^ p23_literal_2043914[p23_res7__300] ^ p23_literal_2043916[p23_res7__298] ^ p24_array_index_2048170_comb ^ p24_array_index_2048171_comb ^ p23_res7__292 ^ p23_literal_2043923[p23_res7__290] ^ p23_res7__288 ^ p23_array_index_2048005 ^ p23_array_index_2047977 ^ p23_array_index_2047948 ^ p23_literal_2043914[p23_array_index_2047855] ^ p23_literal_2043912[p23_array_index_2047856] ^ p23_literal_2043910[p23_array_index_2047857] ^ p23_array_index_2047868;
  assign p24_array_index_2048182_comb = p23_literal_2043920[p23_res7__296];
  assign p24_res7__308_comb = p23_literal_2043910[p24_res7__306_comb] ^ p23_literal_2043912[p24_res7__304_comb] ^ p23_literal_2043914[p24_res7__302_comb] ^ p23_literal_2043916[p23_res7__300] ^ p23_literal_2043918[p23_res7__298] ^ p24_array_index_2048182_comb ^ p23_res7__294 ^ p23_literal_2043923[p23_res7__292] ^ p23_res7__290 ^ p23_array_index_2048018 ^ p23_array_index_2047991 ^ p23_array_index_2047962 ^ p23_array_index_2047933 ^ p23_literal_2043912[p23_array_index_2047855] ^ p23_literal_2043910[p23_array_index_2047856] ^ p23_array_index_2047857;
  assign p24_array_index_2048192_comb = p23_literal_2043920[p23_res7__298];
  assign p24_res7__310_comb = p23_literal_2043910[p24_res7__308_comb] ^ p23_literal_2043912[p24_res7__306_comb] ^ p23_literal_2043914[p24_res7__304_comb] ^ p23_literal_2043916[p24_res7__302_comb] ^ p23_literal_2043918[p23_res7__300] ^ p24_array_index_2048192_comb ^ p23_res7__296 ^ p23_literal_2043923[p23_res7__294] ^ p23_res7__292 ^ p24_array_index_2048148_comb ^ p23_array_index_2048004 ^ p23_array_index_2047976 ^ p23_array_index_2047947 ^ p23_literal_2043912[p23_array_index_2047854] ^ p23_literal_2043910[p23_array_index_2047855] ^ p23_array_index_2047856;
  assign p24_res7__312_comb = p23_literal_2043910[p24_res7__310_comb] ^ p23_literal_2043912[p24_res7__308_comb] ^ p23_literal_2043914[p24_res7__306_comb] ^ p23_literal_2043916[p24_res7__304_comb] ^ p23_literal_2043918[p24_res7__302_comb] ^ p23_literal_2043920[p23_res7__300] ^ p23_res7__298 ^ p23_literal_2043923[p23_res7__296] ^ p23_res7__294 ^ p24_array_index_2048160_comb ^ p23_array_index_2048017 ^ p23_array_index_2047990 ^ p23_array_index_2047961 ^ p23_array_index_2047932 ^ p23_literal_2043910[p23_array_index_2047854] ^ p23_array_index_2047855;
  assign p24_res7__314_comb = p23_literal_2043910[p24_res7__312_comb] ^ p23_literal_2043912[p24_res7__310_comb] ^ p23_literal_2043914[p24_res7__308_comb] ^ p23_literal_2043916[p24_res7__306_comb] ^ p23_literal_2043918[p24_res7__304_comb] ^ p23_literal_2043920[p24_res7__302_comb] ^ p23_res7__300 ^ p23_literal_2043923[p23_res7__298] ^ p23_res7__296 ^ p24_array_index_2048171_comb ^ p24_array_index_2048147_comb ^ p23_array_index_2048003 ^ p23_array_index_2047975 ^ p23_array_index_2047946 ^ p23_literal_2043910[p23_array_index_2047853] ^ p23_array_index_2047854;

  // Registers for pipe stage 24:
  reg [127:0] p24_encoded;
  reg [127:0] p24_bit_slice_2043893;
  reg [127:0] p24_bit_slice_2044018;
  reg [127:0] p24_k3;
  reg [127:0] p24_k2;
  reg [127:0] p24_xor_2047836;
  reg [7:0] p24_array_index_2047852;
  reg [7:0] p24_array_index_2047853;
  reg [7:0] p24_array_index_2047931;
  reg [7:0] p24_res7__288;
  reg [7:0] p24_array_index_2047945;
  reg [7:0] p24_res7__290;
  reg [7:0] p24_array_index_2047960;
  reg [7:0] p24_res7__292;
  reg [7:0] p24_array_index_2047974;
  reg [7:0] p24_res7__294;
  reg [7:0] p24_array_index_2047989;
  reg [7:0] p24_res7__296;
  reg [7:0] p24_array_index_2048002;
  reg [7:0] p24_res7__298;
  reg [7:0] p24_array_index_2048016;
  reg [7:0] p24_res7__300;
  reg [7:0] p24_array_index_2048146;
  reg [7:0] p24_res7__302;
  reg [7:0] p24_array_index_2048159;
  reg [7:0] p24_res7__304;
  reg [7:0] p24_array_index_2048170;
  reg [7:0] p24_res7__306;
  reg [7:0] p24_array_index_2048182;
  reg [7:0] p24_res7__308;
  reg [7:0] p24_array_index_2048192;
  reg [7:0] p24_res7__310;
  reg [7:0] p24_res7__312;
  reg [7:0] p24_res7__314;
  reg [7:0] p25_literal_2043896[256];
  reg [7:0] p25_literal_2043910[256];
  reg [7:0] p25_literal_2043912[256];
  reg [7:0] p25_literal_2043914[256];
  reg [7:0] p25_literal_2043916[256];
  reg [7:0] p25_literal_2043918[256];
  reg [7:0] p25_literal_2043920[256];
  reg [7:0] p25_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p24_encoded <= p23_encoded;
    p24_bit_slice_2043893 <= p23_bit_slice_2043893;
    p24_bit_slice_2044018 <= p23_bit_slice_2044018;
    p24_k3 <= p23_k3;
    p24_k2 <= p23_k2;
    p24_xor_2047836 <= p23_xor_2047836;
    p24_array_index_2047852 <= p23_array_index_2047852;
    p24_array_index_2047853 <= p23_array_index_2047853;
    p24_array_index_2047931 <= p23_array_index_2047931;
    p24_res7__288 <= p23_res7__288;
    p24_array_index_2047945 <= p23_array_index_2047945;
    p24_res7__290 <= p23_res7__290;
    p24_array_index_2047960 <= p23_array_index_2047960;
    p24_res7__292 <= p23_res7__292;
    p24_array_index_2047974 <= p23_array_index_2047974;
    p24_res7__294 <= p23_res7__294;
    p24_array_index_2047989 <= p23_array_index_2047989;
    p24_res7__296 <= p23_res7__296;
    p24_array_index_2048002 <= p23_array_index_2048002;
    p24_res7__298 <= p23_res7__298;
    p24_array_index_2048016 <= p23_array_index_2048016;
    p24_res7__300 <= p23_res7__300;
    p24_array_index_2048146 <= p24_array_index_2048146_comb;
    p24_res7__302 <= p24_res7__302_comb;
    p24_array_index_2048159 <= p24_array_index_2048159_comb;
    p24_res7__304 <= p24_res7__304_comb;
    p24_array_index_2048170 <= p24_array_index_2048170_comb;
    p24_res7__306 <= p24_res7__306_comb;
    p24_array_index_2048182 <= p24_array_index_2048182_comb;
    p24_res7__308 <= p24_res7__308_comb;
    p24_array_index_2048192 <= p24_array_index_2048192_comb;
    p24_res7__310 <= p24_res7__310_comb;
    p24_res7__312 <= p24_res7__312_comb;
    p24_res7__314 <= p24_res7__314_comb;
    p25_literal_2043896 <= p24_literal_2043896;
    p25_literal_2043910 <= p24_literal_2043910;
    p25_literal_2043912 <= p24_literal_2043912;
    p25_literal_2043914 <= p24_literal_2043914;
    p25_literal_2043916 <= p24_literal_2043916;
    p25_literal_2043918 <= p24_literal_2043918;
    p25_literal_2043920 <= p24_literal_2043920;
    p25_literal_2043923 <= p24_literal_2043923;
  end

  // ===== Pipe stage 25:
  wire [7:0] p25_res7__316_comb;
  wire [7:0] p25_res7__318_comb;
  wire [127:0] p25_res__9_comb;
  wire [127:0] p25_xor_2048316_comb;
  wire [127:0] p25_addedKey__42_comb;
  wire [7:0] p25_array_index_2048332_comb;
  wire [7:0] p25_array_index_2048333_comb;
  wire [7:0] p25_array_index_2048334_comb;
  wire [7:0] p25_array_index_2048335_comb;
  wire [7:0] p25_array_index_2048336_comb;
  wire [7:0] p25_array_index_2048337_comb;
  wire [7:0] p25_array_index_2048339_comb;
  wire [7:0] p25_array_index_2048341_comb;
  wire [7:0] p25_array_index_2048342_comb;
  wire [7:0] p25_array_index_2048343_comb;
  wire [7:0] p25_array_index_2048344_comb;
  wire [7:0] p25_array_index_2048345_comb;
  wire [7:0] p25_array_index_2048346_comb;
  wire [7:0] p25_array_index_2048348_comb;
  wire [7:0] p25_array_index_2048349_comb;
  wire [7:0] p25_array_index_2048350_comb;
  wire [7:0] p25_array_index_2048351_comb;
  wire [7:0] p25_array_index_2048352_comb;
  wire [7:0] p25_array_index_2048353_comb;
  wire [7:0] p25_array_index_2048354_comb;
  wire [7:0] p25_array_index_2048356_comb;
  wire [7:0] p25_res7__320_comb;
  wire [7:0] p25_array_index_2048365_comb;
  wire [7:0] p25_array_index_2048366_comb;
  wire [7:0] p25_array_index_2048367_comb;
  wire [7:0] p25_array_index_2048368_comb;
  wire [7:0] p25_array_index_2048369_comb;
  wire [7:0] p25_array_index_2048370_comb;
  wire [7:0] p25_res7__322_comb;
  wire [7:0] p25_array_index_2048380_comb;
  wire [7:0] p25_array_index_2048381_comb;
  wire [7:0] p25_array_index_2048382_comb;
  wire [7:0] p25_array_index_2048383_comb;
  wire [7:0] p25_array_index_2048384_comb;
  wire [7:0] p25_res7__324_comb;
  wire [7:0] p25_array_index_2048394_comb;
  wire [7:0] p25_array_index_2048395_comb;
  wire [7:0] p25_array_index_2048396_comb;
  wire [7:0] p25_array_index_2048397_comb;
  wire [7:0] p25_array_index_2048398_comb;
  wire [7:0] p25_res7__326_comb;
  assign p25_res7__316_comb = p24_literal_2043910[p24_res7__314] ^ p24_literal_2043912[p24_res7__312] ^ p24_literal_2043914[p24_res7__310] ^ p24_literal_2043916[p24_res7__308] ^ p24_literal_2043918[p24_res7__306] ^ p24_literal_2043920[p24_res7__304] ^ p24_res7__302 ^ p24_literal_2043923[p24_res7__300] ^ p24_res7__298 ^ p24_array_index_2048182 ^ p24_array_index_2048159 ^ p24_array_index_2048016 ^ p24_array_index_2047989 ^ p24_array_index_2047960 ^ p24_array_index_2047931 ^ p24_array_index_2047853;
  assign p25_res7__318_comb = p24_literal_2043910[p25_res7__316_comb] ^ p24_literal_2043912[p24_res7__314] ^ p24_literal_2043914[p24_res7__312] ^ p24_literal_2043916[p24_res7__310] ^ p24_literal_2043918[p24_res7__308] ^ p24_literal_2043920[p24_res7__306] ^ p24_res7__304 ^ p24_literal_2043923[p24_res7__302] ^ p24_res7__300 ^ p24_array_index_2048192 ^ p24_array_index_2048170 ^ p24_array_index_2048146 ^ p24_array_index_2048002 ^ p24_array_index_2047974 ^ p24_array_index_2047945 ^ p24_array_index_2047852;
  assign p25_res__9_comb = {p25_res7__318_comb, p25_res7__316_comb, p24_res7__314, p24_res7__312, p24_res7__310, p24_res7__308, p24_res7__306, p24_res7__304, p24_res7__302, p24_res7__300, p24_res7__298, p24_res7__296, p24_res7__294, p24_res7__292, p24_res7__290, p24_res7__288};
  assign p25_xor_2048316_comb = p25_res__9_comb ^ p24_k2;
  assign p25_addedKey__42_comb = p25_xor_2048316_comb ^ 128'h447c_ac80_52dd_d882_4a92_a5b0_83e5_550b;
  assign p25_array_index_2048332_comb = p24_literal_2043896[p25_addedKey__42_comb[127:120]];
  assign p25_array_index_2048333_comb = p24_literal_2043896[p25_addedKey__42_comb[119:112]];
  assign p25_array_index_2048334_comb = p24_literal_2043896[p25_addedKey__42_comb[111:104]];
  assign p25_array_index_2048335_comb = p24_literal_2043896[p25_addedKey__42_comb[103:96]];
  assign p25_array_index_2048336_comb = p24_literal_2043896[p25_addedKey__42_comb[95:88]];
  assign p25_array_index_2048337_comb = p24_literal_2043896[p25_addedKey__42_comb[87:80]];
  assign p25_array_index_2048339_comb = p24_literal_2043896[p25_addedKey__42_comb[71:64]];
  assign p25_array_index_2048341_comb = p24_literal_2043896[p25_addedKey__42_comb[55:48]];
  assign p25_array_index_2048342_comb = p24_literal_2043896[p25_addedKey__42_comb[47:40]];
  assign p25_array_index_2048343_comb = p24_literal_2043896[p25_addedKey__42_comb[39:32]];
  assign p25_array_index_2048344_comb = p24_literal_2043896[p25_addedKey__42_comb[31:24]];
  assign p25_array_index_2048345_comb = p24_literal_2043896[p25_addedKey__42_comb[23:16]];
  assign p25_array_index_2048346_comb = p24_literal_2043896[p25_addedKey__42_comb[15:8]];
  assign p25_array_index_2048348_comb = p24_literal_2043910[p25_array_index_2048332_comb];
  assign p25_array_index_2048349_comb = p24_literal_2043912[p25_array_index_2048333_comb];
  assign p25_array_index_2048350_comb = p24_literal_2043914[p25_array_index_2048334_comb];
  assign p25_array_index_2048351_comb = p24_literal_2043916[p25_array_index_2048335_comb];
  assign p25_array_index_2048352_comb = p24_literal_2043918[p25_array_index_2048336_comb];
  assign p25_array_index_2048353_comb = p24_literal_2043920[p25_array_index_2048337_comb];
  assign p25_array_index_2048354_comb = p24_literal_2043896[p25_addedKey__42_comb[79:72]];
  assign p25_array_index_2048356_comb = p24_literal_2043896[p25_addedKey__42_comb[63:56]];
  assign p25_res7__320_comb = p25_array_index_2048348_comb ^ p25_array_index_2048349_comb ^ p25_array_index_2048350_comb ^ p25_array_index_2048351_comb ^ p25_array_index_2048352_comb ^ p25_array_index_2048353_comb ^ p25_array_index_2048354_comb ^ p24_literal_2043923[p25_array_index_2048339_comb] ^ p25_array_index_2048356_comb ^ p24_literal_2043920[p25_array_index_2048341_comb] ^ p24_literal_2043918[p25_array_index_2048342_comb] ^ p24_literal_2043916[p25_array_index_2048343_comb] ^ p24_literal_2043914[p25_array_index_2048344_comb] ^ p24_literal_2043912[p25_array_index_2048345_comb] ^ p24_literal_2043910[p25_array_index_2048346_comb] ^ p24_literal_2043896[p25_addedKey__42_comb[7:0]];
  assign p25_array_index_2048365_comb = p24_literal_2043910[p25_res7__320_comb];
  assign p25_array_index_2048366_comb = p24_literal_2043912[p25_array_index_2048332_comb];
  assign p25_array_index_2048367_comb = p24_literal_2043914[p25_array_index_2048333_comb];
  assign p25_array_index_2048368_comb = p24_literal_2043916[p25_array_index_2048334_comb];
  assign p25_array_index_2048369_comb = p24_literal_2043918[p25_array_index_2048335_comb];
  assign p25_array_index_2048370_comb = p24_literal_2043920[p25_array_index_2048336_comb];
  assign p25_res7__322_comb = p25_array_index_2048365_comb ^ p25_array_index_2048366_comb ^ p25_array_index_2048367_comb ^ p25_array_index_2048368_comb ^ p25_array_index_2048369_comb ^ p25_array_index_2048370_comb ^ p25_array_index_2048337_comb ^ p24_literal_2043923[p25_array_index_2048354_comb] ^ p25_array_index_2048339_comb ^ p24_literal_2043920[p25_array_index_2048356_comb] ^ p24_literal_2043918[p25_array_index_2048341_comb] ^ p24_literal_2043916[p25_array_index_2048342_comb] ^ p24_literal_2043914[p25_array_index_2048343_comb] ^ p24_literal_2043912[p25_array_index_2048344_comb] ^ p24_literal_2043910[p25_array_index_2048345_comb] ^ p25_array_index_2048346_comb;
  assign p25_array_index_2048380_comb = p24_literal_2043912[p25_res7__320_comb];
  assign p25_array_index_2048381_comb = p24_literal_2043914[p25_array_index_2048332_comb];
  assign p25_array_index_2048382_comb = p24_literal_2043916[p25_array_index_2048333_comb];
  assign p25_array_index_2048383_comb = p24_literal_2043918[p25_array_index_2048334_comb];
  assign p25_array_index_2048384_comb = p24_literal_2043920[p25_array_index_2048335_comb];
  assign p25_res7__324_comb = p24_literal_2043910[p25_res7__322_comb] ^ p25_array_index_2048380_comb ^ p25_array_index_2048381_comb ^ p25_array_index_2048382_comb ^ p25_array_index_2048383_comb ^ p25_array_index_2048384_comb ^ p25_array_index_2048336_comb ^ p24_literal_2043923[p25_array_index_2048337_comb] ^ p25_array_index_2048354_comb ^ p24_literal_2043920[p25_array_index_2048339_comb] ^ p24_literal_2043918[p25_array_index_2048356_comb] ^ p24_literal_2043916[p25_array_index_2048341_comb] ^ p24_literal_2043914[p25_array_index_2048342_comb] ^ p24_literal_2043912[p25_array_index_2048343_comb] ^ p24_literal_2043910[p25_array_index_2048344_comb] ^ p25_array_index_2048345_comb;
  assign p25_array_index_2048394_comb = p24_literal_2043912[p25_res7__322_comb];
  assign p25_array_index_2048395_comb = p24_literal_2043914[p25_res7__320_comb];
  assign p25_array_index_2048396_comb = p24_literal_2043916[p25_array_index_2048332_comb];
  assign p25_array_index_2048397_comb = p24_literal_2043918[p25_array_index_2048333_comb];
  assign p25_array_index_2048398_comb = p24_literal_2043920[p25_array_index_2048334_comb];
  assign p25_res7__326_comb = p24_literal_2043910[p25_res7__324_comb] ^ p25_array_index_2048394_comb ^ p25_array_index_2048395_comb ^ p25_array_index_2048396_comb ^ p25_array_index_2048397_comb ^ p25_array_index_2048398_comb ^ p25_array_index_2048335_comb ^ p24_literal_2043923[p25_array_index_2048336_comb] ^ p25_array_index_2048337_comb ^ p24_literal_2043920[p25_array_index_2048354_comb] ^ p24_literal_2043918[p25_array_index_2048339_comb] ^ p24_literal_2043916[p25_array_index_2048356_comb] ^ p24_literal_2043914[p25_array_index_2048341_comb] ^ p24_literal_2043912[p25_array_index_2048342_comb] ^ p24_literal_2043910[p25_array_index_2048343_comb] ^ p25_array_index_2048344_comb;

  // Registers for pipe stage 25:
  reg [127:0] p25_encoded;
  reg [127:0] p25_bit_slice_2043893;
  reg [127:0] p25_bit_slice_2044018;
  reg [127:0] p25_k3;
  reg [127:0] p25_k2;
  reg [127:0] p25_xor_2047836;
  reg [127:0] p25_xor_2048316;
  reg [7:0] p25_array_index_2048332;
  reg [7:0] p25_array_index_2048333;
  reg [7:0] p25_array_index_2048334;
  reg [7:0] p25_array_index_2048335;
  reg [7:0] p25_array_index_2048336;
  reg [7:0] p25_array_index_2048337;
  reg [7:0] p25_array_index_2048339;
  reg [7:0] p25_array_index_2048341;
  reg [7:0] p25_array_index_2048342;
  reg [7:0] p25_array_index_2048343;
  reg [7:0] p25_array_index_2048348;
  reg [7:0] p25_array_index_2048349;
  reg [7:0] p25_array_index_2048350;
  reg [7:0] p25_array_index_2048351;
  reg [7:0] p25_array_index_2048352;
  reg [7:0] p25_array_index_2048353;
  reg [7:0] p25_array_index_2048354;
  reg [7:0] p25_array_index_2048356;
  reg [7:0] p25_res7__320;
  reg [7:0] p25_array_index_2048365;
  reg [7:0] p25_array_index_2048366;
  reg [7:0] p25_array_index_2048367;
  reg [7:0] p25_array_index_2048368;
  reg [7:0] p25_array_index_2048369;
  reg [7:0] p25_array_index_2048370;
  reg [7:0] p25_res7__322;
  reg [7:0] p25_array_index_2048380;
  reg [7:0] p25_array_index_2048381;
  reg [7:0] p25_array_index_2048382;
  reg [7:0] p25_array_index_2048383;
  reg [7:0] p25_array_index_2048384;
  reg [7:0] p25_res7__324;
  reg [7:0] p25_array_index_2048394;
  reg [7:0] p25_array_index_2048395;
  reg [7:0] p25_array_index_2048396;
  reg [7:0] p25_array_index_2048397;
  reg [7:0] p25_array_index_2048398;
  reg [7:0] p25_res7__326;
  reg [7:0] p26_literal_2043896[256];
  reg [7:0] p26_literal_2043910[256];
  reg [7:0] p26_literal_2043912[256];
  reg [7:0] p26_literal_2043914[256];
  reg [7:0] p26_literal_2043916[256];
  reg [7:0] p26_literal_2043918[256];
  reg [7:0] p26_literal_2043920[256];
  reg [7:0] p26_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p25_encoded <= p24_encoded;
    p25_bit_slice_2043893 <= p24_bit_slice_2043893;
    p25_bit_slice_2044018 <= p24_bit_slice_2044018;
    p25_k3 <= p24_k3;
    p25_k2 <= p24_k2;
    p25_xor_2047836 <= p24_xor_2047836;
    p25_xor_2048316 <= p25_xor_2048316_comb;
    p25_array_index_2048332 <= p25_array_index_2048332_comb;
    p25_array_index_2048333 <= p25_array_index_2048333_comb;
    p25_array_index_2048334 <= p25_array_index_2048334_comb;
    p25_array_index_2048335 <= p25_array_index_2048335_comb;
    p25_array_index_2048336 <= p25_array_index_2048336_comb;
    p25_array_index_2048337 <= p25_array_index_2048337_comb;
    p25_array_index_2048339 <= p25_array_index_2048339_comb;
    p25_array_index_2048341 <= p25_array_index_2048341_comb;
    p25_array_index_2048342 <= p25_array_index_2048342_comb;
    p25_array_index_2048343 <= p25_array_index_2048343_comb;
    p25_array_index_2048348 <= p25_array_index_2048348_comb;
    p25_array_index_2048349 <= p25_array_index_2048349_comb;
    p25_array_index_2048350 <= p25_array_index_2048350_comb;
    p25_array_index_2048351 <= p25_array_index_2048351_comb;
    p25_array_index_2048352 <= p25_array_index_2048352_comb;
    p25_array_index_2048353 <= p25_array_index_2048353_comb;
    p25_array_index_2048354 <= p25_array_index_2048354_comb;
    p25_array_index_2048356 <= p25_array_index_2048356_comb;
    p25_res7__320 <= p25_res7__320_comb;
    p25_array_index_2048365 <= p25_array_index_2048365_comb;
    p25_array_index_2048366 <= p25_array_index_2048366_comb;
    p25_array_index_2048367 <= p25_array_index_2048367_comb;
    p25_array_index_2048368 <= p25_array_index_2048368_comb;
    p25_array_index_2048369 <= p25_array_index_2048369_comb;
    p25_array_index_2048370 <= p25_array_index_2048370_comb;
    p25_res7__322 <= p25_res7__322_comb;
    p25_array_index_2048380 <= p25_array_index_2048380_comb;
    p25_array_index_2048381 <= p25_array_index_2048381_comb;
    p25_array_index_2048382 <= p25_array_index_2048382_comb;
    p25_array_index_2048383 <= p25_array_index_2048383_comb;
    p25_array_index_2048384 <= p25_array_index_2048384_comb;
    p25_res7__324 <= p25_res7__324_comb;
    p25_array_index_2048394 <= p25_array_index_2048394_comb;
    p25_array_index_2048395 <= p25_array_index_2048395_comb;
    p25_array_index_2048396 <= p25_array_index_2048396_comb;
    p25_array_index_2048397 <= p25_array_index_2048397_comb;
    p25_array_index_2048398 <= p25_array_index_2048398_comb;
    p25_res7__326 <= p25_res7__326_comb;
    p26_literal_2043896 <= p25_literal_2043896;
    p26_literal_2043910 <= p25_literal_2043910;
    p26_literal_2043912 <= p25_literal_2043912;
    p26_literal_2043914 <= p25_literal_2043914;
    p26_literal_2043916 <= p25_literal_2043916;
    p26_literal_2043918 <= p25_literal_2043918;
    p26_literal_2043920 <= p25_literal_2043920;
    p26_literal_2043923 <= p25_literal_2043923;
  end

  // ===== Pipe stage 26:
  wire [7:0] p26_array_index_2048515_comb;
  wire [7:0] p26_array_index_2048516_comb;
  wire [7:0] p26_array_index_2048517_comb;
  wire [7:0] p26_array_index_2048518_comb;
  wire [7:0] p26_res7__328_comb;
  wire [7:0] p26_array_index_2048528_comb;
  wire [7:0] p26_array_index_2048529_comb;
  wire [7:0] p26_array_index_2048530_comb;
  wire [7:0] p26_array_index_2048531_comb;
  wire [7:0] p26_res7__330_comb;
  wire [7:0] p26_array_index_2048542_comb;
  wire [7:0] p26_array_index_2048543_comb;
  wire [7:0] p26_array_index_2048544_comb;
  wire [7:0] p26_res7__332_comb;
  wire [7:0] p26_array_index_2048554_comb;
  wire [7:0] p26_array_index_2048555_comb;
  wire [7:0] p26_array_index_2048556_comb;
  wire [7:0] p26_res7__334_comb;
  wire [7:0] p26_array_index_2048567_comb;
  wire [7:0] p26_array_index_2048568_comb;
  wire [7:0] p26_res7__336_comb;
  wire [7:0] p26_array_index_2048578_comb;
  wire [7:0] p26_array_index_2048579_comb;
  wire [7:0] p26_res7__338_comb;
  wire [7:0] p26_array_index_2048590_comb;
  wire [7:0] p26_res7__340_comb;
  assign p26_array_index_2048515_comb = p25_literal_2043914[p25_res7__322];
  assign p26_array_index_2048516_comb = p25_literal_2043916[p25_res7__320];
  assign p26_array_index_2048517_comb = p25_literal_2043918[p25_array_index_2048332];
  assign p26_array_index_2048518_comb = p25_literal_2043920[p25_array_index_2048333];
  assign p26_res7__328_comb = p25_literal_2043910[p25_res7__326] ^ p25_literal_2043912[p25_res7__324] ^ p26_array_index_2048515_comb ^ p26_array_index_2048516_comb ^ p26_array_index_2048517_comb ^ p26_array_index_2048518_comb ^ p25_array_index_2048334 ^ p25_literal_2043923[p25_array_index_2048335] ^ p25_array_index_2048336 ^ p25_array_index_2048353 ^ p25_literal_2043918[p25_array_index_2048354] ^ p25_literal_2043916[p25_array_index_2048339] ^ p25_literal_2043914[p25_array_index_2048356] ^ p25_literal_2043912[p25_array_index_2048341] ^ p25_literal_2043910[p25_array_index_2048342] ^ p25_array_index_2048343;
  assign p26_array_index_2048528_comb = p25_literal_2043914[p25_res7__324];
  assign p26_array_index_2048529_comb = p25_literal_2043916[p25_res7__322];
  assign p26_array_index_2048530_comb = p25_literal_2043918[p25_res7__320];
  assign p26_array_index_2048531_comb = p25_literal_2043920[p25_array_index_2048332];
  assign p26_res7__330_comb = p25_literal_2043910[p26_res7__328_comb] ^ p25_literal_2043912[p25_res7__326] ^ p26_array_index_2048528_comb ^ p26_array_index_2048529_comb ^ p26_array_index_2048530_comb ^ p26_array_index_2048531_comb ^ p25_array_index_2048333 ^ p25_literal_2043923[p25_array_index_2048334] ^ p25_array_index_2048335 ^ p25_array_index_2048370 ^ p25_literal_2043918[p25_array_index_2048337] ^ p25_literal_2043916[p25_array_index_2048354] ^ p25_literal_2043914[p25_array_index_2048339] ^ p25_literal_2043912[p25_array_index_2048356] ^ p25_literal_2043910[p25_array_index_2048341] ^ p25_array_index_2048342;
  assign p26_array_index_2048542_comb = p25_literal_2043916[p25_res7__324];
  assign p26_array_index_2048543_comb = p25_literal_2043918[p25_res7__322];
  assign p26_array_index_2048544_comb = p25_literal_2043920[p25_res7__320];
  assign p26_res7__332_comb = p25_literal_2043910[p26_res7__330_comb] ^ p25_literal_2043912[p26_res7__328_comb] ^ p25_literal_2043914[p25_res7__326] ^ p26_array_index_2048542_comb ^ p26_array_index_2048543_comb ^ p26_array_index_2048544_comb ^ p25_array_index_2048332 ^ p25_literal_2043923[p25_array_index_2048333] ^ p25_array_index_2048334 ^ p25_array_index_2048384 ^ p25_array_index_2048352 ^ p25_literal_2043916[p25_array_index_2048337] ^ p25_literal_2043914[p25_array_index_2048354] ^ p25_literal_2043912[p25_array_index_2048339] ^ p25_literal_2043910[p25_array_index_2048356] ^ p25_array_index_2048341;
  assign p26_array_index_2048554_comb = p25_literal_2043916[p25_res7__326];
  assign p26_array_index_2048555_comb = p25_literal_2043918[p25_res7__324];
  assign p26_array_index_2048556_comb = p25_literal_2043920[p25_res7__322];
  assign p26_res7__334_comb = p25_literal_2043910[p26_res7__332_comb] ^ p25_literal_2043912[p26_res7__330_comb] ^ p25_literal_2043914[p26_res7__328_comb] ^ p26_array_index_2048554_comb ^ p26_array_index_2048555_comb ^ p26_array_index_2048556_comb ^ p25_res7__320 ^ p25_literal_2043923[p25_array_index_2048332] ^ p25_array_index_2048333 ^ p25_array_index_2048398 ^ p25_array_index_2048369 ^ p25_literal_2043916[p25_array_index_2048336] ^ p25_literal_2043914[p25_array_index_2048337] ^ p25_literal_2043912[p25_array_index_2048354] ^ p25_literal_2043910[p25_array_index_2048339] ^ p25_array_index_2048356;
  assign p26_array_index_2048567_comb = p25_literal_2043918[p25_res7__326];
  assign p26_array_index_2048568_comb = p25_literal_2043920[p25_res7__324];
  assign p26_res7__336_comb = p25_literal_2043910[p26_res7__334_comb] ^ p25_literal_2043912[p26_res7__332_comb] ^ p25_literal_2043914[p26_res7__330_comb] ^ p25_literal_2043916[p26_res7__328_comb] ^ p26_array_index_2048567_comb ^ p26_array_index_2048568_comb ^ p25_res7__322 ^ p25_literal_2043923[p25_res7__320] ^ p25_array_index_2048332 ^ p26_array_index_2048518_comb ^ p25_array_index_2048383 ^ p25_array_index_2048351 ^ p25_literal_2043914[p25_array_index_2048336] ^ p25_literal_2043912[p25_array_index_2048337] ^ p25_literal_2043910[p25_array_index_2048354] ^ p25_array_index_2048339;
  assign p26_array_index_2048578_comb = p25_literal_2043918[p26_res7__328_comb];
  assign p26_array_index_2048579_comb = p25_literal_2043920[p25_res7__326];
  assign p26_res7__338_comb = p25_literal_2043910[p26_res7__336_comb] ^ p25_literal_2043912[p26_res7__334_comb] ^ p25_literal_2043914[p26_res7__332_comb] ^ p25_literal_2043916[p26_res7__330_comb] ^ p26_array_index_2048578_comb ^ p26_array_index_2048579_comb ^ p25_res7__324 ^ p25_literal_2043923[p25_res7__322] ^ p25_res7__320 ^ p26_array_index_2048531_comb ^ p25_array_index_2048397 ^ p25_array_index_2048368 ^ p25_literal_2043914[p25_array_index_2048335] ^ p25_literal_2043912[p25_array_index_2048336] ^ p25_literal_2043910[p25_array_index_2048337] ^ p25_array_index_2048354;
  assign p26_array_index_2048590_comb = p25_literal_2043920[p26_res7__328_comb];
  assign p26_res7__340_comb = p25_literal_2043910[p26_res7__338_comb] ^ p25_literal_2043912[p26_res7__336_comb] ^ p25_literal_2043914[p26_res7__334_comb] ^ p25_literal_2043916[p26_res7__332_comb] ^ p25_literal_2043918[p26_res7__330_comb] ^ p26_array_index_2048590_comb ^ p25_res7__326 ^ p25_literal_2043923[p25_res7__324] ^ p25_res7__322 ^ p26_array_index_2048544_comb ^ p26_array_index_2048517_comb ^ p25_array_index_2048382 ^ p25_array_index_2048350 ^ p25_literal_2043912[p25_array_index_2048335] ^ p25_literal_2043910[p25_array_index_2048336] ^ p25_array_index_2048337;

  // Registers for pipe stage 26:
  reg [127:0] p26_encoded;
  reg [127:0] p26_bit_slice_2043893;
  reg [127:0] p26_bit_slice_2044018;
  reg [127:0] p26_k3;
  reg [127:0] p26_k2;
  reg [127:0] p26_xor_2047836;
  reg [127:0] p26_xor_2048316;
  reg [7:0] p26_array_index_2048332;
  reg [7:0] p26_array_index_2048333;
  reg [7:0] p26_array_index_2048334;
  reg [7:0] p26_array_index_2048335;
  reg [7:0] p26_array_index_2048336;
  reg [7:0] p26_array_index_2048348;
  reg [7:0] p26_array_index_2048349;
  reg [7:0] p26_res7__320;
  reg [7:0] p26_array_index_2048365;
  reg [7:0] p26_array_index_2048366;
  reg [7:0] p26_array_index_2048367;
  reg [7:0] p26_res7__322;
  reg [7:0] p26_array_index_2048380;
  reg [7:0] p26_array_index_2048381;
  reg [7:0] p26_res7__324;
  reg [7:0] p26_array_index_2048394;
  reg [7:0] p26_array_index_2048395;
  reg [7:0] p26_array_index_2048396;
  reg [7:0] p26_res7__326;
  reg [7:0] p26_array_index_2048515;
  reg [7:0] p26_array_index_2048516;
  reg [7:0] p26_res7__328;
  reg [7:0] p26_array_index_2048528;
  reg [7:0] p26_array_index_2048529;
  reg [7:0] p26_array_index_2048530;
  reg [7:0] p26_res7__330;
  reg [7:0] p26_array_index_2048542;
  reg [7:0] p26_array_index_2048543;
  reg [7:0] p26_res7__332;
  reg [7:0] p26_array_index_2048554;
  reg [7:0] p26_array_index_2048555;
  reg [7:0] p26_array_index_2048556;
  reg [7:0] p26_res7__334;
  reg [7:0] p26_array_index_2048567;
  reg [7:0] p26_array_index_2048568;
  reg [7:0] p26_res7__336;
  reg [7:0] p26_array_index_2048578;
  reg [7:0] p26_array_index_2048579;
  reg [7:0] p26_res7__338;
  reg [7:0] p26_array_index_2048590;
  reg [7:0] p26_res7__340;
  reg [7:0] p27_literal_2043896[256];
  reg [7:0] p27_literal_2043910[256];
  reg [7:0] p27_literal_2043912[256];
  reg [7:0] p27_literal_2043914[256];
  reg [7:0] p27_literal_2043916[256];
  reg [7:0] p27_literal_2043918[256];
  reg [7:0] p27_literal_2043920[256];
  reg [7:0] p27_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p26_encoded <= p25_encoded;
    p26_bit_slice_2043893 <= p25_bit_slice_2043893;
    p26_bit_slice_2044018 <= p25_bit_slice_2044018;
    p26_k3 <= p25_k3;
    p26_k2 <= p25_k2;
    p26_xor_2047836 <= p25_xor_2047836;
    p26_xor_2048316 <= p25_xor_2048316;
    p26_array_index_2048332 <= p25_array_index_2048332;
    p26_array_index_2048333 <= p25_array_index_2048333;
    p26_array_index_2048334 <= p25_array_index_2048334;
    p26_array_index_2048335 <= p25_array_index_2048335;
    p26_array_index_2048336 <= p25_array_index_2048336;
    p26_array_index_2048348 <= p25_array_index_2048348;
    p26_array_index_2048349 <= p25_array_index_2048349;
    p26_res7__320 <= p25_res7__320;
    p26_array_index_2048365 <= p25_array_index_2048365;
    p26_array_index_2048366 <= p25_array_index_2048366;
    p26_array_index_2048367 <= p25_array_index_2048367;
    p26_res7__322 <= p25_res7__322;
    p26_array_index_2048380 <= p25_array_index_2048380;
    p26_array_index_2048381 <= p25_array_index_2048381;
    p26_res7__324 <= p25_res7__324;
    p26_array_index_2048394 <= p25_array_index_2048394;
    p26_array_index_2048395 <= p25_array_index_2048395;
    p26_array_index_2048396 <= p25_array_index_2048396;
    p26_res7__326 <= p25_res7__326;
    p26_array_index_2048515 <= p26_array_index_2048515_comb;
    p26_array_index_2048516 <= p26_array_index_2048516_comb;
    p26_res7__328 <= p26_res7__328_comb;
    p26_array_index_2048528 <= p26_array_index_2048528_comb;
    p26_array_index_2048529 <= p26_array_index_2048529_comb;
    p26_array_index_2048530 <= p26_array_index_2048530_comb;
    p26_res7__330 <= p26_res7__330_comb;
    p26_array_index_2048542 <= p26_array_index_2048542_comb;
    p26_array_index_2048543 <= p26_array_index_2048543_comb;
    p26_res7__332 <= p26_res7__332_comb;
    p26_array_index_2048554 <= p26_array_index_2048554_comb;
    p26_array_index_2048555 <= p26_array_index_2048555_comb;
    p26_array_index_2048556 <= p26_array_index_2048556_comb;
    p26_res7__334 <= p26_res7__334_comb;
    p26_array_index_2048567 <= p26_array_index_2048567_comb;
    p26_array_index_2048568 <= p26_array_index_2048568_comb;
    p26_res7__336 <= p26_res7__336_comb;
    p26_array_index_2048578 <= p26_array_index_2048578_comb;
    p26_array_index_2048579 <= p26_array_index_2048579_comb;
    p26_res7__338 <= p26_res7__338_comb;
    p26_array_index_2048590 <= p26_array_index_2048590_comb;
    p26_res7__340 <= p26_res7__340_comb;
    p27_literal_2043896 <= p26_literal_2043896;
    p27_literal_2043910 <= p26_literal_2043910;
    p27_literal_2043912 <= p26_literal_2043912;
    p27_literal_2043914 <= p26_literal_2043914;
    p27_literal_2043916 <= p26_literal_2043916;
    p27_literal_2043918 <= p26_literal_2043918;
    p27_literal_2043920 <= p26_literal_2043920;
    p27_literal_2043923 <= p26_literal_2043923;
  end

  // ===== Pipe stage 27:
  wire [7:0] p27_array_index_2048712_comb;
  wire [7:0] p27_res7__342_comb;
  wire [7:0] p27_res7__344_comb;
  wire [7:0] p27_res7__346_comb;
  wire [7:0] p27_res7__348_comb;
  wire [7:0] p27_res7__350_comb;
  wire [127:0] p27_res__10_comb;
  wire [127:0] p27_xor_2048752_comb;
  wire [127:0] p27_addedKey__43_comb;
  wire [7:0] p27_array_index_2048768_comb;
  wire [7:0] p27_array_index_2048769_comb;
  wire [7:0] p27_array_index_2048770_comb;
  wire [7:0] p27_array_index_2048771_comb;
  wire [7:0] p27_array_index_2048772_comb;
  wire [7:0] p27_array_index_2048773_comb;
  wire [7:0] p27_array_index_2048775_comb;
  wire [7:0] p27_array_index_2048777_comb;
  wire [7:0] p27_array_index_2048778_comb;
  wire [7:0] p27_array_index_2048779_comb;
  wire [7:0] p27_array_index_2048780_comb;
  wire [7:0] p27_array_index_2048781_comb;
  wire [7:0] p27_array_index_2048782_comb;
  wire [7:0] p27_array_index_2048784_comb;
  wire [7:0] p27_array_index_2048785_comb;
  wire [7:0] p27_array_index_2048786_comb;
  wire [7:0] p27_array_index_2048787_comb;
  wire [7:0] p27_array_index_2048788_comb;
  wire [7:0] p27_array_index_2048789_comb;
  wire [7:0] p27_array_index_2048790_comb;
  wire [7:0] p27_array_index_2048792_comb;
  wire [7:0] p27_res7__352_comb;
  assign p27_array_index_2048712_comb = p26_literal_2043920[p26_res7__330];
  assign p27_res7__342_comb = p26_literal_2043910[p26_res7__340] ^ p26_literal_2043912[p26_res7__338] ^ p26_literal_2043914[p26_res7__336] ^ p26_literal_2043916[p26_res7__334] ^ p26_literal_2043918[p26_res7__332] ^ p27_array_index_2048712_comb ^ p26_res7__328 ^ p26_literal_2043923[p26_res7__326] ^ p26_res7__324 ^ p26_array_index_2048556 ^ p26_array_index_2048530 ^ p26_array_index_2048396 ^ p26_array_index_2048367 ^ p26_literal_2043912[p26_array_index_2048334] ^ p26_literal_2043910[p26_array_index_2048335] ^ p26_array_index_2048336;
  assign p27_res7__344_comb = p26_literal_2043910[p27_res7__342_comb] ^ p26_literal_2043912[p26_res7__340] ^ p26_literal_2043914[p26_res7__338] ^ p26_literal_2043916[p26_res7__336] ^ p26_literal_2043918[p26_res7__334] ^ p26_literal_2043920[p26_res7__332] ^ p26_res7__330 ^ p26_literal_2043923[p26_res7__328] ^ p26_res7__326 ^ p26_array_index_2048568 ^ p26_array_index_2048543 ^ p26_array_index_2048516 ^ p26_array_index_2048381 ^ p26_array_index_2048349 ^ p26_literal_2043910[p26_array_index_2048334] ^ p26_array_index_2048335;
  assign p27_res7__346_comb = p26_literal_2043910[p27_res7__344_comb] ^ p26_literal_2043912[p27_res7__342_comb] ^ p26_literal_2043914[p26_res7__340] ^ p26_literal_2043916[p26_res7__338] ^ p26_literal_2043918[p26_res7__336] ^ p26_literal_2043920[p26_res7__334] ^ p26_res7__332 ^ p26_literal_2043923[p26_res7__330] ^ p26_res7__328 ^ p26_array_index_2048579 ^ p26_array_index_2048555 ^ p26_array_index_2048529 ^ p26_array_index_2048395 ^ p26_array_index_2048366 ^ p26_literal_2043910[p26_array_index_2048333] ^ p26_array_index_2048334;
  assign p27_res7__348_comb = p26_literal_2043910[p27_res7__346_comb] ^ p26_literal_2043912[p27_res7__344_comb] ^ p26_literal_2043914[p27_res7__342_comb] ^ p26_literal_2043916[p26_res7__340] ^ p26_literal_2043918[p26_res7__338] ^ p26_literal_2043920[p26_res7__336] ^ p26_res7__334 ^ p26_literal_2043923[p26_res7__332] ^ p26_res7__330 ^ p26_array_index_2048590 ^ p26_array_index_2048567 ^ p26_array_index_2048542 ^ p26_array_index_2048515 ^ p26_array_index_2048380 ^ p26_array_index_2048348 ^ p26_array_index_2048333;
  assign p27_res7__350_comb = p26_literal_2043910[p27_res7__348_comb] ^ p26_literal_2043912[p27_res7__346_comb] ^ p26_literal_2043914[p27_res7__344_comb] ^ p26_literal_2043916[p27_res7__342_comb] ^ p26_literal_2043918[p26_res7__340] ^ p26_literal_2043920[p26_res7__338] ^ p26_res7__336 ^ p26_literal_2043923[p26_res7__334] ^ p26_res7__332 ^ p27_array_index_2048712_comb ^ p26_array_index_2048578 ^ p26_array_index_2048554 ^ p26_array_index_2048528 ^ p26_array_index_2048394 ^ p26_array_index_2048365 ^ p26_array_index_2048332;
  assign p27_res__10_comb = {p27_res7__350_comb, p27_res7__348_comb, p27_res7__346_comb, p27_res7__344_comb, p27_res7__342_comb, p26_res7__340, p26_res7__338, p26_res7__336, p26_res7__334, p26_res7__332, p26_res7__330, p26_res7__328, p26_res7__326, p26_res7__324, p26_res7__322, p26_res7__320};
  assign p27_xor_2048752_comb = p27_res__10_comb ^ p26_xor_2047836;
  assign p27_addedKey__43_comb = p27_xor_2048752_comb ^ 128'h8d94_2d1d_95e6_7d2c_1a67_10c0_d5ff_3f0c;
  assign p27_array_index_2048768_comb = p26_literal_2043896[p27_addedKey__43_comb[127:120]];
  assign p27_array_index_2048769_comb = p26_literal_2043896[p27_addedKey__43_comb[119:112]];
  assign p27_array_index_2048770_comb = p26_literal_2043896[p27_addedKey__43_comb[111:104]];
  assign p27_array_index_2048771_comb = p26_literal_2043896[p27_addedKey__43_comb[103:96]];
  assign p27_array_index_2048772_comb = p26_literal_2043896[p27_addedKey__43_comb[95:88]];
  assign p27_array_index_2048773_comb = p26_literal_2043896[p27_addedKey__43_comb[87:80]];
  assign p27_array_index_2048775_comb = p26_literal_2043896[p27_addedKey__43_comb[71:64]];
  assign p27_array_index_2048777_comb = p26_literal_2043896[p27_addedKey__43_comb[55:48]];
  assign p27_array_index_2048778_comb = p26_literal_2043896[p27_addedKey__43_comb[47:40]];
  assign p27_array_index_2048779_comb = p26_literal_2043896[p27_addedKey__43_comb[39:32]];
  assign p27_array_index_2048780_comb = p26_literal_2043896[p27_addedKey__43_comb[31:24]];
  assign p27_array_index_2048781_comb = p26_literal_2043896[p27_addedKey__43_comb[23:16]];
  assign p27_array_index_2048782_comb = p26_literal_2043896[p27_addedKey__43_comb[15:8]];
  assign p27_array_index_2048784_comb = p26_literal_2043910[p27_array_index_2048768_comb];
  assign p27_array_index_2048785_comb = p26_literal_2043912[p27_array_index_2048769_comb];
  assign p27_array_index_2048786_comb = p26_literal_2043914[p27_array_index_2048770_comb];
  assign p27_array_index_2048787_comb = p26_literal_2043916[p27_array_index_2048771_comb];
  assign p27_array_index_2048788_comb = p26_literal_2043918[p27_array_index_2048772_comb];
  assign p27_array_index_2048789_comb = p26_literal_2043920[p27_array_index_2048773_comb];
  assign p27_array_index_2048790_comb = p26_literal_2043896[p27_addedKey__43_comb[79:72]];
  assign p27_array_index_2048792_comb = p26_literal_2043896[p27_addedKey__43_comb[63:56]];
  assign p27_res7__352_comb = p27_array_index_2048784_comb ^ p27_array_index_2048785_comb ^ p27_array_index_2048786_comb ^ p27_array_index_2048787_comb ^ p27_array_index_2048788_comb ^ p27_array_index_2048789_comb ^ p27_array_index_2048790_comb ^ p26_literal_2043923[p27_array_index_2048775_comb] ^ p27_array_index_2048792_comb ^ p26_literal_2043920[p27_array_index_2048777_comb] ^ p26_literal_2043918[p27_array_index_2048778_comb] ^ p26_literal_2043916[p27_array_index_2048779_comb] ^ p26_literal_2043914[p27_array_index_2048780_comb] ^ p26_literal_2043912[p27_array_index_2048781_comb] ^ p26_literal_2043910[p27_array_index_2048782_comb] ^ p26_literal_2043896[p27_addedKey__43_comb[7:0]];

  // Registers for pipe stage 27:
  reg [127:0] p27_encoded;
  reg [127:0] p27_bit_slice_2043893;
  reg [127:0] p27_bit_slice_2044018;
  reg [127:0] p27_k3;
  reg [127:0] p27_k2;
  reg [127:0] p27_xor_2048316;
  reg [127:0] p27_xor_2048752;
  reg [7:0] p27_array_index_2048768;
  reg [7:0] p27_array_index_2048769;
  reg [7:0] p27_array_index_2048770;
  reg [7:0] p27_array_index_2048771;
  reg [7:0] p27_array_index_2048772;
  reg [7:0] p27_array_index_2048773;
  reg [7:0] p27_array_index_2048775;
  reg [7:0] p27_array_index_2048777;
  reg [7:0] p27_array_index_2048778;
  reg [7:0] p27_array_index_2048779;
  reg [7:0] p27_array_index_2048780;
  reg [7:0] p27_array_index_2048781;
  reg [7:0] p27_array_index_2048782;
  reg [7:0] p27_array_index_2048784;
  reg [7:0] p27_array_index_2048785;
  reg [7:0] p27_array_index_2048786;
  reg [7:0] p27_array_index_2048787;
  reg [7:0] p27_array_index_2048788;
  reg [7:0] p27_array_index_2048789;
  reg [7:0] p27_array_index_2048790;
  reg [7:0] p27_array_index_2048792;
  reg [7:0] p27_res7__352;
  reg [7:0] p28_literal_2043896[256];
  reg [7:0] p28_literal_2043910[256];
  reg [7:0] p28_literal_2043912[256];
  reg [7:0] p28_literal_2043914[256];
  reg [7:0] p28_literal_2043916[256];
  reg [7:0] p28_literal_2043918[256];
  reg [7:0] p28_literal_2043920[256];
  reg [7:0] p28_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p27_encoded <= p26_encoded;
    p27_bit_slice_2043893 <= p26_bit_slice_2043893;
    p27_bit_slice_2044018 <= p26_bit_slice_2044018;
    p27_k3 <= p26_k3;
    p27_k2 <= p26_k2;
    p27_xor_2048316 <= p26_xor_2048316;
    p27_xor_2048752 <= p27_xor_2048752_comb;
    p27_array_index_2048768 <= p27_array_index_2048768_comb;
    p27_array_index_2048769 <= p27_array_index_2048769_comb;
    p27_array_index_2048770 <= p27_array_index_2048770_comb;
    p27_array_index_2048771 <= p27_array_index_2048771_comb;
    p27_array_index_2048772 <= p27_array_index_2048772_comb;
    p27_array_index_2048773 <= p27_array_index_2048773_comb;
    p27_array_index_2048775 <= p27_array_index_2048775_comb;
    p27_array_index_2048777 <= p27_array_index_2048777_comb;
    p27_array_index_2048778 <= p27_array_index_2048778_comb;
    p27_array_index_2048779 <= p27_array_index_2048779_comb;
    p27_array_index_2048780 <= p27_array_index_2048780_comb;
    p27_array_index_2048781 <= p27_array_index_2048781_comb;
    p27_array_index_2048782 <= p27_array_index_2048782_comb;
    p27_array_index_2048784 <= p27_array_index_2048784_comb;
    p27_array_index_2048785 <= p27_array_index_2048785_comb;
    p27_array_index_2048786 <= p27_array_index_2048786_comb;
    p27_array_index_2048787 <= p27_array_index_2048787_comb;
    p27_array_index_2048788 <= p27_array_index_2048788_comb;
    p27_array_index_2048789 <= p27_array_index_2048789_comb;
    p27_array_index_2048790 <= p27_array_index_2048790_comb;
    p27_array_index_2048792 <= p27_array_index_2048792_comb;
    p27_res7__352 <= p27_res7__352_comb;
    p28_literal_2043896 <= p27_literal_2043896;
    p28_literal_2043910 <= p27_literal_2043910;
    p28_literal_2043912 <= p27_literal_2043912;
    p28_literal_2043914 <= p27_literal_2043914;
    p28_literal_2043916 <= p27_literal_2043916;
    p28_literal_2043918 <= p27_literal_2043918;
    p28_literal_2043920 <= p27_literal_2043920;
    p28_literal_2043923 <= p27_literal_2043923;
  end

  // ===== Pipe stage 28:
  wire [7:0] p28_array_index_2048875_comb;
  wire [7:0] p28_array_index_2048876_comb;
  wire [7:0] p28_array_index_2048877_comb;
  wire [7:0] p28_array_index_2048878_comb;
  wire [7:0] p28_array_index_2048879_comb;
  wire [7:0] p28_array_index_2048880_comb;
  wire [7:0] p28_res7__354_comb;
  wire [7:0] p28_array_index_2048890_comb;
  wire [7:0] p28_array_index_2048891_comb;
  wire [7:0] p28_array_index_2048892_comb;
  wire [7:0] p28_array_index_2048893_comb;
  wire [7:0] p28_array_index_2048894_comb;
  wire [7:0] p28_res7__356_comb;
  wire [7:0] p28_array_index_2048904_comb;
  wire [7:0] p28_array_index_2048905_comb;
  wire [7:0] p28_array_index_2048906_comb;
  wire [7:0] p28_array_index_2048907_comb;
  wire [7:0] p28_array_index_2048908_comb;
  wire [7:0] p28_res7__358_comb;
  wire [7:0] p28_array_index_2048919_comb;
  wire [7:0] p28_array_index_2048920_comb;
  wire [7:0] p28_array_index_2048921_comb;
  wire [7:0] p28_array_index_2048922_comb;
  wire [7:0] p28_res7__360_comb;
  wire [7:0] p28_array_index_2048932_comb;
  wire [7:0] p28_array_index_2048933_comb;
  wire [7:0] p28_array_index_2048934_comb;
  wire [7:0] p28_array_index_2048935_comb;
  wire [7:0] p28_res7__362_comb;
  wire [7:0] p28_array_index_2048946_comb;
  wire [7:0] p28_array_index_2048947_comb;
  wire [7:0] p28_array_index_2048948_comb;
  wire [7:0] p28_res7__364_comb;
  wire [7:0] p28_array_index_2048958_comb;
  wire [7:0] p28_array_index_2048959_comb;
  wire [7:0] p28_array_index_2048960_comb;
  wire [7:0] p28_res7__366_comb;
  assign p28_array_index_2048875_comb = p27_literal_2043910[p27_res7__352];
  assign p28_array_index_2048876_comb = p27_literal_2043912[p27_array_index_2048768];
  assign p28_array_index_2048877_comb = p27_literal_2043914[p27_array_index_2048769];
  assign p28_array_index_2048878_comb = p27_literal_2043916[p27_array_index_2048770];
  assign p28_array_index_2048879_comb = p27_literal_2043918[p27_array_index_2048771];
  assign p28_array_index_2048880_comb = p27_literal_2043920[p27_array_index_2048772];
  assign p28_res7__354_comb = p28_array_index_2048875_comb ^ p28_array_index_2048876_comb ^ p28_array_index_2048877_comb ^ p28_array_index_2048878_comb ^ p28_array_index_2048879_comb ^ p28_array_index_2048880_comb ^ p27_array_index_2048773 ^ p27_literal_2043923[p27_array_index_2048790] ^ p27_array_index_2048775 ^ p27_literal_2043920[p27_array_index_2048792] ^ p27_literal_2043918[p27_array_index_2048777] ^ p27_literal_2043916[p27_array_index_2048778] ^ p27_literal_2043914[p27_array_index_2048779] ^ p27_literal_2043912[p27_array_index_2048780] ^ p27_literal_2043910[p27_array_index_2048781] ^ p27_array_index_2048782;
  assign p28_array_index_2048890_comb = p27_literal_2043912[p27_res7__352];
  assign p28_array_index_2048891_comb = p27_literal_2043914[p27_array_index_2048768];
  assign p28_array_index_2048892_comb = p27_literal_2043916[p27_array_index_2048769];
  assign p28_array_index_2048893_comb = p27_literal_2043918[p27_array_index_2048770];
  assign p28_array_index_2048894_comb = p27_literal_2043920[p27_array_index_2048771];
  assign p28_res7__356_comb = p27_literal_2043910[p28_res7__354_comb] ^ p28_array_index_2048890_comb ^ p28_array_index_2048891_comb ^ p28_array_index_2048892_comb ^ p28_array_index_2048893_comb ^ p28_array_index_2048894_comb ^ p27_array_index_2048772 ^ p27_literal_2043923[p27_array_index_2048773] ^ p27_array_index_2048790 ^ p27_literal_2043920[p27_array_index_2048775] ^ p27_literal_2043918[p27_array_index_2048792] ^ p27_literal_2043916[p27_array_index_2048777] ^ p27_literal_2043914[p27_array_index_2048778] ^ p27_literal_2043912[p27_array_index_2048779] ^ p27_literal_2043910[p27_array_index_2048780] ^ p27_array_index_2048781;
  assign p28_array_index_2048904_comb = p27_literal_2043912[p28_res7__354_comb];
  assign p28_array_index_2048905_comb = p27_literal_2043914[p27_res7__352];
  assign p28_array_index_2048906_comb = p27_literal_2043916[p27_array_index_2048768];
  assign p28_array_index_2048907_comb = p27_literal_2043918[p27_array_index_2048769];
  assign p28_array_index_2048908_comb = p27_literal_2043920[p27_array_index_2048770];
  assign p28_res7__358_comb = p27_literal_2043910[p28_res7__356_comb] ^ p28_array_index_2048904_comb ^ p28_array_index_2048905_comb ^ p28_array_index_2048906_comb ^ p28_array_index_2048907_comb ^ p28_array_index_2048908_comb ^ p27_array_index_2048771 ^ p27_literal_2043923[p27_array_index_2048772] ^ p27_array_index_2048773 ^ p27_literal_2043920[p27_array_index_2048790] ^ p27_literal_2043918[p27_array_index_2048775] ^ p27_literal_2043916[p27_array_index_2048792] ^ p27_literal_2043914[p27_array_index_2048777] ^ p27_literal_2043912[p27_array_index_2048778] ^ p27_literal_2043910[p27_array_index_2048779] ^ p27_array_index_2048780;
  assign p28_array_index_2048919_comb = p27_literal_2043914[p28_res7__354_comb];
  assign p28_array_index_2048920_comb = p27_literal_2043916[p27_res7__352];
  assign p28_array_index_2048921_comb = p27_literal_2043918[p27_array_index_2048768];
  assign p28_array_index_2048922_comb = p27_literal_2043920[p27_array_index_2048769];
  assign p28_res7__360_comb = p27_literal_2043910[p28_res7__358_comb] ^ p27_literal_2043912[p28_res7__356_comb] ^ p28_array_index_2048919_comb ^ p28_array_index_2048920_comb ^ p28_array_index_2048921_comb ^ p28_array_index_2048922_comb ^ p27_array_index_2048770 ^ p27_literal_2043923[p27_array_index_2048771] ^ p27_array_index_2048772 ^ p27_array_index_2048789 ^ p27_literal_2043918[p27_array_index_2048790] ^ p27_literal_2043916[p27_array_index_2048775] ^ p27_literal_2043914[p27_array_index_2048792] ^ p27_literal_2043912[p27_array_index_2048777] ^ p27_literal_2043910[p27_array_index_2048778] ^ p27_array_index_2048779;
  assign p28_array_index_2048932_comb = p27_literal_2043914[p28_res7__356_comb];
  assign p28_array_index_2048933_comb = p27_literal_2043916[p28_res7__354_comb];
  assign p28_array_index_2048934_comb = p27_literal_2043918[p27_res7__352];
  assign p28_array_index_2048935_comb = p27_literal_2043920[p27_array_index_2048768];
  assign p28_res7__362_comb = p27_literal_2043910[p28_res7__360_comb] ^ p27_literal_2043912[p28_res7__358_comb] ^ p28_array_index_2048932_comb ^ p28_array_index_2048933_comb ^ p28_array_index_2048934_comb ^ p28_array_index_2048935_comb ^ p27_array_index_2048769 ^ p27_literal_2043923[p27_array_index_2048770] ^ p27_array_index_2048771 ^ p28_array_index_2048880_comb ^ p27_literal_2043918[p27_array_index_2048773] ^ p27_literal_2043916[p27_array_index_2048790] ^ p27_literal_2043914[p27_array_index_2048775] ^ p27_literal_2043912[p27_array_index_2048792] ^ p27_literal_2043910[p27_array_index_2048777] ^ p27_array_index_2048778;
  assign p28_array_index_2048946_comb = p27_literal_2043916[p28_res7__356_comb];
  assign p28_array_index_2048947_comb = p27_literal_2043918[p28_res7__354_comb];
  assign p28_array_index_2048948_comb = p27_literal_2043920[p27_res7__352];
  assign p28_res7__364_comb = p27_literal_2043910[p28_res7__362_comb] ^ p27_literal_2043912[p28_res7__360_comb] ^ p27_literal_2043914[p28_res7__358_comb] ^ p28_array_index_2048946_comb ^ p28_array_index_2048947_comb ^ p28_array_index_2048948_comb ^ p27_array_index_2048768 ^ p27_literal_2043923[p27_array_index_2048769] ^ p27_array_index_2048770 ^ p28_array_index_2048894_comb ^ p27_array_index_2048788 ^ p27_literal_2043916[p27_array_index_2048773] ^ p27_literal_2043914[p27_array_index_2048790] ^ p27_literal_2043912[p27_array_index_2048775] ^ p27_literal_2043910[p27_array_index_2048792] ^ p27_array_index_2048777;
  assign p28_array_index_2048958_comb = p27_literal_2043916[p28_res7__358_comb];
  assign p28_array_index_2048959_comb = p27_literal_2043918[p28_res7__356_comb];
  assign p28_array_index_2048960_comb = p27_literal_2043920[p28_res7__354_comb];
  assign p28_res7__366_comb = p27_literal_2043910[p28_res7__364_comb] ^ p27_literal_2043912[p28_res7__362_comb] ^ p27_literal_2043914[p28_res7__360_comb] ^ p28_array_index_2048958_comb ^ p28_array_index_2048959_comb ^ p28_array_index_2048960_comb ^ p27_res7__352 ^ p27_literal_2043923[p27_array_index_2048768] ^ p27_array_index_2048769 ^ p28_array_index_2048908_comb ^ p28_array_index_2048879_comb ^ p27_literal_2043916[p27_array_index_2048772] ^ p27_literal_2043914[p27_array_index_2048773] ^ p27_literal_2043912[p27_array_index_2048790] ^ p27_literal_2043910[p27_array_index_2048775] ^ p27_array_index_2048792;

  // Registers for pipe stage 28:
  reg [127:0] p28_encoded;
  reg [127:0] p28_bit_slice_2043893;
  reg [127:0] p28_bit_slice_2044018;
  reg [127:0] p28_k3;
  reg [127:0] p28_k2;
  reg [127:0] p28_xor_2048316;
  reg [127:0] p28_xor_2048752;
  reg [7:0] p28_array_index_2048768;
  reg [7:0] p28_array_index_2048769;
  reg [7:0] p28_array_index_2048770;
  reg [7:0] p28_array_index_2048771;
  reg [7:0] p28_array_index_2048772;
  reg [7:0] p28_array_index_2048773;
  reg [7:0] p28_array_index_2048775;
  reg [7:0] p28_array_index_2048784;
  reg [7:0] p28_array_index_2048785;
  reg [7:0] p28_array_index_2048786;
  reg [7:0] p28_array_index_2048787;
  reg [7:0] p28_array_index_2048790;
  reg [7:0] p28_res7__352;
  reg [7:0] p28_array_index_2048875;
  reg [7:0] p28_array_index_2048876;
  reg [7:0] p28_array_index_2048877;
  reg [7:0] p28_array_index_2048878;
  reg [7:0] p28_res7__354;
  reg [7:0] p28_array_index_2048890;
  reg [7:0] p28_array_index_2048891;
  reg [7:0] p28_array_index_2048892;
  reg [7:0] p28_array_index_2048893;
  reg [7:0] p28_res7__356;
  reg [7:0] p28_array_index_2048904;
  reg [7:0] p28_array_index_2048905;
  reg [7:0] p28_array_index_2048906;
  reg [7:0] p28_array_index_2048907;
  reg [7:0] p28_res7__358;
  reg [7:0] p28_array_index_2048919;
  reg [7:0] p28_array_index_2048920;
  reg [7:0] p28_array_index_2048921;
  reg [7:0] p28_array_index_2048922;
  reg [7:0] p28_res7__360;
  reg [7:0] p28_array_index_2048932;
  reg [7:0] p28_array_index_2048933;
  reg [7:0] p28_array_index_2048934;
  reg [7:0] p28_array_index_2048935;
  reg [7:0] p28_res7__362;
  reg [7:0] p28_array_index_2048946;
  reg [7:0] p28_array_index_2048947;
  reg [7:0] p28_array_index_2048948;
  reg [7:0] p28_res7__364;
  reg [7:0] p28_array_index_2048958;
  reg [7:0] p28_array_index_2048959;
  reg [7:0] p28_array_index_2048960;
  reg [7:0] p28_res7__366;
  reg [7:0] p29_literal_2043896[256];
  reg [7:0] p29_literal_2043910[256];
  reg [7:0] p29_literal_2043912[256];
  reg [7:0] p29_literal_2043914[256];
  reg [7:0] p29_literal_2043916[256];
  reg [7:0] p29_literal_2043918[256];
  reg [7:0] p29_literal_2043920[256];
  reg [7:0] p29_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p28_encoded <= p27_encoded;
    p28_bit_slice_2043893 <= p27_bit_slice_2043893;
    p28_bit_slice_2044018 <= p27_bit_slice_2044018;
    p28_k3 <= p27_k3;
    p28_k2 <= p27_k2;
    p28_xor_2048316 <= p27_xor_2048316;
    p28_xor_2048752 <= p27_xor_2048752;
    p28_array_index_2048768 <= p27_array_index_2048768;
    p28_array_index_2048769 <= p27_array_index_2048769;
    p28_array_index_2048770 <= p27_array_index_2048770;
    p28_array_index_2048771 <= p27_array_index_2048771;
    p28_array_index_2048772 <= p27_array_index_2048772;
    p28_array_index_2048773 <= p27_array_index_2048773;
    p28_array_index_2048775 <= p27_array_index_2048775;
    p28_array_index_2048784 <= p27_array_index_2048784;
    p28_array_index_2048785 <= p27_array_index_2048785;
    p28_array_index_2048786 <= p27_array_index_2048786;
    p28_array_index_2048787 <= p27_array_index_2048787;
    p28_array_index_2048790 <= p27_array_index_2048790;
    p28_res7__352 <= p27_res7__352;
    p28_array_index_2048875 <= p28_array_index_2048875_comb;
    p28_array_index_2048876 <= p28_array_index_2048876_comb;
    p28_array_index_2048877 <= p28_array_index_2048877_comb;
    p28_array_index_2048878 <= p28_array_index_2048878_comb;
    p28_res7__354 <= p28_res7__354_comb;
    p28_array_index_2048890 <= p28_array_index_2048890_comb;
    p28_array_index_2048891 <= p28_array_index_2048891_comb;
    p28_array_index_2048892 <= p28_array_index_2048892_comb;
    p28_array_index_2048893 <= p28_array_index_2048893_comb;
    p28_res7__356 <= p28_res7__356_comb;
    p28_array_index_2048904 <= p28_array_index_2048904_comb;
    p28_array_index_2048905 <= p28_array_index_2048905_comb;
    p28_array_index_2048906 <= p28_array_index_2048906_comb;
    p28_array_index_2048907 <= p28_array_index_2048907_comb;
    p28_res7__358 <= p28_res7__358_comb;
    p28_array_index_2048919 <= p28_array_index_2048919_comb;
    p28_array_index_2048920 <= p28_array_index_2048920_comb;
    p28_array_index_2048921 <= p28_array_index_2048921_comb;
    p28_array_index_2048922 <= p28_array_index_2048922_comb;
    p28_res7__360 <= p28_res7__360_comb;
    p28_array_index_2048932 <= p28_array_index_2048932_comb;
    p28_array_index_2048933 <= p28_array_index_2048933_comb;
    p28_array_index_2048934 <= p28_array_index_2048934_comb;
    p28_array_index_2048935 <= p28_array_index_2048935_comb;
    p28_res7__362 <= p28_res7__362_comb;
    p28_array_index_2048946 <= p28_array_index_2048946_comb;
    p28_array_index_2048947 <= p28_array_index_2048947_comb;
    p28_array_index_2048948 <= p28_array_index_2048948_comb;
    p28_res7__364 <= p28_res7__364_comb;
    p28_array_index_2048958 <= p28_array_index_2048958_comb;
    p28_array_index_2048959 <= p28_array_index_2048959_comb;
    p28_array_index_2048960 <= p28_array_index_2048960_comb;
    p28_res7__366 <= p28_res7__366_comb;
    p29_literal_2043896 <= p28_literal_2043896;
    p29_literal_2043910 <= p28_literal_2043910;
    p29_literal_2043912 <= p28_literal_2043912;
    p29_literal_2043914 <= p28_literal_2043914;
    p29_literal_2043916 <= p28_literal_2043916;
    p29_literal_2043918 <= p28_literal_2043918;
    p29_literal_2043920 <= p28_literal_2043920;
    p29_literal_2043923 <= p28_literal_2043923;
  end

  // ===== Pipe stage 29:
  wire [7:0] p29_array_index_2049093_comb;
  wire [7:0] p29_array_index_2049094_comb;
  wire [7:0] p29_res7__368_comb;
  wire [7:0] p29_array_index_2049104_comb;
  wire [7:0] p29_array_index_2049105_comb;
  wire [7:0] p29_res7__370_comb;
  wire [7:0] p29_array_index_2049116_comb;
  wire [7:0] p29_res7__372_comb;
  wire [7:0] p29_array_index_2049126_comb;
  wire [7:0] p29_res7__374_comb;
  wire [7:0] p29_res7__376_comb;
  wire [7:0] p29_res7__378_comb;
  wire [7:0] p29_res7__380_comb;
  assign p29_array_index_2049093_comb = p28_literal_2043918[p28_res7__358];
  assign p29_array_index_2049094_comb = p28_literal_2043920[p28_res7__356];
  assign p29_res7__368_comb = p28_literal_2043910[p28_res7__366] ^ p28_literal_2043912[p28_res7__364] ^ p28_literal_2043914[p28_res7__362] ^ p28_literal_2043916[p28_res7__360] ^ p29_array_index_2049093_comb ^ p29_array_index_2049094_comb ^ p28_res7__354 ^ p28_literal_2043923[p28_res7__352] ^ p28_array_index_2048768 ^ p28_array_index_2048922 ^ p28_array_index_2048893 ^ p28_array_index_2048787 ^ p28_literal_2043914[p28_array_index_2048772] ^ p28_literal_2043912[p28_array_index_2048773] ^ p28_literal_2043910[p28_array_index_2048790] ^ p28_array_index_2048775;
  assign p29_array_index_2049104_comb = p28_literal_2043918[p28_res7__360];
  assign p29_array_index_2049105_comb = p28_literal_2043920[p28_res7__358];
  assign p29_res7__370_comb = p28_literal_2043910[p29_res7__368_comb] ^ p28_literal_2043912[p28_res7__366] ^ p28_literal_2043914[p28_res7__364] ^ p28_literal_2043916[p28_res7__362] ^ p29_array_index_2049104_comb ^ p29_array_index_2049105_comb ^ p28_res7__356 ^ p28_literal_2043923[p28_res7__354] ^ p28_res7__352 ^ p28_array_index_2048935 ^ p28_array_index_2048907 ^ p28_array_index_2048878 ^ p28_literal_2043914[p28_array_index_2048771] ^ p28_literal_2043912[p28_array_index_2048772] ^ p28_literal_2043910[p28_array_index_2048773] ^ p28_array_index_2048790;
  assign p29_array_index_2049116_comb = p28_literal_2043920[p28_res7__360];
  assign p29_res7__372_comb = p28_literal_2043910[p29_res7__370_comb] ^ p28_literal_2043912[p29_res7__368_comb] ^ p28_literal_2043914[p28_res7__366] ^ p28_literal_2043916[p28_res7__364] ^ p28_literal_2043918[p28_res7__362] ^ p29_array_index_2049116_comb ^ p28_res7__358 ^ p28_literal_2043923[p28_res7__356] ^ p28_res7__354 ^ p28_array_index_2048948 ^ p28_array_index_2048921 ^ p28_array_index_2048892 ^ p28_array_index_2048786 ^ p28_literal_2043912[p28_array_index_2048771] ^ p28_literal_2043910[p28_array_index_2048772] ^ p28_array_index_2048773;
  assign p29_array_index_2049126_comb = p28_literal_2043920[p28_res7__362];
  assign p29_res7__374_comb = p28_literal_2043910[p29_res7__372_comb] ^ p28_literal_2043912[p29_res7__370_comb] ^ p28_literal_2043914[p29_res7__368_comb] ^ p28_literal_2043916[p28_res7__366] ^ p28_literal_2043918[p28_res7__364] ^ p29_array_index_2049126_comb ^ p28_res7__360 ^ p28_literal_2043923[p28_res7__358] ^ p28_res7__356 ^ p28_array_index_2048960 ^ p28_array_index_2048934 ^ p28_array_index_2048906 ^ p28_array_index_2048877 ^ p28_literal_2043912[p28_array_index_2048770] ^ p28_literal_2043910[p28_array_index_2048771] ^ p28_array_index_2048772;
  assign p29_res7__376_comb = p28_literal_2043910[p29_res7__374_comb] ^ p28_literal_2043912[p29_res7__372_comb] ^ p28_literal_2043914[p29_res7__370_comb] ^ p28_literal_2043916[p29_res7__368_comb] ^ p28_literal_2043918[p28_res7__366] ^ p28_literal_2043920[p28_res7__364] ^ p28_res7__362 ^ p28_literal_2043923[p28_res7__360] ^ p28_res7__358 ^ p29_array_index_2049094_comb ^ p28_array_index_2048947 ^ p28_array_index_2048920 ^ p28_array_index_2048891 ^ p28_array_index_2048785 ^ p28_literal_2043910[p28_array_index_2048770] ^ p28_array_index_2048771;
  assign p29_res7__378_comb = p28_literal_2043910[p29_res7__376_comb] ^ p28_literal_2043912[p29_res7__374_comb] ^ p28_literal_2043914[p29_res7__372_comb] ^ p28_literal_2043916[p29_res7__370_comb] ^ p28_literal_2043918[p29_res7__368_comb] ^ p28_literal_2043920[p28_res7__366] ^ p28_res7__364 ^ p28_literal_2043923[p28_res7__362] ^ p28_res7__360 ^ p29_array_index_2049105_comb ^ p28_array_index_2048959 ^ p28_array_index_2048933 ^ p28_array_index_2048905 ^ p28_array_index_2048876 ^ p28_literal_2043910[p28_array_index_2048769] ^ p28_array_index_2048770;
  assign p29_res7__380_comb = p28_literal_2043910[p29_res7__378_comb] ^ p28_literal_2043912[p29_res7__376_comb] ^ p28_literal_2043914[p29_res7__374_comb] ^ p28_literal_2043916[p29_res7__372_comb] ^ p28_literal_2043918[p29_res7__370_comb] ^ p28_literal_2043920[p29_res7__368_comb] ^ p28_res7__366 ^ p28_literal_2043923[p28_res7__364] ^ p28_res7__362 ^ p29_array_index_2049116_comb ^ p29_array_index_2049093_comb ^ p28_array_index_2048946 ^ p28_array_index_2048919 ^ p28_array_index_2048890 ^ p28_array_index_2048784 ^ p28_array_index_2048769;

  // Registers for pipe stage 29:
  reg [127:0] p29_encoded;
  reg [127:0] p29_bit_slice_2043893;
  reg [127:0] p29_bit_slice_2044018;
  reg [127:0] p29_k3;
  reg [127:0] p29_k2;
  reg [127:0] p29_xor_2048316;
  reg [127:0] p29_xor_2048752;
  reg [7:0] p29_array_index_2048768;
  reg [7:0] p29_res7__352;
  reg [7:0] p29_array_index_2048875;
  reg [7:0] p29_res7__354;
  reg [7:0] p29_res7__356;
  reg [7:0] p29_array_index_2048904;
  reg [7:0] p29_res7__358;
  reg [7:0] p29_res7__360;
  reg [7:0] p29_array_index_2048932;
  reg [7:0] p29_res7__362;
  reg [7:0] p29_res7__364;
  reg [7:0] p29_array_index_2048958;
  reg [7:0] p29_res7__366;
  reg [7:0] p29_res7__368;
  reg [7:0] p29_array_index_2049104;
  reg [7:0] p29_res7__370;
  reg [7:0] p29_res7__372;
  reg [7:0] p29_array_index_2049126;
  reg [7:0] p29_res7__374;
  reg [7:0] p29_res7__376;
  reg [7:0] p29_res7__378;
  reg [7:0] p29_res7__380;
  reg [7:0] p30_literal_2043896[256];
  reg [7:0] p30_literal_2043910[256];
  reg [7:0] p30_literal_2043912[256];
  reg [7:0] p30_literal_2043914[256];
  reg [7:0] p30_literal_2043916[256];
  reg [7:0] p30_literal_2043918[256];
  reg [7:0] p30_literal_2043920[256];
  reg [7:0] p30_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p29_encoded <= p28_encoded;
    p29_bit_slice_2043893 <= p28_bit_slice_2043893;
    p29_bit_slice_2044018 <= p28_bit_slice_2044018;
    p29_k3 <= p28_k3;
    p29_k2 <= p28_k2;
    p29_xor_2048316 <= p28_xor_2048316;
    p29_xor_2048752 <= p28_xor_2048752;
    p29_array_index_2048768 <= p28_array_index_2048768;
    p29_res7__352 <= p28_res7__352;
    p29_array_index_2048875 <= p28_array_index_2048875;
    p29_res7__354 <= p28_res7__354;
    p29_res7__356 <= p28_res7__356;
    p29_array_index_2048904 <= p28_array_index_2048904;
    p29_res7__358 <= p28_res7__358;
    p29_res7__360 <= p28_res7__360;
    p29_array_index_2048932 <= p28_array_index_2048932;
    p29_res7__362 <= p28_res7__362;
    p29_res7__364 <= p28_res7__364;
    p29_array_index_2048958 <= p28_array_index_2048958;
    p29_res7__366 <= p28_res7__366;
    p29_res7__368 <= p29_res7__368_comb;
    p29_array_index_2049104 <= p29_array_index_2049104_comb;
    p29_res7__370 <= p29_res7__370_comb;
    p29_res7__372 <= p29_res7__372_comb;
    p29_array_index_2049126 <= p29_array_index_2049126_comb;
    p29_res7__374 <= p29_res7__374_comb;
    p29_res7__376 <= p29_res7__376_comb;
    p29_res7__378 <= p29_res7__378_comb;
    p29_res7__380 <= p29_res7__380_comb;
    p30_literal_2043896 <= p29_literal_2043896;
    p30_literal_2043910 <= p29_literal_2043910;
    p30_literal_2043912 <= p29_literal_2043912;
    p30_literal_2043914 <= p29_literal_2043914;
    p30_literal_2043916 <= p29_literal_2043916;
    p30_literal_2043918 <= p29_literal_2043918;
    p30_literal_2043920 <= p29_literal_2043920;
    p30_literal_2043923 <= p29_literal_2043923;
  end

  // ===== Pipe stage 30:
  wire [7:0] p30_res7__382_comb;
  wire [127:0] p30_res__11_comb;
  wire [127:0] p30_xor_2049240_comb;
  wire [127:0] p30_addedKey__44_comb;
  wire [7:0] p30_array_index_2049256_comb;
  wire [7:0] p30_array_index_2049257_comb;
  wire [7:0] p30_array_index_2049258_comb;
  wire [7:0] p30_array_index_2049259_comb;
  wire [7:0] p30_array_index_2049260_comb;
  wire [7:0] p30_array_index_2049261_comb;
  wire [7:0] p30_array_index_2049263_comb;
  wire [7:0] p30_array_index_2049265_comb;
  wire [7:0] p30_array_index_2049266_comb;
  wire [7:0] p30_array_index_2049267_comb;
  wire [7:0] p30_array_index_2049268_comb;
  wire [7:0] p30_array_index_2049269_comb;
  wire [7:0] p30_array_index_2049270_comb;
  wire [7:0] p30_array_index_2049272_comb;
  wire [7:0] p30_array_index_2049273_comb;
  wire [7:0] p30_array_index_2049274_comb;
  wire [7:0] p30_array_index_2049275_comb;
  wire [7:0] p30_array_index_2049276_comb;
  wire [7:0] p30_array_index_2049277_comb;
  wire [7:0] p30_array_index_2049278_comb;
  wire [7:0] p30_array_index_2049280_comb;
  wire [7:0] p30_res7__384_comb;
  wire [7:0] p30_array_index_2049289_comb;
  wire [7:0] p30_array_index_2049290_comb;
  wire [7:0] p30_array_index_2049291_comb;
  wire [7:0] p30_array_index_2049292_comb;
  wire [7:0] p30_array_index_2049293_comb;
  wire [7:0] p30_array_index_2049294_comb;
  wire [7:0] p30_res7__386_comb;
  wire [7:0] p30_array_index_2049304_comb;
  wire [7:0] p30_array_index_2049305_comb;
  wire [7:0] p30_array_index_2049306_comb;
  wire [7:0] p30_array_index_2049307_comb;
  wire [7:0] p30_array_index_2049308_comb;
  wire [7:0] p30_res7__388_comb;
  wire [7:0] p30_array_index_2049318_comb;
  wire [7:0] p30_array_index_2049319_comb;
  wire [7:0] p30_array_index_2049320_comb;
  wire [7:0] p30_array_index_2049321_comb;
  wire [7:0] p30_array_index_2049322_comb;
  wire [7:0] p30_res7__390_comb;
  wire [7:0] p30_array_index_2049333_comb;
  wire [7:0] p30_array_index_2049334_comb;
  wire [7:0] p30_array_index_2049335_comb;
  wire [7:0] p30_array_index_2049336_comb;
  wire [7:0] p30_res7__392_comb;
  assign p30_res7__382_comb = p29_literal_2043910[p29_res7__380] ^ p29_literal_2043912[p29_res7__378] ^ p29_literal_2043914[p29_res7__376] ^ p29_literal_2043916[p29_res7__374] ^ p29_literal_2043918[p29_res7__372] ^ p29_literal_2043920[p29_res7__370] ^ p29_res7__368 ^ p29_literal_2043923[p29_res7__366] ^ p29_res7__364 ^ p29_array_index_2049126 ^ p29_array_index_2049104 ^ p29_array_index_2048958 ^ p29_array_index_2048932 ^ p29_array_index_2048904 ^ p29_array_index_2048875 ^ p29_array_index_2048768;
  assign p30_res__11_comb = {p30_res7__382_comb, p29_res7__380, p29_res7__378, p29_res7__376, p29_res7__374, p29_res7__372, p29_res7__370, p29_res7__368, p29_res7__366, p29_res7__364, p29_res7__362, p29_res7__360, p29_res7__358, p29_res7__356, p29_res7__354, p29_res7__352};
  assign p30_xor_2049240_comb = p30_res__11_comb ^ p29_xor_2048316;
  assign p30_addedKey__44_comb = p30_xor_2049240_comb ^ 128'he336_5b6f_f9ae_0794_4740_add0_087b_ab0d;
  assign p30_array_index_2049256_comb = p29_literal_2043896[p30_addedKey__44_comb[127:120]];
  assign p30_array_index_2049257_comb = p29_literal_2043896[p30_addedKey__44_comb[119:112]];
  assign p30_array_index_2049258_comb = p29_literal_2043896[p30_addedKey__44_comb[111:104]];
  assign p30_array_index_2049259_comb = p29_literal_2043896[p30_addedKey__44_comb[103:96]];
  assign p30_array_index_2049260_comb = p29_literal_2043896[p30_addedKey__44_comb[95:88]];
  assign p30_array_index_2049261_comb = p29_literal_2043896[p30_addedKey__44_comb[87:80]];
  assign p30_array_index_2049263_comb = p29_literal_2043896[p30_addedKey__44_comb[71:64]];
  assign p30_array_index_2049265_comb = p29_literal_2043896[p30_addedKey__44_comb[55:48]];
  assign p30_array_index_2049266_comb = p29_literal_2043896[p30_addedKey__44_comb[47:40]];
  assign p30_array_index_2049267_comb = p29_literal_2043896[p30_addedKey__44_comb[39:32]];
  assign p30_array_index_2049268_comb = p29_literal_2043896[p30_addedKey__44_comb[31:24]];
  assign p30_array_index_2049269_comb = p29_literal_2043896[p30_addedKey__44_comb[23:16]];
  assign p30_array_index_2049270_comb = p29_literal_2043896[p30_addedKey__44_comb[15:8]];
  assign p30_array_index_2049272_comb = p29_literal_2043910[p30_array_index_2049256_comb];
  assign p30_array_index_2049273_comb = p29_literal_2043912[p30_array_index_2049257_comb];
  assign p30_array_index_2049274_comb = p29_literal_2043914[p30_array_index_2049258_comb];
  assign p30_array_index_2049275_comb = p29_literal_2043916[p30_array_index_2049259_comb];
  assign p30_array_index_2049276_comb = p29_literal_2043918[p30_array_index_2049260_comb];
  assign p30_array_index_2049277_comb = p29_literal_2043920[p30_array_index_2049261_comb];
  assign p30_array_index_2049278_comb = p29_literal_2043896[p30_addedKey__44_comb[79:72]];
  assign p30_array_index_2049280_comb = p29_literal_2043896[p30_addedKey__44_comb[63:56]];
  assign p30_res7__384_comb = p30_array_index_2049272_comb ^ p30_array_index_2049273_comb ^ p30_array_index_2049274_comb ^ p30_array_index_2049275_comb ^ p30_array_index_2049276_comb ^ p30_array_index_2049277_comb ^ p30_array_index_2049278_comb ^ p29_literal_2043923[p30_array_index_2049263_comb] ^ p30_array_index_2049280_comb ^ p29_literal_2043920[p30_array_index_2049265_comb] ^ p29_literal_2043918[p30_array_index_2049266_comb] ^ p29_literal_2043916[p30_array_index_2049267_comb] ^ p29_literal_2043914[p30_array_index_2049268_comb] ^ p29_literal_2043912[p30_array_index_2049269_comb] ^ p29_literal_2043910[p30_array_index_2049270_comb] ^ p29_literal_2043896[p30_addedKey__44_comb[7:0]];
  assign p30_array_index_2049289_comb = p29_literal_2043910[p30_res7__384_comb];
  assign p30_array_index_2049290_comb = p29_literal_2043912[p30_array_index_2049256_comb];
  assign p30_array_index_2049291_comb = p29_literal_2043914[p30_array_index_2049257_comb];
  assign p30_array_index_2049292_comb = p29_literal_2043916[p30_array_index_2049258_comb];
  assign p30_array_index_2049293_comb = p29_literal_2043918[p30_array_index_2049259_comb];
  assign p30_array_index_2049294_comb = p29_literal_2043920[p30_array_index_2049260_comb];
  assign p30_res7__386_comb = p30_array_index_2049289_comb ^ p30_array_index_2049290_comb ^ p30_array_index_2049291_comb ^ p30_array_index_2049292_comb ^ p30_array_index_2049293_comb ^ p30_array_index_2049294_comb ^ p30_array_index_2049261_comb ^ p29_literal_2043923[p30_array_index_2049278_comb] ^ p30_array_index_2049263_comb ^ p29_literal_2043920[p30_array_index_2049280_comb] ^ p29_literal_2043918[p30_array_index_2049265_comb] ^ p29_literal_2043916[p30_array_index_2049266_comb] ^ p29_literal_2043914[p30_array_index_2049267_comb] ^ p29_literal_2043912[p30_array_index_2049268_comb] ^ p29_literal_2043910[p30_array_index_2049269_comb] ^ p30_array_index_2049270_comb;
  assign p30_array_index_2049304_comb = p29_literal_2043912[p30_res7__384_comb];
  assign p30_array_index_2049305_comb = p29_literal_2043914[p30_array_index_2049256_comb];
  assign p30_array_index_2049306_comb = p29_literal_2043916[p30_array_index_2049257_comb];
  assign p30_array_index_2049307_comb = p29_literal_2043918[p30_array_index_2049258_comb];
  assign p30_array_index_2049308_comb = p29_literal_2043920[p30_array_index_2049259_comb];
  assign p30_res7__388_comb = p29_literal_2043910[p30_res7__386_comb] ^ p30_array_index_2049304_comb ^ p30_array_index_2049305_comb ^ p30_array_index_2049306_comb ^ p30_array_index_2049307_comb ^ p30_array_index_2049308_comb ^ p30_array_index_2049260_comb ^ p29_literal_2043923[p30_array_index_2049261_comb] ^ p30_array_index_2049278_comb ^ p29_literal_2043920[p30_array_index_2049263_comb] ^ p29_literal_2043918[p30_array_index_2049280_comb] ^ p29_literal_2043916[p30_array_index_2049265_comb] ^ p29_literal_2043914[p30_array_index_2049266_comb] ^ p29_literal_2043912[p30_array_index_2049267_comb] ^ p29_literal_2043910[p30_array_index_2049268_comb] ^ p30_array_index_2049269_comb;
  assign p30_array_index_2049318_comb = p29_literal_2043912[p30_res7__386_comb];
  assign p30_array_index_2049319_comb = p29_literal_2043914[p30_res7__384_comb];
  assign p30_array_index_2049320_comb = p29_literal_2043916[p30_array_index_2049256_comb];
  assign p30_array_index_2049321_comb = p29_literal_2043918[p30_array_index_2049257_comb];
  assign p30_array_index_2049322_comb = p29_literal_2043920[p30_array_index_2049258_comb];
  assign p30_res7__390_comb = p29_literal_2043910[p30_res7__388_comb] ^ p30_array_index_2049318_comb ^ p30_array_index_2049319_comb ^ p30_array_index_2049320_comb ^ p30_array_index_2049321_comb ^ p30_array_index_2049322_comb ^ p30_array_index_2049259_comb ^ p29_literal_2043923[p30_array_index_2049260_comb] ^ p30_array_index_2049261_comb ^ p29_literal_2043920[p30_array_index_2049278_comb] ^ p29_literal_2043918[p30_array_index_2049263_comb] ^ p29_literal_2043916[p30_array_index_2049280_comb] ^ p29_literal_2043914[p30_array_index_2049265_comb] ^ p29_literal_2043912[p30_array_index_2049266_comb] ^ p29_literal_2043910[p30_array_index_2049267_comb] ^ p30_array_index_2049268_comb;
  assign p30_array_index_2049333_comb = p29_literal_2043914[p30_res7__386_comb];
  assign p30_array_index_2049334_comb = p29_literal_2043916[p30_res7__384_comb];
  assign p30_array_index_2049335_comb = p29_literal_2043918[p30_array_index_2049256_comb];
  assign p30_array_index_2049336_comb = p29_literal_2043920[p30_array_index_2049257_comb];
  assign p30_res7__392_comb = p29_literal_2043910[p30_res7__390_comb] ^ p29_literal_2043912[p30_res7__388_comb] ^ p30_array_index_2049333_comb ^ p30_array_index_2049334_comb ^ p30_array_index_2049335_comb ^ p30_array_index_2049336_comb ^ p30_array_index_2049258_comb ^ p29_literal_2043923[p30_array_index_2049259_comb] ^ p30_array_index_2049260_comb ^ p30_array_index_2049277_comb ^ p29_literal_2043918[p30_array_index_2049278_comb] ^ p29_literal_2043916[p30_array_index_2049263_comb] ^ p29_literal_2043914[p30_array_index_2049280_comb] ^ p29_literal_2043912[p30_array_index_2049265_comb] ^ p29_literal_2043910[p30_array_index_2049266_comb] ^ p30_array_index_2049267_comb;

  // Registers for pipe stage 30:
  reg [127:0] p30_encoded;
  reg [127:0] p30_bit_slice_2043893;
  reg [127:0] p30_bit_slice_2044018;
  reg [127:0] p30_k3;
  reg [127:0] p30_k2;
  reg [127:0] p30_xor_2048752;
  reg [127:0] p30_xor_2049240;
  reg [7:0] p30_array_index_2049256;
  reg [7:0] p30_array_index_2049257;
  reg [7:0] p30_array_index_2049258;
  reg [7:0] p30_array_index_2049259;
  reg [7:0] p30_array_index_2049260;
  reg [7:0] p30_array_index_2049261;
  reg [7:0] p30_array_index_2049263;
  reg [7:0] p30_array_index_2049265;
  reg [7:0] p30_array_index_2049266;
  reg [7:0] p30_array_index_2049272;
  reg [7:0] p30_array_index_2049273;
  reg [7:0] p30_array_index_2049274;
  reg [7:0] p30_array_index_2049275;
  reg [7:0] p30_array_index_2049276;
  reg [7:0] p30_array_index_2049278;
  reg [7:0] p30_array_index_2049280;
  reg [7:0] p30_res7__384;
  reg [7:0] p30_array_index_2049289;
  reg [7:0] p30_array_index_2049290;
  reg [7:0] p30_array_index_2049291;
  reg [7:0] p30_array_index_2049292;
  reg [7:0] p30_array_index_2049293;
  reg [7:0] p30_array_index_2049294;
  reg [7:0] p30_res7__386;
  reg [7:0] p30_array_index_2049304;
  reg [7:0] p30_array_index_2049305;
  reg [7:0] p30_array_index_2049306;
  reg [7:0] p30_array_index_2049307;
  reg [7:0] p30_array_index_2049308;
  reg [7:0] p30_res7__388;
  reg [7:0] p30_array_index_2049318;
  reg [7:0] p30_array_index_2049319;
  reg [7:0] p30_array_index_2049320;
  reg [7:0] p30_array_index_2049321;
  reg [7:0] p30_array_index_2049322;
  reg [7:0] p30_res7__390;
  reg [7:0] p30_array_index_2049333;
  reg [7:0] p30_array_index_2049334;
  reg [7:0] p30_array_index_2049335;
  reg [7:0] p30_array_index_2049336;
  reg [7:0] p30_res7__392;
  reg [7:0] p31_literal_2043896[256];
  reg [7:0] p31_literal_2043910[256];
  reg [7:0] p31_literal_2043912[256];
  reg [7:0] p31_literal_2043914[256];
  reg [7:0] p31_literal_2043916[256];
  reg [7:0] p31_literal_2043918[256];
  reg [7:0] p31_literal_2043920[256];
  reg [7:0] p31_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p30_encoded <= p29_encoded;
    p30_bit_slice_2043893 <= p29_bit_slice_2043893;
    p30_bit_slice_2044018 <= p29_bit_slice_2044018;
    p30_k3 <= p29_k3;
    p30_k2 <= p29_k2;
    p30_xor_2048752 <= p29_xor_2048752;
    p30_xor_2049240 <= p30_xor_2049240_comb;
    p30_array_index_2049256 <= p30_array_index_2049256_comb;
    p30_array_index_2049257 <= p30_array_index_2049257_comb;
    p30_array_index_2049258 <= p30_array_index_2049258_comb;
    p30_array_index_2049259 <= p30_array_index_2049259_comb;
    p30_array_index_2049260 <= p30_array_index_2049260_comb;
    p30_array_index_2049261 <= p30_array_index_2049261_comb;
    p30_array_index_2049263 <= p30_array_index_2049263_comb;
    p30_array_index_2049265 <= p30_array_index_2049265_comb;
    p30_array_index_2049266 <= p30_array_index_2049266_comb;
    p30_array_index_2049272 <= p30_array_index_2049272_comb;
    p30_array_index_2049273 <= p30_array_index_2049273_comb;
    p30_array_index_2049274 <= p30_array_index_2049274_comb;
    p30_array_index_2049275 <= p30_array_index_2049275_comb;
    p30_array_index_2049276 <= p30_array_index_2049276_comb;
    p30_array_index_2049278 <= p30_array_index_2049278_comb;
    p30_array_index_2049280 <= p30_array_index_2049280_comb;
    p30_res7__384 <= p30_res7__384_comb;
    p30_array_index_2049289 <= p30_array_index_2049289_comb;
    p30_array_index_2049290 <= p30_array_index_2049290_comb;
    p30_array_index_2049291 <= p30_array_index_2049291_comb;
    p30_array_index_2049292 <= p30_array_index_2049292_comb;
    p30_array_index_2049293 <= p30_array_index_2049293_comb;
    p30_array_index_2049294 <= p30_array_index_2049294_comb;
    p30_res7__386 <= p30_res7__386_comb;
    p30_array_index_2049304 <= p30_array_index_2049304_comb;
    p30_array_index_2049305 <= p30_array_index_2049305_comb;
    p30_array_index_2049306 <= p30_array_index_2049306_comb;
    p30_array_index_2049307 <= p30_array_index_2049307_comb;
    p30_array_index_2049308 <= p30_array_index_2049308_comb;
    p30_res7__388 <= p30_res7__388_comb;
    p30_array_index_2049318 <= p30_array_index_2049318_comb;
    p30_array_index_2049319 <= p30_array_index_2049319_comb;
    p30_array_index_2049320 <= p30_array_index_2049320_comb;
    p30_array_index_2049321 <= p30_array_index_2049321_comb;
    p30_array_index_2049322 <= p30_array_index_2049322_comb;
    p30_res7__390 <= p30_res7__390_comb;
    p30_array_index_2049333 <= p30_array_index_2049333_comb;
    p30_array_index_2049334 <= p30_array_index_2049334_comb;
    p30_array_index_2049335 <= p30_array_index_2049335_comb;
    p30_array_index_2049336 <= p30_array_index_2049336_comb;
    p30_res7__392 <= p30_res7__392_comb;
    p31_literal_2043896 <= p30_literal_2043896;
    p31_literal_2043910 <= p30_literal_2043910;
    p31_literal_2043912 <= p30_literal_2043912;
    p31_literal_2043914 <= p30_literal_2043914;
    p31_literal_2043916 <= p30_literal_2043916;
    p31_literal_2043918 <= p30_literal_2043918;
    p31_literal_2043920 <= p30_literal_2043920;
    p31_literal_2043923 <= p30_literal_2043923;
  end

  // ===== Pipe stage 31:
  wire [7:0] p31_array_index_2049458_comb;
  wire [7:0] p31_array_index_2049459_comb;
  wire [7:0] p31_array_index_2049460_comb;
  wire [7:0] p31_array_index_2049461_comb;
  wire [7:0] p31_res7__394_comb;
  wire [7:0] p31_array_index_2049472_comb;
  wire [7:0] p31_array_index_2049473_comb;
  wire [7:0] p31_array_index_2049474_comb;
  wire [7:0] p31_res7__396_comb;
  wire [7:0] p31_array_index_2049484_comb;
  wire [7:0] p31_array_index_2049485_comb;
  wire [7:0] p31_array_index_2049486_comb;
  wire [7:0] p31_res7__398_comb;
  wire [7:0] p31_array_index_2049497_comb;
  wire [7:0] p31_array_index_2049498_comb;
  wire [7:0] p31_res7__400_comb;
  wire [7:0] p31_array_index_2049508_comb;
  wire [7:0] p31_array_index_2049509_comb;
  wire [7:0] p31_res7__402_comb;
  wire [7:0] p31_array_index_2049520_comb;
  wire [7:0] p31_res7__404_comb;
  wire [7:0] p31_array_index_2049530_comb;
  wire [7:0] p31_res7__406_comb;
  assign p31_array_index_2049458_comb = p30_literal_2043914[p30_res7__388];
  assign p31_array_index_2049459_comb = p30_literal_2043916[p30_res7__386];
  assign p31_array_index_2049460_comb = p30_literal_2043918[p30_res7__384];
  assign p31_array_index_2049461_comb = p30_literal_2043920[p30_array_index_2049256];
  assign p31_res7__394_comb = p30_literal_2043910[p30_res7__392] ^ p30_literal_2043912[p30_res7__390] ^ p31_array_index_2049458_comb ^ p31_array_index_2049459_comb ^ p31_array_index_2049460_comb ^ p31_array_index_2049461_comb ^ p30_array_index_2049257 ^ p30_literal_2043923[p30_array_index_2049258] ^ p30_array_index_2049259 ^ p30_array_index_2049294 ^ p30_literal_2043918[p30_array_index_2049261] ^ p30_literal_2043916[p30_array_index_2049278] ^ p30_literal_2043914[p30_array_index_2049263] ^ p30_literal_2043912[p30_array_index_2049280] ^ p30_literal_2043910[p30_array_index_2049265] ^ p30_array_index_2049266;
  assign p31_array_index_2049472_comb = p30_literal_2043916[p30_res7__388];
  assign p31_array_index_2049473_comb = p30_literal_2043918[p30_res7__386];
  assign p31_array_index_2049474_comb = p30_literal_2043920[p30_res7__384];
  assign p31_res7__396_comb = p30_literal_2043910[p31_res7__394_comb] ^ p30_literal_2043912[p30_res7__392] ^ p30_literal_2043914[p30_res7__390] ^ p31_array_index_2049472_comb ^ p31_array_index_2049473_comb ^ p31_array_index_2049474_comb ^ p30_array_index_2049256 ^ p30_literal_2043923[p30_array_index_2049257] ^ p30_array_index_2049258 ^ p30_array_index_2049308 ^ p30_array_index_2049276 ^ p30_literal_2043916[p30_array_index_2049261] ^ p30_literal_2043914[p30_array_index_2049278] ^ p30_literal_2043912[p30_array_index_2049263] ^ p30_literal_2043910[p30_array_index_2049280] ^ p30_array_index_2049265;
  assign p31_array_index_2049484_comb = p30_literal_2043916[p30_res7__390];
  assign p31_array_index_2049485_comb = p30_literal_2043918[p30_res7__388];
  assign p31_array_index_2049486_comb = p30_literal_2043920[p30_res7__386];
  assign p31_res7__398_comb = p30_literal_2043910[p31_res7__396_comb] ^ p30_literal_2043912[p31_res7__394_comb] ^ p30_literal_2043914[p30_res7__392] ^ p31_array_index_2049484_comb ^ p31_array_index_2049485_comb ^ p31_array_index_2049486_comb ^ p30_res7__384 ^ p30_literal_2043923[p30_array_index_2049256] ^ p30_array_index_2049257 ^ p30_array_index_2049322 ^ p30_array_index_2049293 ^ p30_literal_2043916[p30_array_index_2049260] ^ p30_literal_2043914[p30_array_index_2049261] ^ p30_literal_2043912[p30_array_index_2049278] ^ p30_literal_2043910[p30_array_index_2049263] ^ p30_array_index_2049280;
  assign p31_array_index_2049497_comb = p30_literal_2043918[p30_res7__390];
  assign p31_array_index_2049498_comb = p30_literal_2043920[p30_res7__388];
  assign p31_res7__400_comb = p30_literal_2043910[p31_res7__398_comb] ^ p30_literal_2043912[p31_res7__396_comb] ^ p30_literal_2043914[p31_res7__394_comb] ^ p30_literal_2043916[p30_res7__392] ^ p31_array_index_2049497_comb ^ p31_array_index_2049498_comb ^ p30_res7__386 ^ p30_literal_2043923[p30_res7__384] ^ p30_array_index_2049256 ^ p30_array_index_2049336 ^ p30_array_index_2049307 ^ p30_array_index_2049275 ^ p30_literal_2043914[p30_array_index_2049260] ^ p30_literal_2043912[p30_array_index_2049261] ^ p30_literal_2043910[p30_array_index_2049278] ^ p30_array_index_2049263;
  assign p31_array_index_2049508_comb = p30_literal_2043918[p30_res7__392];
  assign p31_array_index_2049509_comb = p30_literal_2043920[p30_res7__390];
  assign p31_res7__402_comb = p30_literal_2043910[p31_res7__400_comb] ^ p30_literal_2043912[p31_res7__398_comb] ^ p30_literal_2043914[p31_res7__396_comb] ^ p30_literal_2043916[p31_res7__394_comb] ^ p31_array_index_2049508_comb ^ p31_array_index_2049509_comb ^ p30_res7__388 ^ p30_literal_2043923[p30_res7__386] ^ p30_res7__384 ^ p31_array_index_2049461_comb ^ p30_array_index_2049321 ^ p30_array_index_2049292 ^ p30_literal_2043914[p30_array_index_2049259] ^ p30_literal_2043912[p30_array_index_2049260] ^ p30_literal_2043910[p30_array_index_2049261] ^ p30_array_index_2049278;
  assign p31_array_index_2049520_comb = p30_literal_2043920[p30_res7__392];
  assign p31_res7__404_comb = p30_literal_2043910[p31_res7__402_comb] ^ p30_literal_2043912[p31_res7__400_comb] ^ p30_literal_2043914[p31_res7__398_comb] ^ p30_literal_2043916[p31_res7__396_comb] ^ p30_literal_2043918[p31_res7__394_comb] ^ p31_array_index_2049520_comb ^ p30_res7__390 ^ p30_literal_2043923[p30_res7__388] ^ p30_res7__386 ^ p31_array_index_2049474_comb ^ p30_array_index_2049335 ^ p30_array_index_2049306 ^ p30_array_index_2049274 ^ p30_literal_2043912[p30_array_index_2049259] ^ p30_literal_2043910[p30_array_index_2049260] ^ p30_array_index_2049261;
  assign p31_array_index_2049530_comb = p30_literal_2043920[p31_res7__394_comb];
  assign p31_res7__406_comb = p30_literal_2043910[p31_res7__404_comb] ^ p30_literal_2043912[p31_res7__402_comb] ^ p30_literal_2043914[p31_res7__400_comb] ^ p30_literal_2043916[p31_res7__398_comb] ^ p30_literal_2043918[p31_res7__396_comb] ^ p31_array_index_2049530_comb ^ p30_res7__392 ^ p30_literal_2043923[p30_res7__390] ^ p30_res7__388 ^ p31_array_index_2049486_comb ^ p31_array_index_2049460_comb ^ p30_array_index_2049320 ^ p30_array_index_2049291 ^ p30_literal_2043912[p30_array_index_2049258] ^ p30_literal_2043910[p30_array_index_2049259] ^ p30_array_index_2049260;

  // Registers for pipe stage 31:
  reg [127:0] p31_encoded;
  reg [127:0] p31_bit_slice_2043893;
  reg [127:0] p31_bit_slice_2044018;
  reg [127:0] p31_k3;
  reg [127:0] p31_k2;
  reg [127:0] p31_xor_2048752;
  reg [127:0] p31_xor_2049240;
  reg [7:0] p31_array_index_2049256;
  reg [7:0] p31_array_index_2049257;
  reg [7:0] p31_array_index_2049258;
  reg [7:0] p31_array_index_2049259;
  reg [7:0] p31_array_index_2049272;
  reg [7:0] p31_array_index_2049273;
  reg [7:0] p31_res7__384;
  reg [7:0] p31_array_index_2049289;
  reg [7:0] p31_array_index_2049290;
  reg [7:0] p31_res7__386;
  reg [7:0] p31_array_index_2049304;
  reg [7:0] p31_array_index_2049305;
  reg [7:0] p31_res7__388;
  reg [7:0] p31_array_index_2049318;
  reg [7:0] p31_array_index_2049319;
  reg [7:0] p31_res7__390;
  reg [7:0] p31_array_index_2049333;
  reg [7:0] p31_array_index_2049334;
  reg [7:0] p31_res7__392;
  reg [7:0] p31_array_index_2049458;
  reg [7:0] p31_array_index_2049459;
  reg [7:0] p31_res7__394;
  reg [7:0] p31_array_index_2049472;
  reg [7:0] p31_array_index_2049473;
  reg [7:0] p31_res7__396;
  reg [7:0] p31_array_index_2049484;
  reg [7:0] p31_array_index_2049485;
  reg [7:0] p31_res7__398;
  reg [7:0] p31_array_index_2049497;
  reg [7:0] p31_array_index_2049498;
  reg [7:0] p31_res7__400;
  reg [7:0] p31_array_index_2049508;
  reg [7:0] p31_array_index_2049509;
  reg [7:0] p31_res7__402;
  reg [7:0] p31_array_index_2049520;
  reg [7:0] p31_res7__404;
  reg [7:0] p31_array_index_2049530;
  reg [7:0] p31_res7__406;
  reg [7:0] p32_literal_2043896[256];
  reg [7:0] p32_literal_2043910[256];
  reg [7:0] p32_literal_2043912[256];
  reg [7:0] p32_literal_2043914[256];
  reg [7:0] p32_literal_2043916[256];
  reg [7:0] p32_literal_2043918[256];
  reg [7:0] p32_literal_2043920[256];
  reg [7:0] p32_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p31_encoded <= p30_encoded;
    p31_bit_slice_2043893 <= p30_bit_slice_2043893;
    p31_bit_slice_2044018 <= p30_bit_slice_2044018;
    p31_k3 <= p30_k3;
    p31_k2 <= p30_k2;
    p31_xor_2048752 <= p30_xor_2048752;
    p31_xor_2049240 <= p30_xor_2049240;
    p31_array_index_2049256 <= p30_array_index_2049256;
    p31_array_index_2049257 <= p30_array_index_2049257;
    p31_array_index_2049258 <= p30_array_index_2049258;
    p31_array_index_2049259 <= p30_array_index_2049259;
    p31_array_index_2049272 <= p30_array_index_2049272;
    p31_array_index_2049273 <= p30_array_index_2049273;
    p31_res7__384 <= p30_res7__384;
    p31_array_index_2049289 <= p30_array_index_2049289;
    p31_array_index_2049290 <= p30_array_index_2049290;
    p31_res7__386 <= p30_res7__386;
    p31_array_index_2049304 <= p30_array_index_2049304;
    p31_array_index_2049305 <= p30_array_index_2049305;
    p31_res7__388 <= p30_res7__388;
    p31_array_index_2049318 <= p30_array_index_2049318;
    p31_array_index_2049319 <= p30_array_index_2049319;
    p31_res7__390 <= p30_res7__390;
    p31_array_index_2049333 <= p30_array_index_2049333;
    p31_array_index_2049334 <= p30_array_index_2049334;
    p31_res7__392 <= p30_res7__392;
    p31_array_index_2049458 <= p31_array_index_2049458_comb;
    p31_array_index_2049459 <= p31_array_index_2049459_comb;
    p31_res7__394 <= p31_res7__394_comb;
    p31_array_index_2049472 <= p31_array_index_2049472_comb;
    p31_array_index_2049473 <= p31_array_index_2049473_comb;
    p31_res7__396 <= p31_res7__396_comb;
    p31_array_index_2049484 <= p31_array_index_2049484_comb;
    p31_array_index_2049485 <= p31_array_index_2049485_comb;
    p31_res7__398 <= p31_res7__398_comb;
    p31_array_index_2049497 <= p31_array_index_2049497_comb;
    p31_array_index_2049498 <= p31_array_index_2049498_comb;
    p31_res7__400 <= p31_res7__400_comb;
    p31_array_index_2049508 <= p31_array_index_2049508_comb;
    p31_array_index_2049509 <= p31_array_index_2049509_comb;
    p31_res7__402 <= p31_res7__402_comb;
    p31_array_index_2049520 <= p31_array_index_2049520_comb;
    p31_res7__404 <= p31_res7__404_comb;
    p31_array_index_2049530 <= p31_array_index_2049530_comb;
    p31_res7__406 <= p31_res7__406_comb;
    p32_literal_2043896 <= p31_literal_2043896;
    p32_literal_2043910 <= p31_literal_2043910;
    p32_literal_2043912 <= p31_literal_2043912;
    p32_literal_2043914 <= p31_literal_2043914;
    p32_literal_2043916 <= p31_literal_2043916;
    p32_literal_2043918 <= p31_literal_2043918;
    p32_literal_2043920 <= p31_literal_2043920;
    p32_literal_2043923 <= p31_literal_2043923;
  end

  // ===== Pipe stage 32:
  wire [7:0] p32_res7__408_comb;
  wire [7:0] p32_res7__410_comb;
  wire [7:0] p32_res7__412_comb;
  wire [7:0] p32_res7__414_comb;
  wire [127:0] p32_res__12_comb;
  wire [127:0] p32_xor_2049676_comb;
  wire [127:0] p32_addedKey__45_comb;
  wire [7:0] p32_array_index_2049692_comb;
  wire [7:0] p32_array_index_2049693_comb;
  wire [7:0] p32_array_index_2049694_comb;
  wire [7:0] p32_array_index_2049695_comb;
  wire [7:0] p32_array_index_2049696_comb;
  wire [7:0] p32_array_index_2049697_comb;
  wire [7:0] p32_array_index_2049699_comb;
  wire [7:0] p32_array_index_2049701_comb;
  wire [7:0] p32_array_index_2049702_comb;
  wire [7:0] p32_array_index_2049703_comb;
  wire [7:0] p32_array_index_2049704_comb;
  wire [7:0] p32_array_index_2049705_comb;
  wire [7:0] p32_array_index_2049706_comb;
  wire [7:0] p32_array_index_2049708_comb;
  wire [7:0] p32_array_index_2049709_comb;
  wire [7:0] p32_array_index_2049710_comb;
  wire [7:0] p32_array_index_2049711_comb;
  wire [7:0] p32_array_index_2049712_comb;
  wire [7:0] p32_array_index_2049713_comb;
  wire [7:0] p32_array_index_2049714_comb;
  wire [7:0] p32_array_index_2049716_comb;
  wire [7:0] p32_res7__416_comb;
  wire [7:0] p32_array_index_2049725_comb;
  wire [7:0] p32_array_index_2049726_comb;
  wire [7:0] p32_array_index_2049727_comb;
  wire [7:0] p32_array_index_2049728_comb;
  wire [7:0] p32_array_index_2049729_comb;
  wire [7:0] p32_array_index_2049730_comb;
  wire [7:0] p32_res7__418_comb;
  assign p32_res7__408_comb = p31_literal_2043910[p31_res7__406] ^ p31_literal_2043912[p31_res7__404] ^ p31_literal_2043914[p31_res7__402] ^ p31_literal_2043916[p31_res7__400] ^ p31_literal_2043918[p31_res7__398] ^ p31_literal_2043920[p31_res7__396] ^ p31_res7__394 ^ p31_literal_2043923[p31_res7__392] ^ p31_res7__390 ^ p31_array_index_2049498 ^ p31_array_index_2049473 ^ p31_array_index_2049334 ^ p31_array_index_2049305 ^ p31_array_index_2049273 ^ p31_literal_2043910[p31_array_index_2049258] ^ p31_array_index_2049259;
  assign p32_res7__410_comb = p31_literal_2043910[p32_res7__408_comb] ^ p31_literal_2043912[p31_res7__406] ^ p31_literal_2043914[p31_res7__404] ^ p31_literal_2043916[p31_res7__402] ^ p31_literal_2043918[p31_res7__400] ^ p31_literal_2043920[p31_res7__398] ^ p31_res7__396 ^ p31_literal_2043923[p31_res7__394] ^ p31_res7__392 ^ p31_array_index_2049509 ^ p31_array_index_2049485 ^ p31_array_index_2049459 ^ p31_array_index_2049319 ^ p31_array_index_2049290 ^ p31_literal_2043910[p31_array_index_2049257] ^ p31_array_index_2049258;
  assign p32_res7__412_comb = p31_literal_2043910[p32_res7__410_comb] ^ p31_literal_2043912[p32_res7__408_comb] ^ p31_literal_2043914[p31_res7__406] ^ p31_literal_2043916[p31_res7__404] ^ p31_literal_2043918[p31_res7__402] ^ p31_literal_2043920[p31_res7__400] ^ p31_res7__398 ^ p31_literal_2043923[p31_res7__396] ^ p31_res7__394 ^ p31_array_index_2049520 ^ p31_array_index_2049497 ^ p31_array_index_2049472 ^ p31_array_index_2049333 ^ p31_array_index_2049304 ^ p31_array_index_2049272 ^ p31_array_index_2049257;
  assign p32_res7__414_comb = p31_literal_2043910[p32_res7__412_comb] ^ p31_literal_2043912[p32_res7__410_comb] ^ p31_literal_2043914[p32_res7__408_comb] ^ p31_literal_2043916[p31_res7__406] ^ p31_literal_2043918[p31_res7__404] ^ p31_literal_2043920[p31_res7__402] ^ p31_res7__400 ^ p31_literal_2043923[p31_res7__398] ^ p31_res7__396 ^ p31_array_index_2049530 ^ p31_array_index_2049508 ^ p31_array_index_2049484 ^ p31_array_index_2049458 ^ p31_array_index_2049318 ^ p31_array_index_2049289 ^ p31_array_index_2049256;
  assign p32_res__12_comb = {p32_res7__414_comb, p32_res7__412_comb, p32_res7__410_comb, p32_res7__408_comb, p31_res7__406, p31_res7__404, p31_res7__402, p31_res7__400, p31_res7__398, p31_res7__396, p31_res7__394, p31_res7__392, p31_res7__390, p31_res7__388, p31_res7__386, p31_res7__384};
  assign p32_xor_2049676_comb = p32_res__12_comb ^ p31_xor_2048752;
  assign p32_addedKey__45_comb = p32_xor_2049676_comb ^ 128'h5113_c1f9_4d76_899f_a029_a9e0_ac34_d40e;
  assign p32_array_index_2049692_comb = p31_literal_2043896[p32_addedKey__45_comb[127:120]];
  assign p32_array_index_2049693_comb = p31_literal_2043896[p32_addedKey__45_comb[119:112]];
  assign p32_array_index_2049694_comb = p31_literal_2043896[p32_addedKey__45_comb[111:104]];
  assign p32_array_index_2049695_comb = p31_literal_2043896[p32_addedKey__45_comb[103:96]];
  assign p32_array_index_2049696_comb = p31_literal_2043896[p32_addedKey__45_comb[95:88]];
  assign p32_array_index_2049697_comb = p31_literal_2043896[p32_addedKey__45_comb[87:80]];
  assign p32_array_index_2049699_comb = p31_literal_2043896[p32_addedKey__45_comb[71:64]];
  assign p32_array_index_2049701_comb = p31_literal_2043896[p32_addedKey__45_comb[55:48]];
  assign p32_array_index_2049702_comb = p31_literal_2043896[p32_addedKey__45_comb[47:40]];
  assign p32_array_index_2049703_comb = p31_literal_2043896[p32_addedKey__45_comb[39:32]];
  assign p32_array_index_2049704_comb = p31_literal_2043896[p32_addedKey__45_comb[31:24]];
  assign p32_array_index_2049705_comb = p31_literal_2043896[p32_addedKey__45_comb[23:16]];
  assign p32_array_index_2049706_comb = p31_literal_2043896[p32_addedKey__45_comb[15:8]];
  assign p32_array_index_2049708_comb = p31_literal_2043910[p32_array_index_2049692_comb];
  assign p32_array_index_2049709_comb = p31_literal_2043912[p32_array_index_2049693_comb];
  assign p32_array_index_2049710_comb = p31_literal_2043914[p32_array_index_2049694_comb];
  assign p32_array_index_2049711_comb = p31_literal_2043916[p32_array_index_2049695_comb];
  assign p32_array_index_2049712_comb = p31_literal_2043918[p32_array_index_2049696_comb];
  assign p32_array_index_2049713_comb = p31_literal_2043920[p32_array_index_2049697_comb];
  assign p32_array_index_2049714_comb = p31_literal_2043896[p32_addedKey__45_comb[79:72]];
  assign p32_array_index_2049716_comb = p31_literal_2043896[p32_addedKey__45_comb[63:56]];
  assign p32_res7__416_comb = p32_array_index_2049708_comb ^ p32_array_index_2049709_comb ^ p32_array_index_2049710_comb ^ p32_array_index_2049711_comb ^ p32_array_index_2049712_comb ^ p32_array_index_2049713_comb ^ p32_array_index_2049714_comb ^ p31_literal_2043923[p32_array_index_2049699_comb] ^ p32_array_index_2049716_comb ^ p31_literal_2043920[p32_array_index_2049701_comb] ^ p31_literal_2043918[p32_array_index_2049702_comb] ^ p31_literal_2043916[p32_array_index_2049703_comb] ^ p31_literal_2043914[p32_array_index_2049704_comb] ^ p31_literal_2043912[p32_array_index_2049705_comb] ^ p31_literal_2043910[p32_array_index_2049706_comb] ^ p31_literal_2043896[p32_addedKey__45_comb[7:0]];
  assign p32_array_index_2049725_comb = p31_literal_2043910[p32_res7__416_comb];
  assign p32_array_index_2049726_comb = p31_literal_2043912[p32_array_index_2049692_comb];
  assign p32_array_index_2049727_comb = p31_literal_2043914[p32_array_index_2049693_comb];
  assign p32_array_index_2049728_comb = p31_literal_2043916[p32_array_index_2049694_comb];
  assign p32_array_index_2049729_comb = p31_literal_2043918[p32_array_index_2049695_comb];
  assign p32_array_index_2049730_comb = p31_literal_2043920[p32_array_index_2049696_comb];
  assign p32_res7__418_comb = p32_array_index_2049725_comb ^ p32_array_index_2049726_comb ^ p32_array_index_2049727_comb ^ p32_array_index_2049728_comb ^ p32_array_index_2049729_comb ^ p32_array_index_2049730_comb ^ p32_array_index_2049697_comb ^ p31_literal_2043923[p32_array_index_2049714_comb] ^ p32_array_index_2049699_comb ^ p31_literal_2043920[p32_array_index_2049716_comb] ^ p31_literal_2043918[p32_array_index_2049701_comb] ^ p31_literal_2043916[p32_array_index_2049702_comb] ^ p31_literal_2043914[p32_array_index_2049703_comb] ^ p31_literal_2043912[p32_array_index_2049704_comb] ^ p31_literal_2043910[p32_array_index_2049705_comb] ^ p32_array_index_2049706_comb;

  // Registers for pipe stage 32:
  reg [127:0] p32_encoded;
  reg [127:0] p32_bit_slice_2043893;
  reg [127:0] p32_bit_slice_2044018;
  reg [127:0] p32_k3;
  reg [127:0] p32_k2;
  reg [127:0] p32_xor_2049240;
  reg [127:0] p32_xor_2049676;
  reg [7:0] p32_array_index_2049692;
  reg [7:0] p32_array_index_2049693;
  reg [7:0] p32_array_index_2049694;
  reg [7:0] p32_array_index_2049695;
  reg [7:0] p32_array_index_2049696;
  reg [7:0] p32_array_index_2049697;
  reg [7:0] p32_array_index_2049699;
  reg [7:0] p32_array_index_2049701;
  reg [7:0] p32_array_index_2049702;
  reg [7:0] p32_array_index_2049703;
  reg [7:0] p32_array_index_2049704;
  reg [7:0] p32_array_index_2049705;
  reg [7:0] p32_array_index_2049708;
  reg [7:0] p32_array_index_2049709;
  reg [7:0] p32_array_index_2049710;
  reg [7:0] p32_array_index_2049711;
  reg [7:0] p32_array_index_2049712;
  reg [7:0] p32_array_index_2049713;
  reg [7:0] p32_array_index_2049714;
  reg [7:0] p32_array_index_2049716;
  reg [7:0] p32_res7__416;
  reg [7:0] p32_array_index_2049725;
  reg [7:0] p32_array_index_2049726;
  reg [7:0] p32_array_index_2049727;
  reg [7:0] p32_array_index_2049728;
  reg [7:0] p32_array_index_2049729;
  reg [7:0] p32_array_index_2049730;
  reg [7:0] p32_res7__418;
  reg [7:0] p33_literal_2043896[256];
  reg [7:0] p33_literal_2043910[256];
  reg [7:0] p33_literal_2043912[256];
  reg [7:0] p33_literal_2043914[256];
  reg [7:0] p33_literal_2043916[256];
  reg [7:0] p33_literal_2043918[256];
  reg [7:0] p33_literal_2043920[256];
  reg [7:0] p33_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p32_encoded <= p31_encoded;
    p32_bit_slice_2043893 <= p31_bit_slice_2043893;
    p32_bit_slice_2044018 <= p31_bit_slice_2044018;
    p32_k3 <= p31_k3;
    p32_k2 <= p31_k2;
    p32_xor_2049240 <= p31_xor_2049240;
    p32_xor_2049676 <= p32_xor_2049676_comb;
    p32_array_index_2049692 <= p32_array_index_2049692_comb;
    p32_array_index_2049693 <= p32_array_index_2049693_comb;
    p32_array_index_2049694 <= p32_array_index_2049694_comb;
    p32_array_index_2049695 <= p32_array_index_2049695_comb;
    p32_array_index_2049696 <= p32_array_index_2049696_comb;
    p32_array_index_2049697 <= p32_array_index_2049697_comb;
    p32_array_index_2049699 <= p32_array_index_2049699_comb;
    p32_array_index_2049701 <= p32_array_index_2049701_comb;
    p32_array_index_2049702 <= p32_array_index_2049702_comb;
    p32_array_index_2049703 <= p32_array_index_2049703_comb;
    p32_array_index_2049704 <= p32_array_index_2049704_comb;
    p32_array_index_2049705 <= p32_array_index_2049705_comb;
    p32_array_index_2049708 <= p32_array_index_2049708_comb;
    p32_array_index_2049709 <= p32_array_index_2049709_comb;
    p32_array_index_2049710 <= p32_array_index_2049710_comb;
    p32_array_index_2049711 <= p32_array_index_2049711_comb;
    p32_array_index_2049712 <= p32_array_index_2049712_comb;
    p32_array_index_2049713 <= p32_array_index_2049713_comb;
    p32_array_index_2049714 <= p32_array_index_2049714_comb;
    p32_array_index_2049716 <= p32_array_index_2049716_comb;
    p32_res7__416 <= p32_res7__416_comb;
    p32_array_index_2049725 <= p32_array_index_2049725_comb;
    p32_array_index_2049726 <= p32_array_index_2049726_comb;
    p32_array_index_2049727 <= p32_array_index_2049727_comb;
    p32_array_index_2049728 <= p32_array_index_2049728_comb;
    p32_array_index_2049729 <= p32_array_index_2049729_comb;
    p32_array_index_2049730 <= p32_array_index_2049730_comb;
    p32_res7__418 <= p32_res7__418_comb;
    p33_literal_2043896 <= p32_literal_2043896;
    p33_literal_2043910 <= p32_literal_2043910;
    p33_literal_2043912 <= p32_literal_2043912;
    p33_literal_2043914 <= p32_literal_2043914;
    p33_literal_2043916 <= p32_literal_2043916;
    p33_literal_2043918 <= p32_literal_2043918;
    p33_literal_2043920 <= p32_literal_2043920;
    p33_literal_2043923 <= p32_literal_2043923;
  end

  // ===== Pipe stage 33:
  wire [7:0] p33_array_index_2049826_comb;
  wire [7:0] p33_array_index_2049827_comb;
  wire [7:0] p33_array_index_2049828_comb;
  wire [7:0] p33_array_index_2049829_comb;
  wire [7:0] p33_array_index_2049830_comb;
  wire [7:0] p33_res7__420_comb;
  wire [7:0] p33_array_index_2049840_comb;
  wire [7:0] p33_array_index_2049841_comb;
  wire [7:0] p33_array_index_2049842_comb;
  wire [7:0] p33_array_index_2049843_comb;
  wire [7:0] p33_array_index_2049844_comb;
  wire [7:0] p33_res7__422_comb;
  wire [7:0] p33_array_index_2049855_comb;
  wire [7:0] p33_array_index_2049856_comb;
  wire [7:0] p33_array_index_2049857_comb;
  wire [7:0] p33_array_index_2049858_comb;
  wire [7:0] p33_res7__424_comb;
  wire [7:0] p33_array_index_2049868_comb;
  wire [7:0] p33_array_index_2049869_comb;
  wire [7:0] p33_array_index_2049870_comb;
  wire [7:0] p33_array_index_2049871_comb;
  wire [7:0] p33_res7__426_comb;
  wire [7:0] p33_array_index_2049882_comb;
  wire [7:0] p33_array_index_2049883_comb;
  wire [7:0] p33_array_index_2049884_comb;
  wire [7:0] p33_res7__428_comb;
  wire [7:0] p33_array_index_2049894_comb;
  wire [7:0] p33_array_index_2049895_comb;
  wire [7:0] p33_array_index_2049896_comb;
  wire [7:0] p33_res7__430_comb;
  wire [7:0] p33_array_index_2049907_comb;
  wire [7:0] p33_array_index_2049908_comb;
  wire [7:0] p33_res7__432_comb;
  assign p33_array_index_2049826_comb = p32_literal_2043912[p32_res7__416];
  assign p33_array_index_2049827_comb = p32_literal_2043914[p32_array_index_2049692];
  assign p33_array_index_2049828_comb = p32_literal_2043916[p32_array_index_2049693];
  assign p33_array_index_2049829_comb = p32_literal_2043918[p32_array_index_2049694];
  assign p33_array_index_2049830_comb = p32_literal_2043920[p32_array_index_2049695];
  assign p33_res7__420_comb = p32_literal_2043910[p32_res7__418] ^ p33_array_index_2049826_comb ^ p33_array_index_2049827_comb ^ p33_array_index_2049828_comb ^ p33_array_index_2049829_comb ^ p33_array_index_2049830_comb ^ p32_array_index_2049696 ^ p32_literal_2043923[p32_array_index_2049697] ^ p32_array_index_2049714 ^ p32_literal_2043920[p32_array_index_2049699] ^ p32_literal_2043918[p32_array_index_2049716] ^ p32_literal_2043916[p32_array_index_2049701] ^ p32_literal_2043914[p32_array_index_2049702] ^ p32_literal_2043912[p32_array_index_2049703] ^ p32_literal_2043910[p32_array_index_2049704] ^ p32_array_index_2049705;
  assign p33_array_index_2049840_comb = p32_literal_2043912[p32_res7__418];
  assign p33_array_index_2049841_comb = p32_literal_2043914[p32_res7__416];
  assign p33_array_index_2049842_comb = p32_literal_2043916[p32_array_index_2049692];
  assign p33_array_index_2049843_comb = p32_literal_2043918[p32_array_index_2049693];
  assign p33_array_index_2049844_comb = p32_literal_2043920[p32_array_index_2049694];
  assign p33_res7__422_comb = p32_literal_2043910[p33_res7__420_comb] ^ p33_array_index_2049840_comb ^ p33_array_index_2049841_comb ^ p33_array_index_2049842_comb ^ p33_array_index_2049843_comb ^ p33_array_index_2049844_comb ^ p32_array_index_2049695 ^ p32_literal_2043923[p32_array_index_2049696] ^ p32_array_index_2049697 ^ p32_literal_2043920[p32_array_index_2049714] ^ p32_literal_2043918[p32_array_index_2049699] ^ p32_literal_2043916[p32_array_index_2049716] ^ p32_literal_2043914[p32_array_index_2049701] ^ p32_literal_2043912[p32_array_index_2049702] ^ p32_literal_2043910[p32_array_index_2049703] ^ p32_array_index_2049704;
  assign p33_array_index_2049855_comb = p32_literal_2043914[p32_res7__418];
  assign p33_array_index_2049856_comb = p32_literal_2043916[p32_res7__416];
  assign p33_array_index_2049857_comb = p32_literal_2043918[p32_array_index_2049692];
  assign p33_array_index_2049858_comb = p32_literal_2043920[p32_array_index_2049693];
  assign p33_res7__424_comb = p32_literal_2043910[p33_res7__422_comb] ^ p32_literal_2043912[p33_res7__420_comb] ^ p33_array_index_2049855_comb ^ p33_array_index_2049856_comb ^ p33_array_index_2049857_comb ^ p33_array_index_2049858_comb ^ p32_array_index_2049694 ^ p32_literal_2043923[p32_array_index_2049695] ^ p32_array_index_2049696 ^ p32_array_index_2049713 ^ p32_literal_2043918[p32_array_index_2049714] ^ p32_literal_2043916[p32_array_index_2049699] ^ p32_literal_2043914[p32_array_index_2049716] ^ p32_literal_2043912[p32_array_index_2049701] ^ p32_literal_2043910[p32_array_index_2049702] ^ p32_array_index_2049703;
  assign p33_array_index_2049868_comb = p32_literal_2043914[p33_res7__420_comb];
  assign p33_array_index_2049869_comb = p32_literal_2043916[p32_res7__418];
  assign p33_array_index_2049870_comb = p32_literal_2043918[p32_res7__416];
  assign p33_array_index_2049871_comb = p32_literal_2043920[p32_array_index_2049692];
  assign p33_res7__426_comb = p32_literal_2043910[p33_res7__424_comb] ^ p32_literal_2043912[p33_res7__422_comb] ^ p33_array_index_2049868_comb ^ p33_array_index_2049869_comb ^ p33_array_index_2049870_comb ^ p33_array_index_2049871_comb ^ p32_array_index_2049693 ^ p32_literal_2043923[p32_array_index_2049694] ^ p32_array_index_2049695 ^ p32_array_index_2049730 ^ p32_literal_2043918[p32_array_index_2049697] ^ p32_literal_2043916[p32_array_index_2049714] ^ p32_literal_2043914[p32_array_index_2049699] ^ p32_literal_2043912[p32_array_index_2049716] ^ p32_literal_2043910[p32_array_index_2049701] ^ p32_array_index_2049702;
  assign p33_array_index_2049882_comb = p32_literal_2043916[p33_res7__420_comb];
  assign p33_array_index_2049883_comb = p32_literal_2043918[p32_res7__418];
  assign p33_array_index_2049884_comb = p32_literal_2043920[p32_res7__416];
  assign p33_res7__428_comb = p32_literal_2043910[p33_res7__426_comb] ^ p32_literal_2043912[p33_res7__424_comb] ^ p32_literal_2043914[p33_res7__422_comb] ^ p33_array_index_2049882_comb ^ p33_array_index_2049883_comb ^ p33_array_index_2049884_comb ^ p32_array_index_2049692 ^ p32_literal_2043923[p32_array_index_2049693] ^ p32_array_index_2049694 ^ p33_array_index_2049830_comb ^ p32_array_index_2049712 ^ p32_literal_2043916[p32_array_index_2049697] ^ p32_literal_2043914[p32_array_index_2049714] ^ p32_literal_2043912[p32_array_index_2049699] ^ p32_literal_2043910[p32_array_index_2049716] ^ p32_array_index_2049701;
  assign p33_array_index_2049894_comb = p32_literal_2043916[p33_res7__422_comb];
  assign p33_array_index_2049895_comb = p32_literal_2043918[p33_res7__420_comb];
  assign p33_array_index_2049896_comb = p32_literal_2043920[p32_res7__418];
  assign p33_res7__430_comb = p32_literal_2043910[p33_res7__428_comb] ^ p32_literal_2043912[p33_res7__426_comb] ^ p32_literal_2043914[p33_res7__424_comb] ^ p33_array_index_2049894_comb ^ p33_array_index_2049895_comb ^ p33_array_index_2049896_comb ^ p32_res7__416 ^ p32_literal_2043923[p32_array_index_2049692] ^ p32_array_index_2049693 ^ p33_array_index_2049844_comb ^ p32_array_index_2049729 ^ p32_literal_2043916[p32_array_index_2049696] ^ p32_literal_2043914[p32_array_index_2049697] ^ p32_literal_2043912[p32_array_index_2049714] ^ p32_literal_2043910[p32_array_index_2049699] ^ p32_array_index_2049716;
  assign p33_array_index_2049907_comb = p32_literal_2043918[p33_res7__422_comb];
  assign p33_array_index_2049908_comb = p32_literal_2043920[p33_res7__420_comb];
  assign p33_res7__432_comb = p32_literal_2043910[p33_res7__430_comb] ^ p32_literal_2043912[p33_res7__428_comb] ^ p32_literal_2043914[p33_res7__426_comb] ^ p32_literal_2043916[p33_res7__424_comb] ^ p33_array_index_2049907_comb ^ p33_array_index_2049908_comb ^ p32_res7__418 ^ p32_literal_2043923[p32_res7__416] ^ p32_array_index_2049692 ^ p33_array_index_2049858_comb ^ p33_array_index_2049829_comb ^ p32_array_index_2049711 ^ p32_literal_2043914[p32_array_index_2049696] ^ p32_literal_2043912[p32_array_index_2049697] ^ p32_literal_2043910[p32_array_index_2049714] ^ p32_array_index_2049699;

  // Registers for pipe stage 33:
  reg [127:0] p33_encoded;
  reg [127:0] p33_bit_slice_2043893;
  reg [127:0] p33_bit_slice_2044018;
  reg [127:0] p33_k3;
  reg [127:0] p33_k2;
  reg [127:0] p33_xor_2049240;
  reg [127:0] p33_xor_2049676;
  reg [7:0] p33_array_index_2049692;
  reg [7:0] p33_array_index_2049693;
  reg [7:0] p33_array_index_2049694;
  reg [7:0] p33_array_index_2049695;
  reg [7:0] p33_array_index_2049696;
  reg [7:0] p33_array_index_2049697;
  reg [7:0] p33_array_index_2049708;
  reg [7:0] p33_array_index_2049709;
  reg [7:0] p33_array_index_2049710;
  reg [7:0] p33_array_index_2049714;
  reg [7:0] p33_res7__416;
  reg [7:0] p33_array_index_2049725;
  reg [7:0] p33_array_index_2049726;
  reg [7:0] p33_array_index_2049727;
  reg [7:0] p33_array_index_2049728;
  reg [7:0] p33_res7__418;
  reg [7:0] p33_array_index_2049826;
  reg [7:0] p33_array_index_2049827;
  reg [7:0] p33_array_index_2049828;
  reg [7:0] p33_res7__420;
  reg [7:0] p33_array_index_2049840;
  reg [7:0] p33_array_index_2049841;
  reg [7:0] p33_array_index_2049842;
  reg [7:0] p33_array_index_2049843;
  reg [7:0] p33_res7__422;
  reg [7:0] p33_array_index_2049855;
  reg [7:0] p33_array_index_2049856;
  reg [7:0] p33_array_index_2049857;
  reg [7:0] p33_res7__424;
  reg [7:0] p33_array_index_2049868;
  reg [7:0] p33_array_index_2049869;
  reg [7:0] p33_array_index_2049870;
  reg [7:0] p33_array_index_2049871;
  reg [7:0] p33_res7__426;
  reg [7:0] p33_array_index_2049882;
  reg [7:0] p33_array_index_2049883;
  reg [7:0] p33_array_index_2049884;
  reg [7:0] p33_res7__428;
  reg [7:0] p33_array_index_2049894;
  reg [7:0] p33_array_index_2049895;
  reg [7:0] p33_array_index_2049896;
  reg [7:0] p33_res7__430;
  reg [7:0] p33_array_index_2049907;
  reg [7:0] p33_array_index_2049908;
  reg [7:0] p33_res7__432;
  reg [7:0] p34_literal_2043896[256];
  reg [7:0] p34_literal_2043910[256];
  reg [7:0] p34_literal_2043912[256];
  reg [7:0] p34_literal_2043914[256];
  reg [7:0] p34_literal_2043916[256];
  reg [7:0] p34_literal_2043918[256];
  reg [7:0] p34_literal_2043920[256];
  reg [7:0] p34_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p33_encoded <= p32_encoded;
    p33_bit_slice_2043893 <= p32_bit_slice_2043893;
    p33_bit_slice_2044018 <= p32_bit_slice_2044018;
    p33_k3 <= p32_k3;
    p33_k2 <= p32_k2;
    p33_xor_2049240 <= p32_xor_2049240;
    p33_xor_2049676 <= p32_xor_2049676;
    p33_array_index_2049692 <= p32_array_index_2049692;
    p33_array_index_2049693 <= p32_array_index_2049693;
    p33_array_index_2049694 <= p32_array_index_2049694;
    p33_array_index_2049695 <= p32_array_index_2049695;
    p33_array_index_2049696 <= p32_array_index_2049696;
    p33_array_index_2049697 <= p32_array_index_2049697;
    p33_array_index_2049708 <= p32_array_index_2049708;
    p33_array_index_2049709 <= p32_array_index_2049709;
    p33_array_index_2049710 <= p32_array_index_2049710;
    p33_array_index_2049714 <= p32_array_index_2049714;
    p33_res7__416 <= p32_res7__416;
    p33_array_index_2049725 <= p32_array_index_2049725;
    p33_array_index_2049726 <= p32_array_index_2049726;
    p33_array_index_2049727 <= p32_array_index_2049727;
    p33_array_index_2049728 <= p32_array_index_2049728;
    p33_res7__418 <= p32_res7__418;
    p33_array_index_2049826 <= p33_array_index_2049826_comb;
    p33_array_index_2049827 <= p33_array_index_2049827_comb;
    p33_array_index_2049828 <= p33_array_index_2049828_comb;
    p33_res7__420 <= p33_res7__420_comb;
    p33_array_index_2049840 <= p33_array_index_2049840_comb;
    p33_array_index_2049841 <= p33_array_index_2049841_comb;
    p33_array_index_2049842 <= p33_array_index_2049842_comb;
    p33_array_index_2049843 <= p33_array_index_2049843_comb;
    p33_res7__422 <= p33_res7__422_comb;
    p33_array_index_2049855 <= p33_array_index_2049855_comb;
    p33_array_index_2049856 <= p33_array_index_2049856_comb;
    p33_array_index_2049857 <= p33_array_index_2049857_comb;
    p33_res7__424 <= p33_res7__424_comb;
    p33_array_index_2049868 <= p33_array_index_2049868_comb;
    p33_array_index_2049869 <= p33_array_index_2049869_comb;
    p33_array_index_2049870 <= p33_array_index_2049870_comb;
    p33_array_index_2049871 <= p33_array_index_2049871_comb;
    p33_res7__426 <= p33_res7__426_comb;
    p33_array_index_2049882 <= p33_array_index_2049882_comb;
    p33_array_index_2049883 <= p33_array_index_2049883_comb;
    p33_array_index_2049884 <= p33_array_index_2049884_comb;
    p33_res7__428 <= p33_res7__428_comb;
    p33_array_index_2049894 <= p33_array_index_2049894_comb;
    p33_array_index_2049895 <= p33_array_index_2049895_comb;
    p33_array_index_2049896 <= p33_array_index_2049896_comb;
    p33_res7__430 <= p33_res7__430_comb;
    p33_array_index_2049907 <= p33_array_index_2049907_comb;
    p33_array_index_2049908 <= p33_array_index_2049908_comb;
    p33_res7__432 <= p33_res7__432_comb;
    p34_literal_2043896 <= p33_literal_2043896;
    p34_literal_2043910 <= p33_literal_2043910;
    p34_literal_2043912 <= p33_literal_2043912;
    p34_literal_2043914 <= p33_literal_2043914;
    p34_literal_2043916 <= p33_literal_2043916;
    p34_literal_2043918 <= p33_literal_2043918;
    p34_literal_2043920 <= p33_literal_2043920;
    p34_literal_2043923 <= p33_literal_2043923;
  end

  // ===== Pipe stage 34:
  wire [7:0] p34_array_index_2050038_comb;
  wire [7:0] p34_array_index_2050039_comb;
  wire [7:0] p34_res7__434_comb;
  wire [7:0] p34_array_index_2050050_comb;
  wire [7:0] p34_res7__436_comb;
  wire [7:0] p34_array_index_2050060_comb;
  wire [7:0] p34_res7__438_comb;
  wire [7:0] p34_res7__440_comb;
  wire [7:0] p34_res7__442_comb;
  wire [7:0] p34_res7__444_comb;
  wire [7:0] p34_res7__446_comb;
  wire [127:0] p34_res__13_comb;
  assign p34_array_index_2050038_comb = p33_literal_2043918[p33_res7__424];
  assign p34_array_index_2050039_comb = p33_literal_2043920[p33_res7__422];
  assign p34_res7__434_comb = p33_literal_2043910[p33_res7__432] ^ p33_literal_2043912[p33_res7__430] ^ p33_literal_2043914[p33_res7__428] ^ p33_literal_2043916[p33_res7__426] ^ p34_array_index_2050038_comb ^ p34_array_index_2050039_comb ^ p33_res7__420 ^ p33_literal_2043923[p33_res7__418] ^ p33_res7__416 ^ p33_array_index_2049871 ^ p33_array_index_2049843 ^ p33_array_index_2049728 ^ p33_literal_2043914[p33_array_index_2049695] ^ p33_literal_2043912[p33_array_index_2049696] ^ p33_literal_2043910[p33_array_index_2049697] ^ p33_array_index_2049714;
  assign p34_array_index_2050050_comb = p33_literal_2043920[p33_res7__424];
  assign p34_res7__436_comb = p33_literal_2043910[p34_res7__434_comb] ^ p33_literal_2043912[p33_res7__432] ^ p33_literal_2043914[p33_res7__430] ^ p33_literal_2043916[p33_res7__428] ^ p33_literal_2043918[p33_res7__426] ^ p34_array_index_2050050_comb ^ p33_res7__422 ^ p33_literal_2043923[p33_res7__420] ^ p33_res7__418 ^ p33_array_index_2049884 ^ p33_array_index_2049857 ^ p33_array_index_2049828 ^ p33_array_index_2049710 ^ p33_literal_2043912[p33_array_index_2049695] ^ p33_literal_2043910[p33_array_index_2049696] ^ p33_array_index_2049697;
  assign p34_array_index_2050060_comb = p33_literal_2043920[p33_res7__426];
  assign p34_res7__438_comb = p33_literal_2043910[p34_res7__436_comb] ^ p33_literal_2043912[p34_res7__434_comb] ^ p33_literal_2043914[p33_res7__432] ^ p33_literal_2043916[p33_res7__430] ^ p33_literal_2043918[p33_res7__428] ^ p34_array_index_2050060_comb ^ p33_res7__424 ^ p33_literal_2043923[p33_res7__422] ^ p33_res7__420 ^ p33_array_index_2049896 ^ p33_array_index_2049870 ^ p33_array_index_2049842 ^ p33_array_index_2049727 ^ p33_literal_2043912[p33_array_index_2049694] ^ p33_literal_2043910[p33_array_index_2049695] ^ p33_array_index_2049696;
  assign p34_res7__440_comb = p33_literal_2043910[p34_res7__438_comb] ^ p33_literal_2043912[p34_res7__436_comb] ^ p33_literal_2043914[p34_res7__434_comb] ^ p33_literal_2043916[p33_res7__432] ^ p33_literal_2043918[p33_res7__430] ^ p33_literal_2043920[p33_res7__428] ^ p33_res7__426 ^ p33_literal_2043923[p33_res7__424] ^ p33_res7__422 ^ p33_array_index_2049908 ^ p33_array_index_2049883 ^ p33_array_index_2049856 ^ p33_array_index_2049827 ^ p33_array_index_2049709 ^ p33_literal_2043910[p33_array_index_2049694] ^ p33_array_index_2049695;
  assign p34_res7__442_comb = p33_literal_2043910[p34_res7__440_comb] ^ p33_literal_2043912[p34_res7__438_comb] ^ p33_literal_2043914[p34_res7__436_comb] ^ p33_literal_2043916[p34_res7__434_comb] ^ p33_literal_2043918[p33_res7__432] ^ p33_literal_2043920[p33_res7__430] ^ p33_res7__428 ^ p33_literal_2043923[p33_res7__426] ^ p33_res7__424 ^ p34_array_index_2050039_comb ^ p33_array_index_2049895 ^ p33_array_index_2049869 ^ p33_array_index_2049841 ^ p33_array_index_2049726 ^ p33_literal_2043910[p33_array_index_2049693] ^ p33_array_index_2049694;
  assign p34_res7__444_comb = p33_literal_2043910[p34_res7__442_comb] ^ p33_literal_2043912[p34_res7__440_comb] ^ p33_literal_2043914[p34_res7__438_comb] ^ p33_literal_2043916[p34_res7__436_comb] ^ p33_literal_2043918[p34_res7__434_comb] ^ p33_literal_2043920[p33_res7__432] ^ p33_res7__430 ^ p33_literal_2043923[p33_res7__428] ^ p33_res7__426 ^ p34_array_index_2050050_comb ^ p33_array_index_2049907 ^ p33_array_index_2049882 ^ p33_array_index_2049855 ^ p33_array_index_2049826 ^ p33_array_index_2049708 ^ p33_array_index_2049693;
  assign p34_res7__446_comb = p33_literal_2043910[p34_res7__444_comb] ^ p33_literal_2043912[p34_res7__442_comb] ^ p33_literal_2043914[p34_res7__440_comb] ^ p33_literal_2043916[p34_res7__438_comb] ^ p33_literal_2043918[p34_res7__436_comb] ^ p33_literal_2043920[p34_res7__434_comb] ^ p33_res7__432 ^ p33_literal_2043923[p33_res7__430] ^ p33_res7__428 ^ p34_array_index_2050060_comb ^ p34_array_index_2050038_comb ^ p33_array_index_2049894 ^ p33_array_index_2049868 ^ p33_array_index_2049840 ^ p33_array_index_2049725 ^ p33_array_index_2049692;
  assign p34_res__13_comb = {p34_res7__446_comb, p34_res7__444_comb, p34_res7__442_comb, p34_res7__440_comb, p34_res7__438_comb, p34_res7__436_comb, p34_res7__434_comb, p33_res7__432, p33_res7__430, p33_res7__428, p33_res7__426, p33_res7__424, p33_res7__422, p33_res7__420, p33_res7__418, p33_res7__416};

  // Registers for pipe stage 34:
  reg [127:0] p34_encoded;
  reg [127:0] p34_bit_slice_2043893;
  reg [127:0] p34_bit_slice_2044018;
  reg [127:0] p34_k3;
  reg [127:0] p34_k2;
  reg [127:0] p34_xor_2049240;
  reg [127:0] p34_xor_2049676;
  reg [127:0] p34_res__13;
  reg [7:0] p35_literal_2043896[256];
  reg [7:0] p35_literal_2043910[256];
  reg [7:0] p35_literal_2043912[256];
  reg [7:0] p35_literal_2043914[256];
  reg [7:0] p35_literal_2043916[256];
  reg [7:0] p35_literal_2043918[256];
  reg [7:0] p35_literal_2043920[256];
  reg [7:0] p35_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p34_encoded <= p33_encoded;
    p34_bit_slice_2043893 <= p33_bit_slice_2043893;
    p34_bit_slice_2044018 <= p33_bit_slice_2044018;
    p34_k3 <= p33_k3;
    p34_k2 <= p33_k2;
    p34_xor_2049240 <= p33_xor_2049240;
    p34_xor_2049676 <= p33_xor_2049676;
    p34_res__13 <= p34_res__13_comb;
    p35_literal_2043896 <= p34_literal_2043896;
    p35_literal_2043910 <= p34_literal_2043910;
    p35_literal_2043912 <= p34_literal_2043912;
    p35_literal_2043914 <= p34_literal_2043914;
    p35_literal_2043916 <= p34_literal_2043916;
    p35_literal_2043918 <= p34_literal_2043918;
    p35_literal_2043920 <= p34_literal_2043920;
    p35_literal_2043923 <= p34_literal_2043923;
  end

  // ===== Pipe stage 35:
  wire [127:0] p35_xor_2050132_comb;
  wire [127:0] p35_addedKey__46_comb;
  wire [7:0] p35_array_index_2050148_comb;
  wire [7:0] p35_array_index_2050149_comb;
  wire [7:0] p35_array_index_2050150_comb;
  wire [7:0] p35_array_index_2050151_comb;
  wire [7:0] p35_array_index_2050152_comb;
  wire [7:0] p35_array_index_2050153_comb;
  wire [7:0] p35_array_index_2050155_comb;
  wire [7:0] p35_array_index_2050157_comb;
  wire [7:0] p35_array_index_2050158_comb;
  wire [7:0] p35_array_index_2050159_comb;
  wire [7:0] p35_array_index_2050160_comb;
  wire [7:0] p35_array_index_2050161_comb;
  wire [7:0] p35_array_index_2050162_comb;
  wire [7:0] p35_array_index_2050164_comb;
  wire [7:0] p35_array_index_2050165_comb;
  wire [7:0] p35_array_index_2050166_comb;
  wire [7:0] p35_array_index_2050167_comb;
  wire [7:0] p35_array_index_2050168_comb;
  wire [7:0] p35_array_index_2050169_comb;
  wire [7:0] p35_array_index_2050170_comb;
  wire [7:0] p35_array_index_2050172_comb;
  wire [7:0] p35_res7__448_comb;
  wire [7:0] p35_array_index_2050181_comb;
  wire [7:0] p35_array_index_2050182_comb;
  wire [7:0] p35_array_index_2050183_comb;
  wire [7:0] p35_array_index_2050184_comb;
  wire [7:0] p35_array_index_2050185_comb;
  wire [7:0] p35_array_index_2050186_comb;
  wire [7:0] p35_res7__450_comb;
  wire [7:0] p35_array_index_2050196_comb;
  wire [7:0] p35_array_index_2050197_comb;
  wire [7:0] p35_array_index_2050198_comb;
  wire [7:0] p35_array_index_2050199_comb;
  wire [7:0] p35_array_index_2050200_comb;
  wire [7:0] p35_res7__452_comb;
  wire [7:0] p35_array_index_2050210_comb;
  wire [7:0] p35_array_index_2050211_comb;
  wire [7:0] p35_array_index_2050212_comb;
  wire [7:0] p35_array_index_2050213_comb;
  wire [7:0] p35_array_index_2050214_comb;
  wire [7:0] p35_res7__454_comb;
  wire [7:0] p35_array_index_2050225_comb;
  wire [7:0] p35_array_index_2050226_comb;
  wire [7:0] p35_array_index_2050227_comb;
  wire [7:0] p35_array_index_2050228_comb;
  wire [7:0] p35_res7__456_comb;
  wire [7:0] p35_array_index_2050238_comb;
  wire [7:0] p35_array_index_2050239_comb;
  wire [7:0] p35_array_index_2050240_comb;
  wire [7:0] p35_array_index_2050241_comb;
  wire [7:0] p35_res7__458_comb;
  assign p35_xor_2050132_comb = p34_res__13 ^ p34_xor_2049240;
  assign p35_addedKey__46_comb = p35_xor_2050132_comb ^ 128'h3fb1_b78b_213e_f327_fd0e_14f0_71b0_400f;
  assign p35_array_index_2050148_comb = p34_literal_2043896[p35_addedKey__46_comb[127:120]];
  assign p35_array_index_2050149_comb = p34_literal_2043896[p35_addedKey__46_comb[119:112]];
  assign p35_array_index_2050150_comb = p34_literal_2043896[p35_addedKey__46_comb[111:104]];
  assign p35_array_index_2050151_comb = p34_literal_2043896[p35_addedKey__46_comb[103:96]];
  assign p35_array_index_2050152_comb = p34_literal_2043896[p35_addedKey__46_comb[95:88]];
  assign p35_array_index_2050153_comb = p34_literal_2043896[p35_addedKey__46_comb[87:80]];
  assign p35_array_index_2050155_comb = p34_literal_2043896[p35_addedKey__46_comb[71:64]];
  assign p35_array_index_2050157_comb = p34_literal_2043896[p35_addedKey__46_comb[55:48]];
  assign p35_array_index_2050158_comb = p34_literal_2043896[p35_addedKey__46_comb[47:40]];
  assign p35_array_index_2050159_comb = p34_literal_2043896[p35_addedKey__46_comb[39:32]];
  assign p35_array_index_2050160_comb = p34_literal_2043896[p35_addedKey__46_comb[31:24]];
  assign p35_array_index_2050161_comb = p34_literal_2043896[p35_addedKey__46_comb[23:16]];
  assign p35_array_index_2050162_comb = p34_literal_2043896[p35_addedKey__46_comb[15:8]];
  assign p35_array_index_2050164_comb = p34_literal_2043910[p35_array_index_2050148_comb];
  assign p35_array_index_2050165_comb = p34_literal_2043912[p35_array_index_2050149_comb];
  assign p35_array_index_2050166_comb = p34_literal_2043914[p35_array_index_2050150_comb];
  assign p35_array_index_2050167_comb = p34_literal_2043916[p35_array_index_2050151_comb];
  assign p35_array_index_2050168_comb = p34_literal_2043918[p35_array_index_2050152_comb];
  assign p35_array_index_2050169_comb = p34_literal_2043920[p35_array_index_2050153_comb];
  assign p35_array_index_2050170_comb = p34_literal_2043896[p35_addedKey__46_comb[79:72]];
  assign p35_array_index_2050172_comb = p34_literal_2043896[p35_addedKey__46_comb[63:56]];
  assign p35_res7__448_comb = p35_array_index_2050164_comb ^ p35_array_index_2050165_comb ^ p35_array_index_2050166_comb ^ p35_array_index_2050167_comb ^ p35_array_index_2050168_comb ^ p35_array_index_2050169_comb ^ p35_array_index_2050170_comb ^ p34_literal_2043923[p35_array_index_2050155_comb] ^ p35_array_index_2050172_comb ^ p34_literal_2043920[p35_array_index_2050157_comb] ^ p34_literal_2043918[p35_array_index_2050158_comb] ^ p34_literal_2043916[p35_array_index_2050159_comb] ^ p34_literal_2043914[p35_array_index_2050160_comb] ^ p34_literal_2043912[p35_array_index_2050161_comb] ^ p34_literal_2043910[p35_array_index_2050162_comb] ^ p34_literal_2043896[p35_addedKey__46_comb[7:0]];
  assign p35_array_index_2050181_comb = p34_literal_2043910[p35_res7__448_comb];
  assign p35_array_index_2050182_comb = p34_literal_2043912[p35_array_index_2050148_comb];
  assign p35_array_index_2050183_comb = p34_literal_2043914[p35_array_index_2050149_comb];
  assign p35_array_index_2050184_comb = p34_literal_2043916[p35_array_index_2050150_comb];
  assign p35_array_index_2050185_comb = p34_literal_2043918[p35_array_index_2050151_comb];
  assign p35_array_index_2050186_comb = p34_literal_2043920[p35_array_index_2050152_comb];
  assign p35_res7__450_comb = p35_array_index_2050181_comb ^ p35_array_index_2050182_comb ^ p35_array_index_2050183_comb ^ p35_array_index_2050184_comb ^ p35_array_index_2050185_comb ^ p35_array_index_2050186_comb ^ p35_array_index_2050153_comb ^ p34_literal_2043923[p35_array_index_2050170_comb] ^ p35_array_index_2050155_comb ^ p34_literal_2043920[p35_array_index_2050172_comb] ^ p34_literal_2043918[p35_array_index_2050157_comb] ^ p34_literal_2043916[p35_array_index_2050158_comb] ^ p34_literal_2043914[p35_array_index_2050159_comb] ^ p34_literal_2043912[p35_array_index_2050160_comb] ^ p34_literal_2043910[p35_array_index_2050161_comb] ^ p35_array_index_2050162_comb;
  assign p35_array_index_2050196_comb = p34_literal_2043912[p35_res7__448_comb];
  assign p35_array_index_2050197_comb = p34_literal_2043914[p35_array_index_2050148_comb];
  assign p35_array_index_2050198_comb = p34_literal_2043916[p35_array_index_2050149_comb];
  assign p35_array_index_2050199_comb = p34_literal_2043918[p35_array_index_2050150_comb];
  assign p35_array_index_2050200_comb = p34_literal_2043920[p35_array_index_2050151_comb];
  assign p35_res7__452_comb = p34_literal_2043910[p35_res7__450_comb] ^ p35_array_index_2050196_comb ^ p35_array_index_2050197_comb ^ p35_array_index_2050198_comb ^ p35_array_index_2050199_comb ^ p35_array_index_2050200_comb ^ p35_array_index_2050152_comb ^ p34_literal_2043923[p35_array_index_2050153_comb] ^ p35_array_index_2050170_comb ^ p34_literal_2043920[p35_array_index_2050155_comb] ^ p34_literal_2043918[p35_array_index_2050172_comb] ^ p34_literal_2043916[p35_array_index_2050157_comb] ^ p34_literal_2043914[p35_array_index_2050158_comb] ^ p34_literal_2043912[p35_array_index_2050159_comb] ^ p34_literal_2043910[p35_array_index_2050160_comb] ^ p35_array_index_2050161_comb;
  assign p35_array_index_2050210_comb = p34_literal_2043912[p35_res7__450_comb];
  assign p35_array_index_2050211_comb = p34_literal_2043914[p35_res7__448_comb];
  assign p35_array_index_2050212_comb = p34_literal_2043916[p35_array_index_2050148_comb];
  assign p35_array_index_2050213_comb = p34_literal_2043918[p35_array_index_2050149_comb];
  assign p35_array_index_2050214_comb = p34_literal_2043920[p35_array_index_2050150_comb];
  assign p35_res7__454_comb = p34_literal_2043910[p35_res7__452_comb] ^ p35_array_index_2050210_comb ^ p35_array_index_2050211_comb ^ p35_array_index_2050212_comb ^ p35_array_index_2050213_comb ^ p35_array_index_2050214_comb ^ p35_array_index_2050151_comb ^ p34_literal_2043923[p35_array_index_2050152_comb] ^ p35_array_index_2050153_comb ^ p34_literal_2043920[p35_array_index_2050170_comb] ^ p34_literal_2043918[p35_array_index_2050155_comb] ^ p34_literal_2043916[p35_array_index_2050172_comb] ^ p34_literal_2043914[p35_array_index_2050157_comb] ^ p34_literal_2043912[p35_array_index_2050158_comb] ^ p34_literal_2043910[p35_array_index_2050159_comb] ^ p35_array_index_2050160_comb;
  assign p35_array_index_2050225_comb = p34_literal_2043914[p35_res7__450_comb];
  assign p35_array_index_2050226_comb = p34_literal_2043916[p35_res7__448_comb];
  assign p35_array_index_2050227_comb = p34_literal_2043918[p35_array_index_2050148_comb];
  assign p35_array_index_2050228_comb = p34_literal_2043920[p35_array_index_2050149_comb];
  assign p35_res7__456_comb = p34_literal_2043910[p35_res7__454_comb] ^ p34_literal_2043912[p35_res7__452_comb] ^ p35_array_index_2050225_comb ^ p35_array_index_2050226_comb ^ p35_array_index_2050227_comb ^ p35_array_index_2050228_comb ^ p35_array_index_2050150_comb ^ p34_literal_2043923[p35_array_index_2050151_comb] ^ p35_array_index_2050152_comb ^ p35_array_index_2050169_comb ^ p34_literal_2043918[p35_array_index_2050170_comb] ^ p34_literal_2043916[p35_array_index_2050155_comb] ^ p34_literal_2043914[p35_array_index_2050172_comb] ^ p34_literal_2043912[p35_array_index_2050157_comb] ^ p34_literal_2043910[p35_array_index_2050158_comb] ^ p35_array_index_2050159_comb;
  assign p35_array_index_2050238_comb = p34_literal_2043914[p35_res7__452_comb];
  assign p35_array_index_2050239_comb = p34_literal_2043916[p35_res7__450_comb];
  assign p35_array_index_2050240_comb = p34_literal_2043918[p35_res7__448_comb];
  assign p35_array_index_2050241_comb = p34_literal_2043920[p35_array_index_2050148_comb];
  assign p35_res7__458_comb = p34_literal_2043910[p35_res7__456_comb] ^ p34_literal_2043912[p35_res7__454_comb] ^ p35_array_index_2050238_comb ^ p35_array_index_2050239_comb ^ p35_array_index_2050240_comb ^ p35_array_index_2050241_comb ^ p35_array_index_2050149_comb ^ p34_literal_2043923[p35_array_index_2050150_comb] ^ p35_array_index_2050151_comb ^ p35_array_index_2050186_comb ^ p34_literal_2043918[p35_array_index_2050153_comb] ^ p34_literal_2043916[p35_array_index_2050170_comb] ^ p34_literal_2043914[p35_array_index_2050155_comb] ^ p34_literal_2043912[p35_array_index_2050172_comb] ^ p34_literal_2043910[p35_array_index_2050157_comb] ^ p35_array_index_2050158_comb;

  // Registers for pipe stage 35:
  reg [127:0] p35_encoded;
  reg [127:0] p35_bit_slice_2043893;
  reg [127:0] p35_bit_slice_2044018;
  reg [127:0] p35_k3;
  reg [127:0] p35_k2;
  reg [127:0] p35_xor_2049676;
  reg [127:0] p35_xor_2050132;
  reg [7:0] p35_array_index_2050148;
  reg [7:0] p35_array_index_2050149;
  reg [7:0] p35_array_index_2050150;
  reg [7:0] p35_array_index_2050151;
  reg [7:0] p35_array_index_2050152;
  reg [7:0] p35_array_index_2050153;
  reg [7:0] p35_array_index_2050155;
  reg [7:0] p35_array_index_2050157;
  reg [7:0] p35_array_index_2050164;
  reg [7:0] p35_array_index_2050165;
  reg [7:0] p35_array_index_2050166;
  reg [7:0] p35_array_index_2050167;
  reg [7:0] p35_array_index_2050168;
  reg [7:0] p35_array_index_2050170;
  reg [7:0] p35_array_index_2050172;
  reg [7:0] p35_res7__448;
  reg [7:0] p35_array_index_2050181;
  reg [7:0] p35_array_index_2050182;
  reg [7:0] p35_array_index_2050183;
  reg [7:0] p35_array_index_2050184;
  reg [7:0] p35_array_index_2050185;
  reg [7:0] p35_res7__450;
  reg [7:0] p35_array_index_2050196;
  reg [7:0] p35_array_index_2050197;
  reg [7:0] p35_array_index_2050198;
  reg [7:0] p35_array_index_2050199;
  reg [7:0] p35_array_index_2050200;
  reg [7:0] p35_res7__452;
  reg [7:0] p35_array_index_2050210;
  reg [7:0] p35_array_index_2050211;
  reg [7:0] p35_array_index_2050212;
  reg [7:0] p35_array_index_2050213;
  reg [7:0] p35_array_index_2050214;
  reg [7:0] p35_res7__454;
  reg [7:0] p35_array_index_2050225;
  reg [7:0] p35_array_index_2050226;
  reg [7:0] p35_array_index_2050227;
  reg [7:0] p35_array_index_2050228;
  reg [7:0] p35_res7__456;
  reg [7:0] p35_array_index_2050238;
  reg [7:0] p35_array_index_2050239;
  reg [7:0] p35_array_index_2050240;
  reg [7:0] p35_array_index_2050241;
  reg [7:0] p35_res7__458;
  reg [7:0] p36_literal_2043896[256];
  reg [7:0] p36_literal_2043910[256];
  reg [7:0] p36_literal_2043912[256];
  reg [7:0] p36_literal_2043914[256];
  reg [7:0] p36_literal_2043916[256];
  reg [7:0] p36_literal_2043918[256];
  reg [7:0] p36_literal_2043920[256];
  reg [7:0] p36_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p35_encoded <= p34_encoded;
    p35_bit_slice_2043893 <= p34_bit_slice_2043893;
    p35_bit_slice_2044018 <= p34_bit_slice_2044018;
    p35_k3 <= p34_k3;
    p35_k2 <= p34_k2;
    p35_xor_2049676 <= p34_xor_2049676;
    p35_xor_2050132 <= p35_xor_2050132_comb;
    p35_array_index_2050148 <= p35_array_index_2050148_comb;
    p35_array_index_2050149 <= p35_array_index_2050149_comb;
    p35_array_index_2050150 <= p35_array_index_2050150_comb;
    p35_array_index_2050151 <= p35_array_index_2050151_comb;
    p35_array_index_2050152 <= p35_array_index_2050152_comb;
    p35_array_index_2050153 <= p35_array_index_2050153_comb;
    p35_array_index_2050155 <= p35_array_index_2050155_comb;
    p35_array_index_2050157 <= p35_array_index_2050157_comb;
    p35_array_index_2050164 <= p35_array_index_2050164_comb;
    p35_array_index_2050165 <= p35_array_index_2050165_comb;
    p35_array_index_2050166 <= p35_array_index_2050166_comb;
    p35_array_index_2050167 <= p35_array_index_2050167_comb;
    p35_array_index_2050168 <= p35_array_index_2050168_comb;
    p35_array_index_2050170 <= p35_array_index_2050170_comb;
    p35_array_index_2050172 <= p35_array_index_2050172_comb;
    p35_res7__448 <= p35_res7__448_comb;
    p35_array_index_2050181 <= p35_array_index_2050181_comb;
    p35_array_index_2050182 <= p35_array_index_2050182_comb;
    p35_array_index_2050183 <= p35_array_index_2050183_comb;
    p35_array_index_2050184 <= p35_array_index_2050184_comb;
    p35_array_index_2050185 <= p35_array_index_2050185_comb;
    p35_res7__450 <= p35_res7__450_comb;
    p35_array_index_2050196 <= p35_array_index_2050196_comb;
    p35_array_index_2050197 <= p35_array_index_2050197_comb;
    p35_array_index_2050198 <= p35_array_index_2050198_comb;
    p35_array_index_2050199 <= p35_array_index_2050199_comb;
    p35_array_index_2050200 <= p35_array_index_2050200_comb;
    p35_res7__452 <= p35_res7__452_comb;
    p35_array_index_2050210 <= p35_array_index_2050210_comb;
    p35_array_index_2050211 <= p35_array_index_2050211_comb;
    p35_array_index_2050212 <= p35_array_index_2050212_comb;
    p35_array_index_2050213 <= p35_array_index_2050213_comb;
    p35_array_index_2050214 <= p35_array_index_2050214_comb;
    p35_res7__454 <= p35_res7__454_comb;
    p35_array_index_2050225 <= p35_array_index_2050225_comb;
    p35_array_index_2050226 <= p35_array_index_2050226_comb;
    p35_array_index_2050227 <= p35_array_index_2050227_comb;
    p35_array_index_2050228 <= p35_array_index_2050228_comb;
    p35_res7__456 <= p35_res7__456_comb;
    p35_array_index_2050238 <= p35_array_index_2050238_comb;
    p35_array_index_2050239 <= p35_array_index_2050239_comb;
    p35_array_index_2050240 <= p35_array_index_2050240_comb;
    p35_array_index_2050241 <= p35_array_index_2050241_comb;
    p35_res7__458 <= p35_res7__458_comb;
    p36_literal_2043896 <= p35_literal_2043896;
    p36_literal_2043910 <= p35_literal_2043910;
    p36_literal_2043912 <= p35_literal_2043912;
    p36_literal_2043914 <= p35_literal_2043914;
    p36_literal_2043916 <= p35_literal_2043916;
    p36_literal_2043918 <= p35_literal_2043918;
    p36_literal_2043920 <= p35_literal_2043920;
    p36_literal_2043923 <= p35_literal_2043923;
  end

  // ===== Pipe stage 36:
  wire [7:0] p36_array_index_2050370_comb;
  wire [7:0] p36_array_index_2050371_comb;
  wire [7:0] p36_array_index_2050372_comb;
  wire [7:0] p36_res7__460_comb;
  wire [7:0] p36_array_index_2050382_comb;
  wire [7:0] p36_array_index_2050383_comb;
  wire [7:0] p36_array_index_2050384_comb;
  wire [7:0] p36_res7__462_comb;
  wire [7:0] p36_array_index_2050395_comb;
  wire [7:0] p36_array_index_2050396_comb;
  wire [7:0] p36_res7__464_comb;
  wire [7:0] p36_array_index_2050406_comb;
  wire [7:0] p36_array_index_2050407_comb;
  wire [7:0] p36_res7__466_comb;
  wire [7:0] p36_array_index_2050418_comb;
  wire [7:0] p36_res7__468_comb;
  wire [7:0] p36_array_index_2050428_comb;
  wire [7:0] p36_res7__470_comb;
  wire [7:0] p36_res7__472_comb;
  assign p36_array_index_2050370_comb = p35_literal_2043916[p35_res7__452];
  assign p36_array_index_2050371_comb = p35_literal_2043918[p35_res7__450];
  assign p36_array_index_2050372_comb = p35_literal_2043920[p35_res7__448];
  assign p36_res7__460_comb = p35_literal_2043910[p35_res7__458] ^ p35_literal_2043912[p35_res7__456] ^ p35_literal_2043914[p35_res7__454] ^ p36_array_index_2050370_comb ^ p36_array_index_2050371_comb ^ p36_array_index_2050372_comb ^ p35_array_index_2050148 ^ p35_literal_2043923[p35_array_index_2050149] ^ p35_array_index_2050150 ^ p35_array_index_2050200 ^ p35_array_index_2050168 ^ p35_literal_2043916[p35_array_index_2050153] ^ p35_literal_2043914[p35_array_index_2050170] ^ p35_literal_2043912[p35_array_index_2050155] ^ p35_literal_2043910[p35_array_index_2050172] ^ p35_array_index_2050157;
  assign p36_array_index_2050382_comb = p35_literal_2043916[p35_res7__454];
  assign p36_array_index_2050383_comb = p35_literal_2043918[p35_res7__452];
  assign p36_array_index_2050384_comb = p35_literal_2043920[p35_res7__450];
  assign p36_res7__462_comb = p35_literal_2043910[p36_res7__460_comb] ^ p35_literal_2043912[p35_res7__458] ^ p35_literal_2043914[p35_res7__456] ^ p36_array_index_2050382_comb ^ p36_array_index_2050383_comb ^ p36_array_index_2050384_comb ^ p35_res7__448 ^ p35_literal_2043923[p35_array_index_2050148] ^ p35_array_index_2050149 ^ p35_array_index_2050214 ^ p35_array_index_2050185 ^ p35_literal_2043916[p35_array_index_2050152] ^ p35_literal_2043914[p35_array_index_2050153] ^ p35_literal_2043912[p35_array_index_2050170] ^ p35_literal_2043910[p35_array_index_2050155] ^ p35_array_index_2050172;
  assign p36_array_index_2050395_comb = p35_literal_2043918[p35_res7__454];
  assign p36_array_index_2050396_comb = p35_literal_2043920[p35_res7__452];
  assign p36_res7__464_comb = p35_literal_2043910[p36_res7__462_comb] ^ p35_literal_2043912[p36_res7__460_comb] ^ p35_literal_2043914[p35_res7__458] ^ p35_literal_2043916[p35_res7__456] ^ p36_array_index_2050395_comb ^ p36_array_index_2050396_comb ^ p35_res7__450 ^ p35_literal_2043923[p35_res7__448] ^ p35_array_index_2050148 ^ p35_array_index_2050228 ^ p35_array_index_2050199 ^ p35_array_index_2050167 ^ p35_literal_2043914[p35_array_index_2050152] ^ p35_literal_2043912[p35_array_index_2050153] ^ p35_literal_2043910[p35_array_index_2050170] ^ p35_array_index_2050155;
  assign p36_array_index_2050406_comb = p35_literal_2043918[p35_res7__456];
  assign p36_array_index_2050407_comb = p35_literal_2043920[p35_res7__454];
  assign p36_res7__466_comb = p35_literal_2043910[p36_res7__464_comb] ^ p35_literal_2043912[p36_res7__462_comb] ^ p35_literal_2043914[p36_res7__460_comb] ^ p35_literal_2043916[p35_res7__458] ^ p36_array_index_2050406_comb ^ p36_array_index_2050407_comb ^ p35_res7__452 ^ p35_literal_2043923[p35_res7__450] ^ p35_res7__448 ^ p35_array_index_2050241 ^ p35_array_index_2050213 ^ p35_array_index_2050184 ^ p35_literal_2043914[p35_array_index_2050151] ^ p35_literal_2043912[p35_array_index_2050152] ^ p35_literal_2043910[p35_array_index_2050153] ^ p35_array_index_2050170;
  assign p36_array_index_2050418_comb = p35_literal_2043920[p35_res7__456];
  assign p36_res7__468_comb = p35_literal_2043910[p36_res7__466_comb] ^ p35_literal_2043912[p36_res7__464_comb] ^ p35_literal_2043914[p36_res7__462_comb] ^ p35_literal_2043916[p36_res7__460_comb] ^ p35_literal_2043918[p35_res7__458] ^ p36_array_index_2050418_comb ^ p35_res7__454 ^ p35_literal_2043923[p35_res7__452] ^ p35_res7__450 ^ p36_array_index_2050372_comb ^ p35_array_index_2050227 ^ p35_array_index_2050198 ^ p35_array_index_2050166 ^ p35_literal_2043912[p35_array_index_2050151] ^ p35_literal_2043910[p35_array_index_2050152] ^ p35_array_index_2050153;
  assign p36_array_index_2050428_comb = p35_literal_2043920[p35_res7__458];
  assign p36_res7__470_comb = p35_literal_2043910[p36_res7__468_comb] ^ p35_literal_2043912[p36_res7__466_comb] ^ p35_literal_2043914[p36_res7__464_comb] ^ p35_literal_2043916[p36_res7__462_comb] ^ p35_literal_2043918[p36_res7__460_comb] ^ p36_array_index_2050428_comb ^ p35_res7__456 ^ p35_literal_2043923[p35_res7__454] ^ p35_res7__452 ^ p36_array_index_2050384_comb ^ p35_array_index_2050240 ^ p35_array_index_2050212 ^ p35_array_index_2050183 ^ p35_literal_2043912[p35_array_index_2050150] ^ p35_literal_2043910[p35_array_index_2050151] ^ p35_array_index_2050152;
  assign p36_res7__472_comb = p35_literal_2043910[p36_res7__470_comb] ^ p35_literal_2043912[p36_res7__468_comb] ^ p35_literal_2043914[p36_res7__466_comb] ^ p35_literal_2043916[p36_res7__464_comb] ^ p35_literal_2043918[p36_res7__462_comb] ^ p35_literal_2043920[p36_res7__460_comb] ^ p35_res7__458 ^ p35_literal_2043923[p35_res7__456] ^ p35_res7__454 ^ p36_array_index_2050396_comb ^ p36_array_index_2050371_comb ^ p35_array_index_2050226 ^ p35_array_index_2050197 ^ p35_array_index_2050165 ^ p35_literal_2043910[p35_array_index_2050150] ^ p35_array_index_2050151;

  // Registers for pipe stage 36:
  reg [127:0] p36_encoded;
  reg [127:0] p36_bit_slice_2043893;
  reg [127:0] p36_bit_slice_2044018;
  reg [127:0] p36_k3;
  reg [127:0] p36_k2;
  reg [127:0] p36_xor_2049676;
  reg [127:0] p36_xor_2050132;
  reg [7:0] p36_array_index_2050148;
  reg [7:0] p36_array_index_2050149;
  reg [7:0] p36_array_index_2050150;
  reg [7:0] p36_array_index_2050164;
  reg [7:0] p36_res7__448;
  reg [7:0] p36_array_index_2050181;
  reg [7:0] p36_array_index_2050182;
  reg [7:0] p36_res7__450;
  reg [7:0] p36_array_index_2050196;
  reg [7:0] p36_res7__452;
  reg [7:0] p36_array_index_2050210;
  reg [7:0] p36_array_index_2050211;
  reg [7:0] p36_res7__454;
  reg [7:0] p36_array_index_2050225;
  reg [7:0] p36_res7__456;
  reg [7:0] p36_array_index_2050238;
  reg [7:0] p36_array_index_2050239;
  reg [7:0] p36_res7__458;
  reg [7:0] p36_array_index_2050370;
  reg [7:0] p36_res7__460;
  reg [7:0] p36_array_index_2050382;
  reg [7:0] p36_array_index_2050383;
  reg [7:0] p36_res7__462;
  reg [7:0] p36_array_index_2050395;
  reg [7:0] p36_res7__464;
  reg [7:0] p36_array_index_2050406;
  reg [7:0] p36_array_index_2050407;
  reg [7:0] p36_res7__466;
  reg [7:0] p36_array_index_2050418;
  reg [7:0] p36_res7__468;
  reg [7:0] p36_array_index_2050428;
  reg [7:0] p36_res7__470;
  reg [7:0] p36_res7__472;
  reg [7:0] p37_literal_2043896[256];
  reg [7:0] p37_literal_2043910[256];
  reg [7:0] p37_literal_2043912[256];
  reg [7:0] p37_literal_2043914[256];
  reg [7:0] p37_literal_2043916[256];
  reg [7:0] p37_literal_2043918[256];
  reg [7:0] p37_literal_2043920[256];
  reg [7:0] p37_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p36_encoded <= p35_encoded;
    p36_bit_slice_2043893 <= p35_bit_slice_2043893;
    p36_bit_slice_2044018 <= p35_bit_slice_2044018;
    p36_k3 <= p35_k3;
    p36_k2 <= p35_k2;
    p36_xor_2049676 <= p35_xor_2049676;
    p36_xor_2050132 <= p35_xor_2050132;
    p36_array_index_2050148 <= p35_array_index_2050148;
    p36_array_index_2050149 <= p35_array_index_2050149;
    p36_array_index_2050150 <= p35_array_index_2050150;
    p36_array_index_2050164 <= p35_array_index_2050164;
    p36_res7__448 <= p35_res7__448;
    p36_array_index_2050181 <= p35_array_index_2050181;
    p36_array_index_2050182 <= p35_array_index_2050182;
    p36_res7__450 <= p35_res7__450;
    p36_array_index_2050196 <= p35_array_index_2050196;
    p36_res7__452 <= p35_res7__452;
    p36_array_index_2050210 <= p35_array_index_2050210;
    p36_array_index_2050211 <= p35_array_index_2050211;
    p36_res7__454 <= p35_res7__454;
    p36_array_index_2050225 <= p35_array_index_2050225;
    p36_res7__456 <= p35_res7__456;
    p36_array_index_2050238 <= p35_array_index_2050238;
    p36_array_index_2050239 <= p35_array_index_2050239;
    p36_res7__458 <= p35_res7__458;
    p36_array_index_2050370 <= p36_array_index_2050370_comb;
    p36_res7__460 <= p36_res7__460_comb;
    p36_array_index_2050382 <= p36_array_index_2050382_comb;
    p36_array_index_2050383 <= p36_array_index_2050383_comb;
    p36_res7__462 <= p36_res7__462_comb;
    p36_array_index_2050395 <= p36_array_index_2050395_comb;
    p36_res7__464 <= p36_res7__464_comb;
    p36_array_index_2050406 <= p36_array_index_2050406_comb;
    p36_array_index_2050407 <= p36_array_index_2050407_comb;
    p36_res7__466 <= p36_res7__466_comb;
    p36_array_index_2050418 <= p36_array_index_2050418_comb;
    p36_res7__468 <= p36_res7__468_comb;
    p36_array_index_2050428 <= p36_array_index_2050428_comb;
    p36_res7__470 <= p36_res7__470_comb;
    p36_res7__472 <= p36_res7__472_comb;
    p37_literal_2043896 <= p36_literal_2043896;
    p37_literal_2043910 <= p36_literal_2043910;
    p37_literal_2043912 <= p36_literal_2043912;
    p37_literal_2043914 <= p36_literal_2043914;
    p37_literal_2043916 <= p36_literal_2043916;
    p37_literal_2043918 <= p36_literal_2043918;
    p37_literal_2043920 <= p36_literal_2043920;
    p37_literal_2043923 <= p36_literal_2043923;
  end

  // ===== Pipe stage 37:
  wire [7:0] p37_res7__474_comb;
  wire [7:0] p37_res7__476_comb;
  wire [7:0] p37_res7__478_comb;
  wire [127:0] p37_res__14_comb;
  wire [127:0] p37_k5_comb;
  wire [127:0] p37_addedKey__47_comb;
  wire [7:0] p37_array_index_2050580_comb;
  wire [7:0] p37_array_index_2050581_comb;
  wire [7:0] p37_array_index_2050582_comb;
  wire [7:0] p37_array_index_2050583_comb;
  wire [7:0] p37_array_index_2050584_comb;
  wire [7:0] p37_array_index_2050585_comb;
  wire [7:0] p37_array_index_2050587_comb;
  wire [7:0] p37_array_index_2050589_comb;
  wire [7:0] p37_array_index_2050590_comb;
  wire [7:0] p37_array_index_2050591_comb;
  wire [7:0] p37_array_index_2050592_comb;
  wire [7:0] p37_array_index_2050593_comb;
  wire [7:0] p37_array_index_2050594_comb;
  wire [7:0] p37_array_index_2050596_comb;
  wire [7:0] p37_array_index_2050597_comb;
  wire [7:0] p37_array_index_2050598_comb;
  wire [7:0] p37_array_index_2050599_comb;
  wire [7:0] p37_array_index_2050600_comb;
  wire [7:0] p37_array_index_2050601_comb;
  wire [7:0] p37_array_index_2050602_comb;
  wire [7:0] p37_array_index_2050604_comb;
  wire [7:0] p37_res7__480_comb;
  wire [7:0] p37_array_index_2050613_comb;
  wire [7:0] p37_array_index_2050614_comb;
  wire [7:0] p37_array_index_2050615_comb;
  wire [7:0] p37_array_index_2050616_comb;
  wire [7:0] p37_array_index_2050617_comb;
  wire [7:0] p37_array_index_2050618_comb;
  wire [7:0] p37_res7__482_comb;
  wire [7:0] p37_array_index_2050628_comb;
  wire [7:0] p37_array_index_2050629_comb;
  wire [7:0] p37_array_index_2050630_comb;
  wire [7:0] p37_array_index_2050631_comb;
  wire [7:0] p37_array_index_2050632_comb;
  wire [7:0] p37_res7__484_comb;
  assign p37_res7__474_comb = p36_literal_2043910[p36_res7__472] ^ p36_literal_2043912[p36_res7__470] ^ p36_literal_2043914[p36_res7__468] ^ p36_literal_2043916[p36_res7__466] ^ p36_literal_2043918[p36_res7__464] ^ p36_literal_2043920[p36_res7__462] ^ p36_res7__460 ^ p36_literal_2043923[p36_res7__458] ^ p36_res7__456 ^ p36_array_index_2050407 ^ p36_array_index_2050383 ^ p36_array_index_2050239 ^ p36_array_index_2050211 ^ p36_array_index_2050182 ^ p36_literal_2043910[p36_array_index_2050149] ^ p36_array_index_2050150;
  assign p37_res7__476_comb = p36_literal_2043910[p37_res7__474_comb] ^ p36_literal_2043912[p36_res7__472] ^ p36_literal_2043914[p36_res7__470] ^ p36_literal_2043916[p36_res7__468] ^ p36_literal_2043918[p36_res7__466] ^ p36_literal_2043920[p36_res7__464] ^ p36_res7__462 ^ p36_literal_2043923[p36_res7__460] ^ p36_res7__458 ^ p36_array_index_2050418 ^ p36_array_index_2050395 ^ p36_array_index_2050370 ^ p36_array_index_2050225 ^ p36_array_index_2050196 ^ p36_array_index_2050164 ^ p36_array_index_2050149;
  assign p37_res7__478_comb = p36_literal_2043910[p37_res7__476_comb] ^ p36_literal_2043912[p37_res7__474_comb] ^ p36_literal_2043914[p36_res7__472] ^ p36_literal_2043916[p36_res7__470] ^ p36_literal_2043918[p36_res7__468] ^ p36_literal_2043920[p36_res7__466] ^ p36_res7__464 ^ p36_literal_2043923[p36_res7__462] ^ p36_res7__460 ^ p36_array_index_2050428 ^ p36_array_index_2050406 ^ p36_array_index_2050382 ^ p36_array_index_2050238 ^ p36_array_index_2050210 ^ p36_array_index_2050181 ^ p36_array_index_2050148;
  assign p37_res__14_comb = {p37_res7__478_comb, p37_res7__476_comb, p37_res7__474_comb, p36_res7__472, p36_res7__470, p36_res7__468, p36_res7__466, p36_res7__464, p36_res7__462, p36_res7__460, p36_res7__458, p36_res7__456, p36_res7__454, p36_res7__452, p36_res7__450, p36_res7__448};
  assign p37_k5_comb = p37_res__14_comb ^ p36_xor_2049676;
  assign p37_addedKey__47_comb = p37_k5_comb ^ 128'h2fb2_6c2c_0f0a_acd1_9935_81c3_4e97_5410;
  assign p37_array_index_2050580_comb = p36_literal_2043896[p37_addedKey__47_comb[127:120]];
  assign p37_array_index_2050581_comb = p36_literal_2043896[p37_addedKey__47_comb[119:112]];
  assign p37_array_index_2050582_comb = p36_literal_2043896[p37_addedKey__47_comb[111:104]];
  assign p37_array_index_2050583_comb = p36_literal_2043896[p37_addedKey__47_comb[103:96]];
  assign p37_array_index_2050584_comb = p36_literal_2043896[p37_addedKey__47_comb[95:88]];
  assign p37_array_index_2050585_comb = p36_literal_2043896[p37_addedKey__47_comb[87:80]];
  assign p37_array_index_2050587_comb = p36_literal_2043896[p37_addedKey__47_comb[71:64]];
  assign p37_array_index_2050589_comb = p36_literal_2043896[p37_addedKey__47_comb[55:48]];
  assign p37_array_index_2050590_comb = p36_literal_2043896[p37_addedKey__47_comb[47:40]];
  assign p37_array_index_2050591_comb = p36_literal_2043896[p37_addedKey__47_comb[39:32]];
  assign p37_array_index_2050592_comb = p36_literal_2043896[p37_addedKey__47_comb[31:24]];
  assign p37_array_index_2050593_comb = p36_literal_2043896[p37_addedKey__47_comb[23:16]];
  assign p37_array_index_2050594_comb = p36_literal_2043896[p37_addedKey__47_comb[15:8]];
  assign p37_array_index_2050596_comb = p36_literal_2043910[p37_array_index_2050580_comb];
  assign p37_array_index_2050597_comb = p36_literal_2043912[p37_array_index_2050581_comb];
  assign p37_array_index_2050598_comb = p36_literal_2043914[p37_array_index_2050582_comb];
  assign p37_array_index_2050599_comb = p36_literal_2043916[p37_array_index_2050583_comb];
  assign p37_array_index_2050600_comb = p36_literal_2043918[p37_array_index_2050584_comb];
  assign p37_array_index_2050601_comb = p36_literal_2043920[p37_array_index_2050585_comb];
  assign p37_array_index_2050602_comb = p36_literal_2043896[p37_addedKey__47_comb[79:72]];
  assign p37_array_index_2050604_comb = p36_literal_2043896[p37_addedKey__47_comb[63:56]];
  assign p37_res7__480_comb = p37_array_index_2050596_comb ^ p37_array_index_2050597_comb ^ p37_array_index_2050598_comb ^ p37_array_index_2050599_comb ^ p37_array_index_2050600_comb ^ p37_array_index_2050601_comb ^ p37_array_index_2050602_comb ^ p36_literal_2043923[p37_array_index_2050587_comb] ^ p37_array_index_2050604_comb ^ p36_literal_2043920[p37_array_index_2050589_comb] ^ p36_literal_2043918[p37_array_index_2050590_comb] ^ p36_literal_2043916[p37_array_index_2050591_comb] ^ p36_literal_2043914[p37_array_index_2050592_comb] ^ p36_literal_2043912[p37_array_index_2050593_comb] ^ p36_literal_2043910[p37_array_index_2050594_comb] ^ p36_literal_2043896[p37_addedKey__47_comb[7:0]];
  assign p37_array_index_2050613_comb = p36_literal_2043910[p37_res7__480_comb];
  assign p37_array_index_2050614_comb = p36_literal_2043912[p37_array_index_2050580_comb];
  assign p37_array_index_2050615_comb = p36_literal_2043914[p37_array_index_2050581_comb];
  assign p37_array_index_2050616_comb = p36_literal_2043916[p37_array_index_2050582_comb];
  assign p37_array_index_2050617_comb = p36_literal_2043918[p37_array_index_2050583_comb];
  assign p37_array_index_2050618_comb = p36_literal_2043920[p37_array_index_2050584_comb];
  assign p37_res7__482_comb = p37_array_index_2050613_comb ^ p37_array_index_2050614_comb ^ p37_array_index_2050615_comb ^ p37_array_index_2050616_comb ^ p37_array_index_2050617_comb ^ p37_array_index_2050618_comb ^ p37_array_index_2050585_comb ^ p36_literal_2043923[p37_array_index_2050602_comb] ^ p37_array_index_2050587_comb ^ p36_literal_2043920[p37_array_index_2050604_comb] ^ p36_literal_2043918[p37_array_index_2050589_comb] ^ p36_literal_2043916[p37_array_index_2050590_comb] ^ p36_literal_2043914[p37_array_index_2050591_comb] ^ p36_literal_2043912[p37_array_index_2050592_comb] ^ p36_literal_2043910[p37_array_index_2050593_comb] ^ p37_array_index_2050594_comb;
  assign p37_array_index_2050628_comb = p36_literal_2043912[p37_res7__480_comb];
  assign p37_array_index_2050629_comb = p36_literal_2043914[p37_array_index_2050580_comb];
  assign p37_array_index_2050630_comb = p36_literal_2043916[p37_array_index_2050581_comb];
  assign p37_array_index_2050631_comb = p36_literal_2043918[p37_array_index_2050582_comb];
  assign p37_array_index_2050632_comb = p36_literal_2043920[p37_array_index_2050583_comb];
  assign p37_res7__484_comb = p36_literal_2043910[p37_res7__482_comb] ^ p37_array_index_2050628_comb ^ p37_array_index_2050629_comb ^ p37_array_index_2050630_comb ^ p37_array_index_2050631_comb ^ p37_array_index_2050632_comb ^ p37_array_index_2050584_comb ^ p36_literal_2043923[p37_array_index_2050585_comb] ^ p37_array_index_2050602_comb ^ p36_literal_2043920[p37_array_index_2050587_comb] ^ p36_literal_2043918[p37_array_index_2050604_comb] ^ p36_literal_2043916[p37_array_index_2050589_comb] ^ p36_literal_2043914[p37_array_index_2050590_comb] ^ p36_literal_2043912[p37_array_index_2050591_comb] ^ p36_literal_2043910[p37_array_index_2050592_comb] ^ p37_array_index_2050593_comb;

  // Registers for pipe stage 37:
  reg [127:0] p37_encoded;
  reg [127:0] p37_bit_slice_2043893;
  reg [127:0] p37_bit_slice_2044018;
  reg [127:0] p37_k3;
  reg [127:0] p37_k2;
  reg [127:0] p37_xor_2050132;
  reg [127:0] p37_k5;
  reg [7:0] p37_array_index_2050580;
  reg [7:0] p37_array_index_2050581;
  reg [7:0] p37_array_index_2050582;
  reg [7:0] p37_array_index_2050583;
  reg [7:0] p37_array_index_2050584;
  reg [7:0] p37_array_index_2050585;
  reg [7:0] p37_array_index_2050587;
  reg [7:0] p37_array_index_2050589;
  reg [7:0] p37_array_index_2050590;
  reg [7:0] p37_array_index_2050591;
  reg [7:0] p37_array_index_2050592;
  reg [7:0] p37_array_index_2050596;
  reg [7:0] p37_array_index_2050597;
  reg [7:0] p37_array_index_2050598;
  reg [7:0] p37_array_index_2050599;
  reg [7:0] p37_array_index_2050600;
  reg [7:0] p37_array_index_2050601;
  reg [7:0] p37_array_index_2050602;
  reg [7:0] p37_array_index_2050604;
  reg [7:0] p37_res7__480;
  reg [7:0] p37_array_index_2050613;
  reg [7:0] p37_array_index_2050614;
  reg [7:0] p37_array_index_2050615;
  reg [7:0] p37_array_index_2050616;
  reg [7:0] p37_array_index_2050617;
  reg [7:0] p37_array_index_2050618;
  reg [7:0] p37_res7__482;
  reg [7:0] p37_array_index_2050628;
  reg [7:0] p37_array_index_2050629;
  reg [7:0] p37_array_index_2050630;
  reg [7:0] p37_array_index_2050631;
  reg [7:0] p37_array_index_2050632;
  reg [7:0] p37_res7__484;
  reg [7:0] p38_literal_2043896[256];
  reg [7:0] p38_literal_2043910[256];
  reg [7:0] p38_literal_2043912[256];
  reg [7:0] p38_literal_2043914[256];
  reg [7:0] p38_literal_2043916[256];
  reg [7:0] p38_literal_2043918[256];
  reg [7:0] p38_literal_2043920[256];
  reg [7:0] p38_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p37_encoded <= p36_encoded;
    p37_bit_slice_2043893 <= p36_bit_slice_2043893;
    p37_bit_slice_2044018 <= p36_bit_slice_2044018;
    p37_k3 <= p36_k3;
    p37_k2 <= p36_k2;
    p37_xor_2050132 <= p36_xor_2050132;
    p37_k5 <= p37_k5_comb;
    p37_array_index_2050580 <= p37_array_index_2050580_comb;
    p37_array_index_2050581 <= p37_array_index_2050581_comb;
    p37_array_index_2050582 <= p37_array_index_2050582_comb;
    p37_array_index_2050583 <= p37_array_index_2050583_comb;
    p37_array_index_2050584 <= p37_array_index_2050584_comb;
    p37_array_index_2050585 <= p37_array_index_2050585_comb;
    p37_array_index_2050587 <= p37_array_index_2050587_comb;
    p37_array_index_2050589 <= p37_array_index_2050589_comb;
    p37_array_index_2050590 <= p37_array_index_2050590_comb;
    p37_array_index_2050591 <= p37_array_index_2050591_comb;
    p37_array_index_2050592 <= p37_array_index_2050592_comb;
    p37_array_index_2050596 <= p37_array_index_2050596_comb;
    p37_array_index_2050597 <= p37_array_index_2050597_comb;
    p37_array_index_2050598 <= p37_array_index_2050598_comb;
    p37_array_index_2050599 <= p37_array_index_2050599_comb;
    p37_array_index_2050600 <= p37_array_index_2050600_comb;
    p37_array_index_2050601 <= p37_array_index_2050601_comb;
    p37_array_index_2050602 <= p37_array_index_2050602_comb;
    p37_array_index_2050604 <= p37_array_index_2050604_comb;
    p37_res7__480 <= p37_res7__480_comb;
    p37_array_index_2050613 <= p37_array_index_2050613_comb;
    p37_array_index_2050614 <= p37_array_index_2050614_comb;
    p37_array_index_2050615 <= p37_array_index_2050615_comb;
    p37_array_index_2050616 <= p37_array_index_2050616_comb;
    p37_array_index_2050617 <= p37_array_index_2050617_comb;
    p37_array_index_2050618 <= p37_array_index_2050618_comb;
    p37_res7__482 <= p37_res7__482_comb;
    p37_array_index_2050628 <= p37_array_index_2050628_comb;
    p37_array_index_2050629 <= p37_array_index_2050629_comb;
    p37_array_index_2050630 <= p37_array_index_2050630_comb;
    p37_array_index_2050631 <= p37_array_index_2050631_comb;
    p37_array_index_2050632 <= p37_array_index_2050632_comb;
    p37_res7__484 <= p37_res7__484_comb;
    p38_literal_2043896 <= p37_literal_2043896;
    p38_literal_2043910 <= p37_literal_2043910;
    p38_literal_2043912 <= p37_literal_2043912;
    p38_literal_2043914 <= p37_literal_2043914;
    p38_literal_2043916 <= p37_literal_2043916;
    p38_literal_2043918 <= p37_literal_2043918;
    p38_literal_2043920 <= p37_literal_2043920;
    p38_literal_2043923 <= p37_literal_2043923;
  end

  // ===== Pipe stage 38:
  wire [7:0] p38_array_index_2050738_comb;
  wire [7:0] p38_array_index_2050739_comb;
  wire [7:0] p38_array_index_2050740_comb;
  wire [7:0] p38_array_index_2050741_comb;
  wire [7:0] p38_array_index_2050742_comb;
  wire [7:0] p38_res7__486_comb;
  wire [7:0] p38_array_index_2050753_comb;
  wire [7:0] p38_array_index_2050754_comb;
  wire [7:0] p38_array_index_2050755_comb;
  wire [7:0] p38_array_index_2050756_comb;
  wire [7:0] p38_res7__488_comb;
  wire [7:0] p38_array_index_2050766_comb;
  wire [7:0] p38_array_index_2050767_comb;
  wire [7:0] p38_array_index_2050768_comb;
  wire [7:0] p38_array_index_2050769_comb;
  wire [7:0] p38_res7__490_comb;
  wire [7:0] p38_array_index_2050780_comb;
  wire [7:0] p38_array_index_2050781_comb;
  wire [7:0] p38_array_index_2050782_comb;
  wire [7:0] p38_res7__492_comb;
  wire [7:0] p38_array_index_2050792_comb;
  wire [7:0] p38_array_index_2050793_comb;
  wire [7:0] p38_array_index_2050794_comb;
  wire [7:0] p38_res7__494_comb;
  wire [7:0] p38_array_index_2050805_comb;
  wire [7:0] p38_array_index_2050806_comb;
  wire [7:0] p38_res7__496_comb;
  wire [7:0] p38_array_index_2050816_comb;
  wire [7:0] p38_array_index_2050817_comb;
  wire [7:0] p38_res7__498_comb;
  assign p38_array_index_2050738_comb = p37_literal_2043912[p37_res7__482];
  assign p38_array_index_2050739_comb = p37_literal_2043914[p37_res7__480];
  assign p38_array_index_2050740_comb = p37_literal_2043916[p37_array_index_2050580];
  assign p38_array_index_2050741_comb = p37_literal_2043918[p37_array_index_2050581];
  assign p38_array_index_2050742_comb = p37_literal_2043920[p37_array_index_2050582];
  assign p38_res7__486_comb = p37_literal_2043910[p37_res7__484] ^ p38_array_index_2050738_comb ^ p38_array_index_2050739_comb ^ p38_array_index_2050740_comb ^ p38_array_index_2050741_comb ^ p38_array_index_2050742_comb ^ p37_array_index_2050583 ^ p37_literal_2043923[p37_array_index_2050584] ^ p37_array_index_2050585 ^ p37_literal_2043920[p37_array_index_2050602] ^ p37_literal_2043918[p37_array_index_2050587] ^ p37_literal_2043916[p37_array_index_2050604] ^ p37_literal_2043914[p37_array_index_2050589] ^ p37_literal_2043912[p37_array_index_2050590] ^ p37_literal_2043910[p37_array_index_2050591] ^ p37_array_index_2050592;
  assign p38_array_index_2050753_comb = p37_literal_2043914[p37_res7__482];
  assign p38_array_index_2050754_comb = p37_literal_2043916[p37_res7__480];
  assign p38_array_index_2050755_comb = p37_literal_2043918[p37_array_index_2050580];
  assign p38_array_index_2050756_comb = p37_literal_2043920[p37_array_index_2050581];
  assign p38_res7__488_comb = p37_literal_2043910[p38_res7__486_comb] ^ p37_literal_2043912[p37_res7__484] ^ p38_array_index_2050753_comb ^ p38_array_index_2050754_comb ^ p38_array_index_2050755_comb ^ p38_array_index_2050756_comb ^ p37_array_index_2050582 ^ p37_literal_2043923[p37_array_index_2050583] ^ p37_array_index_2050584 ^ p37_array_index_2050601 ^ p37_literal_2043918[p37_array_index_2050602] ^ p37_literal_2043916[p37_array_index_2050587] ^ p37_literal_2043914[p37_array_index_2050604] ^ p37_literal_2043912[p37_array_index_2050589] ^ p37_literal_2043910[p37_array_index_2050590] ^ p37_array_index_2050591;
  assign p38_array_index_2050766_comb = p37_literal_2043914[p37_res7__484];
  assign p38_array_index_2050767_comb = p37_literal_2043916[p37_res7__482];
  assign p38_array_index_2050768_comb = p37_literal_2043918[p37_res7__480];
  assign p38_array_index_2050769_comb = p37_literal_2043920[p37_array_index_2050580];
  assign p38_res7__490_comb = p37_literal_2043910[p38_res7__488_comb] ^ p37_literal_2043912[p38_res7__486_comb] ^ p38_array_index_2050766_comb ^ p38_array_index_2050767_comb ^ p38_array_index_2050768_comb ^ p38_array_index_2050769_comb ^ p37_array_index_2050581 ^ p37_literal_2043923[p37_array_index_2050582] ^ p37_array_index_2050583 ^ p37_array_index_2050618 ^ p37_literal_2043918[p37_array_index_2050585] ^ p37_literal_2043916[p37_array_index_2050602] ^ p37_literal_2043914[p37_array_index_2050587] ^ p37_literal_2043912[p37_array_index_2050604] ^ p37_literal_2043910[p37_array_index_2050589] ^ p37_array_index_2050590;
  assign p38_array_index_2050780_comb = p37_literal_2043916[p37_res7__484];
  assign p38_array_index_2050781_comb = p37_literal_2043918[p37_res7__482];
  assign p38_array_index_2050782_comb = p37_literal_2043920[p37_res7__480];
  assign p38_res7__492_comb = p37_literal_2043910[p38_res7__490_comb] ^ p37_literal_2043912[p38_res7__488_comb] ^ p37_literal_2043914[p38_res7__486_comb] ^ p38_array_index_2050780_comb ^ p38_array_index_2050781_comb ^ p38_array_index_2050782_comb ^ p37_array_index_2050580 ^ p37_literal_2043923[p37_array_index_2050581] ^ p37_array_index_2050582 ^ p37_array_index_2050632 ^ p37_array_index_2050600 ^ p37_literal_2043916[p37_array_index_2050585] ^ p37_literal_2043914[p37_array_index_2050602] ^ p37_literal_2043912[p37_array_index_2050587] ^ p37_literal_2043910[p37_array_index_2050604] ^ p37_array_index_2050589;
  assign p38_array_index_2050792_comb = p37_literal_2043916[p38_res7__486_comb];
  assign p38_array_index_2050793_comb = p37_literal_2043918[p37_res7__484];
  assign p38_array_index_2050794_comb = p37_literal_2043920[p37_res7__482];
  assign p38_res7__494_comb = p37_literal_2043910[p38_res7__492_comb] ^ p37_literal_2043912[p38_res7__490_comb] ^ p37_literal_2043914[p38_res7__488_comb] ^ p38_array_index_2050792_comb ^ p38_array_index_2050793_comb ^ p38_array_index_2050794_comb ^ p37_res7__480 ^ p37_literal_2043923[p37_array_index_2050580] ^ p37_array_index_2050581 ^ p38_array_index_2050742_comb ^ p37_array_index_2050617 ^ p37_literal_2043916[p37_array_index_2050584] ^ p37_literal_2043914[p37_array_index_2050585] ^ p37_literal_2043912[p37_array_index_2050602] ^ p37_literal_2043910[p37_array_index_2050587] ^ p37_array_index_2050604;
  assign p38_array_index_2050805_comb = p37_literal_2043918[p38_res7__486_comb];
  assign p38_array_index_2050806_comb = p37_literal_2043920[p37_res7__484];
  assign p38_res7__496_comb = p37_literal_2043910[p38_res7__494_comb] ^ p37_literal_2043912[p38_res7__492_comb] ^ p37_literal_2043914[p38_res7__490_comb] ^ p37_literal_2043916[p38_res7__488_comb] ^ p38_array_index_2050805_comb ^ p38_array_index_2050806_comb ^ p37_res7__482 ^ p37_literal_2043923[p37_res7__480] ^ p37_array_index_2050580 ^ p38_array_index_2050756_comb ^ p37_array_index_2050631 ^ p37_array_index_2050599 ^ p37_literal_2043914[p37_array_index_2050584] ^ p37_literal_2043912[p37_array_index_2050585] ^ p37_literal_2043910[p37_array_index_2050602] ^ p37_array_index_2050587;
  assign p38_array_index_2050816_comb = p37_literal_2043918[p38_res7__488_comb];
  assign p38_array_index_2050817_comb = p37_literal_2043920[p38_res7__486_comb];
  assign p38_res7__498_comb = p37_literal_2043910[p38_res7__496_comb] ^ p37_literal_2043912[p38_res7__494_comb] ^ p37_literal_2043914[p38_res7__492_comb] ^ p37_literal_2043916[p38_res7__490_comb] ^ p38_array_index_2050816_comb ^ p38_array_index_2050817_comb ^ p37_res7__484 ^ p37_literal_2043923[p37_res7__482] ^ p37_res7__480 ^ p38_array_index_2050769_comb ^ p38_array_index_2050741_comb ^ p37_array_index_2050616 ^ p37_literal_2043914[p37_array_index_2050583] ^ p37_literal_2043912[p37_array_index_2050584] ^ p37_literal_2043910[p37_array_index_2050585] ^ p37_array_index_2050602;

  // Registers for pipe stage 38:
  reg [127:0] p38_encoded;
  reg [127:0] p38_bit_slice_2043893;
  reg [127:0] p38_bit_slice_2044018;
  reg [127:0] p38_k3;
  reg [127:0] p38_k2;
  reg [127:0] p38_xor_2050132;
  reg [127:0] p38_k5;
  reg [7:0] p38_array_index_2050580;
  reg [7:0] p38_array_index_2050581;
  reg [7:0] p38_array_index_2050582;
  reg [7:0] p38_array_index_2050583;
  reg [7:0] p38_array_index_2050584;
  reg [7:0] p38_array_index_2050585;
  reg [7:0] p38_array_index_2050596;
  reg [7:0] p38_array_index_2050597;
  reg [7:0] p38_array_index_2050598;
  reg [7:0] p38_res7__480;
  reg [7:0] p38_array_index_2050613;
  reg [7:0] p38_array_index_2050614;
  reg [7:0] p38_array_index_2050615;
  reg [7:0] p38_res7__482;
  reg [7:0] p38_array_index_2050628;
  reg [7:0] p38_array_index_2050629;
  reg [7:0] p38_array_index_2050630;
  reg [7:0] p38_res7__484;
  reg [7:0] p38_array_index_2050738;
  reg [7:0] p38_array_index_2050739;
  reg [7:0] p38_array_index_2050740;
  reg [7:0] p38_res7__486;
  reg [7:0] p38_array_index_2050753;
  reg [7:0] p38_array_index_2050754;
  reg [7:0] p38_array_index_2050755;
  reg [7:0] p38_res7__488;
  reg [7:0] p38_array_index_2050766;
  reg [7:0] p38_array_index_2050767;
  reg [7:0] p38_array_index_2050768;
  reg [7:0] p38_res7__490;
  reg [7:0] p38_array_index_2050780;
  reg [7:0] p38_array_index_2050781;
  reg [7:0] p38_array_index_2050782;
  reg [7:0] p38_res7__492;
  reg [7:0] p38_array_index_2050792;
  reg [7:0] p38_array_index_2050793;
  reg [7:0] p38_array_index_2050794;
  reg [7:0] p38_res7__494;
  reg [7:0] p38_array_index_2050805;
  reg [7:0] p38_array_index_2050806;
  reg [7:0] p38_res7__496;
  reg [7:0] p38_array_index_2050816;
  reg [7:0] p38_array_index_2050817;
  reg [7:0] p38_res7__498;
  reg [7:0] p39_literal_2043896[256];
  reg [7:0] p39_literal_2043910[256];
  reg [7:0] p39_literal_2043912[256];
  reg [7:0] p39_literal_2043914[256];
  reg [7:0] p39_literal_2043916[256];
  reg [7:0] p39_literal_2043918[256];
  reg [7:0] p39_literal_2043920[256];
  reg [7:0] p39_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p38_encoded <= p37_encoded;
    p38_bit_slice_2043893 <= p37_bit_slice_2043893;
    p38_bit_slice_2044018 <= p37_bit_slice_2044018;
    p38_k3 <= p37_k3;
    p38_k2 <= p37_k2;
    p38_xor_2050132 <= p37_xor_2050132;
    p38_k5 <= p37_k5;
    p38_array_index_2050580 <= p37_array_index_2050580;
    p38_array_index_2050581 <= p37_array_index_2050581;
    p38_array_index_2050582 <= p37_array_index_2050582;
    p38_array_index_2050583 <= p37_array_index_2050583;
    p38_array_index_2050584 <= p37_array_index_2050584;
    p38_array_index_2050585 <= p37_array_index_2050585;
    p38_array_index_2050596 <= p37_array_index_2050596;
    p38_array_index_2050597 <= p37_array_index_2050597;
    p38_array_index_2050598 <= p37_array_index_2050598;
    p38_res7__480 <= p37_res7__480;
    p38_array_index_2050613 <= p37_array_index_2050613;
    p38_array_index_2050614 <= p37_array_index_2050614;
    p38_array_index_2050615 <= p37_array_index_2050615;
    p38_res7__482 <= p37_res7__482;
    p38_array_index_2050628 <= p37_array_index_2050628;
    p38_array_index_2050629 <= p37_array_index_2050629;
    p38_array_index_2050630 <= p37_array_index_2050630;
    p38_res7__484 <= p37_res7__484;
    p38_array_index_2050738 <= p38_array_index_2050738_comb;
    p38_array_index_2050739 <= p38_array_index_2050739_comb;
    p38_array_index_2050740 <= p38_array_index_2050740_comb;
    p38_res7__486 <= p38_res7__486_comb;
    p38_array_index_2050753 <= p38_array_index_2050753_comb;
    p38_array_index_2050754 <= p38_array_index_2050754_comb;
    p38_array_index_2050755 <= p38_array_index_2050755_comb;
    p38_res7__488 <= p38_res7__488_comb;
    p38_array_index_2050766 <= p38_array_index_2050766_comb;
    p38_array_index_2050767 <= p38_array_index_2050767_comb;
    p38_array_index_2050768 <= p38_array_index_2050768_comb;
    p38_res7__490 <= p38_res7__490_comb;
    p38_array_index_2050780 <= p38_array_index_2050780_comb;
    p38_array_index_2050781 <= p38_array_index_2050781_comb;
    p38_array_index_2050782 <= p38_array_index_2050782_comb;
    p38_res7__492 <= p38_res7__492_comb;
    p38_array_index_2050792 <= p38_array_index_2050792_comb;
    p38_array_index_2050793 <= p38_array_index_2050793_comb;
    p38_array_index_2050794 <= p38_array_index_2050794_comb;
    p38_res7__494 <= p38_res7__494_comb;
    p38_array_index_2050805 <= p38_array_index_2050805_comb;
    p38_array_index_2050806 <= p38_array_index_2050806_comb;
    p38_res7__496 <= p38_res7__496_comb;
    p38_array_index_2050816 <= p38_array_index_2050816_comb;
    p38_array_index_2050817 <= p38_array_index_2050817_comb;
    p38_res7__498 <= p38_res7__498_comb;
    p39_literal_2043896 <= p38_literal_2043896;
    p39_literal_2043910 <= p38_literal_2043910;
    p39_literal_2043912 <= p38_literal_2043912;
    p39_literal_2043914 <= p38_literal_2043914;
    p39_literal_2043916 <= p38_literal_2043916;
    p39_literal_2043918 <= p38_literal_2043918;
    p39_literal_2043920 <= p38_literal_2043920;
    p39_literal_2043923 <= p38_literal_2043923;
  end

  // ===== Pipe stage 39:
  wire [7:0] p39_array_index_2050946_comb;
  wire [7:0] p39_res7__500_comb;
  wire [7:0] p39_array_index_2050956_comb;
  wire [7:0] p39_res7__502_comb;
  wire [7:0] p39_res7__504_comb;
  wire [7:0] p39_res7__506_comb;
  wire [7:0] p39_res7__508_comb;
  wire [7:0] p39_res7__510_comb;
  wire [127:0] p39_res__15_comb;
  wire [127:0] p39_k4_comb;
  wire [127:0] p39_addedKey__48_comb;
  wire [7:0] p39_array_index_2051012_comb;
  wire [7:0] p39_array_index_2051013_comb;
  wire [7:0] p39_array_index_2051014_comb;
  wire [7:0] p39_array_index_2051015_comb;
  wire [7:0] p39_array_index_2051016_comb;
  wire [7:0] p39_array_index_2051017_comb;
  wire [7:0] p39_array_index_2051019_comb;
  wire [7:0] p39_array_index_2051021_comb;
  wire [7:0] p39_array_index_2051022_comb;
  wire [7:0] p39_array_index_2051023_comb;
  wire [7:0] p39_array_index_2051024_comb;
  wire [7:0] p39_array_index_2051025_comb;
  wire [7:0] p39_array_index_2051026_comb;
  wire [7:0] p39_array_index_2051028_comb;
  wire [7:0] p39_array_index_2051029_comb;
  wire [7:0] p39_array_index_2051030_comb;
  assign p39_array_index_2050946_comb = p38_literal_2043920[p38_res7__488];
  assign p39_res7__500_comb = p38_literal_2043910[p38_res7__498] ^ p38_literal_2043912[p38_res7__496] ^ p38_literal_2043914[p38_res7__494] ^ p38_literal_2043916[p38_res7__492] ^ p38_literal_2043918[p38_res7__490] ^ p39_array_index_2050946_comb ^ p38_res7__486 ^ p38_literal_2043923[p38_res7__484] ^ p38_res7__482 ^ p38_array_index_2050782 ^ p38_array_index_2050755 ^ p38_array_index_2050630 ^ p38_array_index_2050598 ^ p38_literal_2043912[p38_array_index_2050583] ^ p38_literal_2043910[p38_array_index_2050584] ^ p38_array_index_2050585;
  assign p39_array_index_2050956_comb = p38_literal_2043920[p38_res7__490];
  assign p39_res7__502_comb = p38_literal_2043910[p39_res7__500_comb] ^ p38_literal_2043912[p38_res7__498] ^ p38_literal_2043914[p38_res7__496] ^ p38_literal_2043916[p38_res7__494] ^ p38_literal_2043918[p38_res7__492] ^ p39_array_index_2050956_comb ^ p38_res7__488 ^ p38_literal_2043923[p38_res7__486] ^ p38_res7__484 ^ p38_array_index_2050794 ^ p38_array_index_2050768 ^ p38_array_index_2050740 ^ p38_array_index_2050615 ^ p38_literal_2043912[p38_array_index_2050582] ^ p38_literal_2043910[p38_array_index_2050583] ^ p38_array_index_2050584;
  assign p39_res7__504_comb = p38_literal_2043910[p39_res7__502_comb] ^ p38_literal_2043912[p39_res7__500_comb] ^ p38_literal_2043914[p38_res7__498] ^ p38_literal_2043916[p38_res7__496] ^ p38_literal_2043918[p38_res7__494] ^ p38_literal_2043920[p38_res7__492] ^ p38_res7__490 ^ p38_literal_2043923[p38_res7__488] ^ p38_res7__486 ^ p38_array_index_2050806 ^ p38_array_index_2050781 ^ p38_array_index_2050754 ^ p38_array_index_2050629 ^ p38_array_index_2050597 ^ p38_literal_2043910[p38_array_index_2050582] ^ p38_array_index_2050583;
  assign p39_res7__506_comb = p38_literal_2043910[p39_res7__504_comb] ^ p38_literal_2043912[p39_res7__502_comb] ^ p38_literal_2043914[p39_res7__500_comb] ^ p38_literal_2043916[p38_res7__498] ^ p38_literal_2043918[p38_res7__496] ^ p38_literal_2043920[p38_res7__494] ^ p38_res7__492 ^ p38_literal_2043923[p38_res7__490] ^ p38_res7__488 ^ p38_array_index_2050817 ^ p38_array_index_2050793 ^ p38_array_index_2050767 ^ p38_array_index_2050739 ^ p38_array_index_2050614 ^ p38_literal_2043910[p38_array_index_2050581] ^ p38_array_index_2050582;
  assign p39_res7__508_comb = p38_literal_2043910[p39_res7__506_comb] ^ p38_literal_2043912[p39_res7__504_comb] ^ p38_literal_2043914[p39_res7__502_comb] ^ p38_literal_2043916[p39_res7__500_comb] ^ p38_literal_2043918[p38_res7__498] ^ p38_literal_2043920[p38_res7__496] ^ p38_res7__494 ^ p38_literal_2043923[p38_res7__492] ^ p38_res7__490 ^ p39_array_index_2050946_comb ^ p38_array_index_2050805 ^ p38_array_index_2050780 ^ p38_array_index_2050753 ^ p38_array_index_2050628 ^ p38_array_index_2050596 ^ p38_array_index_2050581;
  assign p39_res7__510_comb = p38_literal_2043910[p39_res7__508_comb] ^ p38_literal_2043912[p39_res7__506_comb] ^ p38_literal_2043914[p39_res7__504_comb] ^ p38_literal_2043916[p39_res7__502_comb] ^ p38_literal_2043918[p39_res7__500_comb] ^ p38_literal_2043920[p38_res7__498] ^ p38_res7__496 ^ p38_literal_2043923[p38_res7__494] ^ p38_res7__492 ^ p39_array_index_2050956_comb ^ p38_array_index_2050816 ^ p38_array_index_2050792 ^ p38_array_index_2050766 ^ p38_array_index_2050738 ^ p38_array_index_2050613 ^ p38_array_index_2050580;
  assign p39_res__15_comb = {p39_res7__510_comb, p39_res7__508_comb, p39_res7__506_comb, p39_res7__504_comb, p39_res7__502_comb, p39_res7__500_comb, p38_res7__498, p38_res7__496, p38_res7__494, p38_res7__492, p38_res7__490, p38_res7__488, p38_res7__486, p38_res7__484, p38_res7__482, p38_res7__480};
  assign p39_k4_comb = p39_res__15_comb ^ p38_xor_2050132;
  assign p39_addedKey__48_comb = p39_k4_comb ^ 128'h4110_1a5e_6342_d669_c412_3cd3_9313_c011;
  assign p39_array_index_2051012_comb = p38_literal_2043896[p39_addedKey__48_comb[127:120]];
  assign p39_array_index_2051013_comb = p38_literal_2043896[p39_addedKey__48_comb[119:112]];
  assign p39_array_index_2051014_comb = p38_literal_2043896[p39_addedKey__48_comb[111:104]];
  assign p39_array_index_2051015_comb = p38_literal_2043896[p39_addedKey__48_comb[103:96]];
  assign p39_array_index_2051016_comb = p38_literal_2043896[p39_addedKey__48_comb[95:88]];
  assign p39_array_index_2051017_comb = p38_literal_2043896[p39_addedKey__48_comb[87:80]];
  assign p39_array_index_2051019_comb = p38_literal_2043896[p39_addedKey__48_comb[71:64]];
  assign p39_array_index_2051021_comb = p38_literal_2043896[p39_addedKey__48_comb[55:48]];
  assign p39_array_index_2051022_comb = p38_literal_2043896[p39_addedKey__48_comb[47:40]];
  assign p39_array_index_2051023_comb = p38_literal_2043896[p39_addedKey__48_comb[39:32]];
  assign p39_array_index_2051024_comb = p38_literal_2043896[p39_addedKey__48_comb[31:24]];
  assign p39_array_index_2051025_comb = p38_literal_2043896[p39_addedKey__48_comb[23:16]];
  assign p39_array_index_2051026_comb = p38_literal_2043896[p39_addedKey__48_comb[15:8]];
  assign p39_array_index_2051028_comb = p38_literal_2043896[p39_addedKey__48_comb[79:72]];
  assign p39_array_index_2051029_comb = p38_literal_2043896[p39_addedKey__48_comb[63:56]];
  assign p39_array_index_2051030_comb = p38_literal_2043896[p39_addedKey__48_comb[7:0]];

  // Registers for pipe stage 39:
  reg [127:0] p39_encoded;
  reg [127:0] p39_bit_slice_2043893;
  reg [127:0] p39_bit_slice_2044018;
  reg [127:0] p39_k3;
  reg [127:0] p39_k2;
  reg [127:0] p39_k5;
  reg [127:0] p39_k4;
  reg [7:0] p39_array_index_2051012;
  reg [7:0] p39_array_index_2051013;
  reg [7:0] p39_array_index_2051014;
  reg [7:0] p39_array_index_2051015;
  reg [7:0] p39_array_index_2051016;
  reg [7:0] p39_array_index_2051017;
  reg [7:0] p39_array_index_2051019;
  reg [7:0] p39_array_index_2051021;
  reg [7:0] p39_array_index_2051022;
  reg [7:0] p39_array_index_2051023;
  reg [7:0] p39_array_index_2051024;
  reg [7:0] p39_array_index_2051025;
  reg [7:0] p39_array_index_2051026;
  reg [7:0] p39_array_index_2051028;
  reg [7:0] p39_array_index_2051029;
  reg [7:0] p39_array_index_2051030;
  reg [7:0] p40_literal_2043896[256];
  reg [7:0] p40_literal_2043910[256];
  reg [7:0] p40_literal_2043912[256];
  reg [7:0] p40_literal_2043914[256];
  reg [7:0] p40_literal_2043916[256];
  reg [7:0] p40_literal_2043918[256];
  reg [7:0] p40_literal_2043920[256];
  reg [7:0] p40_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p39_encoded <= p38_encoded;
    p39_bit_slice_2043893 <= p38_bit_slice_2043893;
    p39_bit_slice_2044018 <= p38_bit_slice_2044018;
    p39_k3 <= p38_k3;
    p39_k2 <= p38_k2;
    p39_k5 <= p38_k5;
    p39_k4 <= p39_k4_comb;
    p39_array_index_2051012 <= p39_array_index_2051012_comb;
    p39_array_index_2051013 <= p39_array_index_2051013_comb;
    p39_array_index_2051014 <= p39_array_index_2051014_comb;
    p39_array_index_2051015 <= p39_array_index_2051015_comb;
    p39_array_index_2051016 <= p39_array_index_2051016_comb;
    p39_array_index_2051017 <= p39_array_index_2051017_comb;
    p39_array_index_2051019 <= p39_array_index_2051019_comb;
    p39_array_index_2051021 <= p39_array_index_2051021_comb;
    p39_array_index_2051022 <= p39_array_index_2051022_comb;
    p39_array_index_2051023 <= p39_array_index_2051023_comb;
    p39_array_index_2051024 <= p39_array_index_2051024_comb;
    p39_array_index_2051025 <= p39_array_index_2051025_comb;
    p39_array_index_2051026 <= p39_array_index_2051026_comb;
    p39_array_index_2051028 <= p39_array_index_2051028_comb;
    p39_array_index_2051029 <= p39_array_index_2051029_comb;
    p39_array_index_2051030 <= p39_array_index_2051030_comb;
    p40_literal_2043896 <= p39_literal_2043896;
    p40_literal_2043910 <= p39_literal_2043910;
    p40_literal_2043912 <= p39_literal_2043912;
    p40_literal_2043914 <= p39_literal_2043914;
    p40_literal_2043916 <= p39_literal_2043916;
    p40_literal_2043918 <= p39_literal_2043918;
    p40_literal_2043920 <= p39_literal_2043920;
    p40_literal_2043923 <= p39_literal_2043923;
  end

  // ===== Pipe stage 40:
  wire [7:0] p40_array_index_2051093_comb;
  wire [7:0] p40_array_index_2051094_comb;
  wire [7:0] p40_array_index_2051095_comb;
  wire [7:0] p40_array_index_2051096_comb;
  wire [7:0] p40_array_index_2051097_comb;
  wire [7:0] p40_array_index_2051098_comb;
  wire [7:0] p40_res7__512_comb;
  wire [7:0] p40_array_index_2051107_comb;
  wire [7:0] p40_array_index_2051108_comb;
  wire [7:0] p40_array_index_2051109_comb;
  wire [7:0] p40_array_index_2051110_comb;
  wire [7:0] p40_array_index_2051111_comb;
  wire [7:0] p40_array_index_2051112_comb;
  wire [7:0] p40_res7__514_comb;
  wire [7:0] p40_array_index_2051122_comb;
  wire [7:0] p40_array_index_2051123_comb;
  wire [7:0] p40_array_index_2051124_comb;
  wire [7:0] p40_array_index_2051125_comb;
  wire [7:0] p40_array_index_2051126_comb;
  wire [7:0] p40_res7__516_comb;
  wire [7:0] p40_array_index_2051136_comb;
  wire [7:0] p40_array_index_2051137_comb;
  wire [7:0] p40_array_index_2051138_comb;
  wire [7:0] p40_array_index_2051139_comb;
  wire [7:0] p40_array_index_2051140_comb;
  wire [7:0] p40_res7__518_comb;
  wire [7:0] p40_array_index_2051151_comb;
  wire [7:0] p40_array_index_2051152_comb;
  wire [7:0] p40_array_index_2051153_comb;
  wire [7:0] p40_array_index_2051154_comb;
  wire [7:0] p40_res7__520_comb;
  wire [7:0] p40_array_index_2051164_comb;
  wire [7:0] p40_array_index_2051165_comb;
  wire [7:0] p40_array_index_2051166_comb;
  wire [7:0] p40_array_index_2051167_comb;
  wire [7:0] p40_res7__522_comb;
  wire [7:0] p40_array_index_2051178_comb;
  wire [7:0] p40_array_index_2051179_comb;
  wire [7:0] p40_array_index_2051180_comb;
  wire [7:0] p40_res7__524_comb;
  assign p40_array_index_2051093_comb = p39_literal_2043910[p39_array_index_2051012];
  assign p40_array_index_2051094_comb = p39_literal_2043912[p39_array_index_2051013];
  assign p40_array_index_2051095_comb = p39_literal_2043914[p39_array_index_2051014];
  assign p40_array_index_2051096_comb = p39_literal_2043916[p39_array_index_2051015];
  assign p40_array_index_2051097_comb = p39_literal_2043918[p39_array_index_2051016];
  assign p40_array_index_2051098_comb = p39_literal_2043920[p39_array_index_2051017];
  assign p40_res7__512_comb = p40_array_index_2051093_comb ^ p40_array_index_2051094_comb ^ p40_array_index_2051095_comb ^ p40_array_index_2051096_comb ^ p40_array_index_2051097_comb ^ p40_array_index_2051098_comb ^ p39_array_index_2051028 ^ p39_literal_2043923[p39_array_index_2051019] ^ p39_array_index_2051029 ^ p39_literal_2043920[p39_array_index_2051021] ^ p39_literal_2043918[p39_array_index_2051022] ^ p39_literal_2043916[p39_array_index_2051023] ^ p39_literal_2043914[p39_array_index_2051024] ^ p39_literal_2043912[p39_array_index_2051025] ^ p39_literal_2043910[p39_array_index_2051026] ^ p39_array_index_2051030;
  assign p40_array_index_2051107_comb = p39_literal_2043910[p40_res7__512_comb];
  assign p40_array_index_2051108_comb = p39_literal_2043912[p39_array_index_2051012];
  assign p40_array_index_2051109_comb = p39_literal_2043914[p39_array_index_2051013];
  assign p40_array_index_2051110_comb = p39_literal_2043916[p39_array_index_2051014];
  assign p40_array_index_2051111_comb = p39_literal_2043918[p39_array_index_2051015];
  assign p40_array_index_2051112_comb = p39_literal_2043920[p39_array_index_2051016];
  assign p40_res7__514_comb = p40_array_index_2051107_comb ^ p40_array_index_2051108_comb ^ p40_array_index_2051109_comb ^ p40_array_index_2051110_comb ^ p40_array_index_2051111_comb ^ p40_array_index_2051112_comb ^ p39_array_index_2051017 ^ p39_literal_2043923[p39_array_index_2051028] ^ p39_array_index_2051019 ^ p39_literal_2043920[p39_array_index_2051029] ^ p39_literal_2043918[p39_array_index_2051021] ^ p39_literal_2043916[p39_array_index_2051022] ^ p39_literal_2043914[p39_array_index_2051023] ^ p39_literal_2043912[p39_array_index_2051024] ^ p39_literal_2043910[p39_array_index_2051025] ^ p39_array_index_2051026;
  assign p40_array_index_2051122_comb = p39_literal_2043912[p40_res7__512_comb];
  assign p40_array_index_2051123_comb = p39_literal_2043914[p39_array_index_2051012];
  assign p40_array_index_2051124_comb = p39_literal_2043916[p39_array_index_2051013];
  assign p40_array_index_2051125_comb = p39_literal_2043918[p39_array_index_2051014];
  assign p40_array_index_2051126_comb = p39_literal_2043920[p39_array_index_2051015];
  assign p40_res7__516_comb = p39_literal_2043910[p40_res7__514_comb] ^ p40_array_index_2051122_comb ^ p40_array_index_2051123_comb ^ p40_array_index_2051124_comb ^ p40_array_index_2051125_comb ^ p40_array_index_2051126_comb ^ p39_array_index_2051016 ^ p39_literal_2043923[p39_array_index_2051017] ^ p39_array_index_2051028 ^ p39_literal_2043920[p39_array_index_2051019] ^ p39_literal_2043918[p39_array_index_2051029] ^ p39_literal_2043916[p39_array_index_2051021] ^ p39_literal_2043914[p39_array_index_2051022] ^ p39_literal_2043912[p39_array_index_2051023] ^ p39_literal_2043910[p39_array_index_2051024] ^ p39_array_index_2051025;
  assign p40_array_index_2051136_comb = p39_literal_2043912[p40_res7__514_comb];
  assign p40_array_index_2051137_comb = p39_literal_2043914[p40_res7__512_comb];
  assign p40_array_index_2051138_comb = p39_literal_2043916[p39_array_index_2051012];
  assign p40_array_index_2051139_comb = p39_literal_2043918[p39_array_index_2051013];
  assign p40_array_index_2051140_comb = p39_literal_2043920[p39_array_index_2051014];
  assign p40_res7__518_comb = p39_literal_2043910[p40_res7__516_comb] ^ p40_array_index_2051136_comb ^ p40_array_index_2051137_comb ^ p40_array_index_2051138_comb ^ p40_array_index_2051139_comb ^ p40_array_index_2051140_comb ^ p39_array_index_2051015 ^ p39_literal_2043923[p39_array_index_2051016] ^ p39_array_index_2051017 ^ p39_literal_2043920[p39_array_index_2051028] ^ p39_literal_2043918[p39_array_index_2051019] ^ p39_literal_2043916[p39_array_index_2051029] ^ p39_literal_2043914[p39_array_index_2051021] ^ p39_literal_2043912[p39_array_index_2051022] ^ p39_literal_2043910[p39_array_index_2051023] ^ p39_array_index_2051024;
  assign p40_array_index_2051151_comb = p39_literal_2043914[p40_res7__514_comb];
  assign p40_array_index_2051152_comb = p39_literal_2043916[p40_res7__512_comb];
  assign p40_array_index_2051153_comb = p39_literal_2043918[p39_array_index_2051012];
  assign p40_array_index_2051154_comb = p39_literal_2043920[p39_array_index_2051013];
  assign p40_res7__520_comb = p39_literal_2043910[p40_res7__518_comb] ^ p39_literal_2043912[p40_res7__516_comb] ^ p40_array_index_2051151_comb ^ p40_array_index_2051152_comb ^ p40_array_index_2051153_comb ^ p40_array_index_2051154_comb ^ p39_array_index_2051014 ^ p39_literal_2043923[p39_array_index_2051015] ^ p39_array_index_2051016 ^ p40_array_index_2051098_comb ^ p39_literal_2043918[p39_array_index_2051028] ^ p39_literal_2043916[p39_array_index_2051019] ^ p39_literal_2043914[p39_array_index_2051029] ^ p39_literal_2043912[p39_array_index_2051021] ^ p39_literal_2043910[p39_array_index_2051022] ^ p39_array_index_2051023;
  assign p40_array_index_2051164_comb = p39_literal_2043914[p40_res7__516_comb];
  assign p40_array_index_2051165_comb = p39_literal_2043916[p40_res7__514_comb];
  assign p40_array_index_2051166_comb = p39_literal_2043918[p40_res7__512_comb];
  assign p40_array_index_2051167_comb = p39_literal_2043920[p39_array_index_2051012];
  assign p40_res7__522_comb = p39_literal_2043910[p40_res7__520_comb] ^ p39_literal_2043912[p40_res7__518_comb] ^ p40_array_index_2051164_comb ^ p40_array_index_2051165_comb ^ p40_array_index_2051166_comb ^ p40_array_index_2051167_comb ^ p39_array_index_2051013 ^ p39_literal_2043923[p39_array_index_2051014] ^ p39_array_index_2051015 ^ p40_array_index_2051112_comb ^ p39_literal_2043918[p39_array_index_2051017] ^ p39_literal_2043916[p39_array_index_2051028] ^ p39_literal_2043914[p39_array_index_2051019] ^ p39_literal_2043912[p39_array_index_2051029] ^ p39_literal_2043910[p39_array_index_2051021] ^ p39_array_index_2051022;
  assign p40_array_index_2051178_comb = p39_literal_2043916[p40_res7__516_comb];
  assign p40_array_index_2051179_comb = p39_literal_2043918[p40_res7__514_comb];
  assign p40_array_index_2051180_comb = p39_literal_2043920[p40_res7__512_comb];
  assign p40_res7__524_comb = p39_literal_2043910[p40_res7__522_comb] ^ p39_literal_2043912[p40_res7__520_comb] ^ p39_literal_2043914[p40_res7__518_comb] ^ p40_array_index_2051178_comb ^ p40_array_index_2051179_comb ^ p40_array_index_2051180_comb ^ p39_array_index_2051012 ^ p39_literal_2043923[p39_array_index_2051013] ^ p39_array_index_2051014 ^ p40_array_index_2051126_comb ^ p40_array_index_2051097_comb ^ p39_literal_2043916[p39_array_index_2051017] ^ p39_literal_2043914[p39_array_index_2051028] ^ p39_literal_2043912[p39_array_index_2051019] ^ p39_literal_2043910[p39_array_index_2051029] ^ p39_array_index_2051021;

  // Registers for pipe stage 40:
  reg [127:0] p40_encoded;
  reg [127:0] p40_bit_slice_2043893;
  reg [127:0] p40_bit_slice_2044018;
  reg [127:0] p40_k3;
  reg [127:0] p40_k2;
  reg [127:0] p40_k5;
  reg [127:0] p40_k4;
  reg [7:0] p40_array_index_2051012;
  reg [7:0] p40_array_index_2051013;
  reg [7:0] p40_array_index_2051014;
  reg [7:0] p40_array_index_2051015;
  reg [7:0] p40_array_index_2051016;
  reg [7:0] p40_array_index_2051017;
  reg [7:0] p40_array_index_2051019;
  reg [7:0] p40_array_index_2051093;
  reg [7:0] p40_array_index_2051094;
  reg [7:0] p40_array_index_2051095;
  reg [7:0] p40_array_index_2051096;
  reg [7:0] p40_array_index_2051028;
  reg [7:0] p40_array_index_2051029;
  reg [7:0] p40_res7__512;
  reg [7:0] p40_array_index_2051107;
  reg [7:0] p40_array_index_2051108;
  reg [7:0] p40_array_index_2051109;
  reg [7:0] p40_array_index_2051110;
  reg [7:0] p40_array_index_2051111;
  reg [7:0] p40_res7__514;
  reg [7:0] p40_array_index_2051122;
  reg [7:0] p40_array_index_2051123;
  reg [7:0] p40_array_index_2051124;
  reg [7:0] p40_array_index_2051125;
  reg [7:0] p40_res7__516;
  reg [7:0] p40_array_index_2051136;
  reg [7:0] p40_array_index_2051137;
  reg [7:0] p40_array_index_2051138;
  reg [7:0] p40_array_index_2051139;
  reg [7:0] p40_array_index_2051140;
  reg [7:0] p40_res7__518;
  reg [7:0] p40_array_index_2051151;
  reg [7:0] p40_array_index_2051152;
  reg [7:0] p40_array_index_2051153;
  reg [7:0] p40_array_index_2051154;
  reg [7:0] p40_res7__520;
  reg [7:0] p40_array_index_2051164;
  reg [7:0] p40_array_index_2051165;
  reg [7:0] p40_array_index_2051166;
  reg [7:0] p40_array_index_2051167;
  reg [7:0] p40_res7__522;
  reg [7:0] p40_array_index_2051178;
  reg [7:0] p40_array_index_2051179;
  reg [7:0] p40_array_index_2051180;
  reg [7:0] p40_res7__524;
  reg [7:0] p41_literal_2043896[256];
  reg [7:0] p41_literal_2043910[256];
  reg [7:0] p41_literal_2043912[256];
  reg [7:0] p41_literal_2043914[256];
  reg [7:0] p41_literal_2043916[256];
  reg [7:0] p41_literal_2043918[256];
  reg [7:0] p41_literal_2043920[256];
  reg [7:0] p41_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p40_encoded <= p39_encoded;
    p40_bit_slice_2043893 <= p39_bit_slice_2043893;
    p40_bit_slice_2044018 <= p39_bit_slice_2044018;
    p40_k3 <= p39_k3;
    p40_k2 <= p39_k2;
    p40_k5 <= p39_k5;
    p40_k4 <= p39_k4;
    p40_array_index_2051012 <= p39_array_index_2051012;
    p40_array_index_2051013 <= p39_array_index_2051013;
    p40_array_index_2051014 <= p39_array_index_2051014;
    p40_array_index_2051015 <= p39_array_index_2051015;
    p40_array_index_2051016 <= p39_array_index_2051016;
    p40_array_index_2051017 <= p39_array_index_2051017;
    p40_array_index_2051019 <= p39_array_index_2051019;
    p40_array_index_2051093 <= p40_array_index_2051093_comb;
    p40_array_index_2051094 <= p40_array_index_2051094_comb;
    p40_array_index_2051095 <= p40_array_index_2051095_comb;
    p40_array_index_2051096 <= p40_array_index_2051096_comb;
    p40_array_index_2051028 <= p39_array_index_2051028;
    p40_array_index_2051029 <= p39_array_index_2051029;
    p40_res7__512 <= p40_res7__512_comb;
    p40_array_index_2051107 <= p40_array_index_2051107_comb;
    p40_array_index_2051108 <= p40_array_index_2051108_comb;
    p40_array_index_2051109 <= p40_array_index_2051109_comb;
    p40_array_index_2051110 <= p40_array_index_2051110_comb;
    p40_array_index_2051111 <= p40_array_index_2051111_comb;
    p40_res7__514 <= p40_res7__514_comb;
    p40_array_index_2051122 <= p40_array_index_2051122_comb;
    p40_array_index_2051123 <= p40_array_index_2051123_comb;
    p40_array_index_2051124 <= p40_array_index_2051124_comb;
    p40_array_index_2051125 <= p40_array_index_2051125_comb;
    p40_res7__516 <= p40_res7__516_comb;
    p40_array_index_2051136 <= p40_array_index_2051136_comb;
    p40_array_index_2051137 <= p40_array_index_2051137_comb;
    p40_array_index_2051138 <= p40_array_index_2051138_comb;
    p40_array_index_2051139 <= p40_array_index_2051139_comb;
    p40_array_index_2051140 <= p40_array_index_2051140_comb;
    p40_res7__518 <= p40_res7__518_comb;
    p40_array_index_2051151 <= p40_array_index_2051151_comb;
    p40_array_index_2051152 <= p40_array_index_2051152_comb;
    p40_array_index_2051153 <= p40_array_index_2051153_comb;
    p40_array_index_2051154 <= p40_array_index_2051154_comb;
    p40_res7__520 <= p40_res7__520_comb;
    p40_array_index_2051164 <= p40_array_index_2051164_comb;
    p40_array_index_2051165 <= p40_array_index_2051165_comb;
    p40_array_index_2051166 <= p40_array_index_2051166_comb;
    p40_array_index_2051167 <= p40_array_index_2051167_comb;
    p40_res7__522 <= p40_res7__522_comb;
    p40_array_index_2051178 <= p40_array_index_2051178_comb;
    p40_array_index_2051179 <= p40_array_index_2051179_comb;
    p40_array_index_2051180 <= p40_array_index_2051180_comb;
    p40_res7__524 <= p40_res7__524_comb;
    p41_literal_2043896 <= p40_literal_2043896;
    p41_literal_2043910 <= p40_literal_2043910;
    p41_literal_2043912 <= p40_literal_2043912;
    p41_literal_2043914 <= p40_literal_2043914;
    p41_literal_2043916 <= p40_literal_2043916;
    p41_literal_2043918 <= p40_literal_2043918;
    p41_literal_2043920 <= p40_literal_2043920;
    p41_literal_2043923 <= p40_literal_2043923;
  end

  // ===== Pipe stage 41:
  wire [7:0] p41_array_index_2051310_comb;
  wire [7:0] p41_array_index_2051311_comb;
  wire [7:0] p41_array_index_2051312_comb;
  wire [7:0] p41_res7__526_comb;
  wire [7:0] p41_array_index_2051323_comb;
  wire [7:0] p41_array_index_2051324_comb;
  wire [7:0] p41_res7__528_comb;
  wire [7:0] p41_array_index_2051334_comb;
  wire [7:0] p41_array_index_2051335_comb;
  wire [7:0] p41_res7__530_comb;
  wire [7:0] p41_array_index_2051346_comb;
  wire [7:0] p41_res7__532_comb;
  wire [7:0] p41_array_index_2051356_comb;
  wire [7:0] p41_res7__534_comb;
  wire [7:0] p41_res7__536_comb;
  wire [7:0] p41_res7__538_comb;
  assign p41_array_index_2051310_comb = p40_literal_2043916[p40_res7__518];
  assign p41_array_index_2051311_comb = p40_literal_2043918[p40_res7__516];
  assign p41_array_index_2051312_comb = p40_literal_2043920[p40_res7__514];
  assign p41_res7__526_comb = p40_literal_2043910[p40_res7__524] ^ p40_literal_2043912[p40_res7__522] ^ p40_literal_2043914[p40_res7__520] ^ p41_array_index_2051310_comb ^ p41_array_index_2051311_comb ^ p41_array_index_2051312_comb ^ p40_res7__512 ^ p40_literal_2043923[p40_array_index_2051012] ^ p40_array_index_2051013 ^ p40_array_index_2051140 ^ p40_array_index_2051111 ^ p40_literal_2043916[p40_array_index_2051016] ^ p40_literal_2043914[p40_array_index_2051017] ^ p40_literal_2043912[p40_array_index_2051028] ^ p40_literal_2043910[p40_array_index_2051019] ^ p40_array_index_2051029;
  assign p41_array_index_2051323_comb = p40_literal_2043918[p40_res7__518];
  assign p41_array_index_2051324_comb = p40_literal_2043920[p40_res7__516];
  assign p41_res7__528_comb = p40_literal_2043910[p41_res7__526_comb] ^ p40_literal_2043912[p40_res7__524] ^ p40_literal_2043914[p40_res7__522] ^ p40_literal_2043916[p40_res7__520] ^ p41_array_index_2051323_comb ^ p41_array_index_2051324_comb ^ p40_res7__514 ^ p40_literal_2043923[p40_res7__512] ^ p40_array_index_2051012 ^ p40_array_index_2051154 ^ p40_array_index_2051125 ^ p40_array_index_2051096 ^ p40_literal_2043914[p40_array_index_2051016] ^ p40_literal_2043912[p40_array_index_2051017] ^ p40_literal_2043910[p40_array_index_2051028] ^ p40_array_index_2051019;
  assign p41_array_index_2051334_comb = p40_literal_2043918[p40_res7__520];
  assign p41_array_index_2051335_comb = p40_literal_2043920[p40_res7__518];
  assign p41_res7__530_comb = p40_literal_2043910[p41_res7__528_comb] ^ p40_literal_2043912[p41_res7__526_comb] ^ p40_literal_2043914[p40_res7__524] ^ p40_literal_2043916[p40_res7__522] ^ p41_array_index_2051334_comb ^ p41_array_index_2051335_comb ^ p40_res7__516 ^ p40_literal_2043923[p40_res7__514] ^ p40_res7__512 ^ p40_array_index_2051167 ^ p40_array_index_2051139 ^ p40_array_index_2051110 ^ p40_literal_2043914[p40_array_index_2051015] ^ p40_literal_2043912[p40_array_index_2051016] ^ p40_literal_2043910[p40_array_index_2051017] ^ p40_array_index_2051028;
  assign p41_array_index_2051346_comb = p40_literal_2043920[p40_res7__520];
  assign p41_res7__532_comb = p40_literal_2043910[p41_res7__530_comb] ^ p40_literal_2043912[p41_res7__528_comb] ^ p40_literal_2043914[p41_res7__526_comb] ^ p40_literal_2043916[p40_res7__524] ^ p40_literal_2043918[p40_res7__522] ^ p41_array_index_2051346_comb ^ p40_res7__518 ^ p40_literal_2043923[p40_res7__516] ^ p40_res7__514 ^ p40_array_index_2051180 ^ p40_array_index_2051153 ^ p40_array_index_2051124 ^ p40_array_index_2051095 ^ p40_literal_2043912[p40_array_index_2051015] ^ p40_literal_2043910[p40_array_index_2051016] ^ p40_array_index_2051017;
  assign p41_array_index_2051356_comb = p40_literal_2043920[p40_res7__522];
  assign p41_res7__534_comb = p40_literal_2043910[p41_res7__532_comb] ^ p40_literal_2043912[p41_res7__530_comb] ^ p40_literal_2043914[p41_res7__528_comb] ^ p40_literal_2043916[p41_res7__526_comb] ^ p40_literal_2043918[p40_res7__524] ^ p41_array_index_2051356_comb ^ p40_res7__520 ^ p40_literal_2043923[p40_res7__518] ^ p40_res7__516 ^ p41_array_index_2051312_comb ^ p40_array_index_2051166 ^ p40_array_index_2051138 ^ p40_array_index_2051109 ^ p40_literal_2043912[p40_array_index_2051014] ^ p40_literal_2043910[p40_array_index_2051015] ^ p40_array_index_2051016;
  assign p41_res7__536_comb = p40_literal_2043910[p41_res7__534_comb] ^ p40_literal_2043912[p41_res7__532_comb] ^ p40_literal_2043914[p41_res7__530_comb] ^ p40_literal_2043916[p41_res7__528_comb] ^ p40_literal_2043918[p41_res7__526_comb] ^ p40_literal_2043920[p40_res7__524] ^ p40_res7__522 ^ p40_literal_2043923[p40_res7__520] ^ p40_res7__518 ^ p41_array_index_2051324_comb ^ p40_array_index_2051179 ^ p40_array_index_2051152 ^ p40_array_index_2051123 ^ p40_array_index_2051094 ^ p40_literal_2043910[p40_array_index_2051014] ^ p40_array_index_2051015;
  assign p41_res7__538_comb = p40_literal_2043910[p41_res7__536_comb] ^ p40_literal_2043912[p41_res7__534_comb] ^ p40_literal_2043914[p41_res7__532_comb] ^ p40_literal_2043916[p41_res7__530_comb] ^ p40_literal_2043918[p41_res7__528_comb] ^ p40_literal_2043920[p41_res7__526_comb] ^ p40_res7__524 ^ p40_literal_2043923[p40_res7__522] ^ p40_res7__520 ^ p41_array_index_2051335_comb ^ p41_array_index_2051311_comb ^ p40_array_index_2051165 ^ p40_array_index_2051137 ^ p40_array_index_2051108 ^ p40_literal_2043910[p40_array_index_2051013] ^ p40_array_index_2051014;

  // Registers for pipe stage 41:
  reg [127:0] p41_encoded;
  reg [127:0] p41_bit_slice_2043893;
  reg [127:0] p41_bit_slice_2044018;
  reg [127:0] p41_k3;
  reg [127:0] p41_k2;
  reg [127:0] p41_k5;
  reg [127:0] p41_k4;
  reg [7:0] p41_array_index_2051012;
  reg [7:0] p41_array_index_2051013;
  reg [7:0] p41_array_index_2051093;
  reg [7:0] p41_res7__512;
  reg [7:0] p41_array_index_2051107;
  reg [7:0] p41_res7__514;
  reg [7:0] p41_array_index_2051122;
  reg [7:0] p41_res7__516;
  reg [7:0] p41_array_index_2051136;
  reg [7:0] p41_res7__518;
  reg [7:0] p41_array_index_2051151;
  reg [7:0] p41_res7__520;
  reg [7:0] p41_array_index_2051164;
  reg [7:0] p41_res7__522;
  reg [7:0] p41_array_index_2051178;
  reg [7:0] p41_res7__524;
  reg [7:0] p41_array_index_2051310;
  reg [7:0] p41_res7__526;
  reg [7:0] p41_array_index_2051323;
  reg [7:0] p41_res7__528;
  reg [7:0] p41_array_index_2051334;
  reg [7:0] p41_res7__530;
  reg [7:0] p41_array_index_2051346;
  reg [7:0] p41_res7__532;
  reg [7:0] p41_array_index_2051356;
  reg [7:0] p41_res7__534;
  reg [7:0] p41_res7__536;
  reg [7:0] p41_res7__538;
  reg [7:0] p42_literal_2043896[256];
  reg [7:0] p42_literal_2043910[256];
  reg [7:0] p42_literal_2043912[256];
  reg [7:0] p42_literal_2043914[256];
  reg [7:0] p42_literal_2043916[256];
  reg [7:0] p42_literal_2043918[256];
  reg [7:0] p42_literal_2043920[256];
  reg [7:0] p42_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p41_encoded <= p40_encoded;
    p41_bit_slice_2043893 <= p40_bit_slice_2043893;
    p41_bit_slice_2044018 <= p40_bit_slice_2044018;
    p41_k3 <= p40_k3;
    p41_k2 <= p40_k2;
    p41_k5 <= p40_k5;
    p41_k4 <= p40_k4;
    p41_array_index_2051012 <= p40_array_index_2051012;
    p41_array_index_2051013 <= p40_array_index_2051013;
    p41_array_index_2051093 <= p40_array_index_2051093;
    p41_res7__512 <= p40_res7__512;
    p41_array_index_2051107 <= p40_array_index_2051107;
    p41_res7__514 <= p40_res7__514;
    p41_array_index_2051122 <= p40_array_index_2051122;
    p41_res7__516 <= p40_res7__516;
    p41_array_index_2051136 <= p40_array_index_2051136;
    p41_res7__518 <= p40_res7__518;
    p41_array_index_2051151 <= p40_array_index_2051151;
    p41_res7__520 <= p40_res7__520;
    p41_array_index_2051164 <= p40_array_index_2051164;
    p41_res7__522 <= p40_res7__522;
    p41_array_index_2051178 <= p40_array_index_2051178;
    p41_res7__524 <= p40_res7__524;
    p41_array_index_2051310 <= p41_array_index_2051310_comb;
    p41_res7__526 <= p41_res7__526_comb;
    p41_array_index_2051323 <= p41_array_index_2051323_comb;
    p41_res7__528 <= p41_res7__528_comb;
    p41_array_index_2051334 <= p41_array_index_2051334_comb;
    p41_res7__530 <= p41_res7__530_comb;
    p41_array_index_2051346 <= p41_array_index_2051346_comb;
    p41_res7__532 <= p41_res7__532_comb;
    p41_array_index_2051356 <= p41_array_index_2051356_comb;
    p41_res7__534 <= p41_res7__534_comb;
    p41_res7__536 <= p41_res7__536_comb;
    p41_res7__538 <= p41_res7__538_comb;
    p42_literal_2043896 <= p41_literal_2043896;
    p42_literal_2043910 <= p41_literal_2043910;
    p42_literal_2043912 <= p41_literal_2043912;
    p42_literal_2043914 <= p41_literal_2043914;
    p42_literal_2043916 <= p41_literal_2043916;
    p42_literal_2043918 <= p41_literal_2043918;
    p42_literal_2043920 <= p41_literal_2043920;
    p42_literal_2043923 <= p41_literal_2043923;
  end

  // ===== Pipe stage 42:
  wire [7:0] p42_res7__540_comb;
  wire [7:0] p42_res7__542_comb;
  wire [127:0] p42_res__16_comb;
  wire [127:0] p42_xor_2051482_comb;
  wire [127:0] p42_addedKey__49_comb;
  wire [7:0] p42_array_index_2051498_comb;
  wire [7:0] p42_array_index_2051499_comb;
  wire [7:0] p42_array_index_2051500_comb;
  wire [7:0] p42_array_index_2051501_comb;
  wire [7:0] p42_array_index_2051502_comb;
  wire [7:0] p42_array_index_2051503_comb;
  wire [7:0] p42_array_index_2051505_comb;
  wire [7:0] p42_array_index_2051507_comb;
  wire [7:0] p42_array_index_2051508_comb;
  wire [7:0] p42_array_index_2051509_comb;
  wire [7:0] p42_array_index_2051510_comb;
  wire [7:0] p42_array_index_2051511_comb;
  wire [7:0] p42_array_index_2051512_comb;
  wire [7:0] p42_array_index_2051514_comb;
  wire [7:0] p42_array_index_2051515_comb;
  wire [7:0] p42_array_index_2051516_comb;
  wire [7:0] p42_array_index_2051517_comb;
  wire [7:0] p42_array_index_2051518_comb;
  wire [7:0] p42_array_index_2051519_comb;
  wire [7:0] p42_array_index_2051520_comb;
  wire [7:0] p42_array_index_2051522_comb;
  wire [7:0] p42_res7__544_comb;
  wire [7:0] p42_array_index_2051531_comb;
  wire [7:0] p42_array_index_2051532_comb;
  wire [7:0] p42_array_index_2051533_comb;
  wire [7:0] p42_array_index_2051534_comb;
  wire [7:0] p42_array_index_2051535_comb;
  wire [7:0] p42_array_index_2051536_comb;
  wire [7:0] p42_res7__546_comb;
  wire [7:0] p42_array_index_2051546_comb;
  wire [7:0] p42_array_index_2051547_comb;
  wire [7:0] p42_array_index_2051548_comb;
  wire [7:0] p42_array_index_2051549_comb;
  wire [7:0] p42_array_index_2051550_comb;
  wire [7:0] p42_res7__548_comb;
  wire [7:0] p42_array_index_2051560_comb;
  wire [7:0] p42_array_index_2051561_comb;
  wire [7:0] p42_array_index_2051562_comb;
  wire [7:0] p42_array_index_2051563_comb;
  wire [7:0] p42_array_index_2051564_comb;
  wire [7:0] p42_res7__550_comb;
  assign p42_res7__540_comb = p41_literal_2043910[p41_res7__538] ^ p41_literal_2043912[p41_res7__536] ^ p41_literal_2043914[p41_res7__534] ^ p41_literal_2043916[p41_res7__532] ^ p41_literal_2043918[p41_res7__530] ^ p41_literal_2043920[p41_res7__528] ^ p41_res7__526 ^ p41_literal_2043923[p41_res7__524] ^ p41_res7__522 ^ p41_array_index_2051346 ^ p41_array_index_2051323 ^ p41_array_index_2051178 ^ p41_array_index_2051151 ^ p41_array_index_2051122 ^ p41_array_index_2051093 ^ p41_array_index_2051013;
  assign p42_res7__542_comb = p41_literal_2043910[p42_res7__540_comb] ^ p41_literal_2043912[p41_res7__538] ^ p41_literal_2043914[p41_res7__536] ^ p41_literal_2043916[p41_res7__534] ^ p41_literal_2043918[p41_res7__532] ^ p41_literal_2043920[p41_res7__530] ^ p41_res7__528 ^ p41_literal_2043923[p41_res7__526] ^ p41_res7__524 ^ p41_array_index_2051356 ^ p41_array_index_2051334 ^ p41_array_index_2051310 ^ p41_array_index_2051164 ^ p41_array_index_2051136 ^ p41_array_index_2051107 ^ p41_array_index_2051012;
  assign p42_res__16_comb = {p42_res7__542_comb, p42_res7__540_comb, p41_res7__538, p41_res7__536, p41_res7__534, p41_res7__532, p41_res7__530, p41_res7__528, p41_res7__526, p41_res7__524, p41_res7__522, p41_res7__520, p41_res7__518, p41_res7__516, p41_res7__514, p41_res7__512};
  assign p42_xor_2051482_comb = p42_res__16_comb ^ p41_k5;
  assign p42_addedKey__49_comb = p42_xor_2051482_comb ^ 128'hf335_80c8_d79a_5862_237b_38e3_375c_bf12;
  assign p42_array_index_2051498_comb = p41_literal_2043896[p42_addedKey__49_comb[127:120]];
  assign p42_array_index_2051499_comb = p41_literal_2043896[p42_addedKey__49_comb[119:112]];
  assign p42_array_index_2051500_comb = p41_literal_2043896[p42_addedKey__49_comb[111:104]];
  assign p42_array_index_2051501_comb = p41_literal_2043896[p42_addedKey__49_comb[103:96]];
  assign p42_array_index_2051502_comb = p41_literal_2043896[p42_addedKey__49_comb[95:88]];
  assign p42_array_index_2051503_comb = p41_literal_2043896[p42_addedKey__49_comb[87:80]];
  assign p42_array_index_2051505_comb = p41_literal_2043896[p42_addedKey__49_comb[71:64]];
  assign p42_array_index_2051507_comb = p41_literal_2043896[p42_addedKey__49_comb[55:48]];
  assign p42_array_index_2051508_comb = p41_literal_2043896[p42_addedKey__49_comb[47:40]];
  assign p42_array_index_2051509_comb = p41_literal_2043896[p42_addedKey__49_comb[39:32]];
  assign p42_array_index_2051510_comb = p41_literal_2043896[p42_addedKey__49_comb[31:24]];
  assign p42_array_index_2051511_comb = p41_literal_2043896[p42_addedKey__49_comb[23:16]];
  assign p42_array_index_2051512_comb = p41_literal_2043896[p42_addedKey__49_comb[15:8]];
  assign p42_array_index_2051514_comb = p41_literal_2043910[p42_array_index_2051498_comb];
  assign p42_array_index_2051515_comb = p41_literal_2043912[p42_array_index_2051499_comb];
  assign p42_array_index_2051516_comb = p41_literal_2043914[p42_array_index_2051500_comb];
  assign p42_array_index_2051517_comb = p41_literal_2043916[p42_array_index_2051501_comb];
  assign p42_array_index_2051518_comb = p41_literal_2043918[p42_array_index_2051502_comb];
  assign p42_array_index_2051519_comb = p41_literal_2043920[p42_array_index_2051503_comb];
  assign p42_array_index_2051520_comb = p41_literal_2043896[p42_addedKey__49_comb[79:72]];
  assign p42_array_index_2051522_comb = p41_literal_2043896[p42_addedKey__49_comb[63:56]];
  assign p42_res7__544_comb = p42_array_index_2051514_comb ^ p42_array_index_2051515_comb ^ p42_array_index_2051516_comb ^ p42_array_index_2051517_comb ^ p42_array_index_2051518_comb ^ p42_array_index_2051519_comb ^ p42_array_index_2051520_comb ^ p41_literal_2043923[p42_array_index_2051505_comb] ^ p42_array_index_2051522_comb ^ p41_literal_2043920[p42_array_index_2051507_comb] ^ p41_literal_2043918[p42_array_index_2051508_comb] ^ p41_literal_2043916[p42_array_index_2051509_comb] ^ p41_literal_2043914[p42_array_index_2051510_comb] ^ p41_literal_2043912[p42_array_index_2051511_comb] ^ p41_literal_2043910[p42_array_index_2051512_comb] ^ p41_literal_2043896[p42_addedKey__49_comb[7:0]];
  assign p42_array_index_2051531_comb = p41_literal_2043910[p42_res7__544_comb];
  assign p42_array_index_2051532_comb = p41_literal_2043912[p42_array_index_2051498_comb];
  assign p42_array_index_2051533_comb = p41_literal_2043914[p42_array_index_2051499_comb];
  assign p42_array_index_2051534_comb = p41_literal_2043916[p42_array_index_2051500_comb];
  assign p42_array_index_2051535_comb = p41_literal_2043918[p42_array_index_2051501_comb];
  assign p42_array_index_2051536_comb = p41_literal_2043920[p42_array_index_2051502_comb];
  assign p42_res7__546_comb = p42_array_index_2051531_comb ^ p42_array_index_2051532_comb ^ p42_array_index_2051533_comb ^ p42_array_index_2051534_comb ^ p42_array_index_2051535_comb ^ p42_array_index_2051536_comb ^ p42_array_index_2051503_comb ^ p41_literal_2043923[p42_array_index_2051520_comb] ^ p42_array_index_2051505_comb ^ p41_literal_2043920[p42_array_index_2051522_comb] ^ p41_literal_2043918[p42_array_index_2051507_comb] ^ p41_literal_2043916[p42_array_index_2051508_comb] ^ p41_literal_2043914[p42_array_index_2051509_comb] ^ p41_literal_2043912[p42_array_index_2051510_comb] ^ p41_literal_2043910[p42_array_index_2051511_comb] ^ p42_array_index_2051512_comb;
  assign p42_array_index_2051546_comb = p41_literal_2043912[p42_res7__544_comb];
  assign p42_array_index_2051547_comb = p41_literal_2043914[p42_array_index_2051498_comb];
  assign p42_array_index_2051548_comb = p41_literal_2043916[p42_array_index_2051499_comb];
  assign p42_array_index_2051549_comb = p41_literal_2043918[p42_array_index_2051500_comb];
  assign p42_array_index_2051550_comb = p41_literal_2043920[p42_array_index_2051501_comb];
  assign p42_res7__548_comb = p41_literal_2043910[p42_res7__546_comb] ^ p42_array_index_2051546_comb ^ p42_array_index_2051547_comb ^ p42_array_index_2051548_comb ^ p42_array_index_2051549_comb ^ p42_array_index_2051550_comb ^ p42_array_index_2051502_comb ^ p41_literal_2043923[p42_array_index_2051503_comb] ^ p42_array_index_2051520_comb ^ p41_literal_2043920[p42_array_index_2051505_comb] ^ p41_literal_2043918[p42_array_index_2051522_comb] ^ p41_literal_2043916[p42_array_index_2051507_comb] ^ p41_literal_2043914[p42_array_index_2051508_comb] ^ p41_literal_2043912[p42_array_index_2051509_comb] ^ p41_literal_2043910[p42_array_index_2051510_comb] ^ p42_array_index_2051511_comb;
  assign p42_array_index_2051560_comb = p41_literal_2043912[p42_res7__546_comb];
  assign p42_array_index_2051561_comb = p41_literal_2043914[p42_res7__544_comb];
  assign p42_array_index_2051562_comb = p41_literal_2043916[p42_array_index_2051498_comb];
  assign p42_array_index_2051563_comb = p41_literal_2043918[p42_array_index_2051499_comb];
  assign p42_array_index_2051564_comb = p41_literal_2043920[p42_array_index_2051500_comb];
  assign p42_res7__550_comb = p41_literal_2043910[p42_res7__548_comb] ^ p42_array_index_2051560_comb ^ p42_array_index_2051561_comb ^ p42_array_index_2051562_comb ^ p42_array_index_2051563_comb ^ p42_array_index_2051564_comb ^ p42_array_index_2051501_comb ^ p41_literal_2043923[p42_array_index_2051502_comb] ^ p42_array_index_2051503_comb ^ p41_literal_2043920[p42_array_index_2051520_comb] ^ p41_literal_2043918[p42_array_index_2051505_comb] ^ p41_literal_2043916[p42_array_index_2051522_comb] ^ p41_literal_2043914[p42_array_index_2051507_comb] ^ p41_literal_2043912[p42_array_index_2051508_comb] ^ p41_literal_2043910[p42_array_index_2051509_comb] ^ p42_array_index_2051510_comb;

  // Registers for pipe stage 42:
  reg [127:0] p42_encoded;
  reg [127:0] p42_bit_slice_2043893;
  reg [127:0] p42_bit_slice_2044018;
  reg [127:0] p42_k3;
  reg [127:0] p42_k2;
  reg [127:0] p42_k5;
  reg [127:0] p42_k4;
  reg [127:0] p42_xor_2051482;
  reg [7:0] p42_array_index_2051498;
  reg [7:0] p42_array_index_2051499;
  reg [7:0] p42_array_index_2051500;
  reg [7:0] p42_array_index_2051501;
  reg [7:0] p42_array_index_2051502;
  reg [7:0] p42_array_index_2051503;
  reg [7:0] p42_array_index_2051505;
  reg [7:0] p42_array_index_2051507;
  reg [7:0] p42_array_index_2051508;
  reg [7:0] p42_array_index_2051509;
  reg [7:0] p42_array_index_2051514;
  reg [7:0] p42_array_index_2051515;
  reg [7:0] p42_array_index_2051516;
  reg [7:0] p42_array_index_2051517;
  reg [7:0] p42_array_index_2051518;
  reg [7:0] p42_array_index_2051519;
  reg [7:0] p42_array_index_2051520;
  reg [7:0] p42_array_index_2051522;
  reg [7:0] p42_res7__544;
  reg [7:0] p42_array_index_2051531;
  reg [7:0] p42_array_index_2051532;
  reg [7:0] p42_array_index_2051533;
  reg [7:0] p42_array_index_2051534;
  reg [7:0] p42_array_index_2051535;
  reg [7:0] p42_array_index_2051536;
  reg [7:0] p42_res7__546;
  reg [7:0] p42_array_index_2051546;
  reg [7:0] p42_array_index_2051547;
  reg [7:0] p42_array_index_2051548;
  reg [7:0] p42_array_index_2051549;
  reg [7:0] p42_array_index_2051550;
  reg [7:0] p42_res7__548;
  reg [7:0] p42_array_index_2051560;
  reg [7:0] p42_array_index_2051561;
  reg [7:0] p42_array_index_2051562;
  reg [7:0] p42_array_index_2051563;
  reg [7:0] p42_array_index_2051564;
  reg [7:0] p42_res7__550;
  reg [7:0] p43_literal_2043896[256];
  reg [7:0] p43_literal_2043910[256];
  reg [7:0] p43_literal_2043912[256];
  reg [7:0] p43_literal_2043914[256];
  reg [7:0] p43_literal_2043916[256];
  reg [7:0] p43_literal_2043918[256];
  reg [7:0] p43_literal_2043920[256];
  reg [7:0] p43_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p42_encoded <= p41_encoded;
    p42_bit_slice_2043893 <= p41_bit_slice_2043893;
    p42_bit_slice_2044018 <= p41_bit_slice_2044018;
    p42_k3 <= p41_k3;
    p42_k2 <= p41_k2;
    p42_k5 <= p41_k5;
    p42_k4 <= p41_k4;
    p42_xor_2051482 <= p42_xor_2051482_comb;
    p42_array_index_2051498 <= p42_array_index_2051498_comb;
    p42_array_index_2051499 <= p42_array_index_2051499_comb;
    p42_array_index_2051500 <= p42_array_index_2051500_comb;
    p42_array_index_2051501 <= p42_array_index_2051501_comb;
    p42_array_index_2051502 <= p42_array_index_2051502_comb;
    p42_array_index_2051503 <= p42_array_index_2051503_comb;
    p42_array_index_2051505 <= p42_array_index_2051505_comb;
    p42_array_index_2051507 <= p42_array_index_2051507_comb;
    p42_array_index_2051508 <= p42_array_index_2051508_comb;
    p42_array_index_2051509 <= p42_array_index_2051509_comb;
    p42_array_index_2051514 <= p42_array_index_2051514_comb;
    p42_array_index_2051515 <= p42_array_index_2051515_comb;
    p42_array_index_2051516 <= p42_array_index_2051516_comb;
    p42_array_index_2051517 <= p42_array_index_2051517_comb;
    p42_array_index_2051518 <= p42_array_index_2051518_comb;
    p42_array_index_2051519 <= p42_array_index_2051519_comb;
    p42_array_index_2051520 <= p42_array_index_2051520_comb;
    p42_array_index_2051522 <= p42_array_index_2051522_comb;
    p42_res7__544 <= p42_res7__544_comb;
    p42_array_index_2051531 <= p42_array_index_2051531_comb;
    p42_array_index_2051532 <= p42_array_index_2051532_comb;
    p42_array_index_2051533 <= p42_array_index_2051533_comb;
    p42_array_index_2051534 <= p42_array_index_2051534_comb;
    p42_array_index_2051535 <= p42_array_index_2051535_comb;
    p42_array_index_2051536 <= p42_array_index_2051536_comb;
    p42_res7__546 <= p42_res7__546_comb;
    p42_array_index_2051546 <= p42_array_index_2051546_comb;
    p42_array_index_2051547 <= p42_array_index_2051547_comb;
    p42_array_index_2051548 <= p42_array_index_2051548_comb;
    p42_array_index_2051549 <= p42_array_index_2051549_comb;
    p42_array_index_2051550 <= p42_array_index_2051550_comb;
    p42_res7__548 <= p42_res7__548_comb;
    p42_array_index_2051560 <= p42_array_index_2051560_comb;
    p42_array_index_2051561 <= p42_array_index_2051561_comb;
    p42_array_index_2051562 <= p42_array_index_2051562_comb;
    p42_array_index_2051563 <= p42_array_index_2051563_comb;
    p42_array_index_2051564 <= p42_array_index_2051564_comb;
    p42_res7__550 <= p42_res7__550_comb;
    p43_literal_2043896 <= p42_literal_2043896;
    p43_literal_2043910 <= p42_literal_2043910;
    p43_literal_2043912 <= p42_literal_2043912;
    p43_literal_2043914 <= p42_literal_2043914;
    p43_literal_2043916 <= p42_literal_2043916;
    p43_literal_2043918 <= p42_literal_2043918;
    p43_literal_2043920 <= p42_literal_2043920;
    p43_literal_2043923 <= p42_literal_2043923;
  end

  // ===== Pipe stage 43:
  wire [7:0] p43_array_index_2051683_comb;
  wire [7:0] p43_array_index_2051684_comb;
  wire [7:0] p43_array_index_2051685_comb;
  wire [7:0] p43_array_index_2051686_comb;
  wire [7:0] p43_res7__552_comb;
  wire [7:0] p43_array_index_2051696_comb;
  wire [7:0] p43_array_index_2051697_comb;
  wire [7:0] p43_array_index_2051698_comb;
  wire [7:0] p43_array_index_2051699_comb;
  wire [7:0] p43_res7__554_comb;
  wire [7:0] p43_array_index_2051710_comb;
  wire [7:0] p43_array_index_2051711_comb;
  wire [7:0] p43_array_index_2051712_comb;
  wire [7:0] p43_res7__556_comb;
  wire [7:0] p43_array_index_2051722_comb;
  wire [7:0] p43_array_index_2051723_comb;
  wire [7:0] p43_array_index_2051724_comb;
  wire [7:0] p43_res7__558_comb;
  wire [7:0] p43_array_index_2051735_comb;
  wire [7:0] p43_array_index_2051736_comb;
  wire [7:0] p43_res7__560_comb;
  wire [7:0] p43_array_index_2051746_comb;
  wire [7:0] p43_array_index_2051747_comb;
  wire [7:0] p43_res7__562_comb;
  wire [7:0] p43_array_index_2051758_comb;
  wire [7:0] p43_res7__564_comb;
  assign p43_array_index_2051683_comb = p42_literal_2043914[p42_res7__546];
  assign p43_array_index_2051684_comb = p42_literal_2043916[p42_res7__544];
  assign p43_array_index_2051685_comb = p42_literal_2043918[p42_array_index_2051498];
  assign p43_array_index_2051686_comb = p42_literal_2043920[p42_array_index_2051499];
  assign p43_res7__552_comb = p42_literal_2043910[p42_res7__550] ^ p42_literal_2043912[p42_res7__548] ^ p43_array_index_2051683_comb ^ p43_array_index_2051684_comb ^ p43_array_index_2051685_comb ^ p43_array_index_2051686_comb ^ p42_array_index_2051500 ^ p42_literal_2043923[p42_array_index_2051501] ^ p42_array_index_2051502 ^ p42_array_index_2051519 ^ p42_literal_2043918[p42_array_index_2051520] ^ p42_literal_2043916[p42_array_index_2051505] ^ p42_literal_2043914[p42_array_index_2051522] ^ p42_literal_2043912[p42_array_index_2051507] ^ p42_literal_2043910[p42_array_index_2051508] ^ p42_array_index_2051509;
  assign p43_array_index_2051696_comb = p42_literal_2043914[p42_res7__548];
  assign p43_array_index_2051697_comb = p42_literal_2043916[p42_res7__546];
  assign p43_array_index_2051698_comb = p42_literal_2043918[p42_res7__544];
  assign p43_array_index_2051699_comb = p42_literal_2043920[p42_array_index_2051498];
  assign p43_res7__554_comb = p42_literal_2043910[p43_res7__552_comb] ^ p42_literal_2043912[p42_res7__550] ^ p43_array_index_2051696_comb ^ p43_array_index_2051697_comb ^ p43_array_index_2051698_comb ^ p43_array_index_2051699_comb ^ p42_array_index_2051499 ^ p42_literal_2043923[p42_array_index_2051500] ^ p42_array_index_2051501 ^ p42_array_index_2051536 ^ p42_literal_2043918[p42_array_index_2051503] ^ p42_literal_2043916[p42_array_index_2051520] ^ p42_literal_2043914[p42_array_index_2051505] ^ p42_literal_2043912[p42_array_index_2051522] ^ p42_literal_2043910[p42_array_index_2051507] ^ p42_array_index_2051508;
  assign p43_array_index_2051710_comb = p42_literal_2043916[p42_res7__548];
  assign p43_array_index_2051711_comb = p42_literal_2043918[p42_res7__546];
  assign p43_array_index_2051712_comb = p42_literal_2043920[p42_res7__544];
  assign p43_res7__556_comb = p42_literal_2043910[p43_res7__554_comb] ^ p42_literal_2043912[p43_res7__552_comb] ^ p42_literal_2043914[p42_res7__550] ^ p43_array_index_2051710_comb ^ p43_array_index_2051711_comb ^ p43_array_index_2051712_comb ^ p42_array_index_2051498 ^ p42_literal_2043923[p42_array_index_2051499] ^ p42_array_index_2051500 ^ p42_array_index_2051550 ^ p42_array_index_2051518 ^ p42_literal_2043916[p42_array_index_2051503] ^ p42_literal_2043914[p42_array_index_2051520] ^ p42_literal_2043912[p42_array_index_2051505] ^ p42_literal_2043910[p42_array_index_2051522] ^ p42_array_index_2051507;
  assign p43_array_index_2051722_comb = p42_literal_2043916[p42_res7__550];
  assign p43_array_index_2051723_comb = p42_literal_2043918[p42_res7__548];
  assign p43_array_index_2051724_comb = p42_literal_2043920[p42_res7__546];
  assign p43_res7__558_comb = p42_literal_2043910[p43_res7__556_comb] ^ p42_literal_2043912[p43_res7__554_comb] ^ p42_literal_2043914[p43_res7__552_comb] ^ p43_array_index_2051722_comb ^ p43_array_index_2051723_comb ^ p43_array_index_2051724_comb ^ p42_res7__544 ^ p42_literal_2043923[p42_array_index_2051498] ^ p42_array_index_2051499 ^ p42_array_index_2051564 ^ p42_array_index_2051535 ^ p42_literal_2043916[p42_array_index_2051502] ^ p42_literal_2043914[p42_array_index_2051503] ^ p42_literal_2043912[p42_array_index_2051520] ^ p42_literal_2043910[p42_array_index_2051505] ^ p42_array_index_2051522;
  assign p43_array_index_2051735_comb = p42_literal_2043918[p42_res7__550];
  assign p43_array_index_2051736_comb = p42_literal_2043920[p42_res7__548];
  assign p43_res7__560_comb = p42_literal_2043910[p43_res7__558_comb] ^ p42_literal_2043912[p43_res7__556_comb] ^ p42_literal_2043914[p43_res7__554_comb] ^ p42_literal_2043916[p43_res7__552_comb] ^ p43_array_index_2051735_comb ^ p43_array_index_2051736_comb ^ p42_res7__546 ^ p42_literal_2043923[p42_res7__544] ^ p42_array_index_2051498 ^ p43_array_index_2051686_comb ^ p42_array_index_2051549 ^ p42_array_index_2051517 ^ p42_literal_2043914[p42_array_index_2051502] ^ p42_literal_2043912[p42_array_index_2051503] ^ p42_literal_2043910[p42_array_index_2051520] ^ p42_array_index_2051505;
  assign p43_array_index_2051746_comb = p42_literal_2043918[p43_res7__552_comb];
  assign p43_array_index_2051747_comb = p42_literal_2043920[p42_res7__550];
  assign p43_res7__562_comb = p42_literal_2043910[p43_res7__560_comb] ^ p42_literal_2043912[p43_res7__558_comb] ^ p42_literal_2043914[p43_res7__556_comb] ^ p42_literal_2043916[p43_res7__554_comb] ^ p43_array_index_2051746_comb ^ p43_array_index_2051747_comb ^ p42_res7__548 ^ p42_literal_2043923[p42_res7__546] ^ p42_res7__544 ^ p43_array_index_2051699_comb ^ p42_array_index_2051563 ^ p42_array_index_2051534 ^ p42_literal_2043914[p42_array_index_2051501] ^ p42_literal_2043912[p42_array_index_2051502] ^ p42_literal_2043910[p42_array_index_2051503] ^ p42_array_index_2051520;
  assign p43_array_index_2051758_comb = p42_literal_2043920[p43_res7__552_comb];
  assign p43_res7__564_comb = p42_literal_2043910[p43_res7__562_comb] ^ p42_literal_2043912[p43_res7__560_comb] ^ p42_literal_2043914[p43_res7__558_comb] ^ p42_literal_2043916[p43_res7__556_comb] ^ p42_literal_2043918[p43_res7__554_comb] ^ p43_array_index_2051758_comb ^ p42_res7__550 ^ p42_literal_2043923[p42_res7__548] ^ p42_res7__546 ^ p43_array_index_2051712_comb ^ p43_array_index_2051685_comb ^ p42_array_index_2051548 ^ p42_array_index_2051516 ^ p42_literal_2043912[p42_array_index_2051501] ^ p42_literal_2043910[p42_array_index_2051502] ^ p42_array_index_2051503;

  // Registers for pipe stage 43:
  reg [127:0] p43_encoded;
  reg [127:0] p43_bit_slice_2043893;
  reg [127:0] p43_bit_slice_2044018;
  reg [127:0] p43_k3;
  reg [127:0] p43_k2;
  reg [127:0] p43_k5;
  reg [127:0] p43_k4;
  reg [127:0] p43_xor_2051482;
  reg [7:0] p43_array_index_2051498;
  reg [7:0] p43_array_index_2051499;
  reg [7:0] p43_array_index_2051500;
  reg [7:0] p43_array_index_2051501;
  reg [7:0] p43_array_index_2051502;
  reg [7:0] p43_array_index_2051514;
  reg [7:0] p43_array_index_2051515;
  reg [7:0] p43_res7__544;
  reg [7:0] p43_array_index_2051531;
  reg [7:0] p43_array_index_2051532;
  reg [7:0] p43_array_index_2051533;
  reg [7:0] p43_res7__546;
  reg [7:0] p43_array_index_2051546;
  reg [7:0] p43_array_index_2051547;
  reg [7:0] p43_res7__548;
  reg [7:0] p43_array_index_2051560;
  reg [7:0] p43_array_index_2051561;
  reg [7:0] p43_array_index_2051562;
  reg [7:0] p43_res7__550;
  reg [7:0] p43_array_index_2051683;
  reg [7:0] p43_array_index_2051684;
  reg [7:0] p43_res7__552;
  reg [7:0] p43_array_index_2051696;
  reg [7:0] p43_array_index_2051697;
  reg [7:0] p43_array_index_2051698;
  reg [7:0] p43_res7__554;
  reg [7:0] p43_array_index_2051710;
  reg [7:0] p43_array_index_2051711;
  reg [7:0] p43_res7__556;
  reg [7:0] p43_array_index_2051722;
  reg [7:0] p43_array_index_2051723;
  reg [7:0] p43_array_index_2051724;
  reg [7:0] p43_res7__558;
  reg [7:0] p43_array_index_2051735;
  reg [7:0] p43_array_index_2051736;
  reg [7:0] p43_res7__560;
  reg [7:0] p43_array_index_2051746;
  reg [7:0] p43_array_index_2051747;
  reg [7:0] p43_res7__562;
  reg [7:0] p43_array_index_2051758;
  reg [7:0] p43_res7__564;
  reg [7:0] p44_literal_2043896[256];
  reg [7:0] p44_literal_2043910[256];
  reg [7:0] p44_literal_2043912[256];
  reg [7:0] p44_literal_2043914[256];
  reg [7:0] p44_literal_2043916[256];
  reg [7:0] p44_literal_2043918[256];
  reg [7:0] p44_literal_2043920[256];
  reg [7:0] p44_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p43_encoded <= p42_encoded;
    p43_bit_slice_2043893 <= p42_bit_slice_2043893;
    p43_bit_slice_2044018 <= p42_bit_slice_2044018;
    p43_k3 <= p42_k3;
    p43_k2 <= p42_k2;
    p43_k5 <= p42_k5;
    p43_k4 <= p42_k4;
    p43_xor_2051482 <= p42_xor_2051482;
    p43_array_index_2051498 <= p42_array_index_2051498;
    p43_array_index_2051499 <= p42_array_index_2051499;
    p43_array_index_2051500 <= p42_array_index_2051500;
    p43_array_index_2051501 <= p42_array_index_2051501;
    p43_array_index_2051502 <= p42_array_index_2051502;
    p43_array_index_2051514 <= p42_array_index_2051514;
    p43_array_index_2051515 <= p42_array_index_2051515;
    p43_res7__544 <= p42_res7__544;
    p43_array_index_2051531 <= p42_array_index_2051531;
    p43_array_index_2051532 <= p42_array_index_2051532;
    p43_array_index_2051533 <= p42_array_index_2051533;
    p43_res7__546 <= p42_res7__546;
    p43_array_index_2051546 <= p42_array_index_2051546;
    p43_array_index_2051547 <= p42_array_index_2051547;
    p43_res7__548 <= p42_res7__548;
    p43_array_index_2051560 <= p42_array_index_2051560;
    p43_array_index_2051561 <= p42_array_index_2051561;
    p43_array_index_2051562 <= p42_array_index_2051562;
    p43_res7__550 <= p42_res7__550;
    p43_array_index_2051683 <= p43_array_index_2051683_comb;
    p43_array_index_2051684 <= p43_array_index_2051684_comb;
    p43_res7__552 <= p43_res7__552_comb;
    p43_array_index_2051696 <= p43_array_index_2051696_comb;
    p43_array_index_2051697 <= p43_array_index_2051697_comb;
    p43_array_index_2051698 <= p43_array_index_2051698_comb;
    p43_res7__554 <= p43_res7__554_comb;
    p43_array_index_2051710 <= p43_array_index_2051710_comb;
    p43_array_index_2051711 <= p43_array_index_2051711_comb;
    p43_res7__556 <= p43_res7__556_comb;
    p43_array_index_2051722 <= p43_array_index_2051722_comb;
    p43_array_index_2051723 <= p43_array_index_2051723_comb;
    p43_array_index_2051724 <= p43_array_index_2051724_comb;
    p43_res7__558 <= p43_res7__558_comb;
    p43_array_index_2051735 <= p43_array_index_2051735_comb;
    p43_array_index_2051736 <= p43_array_index_2051736_comb;
    p43_res7__560 <= p43_res7__560_comb;
    p43_array_index_2051746 <= p43_array_index_2051746_comb;
    p43_array_index_2051747 <= p43_array_index_2051747_comb;
    p43_res7__562 <= p43_res7__562_comb;
    p43_array_index_2051758 <= p43_array_index_2051758_comb;
    p43_res7__564 <= p43_res7__564_comb;
    p44_literal_2043896 <= p43_literal_2043896;
    p44_literal_2043910 <= p43_literal_2043910;
    p44_literal_2043912 <= p43_literal_2043912;
    p44_literal_2043914 <= p43_literal_2043914;
    p44_literal_2043916 <= p43_literal_2043916;
    p44_literal_2043918 <= p43_literal_2043918;
    p44_literal_2043920 <= p43_literal_2043920;
    p44_literal_2043923 <= p43_literal_2043923;
  end

  // ===== Pipe stage 44:
  wire [7:0] p44_array_index_2051882_comb;
  wire [7:0] p44_res7__566_comb;
  wire [7:0] p44_res7__568_comb;
  wire [7:0] p44_res7__570_comb;
  wire [7:0] p44_res7__572_comb;
  wire [7:0] p44_res7__574_comb;
  wire [127:0] p44_res__17_comb;
  wire [127:0] p44_xor_2051922_comb;
  wire [127:0] p44_addedKey__50_comb;
  wire [7:0] p44_array_index_2051938_comb;
  wire [7:0] p44_array_index_2051939_comb;
  wire [7:0] p44_array_index_2051940_comb;
  wire [7:0] p44_array_index_2051941_comb;
  wire [7:0] p44_array_index_2051942_comb;
  wire [7:0] p44_array_index_2051943_comb;
  wire [7:0] p44_array_index_2051945_comb;
  wire [7:0] p44_array_index_2051947_comb;
  wire [7:0] p44_array_index_2051948_comb;
  wire [7:0] p44_array_index_2051949_comb;
  wire [7:0] p44_array_index_2051950_comb;
  wire [7:0] p44_array_index_2051951_comb;
  wire [7:0] p44_array_index_2051952_comb;
  wire [7:0] p44_array_index_2051954_comb;
  wire [7:0] p44_array_index_2051955_comb;
  wire [7:0] p44_array_index_2051956_comb;
  wire [7:0] p44_array_index_2051957_comb;
  wire [7:0] p44_array_index_2051958_comb;
  wire [7:0] p44_array_index_2051959_comb;
  wire [7:0] p44_array_index_2051960_comb;
  wire [7:0] p44_array_index_2051962_comb;
  wire [7:0] p44_res7__576_comb;
  assign p44_array_index_2051882_comb = p43_literal_2043920[p43_res7__554];
  assign p44_res7__566_comb = p43_literal_2043910[p43_res7__564] ^ p43_literal_2043912[p43_res7__562] ^ p43_literal_2043914[p43_res7__560] ^ p43_literal_2043916[p43_res7__558] ^ p43_literal_2043918[p43_res7__556] ^ p44_array_index_2051882_comb ^ p43_res7__552 ^ p43_literal_2043923[p43_res7__550] ^ p43_res7__548 ^ p43_array_index_2051724 ^ p43_array_index_2051698 ^ p43_array_index_2051562 ^ p43_array_index_2051533 ^ p43_literal_2043912[p43_array_index_2051500] ^ p43_literal_2043910[p43_array_index_2051501] ^ p43_array_index_2051502;
  assign p44_res7__568_comb = p43_literal_2043910[p44_res7__566_comb] ^ p43_literal_2043912[p43_res7__564] ^ p43_literal_2043914[p43_res7__562] ^ p43_literal_2043916[p43_res7__560] ^ p43_literal_2043918[p43_res7__558] ^ p43_literal_2043920[p43_res7__556] ^ p43_res7__554 ^ p43_literal_2043923[p43_res7__552] ^ p43_res7__550 ^ p43_array_index_2051736 ^ p43_array_index_2051711 ^ p43_array_index_2051684 ^ p43_array_index_2051547 ^ p43_array_index_2051515 ^ p43_literal_2043910[p43_array_index_2051500] ^ p43_array_index_2051501;
  assign p44_res7__570_comb = p43_literal_2043910[p44_res7__568_comb] ^ p43_literal_2043912[p44_res7__566_comb] ^ p43_literal_2043914[p43_res7__564] ^ p43_literal_2043916[p43_res7__562] ^ p43_literal_2043918[p43_res7__560] ^ p43_literal_2043920[p43_res7__558] ^ p43_res7__556 ^ p43_literal_2043923[p43_res7__554] ^ p43_res7__552 ^ p43_array_index_2051747 ^ p43_array_index_2051723 ^ p43_array_index_2051697 ^ p43_array_index_2051561 ^ p43_array_index_2051532 ^ p43_literal_2043910[p43_array_index_2051499] ^ p43_array_index_2051500;
  assign p44_res7__572_comb = p43_literal_2043910[p44_res7__570_comb] ^ p43_literal_2043912[p44_res7__568_comb] ^ p43_literal_2043914[p44_res7__566_comb] ^ p43_literal_2043916[p43_res7__564] ^ p43_literal_2043918[p43_res7__562] ^ p43_literal_2043920[p43_res7__560] ^ p43_res7__558 ^ p43_literal_2043923[p43_res7__556] ^ p43_res7__554 ^ p43_array_index_2051758 ^ p43_array_index_2051735 ^ p43_array_index_2051710 ^ p43_array_index_2051683 ^ p43_array_index_2051546 ^ p43_array_index_2051514 ^ p43_array_index_2051499;
  assign p44_res7__574_comb = p43_literal_2043910[p44_res7__572_comb] ^ p43_literal_2043912[p44_res7__570_comb] ^ p43_literal_2043914[p44_res7__568_comb] ^ p43_literal_2043916[p44_res7__566_comb] ^ p43_literal_2043918[p43_res7__564] ^ p43_literal_2043920[p43_res7__562] ^ p43_res7__560 ^ p43_literal_2043923[p43_res7__558] ^ p43_res7__556 ^ p44_array_index_2051882_comb ^ p43_array_index_2051746 ^ p43_array_index_2051722 ^ p43_array_index_2051696 ^ p43_array_index_2051560 ^ p43_array_index_2051531 ^ p43_array_index_2051498;
  assign p44_res__17_comb = {p44_res7__574_comb, p44_res7__572_comb, p44_res7__570_comb, p44_res7__568_comb, p44_res7__566_comb, p43_res7__564, p43_res7__562, p43_res7__560, p43_res7__558, p43_res7__556, p43_res7__554, p43_res7__552, p43_res7__550, p43_res7__548, p43_res7__546, p43_res7__544};
  assign p44_xor_2051922_comb = p44_res__17_comb ^ p43_k4;
  assign p44_addedKey__50_comb = p44_xor_2051922_comb ^ 128'h9d97_f6ba_bbd2_22da_7e5c_85f3_ead8_2b13;
  assign p44_array_index_2051938_comb = p43_literal_2043896[p44_addedKey__50_comb[127:120]];
  assign p44_array_index_2051939_comb = p43_literal_2043896[p44_addedKey__50_comb[119:112]];
  assign p44_array_index_2051940_comb = p43_literal_2043896[p44_addedKey__50_comb[111:104]];
  assign p44_array_index_2051941_comb = p43_literal_2043896[p44_addedKey__50_comb[103:96]];
  assign p44_array_index_2051942_comb = p43_literal_2043896[p44_addedKey__50_comb[95:88]];
  assign p44_array_index_2051943_comb = p43_literal_2043896[p44_addedKey__50_comb[87:80]];
  assign p44_array_index_2051945_comb = p43_literal_2043896[p44_addedKey__50_comb[71:64]];
  assign p44_array_index_2051947_comb = p43_literal_2043896[p44_addedKey__50_comb[55:48]];
  assign p44_array_index_2051948_comb = p43_literal_2043896[p44_addedKey__50_comb[47:40]];
  assign p44_array_index_2051949_comb = p43_literal_2043896[p44_addedKey__50_comb[39:32]];
  assign p44_array_index_2051950_comb = p43_literal_2043896[p44_addedKey__50_comb[31:24]];
  assign p44_array_index_2051951_comb = p43_literal_2043896[p44_addedKey__50_comb[23:16]];
  assign p44_array_index_2051952_comb = p43_literal_2043896[p44_addedKey__50_comb[15:8]];
  assign p44_array_index_2051954_comb = p43_literal_2043910[p44_array_index_2051938_comb];
  assign p44_array_index_2051955_comb = p43_literal_2043912[p44_array_index_2051939_comb];
  assign p44_array_index_2051956_comb = p43_literal_2043914[p44_array_index_2051940_comb];
  assign p44_array_index_2051957_comb = p43_literal_2043916[p44_array_index_2051941_comb];
  assign p44_array_index_2051958_comb = p43_literal_2043918[p44_array_index_2051942_comb];
  assign p44_array_index_2051959_comb = p43_literal_2043920[p44_array_index_2051943_comb];
  assign p44_array_index_2051960_comb = p43_literal_2043896[p44_addedKey__50_comb[79:72]];
  assign p44_array_index_2051962_comb = p43_literal_2043896[p44_addedKey__50_comb[63:56]];
  assign p44_res7__576_comb = p44_array_index_2051954_comb ^ p44_array_index_2051955_comb ^ p44_array_index_2051956_comb ^ p44_array_index_2051957_comb ^ p44_array_index_2051958_comb ^ p44_array_index_2051959_comb ^ p44_array_index_2051960_comb ^ p43_literal_2043923[p44_array_index_2051945_comb] ^ p44_array_index_2051962_comb ^ p43_literal_2043920[p44_array_index_2051947_comb] ^ p43_literal_2043918[p44_array_index_2051948_comb] ^ p43_literal_2043916[p44_array_index_2051949_comb] ^ p43_literal_2043914[p44_array_index_2051950_comb] ^ p43_literal_2043912[p44_array_index_2051951_comb] ^ p43_literal_2043910[p44_array_index_2051952_comb] ^ p43_literal_2043896[p44_addedKey__50_comb[7:0]];

  // Registers for pipe stage 44:
  reg [127:0] p44_encoded;
  reg [127:0] p44_bit_slice_2043893;
  reg [127:0] p44_bit_slice_2044018;
  reg [127:0] p44_k3;
  reg [127:0] p44_k2;
  reg [127:0] p44_k5;
  reg [127:0] p44_k4;
  reg [127:0] p44_xor_2051482;
  reg [127:0] p44_xor_2051922;
  reg [7:0] p44_array_index_2051938;
  reg [7:0] p44_array_index_2051939;
  reg [7:0] p44_array_index_2051940;
  reg [7:0] p44_array_index_2051941;
  reg [7:0] p44_array_index_2051942;
  reg [7:0] p44_array_index_2051943;
  reg [7:0] p44_array_index_2051945;
  reg [7:0] p44_array_index_2051947;
  reg [7:0] p44_array_index_2051948;
  reg [7:0] p44_array_index_2051949;
  reg [7:0] p44_array_index_2051950;
  reg [7:0] p44_array_index_2051951;
  reg [7:0] p44_array_index_2051952;
  reg [7:0] p44_array_index_2051954;
  reg [7:0] p44_array_index_2051955;
  reg [7:0] p44_array_index_2051956;
  reg [7:0] p44_array_index_2051957;
  reg [7:0] p44_array_index_2051958;
  reg [7:0] p44_array_index_2051959;
  reg [7:0] p44_array_index_2051960;
  reg [7:0] p44_array_index_2051962;
  reg [7:0] p44_res7__576;
  reg [7:0] p45_literal_2043896[256];
  reg [7:0] p45_literal_2043910[256];
  reg [7:0] p45_literal_2043912[256];
  reg [7:0] p45_literal_2043914[256];
  reg [7:0] p45_literal_2043916[256];
  reg [7:0] p45_literal_2043918[256];
  reg [7:0] p45_literal_2043920[256];
  reg [7:0] p45_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p44_encoded <= p43_encoded;
    p44_bit_slice_2043893 <= p43_bit_slice_2043893;
    p44_bit_slice_2044018 <= p43_bit_slice_2044018;
    p44_k3 <= p43_k3;
    p44_k2 <= p43_k2;
    p44_k5 <= p43_k5;
    p44_k4 <= p43_k4;
    p44_xor_2051482 <= p43_xor_2051482;
    p44_xor_2051922 <= p44_xor_2051922_comb;
    p44_array_index_2051938 <= p44_array_index_2051938_comb;
    p44_array_index_2051939 <= p44_array_index_2051939_comb;
    p44_array_index_2051940 <= p44_array_index_2051940_comb;
    p44_array_index_2051941 <= p44_array_index_2051941_comb;
    p44_array_index_2051942 <= p44_array_index_2051942_comb;
    p44_array_index_2051943 <= p44_array_index_2051943_comb;
    p44_array_index_2051945 <= p44_array_index_2051945_comb;
    p44_array_index_2051947 <= p44_array_index_2051947_comb;
    p44_array_index_2051948 <= p44_array_index_2051948_comb;
    p44_array_index_2051949 <= p44_array_index_2051949_comb;
    p44_array_index_2051950 <= p44_array_index_2051950_comb;
    p44_array_index_2051951 <= p44_array_index_2051951_comb;
    p44_array_index_2051952 <= p44_array_index_2051952_comb;
    p44_array_index_2051954 <= p44_array_index_2051954_comb;
    p44_array_index_2051955 <= p44_array_index_2051955_comb;
    p44_array_index_2051956 <= p44_array_index_2051956_comb;
    p44_array_index_2051957 <= p44_array_index_2051957_comb;
    p44_array_index_2051958 <= p44_array_index_2051958_comb;
    p44_array_index_2051959 <= p44_array_index_2051959_comb;
    p44_array_index_2051960 <= p44_array_index_2051960_comb;
    p44_array_index_2051962 <= p44_array_index_2051962_comb;
    p44_res7__576 <= p44_res7__576_comb;
    p45_literal_2043896 <= p44_literal_2043896;
    p45_literal_2043910 <= p44_literal_2043910;
    p45_literal_2043912 <= p44_literal_2043912;
    p45_literal_2043914 <= p44_literal_2043914;
    p45_literal_2043916 <= p44_literal_2043916;
    p45_literal_2043918 <= p44_literal_2043918;
    p45_literal_2043920 <= p44_literal_2043920;
    p45_literal_2043923 <= p44_literal_2043923;
  end

  // ===== Pipe stage 45:
  wire [7:0] p45_array_index_2052049_comb;
  wire [7:0] p45_array_index_2052050_comb;
  wire [7:0] p45_array_index_2052051_comb;
  wire [7:0] p45_array_index_2052052_comb;
  wire [7:0] p45_array_index_2052053_comb;
  wire [7:0] p45_array_index_2052054_comb;
  wire [7:0] p45_res7__578_comb;
  wire [7:0] p45_array_index_2052064_comb;
  wire [7:0] p45_array_index_2052065_comb;
  wire [7:0] p45_array_index_2052066_comb;
  wire [7:0] p45_array_index_2052067_comb;
  wire [7:0] p45_array_index_2052068_comb;
  wire [7:0] p45_res7__580_comb;
  wire [7:0] p45_array_index_2052078_comb;
  wire [7:0] p45_array_index_2052079_comb;
  wire [7:0] p45_array_index_2052080_comb;
  wire [7:0] p45_array_index_2052081_comb;
  wire [7:0] p45_array_index_2052082_comb;
  wire [7:0] p45_res7__582_comb;
  wire [7:0] p45_array_index_2052093_comb;
  wire [7:0] p45_array_index_2052094_comb;
  wire [7:0] p45_array_index_2052095_comb;
  wire [7:0] p45_array_index_2052096_comb;
  wire [7:0] p45_res7__584_comb;
  wire [7:0] p45_array_index_2052106_comb;
  wire [7:0] p45_array_index_2052107_comb;
  wire [7:0] p45_array_index_2052108_comb;
  wire [7:0] p45_array_index_2052109_comb;
  wire [7:0] p45_res7__586_comb;
  wire [7:0] p45_array_index_2052120_comb;
  wire [7:0] p45_array_index_2052121_comb;
  wire [7:0] p45_array_index_2052122_comb;
  wire [7:0] p45_res7__588_comb;
  wire [7:0] p45_array_index_2052132_comb;
  wire [7:0] p45_array_index_2052133_comb;
  wire [7:0] p45_array_index_2052134_comb;
  wire [7:0] p45_res7__590_comb;
  assign p45_array_index_2052049_comb = p44_literal_2043910[p44_res7__576];
  assign p45_array_index_2052050_comb = p44_literal_2043912[p44_array_index_2051938];
  assign p45_array_index_2052051_comb = p44_literal_2043914[p44_array_index_2051939];
  assign p45_array_index_2052052_comb = p44_literal_2043916[p44_array_index_2051940];
  assign p45_array_index_2052053_comb = p44_literal_2043918[p44_array_index_2051941];
  assign p45_array_index_2052054_comb = p44_literal_2043920[p44_array_index_2051942];
  assign p45_res7__578_comb = p45_array_index_2052049_comb ^ p45_array_index_2052050_comb ^ p45_array_index_2052051_comb ^ p45_array_index_2052052_comb ^ p45_array_index_2052053_comb ^ p45_array_index_2052054_comb ^ p44_array_index_2051943 ^ p44_literal_2043923[p44_array_index_2051960] ^ p44_array_index_2051945 ^ p44_literal_2043920[p44_array_index_2051962] ^ p44_literal_2043918[p44_array_index_2051947] ^ p44_literal_2043916[p44_array_index_2051948] ^ p44_literal_2043914[p44_array_index_2051949] ^ p44_literal_2043912[p44_array_index_2051950] ^ p44_literal_2043910[p44_array_index_2051951] ^ p44_array_index_2051952;
  assign p45_array_index_2052064_comb = p44_literal_2043912[p44_res7__576];
  assign p45_array_index_2052065_comb = p44_literal_2043914[p44_array_index_2051938];
  assign p45_array_index_2052066_comb = p44_literal_2043916[p44_array_index_2051939];
  assign p45_array_index_2052067_comb = p44_literal_2043918[p44_array_index_2051940];
  assign p45_array_index_2052068_comb = p44_literal_2043920[p44_array_index_2051941];
  assign p45_res7__580_comb = p44_literal_2043910[p45_res7__578_comb] ^ p45_array_index_2052064_comb ^ p45_array_index_2052065_comb ^ p45_array_index_2052066_comb ^ p45_array_index_2052067_comb ^ p45_array_index_2052068_comb ^ p44_array_index_2051942 ^ p44_literal_2043923[p44_array_index_2051943] ^ p44_array_index_2051960 ^ p44_literal_2043920[p44_array_index_2051945] ^ p44_literal_2043918[p44_array_index_2051962] ^ p44_literal_2043916[p44_array_index_2051947] ^ p44_literal_2043914[p44_array_index_2051948] ^ p44_literal_2043912[p44_array_index_2051949] ^ p44_literal_2043910[p44_array_index_2051950] ^ p44_array_index_2051951;
  assign p45_array_index_2052078_comb = p44_literal_2043912[p45_res7__578_comb];
  assign p45_array_index_2052079_comb = p44_literal_2043914[p44_res7__576];
  assign p45_array_index_2052080_comb = p44_literal_2043916[p44_array_index_2051938];
  assign p45_array_index_2052081_comb = p44_literal_2043918[p44_array_index_2051939];
  assign p45_array_index_2052082_comb = p44_literal_2043920[p44_array_index_2051940];
  assign p45_res7__582_comb = p44_literal_2043910[p45_res7__580_comb] ^ p45_array_index_2052078_comb ^ p45_array_index_2052079_comb ^ p45_array_index_2052080_comb ^ p45_array_index_2052081_comb ^ p45_array_index_2052082_comb ^ p44_array_index_2051941 ^ p44_literal_2043923[p44_array_index_2051942] ^ p44_array_index_2051943 ^ p44_literal_2043920[p44_array_index_2051960] ^ p44_literal_2043918[p44_array_index_2051945] ^ p44_literal_2043916[p44_array_index_2051962] ^ p44_literal_2043914[p44_array_index_2051947] ^ p44_literal_2043912[p44_array_index_2051948] ^ p44_literal_2043910[p44_array_index_2051949] ^ p44_array_index_2051950;
  assign p45_array_index_2052093_comb = p44_literal_2043914[p45_res7__578_comb];
  assign p45_array_index_2052094_comb = p44_literal_2043916[p44_res7__576];
  assign p45_array_index_2052095_comb = p44_literal_2043918[p44_array_index_2051938];
  assign p45_array_index_2052096_comb = p44_literal_2043920[p44_array_index_2051939];
  assign p45_res7__584_comb = p44_literal_2043910[p45_res7__582_comb] ^ p44_literal_2043912[p45_res7__580_comb] ^ p45_array_index_2052093_comb ^ p45_array_index_2052094_comb ^ p45_array_index_2052095_comb ^ p45_array_index_2052096_comb ^ p44_array_index_2051940 ^ p44_literal_2043923[p44_array_index_2051941] ^ p44_array_index_2051942 ^ p44_array_index_2051959 ^ p44_literal_2043918[p44_array_index_2051960] ^ p44_literal_2043916[p44_array_index_2051945] ^ p44_literal_2043914[p44_array_index_2051962] ^ p44_literal_2043912[p44_array_index_2051947] ^ p44_literal_2043910[p44_array_index_2051948] ^ p44_array_index_2051949;
  assign p45_array_index_2052106_comb = p44_literal_2043914[p45_res7__580_comb];
  assign p45_array_index_2052107_comb = p44_literal_2043916[p45_res7__578_comb];
  assign p45_array_index_2052108_comb = p44_literal_2043918[p44_res7__576];
  assign p45_array_index_2052109_comb = p44_literal_2043920[p44_array_index_2051938];
  assign p45_res7__586_comb = p44_literal_2043910[p45_res7__584_comb] ^ p44_literal_2043912[p45_res7__582_comb] ^ p45_array_index_2052106_comb ^ p45_array_index_2052107_comb ^ p45_array_index_2052108_comb ^ p45_array_index_2052109_comb ^ p44_array_index_2051939 ^ p44_literal_2043923[p44_array_index_2051940] ^ p44_array_index_2051941 ^ p45_array_index_2052054_comb ^ p44_literal_2043918[p44_array_index_2051943] ^ p44_literal_2043916[p44_array_index_2051960] ^ p44_literal_2043914[p44_array_index_2051945] ^ p44_literal_2043912[p44_array_index_2051962] ^ p44_literal_2043910[p44_array_index_2051947] ^ p44_array_index_2051948;
  assign p45_array_index_2052120_comb = p44_literal_2043916[p45_res7__580_comb];
  assign p45_array_index_2052121_comb = p44_literal_2043918[p45_res7__578_comb];
  assign p45_array_index_2052122_comb = p44_literal_2043920[p44_res7__576];
  assign p45_res7__588_comb = p44_literal_2043910[p45_res7__586_comb] ^ p44_literal_2043912[p45_res7__584_comb] ^ p44_literal_2043914[p45_res7__582_comb] ^ p45_array_index_2052120_comb ^ p45_array_index_2052121_comb ^ p45_array_index_2052122_comb ^ p44_array_index_2051938 ^ p44_literal_2043923[p44_array_index_2051939] ^ p44_array_index_2051940 ^ p45_array_index_2052068_comb ^ p44_array_index_2051958 ^ p44_literal_2043916[p44_array_index_2051943] ^ p44_literal_2043914[p44_array_index_2051960] ^ p44_literal_2043912[p44_array_index_2051945] ^ p44_literal_2043910[p44_array_index_2051962] ^ p44_array_index_2051947;
  assign p45_array_index_2052132_comb = p44_literal_2043916[p45_res7__582_comb];
  assign p45_array_index_2052133_comb = p44_literal_2043918[p45_res7__580_comb];
  assign p45_array_index_2052134_comb = p44_literal_2043920[p45_res7__578_comb];
  assign p45_res7__590_comb = p44_literal_2043910[p45_res7__588_comb] ^ p44_literal_2043912[p45_res7__586_comb] ^ p44_literal_2043914[p45_res7__584_comb] ^ p45_array_index_2052132_comb ^ p45_array_index_2052133_comb ^ p45_array_index_2052134_comb ^ p44_res7__576 ^ p44_literal_2043923[p44_array_index_2051938] ^ p44_array_index_2051939 ^ p45_array_index_2052082_comb ^ p45_array_index_2052053_comb ^ p44_literal_2043916[p44_array_index_2051942] ^ p44_literal_2043914[p44_array_index_2051943] ^ p44_literal_2043912[p44_array_index_2051960] ^ p44_literal_2043910[p44_array_index_2051945] ^ p44_array_index_2051962;

  // Registers for pipe stage 45:
  reg [127:0] p45_encoded;
  reg [127:0] p45_bit_slice_2043893;
  reg [127:0] p45_bit_slice_2044018;
  reg [127:0] p45_k3;
  reg [127:0] p45_k2;
  reg [127:0] p45_k5;
  reg [127:0] p45_k4;
  reg [127:0] p45_xor_2051482;
  reg [127:0] p45_xor_2051922;
  reg [7:0] p45_array_index_2051938;
  reg [7:0] p45_array_index_2051939;
  reg [7:0] p45_array_index_2051940;
  reg [7:0] p45_array_index_2051941;
  reg [7:0] p45_array_index_2051942;
  reg [7:0] p45_array_index_2051943;
  reg [7:0] p45_array_index_2051945;
  reg [7:0] p45_array_index_2051954;
  reg [7:0] p45_array_index_2051955;
  reg [7:0] p45_array_index_2051956;
  reg [7:0] p45_array_index_2051957;
  reg [7:0] p45_array_index_2051960;
  reg [7:0] p45_res7__576;
  reg [7:0] p45_array_index_2052049;
  reg [7:0] p45_array_index_2052050;
  reg [7:0] p45_array_index_2052051;
  reg [7:0] p45_array_index_2052052;
  reg [7:0] p45_res7__578;
  reg [7:0] p45_array_index_2052064;
  reg [7:0] p45_array_index_2052065;
  reg [7:0] p45_array_index_2052066;
  reg [7:0] p45_array_index_2052067;
  reg [7:0] p45_res7__580;
  reg [7:0] p45_array_index_2052078;
  reg [7:0] p45_array_index_2052079;
  reg [7:0] p45_array_index_2052080;
  reg [7:0] p45_array_index_2052081;
  reg [7:0] p45_res7__582;
  reg [7:0] p45_array_index_2052093;
  reg [7:0] p45_array_index_2052094;
  reg [7:0] p45_array_index_2052095;
  reg [7:0] p45_array_index_2052096;
  reg [7:0] p45_res7__584;
  reg [7:0] p45_array_index_2052106;
  reg [7:0] p45_array_index_2052107;
  reg [7:0] p45_array_index_2052108;
  reg [7:0] p45_array_index_2052109;
  reg [7:0] p45_res7__586;
  reg [7:0] p45_array_index_2052120;
  reg [7:0] p45_array_index_2052121;
  reg [7:0] p45_array_index_2052122;
  reg [7:0] p45_res7__588;
  reg [7:0] p45_array_index_2052132;
  reg [7:0] p45_array_index_2052133;
  reg [7:0] p45_array_index_2052134;
  reg [7:0] p45_res7__590;
  reg [7:0] p46_literal_2043896[256];
  reg [7:0] p46_literal_2043910[256];
  reg [7:0] p46_literal_2043912[256];
  reg [7:0] p46_literal_2043914[256];
  reg [7:0] p46_literal_2043916[256];
  reg [7:0] p46_literal_2043918[256];
  reg [7:0] p46_literal_2043920[256];
  reg [7:0] p46_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p45_encoded <= p44_encoded;
    p45_bit_slice_2043893 <= p44_bit_slice_2043893;
    p45_bit_slice_2044018 <= p44_bit_slice_2044018;
    p45_k3 <= p44_k3;
    p45_k2 <= p44_k2;
    p45_k5 <= p44_k5;
    p45_k4 <= p44_k4;
    p45_xor_2051482 <= p44_xor_2051482;
    p45_xor_2051922 <= p44_xor_2051922;
    p45_array_index_2051938 <= p44_array_index_2051938;
    p45_array_index_2051939 <= p44_array_index_2051939;
    p45_array_index_2051940 <= p44_array_index_2051940;
    p45_array_index_2051941 <= p44_array_index_2051941;
    p45_array_index_2051942 <= p44_array_index_2051942;
    p45_array_index_2051943 <= p44_array_index_2051943;
    p45_array_index_2051945 <= p44_array_index_2051945;
    p45_array_index_2051954 <= p44_array_index_2051954;
    p45_array_index_2051955 <= p44_array_index_2051955;
    p45_array_index_2051956 <= p44_array_index_2051956;
    p45_array_index_2051957 <= p44_array_index_2051957;
    p45_array_index_2051960 <= p44_array_index_2051960;
    p45_res7__576 <= p44_res7__576;
    p45_array_index_2052049 <= p45_array_index_2052049_comb;
    p45_array_index_2052050 <= p45_array_index_2052050_comb;
    p45_array_index_2052051 <= p45_array_index_2052051_comb;
    p45_array_index_2052052 <= p45_array_index_2052052_comb;
    p45_res7__578 <= p45_res7__578_comb;
    p45_array_index_2052064 <= p45_array_index_2052064_comb;
    p45_array_index_2052065 <= p45_array_index_2052065_comb;
    p45_array_index_2052066 <= p45_array_index_2052066_comb;
    p45_array_index_2052067 <= p45_array_index_2052067_comb;
    p45_res7__580 <= p45_res7__580_comb;
    p45_array_index_2052078 <= p45_array_index_2052078_comb;
    p45_array_index_2052079 <= p45_array_index_2052079_comb;
    p45_array_index_2052080 <= p45_array_index_2052080_comb;
    p45_array_index_2052081 <= p45_array_index_2052081_comb;
    p45_res7__582 <= p45_res7__582_comb;
    p45_array_index_2052093 <= p45_array_index_2052093_comb;
    p45_array_index_2052094 <= p45_array_index_2052094_comb;
    p45_array_index_2052095 <= p45_array_index_2052095_comb;
    p45_array_index_2052096 <= p45_array_index_2052096_comb;
    p45_res7__584 <= p45_res7__584_comb;
    p45_array_index_2052106 <= p45_array_index_2052106_comb;
    p45_array_index_2052107 <= p45_array_index_2052107_comb;
    p45_array_index_2052108 <= p45_array_index_2052108_comb;
    p45_array_index_2052109 <= p45_array_index_2052109_comb;
    p45_res7__586 <= p45_res7__586_comb;
    p45_array_index_2052120 <= p45_array_index_2052120_comb;
    p45_array_index_2052121 <= p45_array_index_2052121_comb;
    p45_array_index_2052122 <= p45_array_index_2052122_comb;
    p45_res7__588 <= p45_res7__588_comb;
    p45_array_index_2052132 <= p45_array_index_2052132_comb;
    p45_array_index_2052133 <= p45_array_index_2052133_comb;
    p45_array_index_2052134 <= p45_array_index_2052134_comb;
    p45_res7__590 <= p45_res7__590_comb;
    p46_literal_2043896 <= p45_literal_2043896;
    p46_literal_2043910 <= p45_literal_2043910;
    p46_literal_2043912 <= p45_literal_2043912;
    p46_literal_2043914 <= p45_literal_2043914;
    p46_literal_2043916 <= p45_literal_2043916;
    p46_literal_2043918 <= p45_literal_2043918;
    p46_literal_2043920 <= p45_literal_2043920;
    p46_literal_2043923 <= p45_literal_2043923;
  end

  // ===== Pipe stage 46:
  wire [7:0] p46_array_index_2052271_comb;
  wire [7:0] p46_array_index_2052272_comb;
  wire [7:0] p46_res7__592_comb;
  wire [7:0] p46_array_index_2052282_comb;
  wire [7:0] p46_array_index_2052283_comb;
  wire [7:0] p46_res7__594_comb;
  wire [7:0] p46_array_index_2052294_comb;
  wire [7:0] p46_res7__596_comb;
  wire [7:0] p46_array_index_2052304_comb;
  wire [7:0] p46_res7__598_comb;
  wire [7:0] p46_res7__600_comb;
  wire [7:0] p46_res7__602_comb;
  wire [7:0] p46_res7__604_comb;
  assign p46_array_index_2052271_comb = p45_literal_2043918[p45_res7__582];
  assign p46_array_index_2052272_comb = p45_literal_2043920[p45_res7__580];
  assign p46_res7__592_comb = p45_literal_2043910[p45_res7__590] ^ p45_literal_2043912[p45_res7__588] ^ p45_literal_2043914[p45_res7__586] ^ p45_literal_2043916[p45_res7__584] ^ p46_array_index_2052271_comb ^ p46_array_index_2052272_comb ^ p45_res7__578 ^ p45_literal_2043923[p45_res7__576] ^ p45_array_index_2051938 ^ p45_array_index_2052096 ^ p45_array_index_2052067 ^ p45_array_index_2051957 ^ p45_literal_2043914[p45_array_index_2051942] ^ p45_literal_2043912[p45_array_index_2051943] ^ p45_literal_2043910[p45_array_index_2051960] ^ p45_array_index_2051945;
  assign p46_array_index_2052282_comb = p45_literal_2043918[p45_res7__584];
  assign p46_array_index_2052283_comb = p45_literal_2043920[p45_res7__582];
  assign p46_res7__594_comb = p45_literal_2043910[p46_res7__592_comb] ^ p45_literal_2043912[p45_res7__590] ^ p45_literal_2043914[p45_res7__588] ^ p45_literal_2043916[p45_res7__586] ^ p46_array_index_2052282_comb ^ p46_array_index_2052283_comb ^ p45_res7__580 ^ p45_literal_2043923[p45_res7__578] ^ p45_res7__576 ^ p45_array_index_2052109 ^ p45_array_index_2052081 ^ p45_array_index_2052052 ^ p45_literal_2043914[p45_array_index_2051941] ^ p45_literal_2043912[p45_array_index_2051942] ^ p45_literal_2043910[p45_array_index_2051943] ^ p45_array_index_2051960;
  assign p46_array_index_2052294_comb = p45_literal_2043920[p45_res7__584];
  assign p46_res7__596_comb = p45_literal_2043910[p46_res7__594_comb] ^ p45_literal_2043912[p46_res7__592_comb] ^ p45_literal_2043914[p45_res7__590] ^ p45_literal_2043916[p45_res7__588] ^ p45_literal_2043918[p45_res7__586] ^ p46_array_index_2052294_comb ^ p45_res7__582 ^ p45_literal_2043923[p45_res7__580] ^ p45_res7__578 ^ p45_array_index_2052122 ^ p45_array_index_2052095 ^ p45_array_index_2052066 ^ p45_array_index_2051956 ^ p45_literal_2043912[p45_array_index_2051941] ^ p45_literal_2043910[p45_array_index_2051942] ^ p45_array_index_2051943;
  assign p46_array_index_2052304_comb = p45_literal_2043920[p45_res7__586];
  assign p46_res7__598_comb = p45_literal_2043910[p46_res7__596_comb] ^ p45_literal_2043912[p46_res7__594_comb] ^ p45_literal_2043914[p46_res7__592_comb] ^ p45_literal_2043916[p45_res7__590] ^ p45_literal_2043918[p45_res7__588] ^ p46_array_index_2052304_comb ^ p45_res7__584 ^ p45_literal_2043923[p45_res7__582] ^ p45_res7__580 ^ p45_array_index_2052134 ^ p45_array_index_2052108 ^ p45_array_index_2052080 ^ p45_array_index_2052051 ^ p45_literal_2043912[p45_array_index_2051940] ^ p45_literal_2043910[p45_array_index_2051941] ^ p45_array_index_2051942;
  assign p46_res7__600_comb = p45_literal_2043910[p46_res7__598_comb] ^ p45_literal_2043912[p46_res7__596_comb] ^ p45_literal_2043914[p46_res7__594_comb] ^ p45_literal_2043916[p46_res7__592_comb] ^ p45_literal_2043918[p45_res7__590] ^ p45_literal_2043920[p45_res7__588] ^ p45_res7__586 ^ p45_literal_2043923[p45_res7__584] ^ p45_res7__582 ^ p46_array_index_2052272_comb ^ p45_array_index_2052121 ^ p45_array_index_2052094 ^ p45_array_index_2052065 ^ p45_array_index_2051955 ^ p45_literal_2043910[p45_array_index_2051940] ^ p45_array_index_2051941;
  assign p46_res7__602_comb = p45_literal_2043910[p46_res7__600_comb] ^ p45_literal_2043912[p46_res7__598_comb] ^ p45_literal_2043914[p46_res7__596_comb] ^ p45_literal_2043916[p46_res7__594_comb] ^ p45_literal_2043918[p46_res7__592_comb] ^ p45_literal_2043920[p45_res7__590] ^ p45_res7__588 ^ p45_literal_2043923[p45_res7__586] ^ p45_res7__584 ^ p46_array_index_2052283_comb ^ p45_array_index_2052133 ^ p45_array_index_2052107 ^ p45_array_index_2052079 ^ p45_array_index_2052050 ^ p45_literal_2043910[p45_array_index_2051939] ^ p45_array_index_2051940;
  assign p46_res7__604_comb = p45_literal_2043910[p46_res7__602_comb] ^ p45_literal_2043912[p46_res7__600_comb] ^ p45_literal_2043914[p46_res7__598_comb] ^ p45_literal_2043916[p46_res7__596_comb] ^ p45_literal_2043918[p46_res7__594_comb] ^ p45_literal_2043920[p46_res7__592_comb] ^ p45_res7__590 ^ p45_literal_2043923[p45_res7__588] ^ p45_res7__586 ^ p46_array_index_2052294_comb ^ p46_array_index_2052271_comb ^ p45_array_index_2052120 ^ p45_array_index_2052093 ^ p45_array_index_2052064 ^ p45_array_index_2051954 ^ p45_array_index_2051939;

  // Registers for pipe stage 46:
  reg [127:0] p46_encoded;
  reg [127:0] p46_bit_slice_2043893;
  reg [127:0] p46_bit_slice_2044018;
  reg [127:0] p46_k3;
  reg [127:0] p46_k2;
  reg [127:0] p46_k5;
  reg [127:0] p46_k4;
  reg [127:0] p46_xor_2051482;
  reg [127:0] p46_xor_2051922;
  reg [7:0] p46_array_index_2051938;
  reg [7:0] p46_res7__576;
  reg [7:0] p46_array_index_2052049;
  reg [7:0] p46_res7__578;
  reg [7:0] p46_res7__580;
  reg [7:0] p46_array_index_2052078;
  reg [7:0] p46_res7__582;
  reg [7:0] p46_res7__584;
  reg [7:0] p46_array_index_2052106;
  reg [7:0] p46_res7__586;
  reg [7:0] p46_res7__588;
  reg [7:0] p46_array_index_2052132;
  reg [7:0] p46_res7__590;
  reg [7:0] p46_res7__592;
  reg [7:0] p46_array_index_2052282;
  reg [7:0] p46_res7__594;
  reg [7:0] p46_res7__596;
  reg [7:0] p46_array_index_2052304;
  reg [7:0] p46_res7__598;
  reg [7:0] p46_res7__600;
  reg [7:0] p46_res7__602;
  reg [7:0] p46_res7__604;
  reg [7:0] p47_literal_2043896[256];
  reg [7:0] p47_literal_2043910[256];
  reg [7:0] p47_literal_2043912[256];
  reg [7:0] p47_literal_2043914[256];
  reg [7:0] p47_literal_2043916[256];
  reg [7:0] p47_literal_2043918[256];
  reg [7:0] p47_literal_2043920[256];
  reg [7:0] p47_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p46_encoded <= p45_encoded;
    p46_bit_slice_2043893 <= p45_bit_slice_2043893;
    p46_bit_slice_2044018 <= p45_bit_slice_2044018;
    p46_k3 <= p45_k3;
    p46_k2 <= p45_k2;
    p46_k5 <= p45_k5;
    p46_k4 <= p45_k4;
    p46_xor_2051482 <= p45_xor_2051482;
    p46_xor_2051922 <= p45_xor_2051922;
    p46_array_index_2051938 <= p45_array_index_2051938;
    p46_res7__576 <= p45_res7__576;
    p46_array_index_2052049 <= p45_array_index_2052049;
    p46_res7__578 <= p45_res7__578;
    p46_res7__580 <= p45_res7__580;
    p46_array_index_2052078 <= p45_array_index_2052078;
    p46_res7__582 <= p45_res7__582;
    p46_res7__584 <= p45_res7__584;
    p46_array_index_2052106 <= p45_array_index_2052106;
    p46_res7__586 <= p45_res7__586;
    p46_res7__588 <= p45_res7__588;
    p46_array_index_2052132 <= p45_array_index_2052132;
    p46_res7__590 <= p45_res7__590;
    p46_res7__592 <= p46_res7__592_comb;
    p46_array_index_2052282 <= p46_array_index_2052282_comb;
    p46_res7__594 <= p46_res7__594_comb;
    p46_res7__596 <= p46_res7__596_comb;
    p46_array_index_2052304 <= p46_array_index_2052304_comb;
    p46_res7__598 <= p46_res7__598_comb;
    p46_res7__600 <= p46_res7__600_comb;
    p46_res7__602 <= p46_res7__602_comb;
    p46_res7__604 <= p46_res7__604_comb;
    p47_literal_2043896 <= p46_literal_2043896;
    p47_literal_2043910 <= p46_literal_2043910;
    p47_literal_2043912 <= p46_literal_2043912;
    p47_literal_2043914 <= p46_literal_2043914;
    p47_literal_2043916 <= p46_literal_2043916;
    p47_literal_2043918 <= p46_literal_2043918;
    p47_literal_2043920 <= p46_literal_2043920;
    p47_literal_2043923 <= p46_literal_2043923;
  end

  // ===== Pipe stage 47:
  wire [7:0] p47_res7__606_comb;
  wire [127:0] p47_res__18_comb;
  wire [127:0] p47_xor_2052422_comb;
  wire [127:0] p47_addedKey__51_comb;
  wire [7:0] p47_array_index_2052438_comb;
  wire [7:0] p47_array_index_2052439_comb;
  wire [7:0] p47_array_index_2052440_comb;
  wire [7:0] p47_array_index_2052441_comb;
  wire [7:0] p47_array_index_2052442_comb;
  wire [7:0] p47_array_index_2052443_comb;
  wire [7:0] p47_array_index_2052445_comb;
  wire [7:0] p47_array_index_2052447_comb;
  wire [7:0] p47_array_index_2052448_comb;
  wire [7:0] p47_array_index_2052449_comb;
  wire [7:0] p47_array_index_2052450_comb;
  wire [7:0] p47_array_index_2052451_comb;
  wire [7:0] p47_array_index_2052452_comb;
  wire [7:0] p47_array_index_2052454_comb;
  wire [7:0] p47_array_index_2052455_comb;
  wire [7:0] p47_array_index_2052456_comb;
  wire [7:0] p47_array_index_2052457_comb;
  wire [7:0] p47_array_index_2052458_comb;
  wire [7:0] p47_array_index_2052459_comb;
  wire [7:0] p47_array_index_2052460_comb;
  wire [7:0] p47_array_index_2052462_comb;
  wire [7:0] p47_res7__608_comb;
  wire [7:0] p47_array_index_2052471_comb;
  wire [7:0] p47_array_index_2052472_comb;
  wire [7:0] p47_array_index_2052473_comb;
  wire [7:0] p47_array_index_2052474_comb;
  wire [7:0] p47_array_index_2052475_comb;
  wire [7:0] p47_array_index_2052476_comb;
  wire [7:0] p47_res7__610_comb;
  wire [7:0] p47_array_index_2052486_comb;
  wire [7:0] p47_array_index_2052487_comb;
  wire [7:0] p47_array_index_2052488_comb;
  wire [7:0] p47_array_index_2052489_comb;
  wire [7:0] p47_array_index_2052490_comb;
  wire [7:0] p47_res7__612_comb;
  wire [7:0] p47_array_index_2052500_comb;
  wire [7:0] p47_array_index_2052501_comb;
  wire [7:0] p47_array_index_2052502_comb;
  wire [7:0] p47_array_index_2052503_comb;
  wire [7:0] p47_array_index_2052504_comb;
  wire [7:0] p47_res7__614_comb;
  wire [7:0] p47_array_index_2052515_comb;
  wire [7:0] p47_array_index_2052516_comb;
  wire [7:0] p47_array_index_2052517_comb;
  wire [7:0] p47_array_index_2052518_comb;
  wire [7:0] p47_res7__616_comb;
  assign p47_res7__606_comb = p46_literal_2043910[p46_res7__604] ^ p46_literal_2043912[p46_res7__602] ^ p46_literal_2043914[p46_res7__600] ^ p46_literal_2043916[p46_res7__598] ^ p46_literal_2043918[p46_res7__596] ^ p46_literal_2043920[p46_res7__594] ^ p46_res7__592 ^ p46_literal_2043923[p46_res7__590] ^ p46_res7__588 ^ p46_array_index_2052304 ^ p46_array_index_2052282 ^ p46_array_index_2052132 ^ p46_array_index_2052106 ^ p46_array_index_2052078 ^ p46_array_index_2052049 ^ p46_array_index_2051938;
  assign p47_res__18_comb = {p47_res7__606_comb, p46_res7__604, p46_res7__602, p46_res7__600, p46_res7__598, p46_res7__596, p46_res7__594, p46_res7__592, p46_res7__590, p46_res7__588, p46_res7__586, p46_res7__584, p46_res7__582, p46_res7__580, p46_res7__578, p46_res7__576};
  assign p47_xor_2052422_comb = p47_res__18_comb ^ p46_xor_2051482;
  assign p47_addedKey__51_comb = p47_xor_2052422_comb ^ 128'h547f_7727_7ce9_8774_2ea9_3083_bcc2_4114;
  assign p47_array_index_2052438_comb = p46_literal_2043896[p47_addedKey__51_comb[127:120]];
  assign p47_array_index_2052439_comb = p46_literal_2043896[p47_addedKey__51_comb[119:112]];
  assign p47_array_index_2052440_comb = p46_literal_2043896[p47_addedKey__51_comb[111:104]];
  assign p47_array_index_2052441_comb = p46_literal_2043896[p47_addedKey__51_comb[103:96]];
  assign p47_array_index_2052442_comb = p46_literal_2043896[p47_addedKey__51_comb[95:88]];
  assign p47_array_index_2052443_comb = p46_literal_2043896[p47_addedKey__51_comb[87:80]];
  assign p47_array_index_2052445_comb = p46_literal_2043896[p47_addedKey__51_comb[71:64]];
  assign p47_array_index_2052447_comb = p46_literal_2043896[p47_addedKey__51_comb[55:48]];
  assign p47_array_index_2052448_comb = p46_literal_2043896[p47_addedKey__51_comb[47:40]];
  assign p47_array_index_2052449_comb = p46_literal_2043896[p47_addedKey__51_comb[39:32]];
  assign p47_array_index_2052450_comb = p46_literal_2043896[p47_addedKey__51_comb[31:24]];
  assign p47_array_index_2052451_comb = p46_literal_2043896[p47_addedKey__51_comb[23:16]];
  assign p47_array_index_2052452_comb = p46_literal_2043896[p47_addedKey__51_comb[15:8]];
  assign p47_array_index_2052454_comb = p46_literal_2043910[p47_array_index_2052438_comb];
  assign p47_array_index_2052455_comb = p46_literal_2043912[p47_array_index_2052439_comb];
  assign p47_array_index_2052456_comb = p46_literal_2043914[p47_array_index_2052440_comb];
  assign p47_array_index_2052457_comb = p46_literal_2043916[p47_array_index_2052441_comb];
  assign p47_array_index_2052458_comb = p46_literal_2043918[p47_array_index_2052442_comb];
  assign p47_array_index_2052459_comb = p46_literal_2043920[p47_array_index_2052443_comb];
  assign p47_array_index_2052460_comb = p46_literal_2043896[p47_addedKey__51_comb[79:72]];
  assign p47_array_index_2052462_comb = p46_literal_2043896[p47_addedKey__51_comb[63:56]];
  assign p47_res7__608_comb = p47_array_index_2052454_comb ^ p47_array_index_2052455_comb ^ p47_array_index_2052456_comb ^ p47_array_index_2052457_comb ^ p47_array_index_2052458_comb ^ p47_array_index_2052459_comb ^ p47_array_index_2052460_comb ^ p46_literal_2043923[p47_array_index_2052445_comb] ^ p47_array_index_2052462_comb ^ p46_literal_2043920[p47_array_index_2052447_comb] ^ p46_literal_2043918[p47_array_index_2052448_comb] ^ p46_literal_2043916[p47_array_index_2052449_comb] ^ p46_literal_2043914[p47_array_index_2052450_comb] ^ p46_literal_2043912[p47_array_index_2052451_comb] ^ p46_literal_2043910[p47_array_index_2052452_comb] ^ p46_literal_2043896[p47_addedKey__51_comb[7:0]];
  assign p47_array_index_2052471_comb = p46_literal_2043910[p47_res7__608_comb];
  assign p47_array_index_2052472_comb = p46_literal_2043912[p47_array_index_2052438_comb];
  assign p47_array_index_2052473_comb = p46_literal_2043914[p47_array_index_2052439_comb];
  assign p47_array_index_2052474_comb = p46_literal_2043916[p47_array_index_2052440_comb];
  assign p47_array_index_2052475_comb = p46_literal_2043918[p47_array_index_2052441_comb];
  assign p47_array_index_2052476_comb = p46_literal_2043920[p47_array_index_2052442_comb];
  assign p47_res7__610_comb = p47_array_index_2052471_comb ^ p47_array_index_2052472_comb ^ p47_array_index_2052473_comb ^ p47_array_index_2052474_comb ^ p47_array_index_2052475_comb ^ p47_array_index_2052476_comb ^ p47_array_index_2052443_comb ^ p46_literal_2043923[p47_array_index_2052460_comb] ^ p47_array_index_2052445_comb ^ p46_literal_2043920[p47_array_index_2052462_comb] ^ p46_literal_2043918[p47_array_index_2052447_comb] ^ p46_literal_2043916[p47_array_index_2052448_comb] ^ p46_literal_2043914[p47_array_index_2052449_comb] ^ p46_literal_2043912[p47_array_index_2052450_comb] ^ p46_literal_2043910[p47_array_index_2052451_comb] ^ p47_array_index_2052452_comb;
  assign p47_array_index_2052486_comb = p46_literal_2043912[p47_res7__608_comb];
  assign p47_array_index_2052487_comb = p46_literal_2043914[p47_array_index_2052438_comb];
  assign p47_array_index_2052488_comb = p46_literal_2043916[p47_array_index_2052439_comb];
  assign p47_array_index_2052489_comb = p46_literal_2043918[p47_array_index_2052440_comb];
  assign p47_array_index_2052490_comb = p46_literal_2043920[p47_array_index_2052441_comb];
  assign p47_res7__612_comb = p46_literal_2043910[p47_res7__610_comb] ^ p47_array_index_2052486_comb ^ p47_array_index_2052487_comb ^ p47_array_index_2052488_comb ^ p47_array_index_2052489_comb ^ p47_array_index_2052490_comb ^ p47_array_index_2052442_comb ^ p46_literal_2043923[p47_array_index_2052443_comb] ^ p47_array_index_2052460_comb ^ p46_literal_2043920[p47_array_index_2052445_comb] ^ p46_literal_2043918[p47_array_index_2052462_comb] ^ p46_literal_2043916[p47_array_index_2052447_comb] ^ p46_literal_2043914[p47_array_index_2052448_comb] ^ p46_literal_2043912[p47_array_index_2052449_comb] ^ p46_literal_2043910[p47_array_index_2052450_comb] ^ p47_array_index_2052451_comb;
  assign p47_array_index_2052500_comb = p46_literal_2043912[p47_res7__610_comb];
  assign p47_array_index_2052501_comb = p46_literal_2043914[p47_res7__608_comb];
  assign p47_array_index_2052502_comb = p46_literal_2043916[p47_array_index_2052438_comb];
  assign p47_array_index_2052503_comb = p46_literal_2043918[p47_array_index_2052439_comb];
  assign p47_array_index_2052504_comb = p46_literal_2043920[p47_array_index_2052440_comb];
  assign p47_res7__614_comb = p46_literal_2043910[p47_res7__612_comb] ^ p47_array_index_2052500_comb ^ p47_array_index_2052501_comb ^ p47_array_index_2052502_comb ^ p47_array_index_2052503_comb ^ p47_array_index_2052504_comb ^ p47_array_index_2052441_comb ^ p46_literal_2043923[p47_array_index_2052442_comb] ^ p47_array_index_2052443_comb ^ p46_literal_2043920[p47_array_index_2052460_comb] ^ p46_literal_2043918[p47_array_index_2052445_comb] ^ p46_literal_2043916[p47_array_index_2052462_comb] ^ p46_literal_2043914[p47_array_index_2052447_comb] ^ p46_literal_2043912[p47_array_index_2052448_comb] ^ p46_literal_2043910[p47_array_index_2052449_comb] ^ p47_array_index_2052450_comb;
  assign p47_array_index_2052515_comb = p46_literal_2043914[p47_res7__610_comb];
  assign p47_array_index_2052516_comb = p46_literal_2043916[p47_res7__608_comb];
  assign p47_array_index_2052517_comb = p46_literal_2043918[p47_array_index_2052438_comb];
  assign p47_array_index_2052518_comb = p46_literal_2043920[p47_array_index_2052439_comb];
  assign p47_res7__616_comb = p46_literal_2043910[p47_res7__614_comb] ^ p46_literal_2043912[p47_res7__612_comb] ^ p47_array_index_2052515_comb ^ p47_array_index_2052516_comb ^ p47_array_index_2052517_comb ^ p47_array_index_2052518_comb ^ p47_array_index_2052440_comb ^ p46_literal_2043923[p47_array_index_2052441_comb] ^ p47_array_index_2052442_comb ^ p47_array_index_2052459_comb ^ p46_literal_2043918[p47_array_index_2052460_comb] ^ p46_literal_2043916[p47_array_index_2052445_comb] ^ p46_literal_2043914[p47_array_index_2052462_comb] ^ p46_literal_2043912[p47_array_index_2052447_comb] ^ p46_literal_2043910[p47_array_index_2052448_comb] ^ p47_array_index_2052449_comb;

  // Registers for pipe stage 47:
  reg [127:0] p47_encoded;
  reg [127:0] p47_bit_slice_2043893;
  reg [127:0] p47_bit_slice_2044018;
  reg [127:0] p47_k3;
  reg [127:0] p47_k2;
  reg [127:0] p47_k5;
  reg [127:0] p47_k4;
  reg [127:0] p47_xor_2051922;
  reg [127:0] p47_xor_2052422;
  reg [7:0] p47_array_index_2052438;
  reg [7:0] p47_array_index_2052439;
  reg [7:0] p47_array_index_2052440;
  reg [7:0] p47_array_index_2052441;
  reg [7:0] p47_array_index_2052442;
  reg [7:0] p47_array_index_2052443;
  reg [7:0] p47_array_index_2052445;
  reg [7:0] p47_array_index_2052447;
  reg [7:0] p47_array_index_2052448;
  reg [7:0] p47_array_index_2052454;
  reg [7:0] p47_array_index_2052455;
  reg [7:0] p47_array_index_2052456;
  reg [7:0] p47_array_index_2052457;
  reg [7:0] p47_array_index_2052458;
  reg [7:0] p47_array_index_2052460;
  reg [7:0] p47_array_index_2052462;
  reg [7:0] p47_res7__608;
  reg [7:0] p47_array_index_2052471;
  reg [7:0] p47_array_index_2052472;
  reg [7:0] p47_array_index_2052473;
  reg [7:0] p47_array_index_2052474;
  reg [7:0] p47_array_index_2052475;
  reg [7:0] p47_array_index_2052476;
  reg [7:0] p47_res7__610;
  reg [7:0] p47_array_index_2052486;
  reg [7:0] p47_array_index_2052487;
  reg [7:0] p47_array_index_2052488;
  reg [7:0] p47_array_index_2052489;
  reg [7:0] p47_array_index_2052490;
  reg [7:0] p47_res7__612;
  reg [7:0] p47_array_index_2052500;
  reg [7:0] p47_array_index_2052501;
  reg [7:0] p47_array_index_2052502;
  reg [7:0] p47_array_index_2052503;
  reg [7:0] p47_array_index_2052504;
  reg [7:0] p47_res7__614;
  reg [7:0] p47_array_index_2052515;
  reg [7:0] p47_array_index_2052516;
  reg [7:0] p47_array_index_2052517;
  reg [7:0] p47_array_index_2052518;
  reg [7:0] p47_res7__616;
  reg [7:0] p48_literal_2043896[256];
  reg [7:0] p48_literal_2043910[256];
  reg [7:0] p48_literal_2043912[256];
  reg [7:0] p48_literal_2043914[256];
  reg [7:0] p48_literal_2043916[256];
  reg [7:0] p48_literal_2043918[256];
  reg [7:0] p48_literal_2043920[256];
  reg [7:0] p48_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p47_encoded <= p46_encoded;
    p47_bit_slice_2043893 <= p46_bit_slice_2043893;
    p47_bit_slice_2044018 <= p46_bit_slice_2044018;
    p47_k3 <= p46_k3;
    p47_k2 <= p46_k2;
    p47_k5 <= p46_k5;
    p47_k4 <= p46_k4;
    p47_xor_2051922 <= p46_xor_2051922;
    p47_xor_2052422 <= p47_xor_2052422_comb;
    p47_array_index_2052438 <= p47_array_index_2052438_comb;
    p47_array_index_2052439 <= p47_array_index_2052439_comb;
    p47_array_index_2052440 <= p47_array_index_2052440_comb;
    p47_array_index_2052441 <= p47_array_index_2052441_comb;
    p47_array_index_2052442 <= p47_array_index_2052442_comb;
    p47_array_index_2052443 <= p47_array_index_2052443_comb;
    p47_array_index_2052445 <= p47_array_index_2052445_comb;
    p47_array_index_2052447 <= p47_array_index_2052447_comb;
    p47_array_index_2052448 <= p47_array_index_2052448_comb;
    p47_array_index_2052454 <= p47_array_index_2052454_comb;
    p47_array_index_2052455 <= p47_array_index_2052455_comb;
    p47_array_index_2052456 <= p47_array_index_2052456_comb;
    p47_array_index_2052457 <= p47_array_index_2052457_comb;
    p47_array_index_2052458 <= p47_array_index_2052458_comb;
    p47_array_index_2052460 <= p47_array_index_2052460_comb;
    p47_array_index_2052462 <= p47_array_index_2052462_comb;
    p47_res7__608 <= p47_res7__608_comb;
    p47_array_index_2052471 <= p47_array_index_2052471_comb;
    p47_array_index_2052472 <= p47_array_index_2052472_comb;
    p47_array_index_2052473 <= p47_array_index_2052473_comb;
    p47_array_index_2052474 <= p47_array_index_2052474_comb;
    p47_array_index_2052475 <= p47_array_index_2052475_comb;
    p47_array_index_2052476 <= p47_array_index_2052476_comb;
    p47_res7__610 <= p47_res7__610_comb;
    p47_array_index_2052486 <= p47_array_index_2052486_comb;
    p47_array_index_2052487 <= p47_array_index_2052487_comb;
    p47_array_index_2052488 <= p47_array_index_2052488_comb;
    p47_array_index_2052489 <= p47_array_index_2052489_comb;
    p47_array_index_2052490 <= p47_array_index_2052490_comb;
    p47_res7__612 <= p47_res7__612_comb;
    p47_array_index_2052500 <= p47_array_index_2052500_comb;
    p47_array_index_2052501 <= p47_array_index_2052501_comb;
    p47_array_index_2052502 <= p47_array_index_2052502_comb;
    p47_array_index_2052503 <= p47_array_index_2052503_comb;
    p47_array_index_2052504 <= p47_array_index_2052504_comb;
    p47_res7__614 <= p47_res7__614_comb;
    p47_array_index_2052515 <= p47_array_index_2052515_comb;
    p47_array_index_2052516 <= p47_array_index_2052516_comb;
    p47_array_index_2052517 <= p47_array_index_2052517_comb;
    p47_array_index_2052518 <= p47_array_index_2052518_comb;
    p47_res7__616 <= p47_res7__616_comb;
    p48_literal_2043896 <= p47_literal_2043896;
    p48_literal_2043910 <= p47_literal_2043910;
    p48_literal_2043912 <= p47_literal_2043912;
    p48_literal_2043914 <= p47_literal_2043914;
    p48_literal_2043916 <= p47_literal_2043916;
    p48_literal_2043918 <= p47_literal_2043918;
    p48_literal_2043920 <= p47_literal_2043920;
    p48_literal_2043923 <= p47_literal_2043923;
  end

  // ===== Pipe stage 48:
  wire [7:0] p48_array_index_2052644_comb;
  wire [7:0] p48_array_index_2052645_comb;
  wire [7:0] p48_array_index_2052646_comb;
  wire [7:0] p48_array_index_2052647_comb;
  wire [7:0] p48_res7__618_comb;
  wire [7:0] p48_array_index_2052658_comb;
  wire [7:0] p48_array_index_2052659_comb;
  wire [7:0] p48_array_index_2052660_comb;
  wire [7:0] p48_res7__620_comb;
  wire [7:0] p48_array_index_2052670_comb;
  wire [7:0] p48_array_index_2052671_comb;
  wire [7:0] p48_array_index_2052672_comb;
  wire [7:0] p48_res7__622_comb;
  wire [7:0] p48_array_index_2052683_comb;
  wire [7:0] p48_array_index_2052684_comb;
  wire [7:0] p48_res7__624_comb;
  wire [7:0] p48_array_index_2052694_comb;
  wire [7:0] p48_array_index_2052695_comb;
  wire [7:0] p48_res7__626_comb;
  wire [7:0] p48_array_index_2052706_comb;
  wire [7:0] p48_res7__628_comb;
  wire [7:0] p48_array_index_2052716_comb;
  wire [7:0] p48_res7__630_comb;
  assign p48_array_index_2052644_comb = p47_literal_2043914[p47_res7__612];
  assign p48_array_index_2052645_comb = p47_literal_2043916[p47_res7__610];
  assign p48_array_index_2052646_comb = p47_literal_2043918[p47_res7__608];
  assign p48_array_index_2052647_comb = p47_literal_2043920[p47_array_index_2052438];
  assign p48_res7__618_comb = p47_literal_2043910[p47_res7__616] ^ p47_literal_2043912[p47_res7__614] ^ p48_array_index_2052644_comb ^ p48_array_index_2052645_comb ^ p48_array_index_2052646_comb ^ p48_array_index_2052647_comb ^ p47_array_index_2052439 ^ p47_literal_2043923[p47_array_index_2052440] ^ p47_array_index_2052441 ^ p47_array_index_2052476 ^ p47_literal_2043918[p47_array_index_2052443] ^ p47_literal_2043916[p47_array_index_2052460] ^ p47_literal_2043914[p47_array_index_2052445] ^ p47_literal_2043912[p47_array_index_2052462] ^ p47_literal_2043910[p47_array_index_2052447] ^ p47_array_index_2052448;
  assign p48_array_index_2052658_comb = p47_literal_2043916[p47_res7__612];
  assign p48_array_index_2052659_comb = p47_literal_2043918[p47_res7__610];
  assign p48_array_index_2052660_comb = p47_literal_2043920[p47_res7__608];
  assign p48_res7__620_comb = p47_literal_2043910[p48_res7__618_comb] ^ p47_literal_2043912[p47_res7__616] ^ p47_literal_2043914[p47_res7__614] ^ p48_array_index_2052658_comb ^ p48_array_index_2052659_comb ^ p48_array_index_2052660_comb ^ p47_array_index_2052438 ^ p47_literal_2043923[p47_array_index_2052439] ^ p47_array_index_2052440 ^ p47_array_index_2052490 ^ p47_array_index_2052458 ^ p47_literal_2043916[p47_array_index_2052443] ^ p47_literal_2043914[p47_array_index_2052460] ^ p47_literal_2043912[p47_array_index_2052445] ^ p47_literal_2043910[p47_array_index_2052462] ^ p47_array_index_2052447;
  assign p48_array_index_2052670_comb = p47_literal_2043916[p47_res7__614];
  assign p48_array_index_2052671_comb = p47_literal_2043918[p47_res7__612];
  assign p48_array_index_2052672_comb = p47_literal_2043920[p47_res7__610];
  assign p48_res7__622_comb = p47_literal_2043910[p48_res7__620_comb] ^ p47_literal_2043912[p48_res7__618_comb] ^ p47_literal_2043914[p47_res7__616] ^ p48_array_index_2052670_comb ^ p48_array_index_2052671_comb ^ p48_array_index_2052672_comb ^ p47_res7__608 ^ p47_literal_2043923[p47_array_index_2052438] ^ p47_array_index_2052439 ^ p47_array_index_2052504 ^ p47_array_index_2052475 ^ p47_literal_2043916[p47_array_index_2052442] ^ p47_literal_2043914[p47_array_index_2052443] ^ p47_literal_2043912[p47_array_index_2052460] ^ p47_literal_2043910[p47_array_index_2052445] ^ p47_array_index_2052462;
  assign p48_array_index_2052683_comb = p47_literal_2043918[p47_res7__614];
  assign p48_array_index_2052684_comb = p47_literal_2043920[p47_res7__612];
  assign p48_res7__624_comb = p47_literal_2043910[p48_res7__622_comb] ^ p47_literal_2043912[p48_res7__620_comb] ^ p47_literal_2043914[p48_res7__618_comb] ^ p47_literal_2043916[p47_res7__616] ^ p48_array_index_2052683_comb ^ p48_array_index_2052684_comb ^ p47_res7__610 ^ p47_literal_2043923[p47_res7__608] ^ p47_array_index_2052438 ^ p47_array_index_2052518 ^ p47_array_index_2052489 ^ p47_array_index_2052457 ^ p47_literal_2043914[p47_array_index_2052442] ^ p47_literal_2043912[p47_array_index_2052443] ^ p47_literal_2043910[p47_array_index_2052460] ^ p47_array_index_2052445;
  assign p48_array_index_2052694_comb = p47_literal_2043918[p47_res7__616];
  assign p48_array_index_2052695_comb = p47_literal_2043920[p47_res7__614];
  assign p48_res7__626_comb = p47_literal_2043910[p48_res7__624_comb] ^ p47_literal_2043912[p48_res7__622_comb] ^ p47_literal_2043914[p48_res7__620_comb] ^ p47_literal_2043916[p48_res7__618_comb] ^ p48_array_index_2052694_comb ^ p48_array_index_2052695_comb ^ p47_res7__612 ^ p47_literal_2043923[p47_res7__610] ^ p47_res7__608 ^ p48_array_index_2052647_comb ^ p47_array_index_2052503 ^ p47_array_index_2052474 ^ p47_literal_2043914[p47_array_index_2052441] ^ p47_literal_2043912[p47_array_index_2052442] ^ p47_literal_2043910[p47_array_index_2052443] ^ p47_array_index_2052460;
  assign p48_array_index_2052706_comb = p47_literal_2043920[p47_res7__616];
  assign p48_res7__628_comb = p47_literal_2043910[p48_res7__626_comb] ^ p47_literal_2043912[p48_res7__624_comb] ^ p47_literal_2043914[p48_res7__622_comb] ^ p47_literal_2043916[p48_res7__620_comb] ^ p47_literal_2043918[p48_res7__618_comb] ^ p48_array_index_2052706_comb ^ p47_res7__614 ^ p47_literal_2043923[p47_res7__612] ^ p47_res7__610 ^ p48_array_index_2052660_comb ^ p47_array_index_2052517 ^ p47_array_index_2052488 ^ p47_array_index_2052456 ^ p47_literal_2043912[p47_array_index_2052441] ^ p47_literal_2043910[p47_array_index_2052442] ^ p47_array_index_2052443;
  assign p48_array_index_2052716_comb = p47_literal_2043920[p48_res7__618_comb];
  assign p48_res7__630_comb = p47_literal_2043910[p48_res7__628_comb] ^ p47_literal_2043912[p48_res7__626_comb] ^ p47_literal_2043914[p48_res7__624_comb] ^ p47_literal_2043916[p48_res7__622_comb] ^ p47_literal_2043918[p48_res7__620_comb] ^ p48_array_index_2052716_comb ^ p47_res7__616 ^ p47_literal_2043923[p47_res7__614] ^ p47_res7__612 ^ p48_array_index_2052672_comb ^ p48_array_index_2052646_comb ^ p47_array_index_2052502 ^ p47_array_index_2052473 ^ p47_literal_2043912[p47_array_index_2052440] ^ p47_literal_2043910[p47_array_index_2052441] ^ p47_array_index_2052442;

  // Registers for pipe stage 48:
  reg [127:0] p48_encoded;
  reg [127:0] p48_bit_slice_2043893;
  reg [127:0] p48_bit_slice_2044018;
  reg [127:0] p48_k3;
  reg [127:0] p48_k2;
  reg [127:0] p48_k5;
  reg [127:0] p48_k4;
  reg [127:0] p48_xor_2051922;
  reg [127:0] p48_xor_2052422;
  reg [7:0] p48_array_index_2052438;
  reg [7:0] p48_array_index_2052439;
  reg [7:0] p48_array_index_2052440;
  reg [7:0] p48_array_index_2052441;
  reg [7:0] p48_array_index_2052454;
  reg [7:0] p48_array_index_2052455;
  reg [7:0] p48_res7__608;
  reg [7:0] p48_array_index_2052471;
  reg [7:0] p48_array_index_2052472;
  reg [7:0] p48_res7__610;
  reg [7:0] p48_array_index_2052486;
  reg [7:0] p48_array_index_2052487;
  reg [7:0] p48_res7__612;
  reg [7:0] p48_array_index_2052500;
  reg [7:0] p48_array_index_2052501;
  reg [7:0] p48_res7__614;
  reg [7:0] p48_array_index_2052515;
  reg [7:0] p48_array_index_2052516;
  reg [7:0] p48_res7__616;
  reg [7:0] p48_array_index_2052644;
  reg [7:0] p48_array_index_2052645;
  reg [7:0] p48_res7__618;
  reg [7:0] p48_array_index_2052658;
  reg [7:0] p48_array_index_2052659;
  reg [7:0] p48_res7__620;
  reg [7:0] p48_array_index_2052670;
  reg [7:0] p48_array_index_2052671;
  reg [7:0] p48_res7__622;
  reg [7:0] p48_array_index_2052683;
  reg [7:0] p48_array_index_2052684;
  reg [7:0] p48_res7__624;
  reg [7:0] p48_array_index_2052694;
  reg [7:0] p48_array_index_2052695;
  reg [7:0] p48_res7__626;
  reg [7:0] p48_array_index_2052706;
  reg [7:0] p48_res7__628;
  reg [7:0] p48_array_index_2052716;
  reg [7:0] p48_res7__630;
  reg [7:0] p49_literal_2043896[256];
  reg [7:0] p49_literal_2043910[256];
  reg [7:0] p49_literal_2043912[256];
  reg [7:0] p49_literal_2043914[256];
  reg [7:0] p49_literal_2043916[256];
  reg [7:0] p49_literal_2043918[256];
  reg [7:0] p49_literal_2043920[256];
  reg [7:0] p49_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p48_encoded <= p47_encoded;
    p48_bit_slice_2043893 <= p47_bit_slice_2043893;
    p48_bit_slice_2044018 <= p47_bit_slice_2044018;
    p48_k3 <= p47_k3;
    p48_k2 <= p47_k2;
    p48_k5 <= p47_k5;
    p48_k4 <= p47_k4;
    p48_xor_2051922 <= p47_xor_2051922;
    p48_xor_2052422 <= p47_xor_2052422;
    p48_array_index_2052438 <= p47_array_index_2052438;
    p48_array_index_2052439 <= p47_array_index_2052439;
    p48_array_index_2052440 <= p47_array_index_2052440;
    p48_array_index_2052441 <= p47_array_index_2052441;
    p48_array_index_2052454 <= p47_array_index_2052454;
    p48_array_index_2052455 <= p47_array_index_2052455;
    p48_res7__608 <= p47_res7__608;
    p48_array_index_2052471 <= p47_array_index_2052471;
    p48_array_index_2052472 <= p47_array_index_2052472;
    p48_res7__610 <= p47_res7__610;
    p48_array_index_2052486 <= p47_array_index_2052486;
    p48_array_index_2052487 <= p47_array_index_2052487;
    p48_res7__612 <= p47_res7__612;
    p48_array_index_2052500 <= p47_array_index_2052500;
    p48_array_index_2052501 <= p47_array_index_2052501;
    p48_res7__614 <= p47_res7__614;
    p48_array_index_2052515 <= p47_array_index_2052515;
    p48_array_index_2052516 <= p47_array_index_2052516;
    p48_res7__616 <= p47_res7__616;
    p48_array_index_2052644 <= p48_array_index_2052644_comb;
    p48_array_index_2052645 <= p48_array_index_2052645_comb;
    p48_res7__618 <= p48_res7__618_comb;
    p48_array_index_2052658 <= p48_array_index_2052658_comb;
    p48_array_index_2052659 <= p48_array_index_2052659_comb;
    p48_res7__620 <= p48_res7__620_comb;
    p48_array_index_2052670 <= p48_array_index_2052670_comb;
    p48_array_index_2052671 <= p48_array_index_2052671_comb;
    p48_res7__622 <= p48_res7__622_comb;
    p48_array_index_2052683 <= p48_array_index_2052683_comb;
    p48_array_index_2052684 <= p48_array_index_2052684_comb;
    p48_res7__624 <= p48_res7__624_comb;
    p48_array_index_2052694 <= p48_array_index_2052694_comb;
    p48_array_index_2052695 <= p48_array_index_2052695_comb;
    p48_res7__626 <= p48_res7__626_comb;
    p48_array_index_2052706 <= p48_array_index_2052706_comb;
    p48_res7__628 <= p48_res7__628_comb;
    p48_array_index_2052716 <= p48_array_index_2052716_comb;
    p48_res7__630 <= p48_res7__630_comb;
    p49_literal_2043896 <= p48_literal_2043896;
    p49_literal_2043910 <= p48_literal_2043910;
    p49_literal_2043912 <= p48_literal_2043912;
    p49_literal_2043914 <= p48_literal_2043914;
    p49_literal_2043916 <= p48_literal_2043916;
    p49_literal_2043918 <= p48_literal_2043918;
    p49_literal_2043920 <= p48_literal_2043920;
    p49_literal_2043923 <= p48_literal_2043923;
  end

  // ===== Pipe stage 49:
  wire [7:0] p49_res7__632_comb;
  wire [7:0] p49_res7__634_comb;
  wire [7:0] p49_res7__636_comb;
  wire [7:0] p49_res7__638_comb;
  wire [127:0] p49_res__19_comb;
  wire [127:0] p49_xor_2052866_comb;
  wire [127:0] p49_addedKey__52_comb;
  wire [7:0] p49_array_index_2052882_comb;
  wire [7:0] p49_array_index_2052883_comb;
  wire [7:0] p49_array_index_2052884_comb;
  wire [7:0] p49_array_index_2052885_comb;
  wire [7:0] p49_array_index_2052886_comb;
  wire [7:0] p49_array_index_2052887_comb;
  wire [7:0] p49_array_index_2052889_comb;
  wire [7:0] p49_array_index_2052891_comb;
  wire [7:0] p49_array_index_2052892_comb;
  wire [7:0] p49_array_index_2052893_comb;
  wire [7:0] p49_array_index_2052894_comb;
  wire [7:0] p49_array_index_2052895_comb;
  wire [7:0] p49_array_index_2052896_comb;
  wire [7:0] p49_array_index_2052898_comb;
  wire [7:0] p49_array_index_2052899_comb;
  wire [7:0] p49_array_index_2052900_comb;
  wire [7:0] p49_array_index_2052901_comb;
  wire [7:0] p49_array_index_2052902_comb;
  wire [7:0] p49_array_index_2052903_comb;
  wire [7:0] p49_array_index_2052904_comb;
  wire [7:0] p49_array_index_2052906_comb;
  wire [7:0] p49_res7__640_comb;
  wire [7:0] p49_array_index_2052915_comb;
  wire [7:0] p49_array_index_2052916_comb;
  wire [7:0] p49_array_index_2052917_comb;
  wire [7:0] p49_array_index_2052918_comb;
  wire [7:0] p49_array_index_2052919_comb;
  wire [7:0] p49_array_index_2052920_comb;
  wire [7:0] p49_res7__642_comb;
  assign p49_res7__632_comb = p48_literal_2043910[p48_res7__630] ^ p48_literal_2043912[p48_res7__628] ^ p48_literal_2043914[p48_res7__626] ^ p48_literal_2043916[p48_res7__624] ^ p48_literal_2043918[p48_res7__622] ^ p48_literal_2043920[p48_res7__620] ^ p48_res7__618 ^ p48_literal_2043923[p48_res7__616] ^ p48_res7__614 ^ p48_array_index_2052684 ^ p48_array_index_2052659 ^ p48_array_index_2052516 ^ p48_array_index_2052487 ^ p48_array_index_2052455 ^ p48_literal_2043910[p48_array_index_2052440] ^ p48_array_index_2052441;
  assign p49_res7__634_comb = p48_literal_2043910[p49_res7__632_comb] ^ p48_literal_2043912[p48_res7__630] ^ p48_literal_2043914[p48_res7__628] ^ p48_literal_2043916[p48_res7__626] ^ p48_literal_2043918[p48_res7__624] ^ p48_literal_2043920[p48_res7__622] ^ p48_res7__620 ^ p48_literal_2043923[p48_res7__618] ^ p48_res7__616 ^ p48_array_index_2052695 ^ p48_array_index_2052671 ^ p48_array_index_2052645 ^ p48_array_index_2052501 ^ p48_array_index_2052472 ^ p48_literal_2043910[p48_array_index_2052439] ^ p48_array_index_2052440;
  assign p49_res7__636_comb = p48_literal_2043910[p49_res7__634_comb] ^ p48_literal_2043912[p49_res7__632_comb] ^ p48_literal_2043914[p48_res7__630] ^ p48_literal_2043916[p48_res7__628] ^ p48_literal_2043918[p48_res7__626] ^ p48_literal_2043920[p48_res7__624] ^ p48_res7__622 ^ p48_literal_2043923[p48_res7__620] ^ p48_res7__618 ^ p48_array_index_2052706 ^ p48_array_index_2052683 ^ p48_array_index_2052658 ^ p48_array_index_2052515 ^ p48_array_index_2052486 ^ p48_array_index_2052454 ^ p48_array_index_2052439;
  assign p49_res7__638_comb = p48_literal_2043910[p49_res7__636_comb] ^ p48_literal_2043912[p49_res7__634_comb] ^ p48_literal_2043914[p49_res7__632_comb] ^ p48_literal_2043916[p48_res7__630] ^ p48_literal_2043918[p48_res7__628] ^ p48_literal_2043920[p48_res7__626] ^ p48_res7__624 ^ p48_literal_2043923[p48_res7__622] ^ p48_res7__620 ^ p48_array_index_2052716 ^ p48_array_index_2052694 ^ p48_array_index_2052670 ^ p48_array_index_2052644 ^ p48_array_index_2052500 ^ p48_array_index_2052471 ^ p48_array_index_2052438;
  assign p49_res__19_comb = {p49_res7__638_comb, p49_res7__636_comb, p49_res7__634_comb, p49_res7__632_comb, p48_res7__630, p48_res7__628, p48_res7__626, p48_res7__624, p48_res7__622, p48_res7__620, p48_res7__618, p48_res7__616, p48_res7__614, p48_res7__612, p48_res7__610, p48_res7__608};
  assign p49_xor_2052866_comb = p49_res__19_comb ^ p48_xor_2051922;
  assign p49_addedKey__52_comb = p49_xor_2052866_comb ^ 128'h3add_0155_10a1_fdcc_738e_8d93_6146_d515;
  assign p49_array_index_2052882_comb = p48_literal_2043896[p49_addedKey__52_comb[127:120]];
  assign p49_array_index_2052883_comb = p48_literal_2043896[p49_addedKey__52_comb[119:112]];
  assign p49_array_index_2052884_comb = p48_literal_2043896[p49_addedKey__52_comb[111:104]];
  assign p49_array_index_2052885_comb = p48_literal_2043896[p49_addedKey__52_comb[103:96]];
  assign p49_array_index_2052886_comb = p48_literal_2043896[p49_addedKey__52_comb[95:88]];
  assign p49_array_index_2052887_comb = p48_literal_2043896[p49_addedKey__52_comb[87:80]];
  assign p49_array_index_2052889_comb = p48_literal_2043896[p49_addedKey__52_comb[71:64]];
  assign p49_array_index_2052891_comb = p48_literal_2043896[p49_addedKey__52_comb[55:48]];
  assign p49_array_index_2052892_comb = p48_literal_2043896[p49_addedKey__52_comb[47:40]];
  assign p49_array_index_2052893_comb = p48_literal_2043896[p49_addedKey__52_comb[39:32]];
  assign p49_array_index_2052894_comb = p48_literal_2043896[p49_addedKey__52_comb[31:24]];
  assign p49_array_index_2052895_comb = p48_literal_2043896[p49_addedKey__52_comb[23:16]];
  assign p49_array_index_2052896_comb = p48_literal_2043896[p49_addedKey__52_comb[15:8]];
  assign p49_array_index_2052898_comb = p48_literal_2043910[p49_array_index_2052882_comb];
  assign p49_array_index_2052899_comb = p48_literal_2043912[p49_array_index_2052883_comb];
  assign p49_array_index_2052900_comb = p48_literal_2043914[p49_array_index_2052884_comb];
  assign p49_array_index_2052901_comb = p48_literal_2043916[p49_array_index_2052885_comb];
  assign p49_array_index_2052902_comb = p48_literal_2043918[p49_array_index_2052886_comb];
  assign p49_array_index_2052903_comb = p48_literal_2043920[p49_array_index_2052887_comb];
  assign p49_array_index_2052904_comb = p48_literal_2043896[p49_addedKey__52_comb[79:72]];
  assign p49_array_index_2052906_comb = p48_literal_2043896[p49_addedKey__52_comb[63:56]];
  assign p49_res7__640_comb = p49_array_index_2052898_comb ^ p49_array_index_2052899_comb ^ p49_array_index_2052900_comb ^ p49_array_index_2052901_comb ^ p49_array_index_2052902_comb ^ p49_array_index_2052903_comb ^ p49_array_index_2052904_comb ^ p48_literal_2043923[p49_array_index_2052889_comb] ^ p49_array_index_2052906_comb ^ p48_literal_2043920[p49_array_index_2052891_comb] ^ p48_literal_2043918[p49_array_index_2052892_comb] ^ p48_literal_2043916[p49_array_index_2052893_comb] ^ p48_literal_2043914[p49_array_index_2052894_comb] ^ p48_literal_2043912[p49_array_index_2052895_comb] ^ p48_literal_2043910[p49_array_index_2052896_comb] ^ p48_literal_2043896[p49_addedKey__52_comb[7:0]];
  assign p49_array_index_2052915_comb = p48_literal_2043910[p49_res7__640_comb];
  assign p49_array_index_2052916_comb = p48_literal_2043912[p49_array_index_2052882_comb];
  assign p49_array_index_2052917_comb = p48_literal_2043914[p49_array_index_2052883_comb];
  assign p49_array_index_2052918_comb = p48_literal_2043916[p49_array_index_2052884_comb];
  assign p49_array_index_2052919_comb = p48_literal_2043918[p49_array_index_2052885_comb];
  assign p49_array_index_2052920_comb = p48_literal_2043920[p49_array_index_2052886_comb];
  assign p49_res7__642_comb = p49_array_index_2052915_comb ^ p49_array_index_2052916_comb ^ p49_array_index_2052917_comb ^ p49_array_index_2052918_comb ^ p49_array_index_2052919_comb ^ p49_array_index_2052920_comb ^ p49_array_index_2052887_comb ^ p48_literal_2043923[p49_array_index_2052904_comb] ^ p49_array_index_2052889_comb ^ p48_literal_2043920[p49_array_index_2052906_comb] ^ p48_literal_2043918[p49_array_index_2052891_comb] ^ p48_literal_2043916[p49_array_index_2052892_comb] ^ p48_literal_2043914[p49_array_index_2052893_comb] ^ p48_literal_2043912[p49_array_index_2052894_comb] ^ p48_literal_2043910[p49_array_index_2052895_comb] ^ p49_array_index_2052896_comb;

  // Registers for pipe stage 49:
  reg [127:0] p49_encoded;
  reg [127:0] p49_bit_slice_2043893;
  reg [127:0] p49_bit_slice_2044018;
  reg [127:0] p49_k3;
  reg [127:0] p49_k2;
  reg [127:0] p49_k5;
  reg [127:0] p49_k4;
  reg [127:0] p49_xor_2052422;
  reg [127:0] p49_xor_2052866;
  reg [7:0] p49_array_index_2052882;
  reg [7:0] p49_array_index_2052883;
  reg [7:0] p49_array_index_2052884;
  reg [7:0] p49_array_index_2052885;
  reg [7:0] p49_array_index_2052886;
  reg [7:0] p49_array_index_2052887;
  reg [7:0] p49_array_index_2052889;
  reg [7:0] p49_array_index_2052891;
  reg [7:0] p49_array_index_2052892;
  reg [7:0] p49_array_index_2052893;
  reg [7:0] p49_array_index_2052894;
  reg [7:0] p49_array_index_2052895;
  reg [7:0] p49_array_index_2052898;
  reg [7:0] p49_array_index_2052899;
  reg [7:0] p49_array_index_2052900;
  reg [7:0] p49_array_index_2052901;
  reg [7:0] p49_array_index_2052902;
  reg [7:0] p49_array_index_2052903;
  reg [7:0] p49_array_index_2052904;
  reg [7:0] p49_array_index_2052906;
  reg [7:0] p49_res7__640;
  reg [7:0] p49_array_index_2052915;
  reg [7:0] p49_array_index_2052916;
  reg [7:0] p49_array_index_2052917;
  reg [7:0] p49_array_index_2052918;
  reg [7:0] p49_array_index_2052919;
  reg [7:0] p49_array_index_2052920;
  reg [7:0] p49_res7__642;
  reg [7:0] p50_literal_2043896[256];
  reg [7:0] p50_literal_2043910[256];
  reg [7:0] p50_literal_2043912[256];
  reg [7:0] p50_literal_2043914[256];
  reg [7:0] p50_literal_2043916[256];
  reg [7:0] p50_literal_2043918[256];
  reg [7:0] p50_literal_2043920[256];
  reg [7:0] p50_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p49_encoded <= p48_encoded;
    p49_bit_slice_2043893 <= p48_bit_slice_2043893;
    p49_bit_slice_2044018 <= p48_bit_slice_2044018;
    p49_k3 <= p48_k3;
    p49_k2 <= p48_k2;
    p49_k5 <= p48_k5;
    p49_k4 <= p48_k4;
    p49_xor_2052422 <= p48_xor_2052422;
    p49_xor_2052866 <= p49_xor_2052866_comb;
    p49_array_index_2052882 <= p49_array_index_2052882_comb;
    p49_array_index_2052883 <= p49_array_index_2052883_comb;
    p49_array_index_2052884 <= p49_array_index_2052884_comb;
    p49_array_index_2052885 <= p49_array_index_2052885_comb;
    p49_array_index_2052886 <= p49_array_index_2052886_comb;
    p49_array_index_2052887 <= p49_array_index_2052887_comb;
    p49_array_index_2052889 <= p49_array_index_2052889_comb;
    p49_array_index_2052891 <= p49_array_index_2052891_comb;
    p49_array_index_2052892 <= p49_array_index_2052892_comb;
    p49_array_index_2052893 <= p49_array_index_2052893_comb;
    p49_array_index_2052894 <= p49_array_index_2052894_comb;
    p49_array_index_2052895 <= p49_array_index_2052895_comb;
    p49_array_index_2052898 <= p49_array_index_2052898_comb;
    p49_array_index_2052899 <= p49_array_index_2052899_comb;
    p49_array_index_2052900 <= p49_array_index_2052900_comb;
    p49_array_index_2052901 <= p49_array_index_2052901_comb;
    p49_array_index_2052902 <= p49_array_index_2052902_comb;
    p49_array_index_2052903 <= p49_array_index_2052903_comb;
    p49_array_index_2052904 <= p49_array_index_2052904_comb;
    p49_array_index_2052906 <= p49_array_index_2052906_comb;
    p49_res7__640 <= p49_res7__640_comb;
    p49_array_index_2052915 <= p49_array_index_2052915_comb;
    p49_array_index_2052916 <= p49_array_index_2052916_comb;
    p49_array_index_2052917 <= p49_array_index_2052917_comb;
    p49_array_index_2052918 <= p49_array_index_2052918_comb;
    p49_array_index_2052919 <= p49_array_index_2052919_comb;
    p49_array_index_2052920 <= p49_array_index_2052920_comb;
    p49_res7__642 <= p49_res7__642_comb;
    p50_literal_2043896 <= p49_literal_2043896;
    p50_literal_2043910 <= p49_literal_2043910;
    p50_literal_2043912 <= p49_literal_2043912;
    p50_literal_2043914 <= p49_literal_2043914;
    p50_literal_2043916 <= p49_literal_2043916;
    p50_literal_2043918 <= p49_literal_2043918;
    p50_literal_2043920 <= p49_literal_2043920;
    p50_literal_2043923 <= p49_literal_2043923;
  end

  // ===== Pipe stage 50:
  wire [7:0] p50_array_index_2053020_comb;
  wire [7:0] p50_array_index_2053021_comb;
  wire [7:0] p50_array_index_2053022_comb;
  wire [7:0] p50_array_index_2053023_comb;
  wire [7:0] p50_array_index_2053024_comb;
  wire [7:0] p50_res7__644_comb;
  wire [7:0] p50_array_index_2053034_comb;
  wire [7:0] p50_array_index_2053035_comb;
  wire [7:0] p50_array_index_2053036_comb;
  wire [7:0] p50_array_index_2053037_comb;
  wire [7:0] p50_array_index_2053038_comb;
  wire [7:0] p50_res7__646_comb;
  wire [7:0] p50_array_index_2053049_comb;
  wire [7:0] p50_array_index_2053050_comb;
  wire [7:0] p50_array_index_2053051_comb;
  wire [7:0] p50_array_index_2053052_comb;
  wire [7:0] p50_res7__648_comb;
  wire [7:0] p50_array_index_2053062_comb;
  wire [7:0] p50_array_index_2053063_comb;
  wire [7:0] p50_array_index_2053064_comb;
  wire [7:0] p50_array_index_2053065_comb;
  wire [7:0] p50_res7__650_comb;
  wire [7:0] p50_array_index_2053076_comb;
  wire [7:0] p50_array_index_2053077_comb;
  wire [7:0] p50_array_index_2053078_comb;
  wire [7:0] p50_res7__652_comb;
  wire [7:0] p50_array_index_2053088_comb;
  wire [7:0] p50_array_index_2053089_comb;
  wire [7:0] p50_array_index_2053090_comb;
  wire [7:0] p50_res7__654_comb;
  wire [7:0] p50_array_index_2053101_comb;
  wire [7:0] p50_array_index_2053102_comb;
  wire [7:0] p50_res7__656_comb;
  assign p50_array_index_2053020_comb = p49_literal_2043912[p49_res7__640];
  assign p50_array_index_2053021_comb = p49_literal_2043914[p49_array_index_2052882];
  assign p50_array_index_2053022_comb = p49_literal_2043916[p49_array_index_2052883];
  assign p50_array_index_2053023_comb = p49_literal_2043918[p49_array_index_2052884];
  assign p50_array_index_2053024_comb = p49_literal_2043920[p49_array_index_2052885];
  assign p50_res7__644_comb = p49_literal_2043910[p49_res7__642] ^ p50_array_index_2053020_comb ^ p50_array_index_2053021_comb ^ p50_array_index_2053022_comb ^ p50_array_index_2053023_comb ^ p50_array_index_2053024_comb ^ p49_array_index_2052886 ^ p49_literal_2043923[p49_array_index_2052887] ^ p49_array_index_2052904 ^ p49_literal_2043920[p49_array_index_2052889] ^ p49_literal_2043918[p49_array_index_2052906] ^ p49_literal_2043916[p49_array_index_2052891] ^ p49_literal_2043914[p49_array_index_2052892] ^ p49_literal_2043912[p49_array_index_2052893] ^ p49_literal_2043910[p49_array_index_2052894] ^ p49_array_index_2052895;
  assign p50_array_index_2053034_comb = p49_literal_2043912[p49_res7__642];
  assign p50_array_index_2053035_comb = p49_literal_2043914[p49_res7__640];
  assign p50_array_index_2053036_comb = p49_literal_2043916[p49_array_index_2052882];
  assign p50_array_index_2053037_comb = p49_literal_2043918[p49_array_index_2052883];
  assign p50_array_index_2053038_comb = p49_literal_2043920[p49_array_index_2052884];
  assign p50_res7__646_comb = p49_literal_2043910[p50_res7__644_comb] ^ p50_array_index_2053034_comb ^ p50_array_index_2053035_comb ^ p50_array_index_2053036_comb ^ p50_array_index_2053037_comb ^ p50_array_index_2053038_comb ^ p49_array_index_2052885 ^ p49_literal_2043923[p49_array_index_2052886] ^ p49_array_index_2052887 ^ p49_literal_2043920[p49_array_index_2052904] ^ p49_literal_2043918[p49_array_index_2052889] ^ p49_literal_2043916[p49_array_index_2052906] ^ p49_literal_2043914[p49_array_index_2052891] ^ p49_literal_2043912[p49_array_index_2052892] ^ p49_literal_2043910[p49_array_index_2052893] ^ p49_array_index_2052894;
  assign p50_array_index_2053049_comb = p49_literal_2043914[p49_res7__642];
  assign p50_array_index_2053050_comb = p49_literal_2043916[p49_res7__640];
  assign p50_array_index_2053051_comb = p49_literal_2043918[p49_array_index_2052882];
  assign p50_array_index_2053052_comb = p49_literal_2043920[p49_array_index_2052883];
  assign p50_res7__648_comb = p49_literal_2043910[p50_res7__646_comb] ^ p49_literal_2043912[p50_res7__644_comb] ^ p50_array_index_2053049_comb ^ p50_array_index_2053050_comb ^ p50_array_index_2053051_comb ^ p50_array_index_2053052_comb ^ p49_array_index_2052884 ^ p49_literal_2043923[p49_array_index_2052885] ^ p49_array_index_2052886 ^ p49_array_index_2052903 ^ p49_literal_2043918[p49_array_index_2052904] ^ p49_literal_2043916[p49_array_index_2052889] ^ p49_literal_2043914[p49_array_index_2052906] ^ p49_literal_2043912[p49_array_index_2052891] ^ p49_literal_2043910[p49_array_index_2052892] ^ p49_array_index_2052893;
  assign p50_array_index_2053062_comb = p49_literal_2043914[p50_res7__644_comb];
  assign p50_array_index_2053063_comb = p49_literal_2043916[p49_res7__642];
  assign p50_array_index_2053064_comb = p49_literal_2043918[p49_res7__640];
  assign p50_array_index_2053065_comb = p49_literal_2043920[p49_array_index_2052882];
  assign p50_res7__650_comb = p49_literal_2043910[p50_res7__648_comb] ^ p49_literal_2043912[p50_res7__646_comb] ^ p50_array_index_2053062_comb ^ p50_array_index_2053063_comb ^ p50_array_index_2053064_comb ^ p50_array_index_2053065_comb ^ p49_array_index_2052883 ^ p49_literal_2043923[p49_array_index_2052884] ^ p49_array_index_2052885 ^ p49_array_index_2052920 ^ p49_literal_2043918[p49_array_index_2052887] ^ p49_literal_2043916[p49_array_index_2052904] ^ p49_literal_2043914[p49_array_index_2052889] ^ p49_literal_2043912[p49_array_index_2052906] ^ p49_literal_2043910[p49_array_index_2052891] ^ p49_array_index_2052892;
  assign p50_array_index_2053076_comb = p49_literal_2043916[p50_res7__644_comb];
  assign p50_array_index_2053077_comb = p49_literal_2043918[p49_res7__642];
  assign p50_array_index_2053078_comb = p49_literal_2043920[p49_res7__640];
  assign p50_res7__652_comb = p49_literal_2043910[p50_res7__650_comb] ^ p49_literal_2043912[p50_res7__648_comb] ^ p49_literal_2043914[p50_res7__646_comb] ^ p50_array_index_2053076_comb ^ p50_array_index_2053077_comb ^ p50_array_index_2053078_comb ^ p49_array_index_2052882 ^ p49_literal_2043923[p49_array_index_2052883] ^ p49_array_index_2052884 ^ p50_array_index_2053024_comb ^ p49_array_index_2052902 ^ p49_literal_2043916[p49_array_index_2052887] ^ p49_literal_2043914[p49_array_index_2052904] ^ p49_literal_2043912[p49_array_index_2052889] ^ p49_literal_2043910[p49_array_index_2052906] ^ p49_array_index_2052891;
  assign p50_array_index_2053088_comb = p49_literal_2043916[p50_res7__646_comb];
  assign p50_array_index_2053089_comb = p49_literal_2043918[p50_res7__644_comb];
  assign p50_array_index_2053090_comb = p49_literal_2043920[p49_res7__642];
  assign p50_res7__654_comb = p49_literal_2043910[p50_res7__652_comb] ^ p49_literal_2043912[p50_res7__650_comb] ^ p49_literal_2043914[p50_res7__648_comb] ^ p50_array_index_2053088_comb ^ p50_array_index_2053089_comb ^ p50_array_index_2053090_comb ^ p49_res7__640 ^ p49_literal_2043923[p49_array_index_2052882] ^ p49_array_index_2052883 ^ p50_array_index_2053038_comb ^ p49_array_index_2052919 ^ p49_literal_2043916[p49_array_index_2052886] ^ p49_literal_2043914[p49_array_index_2052887] ^ p49_literal_2043912[p49_array_index_2052904] ^ p49_literal_2043910[p49_array_index_2052889] ^ p49_array_index_2052906;
  assign p50_array_index_2053101_comb = p49_literal_2043918[p50_res7__646_comb];
  assign p50_array_index_2053102_comb = p49_literal_2043920[p50_res7__644_comb];
  assign p50_res7__656_comb = p49_literal_2043910[p50_res7__654_comb] ^ p49_literal_2043912[p50_res7__652_comb] ^ p49_literal_2043914[p50_res7__650_comb] ^ p49_literal_2043916[p50_res7__648_comb] ^ p50_array_index_2053101_comb ^ p50_array_index_2053102_comb ^ p49_res7__642 ^ p49_literal_2043923[p49_res7__640] ^ p49_array_index_2052882 ^ p50_array_index_2053052_comb ^ p50_array_index_2053023_comb ^ p49_array_index_2052901 ^ p49_literal_2043914[p49_array_index_2052886] ^ p49_literal_2043912[p49_array_index_2052887] ^ p49_literal_2043910[p49_array_index_2052904] ^ p49_array_index_2052889;

  // Registers for pipe stage 50:
  reg [127:0] p50_encoded;
  reg [127:0] p50_bit_slice_2043893;
  reg [127:0] p50_bit_slice_2044018;
  reg [127:0] p50_k3;
  reg [127:0] p50_k2;
  reg [127:0] p50_k5;
  reg [127:0] p50_k4;
  reg [127:0] p50_xor_2052422;
  reg [127:0] p50_xor_2052866;
  reg [7:0] p50_array_index_2052882;
  reg [7:0] p50_array_index_2052883;
  reg [7:0] p50_array_index_2052884;
  reg [7:0] p50_array_index_2052885;
  reg [7:0] p50_array_index_2052886;
  reg [7:0] p50_array_index_2052887;
  reg [7:0] p50_array_index_2052898;
  reg [7:0] p50_array_index_2052899;
  reg [7:0] p50_array_index_2052900;
  reg [7:0] p50_array_index_2052904;
  reg [7:0] p50_res7__640;
  reg [7:0] p50_array_index_2052915;
  reg [7:0] p50_array_index_2052916;
  reg [7:0] p50_array_index_2052917;
  reg [7:0] p50_array_index_2052918;
  reg [7:0] p50_res7__642;
  reg [7:0] p50_array_index_2053020;
  reg [7:0] p50_array_index_2053021;
  reg [7:0] p50_array_index_2053022;
  reg [7:0] p50_res7__644;
  reg [7:0] p50_array_index_2053034;
  reg [7:0] p50_array_index_2053035;
  reg [7:0] p50_array_index_2053036;
  reg [7:0] p50_array_index_2053037;
  reg [7:0] p50_res7__646;
  reg [7:0] p50_array_index_2053049;
  reg [7:0] p50_array_index_2053050;
  reg [7:0] p50_array_index_2053051;
  reg [7:0] p50_res7__648;
  reg [7:0] p50_array_index_2053062;
  reg [7:0] p50_array_index_2053063;
  reg [7:0] p50_array_index_2053064;
  reg [7:0] p50_array_index_2053065;
  reg [7:0] p50_res7__650;
  reg [7:0] p50_array_index_2053076;
  reg [7:0] p50_array_index_2053077;
  reg [7:0] p50_array_index_2053078;
  reg [7:0] p50_res7__652;
  reg [7:0] p50_array_index_2053088;
  reg [7:0] p50_array_index_2053089;
  reg [7:0] p50_array_index_2053090;
  reg [7:0] p50_res7__654;
  reg [7:0] p50_array_index_2053101;
  reg [7:0] p50_array_index_2053102;
  reg [7:0] p50_res7__656;
  reg [7:0] p51_literal_2043896[256];
  reg [7:0] p51_literal_2043910[256];
  reg [7:0] p51_literal_2043912[256];
  reg [7:0] p51_literal_2043914[256];
  reg [7:0] p51_literal_2043916[256];
  reg [7:0] p51_literal_2043918[256];
  reg [7:0] p51_literal_2043920[256];
  reg [7:0] p51_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p50_encoded <= p49_encoded;
    p50_bit_slice_2043893 <= p49_bit_slice_2043893;
    p50_bit_slice_2044018 <= p49_bit_slice_2044018;
    p50_k3 <= p49_k3;
    p50_k2 <= p49_k2;
    p50_k5 <= p49_k5;
    p50_k4 <= p49_k4;
    p50_xor_2052422 <= p49_xor_2052422;
    p50_xor_2052866 <= p49_xor_2052866;
    p50_array_index_2052882 <= p49_array_index_2052882;
    p50_array_index_2052883 <= p49_array_index_2052883;
    p50_array_index_2052884 <= p49_array_index_2052884;
    p50_array_index_2052885 <= p49_array_index_2052885;
    p50_array_index_2052886 <= p49_array_index_2052886;
    p50_array_index_2052887 <= p49_array_index_2052887;
    p50_array_index_2052898 <= p49_array_index_2052898;
    p50_array_index_2052899 <= p49_array_index_2052899;
    p50_array_index_2052900 <= p49_array_index_2052900;
    p50_array_index_2052904 <= p49_array_index_2052904;
    p50_res7__640 <= p49_res7__640;
    p50_array_index_2052915 <= p49_array_index_2052915;
    p50_array_index_2052916 <= p49_array_index_2052916;
    p50_array_index_2052917 <= p49_array_index_2052917;
    p50_array_index_2052918 <= p49_array_index_2052918;
    p50_res7__642 <= p49_res7__642;
    p50_array_index_2053020 <= p50_array_index_2053020_comb;
    p50_array_index_2053021 <= p50_array_index_2053021_comb;
    p50_array_index_2053022 <= p50_array_index_2053022_comb;
    p50_res7__644 <= p50_res7__644_comb;
    p50_array_index_2053034 <= p50_array_index_2053034_comb;
    p50_array_index_2053035 <= p50_array_index_2053035_comb;
    p50_array_index_2053036 <= p50_array_index_2053036_comb;
    p50_array_index_2053037 <= p50_array_index_2053037_comb;
    p50_res7__646 <= p50_res7__646_comb;
    p50_array_index_2053049 <= p50_array_index_2053049_comb;
    p50_array_index_2053050 <= p50_array_index_2053050_comb;
    p50_array_index_2053051 <= p50_array_index_2053051_comb;
    p50_res7__648 <= p50_res7__648_comb;
    p50_array_index_2053062 <= p50_array_index_2053062_comb;
    p50_array_index_2053063 <= p50_array_index_2053063_comb;
    p50_array_index_2053064 <= p50_array_index_2053064_comb;
    p50_array_index_2053065 <= p50_array_index_2053065_comb;
    p50_res7__650 <= p50_res7__650_comb;
    p50_array_index_2053076 <= p50_array_index_2053076_comb;
    p50_array_index_2053077 <= p50_array_index_2053077_comb;
    p50_array_index_2053078 <= p50_array_index_2053078_comb;
    p50_res7__652 <= p50_res7__652_comb;
    p50_array_index_2053088 <= p50_array_index_2053088_comb;
    p50_array_index_2053089 <= p50_array_index_2053089_comb;
    p50_array_index_2053090 <= p50_array_index_2053090_comb;
    p50_res7__654 <= p50_res7__654_comb;
    p50_array_index_2053101 <= p50_array_index_2053101_comb;
    p50_array_index_2053102 <= p50_array_index_2053102_comb;
    p50_res7__656 <= p50_res7__656_comb;
    p51_literal_2043896 <= p50_literal_2043896;
    p51_literal_2043910 <= p50_literal_2043910;
    p51_literal_2043912 <= p50_literal_2043912;
    p51_literal_2043914 <= p50_literal_2043914;
    p51_literal_2043916 <= p50_literal_2043916;
    p51_literal_2043918 <= p50_literal_2043918;
    p51_literal_2043920 <= p50_literal_2043920;
    p51_literal_2043923 <= p50_literal_2043923;
  end

  // ===== Pipe stage 51:
  wire [7:0] p51_array_index_2053236_comb;
  wire [7:0] p51_array_index_2053237_comb;
  wire [7:0] p51_res7__658_comb;
  wire [7:0] p51_array_index_2053248_comb;
  wire [7:0] p51_res7__660_comb;
  wire [7:0] p51_array_index_2053258_comb;
  wire [7:0] p51_res7__662_comb;
  wire [7:0] p51_res7__664_comb;
  wire [7:0] p51_res7__666_comb;
  wire [7:0] p51_res7__668_comb;
  wire [7:0] p51_res7__670_comb;
  wire [127:0] p51_res__20_comb;
  assign p51_array_index_2053236_comb = p50_literal_2043918[p50_res7__648];
  assign p51_array_index_2053237_comb = p50_literal_2043920[p50_res7__646];
  assign p51_res7__658_comb = p50_literal_2043910[p50_res7__656] ^ p50_literal_2043912[p50_res7__654] ^ p50_literal_2043914[p50_res7__652] ^ p50_literal_2043916[p50_res7__650] ^ p51_array_index_2053236_comb ^ p51_array_index_2053237_comb ^ p50_res7__644 ^ p50_literal_2043923[p50_res7__642] ^ p50_res7__640 ^ p50_array_index_2053065 ^ p50_array_index_2053037 ^ p50_array_index_2052918 ^ p50_literal_2043914[p50_array_index_2052885] ^ p50_literal_2043912[p50_array_index_2052886] ^ p50_literal_2043910[p50_array_index_2052887] ^ p50_array_index_2052904;
  assign p51_array_index_2053248_comb = p50_literal_2043920[p50_res7__648];
  assign p51_res7__660_comb = p50_literal_2043910[p51_res7__658_comb] ^ p50_literal_2043912[p50_res7__656] ^ p50_literal_2043914[p50_res7__654] ^ p50_literal_2043916[p50_res7__652] ^ p50_literal_2043918[p50_res7__650] ^ p51_array_index_2053248_comb ^ p50_res7__646 ^ p50_literal_2043923[p50_res7__644] ^ p50_res7__642 ^ p50_array_index_2053078 ^ p50_array_index_2053051 ^ p50_array_index_2053022 ^ p50_array_index_2052900 ^ p50_literal_2043912[p50_array_index_2052885] ^ p50_literal_2043910[p50_array_index_2052886] ^ p50_array_index_2052887;
  assign p51_array_index_2053258_comb = p50_literal_2043920[p50_res7__650];
  assign p51_res7__662_comb = p50_literal_2043910[p51_res7__660_comb] ^ p50_literal_2043912[p51_res7__658_comb] ^ p50_literal_2043914[p50_res7__656] ^ p50_literal_2043916[p50_res7__654] ^ p50_literal_2043918[p50_res7__652] ^ p51_array_index_2053258_comb ^ p50_res7__648 ^ p50_literal_2043923[p50_res7__646] ^ p50_res7__644 ^ p50_array_index_2053090 ^ p50_array_index_2053064 ^ p50_array_index_2053036 ^ p50_array_index_2052917 ^ p50_literal_2043912[p50_array_index_2052884] ^ p50_literal_2043910[p50_array_index_2052885] ^ p50_array_index_2052886;
  assign p51_res7__664_comb = p50_literal_2043910[p51_res7__662_comb] ^ p50_literal_2043912[p51_res7__660_comb] ^ p50_literal_2043914[p51_res7__658_comb] ^ p50_literal_2043916[p50_res7__656] ^ p50_literal_2043918[p50_res7__654] ^ p50_literal_2043920[p50_res7__652] ^ p50_res7__650 ^ p50_literal_2043923[p50_res7__648] ^ p50_res7__646 ^ p50_array_index_2053102 ^ p50_array_index_2053077 ^ p50_array_index_2053050 ^ p50_array_index_2053021 ^ p50_array_index_2052899 ^ p50_literal_2043910[p50_array_index_2052884] ^ p50_array_index_2052885;
  assign p51_res7__666_comb = p50_literal_2043910[p51_res7__664_comb] ^ p50_literal_2043912[p51_res7__662_comb] ^ p50_literal_2043914[p51_res7__660_comb] ^ p50_literal_2043916[p51_res7__658_comb] ^ p50_literal_2043918[p50_res7__656] ^ p50_literal_2043920[p50_res7__654] ^ p50_res7__652 ^ p50_literal_2043923[p50_res7__650] ^ p50_res7__648 ^ p51_array_index_2053237_comb ^ p50_array_index_2053089 ^ p50_array_index_2053063 ^ p50_array_index_2053035 ^ p50_array_index_2052916 ^ p50_literal_2043910[p50_array_index_2052883] ^ p50_array_index_2052884;
  assign p51_res7__668_comb = p50_literal_2043910[p51_res7__666_comb] ^ p50_literal_2043912[p51_res7__664_comb] ^ p50_literal_2043914[p51_res7__662_comb] ^ p50_literal_2043916[p51_res7__660_comb] ^ p50_literal_2043918[p51_res7__658_comb] ^ p50_literal_2043920[p50_res7__656] ^ p50_res7__654 ^ p50_literal_2043923[p50_res7__652] ^ p50_res7__650 ^ p51_array_index_2053248_comb ^ p50_array_index_2053101 ^ p50_array_index_2053076 ^ p50_array_index_2053049 ^ p50_array_index_2053020 ^ p50_array_index_2052898 ^ p50_array_index_2052883;
  assign p51_res7__670_comb = p50_literal_2043910[p51_res7__668_comb] ^ p50_literal_2043912[p51_res7__666_comb] ^ p50_literal_2043914[p51_res7__664_comb] ^ p50_literal_2043916[p51_res7__662_comb] ^ p50_literal_2043918[p51_res7__660_comb] ^ p50_literal_2043920[p51_res7__658_comb] ^ p50_res7__656 ^ p50_literal_2043923[p50_res7__654] ^ p50_res7__652 ^ p51_array_index_2053258_comb ^ p51_array_index_2053236_comb ^ p50_array_index_2053088 ^ p50_array_index_2053062 ^ p50_array_index_2053034 ^ p50_array_index_2052915 ^ p50_array_index_2052882;
  assign p51_res__20_comb = {p51_res7__670_comb, p51_res7__668_comb, p51_res7__666_comb, p51_res7__664_comb, p51_res7__662_comb, p51_res7__660_comb, p51_res7__658_comb, p50_res7__656, p50_res7__654, p50_res7__652, p50_res7__650, p50_res7__648, p50_res7__646, p50_res7__644, p50_res7__642, p50_res7__640};

  // Registers for pipe stage 51:
  reg [127:0] p51_encoded;
  reg [127:0] p51_bit_slice_2043893;
  reg [127:0] p51_bit_slice_2044018;
  reg [127:0] p51_k3;
  reg [127:0] p51_k2;
  reg [127:0] p51_k5;
  reg [127:0] p51_k4;
  reg [127:0] p51_xor_2052422;
  reg [127:0] p51_xor_2052866;
  reg [127:0] p51_res__20;
  reg [7:0] p52_literal_2043896[256];
  reg [7:0] p52_literal_2043910[256];
  reg [7:0] p52_literal_2043912[256];
  reg [7:0] p52_literal_2043914[256];
  reg [7:0] p52_literal_2043916[256];
  reg [7:0] p52_literal_2043918[256];
  reg [7:0] p52_literal_2043920[256];
  reg [7:0] p52_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p51_encoded <= p50_encoded;
    p51_bit_slice_2043893 <= p50_bit_slice_2043893;
    p51_bit_slice_2044018 <= p50_bit_slice_2044018;
    p51_k3 <= p50_k3;
    p51_k2 <= p50_k2;
    p51_k5 <= p50_k5;
    p51_k4 <= p50_k4;
    p51_xor_2052422 <= p50_xor_2052422;
    p51_xor_2052866 <= p50_xor_2052866;
    p51_res__20 <= p51_res__20_comb;
    p52_literal_2043896 <= p51_literal_2043896;
    p52_literal_2043910 <= p51_literal_2043910;
    p52_literal_2043912 <= p51_literal_2043912;
    p52_literal_2043914 <= p51_literal_2043914;
    p52_literal_2043916 <= p51_literal_2043916;
    p52_literal_2043918 <= p51_literal_2043918;
    p52_literal_2043920 <= p51_literal_2043920;
    p52_literal_2043923 <= p51_literal_2043923;
  end

  // ===== Pipe stage 52:
  wire [127:0] p52_xor_2053334_comb;
  wire [127:0] p52_addedKey__53_comb;
  wire [7:0] p52_array_index_2053350_comb;
  wire [7:0] p52_array_index_2053351_comb;
  wire [7:0] p52_array_index_2053352_comb;
  wire [7:0] p52_array_index_2053353_comb;
  wire [7:0] p52_array_index_2053354_comb;
  wire [7:0] p52_array_index_2053355_comb;
  wire [7:0] p52_array_index_2053357_comb;
  wire [7:0] p52_array_index_2053359_comb;
  wire [7:0] p52_array_index_2053360_comb;
  wire [7:0] p52_array_index_2053361_comb;
  wire [7:0] p52_array_index_2053362_comb;
  wire [7:0] p52_array_index_2053363_comb;
  wire [7:0] p52_array_index_2053364_comb;
  wire [7:0] p52_array_index_2053366_comb;
  wire [7:0] p52_array_index_2053367_comb;
  wire [7:0] p52_array_index_2053368_comb;
  wire [7:0] p52_array_index_2053369_comb;
  wire [7:0] p52_array_index_2053370_comb;
  wire [7:0] p52_array_index_2053371_comb;
  wire [7:0] p52_array_index_2053372_comb;
  wire [7:0] p52_array_index_2053374_comb;
  wire [7:0] p52_res7__672_comb;
  wire [7:0] p52_array_index_2053383_comb;
  wire [7:0] p52_array_index_2053384_comb;
  wire [7:0] p52_array_index_2053385_comb;
  wire [7:0] p52_array_index_2053386_comb;
  wire [7:0] p52_array_index_2053387_comb;
  wire [7:0] p52_array_index_2053388_comb;
  wire [7:0] p52_res7__674_comb;
  wire [7:0] p52_array_index_2053398_comb;
  wire [7:0] p52_array_index_2053399_comb;
  wire [7:0] p52_array_index_2053400_comb;
  wire [7:0] p52_array_index_2053401_comb;
  wire [7:0] p52_array_index_2053402_comb;
  wire [7:0] p52_res7__676_comb;
  wire [7:0] p52_array_index_2053412_comb;
  wire [7:0] p52_array_index_2053413_comb;
  wire [7:0] p52_array_index_2053414_comb;
  wire [7:0] p52_array_index_2053415_comb;
  wire [7:0] p52_array_index_2053416_comb;
  wire [7:0] p52_res7__678_comb;
  wire [7:0] p52_array_index_2053427_comb;
  wire [7:0] p52_array_index_2053428_comb;
  wire [7:0] p52_array_index_2053429_comb;
  wire [7:0] p52_array_index_2053430_comb;
  wire [7:0] p52_res7__680_comb;
  wire [7:0] p52_array_index_2053440_comb;
  wire [7:0] p52_array_index_2053441_comb;
  wire [7:0] p52_array_index_2053442_comb;
  wire [7:0] p52_array_index_2053443_comb;
  wire [7:0] p52_res7__682_comb;
  assign p52_xor_2053334_comb = p51_res__20 ^ p51_xor_2052422;
  assign p52_addedKey__53_comb = p52_xor_2053334_comb ^ 128'h88f8_9bc3_a479_73c7_94e7_89a3_c509_aa16;
  assign p52_array_index_2053350_comb = p51_literal_2043896[p52_addedKey__53_comb[127:120]];
  assign p52_array_index_2053351_comb = p51_literal_2043896[p52_addedKey__53_comb[119:112]];
  assign p52_array_index_2053352_comb = p51_literal_2043896[p52_addedKey__53_comb[111:104]];
  assign p52_array_index_2053353_comb = p51_literal_2043896[p52_addedKey__53_comb[103:96]];
  assign p52_array_index_2053354_comb = p51_literal_2043896[p52_addedKey__53_comb[95:88]];
  assign p52_array_index_2053355_comb = p51_literal_2043896[p52_addedKey__53_comb[87:80]];
  assign p52_array_index_2053357_comb = p51_literal_2043896[p52_addedKey__53_comb[71:64]];
  assign p52_array_index_2053359_comb = p51_literal_2043896[p52_addedKey__53_comb[55:48]];
  assign p52_array_index_2053360_comb = p51_literal_2043896[p52_addedKey__53_comb[47:40]];
  assign p52_array_index_2053361_comb = p51_literal_2043896[p52_addedKey__53_comb[39:32]];
  assign p52_array_index_2053362_comb = p51_literal_2043896[p52_addedKey__53_comb[31:24]];
  assign p52_array_index_2053363_comb = p51_literal_2043896[p52_addedKey__53_comb[23:16]];
  assign p52_array_index_2053364_comb = p51_literal_2043896[p52_addedKey__53_comb[15:8]];
  assign p52_array_index_2053366_comb = p51_literal_2043910[p52_array_index_2053350_comb];
  assign p52_array_index_2053367_comb = p51_literal_2043912[p52_array_index_2053351_comb];
  assign p52_array_index_2053368_comb = p51_literal_2043914[p52_array_index_2053352_comb];
  assign p52_array_index_2053369_comb = p51_literal_2043916[p52_array_index_2053353_comb];
  assign p52_array_index_2053370_comb = p51_literal_2043918[p52_array_index_2053354_comb];
  assign p52_array_index_2053371_comb = p51_literal_2043920[p52_array_index_2053355_comb];
  assign p52_array_index_2053372_comb = p51_literal_2043896[p52_addedKey__53_comb[79:72]];
  assign p52_array_index_2053374_comb = p51_literal_2043896[p52_addedKey__53_comb[63:56]];
  assign p52_res7__672_comb = p52_array_index_2053366_comb ^ p52_array_index_2053367_comb ^ p52_array_index_2053368_comb ^ p52_array_index_2053369_comb ^ p52_array_index_2053370_comb ^ p52_array_index_2053371_comb ^ p52_array_index_2053372_comb ^ p51_literal_2043923[p52_array_index_2053357_comb] ^ p52_array_index_2053374_comb ^ p51_literal_2043920[p52_array_index_2053359_comb] ^ p51_literal_2043918[p52_array_index_2053360_comb] ^ p51_literal_2043916[p52_array_index_2053361_comb] ^ p51_literal_2043914[p52_array_index_2053362_comb] ^ p51_literal_2043912[p52_array_index_2053363_comb] ^ p51_literal_2043910[p52_array_index_2053364_comb] ^ p51_literal_2043896[p52_addedKey__53_comb[7:0]];
  assign p52_array_index_2053383_comb = p51_literal_2043910[p52_res7__672_comb];
  assign p52_array_index_2053384_comb = p51_literal_2043912[p52_array_index_2053350_comb];
  assign p52_array_index_2053385_comb = p51_literal_2043914[p52_array_index_2053351_comb];
  assign p52_array_index_2053386_comb = p51_literal_2043916[p52_array_index_2053352_comb];
  assign p52_array_index_2053387_comb = p51_literal_2043918[p52_array_index_2053353_comb];
  assign p52_array_index_2053388_comb = p51_literal_2043920[p52_array_index_2053354_comb];
  assign p52_res7__674_comb = p52_array_index_2053383_comb ^ p52_array_index_2053384_comb ^ p52_array_index_2053385_comb ^ p52_array_index_2053386_comb ^ p52_array_index_2053387_comb ^ p52_array_index_2053388_comb ^ p52_array_index_2053355_comb ^ p51_literal_2043923[p52_array_index_2053372_comb] ^ p52_array_index_2053357_comb ^ p51_literal_2043920[p52_array_index_2053374_comb] ^ p51_literal_2043918[p52_array_index_2053359_comb] ^ p51_literal_2043916[p52_array_index_2053360_comb] ^ p51_literal_2043914[p52_array_index_2053361_comb] ^ p51_literal_2043912[p52_array_index_2053362_comb] ^ p51_literal_2043910[p52_array_index_2053363_comb] ^ p52_array_index_2053364_comb;
  assign p52_array_index_2053398_comb = p51_literal_2043912[p52_res7__672_comb];
  assign p52_array_index_2053399_comb = p51_literal_2043914[p52_array_index_2053350_comb];
  assign p52_array_index_2053400_comb = p51_literal_2043916[p52_array_index_2053351_comb];
  assign p52_array_index_2053401_comb = p51_literal_2043918[p52_array_index_2053352_comb];
  assign p52_array_index_2053402_comb = p51_literal_2043920[p52_array_index_2053353_comb];
  assign p52_res7__676_comb = p51_literal_2043910[p52_res7__674_comb] ^ p52_array_index_2053398_comb ^ p52_array_index_2053399_comb ^ p52_array_index_2053400_comb ^ p52_array_index_2053401_comb ^ p52_array_index_2053402_comb ^ p52_array_index_2053354_comb ^ p51_literal_2043923[p52_array_index_2053355_comb] ^ p52_array_index_2053372_comb ^ p51_literal_2043920[p52_array_index_2053357_comb] ^ p51_literal_2043918[p52_array_index_2053374_comb] ^ p51_literal_2043916[p52_array_index_2053359_comb] ^ p51_literal_2043914[p52_array_index_2053360_comb] ^ p51_literal_2043912[p52_array_index_2053361_comb] ^ p51_literal_2043910[p52_array_index_2053362_comb] ^ p52_array_index_2053363_comb;
  assign p52_array_index_2053412_comb = p51_literal_2043912[p52_res7__674_comb];
  assign p52_array_index_2053413_comb = p51_literal_2043914[p52_res7__672_comb];
  assign p52_array_index_2053414_comb = p51_literal_2043916[p52_array_index_2053350_comb];
  assign p52_array_index_2053415_comb = p51_literal_2043918[p52_array_index_2053351_comb];
  assign p52_array_index_2053416_comb = p51_literal_2043920[p52_array_index_2053352_comb];
  assign p52_res7__678_comb = p51_literal_2043910[p52_res7__676_comb] ^ p52_array_index_2053412_comb ^ p52_array_index_2053413_comb ^ p52_array_index_2053414_comb ^ p52_array_index_2053415_comb ^ p52_array_index_2053416_comb ^ p52_array_index_2053353_comb ^ p51_literal_2043923[p52_array_index_2053354_comb] ^ p52_array_index_2053355_comb ^ p51_literal_2043920[p52_array_index_2053372_comb] ^ p51_literal_2043918[p52_array_index_2053357_comb] ^ p51_literal_2043916[p52_array_index_2053374_comb] ^ p51_literal_2043914[p52_array_index_2053359_comb] ^ p51_literal_2043912[p52_array_index_2053360_comb] ^ p51_literal_2043910[p52_array_index_2053361_comb] ^ p52_array_index_2053362_comb;
  assign p52_array_index_2053427_comb = p51_literal_2043914[p52_res7__674_comb];
  assign p52_array_index_2053428_comb = p51_literal_2043916[p52_res7__672_comb];
  assign p52_array_index_2053429_comb = p51_literal_2043918[p52_array_index_2053350_comb];
  assign p52_array_index_2053430_comb = p51_literal_2043920[p52_array_index_2053351_comb];
  assign p52_res7__680_comb = p51_literal_2043910[p52_res7__678_comb] ^ p51_literal_2043912[p52_res7__676_comb] ^ p52_array_index_2053427_comb ^ p52_array_index_2053428_comb ^ p52_array_index_2053429_comb ^ p52_array_index_2053430_comb ^ p52_array_index_2053352_comb ^ p51_literal_2043923[p52_array_index_2053353_comb] ^ p52_array_index_2053354_comb ^ p52_array_index_2053371_comb ^ p51_literal_2043918[p52_array_index_2053372_comb] ^ p51_literal_2043916[p52_array_index_2053357_comb] ^ p51_literal_2043914[p52_array_index_2053374_comb] ^ p51_literal_2043912[p52_array_index_2053359_comb] ^ p51_literal_2043910[p52_array_index_2053360_comb] ^ p52_array_index_2053361_comb;
  assign p52_array_index_2053440_comb = p51_literal_2043914[p52_res7__676_comb];
  assign p52_array_index_2053441_comb = p51_literal_2043916[p52_res7__674_comb];
  assign p52_array_index_2053442_comb = p51_literal_2043918[p52_res7__672_comb];
  assign p52_array_index_2053443_comb = p51_literal_2043920[p52_array_index_2053350_comb];
  assign p52_res7__682_comb = p51_literal_2043910[p52_res7__680_comb] ^ p51_literal_2043912[p52_res7__678_comb] ^ p52_array_index_2053440_comb ^ p52_array_index_2053441_comb ^ p52_array_index_2053442_comb ^ p52_array_index_2053443_comb ^ p52_array_index_2053351_comb ^ p51_literal_2043923[p52_array_index_2053352_comb] ^ p52_array_index_2053353_comb ^ p52_array_index_2053388_comb ^ p51_literal_2043918[p52_array_index_2053355_comb] ^ p51_literal_2043916[p52_array_index_2053372_comb] ^ p51_literal_2043914[p52_array_index_2053357_comb] ^ p51_literal_2043912[p52_array_index_2053374_comb] ^ p51_literal_2043910[p52_array_index_2053359_comb] ^ p52_array_index_2053360_comb;

  // Registers for pipe stage 52:
  reg [127:0] p52_encoded;
  reg [127:0] p52_bit_slice_2043893;
  reg [127:0] p52_bit_slice_2044018;
  reg [127:0] p52_k3;
  reg [127:0] p52_k2;
  reg [127:0] p52_k5;
  reg [127:0] p52_k4;
  reg [127:0] p52_xor_2052866;
  reg [127:0] p52_xor_2053334;
  reg [7:0] p52_array_index_2053350;
  reg [7:0] p52_array_index_2053351;
  reg [7:0] p52_array_index_2053352;
  reg [7:0] p52_array_index_2053353;
  reg [7:0] p52_array_index_2053354;
  reg [7:0] p52_array_index_2053355;
  reg [7:0] p52_array_index_2053357;
  reg [7:0] p52_array_index_2053359;
  reg [7:0] p52_array_index_2053366;
  reg [7:0] p52_array_index_2053367;
  reg [7:0] p52_array_index_2053368;
  reg [7:0] p52_array_index_2053369;
  reg [7:0] p52_array_index_2053370;
  reg [7:0] p52_array_index_2053372;
  reg [7:0] p52_array_index_2053374;
  reg [7:0] p52_res7__672;
  reg [7:0] p52_array_index_2053383;
  reg [7:0] p52_array_index_2053384;
  reg [7:0] p52_array_index_2053385;
  reg [7:0] p52_array_index_2053386;
  reg [7:0] p52_array_index_2053387;
  reg [7:0] p52_res7__674;
  reg [7:0] p52_array_index_2053398;
  reg [7:0] p52_array_index_2053399;
  reg [7:0] p52_array_index_2053400;
  reg [7:0] p52_array_index_2053401;
  reg [7:0] p52_array_index_2053402;
  reg [7:0] p52_res7__676;
  reg [7:0] p52_array_index_2053412;
  reg [7:0] p52_array_index_2053413;
  reg [7:0] p52_array_index_2053414;
  reg [7:0] p52_array_index_2053415;
  reg [7:0] p52_array_index_2053416;
  reg [7:0] p52_res7__678;
  reg [7:0] p52_array_index_2053427;
  reg [7:0] p52_array_index_2053428;
  reg [7:0] p52_array_index_2053429;
  reg [7:0] p52_array_index_2053430;
  reg [7:0] p52_res7__680;
  reg [7:0] p52_array_index_2053440;
  reg [7:0] p52_array_index_2053441;
  reg [7:0] p52_array_index_2053442;
  reg [7:0] p52_array_index_2053443;
  reg [7:0] p52_res7__682;
  reg [7:0] p53_literal_2043896[256];
  reg [7:0] p53_literal_2043910[256];
  reg [7:0] p53_literal_2043912[256];
  reg [7:0] p53_literal_2043914[256];
  reg [7:0] p53_literal_2043916[256];
  reg [7:0] p53_literal_2043918[256];
  reg [7:0] p53_literal_2043920[256];
  reg [7:0] p53_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p52_encoded <= p51_encoded;
    p52_bit_slice_2043893 <= p51_bit_slice_2043893;
    p52_bit_slice_2044018 <= p51_bit_slice_2044018;
    p52_k3 <= p51_k3;
    p52_k2 <= p51_k2;
    p52_k5 <= p51_k5;
    p52_k4 <= p51_k4;
    p52_xor_2052866 <= p51_xor_2052866;
    p52_xor_2053334 <= p52_xor_2053334_comb;
    p52_array_index_2053350 <= p52_array_index_2053350_comb;
    p52_array_index_2053351 <= p52_array_index_2053351_comb;
    p52_array_index_2053352 <= p52_array_index_2053352_comb;
    p52_array_index_2053353 <= p52_array_index_2053353_comb;
    p52_array_index_2053354 <= p52_array_index_2053354_comb;
    p52_array_index_2053355 <= p52_array_index_2053355_comb;
    p52_array_index_2053357 <= p52_array_index_2053357_comb;
    p52_array_index_2053359 <= p52_array_index_2053359_comb;
    p52_array_index_2053366 <= p52_array_index_2053366_comb;
    p52_array_index_2053367 <= p52_array_index_2053367_comb;
    p52_array_index_2053368 <= p52_array_index_2053368_comb;
    p52_array_index_2053369 <= p52_array_index_2053369_comb;
    p52_array_index_2053370 <= p52_array_index_2053370_comb;
    p52_array_index_2053372 <= p52_array_index_2053372_comb;
    p52_array_index_2053374 <= p52_array_index_2053374_comb;
    p52_res7__672 <= p52_res7__672_comb;
    p52_array_index_2053383 <= p52_array_index_2053383_comb;
    p52_array_index_2053384 <= p52_array_index_2053384_comb;
    p52_array_index_2053385 <= p52_array_index_2053385_comb;
    p52_array_index_2053386 <= p52_array_index_2053386_comb;
    p52_array_index_2053387 <= p52_array_index_2053387_comb;
    p52_res7__674 <= p52_res7__674_comb;
    p52_array_index_2053398 <= p52_array_index_2053398_comb;
    p52_array_index_2053399 <= p52_array_index_2053399_comb;
    p52_array_index_2053400 <= p52_array_index_2053400_comb;
    p52_array_index_2053401 <= p52_array_index_2053401_comb;
    p52_array_index_2053402 <= p52_array_index_2053402_comb;
    p52_res7__676 <= p52_res7__676_comb;
    p52_array_index_2053412 <= p52_array_index_2053412_comb;
    p52_array_index_2053413 <= p52_array_index_2053413_comb;
    p52_array_index_2053414 <= p52_array_index_2053414_comb;
    p52_array_index_2053415 <= p52_array_index_2053415_comb;
    p52_array_index_2053416 <= p52_array_index_2053416_comb;
    p52_res7__678 <= p52_res7__678_comb;
    p52_array_index_2053427 <= p52_array_index_2053427_comb;
    p52_array_index_2053428 <= p52_array_index_2053428_comb;
    p52_array_index_2053429 <= p52_array_index_2053429_comb;
    p52_array_index_2053430 <= p52_array_index_2053430_comb;
    p52_res7__680 <= p52_res7__680_comb;
    p52_array_index_2053440 <= p52_array_index_2053440_comb;
    p52_array_index_2053441 <= p52_array_index_2053441_comb;
    p52_array_index_2053442 <= p52_array_index_2053442_comb;
    p52_array_index_2053443 <= p52_array_index_2053443_comb;
    p52_res7__682 <= p52_res7__682_comb;
    p53_literal_2043896 <= p52_literal_2043896;
    p53_literal_2043910 <= p52_literal_2043910;
    p53_literal_2043912 <= p52_literal_2043912;
    p53_literal_2043914 <= p52_literal_2043914;
    p53_literal_2043916 <= p52_literal_2043916;
    p53_literal_2043918 <= p52_literal_2043918;
    p53_literal_2043920 <= p52_literal_2043920;
    p53_literal_2043923 <= p52_literal_2043923;
  end

  // ===== Pipe stage 53:
  wire [7:0] p53_array_index_2053576_comb;
  wire [7:0] p53_array_index_2053577_comb;
  wire [7:0] p53_array_index_2053578_comb;
  wire [7:0] p53_res7__684_comb;
  wire [7:0] p53_array_index_2053588_comb;
  wire [7:0] p53_array_index_2053589_comb;
  wire [7:0] p53_array_index_2053590_comb;
  wire [7:0] p53_res7__686_comb;
  wire [7:0] p53_array_index_2053601_comb;
  wire [7:0] p53_array_index_2053602_comb;
  wire [7:0] p53_res7__688_comb;
  wire [7:0] p53_array_index_2053612_comb;
  wire [7:0] p53_array_index_2053613_comb;
  wire [7:0] p53_res7__690_comb;
  wire [7:0] p53_array_index_2053624_comb;
  wire [7:0] p53_res7__692_comb;
  wire [7:0] p53_array_index_2053634_comb;
  wire [7:0] p53_res7__694_comb;
  wire [7:0] p53_res7__696_comb;
  assign p53_array_index_2053576_comb = p52_literal_2043916[p52_res7__676];
  assign p53_array_index_2053577_comb = p52_literal_2043918[p52_res7__674];
  assign p53_array_index_2053578_comb = p52_literal_2043920[p52_res7__672];
  assign p53_res7__684_comb = p52_literal_2043910[p52_res7__682] ^ p52_literal_2043912[p52_res7__680] ^ p52_literal_2043914[p52_res7__678] ^ p53_array_index_2053576_comb ^ p53_array_index_2053577_comb ^ p53_array_index_2053578_comb ^ p52_array_index_2053350 ^ p52_literal_2043923[p52_array_index_2053351] ^ p52_array_index_2053352 ^ p52_array_index_2053402 ^ p52_array_index_2053370 ^ p52_literal_2043916[p52_array_index_2053355] ^ p52_literal_2043914[p52_array_index_2053372] ^ p52_literal_2043912[p52_array_index_2053357] ^ p52_literal_2043910[p52_array_index_2053374] ^ p52_array_index_2053359;
  assign p53_array_index_2053588_comb = p52_literal_2043916[p52_res7__678];
  assign p53_array_index_2053589_comb = p52_literal_2043918[p52_res7__676];
  assign p53_array_index_2053590_comb = p52_literal_2043920[p52_res7__674];
  assign p53_res7__686_comb = p52_literal_2043910[p53_res7__684_comb] ^ p52_literal_2043912[p52_res7__682] ^ p52_literal_2043914[p52_res7__680] ^ p53_array_index_2053588_comb ^ p53_array_index_2053589_comb ^ p53_array_index_2053590_comb ^ p52_res7__672 ^ p52_literal_2043923[p52_array_index_2053350] ^ p52_array_index_2053351 ^ p52_array_index_2053416 ^ p52_array_index_2053387 ^ p52_literal_2043916[p52_array_index_2053354] ^ p52_literal_2043914[p52_array_index_2053355] ^ p52_literal_2043912[p52_array_index_2053372] ^ p52_literal_2043910[p52_array_index_2053357] ^ p52_array_index_2053374;
  assign p53_array_index_2053601_comb = p52_literal_2043918[p52_res7__678];
  assign p53_array_index_2053602_comb = p52_literal_2043920[p52_res7__676];
  assign p53_res7__688_comb = p52_literal_2043910[p53_res7__686_comb] ^ p52_literal_2043912[p53_res7__684_comb] ^ p52_literal_2043914[p52_res7__682] ^ p52_literal_2043916[p52_res7__680] ^ p53_array_index_2053601_comb ^ p53_array_index_2053602_comb ^ p52_res7__674 ^ p52_literal_2043923[p52_res7__672] ^ p52_array_index_2053350 ^ p52_array_index_2053430 ^ p52_array_index_2053401 ^ p52_array_index_2053369 ^ p52_literal_2043914[p52_array_index_2053354] ^ p52_literal_2043912[p52_array_index_2053355] ^ p52_literal_2043910[p52_array_index_2053372] ^ p52_array_index_2053357;
  assign p53_array_index_2053612_comb = p52_literal_2043918[p52_res7__680];
  assign p53_array_index_2053613_comb = p52_literal_2043920[p52_res7__678];
  assign p53_res7__690_comb = p52_literal_2043910[p53_res7__688_comb] ^ p52_literal_2043912[p53_res7__686_comb] ^ p52_literal_2043914[p53_res7__684_comb] ^ p52_literal_2043916[p52_res7__682] ^ p53_array_index_2053612_comb ^ p53_array_index_2053613_comb ^ p52_res7__676 ^ p52_literal_2043923[p52_res7__674] ^ p52_res7__672 ^ p52_array_index_2053443 ^ p52_array_index_2053415 ^ p52_array_index_2053386 ^ p52_literal_2043914[p52_array_index_2053353] ^ p52_literal_2043912[p52_array_index_2053354] ^ p52_literal_2043910[p52_array_index_2053355] ^ p52_array_index_2053372;
  assign p53_array_index_2053624_comb = p52_literal_2043920[p52_res7__680];
  assign p53_res7__692_comb = p52_literal_2043910[p53_res7__690_comb] ^ p52_literal_2043912[p53_res7__688_comb] ^ p52_literal_2043914[p53_res7__686_comb] ^ p52_literal_2043916[p53_res7__684_comb] ^ p52_literal_2043918[p52_res7__682] ^ p53_array_index_2053624_comb ^ p52_res7__678 ^ p52_literal_2043923[p52_res7__676] ^ p52_res7__674 ^ p53_array_index_2053578_comb ^ p52_array_index_2053429 ^ p52_array_index_2053400 ^ p52_array_index_2053368 ^ p52_literal_2043912[p52_array_index_2053353] ^ p52_literal_2043910[p52_array_index_2053354] ^ p52_array_index_2053355;
  assign p53_array_index_2053634_comb = p52_literal_2043920[p52_res7__682];
  assign p53_res7__694_comb = p52_literal_2043910[p53_res7__692_comb] ^ p52_literal_2043912[p53_res7__690_comb] ^ p52_literal_2043914[p53_res7__688_comb] ^ p52_literal_2043916[p53_res7__686_comb] ^ p52_literal_2043918[p53_res7__684_comb] ^ p53_array_index_2053634_comb ^ p52_res7__680 ^ p52_literal_2043923[p52_res7__678] ^ p52_res7__676 ^ p53_array_index_2053590_comb ^ p52_array_index_2053442 ^ p52_array_index_2053414 ^ p52_array_index_2053385 ^ p52_literal_2043912[p52_array_index_2053352] ^ p52_literal_2043910[p52_array_index_2053353] ^ p52_array_index_2053354;
  assign p53_res7__696_comb = p52_literal_2043910[p53_res7__694_comb] ^ p52_literal_2043912[p53_res7__692_comb] ^ p52_literal_2043914[p53_res7__690_comb] ^ p52_literal_2043916[p53_res7__688_comb] ^ p52_literal_2043918[p53_res7__686_comb] ^ p52_literal_2043920[p53_res7__684_comb] ^ p52_res7__682 ^ p52_literal_2043923[p52_res7__680] ^ p52_res7__678 ^ p53_array_index_2053602_comb ^ p53_array_index_2053577_comb ^ p52_array_index_2053428 ^ p52_array_index_2053399 ^ p52_array_index_2053367 ^ p52_literal_2043910[p52_array_index_2053352] ^ p52_array_index_2053353;

  // Registers for pipe stage 53:
  reg [127:0] p53_encoded;
  reg [127:0] p53_bit_slice_2043893;
  reg [127:0] p53_bit_slice_2044018;
  reg [127:0] p53_k3;
  reg [127:0] p53_k2;
  reg [127:0] p53_k5;
  reg [127:0] p53_k4;
  reg [127:0] p53_xor_2052866;
  reg [127:0] p53_xor_2053334;
  reg [7:0] p53_array_index_2053350;
  reg [7:0] p53_array_index_2053351;
  reg [7:0] p53_array_index_2053352;
  reg [7:0] p53_array_index_2053366;
  reg [7:0] p53_res7__672;
  reg [7:0] p53_array_index_2053383;
  reg [7:0] p53_array_index_2053384;
  reg [7:0] p53_res7__674;
  reg [7:0] p53_array_index_2053398;
  reg [7:0] p53_res7__676;
  reg [7:0] p53_array_index_2053412;
  reg [7:0] p53_array_index_2053413;
  reg [7:0] p53_res7__678;
  reg [7:0] p53_array_index_2053427;
  reg [7:0] p53_res7__680;
  reg [7:0] p53_array_index_2053440;
  reg [7:0] p53_array_index_2053441;
  reg [7:0] p53_res7__682;
  reg [7:0] p53_array_index_2053576;
  reg [7:0] p53_res7__684;
  reg [7:0] p53_array_index_2053588;
  reg [7:0] p53_array_index_2053589;
  reg [7:0] p53_res7__686;
  reg [7:0] p53_array_index_2053601;
  reg [7:0] p53_res7__688;
  reg [7:0] p53_array_index_2053612;
  reg [7:0] p53_array_index_2053613;
  reg [7:0] p53_res7__690;
  reg [7:0] p53_array_index_2053624;
  reg [7:0] p53_res7__692;
  reg [7:0] p53_array_index_2053634;
  reg [7:0] p53_res7__694;
  reg [7:0] p53_res7__696;
  reg [7:0] p54_literal_2043896[256];
  reg [7:0] p54_literal_2043910[256];
  reg [7:0] p54_literal_2043912[256];
  reg [7:0] p54_literal_2043914[256];
  reg [7:0] p54_literal_2043916[256];
  reg [7:0] p54_literal_2043918[256];
  reg [7:0] p54_literal_2043920[256];
  reg [7:0] p54_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p53_encoded <= p52_encoded;
    p53_bit_slice_2043893 <= p52_bit_slice_2043893;
    p53_bit_slice_2044018 <= p52_bit_slice_2044018;
    p53_k3 <= p52_k3;
    p53_k2 <= p52_k2;
    p53_k5 <= p52_k5;
    p53_k4 <= p52_k4;
    p53_xor_2052866 <= p52_xor_2052866;
    p53_xor_2053334 <= p52_xor_2053334;
    p53_array_index_2053350 <= p52_array_index_2053350;
    p53_array_index_2053351 <= p52_array_index_2053351;
    p53_array_index_2053352 <= p52_array_index_2053352;
    p53_array_index_2053366 <= p52_array_index_2053366;
    p53_res7__672 <= p52_res7__672;
    p53_array_index_2053383 <= p52_array_index_2053383;
    p53_array_index_2053384 <= p52_array_index_2053384;
    p53_res7__674 <= p52_res7__674;
    p53_array_index_2053398 <= p52_array_index_2053398;
    p53_res7__676 <= p52_res7__676;
    p53_array_index_2053412 <= p52_array_index_2053412;
    p53_array_index_2053413 <= p52_array_index_2053413;
    p53_res7__678 <= p52_res7__678;
    p53_array_index_2053427 <= p52_array_index_2053427;
    p53_res7__680 <= p52_res7__680;
    p53_array_index_2053440 <= p52_array_index_2053440;
    p53_array_index_2053441 <= p52_array_index_2053441;
    p53_res7__682 <= p52_res7__682;
    p53_array_index_2053576 <= p53_array_index_2053576_comb;
    p53_res7__684 <= p53_res7__684_comb;
    p53_array_index_2053588 <= p53_array_index_2053588_comb;
    p53_array_index_2053589 <= p53_array_index_2053589_comb;
    p53_res7__686 <= p53_res7__686_comb;
    p53_array_index_2053601 <= p53_array_index_2053601_comb;
    p53_res7__688 <= p53_res7__688_comb;
    p53_array_index_2053612 <= p53_array_index_2053612_comb;
    p53_array_index_2053613 <= p53_array_index_2053613_comb;
    p53_res7__690 <= p53_res7__690_comb;
    p53_array_index_2053624 <= p53_array_index_2053624_comb;
    p53_res7__692 <= p53_res7__692_comb;
    p53_array_index_2053634 <= p53_array_index_2053634_comb;
    p53_res7__694 <= p53_res7__694_comb;
    p53_res7__696 <= p53_res7__696_comb;
    p54_literal_2043896 <= p53_literal_2043896;
    p54_literal_2043910 <= p53_literal_2043910;
    p54_literal_2043912 <= p53_literal_2043912;
    p54_literal_2043914 <= p53_literal_2043914;
    p54_literal_2043916 <= p53_literal_2043916;
    p54_literal_2043918 <= p53_literal_2043918;
    p54_literal_2043920 <= p53_literal_2043920;
    p54_literal_2043923 <= p53_literal_2043923;
  end

  // ===== Pipe stage 54:
  wire [7:0] p54_res7__698_comb;
  wire [7:0] p54_res7__700_comb;
  wire [7:0] p54_res7__702_comb;
  wire [127:0] p54_res__21_comb;
  wire [127:0] p54_xor_2053774_comb;
  wire [127:0] p54_addedKey__54_comb;
  wire [7:0] p54_array_index_2053790_comb;
  wire [7:0] p54_array_index_2053791_comb;
  wire [7:0] p54_array_index_2053792_comb;
  wire [7:0] p54_array_index_2053793_comb;
  wire [7:0] p54_array_index_2053794_comb;
  wire [7:0] p54_array_index_2053795_comb;
  wire [7:0] p54_array_index_2053797_comb;
  wire [7:0] p54_array_index_2053799_comb;
  wire [7:0] p54_array_index_2053800_comb;
  wire [7:0] p54_array_index_2053801_comb;
  wire [7:0] p54_array_index_2053802_comb;
  wire [7:0] p54_array_index_2053803_comb;
  wire [7:0] p54_array_index_2053804_comb;
  wire [7:0] p54_array_index_2053806_comb;
  wire [7:0] p54_array_index_2053807_comb;
  wire [7:0] p54_array_index_2053808_comb;
  wire [7:0] p54_array_index_2053809_comb;
  wire [7:0] p54_array_index_2053810_comb;
  wire [7:0] p54_array_index_2053811_comb;
  wire [7:0] p54_array_index_2053812_comb;
  wire [7:0] p54_array_index_2053814_comb;
  wire [7:0] p54_res7__704_comb;
  wire [7:0] p54_array_index_2053823_comb;
  wire [7:0] p54_array_index_2053824_comb;
  wire [7:0] p54_array_index_2053825_comb;
  wire [7:0] p54_array_index_2053826_comb;
  wire [7:0] p54_array_index_2053827_comb;
  wire [7:0] p54_array_index_2053828_comb;
  wire [7:0] p54_res7__706_comb;
  wire [7:0] p54_array_index_2053838_comb;
  wire [7:0] p54_array_index_2053839_comb;
  wire [7:0] p54_array_index_2053840_comb;
  wire [7:0] p54_array_index_2053841_comb;
  wire [7:0] p54_array_index_2053842_comb;
  wire [7:0] p54_res7__708_comb;
  assign p54_res7__698_comb = p53_literal_2043910[p53_res7__696] ^ p53_literal_2043912[p53_res7__694] ^ p53_literal_2043914[p53_res7__692] ^ p53_literal_2043916[p53_res7__690] ^ p53_literal_2043918[p53_res7__688] ^ p53_literal_2043920[p53_res7__686] ^ p53_res7__684 ^ p53_literal_2043923[p53_res7__682] ^ p53_res7__680 ^ p53_array_index_2053613 ^ p53_array_index_2053589 ^ p53_array_index_2053441 ^ p53_array_index_2053413 ^ p53_array_index_2053384 ^ p53_literal_2043910[p53_array_index_2053351] ^ p53_array_index_2053352;
  assign p54_res7__700_comb = p53_literal_2043910[p54_res7__698_comb] ^ p53_literal_2043912[p53_res7__696] ^ p53_literal_2043914[p53_res7__694] ^ p53_literal_2043916[p53_res7__692] ^ p53_literal_2043918[p53_res7__690] ^ p53_literal_2043920[p53_res7__688] ^ p53_res7__686 ^ p53_literal_2043923[p53_res7__684] ^ p53_res7__682 ^ p53_array_index_2053624 ^ p53_array_index_2053601 ^ p53_array_index_2053576 ^ p53_array_index_2053427 ^ p53_array_index_2053398 ^ p53_array_index_2053366 ^ p53_array_index_2053351;
  assign p54_res7__702_comb = p53_literal_2043910[p54_res7__700_comb] ^ p53_literal_2043912[p54_res7__698_comb] ^ p53_literal_2043914[p53_res7__696] ^ p53_literal_2043916[p53_res7__694] ^ p53_literal_2043918[p53_res7__692] ^ p53_literal_2043920[p53_res7__690] ^ p53_res7__688 ^ p53_literal_2043923[p53_res7__686] ^ p53_res7__684 ^ p53_array_index_2053634 ^ p53_array_index_2053612 ^ p53_array_index_2053588 ^ p53_array_index_2053440 ^ p53_array_index_2053412 ^ p53_array_index_2053383 ^ p53_array_index_2053350;
  assign p54_res__21_comb = {p54_res7__702_comb, p54_res7__700_comb, p54_res7__698_comb, p53_res7__696, p53_res7__694, p53_res7__692, p53_res7__690, p53_res7__688, p53_res7__686, p53_res7__684, p53_res7__682, p53_res7__680, p53_res7__678, p53_res7__676, p53_res7__674, p53_res7__672};
  assign p54_xor_2053774_comb = p54_res__21_comb ^ p53_xor_2052866;
  assign p54_addedKey__54_comb = p54_xor_2053774_comb ^ 128'he65a_edb1_c831_097f_c9c0_34b3_188d_3e17;
  assign p54_array_index_2053790_comb = p53_literal_2043896[p54_addedKey__54_comb[127:120]];
  assign p54_array_index_2053791_comb = p53_literal_2043896[p54_addedKey__54_comb[119:112]];
  assign p54_array_index_2053792_comb = p53_literal_2043896[p54_addedKey__54_comb[111:104]];
  assign p54_array_index_2053793_comb = p53_literal_2043896[p54_addedKey__54_comb[103:96]];
  assign p54_array_index_2053794_comb = p53_literal_2043896[p54_addedKey__54_comb[95:88]];
  assign p54_array_index_2053795_comb = p53_literal_2043896[p54_addedKey__54_comb[87:80]];
  assign p54_array_index_2053797_comb = p53_literal_2043896[p54_addedKey__54_comb[71:64]];
  assign p54_array_index_2053799_comb = p53_literal_2043896[p54_addedKey__54_comb[55:48]];
  assign p54_array_index_2053800_comb = p53_literal_2043896[p54_addedKey__54_comb[47:40]];
  assign p54_array_index_2053801_comb = p53_literal_2043896[p54_addedKey__54_comb[39:32]];
  assign p54_array_index_2053802_comb = p53_literal_2043896[p54_addedKey__54_comb[31:24]];
  assign p54_array_index_2053803_comb = p53_literal_2043896[p54_addedKey__54_comb[23:16]];
  assign p54_array_index_2053804_comb = p53_literal_2043896[p54_addedKey__54_comb[15:8]];
  assign p54_array_index_2053806_comb = p53_literal_2043910[p54_array_index_2053790_comb];
  assign p54_array_index_2053807_comb = p53_literal_2043912[p54_array_index_2053791_comb];
  assign p54_array_index_2053808_comb = p53_literal_2043914[p54_array_index_2053792_comb];
  assign p54_array_index_2053809_comb = p53_literal_2043916[p54_array_index_2053793_comb];
  assign p54_array_index_2053810_comb = p53_literal_2043918[p54_array_index_2053794_comb];
  assign p54_array_index_2053811_comb = p53_literal_2043920[p54_array_index_2053795_comb];
  assign p54_array_index_2053812_comb = p53_literal_2043896[p54_addedKey__54_comb[79:72]];
  assign p54_array_index_2053814_comb = p53_literal_2043896[p54_addedKey__54_comb[63:56]];
  assign p54_res7__704_comb = p54_array_index_2053806_comb ^ p54_array_index_2053807_comb ^ p54_array_index_2053808_comb ^ p54_array_index_2053809_comb ^ p54_array_index_2053810_comb ^ p54_array_index_2053811_comb ^ p54_array_index_2053812_comb ^ p53_literal_2043923[p54_array_index_2053797_comb] ^ p54_array_index_2053814_comb ^ p53_literal_2043920[p54_array_index_2053799_comb] ^ p53_literal_2043918[p54_array_index_2053800_comb] ^ p53_literal_2043916[p54_array_index_2053801_comb] ^ p53_literal_2043914[p54_array_index_2053802_comb] ^ p53_literal_2043912[p54_array_index_2053803_comb] ^ p53_literal_2043910[p54_array_index_2053804_comb] ^ p53_literal_2043896[p54_addedKey__54_comb[7:0]];
  assign p54_array_index_2053823_comb = p53_literal_2043910[p54_res7__704_comb];
  assign p54_array_index_2053824_comb = p53_literal_2043912[p54_array_index_2053790_comb];
  assign p54_array_index_2053825_comb = p53_literal_2043914[p54_array_index_2053791_comb];
  assign p54_array_index_2053826_comb = p53_literal_2043916[p54_array_index_2053792_comb];
  assign p54_array_index_2053827_comb = p53_literal_2043918[p54_array_index_2053793_comb];
  assign p54_array_index_2053828_comb = p53_literal_2043920[p54_array_index_2053794_comb];
  assign p54_res7__706_comb = p54_array_index_2053823_comb ^ p54_array_index_2053824_comb ^ p54_array_index_2053825_comb ^ p54_array_index_2053826_comb ^ p54_array_index_2053827_comb ^ p54_array_index_2053828_comb ^ p54_array_index_2053795_comb ^ p53_literal_2043923[p54_array_index_2053812_comb] ^ p54_array_index_2053797_comb ^ p53_literal_2043920[p54_array_index_2053814_comb] ^ p53_literal_2043918[p54_array_index_2053799_comb] ^ p53_literal_2043916[p54_array_index_2053800_comb] ^ p53_literal_2043914[p54_array_index_2053801_comb] ^ p53_literal_2043912[p54_array_index_2053802_comb] ^ p53_literal_2043910[p54_array_index_2053803_comb] ^ p54_array_index_2053804_comb;
  assign p54_array_index_2053838_comb = p53_literal_2043912[p54_res7__704_comb];
  assign p54_array_index_2053839_comb = p53_literal_2043914[p54_array_index_2053790_comb];
  assign p54_array_index_2053840_comb = p53_literal_2043916[p54_array_index_2053791_comb];
  assign p54_array_index_2053841_comb = p53_literal_2043918[p54_array_index_2053792_comb];
  assign p54_array_index_2053842_comb = p53_literal_2043920[p54_array_index_2053793_comb];
  assign p54_res7__708_comb = p53_literal_2043910[p54_res7__706_comb] ^ p54_array_index_2053838_comb ^ p54_array_index_2053839_comb ^ p54_array_index_2053840_comb ^ p54_array_index_2053841_comb ^ p54_array_index_2053842_comb ^ p54_array_index_2053794_comb ^ p53_literal_2043923[p54_array_index_2053795_comb] ^ p54_array_index_2053812_comb ^ p53_literal_2043920[p54_array_index_2053797_comb] ^ p53_literal_2043918[p54_array_index_2053814_comb] ^ p53_literal_2043916[p54_array_index_2053799_comb] ^ p53_literal_2043914[p54_array_index_2053800_comb] ^ p53_literal_2043912[p54_array_index_2053801_comb] ^ p53_literal_2043910[p54_array_index_2053802_comb] ^ p54_array_index_2053803_comb;

  // Registers for pipe stage 54:
  reg [127:0] p54_encoded;
  reg [127:0] p54_bit_slice_2043893;
  reg [127:0] p54_bit_slice_2044018;
  reg [127:0] p54_k3;
  reg [127:0] p54_k2;
  reg [127:0] p54_k5;
  reg [127:0] p54_k4;
  reg [127:0] p54_xor_2053334;
  reg [127:0] p54_xor_2053774;
  reg [7:0] p54_array_index_2053790;
  reg [7:0] p54_array_index_2053791;
  reg [7:0] p54_array_index_2053792;
  reg [7:0] p54_array_index_2053793;
  reg [7:0] p54_array_index_2053794;
  reg [7:0] p54_array_index_2053795;
  reg [7:0] p54_array_index_2053797;
  reg [7:0] p54_array_index_2053799;
  reg [7:0] p54_array_index_2053800;
  reg [7:0] p54_array_index_2053801;
  reg [7:0] p54_array_index_2053802;
  reg [7:0] p54_array_index_2053806;
  reg [7:0] p54_array_index_2053807;
  reg [7:0] p54_array_index_2053808;
  reg [7:0] p54_array_index_2053809;
  reg [7:0] p54_array_index_2053810;
  reg [7:0] p54_array_index_2053811;
  reg [7:0] p54_array_index_2053812;
  reg [7:0] p54_array_index_2053814;
  reg [7:0] p54_res7__704;
  reg [7:0] p54_array_index_2053823;
  reg [7:0] p54_array_index_2053824;
  reg [7:0] p54_array_index_2053825;
  reg [7:0] p54_array_index_2053826;
  reg [7:0] p54_array_index_2053827;
  reg [7:0] p54_array_index_2053828;
  reg [7:0] p54_res7__706;
  reg [7:0] p54_array_index_2053838;
  reg [7:0] p54_array_index_2053839;
  reg [7:0] p54_array_index_2053840;
  reg [7:0] p54_array_index_2053841;
  reg [7:0] p54_array_index_2053842;
  reg [7:0] p54_res7__708;
  reg [7:0] p55_literal_2043896[256];
  reg [7:0] p55_literal_2043910[256];
  reg [7:0] p55_literal_2043912[256];
  reg [7:0] p55_literal_2043914[256];
  reg [7:0] p55_literal_2043916[256];
  reg [7:0] p55_literal_2043918[256];
  reg [7:0] p55_literal_2043920[256];
  reg [7:0] p55_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p54_encoded <= p53_encoded;
    p54_bit_slice_2043893 <= p53_bit_slice_2043893;
    p54_bit_slice_2044018 <= p53_bit_slice_2044018;
    p54_k3 <= p53_k3;
    p54_k2 <= p53_k2;
    p54_k5 <= p53_k5;
    p54_k4 <= p53_k4;
    p54_xor_2053334 <= p53_xor_2053334;
    p54_xor_2053774 <= p54_xor_2053774_comb;
    p54_array_index_2053790 <= p54_array_index_2053790_comb;
    p54_array_index_2053791 <= p54_array_index_2053791_comb;
    p54_array_index_2053792 <= p54_array_index_2053792_comb;
    p54_array_index_2053793 <= p54_array_index_2053793_comb;
    p54_array_index_2053794 <= p54_array_index_2053794_comb;
    p54_array_index_2053795 <= p54_array_index_2053795_comb;
    p54_array_index_2053797 <= p54_array_index_2053797_comb;
    p54_array_index_2053799 <= p54_array_index_2053799_comb;
    p54_array_index_2053800 <= p54_array_index_2053800_comb;
    p54_array_index_2053801 <= p54_array_index_2053801_comb;
    p54_array_index_2053802 <= p54_array_index_2053802_comb;
    p54_array_index_2053806 <= p54_array_index_2053806_comb;
    p54_array_index_2053807 <= p54_array_index_2053807_comb;
    p54_array_index_2053808 <= p54_array_index_2053808_comb;
    p54_array_index_2053809 <= p54_array_index_2053809_comb;
    p54_array_index_2053810 <= p54_array_index_2053810_comb;
    p54_array_index_2053811 <= p54_array_index_2053811_comb;
    p54_array_index_2053812 <= p54_array_index_2053812_comb;
    p54_array_index_2053814 <= p54_array_index_2053814_comb;
    p54_res7__704 <= p54_res7__704_comb;
    p54_array_index_2053823 <= p54_array_index_2053823_comb;
    p54_array_index_2053824 <= p54_array_index_2053824_comb;
    p54_array_index_2053825 <= p54_array_index_2053825_comb;
    p54_array_index_2053826 <= p54_array_index_2053826_comb;
    p54_array_index_2053827 <= p54_array_index_2053827_comb;
    p54_array_index_2053828 <= p54_array_index_2053828_comb;
    p54_res7__706 <= p54_res7__706_comb;
    p54_array_index_2053838 <= p54_array_index_2053838_comb;
    p54_array_index_2053839 <= p54_array_index_2053839_comb;
    p54_array_index_2053840 <= p54_array_index_2053840_comb;
    p54_array_index_2053841 <= p54_array_index_2053841_comb;
    p54_array_index_2053842 <= p54_array_index_2053842_comb;
    p54_res7__708 <= p54_res7__708_comb;
    p55_literal_2043896 <= p54_literal_2043896;
    p55_literal_2043910 <= p54_literal_2043910;
    p55_literal_2043912 <= p54_literal_2043912;
    p55_literal_2043914 <= p54_literal_2043914;
    p55_literal_2043916 <= p54_literal_2043916;
    p55_literal_2043918 <= p54_literal_2043918;
    p55_literal_2043920 <= p54_literal_2043920;
    p55_literal_2043923 <= p54_literal_2043923;
  end

  // ===== Pipe stage 55:
  wire [7:0] p55_array_index_2053952_comb;
  wire [7:0] p55_array_index_2053953_comb;
  wire [7:0] p55_array_index_2053954_comb;
  wire [7:0] p55_array_index_2053955_comb;
  wire [7:0] p55_array_index_2053956_comb;
  wire [7:0] p55_res7__710_comb;
  wire [7:0] p55_array_index_2053967_comb;
  wire [7:0] p55_array_index_2053968_comb;
  wire [7:0] p55_array_index_2053969_comb;
  wire [7:0] p55_array_index_2053970_comb;
  wire [7:0] p55_res7__712_comb;
  wire [7:0] p55_array_index_2053980_comb;
  wire [7:0] p55_array_index_2053981_comb;
  wire [7:0] p55_array_index_2053982_comb;
  wire [7:0] p55_array_index_2053983_comb;
  wire [7:0] p55_res7__714_comb;
  wire [7:0] p55_array_index_2053994_comb;
  wire [7:0] p55_array_index_2053995_comb;
  wire [7:0] p55_array_index_2053996_comb;
  wire [7:0] p55_res7__716_comb;
  wire [7:0] p55_array_index_2054006_comb;
  wire [7:0] p55_array_index_2054007_comb;
  wire [7:0] p55_array_index_2054008_comb;
  wire [7:0] p55_res7__718_comb;
  wire [7:0] p55_array_index_2054019_comb;
  wire [7:0] p55_array_index_2054020_comb;
  wire [7:0] p55_res7__720_comb;
  wire [7:0] p55_array_index_2054030_comb;
  wire [7:0] p55_array_index_2054031_comb;
  wire [7:0] p55_res7__722_comb;
  assign p55_array_index_2053952_comb = p54_literal_2043912[p54_res7__706];
  assign p55_array_index_2053953_comb = p54_literal_2043914[p54_res7__704];
  assign p55_array_index_2053954_comb = p54_literal_2043916[p54_array_index_2053790];
  assign p55_array_index_2053955_comb = p54_literal_2043918[p54_array_index_2053791];
  assign p55_array_index_2053956_comb = p54_literal_2043920[p54_array_index_2053792];
  assign p55_res7__710_comb = p54_literal_2043910[p54_res7__708] ^ p55_array_index_2053952_comb ^ p55_array_index_2053953_comb ^ p55_array_index_2053954_comb ^ p55_array_index_2053955_comb ^ p55_array_index_2053956_comb ^ p54_array_index_2053793 ^ p54_literal_2043923[p54_array_index_2053794] ^ p54_array_index_2053795 ^ p54_literal_2043920[p54_array_index_2053812] ^ p54_literal_2043918[p54_array_index_2053797] ^ p54_literal_2043916[p54_array_index_2053814] ^ p54_literal_2043914[p54_array_index_2053799] ^ p54_literal_2043912[p54_array_index_2053800] ^ p54_literal_2043910[p54_array_index_2053801] ^ p54_array_index_2053802;
  assign p55_array_index_2053967_comb = p54_literal_2043914[p54_res7__706];
  assign p55_array_index_2053968_comb = p54_literal_2043916[p54_res7__704];
  assign p55_array_index_2053969_comb = p54_literal_2043918[p54_array_index_2053790];
  assign p55_array_index_2053970_comb = p54_literal_2043920[p54_array_index_2053791];
  assign p55_res7__712_comb = p54_literal_2043910[p55_res7__710_comb] ^ p54_literal_2043912[p54_res7__708] ^ p55_array_index_2053967_comb ^ p55_array_index_2053968_comb ^ p55_array_index_2053969_comb ^ p55_array_index_2053970_comb ^ p54_array_index_2053792 ^ p54_literal_2043923[p54_array_index_2053793] ^ p54_array_index_2053794 ^ p54_array_index_2053811 ^ p54_literal_2043918[p54_array_index_2053812] ^ p54_literal_2043916[p54_array_index_2053797] ^ p54_literal_2043914[p54_array_index_2053814] ^ p54_literal_2043912[p54_array_index_2053799] ^ p54_literal_2043910[p54_array_index_2053800] ^ p54_array_index_2053801;
  assign p55_array_index_2053980_comb = p54_literal_2043914[p54_res7__708];
  assign p55_array_index_2053981_comb = p54_literal_2043916[p54_res7__706];
  assign p55_array_index_2053982_comb = p54_literal_2043918[p54_res7__704];
  assign p55_array_index_2053983_comb = p54_literal_2043920[p54_array_index_2053790];
  assign p55_res7__714_comb = p54_literal_2043910[p55_res7__712_comb] ^ p54_literal_2043912[p55_res7__710_comb] ^ p55_array_index_2053980_comb ^ p55_array_index_2053981_comb ^ p55_array_index_2053982_comb ^ p55_array_index_2053983_comb ^ p54_array_index_2053791 ^ p54_literal_2043923[p54_array_index_2053792] ^ p54_array_index_2053793 ^ p54_array_index_2053828 ^ p54_literal_2043918[p54_array_index_2053795] ^ p54_literal_2043916[p54_array_index_2053812] ^ p54_literal_2043914[p54_array_index_2053797] ^ p54_literal_2043912[p54_array_index_2053814] ^ p54_literal_2043910[p54_array_index_2053799] ^ p54_array_index_2053800;
  assign p55_array_index_2053994_comb = p54_literal_2043916[p54_res7__708];
  assign p55_array_index_2053995_comb = p54_literal_2043918[p54_res7__706];
  assign p55_array_index_2053996_comb = p54_literal_2043920[p54_res7__704];
  assign p55_res7__716_comb = p54_literal_2043910[p55_res7__714_comb] ^ p54_literal_2043912[p55_res7__712_comb] ^ p54_literal_2043914[p55_res7__710_comb] ^ p55_array_index_2053994_comb ^ p55_array_index_2053995_comb ^ p55_array_index_2053996_comb ^ p54_array_index_2053790 ^ p54_literal_2043923[p54_array_index_2053791] ^ p54_array_index_2053792 ^ p54_array_index_2053842 ^ p54_array_index_2053810 ^ p54_literal_2043916[p54_array_index_2053795] ^ p54_literal_2043914[p54_array_index_2053812] ^ p54_literal_2043912[p54_array_index_2053797] ^ p54_literal_2043910[p54_array_index_2053814] ^ p54_array_index_2053799;
  assign p55_array_index_2054006_comb = p54_literal_2043916[p55_res7__710_comb];
  assign p55_array_index_2054007_comb = p54_literal_2043918[p54_res7__708];
  assign p55_array_index_2054008_comb = p54_literal_2043920[p54_res7__706];
  assign p55_res7__718_comb = p54_literal_2043910[p55_res7__716_comb] ^ p54_literal_2043912[p55_res7__714_comb] ^ p54_literal_2043914[p55_res7__712_comb] ^ p55_array_index_2054006_comb ^ p55_array_index_2054007_comb ^ p55_array_index_2054008_comb ^ p54_res7__704 ^ p54_literal_2043923[p54_array_index_2053790] ^ p54_array_index_2053791 ^ p55_array_index_2053956_comb ^ p54_array_index_2053827 ^ p54_literal_2043916[p54_array_index_2053794] ^ p54_literal_2043914[p54_array_index_2053795] ^ p54_literal_2043912[p54_array_index_2053812] ^ p54_literal_2043910[p54_array_index_2053797] ^ p54_array_index_2053814;
  assign p55_array_index_2054019_comb = p54_literal_2043918[p55_res7__710_comb];
  assign p55_array_index_2054020_comb = p54_literal_2043920[p54_res7__708];
  assign p55_res7__720_comb = p54_literal_2043910[p55_res7__718_comb] ^ p54_literal_2043912[p55_res7__716_comb] ^ p54_literal_2043914[p55_res7__714_comb] ^ p54_literal_2043916[p55_res7__712_comb] ^ p55_array_index_2054019_comb ^ p55_array_index_2054020_comb ^ p54_res7__706 ^ p54_literal_2043923[p54_res7__704] ^ p54_array_index_2053790 ^ p55_array_index_2053970_comb ^ p54_array_index_2053841 ^ p54_array_index_2053809 ^ p54_literal_2043914[p54_array_index_2053794] ^ p54_literal_2043912[p54_array_index_2053795] ^ p54_literal_2043910[p54_array_index_2053812] ^ p54_array_index_2053797;
  assign p55_array_index_2054030_comb = p54_literal_2043918[p55_res7__712_comb];
  assign p55_array_index_2054031_comb = p54_literal_2043920[p55_res7__710_comb];
  assign p55_res7__722_comb = p54_literal_2043910[p55_res7__720_comb] ^ p54_literal_2043912[p55_res7__718_comb] ^ p54_literal_2043914[p55_res7__716_comb] ^ p54_literal_2043916[p55_res7__714_comb] ^ p55_array_index_2054030_comb ^ p55_array_index_2054031_comb ^ p54_res7__708 ^ p54_literal_2043923[p54_res7__706] ^ p54_res7__704 ^ p55_array_index_2053983_comb ^ p55_array_index_2053955_comb ^ p54_array_index_2053826 ^ p54_literal_2043914[p54_array_index_2053793] ^ p54_literal_2043912[p54_array_index_2053794] ^ p54_literal_2043910[p54_array_index_2053795] ^ p54_array_index_2053812;

  // Registers for pipe stage 55:
  reg [127:0] p55_encoded;
  reg [127:0] p55_bit_slice_2043893;
  reg [127:0] p55_bit_slice_2044018;
  reg [127:0] p55_k3;
  reg [127:0] p55_k2;
  reg [127:0] p55_k5;
  reg [127:0] p55_k4;
  reg [127:0] p55_xor_2053334;
  reg [127:0] p55_xor_2053774;
  reg [7:0] p55_array_index_2053790;
  reg [7:0] p55_array_index_2053791;
  reg [7:0] p55_array_index_2053792;
  reg [7:0] p55_array_index_2053793;
  reg [7:0] p55_array_index_2053794;
  reg [7:0] p55_array_index_2053795;
  reg [7:0] p55_array_index_2053806;
  reg [7:0] p55_array_index_2053807;
  reg [7:0] p55_array_index_2053808;
  reg [7:0] p55_res7__704;
  reg [7:0] p55_array_index_2053823;
  reg [7:0] p55_array_index_2053824;
  reg [7:0] p55_array_index_2053825;
  reg [7:0] p55_res7__706;
  reg [7:0] p55_array_index_2053838;
  reg [7:0] p55_array_index_2053839;
  reg [7:0] p55_array_index_2053840;
  reg [7:0] p55_res7__708;
  reg [7:0] p55_array_index_2053952;
  reg [7:0] p55_array_index_2053953;
  reg [7:0] p55_array_index_2053954;
  reg [7:0] p55_res7__710;
  reg [7:0] p55_array_index_2053967;
  reg [7:0] p55_array_index_2053968;
  reg [7:0] p55_array_index_2053969;
  reg [7:0] p55_res7__712;
  reg [7:0] p55_array_index_2053980;
  reg [7:0] p55_array_index_2053981;
  reg [7:0] p55_array_index_2053982;
  reg [7:0] p55_res7__714;
  reg [7:0] p55_array_index_2053994;
  reg [7:0] p55_array_index_2053995;
  reg [7:0] p55_array_index_2053996;
  reg [7:0] p55_res7__716;
  reg [7:0] p55_array_index_2054006;
  reg [7:0] p55_array_index_2054007;
  reg [7:0] p55_array_index_2054008;
  reg [7:0] p55_res7__718;
  reg [7:0] p55_array_index_2054019;
  reg [7:0] p55_array_index_2054020;
  reg [7:0] p55_res7__720;
  reg [7:0] p55_array_index_2054030;
  reg [7:0] p55_array_index_2054031;
  reg [7:0] p55_res7__722;
  reg [7:0] p56_literal_2043896[256];
  reg [7:0] p56_literal_2043910[256];
  reg [7:0] p56_literal_2043912[256];
  reg [7:0] p56_literal_2043914[256];
  reg [7:0] p56_literal_2043916[256];
  reg [7:0] p56_literal_2043918[256];
  reg [7:0] p56_literal_2043920[256];
  reg [7:0] p56_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p55_encoded <= p54_encoded;
    p55_bit_slice_2043893 <= p54_bit_slice_2043893;
    p55_bit_slice_2044018 <= p54_bit_slice_2044018;
    p55_k3 <= p54_k3;
    p55_k2 <= p54_k2;
    p55_k5 <= p54_k5;
    p55_k4 <= p54_k4;
    p55_xor_2053334 <= p54_xor_2053334;
    p55_xor_2053774 <= p54_xor_2053774;
    p55_array_index_2053790 <= p54_array_index_2053790;
    p55_array_index_2053791 <= p54_array_index_2053791;
    p55_array_index_2053792 <= p54_array_index_2053792;
    p55_array_index_2053793 <= p54_array_index_2053793;
    p55_array_index_2053794 <= p54_array_index_2053794;
    p55_array_index_2053795 <= p54_array_index_2053795;
    p55_array_index_2053806 <= p54_array_index_2053806;
    p55_array_index_2053807 <= p54_array_index_2053807;
    p55_array_index_2053808 <= p54_array_index_2053808;
    p55_res7__704 <= p54_res7__704;
    p55_array_index_2053823 <= p54_array_index_2053823;
    p55_array_index_2053824 <= p54_array_index_2053824;
    p55_array_index_2053825 <= p54_array_index_2053825;
    p55_res7__706 <= p54_res7__706;
    p55_array_index_2053838 <= p54_array_index_2053838;
    p55_array_index_2053839 <= p54_array_index_2053839;
    p55_array_index_2053840 <= p54_array_index_2053840;
    p55_res7__708 <= p54_res7__708;
    p55_array_index_2053952 <= p55_array_index_2053952_comb;
    p55_array_index_2053953 <= p55_array_index_2053953_comb;
    p55_array_index_2053954 <= p55_array_index_2053954_comb;
    p55_res7__710 <= p55_res7__710_comb;
    p55_array_index_2053967 <= p55_array_index_2053967_comb;
    p55_array_index_2053968 <= p55_array_index_2053968_comb;
    p55_array_index_2053969 <= p55_array_index_2053969_comb;
    p55_res7__712 <= p55_res7__712_comb;
    p55_array_index_2053980 <= p55_array_index_2053980_comb;
    p55_array_index_2053981 <= p55_array_index_2053981_comb;
    p55_array_index_2053982 <= p55_array_index_2053982_comb;
    p55_res7__714 <= p55_res7__714_comb;
    p55_array_index_2053994 <= p55_array_index_2053994_comb;
    p55_array_index_2053995 <= p55_array_index_2053995_comb;
    p55_array_index_2053996 <= p55_array_index_2053996_comb;
    p55_res7__716 <= p55_res7__716_comb;
    p55_array_index_2054006 <= p55_array_index_2054006_comb;
    p55_array_index_2054007 <= p55_array_index_2054007_comb;
    p55_array_index_2054008 <= p55_array_index_2054008_comb;
    p55_res7__718 <= p55_res7__718_comb;
    p55_array_index_2054019 <= p55_array_index_2054019_comb;
    p55_array_index_2054020 <= p55_array_index_2054020_comb;
    p55_res7__720 <= p55_res7__720_comb;
    p55_array_index_2054030 <= p55_array_index_2054030_comb;
    p55_array_index_2054031 <= p55_array_index_2054031_comb;
    p55_res7__722 <= p55_res7__722_comb;
    p56_literal_2043896 <= p55_literal_2043896;
    p56_literal_2043910 <= p55_literal_2043910;
    p56_literal_2043912 <= p55_literal_2043912;
    p56_literal_2043914 <= p55_literal_2043914;
    p56_literal_2043916 <= p55_literal_2043916;
    p56_literal_2043918 <= p55_literal_2043918;
    p56_literal_2043920 <= p55_literal_2043920;
    p56_literal_2043923 <= p55_literal_2043923;
  end

  // ===== Pipe stage 56:
  wire [7:0] p56_array_index_2054164_comb;
  wire [7:0] p56_res7__724_comb;
  wire [7:0] p56_array_index_2054174_comb;
  wire [7:0] p56_res7__726_comb;
  wire [7:0] p56_res7__728_comb;
  wire [7:0] p56_res7__730_comb;
  wire [7:0] p56_res7__732_comb;
  wire [7:0] p56_res7__734_comb;
  wire [127:0] p56_res__22_comb;
  wire [127:0] p56_k7_comb;
  wire [127:0] p56_addedKey__55_comb;
  wire [7:0] p56_array_index_2054230_comb;
  wire [7:0] p56_array_index_2054231_comb;
  wire [7:0] p56_array_index_2054232_comb;
  wire [7:0] p56_array_index_2054233_comb;
  wire [7:0] p56_array_index_2054234_comb;
  wire [7:0] p56_array_index_2054235_comb;
  wire [7:0] p56_array_index_2054237_comb;
  wire [7:0] p56_array_index_2054239_comb;
  wire [7:0] p56_array_index_2054240_comb;
  wire [7:0] p56_array_index_2054241_comb;
  wire [7:0] p56_array_index_2054242_comb;
  wire [7:0] p56_array_index_2054243_comb;
  wire [7:0] p56_array_index_2054244_comb;
  wire [7:0] p56_array_index_2054246_comb;
  wire [7:0] p56_array_index_2054247_comb;
  wire [7:0] p56_array_index_2054248_comb;
  assign p56_array_index_2054164_comb = p55_literal_2043920[p55_res7__712];
  assign p56_res7__724_comb = p55_literal_2043910[p55_res7__722] ^ p55_literal_2043912[p55_res7__720] ^ p55_literal_2043914[p55_res7__718] ^ p55_literal_2043916[p55_res7__716] ^ p55_literal_2043918[p55_res7__714] ^ p56_array_index_2054164_comb ^ p55_res7__710 ^ p55_literal_2043923[p55_res7__708] ^ p55_res7__706 ^ p55_array_index_2053996 ^ p55_array_index_2053969 ^ p55_array_index_2053840 ^ p55_array_index_2053808 ^ p55_literal_2043912[p55_array_index_2053793] ^ p55_literal_2043910[p55_array_index_2053794] ^ p55_array_index_2053795;
  assign p56_array_index_2054174_comb = p55_literal_2043920[p55_res7__714];
  assign p56_res7__726_comb = p55_literal_2043910[p56_res7__724_comb] ^ p55_literal_2043912[p55_res7__722] ^ p55_literal_2043914[p55_res7__720] ^ p55_literal_2043916[p55_res7__718] ^ p55_literal_2043918[p55_res7__716] ^ p56_array_index_2054174_comb ^ p55_res7__712 ^ p55_literal_2043923[p55_res7__710] ^ p55_res7__708 ^ p55_array_index_2054008 ^ p55_array_index_2053982 ^ p55_array_index_2053954 ^ p55_array_index_2053825 ^ p55_literal_2043912[p55_array_index_2053792] ^ p55_literal_2043910[p55_array_index_2053793] ^ p55_array_index_2053794;
  assign p56_res7__728_comb = p55_literal_2043910[p56_res7__726_comb] ^ p55_literal_2043912[p56_res7__724_comb] ^ p55_literal_2043914[p55_res7__722] ^ p55_literal_2043916[p55_res7__720] ^ p55_literal_2043918[p55_res7__718] ^ p55_literal_2043920[p55_res7__716] ^ p55_res7__714 ^ p55_literal_2043923[p55_res7__712] ^ p55_res7__710 ^ p55_array_index_2054020 ^ p55_array_index_2053995 ^ p55_array_index_2053968 ^ p55_array_index_2053839 ^ p55_array_index_2053807 ^ p55_literal_2043910[p55_array_index_2053792] ^ p55_array_index_2053793;
  assign p56_res7__730_comb = p55_literal_2043910[p56_res7__728_comb] ^ p55_literal_2043912[p56_res7__726_comb] ^ p55_literal_2043914[p56_res7__724_comb] ^ p55_literal_2043916[p55_res7__722] ^ p55_literal_2043918[p55_res7__720] ^ p55_literal_2043920[p55_res7__718] ^ p55_res7__716 ^ p55_literal_2043923[p55_res7__714] ^ p55_res7__712 ^ p55_array_index_2054031 ^ p55_array_index_2054007 ^ p55_array_index_2053981 ^ p55_array_index_2053953 ^ p55_array_index_2053824 ^ p55_literal_2043910[p55_array_index_2053791] ^ p55_array_index_2053792;
  assign p56_res7__732_comb = p55_literal_2043910[p56_res7__730_comb] ^ p55_literal_2043912[p56_res7__728_comb] ^ p55_literal_2043914[p56_res7__726_comb] ^ p55_literal_2043916[p56_res7__724_comb] ^ p55_literal_2043918[p55_res7__722] ^ p55_literal_2043920[p55_res7__720] ^ p55_res7__718 ^ p55_literal_2043923[p55_res7__716] ^ p55_res7__714 ^ p56_array_index_2054164_comb ^ p55_array_index_2054019 ^ p55_array_index_2053994 ^ p55_array_index_2053967 ^ p55_array_index_2053838 ^ p55_array_index_2053806 ^ p55_array_index_2053791;
  assign p56_res7__734_comb = p55_literal_2043910[p56_res7__732_comb] ^ p55_literal_2043912[p56_res7__730_comb] ^ p55_literal_2043914[p56_res7__728_comb] ^ p55_literal_2043916[p56_res7__726_comb] ^ p55_literal_2043918[p56_res7__724_comb] ^ p55_literal_2043920[p55_res7__722] ^ p55_res7__720 ^ p55_literal_2043923[p55_res7__718] ^ p55_res7__716 ^ p56_array_index_2054174_comb ^ p55_array_index_2054030 ^ p55_array_index_2054006 ^ p55_array_index_2053980 ^ p55_array_index_2053952 ^ p55_array_index_2053823 ^ p55_array_index_2053790;
  assign p56_res__22_comb = {p56_res7__734_comb, p56_res7__732_comb, p56_res7__730_comb, p56_res7__728_comb, p56_res7__726_comb, p56_res7__724_comb, p55_res7__722, p55_res7__720, p55_res7__718, p55_res7__716, p55_res7__714, p55_res7__712, p55_res7__710, p55_res7__708, p55_res7__706, p55_res7__704};
  assign p56_k7_comb = p56_res__22_comb ^ p55_xor_2053334;
  assign p56_addedKey__55_comb = p56_k7_comb ^ 128'hd9eb_5a3a_e90f_fa58_34ce_2043_693d_7e18;
  assign p56_array_index_2054230_comb = p55_literal_2043896[p56_addedKey__55_comb[127:120]];
  assign p56_array_index_2054231_comb = p55_literal_2043896[p56_addedKey__55_comb[119:112]];
  assign p56_array_index_2054232_comb = p55_literal_2043896[p56_addedKey__55_comb[111:104]];
  assign p56_array_index_2054233_comb = p55_literal_2043896[p56_addedKey__55_comb[103:96]];
  assign p56_array_index_2054234_comb = p55_literal_2043896[p56_addedKey__55_comb[95:88]];
  assign p56_array_index_2054235_comb = p55_literal_2043896[p56_addedKey__55_comb[87:80]];
  assign p56_array_index_2054237_comb = p55_literal_2043896[p56_addedKey__55_comb[71:64]];
  assign p56_array_index_2054239_comb = p55_literal_2043896[p56_addedKey__55_comb[55:48]];
  assign p56_array_index_2054240_comb = p55_literal_2043896[p56_addedKey__55_comb[47:40]];
  assign p56_array_index_2054241_comb = p55_literal_2043896[p56_addedKey__55_comb[39:32]];
  assign p56_array_index_2054242_comb = p55_literal_2043896[p56_addedKey__55_comb[31:24]];
  assign p56_array_index_2054243_comb = p55_literal_2043896[p56_addedKey__55_comb[23:16]];
  assign p56_array_index_2054244_comb = p55_literal_2043896[p56_addedKey__55_comb[15:8]];
  assign p56_array_index_2054246_comb = p55_literal_2043896[p56_addedKey__55_comb[79:72]];
  assign p56_array_index_2054247_comb = p55_literal_2043896[p56_addedKey__55_comb[63:56]];
  assign p56_array_index_2054248_comb = p55_literal_2043896[p56_addedKey__55_comb[7:0]];

  // Registers for pipe stage 56:
  reg [127:0] p56_encoded;
  reg [127:0] p56_bit_slice_2043893;
  reg [127:0] p56_bit_slice_2044018;
  reg [127:0] p56_k3;
  reg [127:0] p56_k2;
  reg [127:0] p56_k5;
  reg [127:0] p56_k4;
  reg [127:0] p56_xor_2053774;
  reg [127:0] p56_k7;
  reg [7:0] p56_array_index_2054230;
  reg [7:0] p56_array_index_2054231;
  reg [7:0] p56_array_index_2054232;
  reg [7:0] p56_array_index_2054233;
  reg [7:0] p56_array_index_2054234;
  reg [7:0] p56_array_index_2054235;
  reg [7:0] p56_array_index_2054237;
  reg [7:0] p56_array_index_2054239;
  reg [7:0] p56_array_index_2054240;
  reg [7:0] p56_array_index_2054241;
  reg [7:0] p56_array_index_2054242;
  reg [7:0] p56_array_index_2054243;
  reg [7:0] p56_array_index_2054244;
  reg [7:0] p56_array_index_2054246;
  reg [7:0] p56_array_index_2054247;
  reg [7:0] p56_array_index_2054248;
  reg [7:0] p57_literal_2043896[256];
  reg [7:0] p57_literal_2043910[256];
  reg [7:0] p57_literal_2043912[256];
  reg [7:0] p57_literal_2043914[256];
  reg [7:0] p57_literal_2043916[256];
  reg [7:0] p57_literal_2043918[256];
  reg [7:0] p57_literal_2043920[256];
  reg [7:0] p57_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p56_encoded <= p55_encoded;
    p56_bit_slice_2043893 <= p55_bit_slice_2043893;
    p56_bit_slice_2044018 <= p55_bit_slice_2044018;
    p56_k3 <= p55_k3;
    p56_k2 <= p55_k2;
    p56_k5 <= p55_k5;
    p56_k4 <= p55_k4;
    p56_xor_2053774 <= p55_xor_2053774;
    p56_k7 <= p56_k7_comb;
    p56_array_index_2054230 <= p56_array_index_2054230_comb;
    p56_array_index_2054231 <= p56_array_index_2054231_comb;
    p56_array_index_2054232 <= p56_array_index_2054232_comb;
    p56_array_index_2054233 <= p56_array_index_2054233_comb;
    p56_array_index_2054234 <= p56_array_index_2054234_comb;
    p56_array_index_2054235 <= p56_array_index_2054235_comb;
    p56_array_index_2054237 <= p56_array_index_2054237_comb;
    p56_array_index_2054239 <= p56_array_index_2054239_comb;
    p56_array_index_2054240 <= p56_array_index_2054240_comb;
    p56_array_index_2054241 <= p56_array_index_2054241_comb;
    p56_array_index_2054242 <= p56_array_index_2054242_comb;
    p56_array_index_2054243 <= p56_array_index_2054243_comb;
    p56_array_index_2054244 <= p56_array_index_2054244_comb;
    p56_array_index_2054246 <= p56_array_index_2054246_comb;
    p56_array_index_2054247 <= p56_array_index_2054247_comb;
    p56_array_index_2054248 <= p56_array_index_2054248_comb;
    p57_literal_2043896 <= p56_literal_2043896;
    p57_literal_2043910 <= p56_literal_2043910;
    p57_literal_2043912 <= p56_literal_2043912;
    p57_literal_2043914 <= p56_literal_2043914;
    p57_literal_2043916 <= p56_literal_2043916;
    p57_literal_2043918 <= p56_literal_2043918;
    p57_literal_2043920 <= p56_literal_2043920;
    p57_literal_2043923 <= p56_literal_2043923;
  end

  // ===== Pipe stage 57:
  wire [7:0] p57_array_index_2054315_comb;
  wire [7:0] p57_array_index_2054316_comb;
  wire [7:0] p57_array_index_2054317_comb;
  wire [7:0] p57_array_index_2054318_comb;
  wire [7:0] p57_array_index_2054319_comb;
  wire [7:0] p57_array_index_2054320_comb;
  wire [7:0] p57_res7__736_comb;
  wire [7:0] p57_array_index_2054329_comb;
  wire [7:0] p57_array_index_2054330_comb;
  wire [7:0] p57_array_index_2054331_comb;
  wire [7:0] p57_array_index_2054332_comb;
  wire [7:0] p57_array_index_2054333_comb;
  wire [7:0] p57_array_index_2054334_comb;
  wire [7:0] p57_res7__738_comb;
  wire [7:0] p57_array_index_2054344_comb;
  wire [7:0] p57_array_index_2054345_comb;
  wire [7:0] p57_array_index_2054346_comb;
  wire [7:0] p57_array_index_2054347_comb;
  wire [7:0] p57_array_index_2054348_comb;
  wire [7:0] p57_res7__740_comb;
  wire [7:0] p57_array_index_2054358_comb;
  wire [7:0] p57_array_index_2054359_comb;
  wire [7:0] p57_array_index_2054360_comb;
  wire [7:0] p57_array_index_2054361_comb;
  wire [7:0] p57_array_index_2054362_comb;
  wire [7:0] p57_res7__742_comb;
  wire [7:0] p57_array_index_2054373_comb;
  wire [7:0] p57_array_index_2054374_comb;
  wire [7:0] p57_array_index_2054375_comb;
  wire [7:0] p57_array_index_2054376_comb;
  wire [7:0] p57_res7__744_comb;
  wire [7:0] p57_array_index_2054386_comb;
  wire [7:0] p57_array_index_2054387_comb;
  wire [7:0] p57_array_index_2054388_comb;
  wire [7:0] p57_array_index_2054389_comb;
  wire [7:0] p57_res7__746_comb;
  wire [7:0] p57_array_index_2054400_comb;
  wire [7:0] p57_array_index_2054401_comb;
  wire [7:0] p57_array_index_2054402_comb;
  wire [7:0] p57_res7__748_comb;
  assign p57_array_index_2054315_comb = p56_literal_2043910[p56_array_index_2054230];
  assign p57_array_index_2054316_comb = p56_literal_2043912[p56_array_index_2054231];
  assign p57_array_index_2054317_comb = p56_literal_2043914[p56_array_index_2054232];
  assign p57_array_index_2054318_comb = p56_literal_2043916[p56_array_index_2054233];
  assign p57_array_index_2054319_comb = p56_literal_2043918[p56_array_index_2054234];
  assign p57_array_index_2054320_comb = p56_literal_2043920[p56_array_index_2054235];
  assign p57_res7__736_comb = p57_array_index_2054315_comb ^ p57_array_index_2054316_comb ^ p57_array_index_2054317_comb ^ p57_array_index_2054318_comb ^ p57_array_index_2054319_comb ^ p57_array_index_2054320_comb ^ p56_array_index_2054246 ^ p56_literal_2043923[p56_array_index_2054237] ^ p56_array_index_2054247 ^ p56_literal_2043920[p56_array_index_2054239] ^ p56_literal_2043918[p56_array_index_2054240] ^ p56_literal_2043916[p56_array_index_2054241] ^ p56_literal_2043914[p56_array_index_2054242] ^ p56_literal_2043912[p56_array_index_2054243] ^ p56_literal_2043910[p56_array_index_2054244] ^ p56_array_index_2054248;
  assign p57_array_index_2054329_comb = p56_literal_2043910[p57_res7__736_comb];
  assign p57_array_index_2054330_comb = p56_literal_2043912[p56_array_index_2054230];
  assign p57_array_index_2054331_comb = p56_literal_2043914[p56_array_index_2054231];
  assign p57_array_index_2054332_comb = p56_literal_2043916[p56_array_index_2054232];
  assign p57_array_index_2054333_comb = p56_literal_2043918[p56_array_index_2054233];
  assign p57_array_index_2054334_comb = p56_literal_2043920[p56_array_index_2054234];
  assign p57_res7__738_comb = p57_array_index_2054329_comb ^ p57_array_index_2054330_comb ^ p57_array_index_2054331_comb ^ p57_array_index_2054332_comb ^ p57_array_index_2054333_comb ^ p57_array_index_2054334_comb ^ p56_array_index_2054235 ^ p56_literal_2043923[p56_array_index_2054246] ^ p56_array_index_2054237 ^ p56_literal_2043920[p56_array_index_2054247] ^ p56_literal_2043918[p56_array_index_2054239] ^ p56_literal_2043916[p56_array_index_2054240] ^ p56_literal_2043914[p56_array_index_2054241] ^ p56_literal_2043912[p56_array_index_2054242] ^ p56_literal_2043910[p56_array_index_2054243] ^ p56_array_index_2054244;
  assign p57_array_index_2054344_comb = p56_literal_2043912[p57_res7__736_comb];
  assign p57_array_index_2054345_comb = p56_literal_2043914[p56_array_index_2054230];
  assign p57_array_index_2054346_comb = p56_literal_2043916[p56_array_index_2054231];
  assign p57_array_index_2054347_comb = p56_literal_2043918[p56_array_index_2054232];
  assign p57_array_index_2054348_comb = p56_literal_2043920[p56_array_index_2054233];
  assign p57_res7__740_comb = p56_literal_2043910[p57_res7__738_comb] ^ p57_array_index_2054344_comb ^ p57_array_index_2054345_comb ^ p57_array_index_2054346_comb ^ p57_array_index_2054347_comb ^ p57_array_index_2054348_comb ^ p56_array_index_2054234 ^ p56_literal_2043923[p56_array_index_2054235] ^ p56_array_index_2054246 ^ p56_literal_2043920[p56_array_index_2054237] ^ p56_literal_2043918[p56_array_index_2054247] ^ p56_literal_2043916[p56_array_index_2054239] ^ p56_literal_2043914[p56_array_index_2054240] ^ p56_literal_2043912[p56_array_index_2054241] ^ p56_literal_2043910[p56_array_index_2054242] ^ p56_array_index_2054243;
  assign p57_array_index_2054358_comb = p56_literal_2043912[p57_res7__738_comb];
  assign p57_array_index_2054359_comb = p56_literal_2043914[p57_res7__736_comb];
  assign p57_array_index_2054360_comb = p56_literal_2043916[p56_array_index_2054230];
  assign p57_array_index_2054361_comb = p56_literal_2043918[p56_array_index_2054231];
  assign p57_array_index_2054362_comb = p56_literal_2043920[p56_array_index_2054232];
  assign p57_res7__742_comb = p56_literal_2043910[p57_res7__740_comb] ^ p57_array_index_2054358_comb ^ p57_array_index_2054359_comb ^ p57_array_index_2054360_comb ^ p57_array_index_2054361_comb ^ p57_array_index_2054362_comb ^ p56_array_index_2054233 ^ p56_literal_2043923[p56_array_index_2054234] ^ p56_array_index_2054235 ^ p56_literal_2043920[p56_array_index_2054246] ^ p56_literal_2043918[p56_array_index_2054237] ^ p56_literal_2043916[p56_array_index_2054247] ^ p56_literal_2043914[p56_array_index_2054239] ^ p56_literal_2043912[p56_array_index_2054240] ^ p56_literal_2043910[p56_array_index_2054241] ^ p56_array_index_2054242;
  assign p57_array_index_2054373_comb = p56_literal_2043914[p57_res7__738_comb];
  assign p57_array_index_2054374_comb = p56_literal_2043916[p57_res7__736_comb];
  assign p57_array_index_2054375_comb = p56_literal_2043918[p56_array_index_2054230];
  assign p57_array_index_2054376_comb = p56_literal_2043920[p56_array_index_2054231];
  assign p57_res7__744_comb = p56_literal_2043910[p57_res7__742_comb] ^ p56_literal_2043912[p57_res7__740_comb] ^ p57_array_index_2054373_comb ^ p57_array_index_2054374_comb ^ p57_array_index_2054375_comb ^ p57_array_index_2054376_comb ^ p56_array_index_2054232 ^ p56_literal_2043923[p56_array_index_2054233] ^ p56_array_index_2054234 ^ p57_array_index_2054320_comb ^ p56_literal_2043918[p56_array_index_2054246] ^ p56_literal_2043916[p56_array_index_2054237] ^ p56_literal_2043914[p56_array_index_2054247] ^ p56_literal_2043912[p56_array_index_2054239] ^ p56_literal_2043910[p56_array_index_2054240] ^ p56_array_index_2054241;
  assign p57_array_index_2054386_comb = p56_literal_2043914[p57_res7__740_comb];
  assign p57_array_index_2054387_comb = p56_literal_2043916[p57_res7__738_comb];
  assign p57_array_index_2054388_comb = p56_literal_2043918[p57_res7__736_comb];
  assign p57_array_index_2054389_comb = p56_literal_2043920[p56_array_index_2054230];
  assign p57_res7__746_comb = p56_literal_2043910[p57_res7__744_comb] ^ p56_literal_2043912[p57_res7__742_comb] ^ p57_array_index_2054386_comb ^ p57_array_index_2054387_comb ^ p57_array_index_2054388_comb ^ p57_array_index_2054389_comb ^ p56_array_index_2054231 ^ p56_literal_2043923[p56_array_index_2054232] ^ p56_array_index_2054233 ^ p57_array_index_2054334_comb ^ p56_literal_2043918[p56_array_index_2054235] ^ p56_literal_2043916[p56_array_index_2054246] ^ p56_literal_2043914[p56_array_index_2054237] ^ p56_literal_2043912[p56_array_index_2054247] ^ p56_literal_2043910[p56_array_index_2054239] ^ p56_array_index_2054240;
  assign p57_array_index_2054400_comb = p56_literal_2043916[p57_res7__740_comb];
  assign p57_array_index_2054401_comb = p56_literal_2043918[p57_res7__738_comb];
  assign p57_array_index_2054402_comb = p56_literal_2043920[p57_res7__736_comb];
  assign p57_res7__748_comb = p56_literal_2043910[p57_res7__746_comb] ^ p56_literal_2043912[p57_res7__744_comb] ^ p56_literal_2043914[p57_res7__742_comb] ^ p57_array_index_2054400_comb ^ p57_array_index_2054401_comb ^ p57_array_index_2054402_comb ^ p56_array_index_2054230 ^ p56_literal_2043923[p56_array_index_2054231] ^ p56_array_index_2054232 ^ p57_array_index_2054348_comb ^ p57_array_index_2054319_comb ^ p56_literal_2043916[p56_array_index_2054235] ^ p56_literal_2043914[p56_array_index_2054246] ^ p56_literal_2043912[p56_array_index_2054237] ^ p56_literal_2043910[p56_array_index_2054247] ^ p56_array_index_2054239;

  // Registers for pipe stage 57:
  reg [127:0] p57_encoded;
  reg [127:0] p57_bit_slice_2043893;
  reg [127:0] p57_bit_slice_2044018;
  reg [127:0] p57_k3;
  reg [127:0] p57_k2;
  reg [127:0] p57_k5;
  reg [127:0] p57_k4;
  reg [127:0] p57_xor_2053774;
  reg [127:0] p57_k7;
  reg [7:0] p57_array_index_2054230;
  reg [7:0] p57_array_index_2054231;
  reg [7:0] p57_array_index_2054232;
  reg [7:0] p57_array_index_2054233;
  reg [7:0] p57_array_index_2054234;
  reg [7:0] p57_array_index_2054235;
  reg [7:0] p57_array_index_2054237;
  reg [7:0] p57_array_index_2054315;
  reg [7:0] p57_array_index_2054316;
  reg [7:0] p57_array_index_2054317;
  reg [7:0] p57_array_index_2054318;
  reg [7:0] p57_array_index_2054246;
  reg [7:0] p57_array_index_2054247;
  reg [7:0] p57_res7__736;
  reg [7:0] p57_array_index_2054329;
  reg [7:0] p57_array_index_2054330;
  reg [7:0] p57_array_index_2054331;
  reg [7:0] p57_array_index_2054332;
  reg [7:0] p57_array_index_2054333;
  reg [7:0] p57_res7__738;
  reg [7:0] p57_array_index_2054344;
  reg [7:0] p57_array_index_2054345;
  reg [7:0] p57_array_index_2054346;
  reg [7:0] p57_array_index_2054347;
  reg [7:0] p57_res7__740;
  reg [7:0] p57_array_index_2054358;
  reg [7:0] p57_array_index_2054359;
  reg [7:0] p57_array_index_2054360;
  reg [7:0] p57_array_index_2054361;
  reg [7:0] p57_array_index_2054362;
  reg [7:0] p57_res7__742;
  reg [7:0] p57_array_index_2054373;
  reg [7:0] p57_array_index_2054374;
  reg [7:0] p57_array_index_2054375;
  reg [7:0] p57_array_index_2054376;
  reg [7:0] p57_res7__744;
  reg [7:0] p57_array_index_2054386;
  reg [7:0] p57_array_index_2054387;
  reg [7:0] p57_array_index_2054388;
  reg [7:0] p57_array_index_2054389;
  reg [7:0] p57_res7__746;
  reg [7:0] p57_array_index_2054400;
  reg [7:0] p57_array_index_2054401;
  reg [7:0] p57_array_index_2054402;
  reg [7:0] p57_res7__748;
  reg [7:0] p58_literal_2043896[256];
  reg [7:0] p58_literal_2043910[256];
  reg [7:0] p58_literal_2043912[256];
  reg [7:0] p58_literal_2043914[256];
  reg [7:0] p58_literal_2043916[256];
  reg [7:0] p58_literal_2043918[256];
  reg [7:0] p58_literal_2043920[256];
  reg [7:0] p58_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p57_encoded <= p56_encoded;
    p57_bit_slice_2043893 <= p56_bit_slice_2043893;
    p57_bit_slice_2044018 <= p56_bit_slice_2044018;
    p57_k3 <= p56_k3;
    p57_k2 <= p56_k2;
    p57_k5 <= p56_k5;
    p57_k4 <= p56_k4;
    p57_xor_2053774 <= p56_xor_2053774;
    p57_k7 <= p56_k7;
    p57_array_index_2054230 <= p56_array_index_2054230;
    p57_array_index_2054231 <= p56_array_index_2054231;
    p57_array_index_2054232 <= p56_array_index_2054232;
    p57_array_index_2054233 <= p56_array_index_2054233;
    p57_array_index_2054234 <= p56_array_index_2054234;
    p57_array_index_2054235 <= p56_array_index_2054235;
    p57_array_index_2054237 <= p56_array_index_2054237;
    p57_array_index_2054315 <= p57_array_index_2054315_comb;
    p57_array_index_2054316 <= p57_array_index_2054316_comb;
    p57_array_index_2054317 <= p57_array_index_2054317_comb;
    p57_array_index_2054318 <= p57_array_index_2054318_comb;
    p57_array_index_2054246 <= p56_array_index_2054246;
    p57_array_index_2054247 <= p56_array_index_2054247;
    p57_res7__736 <= p57_res7__736_comb;
    p57_array_index_2054329 <= p57_array_index_2054329_comb;
    p57_array_index_2054330 <= p57_array_index_2054330_comb;
    p57_array_index_2054331 <= p57_array_index_2054331_comb;
    p57_array_index_2054332 <= p57_array_index_2054332_comb;
    p57_array_index_2054333 <= p57_array_index_2054333_comb;
    p57_res7__738 <= p57_res7__738_comb;
    p57_array_index_2054344 <= p57_array_index_2054344_comb;
    p57_array_index_2054345 <= p57_array_index_2054345_comb;
    p57_array_index_2054346 <= p57_array_index_2054346_comb;
    p57_array_index_2054347 <= p57_array_index_2054347_comb;
    p57_res7__740 <= p57_res7__740_comb;
    p57_array_index_2054358 <= p57_array_index_2054358_comb;
    p57_array_index_2054359 <= p57_array_index_2054359_comb;
    p57_array_index_2054360 <= p57_array_index_2054360_comb;
    p57_array_index_2054361 <= p57_array_index_2054361_comb;
    p57_array_index_2054362 <= p57_array_index_2054362_comb;
    p57_res7__742 <= p57_res7__742_comb;
    p57_array_index_2054373 <= p57_array_index_2054373_comb;
    p57_array_index_2054374 <= p57_array_index_2054374_comb;
    p57_array_index_2054375 <= p57_array_index_2054375_comb;
    p57_array_index_2054376 <= p57_array_index_2054376_comb;
    p57_res7__744 <= p57_res7__744_comb;
    p57_array_index_2054386 <= p57_array_index_2054386_comb;
    p57_array_index_2054387 <= p57_array_index_2054387_comb;
    p57_array_index_2054388 <= p57_array_index_2054388_comb;
    p57_array_index_2054389 <= p57_array_index_2054389_comb;
    p57_res7__746 <= p57_res7__746_comb;
    p57_array_index_2054400 <= p57_array_index_2054400_comb;
    p57_array_index_2054401 <= p57_array_index_2054401_comb;
    p57_array_index_2054402 <= p57_array_index_2054402_comb;
    p57_res7__748 <= p57_res7__748_comb;
    p58_literal_2043896 <= p57_literal_2043896;
    p58_literal_2043910 <= p57_literal_2043910;
    p58_literal_2043912 <= p57_literal_2043912;
    p58_literal_2043914 <= p57_literal_2043914;
    p58_literal_2043916 <= p57_literal_2043916;
    p58_literal_2043918 <= p57_literal_2043918;
    p58_literal_2043920 <= p57_literal_2043920;
    p58_literal_2043923 <= p57_literal_2043923;
  end

  // ===== Pipe stage 58:
  wire [7:0] p58_array_index_2054536_comb;
  wire [7:0] p58_array_index_2054537_comb;
  wire [7:0] p58_array_index_2054538_comb;
  wire [7:0] p58_res7__750_comb;
  wire [7:0] p58_array_index_2054549_comb;
  wire [7:0] p58_array_index_2054550_comb;
  wire [7:0] p58_res7__752_comb;
  wire [7:0] p58_array_index_2054560_comb;
  wire [7:0] p58_array_index_2054561_comb;
  wire [7:0] p58_res7__754_comb;
  wire [7:0] p58_array_index_2054572_comb;
  wire [7:0] p58_res7__756_comb;
  wire [7:0] p58_array_index_2054582_comb;
  wire [7:0] p58_res7__758_comb;
  wire [7:0] p58_res7__760_comb;
  wire [7:0] p58_res7__762_comb;
  assign p58_array_index_2054536_comb = p57_literal_2043916[p57_res7__742];
  assign p58_array_index_2054537_comb = p57_literal_2043918[p57_res7__740];
  assign p58_array_index_2054538_comb = p57_literal_2043920[p57_res7__738];
  assign p58_res7__750_comb = p57_literal_2043910[p57_res7__748] ^ p57_literal_2043912[p57_res7__746] ^ p57_literal_2043914[p57_res7__744] ^ p58_array_index_2054536_comb ^ p58_array_index_2054537_comb ^ p58_array_index_2054538_comb ^ p57_res7__736 ^ p57_literal_2043923[p57_array_index_2054230] ^ p57_array_index_2054231 ^ p57_array_index_2054362 ^ p57_array_index_2054333 ^ p57_literal_2043916[p57_array_index_2054234] ^ p57_literal_2043914[p57_array_index_2054235] ^ p57_literal_2043912[p57_array_index_2054246] ^ p57_literal_2043910[p57_array_index_2054237] ^ p57_array_index_2054247;
  assign p58_array_index_2054549_comb = p57_literal_2043918[p57_res7__742];
  assign p58_array_index_2054550_comb = p57_literal_2043920[p57_res7__740];
  assign p58_res7__752_comb = p57_literal_2043910[p58_res7__750_comb] ^ p57_literal_2043912[p57_res7__748] ^ p57_literal_2043914[p57_res7__746] ^ p57_literal_2043916[p57_res7__744] ^ p58_array_index_2054549_comb ^ p58_array_index_2054550_comb ^ p57_res7__738 ^ p57_literal_2043923[p57_res7__736] ^ p57_array_index_2054230 ^ p57_array_index_2054376 ^ p57_array_index_2054347 ^ p57_array_index_2054318 ^ p57_literal_2043914[p57_array_index_2054234] ^ p57_literal_2043912[p57_array_index_2054235] ^ p57_literal_2043910[p57_array_index_2054246] ^ p57_array_index_2054237;
  assign p58_array_index_2054560_comb = p57_literal_2043918[p57_res7__744];
  assign p58_array_index_2054561_comb = p57_literal_2043920[p57_res7__742];
  assign p58_res7__754_comb = p57_literal_2043910[p58_res7__752_comb] ^ p57_literal_2043912[p58_res7__750_comb] ^ p57_literal_2043914[p57_res7__748] ^ p57_literal_2043916[p57_res7__746] ^ p58_array_index_2054560_comb ^ p58_array_index_2054561_comb ^ p57_res7__740 ^ p57_literal_2043923[p57_res7__738] ^ p57_res7__736 ^ p57_array_index_2054389 ^ p57_array_index_2054361 ^ p57_array_index_2054332 ^ p57_literal_2043914[p57_array_index_2054233] ^ p57_literal_2043912[p57_array_index_2054234] ^ p57_literal_2043910[p57_array_index_2054235] ^ p57_array_index_2054246;
  assign p58_array_index_2054572_comb = p57_literal_2043920[p57_res7__744];
  assign p58_res7__756_comb = p57_literal_2043910[p58_res7__754_comb] ^ p57_literal_2043912[p58_res7__752_comb] ^ p57_literal_2043914[p58_res7__750_comb] ^ p57_literal_2043916[p57_res7__748] ^ p57_literal_2043918[p57_res7__746] ^ p58_array_index_2054572_comb ^ p57_res7__742 ^ p57_literal_2043923[p57_res7__740] ^ p57_res7__738 ^ p57_array_index_2054402 ^ p57_array_index_2054375 ^ p57_array_index_2054346 ^ p57_array_index_2054317 ^ p57_literal_2043912[p57_array_index_2054233] ^ p57_literal_2043910[p57_array_index_2054234] ^ p57_array_index_2054235;
  assign p58_array_index_2054582_comb = p57_literal_2043920[p57_res7__746];
  assign p58_res7__758_comb = p57_literal_2043910[p58_res7__756_comb] ^ p57_literal_2043912[p58_res7__754_comb] ^ p57_literal_2043914[p58_res7__752_comb] ^ p57_literal_2043916[p58_res7__750_comb] ^ p57_literal_2043918[p57_res7__748] ^ p58_array_index_2054582_comb ^ p57_res7__744 ^ p57_literal_2043923[p57_res7__742] ^ p57_res7__740 ^ p58_array_index_2054538_comb ^ p57_array_index_2054388 ^ p57_array_index_2054360 ^ p57_array_index_2054331 ^ p57_literal_2043912[p57_array_index_2054232] ^ p57_literal_2043910[p57_array_index_2054233] ^ p57_array_index_2054234;
  assign p58_res7__760_comb = p57_literal_2043910[p58_res7__758_comb] ^ p57_literal_2043912[p58_res7__756_comb] ^ p57_literal_2043914[p58_res7__754_comb] ^ p57_literal_2043916[p58_res7__752_comb] ^ p57_literal_2043918[p58_res7__750_comb] ^ p57_literal_2043920[p57_res7__748] ^ p57_res7__746 ^ p57_literal_2043923[p57_res7__744] ^ p57_res7__742 ^ p58_array_index_2054550_comb ^ p57_array_index_2054401 ^ p57_array_index_2054374 ^ p57_array_index_2054345 ^ p57_array_index_2054316 ^ p57_literal_2043910[p57_array_index_2054232] ^ p57_array_index_2054233;
  assign p58_res7__762_comb = p57_literal_2043910[p58_res7__760_comb] ^ p57_literal_2043912[p58_res7__758_comb] ^ p57_literal_2043914[p58_res7__756_comb] ^ p57_literal_2043916[p58_res7__754_comb] ^ p57_literal_2043918[p58_res7__752_comb] ^ p57_literal_2043920[p58_res7__750_comb] ^ p57_res7__748 ^ p57_literal_2043923[p57_res7__746] ^ p57_res7__744 ^ p58_array_index_2054561_comb ^ p58_array_index_2054537_comb ^ p57_array_index_2054387 ^ p57_array_index_2054359 ^ p57_array_index_2054330 ^ p57_literal_2043910[p57_array_index_2054231] ^ p57_array_index_2054232;

  // Registers for pipe stage 58:
  reg [127:0] p58_encoded;
  reg [127:0] p58_bit_slice_2043893;
  reg [127:0] p58_bit_slice_2044018;
  reg [127:0] p58_k3;
  reg [127:0] p58_k2;
  reg [127:0] p58_k5;
  reg [127:0] p58_k4;
  reg [127:0] p58_xor_2053774;
  reg [127:0] p58_k7;
  reg [7:0] p58_array_index_2054230;
  reg [7:0] p58_array_index_2054231;
  reg [7:0] p58_array_index_2054315;
  reg [7:0] p58_res7__736;
  reg [7:0] p58_array_index_2054329;
  reg [7:0] p58_res7__738;
  reg [7:0] p58_array_index_2054344;
  reg [7:0] p58_res7__740;
  reg [7:0] p58_array_index_2054358;
  reg [7:0] p58_res7__742;
  reg [7:0] p58_array_index_2054373;
  reg [7:0] p58_res7__744;
  reg [7:0] p58_array_index_2054386;
  reg [7:0] p58_res7__746;
  reg [7:0] p58_array_index_2054400;
  reg [7:0] p58_res7__748;
  reg [7:0] p58_array_index_2054536;
  reg [7:0] p58_res7__750;
  reg [7:0] p58_array_index_2054549;
  reg [7:0] p58_res7__752;
  reg [7:0] p58_array_index_2054560;
  reg [7:0] p58_res7__754;
  reg [7:0] p58_array_index_2054572;
  reg [7:0] p58_res7__756;
  reg [7:0] p58_array_index_2054582;
  reg [7:0] p58_res7__758;
  reg [7:0] p58_res7__760;
  reg [7:0] p58_res7__762;
  reg [7:0] p59_literal_2043896[256];
  reg [7:0] p59_literal_2043910[256];
  reg [7:0] p59_literal_2043912[256];
  reg [7:0] p59_literal_2043914[256];
  reg [7:0] p59_literal_2043916[256];
  reg [7:0] p59_literal_2043918[256];
  reg [7:0] p59_literal_2043920[256];
  reg [7:0] p59_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p58_encoded <= p57_encoded;
    p58_bit_slice_2043893 <= p57_bit_slice_2043893;
    p58_bit_slice_2044018 <= p57_bit_slice_2044018;
    p58_k3 <= p57_k3;
    p58_k2 <= p57_k2;
    p58_k5 <= p57_k5;
    p58_k4 <= p57_k4;
    p58_xor_2053774 <= p57_xor_2053774;
    p58_k7 <= p57_k7;
    p58_array_index_2054230 <= p57_array_index_2054230;
    p58_array_index_2054231 <= p57_array_index_2054231;
    p58_array_index_2054315 <= p57_array_index_2054315;
    p58_res7__736 <= p57_res7__736;
    p58_array_index_2054329 <= p57_array_index_2054329;
    p58_res7__738 <= p57_res7__738;
    p58_array_index_2054344 <= p57_array_index_2054344;
    p58_res7__740 <= p57_res7__740;
    p58_array_index_2054358 <= p57_array_index_2054358;
    p58_res7__742 <= p57_res7__742;
    p58_array_index_2054373 <= p57_array_index_2054373;
    p58_res7__744 <= p57_res7__744;
    p58_array_index_2054386 <= p57_array_index_2054386;
    p58_res7__746 <= p57_res7__746;
    p58_array_index_2054400 <= p57_array_index_2054400;
    p58_res7__748 <= p57_res7__748;
    p58_array_index_2054536 <= p58_array_index_2054536_comb;
    p58_res7__750 <= p58_res7__750_comb;
    p58_array_index_2054549 <= p58_array_index_2054549_comb;
    p58_res7__752 <= p58_res7__752_comb;
    p58_array_index_2054560 <= p58_array_index_2054560_comb;
    p58_res7__754 <= p58_res7__754_comb;
    p58_array_index_2054572 <= p58_array_index_2054572_comb;
    p58_res7__756 <= p58_res7__756_comb;
    p58_array_index_2054582 <= p58_array_index_2054582_comb;
    p58_res7__758 <= p58_res7__758_comb;
    p58_res7__760 <= p58_res7__760_comb;
    p58_res7__762 <= p58_res7__762_comb;
    p59_literal_2043896 <= p58_literal_2043896;
    p59_literal_2043910 <= p58_literal_2043910;
    p59_literal_2043912 <= p58_literal_2043912;
    p59_literal_2043914 <= p58_literal_2043914;
    p59_literal_2043916 <= p58_literal_2043916;
    p59_literal_2043918 <= p58_literal_2043918;
    p59_literal_2043920 <= p58_literal_2043920;
    p59_literal_2043923 <= p58_literal_2043923;
  end

  // ===== Pipe stage 59:
  wire [7:0] p59_res7__764_comb;
  wire [7:0] p59_res7__766_comb;
  wire [127:0] p59_res__23_comb;
  wire [127:0] p59_k6_comb;
  wire [127:0] p59_addedKey__56_comb;
  wire [7:0] p59_array_index_2054728_comb;
  wire [7:0] p59_array_index_2054729_comb;
  wire [7:0] p59_array_index_2054730_comb;
  wire [7:0] p59_array_index_2054731_comb;
  wire [7:0] p59_array_index_2054732_comb;
  wire [7:0] p59_array_index_2054733_comb;
  wire [7:0] p59_array_index_2054735_comb;
  wire [7:0] p59_array_index_2054737_comb;
  wire [7:0] p59_array_index_2054738_comb;
  wire [7:0] p59_array_index_2054739_comb;
  wire [7:0] p59_array_index_2054740_comb;
  wire [7:0] p59_array_index_2054741_comb;
  wire [7:0] p59_array_index_2054742_comb;
  wire [7:0] p59_array_index_2054744_comb;
  wire [7:0] p59_array_index_2054745_comb;
  wire [7:0] p59_array_index_2054746_comb;
  wire [7:0] p59_array_index_2054747_comb;
  wire [7:0] p59_array_index_2054748_comb;
  wire [7:0] p59_array_index_2054749_comb;
  wire [7:0] p59_array_index_2054750_comb;
  wire [7:0] p59_array_index_2054752_comb;
  wire [7:0] p59_res7__768_comb;
  wire [7:0] p59_array_index_2054761_comb;
  wire [7:0] p59_array_index_2054762_comb;
  wire [7:0] p59_array_index_2054763_comb;
  wire [7:0] p59_array_index_2054764_comb;
  wire [7:0] p59_array_index_2054765_comb;
  wire [7:0] p59_array_index_2054766_comb;
  wire [7:0] p59_res7__770_comb;
  wire [7:0] p59_array_index_2054776_comb;
  wire [7:0] p59_array_index_2054777_comb;
  wire [7:0] p59_array_index_2054778_comb;
  wire [7:0] p59_array_index_2054779_comb;
  wire [7:0] p59_array_index_2054780_comb;
  wire [7:0] p59_res7__772_comb;
  wire [7:0] p59_array_index_2054790_comb;
  wire [7:0] p59_array_index_2054791_comb;
  wire [7:0] p59_array_index_2054792_comb;
  wire [7:0] p59_array_index_2054793_comb;
  wire [7:0] p59_array_index_2054794_comb;
  wire [7:0] p59_res7__774_comb;
  assign p59_res7__764_comb = p58_literal_2043910[p58_res7__762] ^ p58_literal_2043912[p58_res7__760] ^ p58_literal_2043914[p58_res7__758] ^ p58_literal_2043916[p58_res7__756] ^ p58_literal_2043918[p58_res7__754] ^ p58_literal_2043920[p58_res7__752] ^ p58_res7__750 ^ p58_literal_2043923[p58_res7__748] ^ p58_res7__746 ^ p58_array_index_2054572 ^ p58_array_index_2054549 ^ p58_array_index_2054400 ^ p58_array_index_2054373 ^ p58_array_index_2054344 ^ p58_array_index_2054315 ^ p58_array_index_2054231;
  assign p59_res7__766_comb = p58_literal_2043910[p59_res7__764_comb] ^ p58_literal_2043912[p58_res7__762] ^ p58_literal_2043914[p58_res7__760] ^ p58_literal_2043916[p58_res7__758] ^ p58_literal_2043918[p58_res7__756] ^ p58_literal_2043920[p58_res7__754] ^ p58_res7__752 ^ p58_literal_2043923[p58_res7__750] ^ p58_res7__748 ^ p58_array_index_2054582 ^ p58_array_index_2054560 ^ p58_array_index_2054536 ^ p58_array_index_2054386 ^ p58_array_index_2054358 ^ p58_array_index_2054329 ^ p58_array_index_2054230;
  assign p59_res__23_comb = {p59_res7__766_comb, p59_res7__764_comb, p58_res7__762, p58_res7__760, p58_res7__758, p58_res7__756, p58_res7__754, p58_res7__752, p58_res7__750, p58_res7__748, p58_res7__746, p58_res7__744, p58_res7__742, p58_res7__740, p58_res7__738, p58_res7__736};
  assign p59_k6_comb = p59_res__23_comb ^ p58_xor_2053774;
  assign p59_addedKey__56_comb = p59_k6_comb ^ 128'hb749_2c48_8547_80e0_69e9_9d53_b4b9_ea19;
  assign p59_array_index_2054728_comb = p58_literal_2043896[p59_addedKey__56_comb[127:120]];
  assign p59_array_index_2054729_comb = p58_literal_2043896[p59_addedKey__56_comb[119:112]];
  assign p59_array_index_2054730_comb = p58_literal_2043896[p59_addedKey__56_comb[111:104]];
  assign p59_array_index_2054731_comb = p58_literal_2043896[p59_addedKey__56_comb[103:96]];
  assign p59_array_index_2054732_comb = p58_literal_2043896[p59_addedKey__56_comb[95:88]];
  assign p59_array_index_2054733_comb = p58_literal_2043896[p59_addedKey__56_comb[87:80]];
  assign p59_array_index_2054735_comb = p58_literal_2043896[p59_addedKey__56_comb[71:64]];
  assign p59_array_index_2054737_comb = p58_literal_2043896[p59_addedKey__56_comb[55:48]];
  assign p59_array_index_2054738_comb = p58_literal_2043896[p59_addedKey__56_comb[47:40]];
  assign p59_array_index_2054739_comb = p58_literal_2043896[p59_addedKey__56_comb[39:32]];
  assign p59_array_index_2054740_comb = p58_literal_2043896[p59_addedKey__56_comb[31:24]];
  assign p59_array_index_2054741_comb = p58_literal_2043896[p59_addedKey__56_comb[23:16]];
  assign p59_array_index_2054742_comb = p58_literal_2043896[p59_addedKey__56_comb[15:8]];
  assign p59_array_index_2054744_comb = p58_literal_2043910[p59_array_index_2054728_comb];
  assign p59_array_index_2054745_comb = p58_literal_2043912[p59_array_index_2054729_comb];
  assign p59_array_index_2054746_comb = p58_literal_2043914[p59_array_index_2054730_comb];
  assign p59_array_index_2054747_comb = p58_literal_2043916[p59_array_index_2054731_comb];
  assign p59_array_index_2054748_comb = p58_literal_2043918[p59_array_index_2054732_comb];
  assign p59_array_index_2054749_comb = p58_literal_2043920[p59_array_index_2054733_comb];
  assign p59_array_index_2054750_comb = p58_literal_2043896[p59_addedKey__56_comb[79:72]];
  assign p59_array_index_2054752_comb = p58_literal_2043896[p59_addedKey__56_comb[63:56]];
  assign p59_res7__768_comb = p59_array_index_2054744_comb ^ p59_array_index_2054745_comb ^ p59_array_index_2054746_comb ^ p59_array_index_2054747_comb ^ p59_array_index_2054748_comb ^ p59_array_index_2054749_comb ^ p59_array_index_2054750_comb ^ p58_literal_2043923[p59_array_index_2054735_comb] ^ p59_array_index_2054752_comb ^ p58_literal_2043920[p59_array_index_2054737_comb] ^ p58_literal_2043918[p59_array_index_2054738_comb] ^ p58_literal_2043916[p59_array_index_2054739_comb] ^ p58_literal_2043914[p59_array_index_2054740_comb] ^ p58_literal_2043912[p59_array_index_2054741_comb] ^ p58_literal_2043910[p59_array_index_2054742_comb] ^ p58_literal_2043896[p59_addedKey__56_comb[7:0]];
  assign p59_array_index_2054761_comb = p58_literal_2043910[p59_res7__768_comb];
  assign p59_array_index_2054762_comb = p58_literal_2043912[p59_array_index_2054728_comb];
  assign p59_array_index_2054763_comb = p58_literal_2043914[p59_array_index_2054729_comb];
  assign p59_array_index_2054764_comb = p58_literal_2043916[p59_array_index_2054730_comb];
  assign p59_array_index_2054765_comb = p58_literal_2043918[p59_array_index_2054731_comb];
  assign p59_array_index_2054766_comb = p58_literal_2043920[p59_array_index_2054732_comb];
  assign p59_res7__770_comb = p59_array_index_2054761_comb ^ p59_array_index_2054762_comb ^ p59_array_index_2054763_comb ^ p59_array_index_2054764_comb ^ p59_array_index_2054765_comb ^ p59_array_index_2054766_comb ^ p59_array_index_2054733_comb ^ p58_literal_2043923[p59_array_index_2054750_comb] ^ p59_array_index_2054735_comb ^ p58_literal_2043920[p59_array_index_2054752_comb] ^ p58_literal_2043918[p59_array_index_2054737_comb] ^ p58_literal_2043916[p59_array_index_2054738_comb] ^ p58_literal_2043914[p59_array_index_2054739_comb] ^ p58_literal_2043912[p59_array_index_2054740_comb] ^ p58_literal_2043910[p59_array_index_2054741_comb] ^ p59_array_index_2054742_comb;
  assign p59_array_index_2054776_comb = p58_literal_2043912[p59_res7__768_comb];
  assign p59_array_index_2054777_comb = p58_literal_2043914[p59_array_index_2054728_comb];
  assign p59_array_index_2054778_comb = p58_literal_2043916[p59_array_index_2054729_comb];
  assign p59_array_index_2054779_comb = p58_literal_2043918[p59_array_index_2054730_comb];
  assign p59_array_index_2054780_comb = p58_literal_2043920[p59_array_index_2054731_comb];
  assign p59_res7__772_comb = p58_literal_2043910[p59_res7__770_comb] ^ p59_array_index_2054776_comb ^ p59_array_index_2054777_comb ^ p59_array_index_2054778_comb ^ p59_array_index_2054779_comb ^ p59_array_index_2054780_comb ^ p59_array_index_2054732_comb ^ p58_literal_2043923[p59_array_index_2054733_comb] ^ p59_array_index_2054750_comb ^ p58_literal_2043920[p59_array_index_2054735_comb] ^ p58_literal_2043918[p59_array_index_2054752_comb] ^ p58_literal_2043916[p59_array_index_2054737_comb] ^ p58_literal_2043914[p59_array_index_2054738_comb] ^ p58_literal_2043912[p59_array_index_2054739_comb] ^ p58_literal_2043910[p59_array_index_2054740_comb] ^ p59_array_index_2054741_comb;
  assign p59_array_index_2054790_comb = p58_literal_2043912[p59_res7__770_comb];
  assign p59_array_index_2054791_comb = p58_literal_2043914[p59_res7__768_comb];
  assign p59_array_index_2054792_comb = p58_literal_2043916[p59_array_index_2054728_comb];
  assign p59_array_index_2054793_comb = p58_literal_2043918[p59_array_index_2054729_comb];
  assign p59_array_index_2054794_comb = p58_literal_2043920[p59_array_index_2054730_comb];
  assign p59_res7__774_comb = p58_literal_2043910[p59_res7__772_comb] ^ p59_array_index_2054790_comb ^ p59_array_index_2054791_comb ^ p59_array_index_2054792_comb ^ p59_array_index_2054793_comb ^ p59_array_index_2054794_comb ^ p59_array_index_2054731_comb ^ p58_literal_2043923[p59_array_index_2054732_comb] ^ p59_array_index_2054733_comb ^ p58_literal_2043920[p59_array_index_2054750_comb] ^ p58_literal_2043918[p59_array_index_2054735_comb] ^ p58_literal_2043916[p59_array_index_2054752_comb] ^ p58_literal_2043914[p59_array_index_2054737_comb] ^ p58_literal_2043912[p59_array_index_2054738_comb] ^ p58_literal_2043910[p59_array_index_2054739_comb] ^ p59_array_index_2054740_comb;

  // Registers for pipe stage 59:
  reg [127:0] p59_encoded;
  reg [127:0] p59_bit_slice_2043893;
  reg [127:0] p59_bit_slice_2044018;
  reg [127:0] p59_k3;
  reg [127:0] p59_k2;
  reg [127:0] p59_k5;
  reg [127:0] p59_k4;
  reg [127:0] p59_k7;
  reg [127:0] p59_k6;
  reg [7:0] p59_array_index_2054728;
  reg [7:0] p59_array_index_2054729;
  reg [7:0] p59_array_index_2054730;
  reg [7:0] p59_array_index_2054731;
  reg [7:0] p59_array_index_2054732;
  reg [7:0] p59_array_index_2054733;
  reg [7:0] p59_array_index_2054735;
  reg [7:0] p59_array_index_2054737;
  reg [7:0] p59_array_index_2054738;
  reg [7:0] p59_array_index_2054739;
  reg [7:0] p59_array_index_2054744;
  reg [7:0] p59_array_index_2054745;
  reg [7:0] p59_array_index_2054746;
  reg [7:0] p59_array_index_2054747;
  reg [7:0] p59_array_index_2054748;
  reg [7:0] p59_array_index_2054749;
  reg [7:0] p59_array_index_2054750;
  reg [7:0] p59_array_index_2054752;
  reg [7:0] p59_res7__768;
  reg [7:0] p59_array_index_2054761;
  reg [7:0] p59_array_index_2054762;
  reg [7:0] p59_array_index_2054763;
  reg [7:0] p59_array_index_2054764;
  reg [7:0] p59_array_index_2054765;
  reg [7:0] p59_array_index_2054766;
  reg [7:0] p59_res7__770;
  reg [7:0] p59_array_index_2054776;
  reg [7:0] p59_array_index_2054777;
  reg [7:0] p59_array_index_2054778;
  reg [7:0] p59_array_index_2054779;
  reg [7:0] p59_array_index_2054780;
  reg [7:0] p59_res7__772;
  reg [7:0] p59_array_index_2054790;
  reg [7:0] p59_array_index_2054791;
  reg [7:0] p59_array_index_2054792;
  reg [7:0] p59_array_index_2054793;
  reg [7:0] p59_array_index_2054794;
  reg [7:0] p59_res7__774;
  reg [7:0] p60_literal_2043896[256];
  reg [7:0] p60_literal_2043910[256];
  reg [7:0] p60_literal_2043912[256];
  reg [7:0] p60_literal_2043914[256];
  reg [7:0] p60_literal_2043916[256];
  reg [7:0] p60_literal_2043918[256];
  reg [7:0] p60_literal_2043920[256];
  reg [7:0] p60_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p59_encoded <= p58_encoded;
    p59_bit_slice_2043893 <= p58_bit_slice_2043893;
    p59_bit_slice_2044018 <= p58_bit_slice_2044018;
    p59_k3 <= p58_k3;
    p59_k2 <= p58_k2;
    p59_k5 <= p58_k5;
    p59_k4 <= p58_k4;
    p59_k7 <= p58_k7;
    p59_k6 <= p59_k6_comb;
    p59_array_index_2054728 <= p59_array_index_2054728_comb;
    p59_array_index_2054729 <= p59_array_index_2054729_comb;
    p59_array_index_2054730 <= p59_array_index_2054730_comb;
    p59_array_index_2054731 <= p59_array_index_2054731_comb;
    p59_array_index_2054732 <= p59_array_index_2054732_comb;
    p59_array_index_2054733 <= p59_array_index_2054733_comb;
    p59_array_index_2054735 <= p59_array_index_2054735_comb;
    p59_array_index_2054737 <= p59_array_index_2054737_comb;
    p59_array_index_2054738 <= p59_array_index_2054738_comb;
    p59_array_index_2054739 <= p59_array_index_2054739_comb;
    p59_array_index_2054744 <= p59_array_index_2054744_comb;
    p59_array_index_2054745 <= p59_array_index_2054745_comb;
    p59_array_index_2054746 <= p59_array_index_2054746_comb;
    p59_array_index_2054747 <= p59_array_index_2054747_comb;
    p59_array_index_2054748 <= p59_array_index_2054748_comb;
    p59_array_index_2054749 <= p59_array_index_2054749_comb;
    p59_array_index_2054750 <= p59_array_index_2054750_comb;
    p59_array_index_2054752 <= p59_array_index_2054752_comb;
    p59_res7__768 <= p59_res7__768_comb;
    p59_array_index_2054761 <= p59_array_index_2054761_comb;
    p59_array_index_2054762 <= p59_array_index_2054762_comb;
    p59_array_index_2054763 <= p59_array_index_2054763_comb;
    p59_array_index_2054764 <= p59_array_index_2054764_comb;
    p59_array_index_2054765 <= p59_array_index_2054765_comb;
    p59_array_index_2054766 <= p59_array_index_2054766_comb;
    p59_res7__770 <= p59_res7__770_comb;
    p59_array_index_2054776 <= p59_array_index_2054776_comb;
    p59_array_index_2054777 <= p59_array_index_2054777_comb;
    p59_array_index_2054778 <= p59_array_index_2054778_comb;
    p59_array_index_2054779 <= p59_array_index_2054779_comb;
    p59_array_index_2054780 <= p59_array_index_2054780_comb;
    p59_res7__772 <= p59_res7__772_comb;
    p59_array_index_2054790 <= p59_array_index_2054790_comb;
    p59_array_index_2054791 <= p59_array_index_2054791_comb;
    p59_array_index_2054792 <= p59_array_index_2054792_comb;
    p59_array_index_2054793 <= p59_array_index_2054793_comb;
    p59_array_index_2054794 <= p59_array_index_2054794_comb;
    p59_res7__774 <= p59_res7__774_comb;
    p60_literal_2043896 <= p59_literal_2043896;
    p60_literal_2043910 <= p59_literal_2043910;
    p60_literal_2043912 <= p59_literal_2043912;
    p60_literal_2043914 <= p59_literal_2043914;
    p60_literal_2043916 <= p59_literal_2043916;
    p60_literal_2043918 <= p59_literal_2043918;
    p60_literal_2043920 <= p59_literal_2043920;
    p60_literal_2043923 <= p59_literal_2043923;
  end

  // ===== Pipe stage 60:
  wire [7:0] p60_array_index_2054915_comb;
  wire [7:0] p60_array_index_2054916_comb;
  wire [7:0] p60_array_index_2054917_comb;
  wire [7:0] p60_array_index_2054918_comb;
  wire [7:0] p60_res7__776_comb;
  wire [7:0] p60_array_index_2054928_comb;
  wire [7:0] p60_array_index_2054929_comb;
  wire [7:0] p60_array_index_2054930_comb;
  wire [7:0] p60_array_index_2054931_comb;
  wire [7:0] p60_res7__778_comb;
  wire [7:0] p60_array_index_2054942_comb;
  wire [7:0] p60_array_index_2054943_comb;
  wire [7:0] p60_array_index_2054944_comb;
  wire [7:0] p60_res7__780_comb;
  wire [7:0] p60_array_index_2054954_comb;
  wire [7:0] p60_array_index_2054955_comb;
  wire [7:0] p60_array_index_2054956_comb;
  wire [7:0] p60_res7__782_comb;
  wire [7:0] p60_array_index_2054967_comb;
  wire [7:0] p60_array_index_2054968_comb;
  wire [7:0] p60_res7__784_comb;
  wire [7:0] p60_array_index_2054978_comb;
  wire [7:0] p60_array_index_2054979_comb;
  wire [7:0] p60_res7__786_comb;
  wire [7:0] p60_array_index_2054990_comb;
  wire [7:0] p60_res7__788_comb;
  assign p60_array_index_2054915_comb = p59_literal_2043914[p59_res7__770];
  assign p60_array_index_2054916_comb = p59_literal_2043916[p59_res7__768];
  assign p60_array_index_2054917_comb = p59_literal_2043918[p59_array_index_2054728];
  assign p60_array_index_2054918_comb = p59_literal_2043920[p59_array_index_2054729];
  assign p60_res7__776_comb = p59_literal_2043910[p59_res7__774] ^ p59_literal_2043912[p59_res7__772] ^ p60_array_index_2054915_comb ^ p60_array_index_2054916_comb ^ p60_array_index_2054917_comb ^ p60_array_index_2054918_comb ^ p59_array_index_2054730 ^ p59_literal_2043923[p59_array_index_2054731] ^ p59_array_index_2054732 ^ p59_array_index_2054749 ^ p59_literal_2043918[p59_array_index_2054750] ^ p59_literal_2043916[p59_array_index_2054735] ^ p59_literal_2043914[p59_array_index_2054752] ^ p59_literal_2043912[p59_array_index_2054737] ^ p59_literal_2043910[p59_array_index_2054738] ^ p59_array_index_2054739;
  assign p60_array_index_2054928_comb = p59_literal_2043914[p59_res7__772];
  assign p60_array_index_2054929_comb = p59_literal_2043916[p59_res7__770];
  assign p60_array_index_2054930_comb = p59_literal_2043918[p59_res7__768];
  assign p60_array_index_2054931_comb = p59_literal_2043920[p59_array_index_2054728];
  assign p60_res7__778_comb = p59_literal_2043910[p60_res7__776_comb] ^ p59_literal_2043912[p59_res7__774] ^ p60_array_index_2054928_comb ^ p60_array_index_2054929_comb ^ p60_array_index_2054930_comb ^ p60_array_index_2054931_comb ^ p59_array_index_2054729 ^ p59_literal_2043923[p59_array_index_2054730] ^ p59_array_index_2054731 ^ p59_array_index_2054766 ^ p59_literal_2043918[p59_array_index_2054733] ^ p59_literal_2043916[p59_array_index_2054750] ^ p59_literal_2043914[p59_array_index_2054735] ^ p59_literal_2043912[p59_array_index_2054752] ^ p59_literal_2043910[p59_array_index_2054737] ^ p59_array_index_2054738;
  assign p60_array_index_2054942_comb = p59_literal_2043916[p59_res7__772];
  assign p60_array_index_2054943_comb = p59_literal_2043918[p59_res7__770];
  assign p60_array_index_2054944_comb = p59_literal_2043920[p59_res7__768];
  assign p60_res7__780_comb = p59_literal_2043910[p60_res7__778_comb] ^ p59_literal_2043912[p60_res7__776_comb] ^ p59_literal_2043914[p59_res7__774] ^ p60_array_index_2054942_comb ^ p60_array_index_2054943_comb ^ p60_array_index_2054944_comb ^ p59_array_index_2054728 ^ p59_literal_2043923[p59_array_index_2054729] ^ p59_array_index_2054730 ^ p59_array_index_2054780 ^ p59_array_index_2054748 ^ p59_literal_2043916[p59_array_index_2054733] ^ p59_literal_2043914[p59_array_index_2054750] ^ p59_literal_2043912[p59_array_index_2054735] ^ p59_literal_2043910[p59_array_index_2054752] ^ p59_array_index_2054737;
  assign p60_array_index_2054954_comb = p59_literal_2043916[p59_res7__774];
  assign p60_array_index_2054955_comb = p59_literal_2043918[p59_res7__772];
  assign p60_array_index_2054956_comb = p59_literal_2043920[p59_res7__770];
  assign p60_res7__782_comb = p59_literal_2043910[p60_res7__780_comb] ^ p59_literal_2043912[p60_res7__778_comb] ^ p59_literal_2043914[p60_res7__776_comb] ^ p60_array_index_2054954_comb ^ p60_array_index_2054955_comb ^ p60_array_index_2054956_comb ^ p59_res7__768 ^ p59_literal_2043923[p59_array_index_2054728] ^ p59_array_index_2054729 ^ p59_array_index_2054794 ^ p59_array_index_2054765 ^ p59_literal_2043916[p59_array_index_2054732] ^ p59_literal_2043914[p59_array_index_2054733] ^ p59_literal_2043912[p59_array_index_2054750] ^ p59_literal_2043910[p59_array_index_2054735] ^ p59_array_index_2054752;
  assign p60_array_index_2054967_comb = p59_literal_2043918[p59_res7__774];
  assign p60_array_index_2054968_comb = p59_literal_2043920[p59_res7__772];
  assign p60_res7__784_comb = p59_literal_2043910[p60_res7__782_comb] ^ p59_literal_2043912[p60_res7__780_comb] ^ p59_literal_2043914[p60_res7__778_comb] ^ p59_literal_2043916[p60_res7__776_comb] ^ p60_array_index_2054967_comb ^ p60_array_index_2054968_comb ^ p59_res7__770 ^ p59_literal_2043923[p59_res7__768] ^ p59_array_index_2054728 ^ p60_array_index_2054918_comb ^ p59_array_index_2054779 ^ p59_array_index_2054747 ^ p59_literal_2043914[p59_array_index_2054732] ^ p59_literal_2043912[p59_array_index_2054733] ^ p59_literal_2043910[p59_array_index_2054750] ^ p59_array_index_2054735;
  assign p60_array_index_2054978_comb = p59_literal_2043918[p60_res7__776_comb];
  assign p60_array_index_2054979_comb = p59_literal_2043920[p59_res7__774];
  assign p60_res7__786_comb = p59_literal_2043910[p60_res7__784_comb] ^ p59_literal_2043912[p60_res7__782_comb] ^ p59_literal_2043914[p60_res7__780_comb] ^ p59_literal_2043916[p60_res7__778_comb] ^ p60_array_index_2054978_comb ^ p60_array_index_2054979_comb ^ p59_res7__772 ^ p59_literal_2043923[p59_res7__770] ^ p59_res7__768 ^ p60_array_index_2054931_comb ^ p59_array_index_2054793 ^ p59_array_index_2054764 ^ p59_literal_2043914[p59_array_index_2054731] ^ p59_literal_2043912[p59_array_index_2054732] ^ p59_literal_2043910[p59_array_index_2054733] ^ p59_array_index_2054750;
  assign p60_array_index_2054990_comb = p59_literal_2043920[p60_res7__776_comb];
  assign p60_res7__788_comb = p59_literal_2043910[p60_res7__786_comb] ^ p59_literal_2043912[p60_res7__784_comb] ^ p59_literal_2043914[p60_res7__782_comb] ^ p59_literal_2043916[p60_res7__780_comb] ^ p59_literal_2043918[p60_res7__778_comb] ^ p60_array_index_2054990_comb ^ p59_res7__774 ^ p59_literal_2043923[p59_res7__772] ^ p59_res7__770 ^ p60_array_index_2054944_comb ^ p60_array_index_2054917_comb ^ p59_array_index_2054778 ^ p59_array_index_2054746 ^ p59_literal_2043912[p59_array_index_2054731] ^ p59_literal_2043910[p59_array_index_2054732] ^ p59_array_index_2054733;

  // Registers for pipe stage 60:
  reg [127:0] p60_encoded;
  reg [127:0] p60_bit_slice_2043893;
  reg [127:0] p60_bit_slice_2044018;
  reg [127:0] p60_k3;
  reg [127:0] p60_k2;
  reg [127:0] p60_k5;
  reg [127:0] p60_k4;
  reg [127:0] p60_k7;
  reg [127:0] p60_k6;
  reg [7:0] p60_array_index_2054728;
  reg [7:0] p60_array_index_2054729;
  reg [7:0] p60_array_index_2054730;
  reg [7:0] p60_array_index_2054731;
  reg [7:0] p60_array_index_2054732;
  reg [7:0] p60_array_index_2054744;
  reg [7:0] p60_array_index_2054745;
  reg [7:0] p60_res7__768;
  reg [7:0] p60_array_index_2054761;
  reg [7:0] p60_array_index_2054762;
  reg [7:0] p60_array_index_2054763;
  reg [7:0] p60_res7__770;
  reg [7:0] p60_array_index_2054776;
  reg [7:0] p60_array_index_2054777;
  reg [7:0] p60_res7__772;
  reg [7:0] p60_array_index_2054790;
  reg [7:0] p60_array_index_2054791;
  reg [7:0] p60_array_index_2054792;
  reg [7:0] p60_res7__774;
  reg [7:0] p60_array_index_2054915;
  reg [7:0] p60_array_index_2054916;
  reg [7:0] p60_res7__776;
  reg [7:0] p60_array_index_2054928;
  reg [7:0] p60_array_index_2054929;
  reg [7:0] p60_array_index_2054930;
  reg [7:0] p60_res7__778;
  reg [7:0] p60_array_index_2054942;
  reg [7:0] p60_array_index_2054943;
  reg [7:0] p60_res7__780;
  reg [7:0] p60_array_index_2054954;
  reg [7:0] p60_array_index_2054955;
  reg [7:0] p60_array_index_2054956;
  reg [7:0] p60_res7__782;
  reg [7:0] p60_array_index_2054967;
  reg [7:0] p60_array_index_2054968;
  reg [7:0] p60_res7__784;
  reg [7:0] p60_array_index_2054978;
  reg [7:0] p60_array_index_2054979;
  reg [7:0] p60_res7__786;
  reg [7:0] p60_array_index_2054990;
  reg [7:0] p60_res7__788;
  reg [7:0] p61_literal_2043896[256];
  reg [7:0] p61_literal_2043910[256];
  reg [7:0] p61_literal_2043912[256];
  reg [7:0] p61_literal_2043914[256];
  reg [7:0] p61_literal_2043916[256];
  reg [7:0] p61_literal_2043918[256];
  reg [7:0] p61_literal_2043920[256];
  reg [7:0] p61_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p60_encoded <= p59_encoded;
    p60_bit_slice_2043893 <= p59_bit_slice_2043893;
    p60_bit_slice_2044018 <= p59_bit_slice_2044018;
    p60_k3 <= p59_k3;
    p60_k2 <= p59_k2;
    p60_k5 <= p59_k5;
    p60_k4 <= p59_k4;
    p60_k7 <= p59_k7;
    p60_k6 <= p59_k6;
    p60_array_index_2054728 <= p59_array_index_2054728;
    p60_array_index_2054729 <= p59_array_index_2054729;
    p60_array_index_2054730 <= p59_array_index_2054730;
    p60_array_index_2054731 <= p59_array_index_2054731;
    p60_array_index_2054732 <= p59_array_index_2054732;
    p60_array_index_2054744 <= p59_array_index_2054744;
    p60_array_index_2054745 <= p59_array_index_2054745;
    p60_res7__768 <= p59_res7__768;
    p60_array_index_2054761 <= p59_array_index_2054761;
    p60_array_index_2054762 <= p59_array_index_2054762;
    p60_array_index_2054763 <= p59_array_index_2054763;
    p60_res7__770 <= p59_res7__770;
    p60_array_index_2054776 <= p59_array_index_2054776;
    p60_array_index_2054777 <= p59_array_index_2054777;
    p60_res7__772 <= p59_res7__772;
    p60_array_index_2054790 <= p59_array_index_2054790;
    p60_array_index_2054791 <= p59_array_index_2054791;
    p60_array_index_2054792 <= p59_array_index_2054792;
    p60_res7__774 <= p59_res7__774;
    p60_array_index_2054915 <= p60_array_index_2054915_comb;
    p60_array_index_2054916 <= p60_array_index_2054916_comb;
    p60_res7__776 <= p60_res7__776_comb;
    p60_array_index_2054928 <= p60_array_index_2054928_comb;
    p60_array_index_2054929 <= p60_array_index_2054929_comb;
    p60_array_index_2054930 <= p60_array_index_2054930_comb;
    p60_res7__778 <= p60_res7__778_comb;
    p60_array_index_2054942 <= p60_array_index_2054942_comb;
    p60_array_index_2054943 <= p60_array_index_2054943_comb;
    p60_res7__780 <= p60_res7__780_comb;
    p60_array_index_2054954 <= p60_array_index_2054954_comb;
    p60_array_index_2054955 <= p60_array_index_2054955_comb;
    p60_array_index_2054956 <= p60_array_index_2054956_comb;
    p60_res7__782 <= p60_res7__782_comb;
    p60_array_index_2054967 <= p60_array_index_2054967_comb;
    p60_array_index_2054968 <= p60_array_index_2054968_comb;
    p60_res7__784 <= p60_res7__784_comb;
    p60_array_index_2054978 <= p60_array_index_2054978_comb;
    p60_array_index_2054979 <= p60_array_index_2054979_comb;
    p60_res7__786 <= p60_res7__786_comb;
    p60_array_index_2054990 <= p60_array_index_2054990_comb;
    p60_res7__788 <= p60_res7__788_comb;
    p61_literal_2043896 <= p60_literal_2043896;
    p61_literal_2043910 <= p60_literal_2043910;
    p61_literal_2043912 <= p60_literal_2043912;
    p61_literal_2043914 <= p60_literal_2043914;
    p61_literal_2043916 <= p60_literal_2043916;
    p61_literal_2043918 <= p60_literal_2043918;
    p61_literal_2043920 <= p60_literal_2043920;
    p61_literal_2043923 <= p60_literal_2043923;
  end

  // ===== Pipe stage 61:
  wire [7:0] p61_array_index_2055116_comb;
  wire [7:0] p61_res7__790_comb;
  wire [7:0] p61_res7__792_comb;
  wire [7:0] p61_res7__794_comb;
  wire [7:0] p61_res7__796_comb;
  wire [7:0] p61_res7__798_comb;
  wire [127:0] p61_res__24_comb;
  wire [127:0] p61_xor_2055156_comb;
  wire [127:0] p61_addedKey__57_comb;
  wire [7:0] p61_array_index_2055172_comb;
  wire [7:0] p61_array_index_2055173_comb;
  wire [7:0] p61_array_index_2055174_comb;
  wire [7:0] p61_array_index_2055175_comb;
  wire [7:0] p61_array_index_2055176_comb;
  wire [7:0] p61_array_index_2055177_comb;
  wire [7:0] p61_array_index_2055179_comb;
  wire [7:0] p61_array_index_2055181_comb;
  wire [7:0] p61_array_index_2055182_comb;
  wire [7:0] p61_array_index_2055183_comb;
  wire [7:0] p61_array_index_2055184_comb;
  wire [7:0] p61_array_index_2055185_comb;
  wire [7:0] p61_array_index_2055186_comb;
  wire [7:0] p61_array_index_2055188_comb;
  wire [7:0] p61_array_index_2055189_comb;
  wire [7:0] p61_array_index_2055190_comb;
  wire [7:0] p61_array_index_2055191_comb;
  wire [7:0] p61_array_index_2055192_comb;
  wire [7:0] p61_array_index_2055193_comb;
  wire [7:0] p61_array_index_2055194_comb;
  wire [7:0] p61_array_index_2055196_comb;
  wire [7:0] p61_res7__800_comb;
  assign p61_array_index_2055116_comb = p60_literal_2043920[p60_res7__778];
  assign p61_res7__790_comb = p60_literal_2043910[p60_res7__788] ^ p60_literal_2043912[p60_res7__786] ^ p60_literal_2043914[p60_res7__784] ^ p60_literal_2043916[p60_res7__782] ^ p60_literal_2043918[p60_res7__780] ^ p61_array_index_2055116_comb ^ p60_res7__776 ^ p60_literal_2043923[p60_res7__774] ^ p60_res7__772 ^ p60_array_index_2054956 ^ p60_array_index_2054930 ^ p60_array_index_2054792 ^ p60_array_index_2054763 ^ p60_literal_2043912[p60_array_index_2054730] ^ p60_literal_2043910[p60_array_index_2054731] ^ p60_array_index_2054732;
  assign p61_res7__792_comb = p60_literal_2043910[p61_res7__790_comb] ^ p60_literal_2043912[p60_res7__788] ^ p60_literal_2043914[p60_res7__786] ^ p60_literal_2043916[p60_res7__784] ^ p60_literal_2043918[p60_res7__782] ^ p60_literal_2043920[p60_res7__780] ^ p60_res7__778 ^ p60_literal_2043923[p60_res7__776] ^ p60_res7__774 ^ p60_array_index_2054968 ^ p60_array_index_2054943 ^ p60_array_index_2054916 ^ p60_array_index_2054777 ^ p60_array_index_2054745 ^ p60_literal_2043910[p60_array_index_2054730] ^ p60_array_index_2054731;
  assign p61_res7__794_comb = p60_literal_2043910[p61_res7__792_comb] ^ p60_literal_2043912[p61_res7__790_comb] ^ p60_literal_2043914[p60_res7__788] ^ p60_literal_2043916[p60_res7__786] ^ p60_literal_2043918[p60_res7__784] ^ p60_literal_2043920[p60_res7__782] ^ p60_res7__780 ^ p60_literal_2043923[p60_res7__778] ^ p60_res7__776 ^ p60_array_index_2054979 ^ p60_array_index_2054955 ^ p60_array_index_2054929 ^ p60_array_index_2054791 ^ p60_array_index_2054762 ^ p60_literal_2043910[p60_array_index_2054729] ^ p60_array_index_2054730;
  assign p61_res7__796_comb = p60_literal_2043910[p61_res7__794_comb] ^ p60_literal_2043912[p61_res7__792_comb] ^ p60_literal_2043914[p61_res7__790_comb] ^ p60_literal_2043916[p60_res7__788] ^ p60_literal_2043918[p60_res7__786] ^ p60_literal_2043920[p60_res7__784] ^ p60_res7__782 ^ p60_literal_2043923[p60_res7__780] ^ p60_res7__778 ^ p60_array_index_2054990 ^ p60_array_index_2054967 ^ p60_array_index_2054942 ^ p60_array_index_2054915 ^ p60_array_index_2054776 ^ p60_array_index_2054744 ^ p60_array_index_2054729;
  assign p61_res7__798_comb = p60_literal_2043910[p61_res7__796_comb] ^ p60_literal_2043912[p61_res7__794_comb] ^ p60_literal_2043914[p61_res7__792_comb] ^ p60_literal_2043916[p61_res7__790_comb] ^ p60_literal_2043918[p60_res7__788] ^ p60_literal_2043920[p60_res7__786] ^ p60_res7__784 ^ p60_literal_2043923[p60_res7__782] ^ p60_res7__780 ^ p61_array_index_2055116_comb ^ p60_array_index_2054978 ^ p60_array_index_2054954 ^ p60_array_index_2054928 ^ p60_array_index_2054790 ^ p60_array_index_2054761 ^ p60_array_index_2054728;
  assign p61_res__24_comb = {p61_res7__798_comb, p61_res7__796_comb, p61_res7__794_comb, p61_res7__792_comb, p61_res7__790_comb, p60_res7__788, p60_res7__786, p60_res7__784, p60_res7__782, p60_res7__780, p60_res7__778, p60_res7__776, p60_res7__774, p60_res7__772, p60_res7__770, p60_res7__768};
  assign p61_xor_2055156_comb = p61_res__24_comb ^ p60_k7;
  assign p61_addedKey__57_comb = p61_xor_2055156_comb ^ 128'h056c_b6de_319f_0eeb_8e80_9963_10f6_951a;
  assign p61_array_index_2055172_comb = p60_literal_2043896[p61_addedKey__57_comb[127:120]];
  assign p61_array_index_2055173_comb = p60_literal_2043896[p61_addedKey__57_comb[119:112]];
  assign p61_array_index_2055174_comb = p60_literal_2043896[p61_addedKey__57_comb[111:104]];
  assign p61_array_index_2055175_comb = p60_literal_2043896[p61_addedKey__57_comb[103:96]];
  assign p61_array_index_2055176_comb = p60_literal_2043896[p61_addedKey__57_comb[95:88]];
  assign p61_array_index_2055177_comb = p60_literal_2043896[p61_addedKey__57_comb[87:80]];
  assign p61_array_index_2055179_comb = p60_literal_2043896[p61_addedKey__57_comb[71:64]];
  assign p61_array_index_2055181_comb = p60_literal_2043896[p61_addedKey__57_comb[55:48]];
  assign p61_array_index_2055182_comb = p60_literal_2043896[p61_addedKey__57_comb[47:40]];
  assign p61_array_index_2055183_comb = p60_literal_2043896[p61_addedKey__57_comb[39:32]];
  assign p61_array_index_2055184_comb = p60_literal_2043896[p61_addedKey__57_comb[31:24]];
  assign p61_array_index_2055185_comb = p60_literal_2043896[p61_addedKey__57_comb[23:16]];
  assign p61_array_index_2055186_comb = p60_literal_2043896[p61_addedKey__57_comb[15:8]];
  assign p61_array_index_2055188_comb = p60_literal_2043910[p61_array_index_2055172_comb];
  assign p61_array_index_2055189_comb = p60_literal_2043912[p61_array_index_2055173_comb];
  assign p61_array_index_2055190_comb = p60_literal_2043914[p61_array_index_2055174_comb];
  assign p61_array_index_2055191_comb = p60_literal_2043916[p61_array_index_2055175_comb];
  assign p61_array_index_2055192_comb = p60_literal_2043918[p61_array_index_2055176_comb];
  assign p61_array_index_2055193_comb = p60_literal_2043920[p61_array_index_2055177_comb];
  assign p61_array_index_2055194_comb = p60_literal_2043896[p61_addedKey__57_comb[79:72]];
  assign p61_array_index_2055196_comb = p60_literal_2043896[p61_addedKey__57_comb[63:56]];
  assign p61_res7__800_comb = p61_array_index_2055188_comb ^ p61_array_index_2055189_comb ^ p61_array_index_2055190_comb ^ p61_array_index_2055191_comb ^ p61_array_index_2055192_comb ^ p61_array_index_2055193_comb ^ p61_array_index_2055194_comb ^ p60_literal_2043923[p61_array_index_2055179_comb] ^ p61_array_index_2055196_comb ^ p60_literal_2043920[p61_array_index_2055181_comb] ^ p60_literal_2043918[p61_array_index_2055182_comb] ^ p60_literal_2043916[p61_array_index_2055183_comb] ^ p60_literal_2043914[p61_array_index_2055184_comb] ^ p60_literal_2043912[p61_array_index_2055185_comb] ^ p60_literal_2043910[p61_array_index_2055186_comb] ^ p60_literal_2043896[p61_addedKey__57_comb[7:0]];

  // Registers for pipe stage 61:
  reg [127:0] p61_encoded;
  reg [127:0] p61_bit_slice_2043893;
  reg [127:0] p61_bit_slice_2044018;
  reg [127:0] p61_k3;
  reg [127:0] p61_k2;
  reg [127:0] p61_k5;
  reg [127:0] p61_k4;
  reg [127:0] p61_k7;
  reg [127:0] p61_k6;
  reg [127:0] p61_xor_2055156;
  reg [7:0] p61_array_index_2055172;
  reg [7:0] p61_array_index_2055173;
  reg [7:0] p61_array_index_2055174;
  reg [7:0] p61_array_index_2055175;
  reg [7:0] p61_array_index_2055176;
  reg [7:0] p61_array_index_2055177;
  reg [7:0] p61_array_index_2055179;
  reg [7:0] p61_array_index_2055181;
  reg [7:0] p61_array_index_2055182;
  reg [7:0] p61_array_index_2055183;
  reg [7:0] p61_array_index_2055184;
  reg [7:0] p61_array_index_2055185;
  reg [7:0] p61_array_index_2055186;
  reg [7:0] p61_array_index_2055188;
  reg [7:0] p61_array_index_2055189;
  reg [7:0] p61_array_index_2055190;
  reg [7:0] p61_array_index_2055191;
  reg [7:0] p61_array_index_2055192;
  reg [7:0] p61_array_index_2055193;
  reg [7:0] p61_array_index_2055194;
  reg [7:0] p61_array_index_2055196;
  reg [7:0] p61_res7__800;
  reg [7:0] p62_literal_2043896[256];
  reg [7:0] p62_literal_2043910[256];
  reg [7:0] p62_literal_2043912[256];
  reg [7:0] p62_literal_2043914[256];
  reg [7:0] p62_literal_2043916[256];
  reg [7:0] p62_literal_2043918[256];
  reg [7:0] p62_literal_2043920[256];
  reg [7:0] p62_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p61_encoded <= p60_encoded;
    p61_bit_slice_2043893 <= p60_bit_slice_2043893;
    p61_bit_slice_2044018 <= p60_bit_slice_2044018;
    p61_k3 <= p60_k3;
    p61_k2 <= p60_k2;
    p61_k5 <= p60_k5;
    p61_k4 <= p60_k4;
    p61_k7 <= p60_k7;
    p61_k6 <= p60_k6;
    p61_xor_2055156 <= p61_xor_2055156_comb;
    p61_array_index_2055172 <= p61_array_index_2055172_comb;
    p61_array_index_2055173 <= p61_array_index_2055173_comb;
    p61_array_index_2055174 <= p61_array_index_2055174_comb;
    p61_array_index_2055175 <= p61_array_index_2055175_comb;
    p61_array_index_2055176 <= p61_array_index_2055176_comb;
    p61_array_index_2055177 <= p61_array_index_2055177_comb;
    p61_array_index_2055179 <= p61_array_index_2055179_comb;
    p61_array_index_2055181 <= p61_array_index_2055181_comb;
    p61_array_index_2055182 <= p61_array_index_2055182_comb;
    p61_array_index_2055183 <= p61_array_index_2055183_comb;
    p61_array_index_2055184 <= p61_array_index_2055184_comb;
    p61_array_index_2055185 <= p61_array_index_2055185_comb;
    p61_array_index_2055186 <= p61_array_index_2055186_comb;
    p61_array_index_2055188 <= p61_array_index_2055188_comb;
    p61_array_index_2055189 <= p61_array_index_2055189_comb;
    p61_array_index_2055190 <= p61_array_index_2055190_comb;
    p61_array_index_2055191 <= p61_array_index_2055191_comb;
    p61_array_index_2055192 <= p61_array_index_2055192_comb;
    p61_array_index_2055193 <= p61_array_index_2055193_comb;
    p61_array_index_2055194 <= p61_array_index_2055194_comb;
    p61_array_index_2055196 <= p61_array_index_2055196_comb;
    p61_res7__800 <= p61_res7__800_comb;
    p62_literal_2043896 <= p61_literal_2043896;
    p62_literal_2043910 <= p61_literal_2043910;
    p62_literal_2043912 <= p61_literal_2043912;
    p62_literal_2043914 <= p61_literal_2043914;
    p62_literal_2043916 <= p61_literal_2043916;
    p62_literal_2043918 <= p61_literal_2043918;
    p62_literal_2043920 <= p61_literal_2043920;
    p62_literal_2043923 <= p61_literal_2043923;
  end

  // ===== Pipe stage 62:
  wire [7:0] p62_array_index_2055285_comb;
  wire [7:0] p62_array_index_2055286_comb;
  wire [7:0] p62_array_index_2055287_comb;
  wire [7:0] p62_array_index_2055288_comb;
  wire [7:0] p62_array_index_2055289_comb;
  wire [7:0] p62_array_index_2055290_comb;
  wire [7:0] p62_res7__802_comb;
  wire [7:0] p62_array_index_2055300_comb;
  wire [7:0] p62_array_index_2055301_comb;
  wire [7:0] p62_array_index_2055302_comb;
  wire [7:0] p62_array_index_2055303_comb;
  wire [7:0] p62_array_index_2055304_comb;
  wire [7:0] p62_res7__804_comb;
  wire [7:0] p62_array_index_2055314_comb;
  wire [7:0] p62_array_index_2055315_comb;
  wire [7:0] p62_array_index_2055316_comb;
  wire [7:0] p62_array_index_2055317_comb;
  wire [7:0] p62_array_index_2055318_comb;
  wire [7:0] p62_res7__806_comb;
  wire [7:0] p62_array_index_2055329_comb;
  wire [7:0] p62_array_index_2055330_comb;
  wire [7:0] p62_array_index_2055331_comb;
  wire [7:0] p62_array_index_2055332_comb;
  wire [7:0] p62_res7__808_comb;
  wire [7:0] p62_array_index_2055342_comb;
  wire [7:0] p62_array_index_2055343_comb;
  wire [7:0] p62_array_index_2055344_comb;
  wire [7:0] p62_array_index_2055345_comb;
  wire [7:0] p62_res7__810_comb;
  wire [7:0] p62_array_index_2055356_comb;
  wire [7:0] p62_array_index_2055357_comb;
  wire [7:0] p62_array_index_2055358_comb;
  wire [7:0] p62_res7__812_comb;
  wire [7:0] p62_array_index_2055368_comb;
  wire [7:0] p62_array_index_2055369_comb;
  wire [7:0] p62_array_index_2055370_comb;
  wire [7:0] p62_res7__814_comb;
  assign p62_array_index_2055285_comb = p61_literal_2043910[p61_res7__800];
  assign p62_array_index_2055286_comb = p61_literal_2043912[p61_array_index_2055172];
  assign p62_array_index_2055287_comb = p61_literal_2043914[p61_array_index_2055173];
  assign p62_array_index_2055288_comb = p61_literal_2043916[p61_array_index_2055174];
  assign p62_array_index_2055289_comb = p61_literal_2043918[p61_array_index_2055175];
  assign p62_array_index_2055290_comb = p61_literal_2043920[p61_array_index_2055176];
  assign p62_res7__802_comb = p62_array_index_2055285_comb ^ p62_array_index_2055286_comb ^ p62_array_index_2055287_comb ^ p62_array_index_2055288_comb ^ p62_array_index_2055289_comb ^ p62_array_index_2055290_comb ^ p61_array_index_2055177 ^ p61_literal_2043923[p61_array_index_2055194] ^ p61_array_index_2055179 ^ p61_literal_2043920[p61_array_index_2055196] ^ p61_literal_2043918[p61_array_index_2055181] ^ p61_literal_2043916[p61_array_index_2055182] ^ p61_literal_2043914[p61_array_index_2055183] ^ p61_literal_2043912[p61_array_index_2055184] ^ p61_literal_2043910[p61_array_index_2055185] ^ p61_array_index_2055186;
  assign p62_array_index_2055300_comb = p61_literal_2043912[p61_res7__800];
  assign p62_array_index_2055301_comb = p61_literal_2043914[p61_array_index_2055172];
  assign p62_array_index_2055302_comb = p61_literal_2043916[p61_array_index_2055173];
  assign p62_array_index_2055303_comb = p61_literal_2043918[p61_array_index_2055174];
  assign p62_array_index_2055304_comb = p61_literal_2043920[p61_array_index_2055175];
  assign p62_res7__804_comb = p61_literal_2043910[p62_res7__802_comb] ^ p62_array_index_2055300_comb ^ p62_array_index_2055301_comb ^ p62_array_index_2055302_comb ^ p62_array_index_2055303_comb ^ p62_array_index_2055304_comb ^ p61_array_index_2055176 ^ p61_literal_2043923[p61_array_index_2055177] ^ p61_array_index_2055194 ^ p61_literal_2043920[p61_array_index_2055179] ^ p61_literal_2043918[p61_array_index_2055196] ^ p61_literal_2043916[p61_array_index_2055181] ^ p61_literal_2043914[p61_array_index_2055182] ^ p61_literal_2043912[p61_array_index_2055183] ^ p61_literal_2043910[p61_array_index_2055184] ^ p61_array_index_2055185;
  assign p62_array_index_2055314_comb = p61_literal_2043912[p62_res7__802_comb];
  assign p62_array_index_2055315_comb = p61_literal_2043914[p61_res7__800];
  assign p62_array_index_2055316_comb = p61_literal_2043916[p61_array_index_2055172];
  assign p62_array_index_2055317_comb = p61_literal_2043918[p61_array_index_2055173];
  assign p62_array_index_2055318_comb = p61_literal_2043920[p61_array_index_2055174];
  assign p62_res7__806_comb = p61_literal_2043910[p62_res7__804_comb] ^ p62_array_index_2055314_comb ^ p62_array_index_2055315_comb ^ p62_array_index_2055316_comb ^ p62_array_index_2055317_comb ^ p62_array_index_2055318_comb ^ p61_array_index_2055175 ^ p61_literal_2043923[p61_array_index_2055176] ^ p61_array_index_2055177 ^ p61_literal_2043920[p61_array_index_2055194] ^ p61_literal_2043918[p61_array_index_2055179] ^ p61_literal_2043916[p61_array_index_2055196] ^ p61_literal_2043914[p61_array_index_2055181] ^ p61_literal_2043912[p61_array_index_2055182] ^ p61_literal_2043910[p61_array_index_2055183] ^ p61_array_index_2055184;
  assign p62_array_index_2055329_comb = p61_literal_2043914[p62_res7__802_comb];
  assign p62_array_index_2055330_comb = p61_literal_2043916[p61_res7__800];
  assign p62_array_index_2055331_comb = p61_literal_2043918[p61_array_index_2055172];
  assign p62_array_index_2055332_comb = p61_literal_2043920[p61_array_index_2055173];
  assign p62_res7__808_comb = p61_literal_2043910[p62_res7__806_comb] ^ p61_literal_2043912[p62_res7__804_comb] ^ p62_array_index_2055329_comb ^ p62_array_index_2055330_comb ^ p62_array_index_2055331_comb ^ p62_array_index_2055332_comb ^ p61_array_index_2055174 ^ p61_literal_2043923[p61_array_index_2055175] ^ p61_array_index_2055176 ^ p61_array_index_2055193 ^ p61_literal_2043918[p61_array_index_2055194] ^ p61_literal_2043916[p61_array_index_2055179] ^ p61_literal_2043914[p61_array_index_2055196] ^ p61_literal_2043912[p61_array_index_2055181] ^ p61_literal_2043910[p61_array_index_2055182] ^ p61_array_index_2055183;
  assign p62_array_index_2055342_comb = p61_literal_2043914[p62_res7__804_comb];
  assign p62_array_index_2055343_comb = p61_literal_2043916[p62_res7__802_comb];
  assign p62_array_index_2055344_comb = p61_literal_2043918[p61_res7__800];
  assign p62_array_index_2055345_comb = p61_literal_2043920[p61_array_index_2055172];
  assign p62_res7__810_comb = p61_literal_2043910[p62_res7__808_comb] ^ p61_literal_2043912[p62_res7__806_comb] ^ p62_array_index_2055342_comb ^ p62_array_index_2055343_comb ^ p62_array_index_2055344_comb ^ p62_array_index_2055345_comb ^ p61_array_index_2055173 ^ p61_literal_2043923[p61_array_index_2055174] ^ p61_array_index_2055175 ^ p62_array_index_2055290_comb ^ p61_literal_2043918[p61_array_index_2055177] ^ p61_literal_2043916[p61_array_index_2055194] ^ p61_literal_2043914[p61_array_index_2055179] ^ p61_literal_2043912[p61_array_index_2055196] ^ p61_literal_2043910[p61_array_index_2055181] ^ p61_array_index_2055182;
  assign p62_array_index_2055356_comb = p61_literal_2043916[p62_res7__804_comb];
  assign p62_array_index_2055357_comb = p61_literal_2043918[p62_res7__802_comb];
  assign p62_array_index_2055358_comb = p61_literal_2043920[p61_res7__800];
  assign p62_res7__812_comb = p61_literal_2043910[p62_res7__810_comb] ^ p61_literal_2043912[p62_res7__808_comb] ^ p61_literal_2043914[p62_res7__806_comb] ^ p62_array_index_2055356_comb ^ p62_array_index_2055357_comb ^ p62_array_index_2055358_comb ^ p61_array_index_2055172 ^ p61_literal_2043923[p61_array_index_2055173] ^ p61_array_index_2055174 ^ p62_array_index_2055304_comb ^ p61_array_index_2055192 ^ p61_literal_2043916[p61_array_index_2055177] ^ p61_literal_2043914[p61_array_index_2055194] ^ p61_literal_2043912[p61_array_index_2055179] ^ p61_literal_2043910[p61_array_index_2055196] ^ p61_array_index_2055181;
  assign p62_array_index_2055368_comb = p61_literal_2043916[p62_res7__806_comb];
  assign p62_array_index_2055369_comb = p61_literal_2043918[p62_res7__804_comb];
  assign p62_array_index_2055370_comb = p61_literal_2043920[p62_res7__802_comb];
  assign p62_res7__814_comb = p61_literal_2043910[p62_res7__812_comb] ^ p61_literal_2043912[p62_res7__810_comb] ^ p61_literal_2043914[p62_res7__808_comb] ^ p62_array_index_2055368_comb ^ p62_array_index_2055369_comb ^ p62_array_index_2055370_comb ^ p61_res7__800 ^ p61_literal_2043923[p61_array_index_2055172] ^ p61_array_index_2055173 ^ p62_array_index_2055318_comb ^ p62_array_index_2055289_comb ^ p61_literal_2043916[p61_array_index_2055176] ^ p61_literal_2043914[p61_array_index_2055177] ^ p61_literal_2043912[p61_array_index_2055194] ^ p61_literal_2043910[p61_array_index_2055179] ^ p61_array_index_2055196;

  // Registers for pipe stage 62:
  reg [127:0] p62_encoded;
  reg [127:0] p62_bit_slice_2043893;
  reg [127:0] p62_bit_slice_2044018;
  reg [127:0] p62_k3;
  reg [127:0] p62_k2;
  reg [127:0] p62_k5;
  reg [127:0] p62_k4;
  reg [127:0] p62_k7;
  reg [127:0] p62_k6;
  reg [127:0] p62_xor_2055156;
  reg [7:0] p62_array_index_2055172;
  reg [7:0] p62_array_index_2055173;
  reg [7:0] p62_array_index_2055174;
  reg [7:0] p62_array_index_2055175;
  reg [7:0] p62_array_index_2055176;
  reg [7:0] p62_array_index_2055177;
  reg [7:0] p62_array_index_2055179;
  reg [7:0] p62_array_index_2055188;
  reg [7:0] p62_array_index_2055189;
  reg [7:0] p62_array_index_2055190;
  reg [7:0] p62_array_index_2055191;
  reg [7:0] p62_array_index_2055194;
  reg [7:0] p62_res7__800;
  reg [7:0] p62_array_index_2055285;
  reg [7:0] p62_array_index_2055286;
  reg [7:0] p62_array_index_2055287;
  reg [7:0] p62_array_index_2055288;
  reg [7:0] p62_res7__802;
  reg [7:0] p62_array_index_2055300;
  reg [7:0] p62_array_index_2055301;
  reg [7:0] p62_array_index_2055302;
  reg [7:0] p62_array_index_2055303;
  reg [7:0] p62_res7__804;
  reg [7:0] p62_array_index_2055314;
  reg [7:0] p62_array_index_2055315;
  reg [7:0] p62_array_index_2055316;
  reg [7:0] p62_array_index_2055317;
  reg [7:0] p62_res7__806;
  reg [7:0] p62_array_index_2055329;
  reg [7:0] p62_array_index_2055330;
  reg [7:0] p62_array_index_2055331;
  reg [7:0] p62_array_index_2055332;
  reg [7:0] p62_res7__808;
  reg [7:0] p62_array_index_2055342;
  reg [7:0] p62_array_index_2055343;
  reg [7:0] p62_array_index_2055344;
  reg [7:0] p62_array_index_2055345;
  reg [7:0] p62_res7__810;
  reg [7:0] p62_array_index_2055356;
  reg [7:0] p62_array_index_2055357;
  reg [7:0] p62_array_index_2055358;
  reg [7:0] p62_res7__812;
  reg [7:0] p62_array_index_2055368;
  reg [7:0] p62_array_index_2055369;
  reg [7:0] p62_array_index_2055370;
  reg [7:0] p62_res7__814;
  reg [7:0] p63_literal_2043896[256];
  reg [7:0] p63_literal_2043910[256];
  reg [7:0] p63_literal_2043912[256];
  reg [7:0] p63_literal_2043914[256];
  reg [7:0] p63_literal_2043916[256];
  reg [7:0] p63_literal_2043918[256];
  reg [7:0] p63_literal_2043920[256];
  reg [7:0] p63_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p62_encoded <= p61_encoded;
    p62_bit_slice_2043893 <= p61_bit_slice_2043893;
    p62_bit_slice_2044018 <= p61_bit_slice_2044018;
    p62_k3 <= p61_k3;
    p62_k2 <= p61_k2;
    p62_k5 <= p61_k5;
    p62_k4 <= p61_k4;
    p62_k7 <= p61_k7;
    p62_k6 <= p61_k6;
    p62_xor_2055156 <= p61_xor_2055156;
    p62_array_index_2055172 <= p61_array_index_2055172;
    p62_array_index_2055173 <= p61_array_index_2055173;
    p62_array_index_2055174 <= p61_array_index_2055174;
    p62_array_index_2055175 <= p61_array_index_2055175;
    p62_array_index_2055176 <= p61_array_index_2055176;
    p62_array_index_2055177 <= p61_array_index_2055177;
    p62_array_index_2055179 <= p61_array_index_2055179;
    p62_array_index_2055188 <= p61_array_index_2055188;
    p62_array_index_2055189 <= p61_array_index_2055189;
    p62_array_index_2055190 <= p61_array_index_2055190;
    p62_array_index_2055191 <= p61_array_index_2055191;
    p62_array_index_2055194 <= p61_array_index_2055194;
    p62_res7__800 <= p61_res7__800;
    p62_array_index_2055285 <= p62_array_index_2055285_comb;
    p62_array_index_2055286 <= p62_array_index_2055286_comb;
    p62_array_index_2055287 <= p62_array_index_2055287_comb;
    p62_array_index_2055288 <= p62_array_index_2055288_comb;
    p62_res7__802 <= p62_res7__802_comb;
    p62_array_index_2055300 <= p62_array_index_2055300_comb;
    p62_array_index_2055301 <= p62_array_index_2055301_comb;
    p62_array_index_2055302 <= p62_array_index_2055302_comb;
    p62_array_index_2055303 <= p62_array_index_2055303_comb;
    p62_res7__804 <= p62_res7__804_comb;
    p62_array_index_2055314 <= p62_array_index_2055314_comb;
    p62_array_index_2055315 <= p62_array_index_2055315_comb;
    p62_array_index_2055316 <= p62_array_index_2055316_comb;
    p62_array_index_2055317 <= p62_array_index_2055317_comb;
    p62_res7__806 <= p62_res7__806_comb;
    p62_array_index_2055329 <= p62_array_index_2055329_comb;
    p62_array_index_2055330 <= p62_array_index_2055330_comb;
    p62_array_index_2055331 <= p62_array_index_2055331_comb;
    p62_array_index_2055332 <= p62_array_index_2055332_comb;
    p62_res7__808 <= p62_res7__808_comb;
    p62_array_index_2055342 <= p62_array_index_2055342_comb;
    p62_array_index_2055343 <= p62_array_index_2055343_comb;
    p62_array_index_2055344 <= p62_array_index_2055344_comb;
    p62_array_index_2055345 <= p62_array_index_2055345_comb;
    p62_res7__810 <= p62_res7__810_comb;
    p62_array_index_2055356 <= p62_array_index_2055356_comb;
    p62_array_index_2055357 <= p62_array_index_2055357_comb;
    p62_array_index_2055358 <= p62_array_index_2055358_comb;
    p62_res7__812 <= p62_res7__812_comb;
    p62_array_index_2055368 <= p62_array_index_2055368_comb;
    p62_array_index_2055369 <= p62_array_index_2055369_comb;
    p62_array_index_2055370 <= p62_array_index_2055370_comb;
    p62_res7__814 <= p62_res7__814_comb;
    p63_literal_2043896 <= p62_literal_2043896;
    p63_literal_2043910 <= p62_literal_2043910;
    p63_literal_2043912 <= p62_literal_2043912;
    p63_literal_2043914 <= p62_literal_2043914;
    p63_literal_2043916 <= p62_literal_2043916;
    p63_literal_2043918 <= p62_literal_2043918;
    p63_literal_2043920 <= p62_literal_2043920;
    p63_literal_2043923 <= p62_literal_2043923;
  end

  // ===== Pipe stage 63:
  wire [7:0] p63_array_index_2055509_comb;
  wire [7:0] p63_array_index_2055510_comb;
  wire [7:0] p63_res7__816_comb;
  wire [7:0] p63_array_index_2055520_comb;
  wire [7:0] p63_array_index_2055521_comb;
  wire [7:0] p63_res7__818_comb;
  wire [7:0] p63_array_index_2055532_comb;
  wire [7:0] p63_res7__820_comb;
  wire [7:0] p63_array_index_2055542_comb;
  wire [7:0] p63_res7__822_comb;
  wire [7:0] p63_res7__824_comb;
  wire [7:0] p63_res7__826_comb;
  wire [7:0] p63_res7__828_comb;
  assign p63_array_index_2055509_comb = p62_literal_2043918[p62_res7__806];
  assign p63_array_index_2055510_comb = p62_literal_2043920[p62_res7__804];
  assign p63_res7__816_comb = p62_literal_2043910[p62_res7__814] ^ p62_literal_2043912[p62_res7__812] ^ p62_literal_2043914[p62_res7__810] ^ p62_literal_2043916[p62_res7__808] ^ p63_array_index_2055509_comb ^ p63_array_index_2055510_comb ^ p62_res7__802 ^ p62_literal_2043923[p62_res7__800] ^ p62_array_index_2055172 ^ p62_array_index_2055332 ^ p62_array_index_2055303 ^ p62_array_index_2055191 ^ p62_literal_2043914[p62_array_index_2055176] ^ p62_literal_2043912[p62_array_index_2055177] ^ p62_literal_2043910[p62_array_index_2055194] ^ p62_array_index_2055179;
  assign p63_array_index_2055520_comb = p62_literal_2043918[p62_res7__808];
  assign p63_array_index_2055521_comb = p62_literal_2043920[p62_res7__806];
  assign p63_res7__818_comb = p62_literal_2043910[p63_res7__816_comb] ^ p62_literal_2043912[p62_res7__814] ^ p62_literal_2043914[p62_res7__812] ^ p62_literal_2043916[p62_res7__810] ^ p63_array_index_2055520_comb ^ p63_array_index_2055521_comb ^ p62_res7__804 ^ p62_literal_2043923[p62_res7__802] ^ p62_res7__800 ^ p62_array_index_2055345 ^ p62_array_index_2055317 ^ p62_array_index_2055288 ^ p62_literal_2043914[p62_array_index_2055175] ^ p62_literal_2043912[p62_array_index_2055176] ^ p62_literal_2043910[p62_array_index_2055177] ^ p62_array_index_2055194;
  assign p63_array_index_2055532_comb = p62_literal_2043920[p62_res7__808];
  assign p63_res7__820_comb = p62_literal_2043910[p63_res7__818_comb] ^ p62_literal_2043912[p63_res7__816_comb] ^ p62_literal_2043914[p62_res7__814] ^ p62_literal_2043916[p62_res7__812] ^ p62_literal_2043918[p62_res7__810] ^ p63_array_index_2055532_comb ^ p62_res7__806 ^ p62_literal_2043923[p62_res7__804] ^ p62_res7__802 ^ p62_array_index_2055358 ^ p62_array_index_2055331 ^ p62_array_index_2055302 ^ p62_array_index_2055190 ^ p62_literal_2043912[p62_array_index_2055175] ^ p62_literal_2043910[p62_array_index_2055176] ^ p62_array_index_2055177;
  assign p63_array_index_2055542_comb = p62_literal_2043920[p62_res7__810];
  assign p63_res7__822_comb = p62_literal_2043910[p63_res7__820_comb] ^ p62_literal_2043912[p63_res7__818_comb] ^ p62_literal_2043914[p63_res7__816_comb] ^ p62_literal_2043916[p62_res7__814] ^ p62_literal_2043918[p62_res7__812] ^ p63_array_index_2055542_comb ^ p62_res7__808 ^ p62_literal_2043923[p62_res7__806] ^ p62_res7__804 ^ p62_array_index_2055370 ^ p62_array_index_2055344 ^ p62_array_index_2055316 ^ p62_array_index_2055287 ^ p62_literal_2043912[p62_array_index_2055174] ^ p62_literal_2043910[p62_array_index_2055175] ^ p62_array_index_2055176;
  assign p63_res7__824_comb = p62_literal_2043910[p63_res7__822_comb] ^ p62_literal_2043912[p63_res7__820_comb] ^ p62_literal_2043914[p63_res7__818_comb] ^ p62_literal_2043916[p63_res7__816_comb] ^ p62_literal_2043918[p62_res7__814] ^ p62_literal_2043920[p62_res7__812] ^ p62_res7__810 ^ p62_literal_2043923[p62_res7__808] ^ p62_res7__806 ^ p63_array_index_2055510_comb ^ p62_array_index_2055357 ^ p62_array_index_2055330 ^ p62_array_index_2055301 ^ p62_array_index_2055189 ^ p62_literal_2043910[p62_array_index_2055174] ^ p62_array_index_2055175;
  assign p63_res7__826_comb = p62_literal_2043910[p63_res7__824_comb] ^ p62_literal_2043912[p63_res7__822_comb] ^ p62_literal_2043914[p63_res7__820_comb] ^ p62_literal_2043916[p63_res7__818_comb] ^ p62_literal_2043918[p63_res7__816_comb] ^ p62_literal_2043920[p62_res7__814] ^ p62_res7__812 ^ p62_literal_2043923[p62_res7__810] ^ p62_res7__808 ^ p63_array_index_2055521_comb ^ p62_array_index_2055369 ^ p62_array_index_2055343 ^ p62_array_index_2055315 ^ p62_array_index_2055286 ^ p62_literal_2043910[p62_array_index_2055173] ^ p62_array_index_2055174;
  assign p63_res7__828_comb = p62_literal_2043910[p63_res7__826_comb] ^ p62_literal_2043912[p63_res7__824_comb] ^ p62_literal_2043914[p63_res7__822_comb] ^ p62_literal_2043916[p63_res7__820_comb] ^ p62_literal_2043918[p63_res7__818_comb] ^ p62_literal_2043920[p63_res7__816_comb] ^ p62_res7__814 ^ p62_literal_2043923[p62_res7__812] ^ p62_res7__810 ^ p63_array_index_2055532_comb ^ p63_array_index_2055509_comb ^ p62_array_index_2055356 ^ p62_array_index_2055329 ^ p62_array_index_2055300 ^ p62_array_index_2055188 ^ p62_array_index_2055173;

  // Registers for pipe stage 63:
  reg [127:0] p63_encoded;
  reg [127:0] p63_bit_slice_2043893;
  reg [127:0] p63_bit_slice_2044018;
  reg [127:0] p63_k3;
  reg [127:0] p63_k2;
  reg [127:0] p63_k5;
  reg [127:0] p63_k4;
  reg [127:0] p63_k7;
  reg [127:0] p63_k6;
  reg [127:0] p63_xor_2055156;
  reg [7:0] p63_array_index_2055172;
  reg [7:0] p63_res7__800;
  reg [7:0] p63_array_index_2055285;
  reg [7:0] p63_res7__802;
  reg [7:0] p63_res7__804;
  reg [7:0] p63_array_index_2055314;
  reg [7:0] p63_res7__806;
  reg [7:0] p63_res7__808;
  reg [7:0] p63_array_index_2055342;
  reg [7:0] p63_res7__810;
  reg [7:0] p63_res7__812;
  reg [7:0] p63_array_index_2055368;
  reg [7:0] p63_res7__814;
  reg [7:0] p63_res7__816;
  reg [7:0] p63_array_index_2055520;
  reg [7:0] p63_res7__818;
  reg [7:0] p63_res7__820;
  reg [7:0] p63_array_index_2055542;
  reg [7:0] p63_res7__822;
  reg [7:0] p63_res7__824;
  reg [7:0] p63_res7__826;
  reg [7:0] p63_res7__828;
  reg [7:0] p64_literal_2043896[256];
  reg [7:0] p64_literal_2043910[256];
  reg [7:0] p64_literal_2043912[256];
  reg [7:0] p64_literal_2043914[256];
  reg [7:0] p64_literal_2043916[256];
  reg [7:0] p64_literal_2043918[256];
  reg [7:0] p64_literal_2043920[256];
  reg [7:0] p64_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p63_encoded <= p62_encoded;
    p63_bit_slice_2043893 <= p62_bit_slice_2043893;
    p63_bit_slice_2044018 <= p62_bit_slice_2044018;
    p63_k3 <= p62_k3;
    p63_k2 <= p62_k2;
    p63_k5 <= p62_k5;
    p63_k4 <= p62_k4;
    p63_k7 <= p62_k7;
    p63_k6 <= p62_k6;
    p63_xor_2055156 <= p62_xor_2055156;
    p63_array_index_2055172 <= p62_array_index_2055172;
    p63_res7__800 <= p62_res7__800;
    p63_array_index_2055285 <= p62_array_index_2055285;
    p63_res7__802 <= p62_res7__802;
    p63_res7__804 <= p62_res7__804;
    p63_array_index_2055314 <= p62_array_index_2055314;
    p63_res7__806 <= p62_res7__806;
    p63_res7__808 <= p62_res7__808;
    p63_array_index_2055342 <= p62_array_index_2055342;
    p63_res7__810 <= p62_res7__810;
    p63_res7__812 <= p62_res7__812;
    p63_array_index_2055368 <= p62_array_index_2055368;
    p63_res7__814 <= p62_res7__814;
    p63_res7__816 <= p63_res7__816_comb;
    p63_array_index_2055520 <= p63_array_index_2055520_comb;
    p63_res7__818 <= p63_res7__818_comb;
    p63_res7__820 <= p63_res7__820_comb;
    p63_array_index_2055542 <= p63_array_index_2055542_comb;
    p63_res7__822 <= p63_res7__822_comb;
    p63_res7__824 <= p63_res7__824_comb;
    p63_res7__826 <= p63_res7__826_comb;
    p63_res7__828 <= p63_res7__828_comb;
    p64_literal_2043896 <= p63_literal_2043896;
    p64_literal_2043910 <= p63_literal_2043910;
    p64_literal_2043912 <= p63_literal_2043912;
    p64_literal_2043914 <= p63_literal_2043914;
    p64_literal_2043916 <= p63_literal_2043916;
    p64_literal_2043918 <= p63_literal_2043918;
    p64_literal_2043920 <= p63_literal_2043920;
    p64_literal_2043923 <= p63_literal_2043923;
  end

  // ===== Pipe stage 64:
  wire [7:0] p64_res7__830_comb;
  wire [127:0] p64_res__25_comb;
  wire [127:0] p64_xor_2055662_comb;
  wire [127:0] p64_addedKey__58_comb;
  wire [7:0] p64_array_index_2055678_comb;
  wire [7:0] p64_array_index_2055679_comb;
  wire [7:0] p64_array_index_2055680_comb;
  wire [7:0] p64_array_index_2055681_comb;
  wire [7:0] p64_array_index_2055682_comb;
  wire [7:0] p64_array_index_2055683_comb;
  wire [7:0] p64_array_index_2055685_comb;
  wire [7:0] p64_array_index_2055687_comb;
  wire [7:0] p64_array_index_2055688_comb;
  wire [7:0] p64_array_index_2055689_comb;
  wire [7:0] p64_array_index_2055690_comb;
  wire [7:0] p64_array_index_2055691_comb;
  wire [7:0] p64_array_index_2055692_comb;
  wire [7:0] p64_array_index_2055694_comb;
  wire [7:0] p64_array_index_2055695_comb;
  wire [7:0] p64_array_index_2055696_comb;
  wire [7:0] p64_array_index_2055697_comb;
  wire [7:0] p64_array_index_2055698_comb;
  wire [7:0] p64_array_index_2055699_comb;
  wire [7:0] p64_array_index_2055700_comb;
  wire [7:0] p64_array_index_2055702_comb;
  wire [7:0] p64_res7__832_comb;
  wire [7:0] p64_array_index_2055711_comb;
  wire [7:0] p64_array_index_2055712_comb;
  wire [7:0] p64_array_index_2055713_comb;
  wire [7:0] p64_array_index_2055714_comb;
  wire [7:0] p64_array_index_2055715_comb;
  wire [7:0] p64_array_index_2055716_comb;
  wire [7:0] p64_res7__834_comb;
  wire [7:0] p64_array_index_2055726_comb;
  wire [7:0] p64_array_index_2055727_comb;
  wire [7:0] p64_array_index_2055728_comb;
  wire [7:0] p64_array_index_2055729_comb;
  wire [7:0] p64_array_index_2055730_comb;
  wire [7:0] p64_res7__836_comb;
  wire [7:0] p64_array_index_2055740_comb;
  wire [7:0] p64_array_index_2055741_comb;
  wire [7:0] p64_array_index_2055742_comb;
  wire [7:0] p64_array_index_2055743_comb;
  wire [7:0] p64_array_index_2055744_comb;
  wire [7:0] p64_res7__838_comb;
  wire [7:0] p64_array_index_2055755_comb;
  wire [7:0] p64_array_index_2055756_comb;
  wire [7:0] p64_array_index_2055757_comb;
  wire [7:0] p64_array_index_2055758_comb;
  wire [7:0] p64_res7__840_comb;
  assign p64_res7__830_comb = p63_literal_2043910[p63_res7__828] ^ p63_literal_2043912[p63_res7__826] ^ p63_literal_2043914[p63_res7__824] ^ p63_literal_2043916[p63_res7__822] ^ p63_literal_2043918[p63_res7__820] ^ p63_literal_2043920[p63_res7__818] ^ p63_res7__816 ^ p63_literal_2043923[p63_res7__814] ^ p63_res7__812 ^ p63_array_index_2055542 ^ p63_array_index_2055520 ^ p63_array_index_2055368 ^ p63_array_index_2055342 ^ p63_array_index_2055314 ^ p63_array_index_2055285 ^ p63_array_index_2055172;
  assign p64_res__25_comb = {p64_res7__830_comb, p63_res7__828, p63_res7__826, p63_res7__824, p63_res7__822, p63_res7__820, p63_res7__818, p63_res7__816, p63_res7__814, p63_res7__812, p63_res7__810, p63_res7__808, p63_res7__806, p63_res7__804, p63_res7__802, p63_res7__800};
  assign p64_xor_2055662_comb = p64_res__25_comb ^ p63_k6;
  assign p64_addedKey__58_comb = p64_xor_2055662_comb ^ 128'h6bce_c0ac_5dd7_7453_d3a7_2473_cd72_011b;
  assign p64_array_index_2055678_comb = p63_literal_2043896[p64_addedKey__58_comb[127:120]];
  assign p64_array_index_2055679_comb = p63_literal_2043896[p64_addedKey__58_comb[119:112]];
  assign p64_array_index_2055680_comb = p63_literal_2043896[p64_addedKey__58_comb[111:104]];
  assign p64_array_index_2055681_comb = p63_literal_2043896[p64_addedKey__58_comb[103:96]];
  assign p64_array_index_2055682_comb = p63_literal_2043896[p64_addedKey__58_comb[95:88]];
  assign p64_array_index_2055683_comb = p63_literal_2043896[p64_addedKey__58_comb[87:80]];
  assign p64_array_index_2055685_comb = p63_literal_2043896[p64_addedKey__58_comb[71:64]];
  assign p64_array_index_2055687_comb = p63_literal_2043896[p64_addedKey__58_comb[55:48]];
  assign p64_array_index_2055688_comb = p63_literal_2043896[p64_addedKey__58_comb[47:40]];
  assign p64_array_index_2055689_comb = p63_literal_2043896[p64_addedKey__58_comb[39:32]];
  assign p64_array_index_2055690_comb = p63_literal_2043896[p64_addedKey__58_comb[31:24]];
  assign p64_array_index_2055691_comb = p63_literal_2043896[p64_addedKey__58_comb[23:16]];
  assign p64_array_index_2055692_comb = p63_literal_2043896[p64_addedKey__58_comb[15:8]];
  assign p64_array_index_2055694_comb = p63_literal_2043910[p64_array_index_2055678_comb];
  assign p64_array_index_2055695_comb = p63_literal_2043912[p64_array_index_2055679_comb];
  assign p64_array_index_2055696_comb = p63_literal_2043914[p64_array_index_2055680_comb];
  assign p64_array_index_2055697_comb = p63_literal_2043916[p64_array_index_2055681_comb];
  assign p64_array_index_2055698_comb = p63_literal_2043918[p64_array_index_2055682_comb];
  assign p64_array_index_2055699_comb = p63_literal_2043920[p64_array_index_2055683_comb];
  assign p64_array_index_2055700_comb = p63_literal_2043896[p64_addedKey__58_comb[79:72]];
  assign p64_array_index_2055702_comb = p63_literal_2043896[p64_addedKey__58_comb[63:56]];
  assign p64_res7__832_comb = p64_array_index_2055694_comb ^ p64_array_index_2055695_comb ^ p64_array_index_2055696_comb ^ p64_array_index_2055697_comb ^ p64_array_index_2055698_comb ^ p64_array_index_2055699_comb ^ p64_array_index_2055700_comb ^ p63_literal_2043923[p64_array_index_2055685_comb] ^ p64_array_index_2055702_comb ^ p63_literal_2043920[p64_array_index_2055687_comb] ^ p63_literal_2043918[p64_array_index_2055688_comb] ^ p63_literal_2043916[p64_array_index_2055689_comb] ^ p63_literal_2043914[p64_array_index_2055690_comb] ^ p63_literal_2043912[p64_array_index_2055691_comb] ^ p63_literal_2043910[p64_array_index_2055692_comb] ^ p63_literal_2043896[p64_addedKey__58_comb[7:0]];
  assign p64_array_index_2055711_comb = p63_literal_2043910[p64_res7__832_comb];
  assign p64_array_index_2055712_comb = p63_literal_2043912[p64_array_index_2055678_comb];
  assign p64_array_index_2055713_comb = p63_literal_2043914[p64_array_index_2055679_comb];
  assign p64_array_index_2055714_comb = p63_literal_2043916[p64_array_index_2055680_comb];
  assign p64_array_index_2055715_comb = p63_literal_2043918[p64_array_index_2055681_comb];
  assign p64_array_index_2055716_comb = p63_literal_2043920[p64_array_index_2055682_comb];
  assign p64_res7__834_comb = p64_array_index_2055711_comb ^ p64_array_index_2055712_comb ^ p64_array_index_2055713_comb ^ p64_array_index_2055714_comb ^ p64_array_index_2055715_comb ^ p64_array_index_2055716_comb ^ p64_array_index_2055683_comb ^ p63_literal_2043923[p64_array_index_2055700_comb] ^ p64_array_index_2055685_comb ^ p63_literal_2043920[p64_array_index_2055702_comb] ^ p63_literal_2043918[p64_array_index_2055687_comb] ^ p63_literal_2043916[p64_array_index_2055688_comb] ^ p63_literal_2043914[p64_array_index_2055689_comb] ^ p63_literal_2043912[p64_array_index_2055690_comb] ^ p63_literal_2043910[p64_array_index_2055691_comb] ^ p64_array_index_2055692_comb;
  assign p64_array_index_2055726_comb = p63_literal_2043912[p64_res7__832_comb];
  assign p64_array_index_2055727_comb = p63_literal_2043914[p64_array_index_2055678_comb];
  assign p64_array_index_2055728_comb = p63_literal_2043916[p64_array_index_2055679_comb];
  assign p64_array_index_2055729_comb = p63_literal_2043918[p64_array_index_2055680_comb];
  assign p64_array_index_2055730_comb = p63_literal_2043920[p64_array_index_2055681_comb];
  assign p64_res7__836_comb = p63_literal_2043910[p64_res7__834_comb] ^ p64_array_index_2055726_comb ^ p64_array_index_2055727_comb ^ p64_array_index_2055728_comb ^ p64_array_index_2055729_comb ^ p64_array_index_2055730_comb ^ p64_array_index_2055682_comb ^ p63_literal_2043923[p64_array_index_2055683_comb] ^ p64_array_index_2055700_comb ^ p63_literal_2043920[p64_array_index_2055685_comb] ^ p63_literal_2043918[p64_array_index_2055702_comb] ^ p63_literal_2043916[p64_array_index_2055687_comb] ^ p63_literal_2043914[p64_array_index_2055688_comb] ^ p63_literal_2043912[p64_array_index_2055689_comb] ^ p63_literal_2043910[p64_array_index_2055690_comb] ^ p64_array_index_2055691_comb;
  assign p64_array_index_2055740_comb = p63_literal_2043912[p64_res7__834_comb];
  assign p64_array_index_2055741_comb = p63_literal_2043914[p64_res7__832_comb];
  assign p64_array_index_2055742_comb = p63_literal_2043916[p64_array_index_2055678_comb];
  assign p64_array_index_2055743_comb = p63_literal_2043918[p64_array_index_2055679_comb];
  assign p64_array_index_2055744_comb = p63_literal_2043920[p64_array_index_2055680_comb];
  assign p64_res7__838_comb = p63_literal_2043910[p64_res7__836_comb] ^ p64_array_index_2055740_comb ^ p64_array_index_2055741_comb ^ p64_array_index_2055742_comb ^ p64_array_index_2055743_comb ^ p64_array_index_2055744_comb ^ p64_array_index_2055681_comb ^ p63_literal_2043923[p64_array_index_2055682_comb] ^ p64_array_index_2055683_comb ^ p63_literal_2043920[p64_array_index_2055700_comb] ^ p63_literal_2043918[p64_array_index_2055685_comb] ^ p63_literal_2043916[p64_array_index_2055702_comb] ^ p63_literal_2043914[p64_array_index_2055687_comb] ^ p63_literal_2043912[p64_array_index_2055688_comb] ^ p63_literal_2043910[p64_array_index_2055689_comb] ^ p64_array_index_2055690_comb;
  assign p64_array_index_2055755_comb = p63_literal_2043914[p64_res7__834_comb];
  assign p64_array_index_2055756_comb = p63_literal_2043916[p64_res7__832_comb];
  assign p64_array_index_2055757_comb = p63_literal_2043918[p64_array_index_2055678_comb];
  assign p64_array_index_2055758_comb = p63_literal_2043920[p64_array_index_2055679_comb];
  assign p64_res7__840_comb = p63_literal_2043910[p64_res7__838_comb] ^ p63_literal_2043912[p64_res7__836_comb] ^ p64_array_index_2055755_comb ^ p64_array_index_2055756_comb ^ p64_array_index_2055757_comb ^ p64_array_index_2055758_comb ^ p64_array_index_2055680_comb ^ p63_literal_2043923[p64_array_index_2055681_comb] ^ p64_array_index_2055682_comb ^ p64_array_index_2055699_comb ^ p63_literal_2043918[p64_array_index_2055700_comb] ^ p63_literal_2043916[p64_array_index_2055685_comb] ^ p63_literal_2043914[p64_array_index_2055702_comb] ^ p63_literal_2043912[p64_array_index_2055687_comb] ^ p63_literal_2043910[p64_array_index_2055688_comb] ^ p64_array_index_2055689_comb;

  // Registers for pipe stage 64:
  reg [127:0] p64_encoded;
  reg [127:0] p64_bit_slice_2043893;
  reg [127:0] p64_bit_slice_2044018;
  reg [127:0] p64_k3;
  reg [127:0] p64_k2;
  reg [127:0] p64_k5;
  reg [127:0] p64_k4;
  reg [127:0] p64_k7;
  reg [127:0] p64_k6;
  reg [127:0] p64_xor_2055156;
  reg [127:0] p64_xor_2055662;
  reg [7:0] p64_array_index_2055678;
  reg [7:0] p64_array_index_2055679;
  reg [7:0] p64_array_index_2055680;
  reg [7:0] p64_array_index_2055681;
  reg [7:0] p64_array_index_2055682;
  reg [7:0] p64_array_index_2055683;
  reg [7:0] p64_array_index_2055685;
  reg [7:0] p64_array_index_2055687;
  reg [7:0] p64_array_index_2055688;
  reg [7:0] p64_array_index_2055694;
  reg [7:0] p64_array_index_2055695;
  reg [7:0] p64_array_index_2055696;
  reg [7:0] p64_array_index_2055697;
  reg [7:0] p64_array_index_2055698;
  reg [7:0] p64_array_index_2055700;
  reg [7:0] p64_array_index_2055702;
  reg [7:0] p64_res7__832;
  reg [7:0] p64_array_index_2055711;
  reg [7:0] p64_array_index_2055712;
  reg [7:0] p64_array_index_2055713;
  reg [7:0] p64_array_index_2055714;
  reg [7:0] p64_array_index_2055715;
  reg [7:0] p64_array_index_2055716;
  reg [7:0] p64_res7__834;
  reg [7:0] p64_array_index_2055726;
  reg [7:0] p64_array_index_2055727;
  reg [7:0] p64_array_index_2055728;
  reg [7:0] p64_array_index_2055729;
  reg [7:0] p64_array_index_2055730;
  reg [7:0] p64_res7__836;
  reg [7:0] p64_array_index_2055740;
  reg [7:0] p64_array_index_2055741;
  reg [7:0] p64_array_index_2055742;
  reg [7:0] p64_array_index_2055743;
  reg [7:0] p64_array_index_2055744;
  reg [7:0] p64_res7__838;
  reg [7:0] p64_array_index_2055755;
  reg [7:0] p64_array_index_2055756;
  reg [7:0] p64_array_index_2055757;
  reg [7:0] p64_array_index_2055758;
  reg [7:0] p64_res7__840;
  reg [7:0] p65_literal_2043896[256];
  reg [7:0] p65_literal_2043910[256];
  reg [7:0] p65_literal_2043912[256];
  reg [7:0] p65_literal_2043914[256];
  reg [7:0] p65_literal_2043916[256];
  reg [7:0] p65_literal_2043918[256];
  reg [7:0] p65_literal_2043920[256];
  reg [7:0] p65_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p64_encoded <= p63_encoded;
    p64_bit_slice_2043893 <= p63_bit_slice_2043893;
    p64_bit_slice_2044018 <= p63_bit_slice_2044018;
    p64_k3 <= p63_k3;
    p64_k2 <= p63_k2;
    p64_k5 <= p63_k5;
    p64_k4 <= p63_k4;
    p64_k7 <= p63_k7;
    p64_k6 <= p63_k6;
    p64_xor_2055156 <= p63_xor_2055156;
    p64_xor_2055662 <= p64_xor_2055662_comb;
    p64_array_index_2055678 <= p64_array_index_2055678_comb;
    p64_array_index_2055679 <= p64_array_index_2055679_comb;
    p64_array_index_2055680 <= p64_array_index_2055680_comb;
    p64_array_index_2055681 <= p64_array_index_2055681_comb;
    p64_array_index_2055682 <= p64_array_index_2055682_comb;
    p64_array_index_2055683 <= p64_array_index_2055683_comb;
    p64_array_index_2055685 <= p64_array_index_2055685_comb;
    p64_array_index_2055687 <= p64_array_index_2055687_comb;
    p64_array_index_2055688 <= p64_array_index_2055688_comb;
    p64_array_index_2055694 <= p64_array_index_2055694_comb;
    p64_array_index_2055695 <= p64_array_index_2055695_comb;
    p64_array_index_2055696 <= p64_array_index_2055696_comb;
    p64_array_index_2055697 <= p64_array_index_2055697_comb;
    p64_array_index_2055698 <= p64_array_index_2055698_comb;
    p64_array_index_2055700 <= p64_array_index_2055700_comb;
    p64_array_index_2055702 <= p64_array_index_2055702_comb;
    p64_res7__832 <= p64_res7__832_comb;
    p64_array_index_2055711 <= p64_array_index_2055711_comb;
    p64_array_index_2055712 <= p64_array_index_2055712_comb;
    p64_array_index_2055713 <= p64_array_index_2055713_comb;
    p64_array_index_2055714 <= p64_array_index_2055714_comb;
    p64_array_index_2055715 <= p64_array_index_2055715_comb;
    p64_array_index_2055716 <= p64_array_index_2055716_comb;
    p64_res7__834 <= p64_res7__834_comb;
    p64_array_index_2055726 <= p64_array_index_2055726_comb;
    p64_array_index_2055727 <= p64_array_index_2055727_comb;
    p64_array_index_2055728 <= p64_array_index_2055728_comb;
    p64_array_index_2055729 <= p64_array_index_2055729_comb;
    p64_array_index_2055730 <= p64_array_index_2055730_comb;
    p64_res7__836 <= p64_res7__836_comb;
    p64_array_index_2055740 <= p64_array_index_2055740_comb;
    p64_array_index_2055741 <= p64_array_index_2055741_comb;
    p64_array_index_2055742 <= p64_array_index_2055742_comb;
    p64_array_index_2055743 <= p64_array_index_2055743_comb;
    p64_array_index_2055744 <= p64_array_index_2055744_comb;
    p64_res7__838 <= p64_res7__838_comb;
    p64_array_index_2055755 <= p64_array_index_2055755_comb;
    p64_array_index_2055756 <= p64_array_index_2055756_comb;
    p64_array_index_2055757 <= p64_array_index_2055757_comb;
    p64_array_index_2055758 <= p64_array_index_2055758_comb;
    p64_res7__840 <= p64_res7__840_comb;
    p65_literal_2043896 <= p64_literal_2043896;
    p65_literal_2043910 <= p64_literal_2043910;
    p65_literal_2043912 <= p64_literal_2043912;
    p65_literal_2043914 <= p64_literal_2043914;
    p65_literal_2043916 <= p64_literal_2043916;
    p65_literal_2043918 <= p64_literal_2043918;
    p65_literal_2043920 <= p64_literal_2043920;
    p65_literal_2043923 <= p64_literal_2043923;
  end

  // ===== Pipe stage 65:
  wire [7:0] p65_array_index_2055888_comb;
  wire [7:0] p65_array_index_2055889_comb;
  wire [7:0] p65_array_index_2055890_comb;
  wire [7:0] p65_array_index_2055891_comb;
  wire [7:0] p65_res7__842_comb;
  wire [7:0] p65_array_index_2055902_comb;
  wire [7:0] p65_array_index_2055903_comb;
  wire [7:0] p65_array_index_2055904_comb;
  wire [7:0] p65_res7__844_comb;
  wire [7:0] p65_array_index_2055914_comb;
  wire [7:0] p65_array_index_2055915_comb;
  wire [7:0] p65_array_index_2055916_comb;
  wire [7:0] p65_res7__846_comb;
  wire [7:0] p65_array_index_2055927_comb;
  wire [7:0] p65_array_index_2055928_comb;
  wire [7:0] p65_res7__848_comb;
  wire [7:0] p65_array_index_2055938_comb;
  wire [7:0] p65_array_index_2055939_comb;
  wire [7:0] p65_res7__850_comb;
  wire [7:0] p65_array_index_2055950_comb;
  wire [7:0] p65_res7__852_comb;
  wire [7:0] p65_array_index_2055960_comb;
  wire [7:0] p65_res7__854_comb;
  assign p65_array_index_2055888_comb = p64_literal_2043914[p64_res7__836];
  assign p65_array_index_2055889_comb = p64_literal_2043916[p64_res7__834];
  assign p65_array_index_2055890_comb = p64_literal_2043918[p64_res7__832];
  assign p65_array_index_2055891_comb = p64_literal_2043920[p64_array_index_2055678];
  assign p65_res7__842_comb = p64_literal_2043910[p64_res7__840] ^ p64_literal_2043912[p64_res7__838] ^ p65_array_index_2055888_comb ^ p65_array_index_2055889_comb ^ p65_array_index_2055890_comb ^ p65_array_index_2055891_comb ^ p64_array_index_2055679 ^ p64_literal_2043923[p64_array_index_2055680] ^ p64_array_index_2055681 ^ p64_array_index_2055716 ^ p64_literal_2043918[p64_array_index_2055683] ^ p64_literal_2043916[p64_array_index_2055700] ^ p64_literal_2043914[p64_array_index_2055685] ^ p64_literal_2043912[p64_array_index_2055702] ^ p64_literal_2043910[p64_array_index_2055687] ^ p64_array_index_2055688;
  assign p65_array_index_2055902_comb = p64_literal_2043916[p64_res7__836];
  assign p65_array_index_2055903_comb = p64_literal_2043918[p64_res7__834];
  assign p65_array_index_2055904_comb = p64_literal_2043920[p64_res7__832];
  assign p65_res7__844_comb = p64_literal_2043910[p65_res7__842_comb] ^ p64_literal_2043912[p64_res7__840] ^ p64_literal_2043914[p64_res7__838] ^ p65_array_index_2055902_comb ^ p65_array_index_2055903_comb ^ p65_array_index_2055904_comb ^ p64_array_index_2055678 ^ p64_literal_2043923[p64_array_index_2055679] ^ p64_array_index_2055680 ^ p64_array_index_2055730 ^ p64_array_index_2055698 ^ p64_literal_2043916[p64_array_index_2055683] ^ p64_literal_2043914[p64_array_index_2055700] ^ p64_literal_2043912[p64_array_index_2055685] ^ p64_literal_2043910[p64_array_index_2055702] ^ p64_array_index_2055687;
  assign p65_array_index_2055914_comb = p64_literal_2043916[p64_res7__838];
  assign p65_array_index_2055915_comb = p64_literal_2043918[p64_res7__836];
  assign p65_array_index_2055916_comb = p64_literal_2043920[p64_res7__834];
  assign p65_res7__846_comb = p64_literal_2043910[p65_res7__844_comb] ^ p64_literal_2043912[p65_res7__842_comb] ^ p64_literal_2043914[p64_res7__840] ^ p65_array_index_2055914_comb ^ p65_array_index_2055915_comb ^ p65_array_index_2055916_comb ^ p64_res7__832 ^ p64_literal_2043923[p64_array_index_2055678] ^ p64_array_index_2055679 ^ p64_array_index_2055744 ^ p64_array_index_2055715 ^ p64_literal_2043916[p64_array_index_2055682] ^ p64_literal_2043914[p64_array_index_2055683] ^ p64_literal_2043912[p64_array_index_2055700] ^ p64_literal_2043910[p64_array_index_2055685] ^ p64_array_index_2055702;
  assign p65_array_index_2055927_comb = p64_literal_2043918[p64_res7__838];
  assign p65_array_index_2055928_comb = p64_literal_2043920[p64_res7__836];
  assign p65_res7__848_comb = p64_literal_2043910[p65_res7__846_comb] ^ p64_literal_2043912[p65_res7__844_comb] ^ p64_literal_2043914[p65_res7__842_comb] ^ p64_literal_2043916[p64_res7__840] ^ p65_array_index_2055927_comb ^ p65_array_index_2055928_comb ^ p64_res7__834 ^ p64_literal_2043923[p64_res7__832] ^ p64_array_index_2055678 ^ p64_array_index_2055758 ^ p64_array_index_2055729 ^ p64_array_index_2055697 ^ p64_literal_2043914[p64_array_index_2055682] ^ p64_literal_2043912[p64_array_index_2055683] ^ p64_literal_2043910[p64_array_index_2055700] ^ p64_array_index_2055685;
  assign p65_array_index_2055938_comb = p64_literal_2043918[p64_res7__840];
  assign p65_array_index_2055939_comb = p64_literal_2043920[p64_res7__838];
  assign p65_res7__850_comb = p64_literal_2043910[p65_res7__848_comb] ^ p64_literal_2043912[p65_res7__846_comb] ^ p64_literal_2043914[p65_res7__844_comb] ^ p64_literal_2043916[p65_res7__842_comb] ^ p65_array_index_2055938_comb ^ p65_array_index_2055939_comb ^ p64_res7__836 ^ p64_literal_2043923[p64_res7__834] ^ p64_res7__832 ^ p65_array_index_2055891_comb ^ p64_array_index_2055743 ^ p64_array_index_2055714 ^ p64_literal_2043914[p64_array_index_2055681] ^ p64_literal_2043912[p64_array_index_2055682] ^ p64_literal_2043910[p64_array_index_2055683] ^ p64_array_index_2055700;
  assign p65_array_index_2055950_comb = p64_literal_2043920[p64_res7__840];
  assign p65_res7__852_comb = p64_literal_2043910[p65_res7__850_comb] ^ p64_literal_2043912[p65_res7__848_comb] ^ p64_literal_2043914[p65_res7__846_comb] ^ p64_literal_2043916[p65_res7__844_comb] ^ p64_literal_2043918[p65_res7__842_comb] ^ p65_array_index_2055950_comb ^ p64_res7__838 ^ p64_literal_2043923[p64_res7__836] ^ p64_res7__834 ^ p65_array_index_2055904_comb ^ p64_array_index_2055757 ^ p64_array_index_2055728 ^ p64_array_index_2055696 ^ p64_literal_2043912[p64_array_index_2055681] ^ p64_literal_2043910[p64_array_index_2055682] ^ p64_array_index_2055683;
  assign p65_array_index_2055960_comb = p64_literal_2043920[p65_res7__842_comb];
  assign p65_res7__854_comb = p64_literal_2043910[p65_res7__852_comb] ^ p64_literal_2043912[p65_res7__850_comb] ^ p64_literal_2043914[p65_res7__848_comb] ^ p64_literal_2043916[p65_res7__846_comb] ^ p64_literal_2043918[p65_res7__844_comb] ^ p65_array_index_2055960_comb ^ p64_res7__840 ^ p64_literal_2043923[p64_res7__838] ^ p64_res7__836 ^ p65_array_index_2055916_comb ^ p65_array_index_2055890_comb ^ p64_array_index_2055742 ^ p64_array_index_2055713 ^ p64_literal_2043912[p64_array_index_2055680] ^ p64_literal_2043910[p64_array_index_2055681] ^ p64_array_index_2055682;

  // Registers for pipe stage 65:
  reg [127:0] p65_encoded;
  reg [127:0] p65_bit_slice_2043893;
  reg [127:0] p65_bit_slice_2044018;
  reg [127:0] p65_k3;
  reg [127:0] p65_k2;
  reg [127:0] p65_k5;
  reg [127:0] p65_k4;
  reg [127:0] p65_k7;
  reg [127:0] p65_k6;
  reg [127:0] p65_xor_2055156;
  reg [127:0] p65_xor_2055662;
  reg [7:0] p65_array_index_2055678;
  reg [7:0] p65_array_index_2055679;
  reg [7:0] p65_array_index_2055680;
  reg [7:0] p65_array_index_2055681;
  reg [7:0] p65_array_index_2055694;
  reg [7:0] p65_array_index_2055695;
  reg [7:0] p65_res7__832;
  reg [7:0] p65_array_index_2055711;
  reg [7:0] p65_array_index_2055712;
  reg [7:0] p65_res7__834;
  reg [7:0] p65_array_index_2055726;
  reg [7:0] p65_array_index_2055727;
  reg [7:0] p65_res7__836;
  reg [7:0] p65_array_index_2055740;
  reg [7:0] p65_array_index_2055741;
  reg [7:0] p65_res7__838;
  reg [7:0] p65_array_index_2055755;
  reg [7:0] p65_array_index_2055756;
  reg [7:0] p65_res7__840;
  reg [7:0] p65_array_index_2055888;
  reg [7:0] p65_array_index_2055889;
  reg [7:0] p65_res7__842;
  reg [7:0] p65_array_index_2055902;
  reg [7:0] p65_array_index_2055903;
  reg [7:0] p65_res7__844;
  reg [7:0] p65_array_index_2055914;
  reg [7:0] p65_array_index_2055915;
  reg [7:0] p65_res7__846;
  reg [7:0] p65_array_index_2055927;
  reg [7:0] p65_array_index_2055928;
  reg [7:0] p65_res7__848;
  reg [7:0] p65_array_index_2055938;
  reg [7:0] p65_array_index_2055939;
  reg [7:0] p65_res7__850;
  reg [7:0] p65_array_index_2055950;
  reg [7:0] p65_res7__852;
  reg [7:0] p65_array_index_2055960;
  reg [7:0] p65_res7__854;
  reg [7:0] p66_literal_2043896[256];
  reg [7:0] p66_literal_2043910[256];
  reg [7:0] p66_literal_2043912[256];
  reg [7:0] p66_literal_2043914[256];
  reg [7:0] p66_literal_2043916[256];
  reg [7:0] p66_literal_2043918[256];
  reg [7:0] p66_literal_2043920[256];
  reg [7:0] p66_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p65_encoded <= p64_encoded;
    p65_bit_slice_2043893 <= p64_bit_slice_2043893;
    p65_bit_slice_2044018 <= p64_bit_slice_2044018;
    p65_k3 <= p64_k3;
    p65_k2 <= p64_k2;
    p65_k5 <= p64_k5;
    p65_k4 <= p64_k4;
    p65_k7 <= p64_k7;
    p65_k6 <= p64_k6;
    p65_xor_2055156 <= p64_xor_2055156;
    p65_xor_2055662 <= p64_xor_2055662;
    p65_array_index_2055678 <= p64_array_index_2055678;
    p65_array_index_2055679 <= p64_array_index_2055679;
    p65_array_index_2055680 <= p64_array_index_2055680;
    p65_array_index_2055681 <= p64_array_index_2055681;
    p65_array_index_2055694 <= p64_array_index_2055694;
    p65_array_index_2055695 <= p64_array_index_2055695;
    p65_res7__832 <= p64_res7__832;
    p65_array_index_2055711 <= p64_array_index_2055711;
    p65_array_index_2055712 <= p64_array_index_2055712;
    p65_res7__834 <= p64_res7__834;
    p65_array_index_2055726 <= p64_array_index_2055726;
    p65_array_index_2055727 <= p64_array_index_2055727;
    p65_res7__836 <= p64_res7__836;
    p65_array_index_2055740 <= p64_array_index_2055740;
    p65_array_index_2055741 <= p64_array_index_2055741;
    p65_res7__838 <= p64_res7__838;
    p65_array_index_2055755 <= p64_array_index_2055755;
    p65_array_index_2055756 <= p64_array_index_2055756;
    p65_res7__840 <= p64_res7__840;
    p65_array_index_2055888 <= p65_array_index_2055888_comb;
    p65_array_index_2055889 <= p65_array_index_2055889_comb;
    p65_res7__842 <= p65_res7__842_comb;
    p65_array_index_2055902 <= p65_array_index_2055902_comb;
    p65_array_index_2055903 <= p65_array_index_2055903_comb;
    p65_res7__844 <= p65_res7__844_comb;
    p65_array_index_2055914 <= p65_array_index_2055914_comb;
    p65_array_index_2055915 <= p65_array_index_2055915_comb;
    p65_res7__846 <= p65_res7__846_comb;
    p65_array_index_2055927 <= p65_array_index_2055927_comb;
    p65_array_index_2055928 <= p65_array_index_2055928_comb;
    p65_res7__848 <= p65_res7__848_comb;
    p65_array_index_2055938 <= p65_array_index_2055938_comb;
    p65_array_index_2055939 <= p65_array_index_2055939_comb;
    p65_res7__850 <= p65_res7__850_comb;
    p65_array_index_2055950 <= p65_array_index_2055950_comb;
    p65_res7__852 <= p65_res7__852_comb;
    p65_array_index_2055960 <= p65_array_index_2055960_comb;
    p65_res7__854 <= p65_res7__854_comb;
    p66_literal_2043896 <= p65_literal_2043896;
    p66_literal_2043910 <= p65_literal_2043910;
    p66_literal_2043912 <= p65_literal_2043912;
    p66_literal_2043914 <= p65_literal_2043914;
    p66_literal_2043916 <= p65_literal_2043916;
    p66_literal_2043918 <= p65_literal_2043918;
    p66_literal_2043920 <= p65_literal_2043920;
    p66_literal_2043923 <= p65_literal_2043923;
  end

  // ===== Pipe stage 66:
  wire [7:0] p66_res7__856_comb;
  wire [7:0] p66_res7__858_comb;
  wire [7:0] p66_res7__860_comb;
  wire [7:0] p66_res7__862_comb;
  wire [127:0] p66_res__26_comb;
  wire [127:0] p66_xor_2056114_comb;
  wire [127:0] p66_addedKey__59_comb;
  wire [7:0] p66_array_index_2056130_comb;
  wire [7:0] p66_array_index_2056131_comb;
  wire [7:0] p66_array_index_2056132_comb;
  wire [7:0] p66_array_index_2056133_comb;
  wire [7:0] p66_array_index_2056134_comb;
  wire [7:0] p66_array_index_2056135_comb;
  wire [7:0] p66_array_index_2056137_comb;
  wire [7:0] p66_array_index_2056139_comb;
  wire [7:0] p66_array_index_2056140_comb;
  wire [7:0] p66_array_index_2056141_comb;
  wire [7:0] p66_array_index_2056142_comb;
  wire [7:0] p66_array_index_2056143_comb;
  wire [7:0] p66_array_index_2056144_comb;
  wire [7:0] p66_array_index_2056146_comb;
  wire [7:0] p66_array_index_2056147_comb;
  wire [7:0] p66_array_index_2056148_comb;
  wire [7:0] p66_array_index_2056149_comb;
  wire [7:0] p66_array_index_2056150_comb;
  wire [7:0] p66_array_index_2056151_comb;
  wire [7:0] p66_array_index_2056152_comb;
  wire [7:0] p66_array_index_2056154_comb;
  wire [7:0] p66_res7__864_comb;
  wire [7:0] p66_array_index_2056163_comb;
  wire [7:0] p66_array_index_2056164_comb;
  wire [7:0] p66_array_index_2056165_comb;
  wire [7:0] p66_array_index_2056166_comb;
  wire [7:0] p66_array_index_2056167_comb;
  wire [7:0] p66_array_index_2056168_comb;
  wire [7:0] p66_res7__866_comb;
  assign p66_res7__856_comb = p65_literal_2043910[p65_res7__854] ^ p65_literal_2043912[p65_res7__852] ^ p65_literal_2043914[p65_res7__850] ^ p65_literal_2043916[p65_res7__848] ^ p65_literal_2043918[p65_res7__846] ^ p65_literal_2043920[p65_res7__844] ^ p65_res7__842 ^ p65_literal_2043923[p65_res7__840] ^ p65_res7__838 ^ p65_array_index_2055928 ^ p65_array_index_2055903 ^ p65_array_index_2055756 ^ p65_array_index_2055727 ^ p65_array_index_2055695 ^ p65_literal_2043910[p65_array_index_2055680] ^ p65_array_index_2055681;
  assign p66_res7__858_comb = p65_literal_2043910[p66_res7__856_comb] ^ p65_literal_2043912[p65_res7__854] ^ p65_literal_2043914[p65_res7__852] ^ p65_literal_2043916[p65_res7__850] ^ p65_literal_2043918[p65_res7__848] ^ p65_literal_2043920[p65_res7__846] ^ p65_res7__844 ^ p65_literal_2043923[p65_res7__842] ^ p65_res7__840 ^ p65_array_index_2055939 ^ p65_array_index_2055915 ^ p65_array_index_2055889 ^ p65_array_index_2055741 ^ p65_array_index_2055712 ^ p65_literal_2043910[p65_array_index_2055679] ^ p65_array_index_2055680;
  assign p66_res7__860_comb = p65_literal_2043910[p66_res7__858_comb] ^ p65_literal_2043912[p66_res7__856_comb] ^ p65_literal_2043914[p65_res7__854] ^ p65_literal_2043916[p65_res7__852] ^ p65_literal_2043918[p65_res7__850] ^ p65_literal_2043920[p65_res7__848] ^ p65_res7__846 ^ p65_literal_2043923[p65_res7__844] ^ p65_res7__842 ^ p65_array_index_2055950 ^ p65_array_index_2055927 ^ p65_array_index_2055902 ^ p65_array_index_2055755 ^ p65_array_index_2055726 ^ p65_array_index_2055694 ^ p65_array_index_2055679;
  assign p66_res7__862_comb = p65_literal_2043910[p66_res7__860_comb] ^ p65_literal_2043912[p66_res7__858_comb] ^ p65_literal_2043914[p66_res7__856_comb] ^ p65_literal_2043916[p65_res7__854] ^ p65_literal_2043918[p65_res7__852] ^ p65_literal_2043920[p65_res7__850] ^ p65_res7__848 ^ p65_literal_2043923[p65_res7__846] ^ p65_res7__844 ^ p65_array_index_2055960 ^ p65_array_index_2055938 ^ p65_array_index_2055914 ^ p65_array_index_2055888 ^ p65_array_index_2055740 ^ p65_array_index_2055711 ^ p65_array_index_2055678;
  assign p66_res__26_comb = {p66_res7__862_comb, p66_res7__860_comb, p66_res7__858_comb, p66_res7__856_comb, p65_res7__854, p65_res7__852, p65_res7__850, p65_res7__848, p65_res7__846, p65_res7__844, p65_res7__842, p65_res7__840, p65_res7__838, p65_res7__836, p65_res7__834, p65_res7__832};
  assign p66_xor_2056114_comb = p66_res__26_comb ^ p65_xor_2055156;
  assign p66_addedKey__59_comb = p66_xor_2056114_comb ^ 128'ha226_4131_9aec_d1fd_8352_9103_9b68_6b1c;
  assign p66_array_index_2056130_comb = p65_literal_2043896[p66_addedKey__59_comb[127:120]];
  assign p66_array_index_2056131_comb = p65_literal_2043896[p66_addedKey__59_comb[119:112]];
  assign p66_array_index_2056132_comb = p65_literal_2043896[p66_addedKey__59_comb[111:104]];
  assign p66_array_index_2056133_comb = p65_literal_2043896[p66_addedKey__59_comb[103:96]];
  assign p66_array_index_2056134_comb = p65_literal_2043896[p66_addedKey__59_comb[95:88]];
  assign p66_array_index_2056135_comb = p65_literal_2043896[p66_addedKey__59_comb[87:80]];
  assign p66_array_index_2056137_comb = p65_literal_2043896[p66_addedKey__59_comb[71:64]];
  assign p66_array_index_2056139_comb = p65_literal_2043896[p66_addedKey__59_comb[55:48]];
  assign p66_array_index_2056140_comb = p65_literal_2043896[p66_addedKey__59_comb[47:40]];
  assign p66_array_index_2056141_comb = p65_literal_2043896[p66_addedKey__59_comb[39:32]];
  assign p66_array_index_2056142_comb = p65_literal_2043896[p66_addedKey__59_comb[31:24]];
  assign p66_array_index_2056143_comb = p65_literal_2043896[p66_addedKey__59_comb[23:16]];
  assign p66_array_index_2056144_comb = p65_literal_2043896[p66_addedKey__59_comb[15:8]];
  assign p66_array_index_2056146_comb = p65_literal_2043910[p66_array_index_2056130_comb];
  assign p66_array_index_2056147_comb = p65_literal_2043912[p66_array_index_2056131_comb];
  assign p66_array_index_2056148_comb = p65_literal_2043914[p66_array_index_2056132_comb];
  assign p66_array_index_2056149_comb = p65_literal_2043916[p66_array_index_2056133_comb];
  assign p66_array_index_2056150_comb = p65_literal_2043918[p66_array_index_2056134_comb];
  assign p66_array_index_2056151_comb = p65_literal_2043920[p66_array_index_2056135_comb];
  assign p66_array_index_2056152_comb = p65_literal_2043896[p66_addedKey__59_comb[79:72]];
  assign p66_array_index_2056154_comb = p65_literal_2043896[p66_addedKey__59_comb[63:56]];
  assign p66_res7__864_comb = p66_array_index_2056146_comb ^ p66_array_index_2056147_comb ^ p66_array_index_2056148_comb ^ p66_array_index_2056149_comb ^ p66_array_index_2056150_comb ^ p66_array_index_2056151_comb ^ p66_array_index_2056152_comb ^ p65_literal_2043923[p66_array_index_2056137_comb] ^ p66_array_index_2056154_comb ^ p65_literal_2043920[p66_array_index_2056139_comb] ^ p65_literal_2043918[p66_array_index_2056140_comb] ^ p65_literal_2043916[p66_array_index_2056141_comb] ^ p65_literal_2043914[p66_array_index_2056142_comb] ^ p65_literal_2043912[p66_array_index_2056143_comb] ^ p65_literal_2043910[p66_array_index_2056144_comb] ^ p65_literal_2043896[p66_addedKey__59_comb[7:0]];
  assign p66_array_index_2056163_comb = p65_literal_2043910[p66_res7__864_comb];
  assign p66_array_index_2056164_comb = p65_literal_2043912[p66_array_index_2056130_comb];
  assign p66_array_index_2056165_comb = p65_literal_2043914[p66_array_index_2056131_comb];
  assign p66_array_index_2056166_comb = p65_literal_2043916[p66_array_index_2056132_comb];
  assign p66_array_index_2056167_comb = p65_literal_2043918[p66_array_index_2056133_comb];
  assign p66_array_index_2056168_comb = p65_literal_2043920[p66_array_index_2056134_comb];
  assign p66_res7__866_comb = p66_array_index_2056163_comb ^ p66_array_index_2056164_comb ^ p66_array_index_2056165_comb ^ p66_array_index_2056166_comb ^ p66_array_index_2056167_comb ^ p66_array_index_2056168_comb ^ p66_array_index_2056135_comb ^ p65_literal_2043923[p66_array_index_2056152_comb] ^ p66_array_index_2056137_comb ^ p65_literal_2043920[p66_array_index_2056154_comb] ^ p65_literal_2043918[p66_array_index_2056139_comb] ^ p65_literal_2043916[p66_array_index_2056140_comb] ^ p65_literal_2043914[p66_array_index_2056141_comb] ^ p65_literal_2043912[p66_array_index_2056142_comb] ^ p65_literal_2043910[p66_array_index_2056143_comb] ^ p66_array_index_2056144_comb;

  // Registers for pipe stage 66:
  reg [127:0] p66_encoded;
  reg [127:0] p66_bit_slice_2043893;
  reg [127:0] p66_bit_slice_2044018;
  reg [127:0] p66_k3;
  reg [127:0] p66_k2;
  reg [127:0] p66_k5;
  reg [127:0] p66_k4;
  reg [127:0] p66_k7;
  reg [127:0] p66_k6;
  reg [127:0] p66_xor_2055662;
  reg [127:0] p66_xor_2056114;
  reg [7:0] p66_array_index_2056130;
  reg [7:0] p66_array_index_2056131;
  reg [7:0] p66_array_index_2056132;
  reg [7:0] p66_array_index_2056133;
  reg [7:0] p66_array_index_2056134;
  reg [7:0] p66_array_index_2056135;
  reg [7:0] p66_array_index_2056137;
  reg [7:0] p66_array_index_2056139;
  reg [7:0] p66_array_index_2056140;
  reg [7:0] p66_array_index_2056141;
  reg [7:0] p66_array_index_2056142;
  reg [7:0] p66_array_index_2056143;
  reg [7:0] p66_array_index_2056146;
  reg [7:0] p66_array_index_2056147;
  reg [7:0] p66_array_index_2056148;
  reg [7:0] p66_array_index_2056149;
  reg [7:0] p66_array_index_2056150;
  reg [7:0] p66_array_index_2056151;
  reg [7:0] p66_array_index_2056152;
  reg [7:0] p66_array_index_2056154;
  reg [7:0] p66_res7__864;
  reg [7:0] p66_array_index_2056163;
  reg [7:0] p66_array_index_2056164;
  reg [7:0] p66_array_index_2056165;
  reg [7:0] p66_array_index_2056166;
  reg [7:0] p66_array_index_2056167;
  reg [7:0] p66_array_index_2056168;
  reg [7:0] p66_res7__866;
  reg [7:0] p67_literal_2043896[256];
  reg [7:0] p67_literal_2043910[256];
  reg [7:0] p67_literal_2043912[256];
  reg [7:0] p67_literal_2043914[256];
  reg [7:0] p67_literal_2043916[256];
  reg [7:0] p67_literal_2043918[256];
  reg [7:0] p67_literal_2043920[256];
  reg [7:0] p67_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p66_encoded <= p65_encoded;
    p66_bit_slice_2043893 <= p65_bit_slice_2043893;
    p66_bit_slice_2044018 <= p65_bit_slice_2044018;
    p66_k3 <= p65_k3;
    p66_k2 <= p65_k2;
    p66_k5 <= p65_k5;
    p66_k4 <= p65_k4;
    p66_k7 <= p65_k7;
    p66_k6 <= p65_k6;
    p66_xor_2055662 <= p65_xor_2055662;
    p66_xor_2056114 <= p66_xor_2056114_comb;
    p66_array_index_2056130 <= p66_array_index_2056130_comb;
    p66_array_index_2056131 <= p66_array_index_2056131_comb;
    p66_array_index_2056132 <= p66_array_index_2056132_comb;
    p66_array_index_2056133 <= p66_array_index_2056133_comb;
    p66_array_index_2056134 <= p66_array_index_2056134_comb;
    p66_array_index_2056135 <= p66_array_index_2056135_comb;
    p66_array_index_2056137 <= p66_array_index_2056137_comb;
    p66_array_index_2056139 <= p66_array_index_2056139_comb;
    p66_array_index_2056140 <= p66_array_index_2056140_comb;
    p66_array_index_2056141 <= p66_array_index_2056141_comb;
    p66_array_index_2056142 <= p66_array_index_2056142_comb;
    p66_array_index_2056143 <= p66_array_index_2056143_comb;
    p66_array_index_2056146 <= p66_array_index_2056146_comb;
    p66_array_index_2056147 <= p66_array_index_2056147_comb;
    p66_array_index_2056148 <= p66_array_index_2056148_comb;
    p66_array_index_2056149 <= p66_array_index_2056149_comb;
    p66_array_index_2056150 <= p66_array_index_2056150_comb;
    p66_array_index_2056151 <= p66_array_index_2056151_comb;
    p66_array_index_2056152 <= p66_array_index_2056152_comb;
    p66_array_index_2056154 <= p66_array_index_2056154_comb;
    p66_res7__864 <= p66_res7__864_comb;
    p66_array_index_2056163 <= p66_array_index_2056163_comb;
    p66_array_index_2056164 <= p66_array_index_2056164_comb;
    p66_array_index_2056165 <= p66_array_index_2056165_comb;
    p66_array_index_2056166 <= p66_array_index_2056166_comb;
    p66_array_index_2056167 <= p66_array_index_2056167_comb;
    p66_array_index_2056168 <= p66_array_index_2056168_comb;
    p66_res7__866 <= p66_res7__866_comb;
    p67_literal_2043896 <= p66_literal_2043896;
    p67_literal_2043910 <= p66_literal_2043910;
    p67_literal_2043912 <= p66_literal_2043912;
    p67_literal_2043914 <= p66_literal_2043914;
    p67_literal_2043916 <= p66_literal_2043916;
    p67_literal_2043918 <= p66_literal_2043918;
    p67_literal_2043920 <= p66_literal_2043920;
    p67_literal_2043923 <= p66_literal_2043923;
  end

  // ===== Pipe stage 67:
  wire [7:0] p67_array_index_2056272_comb;
  wire [7:0] p67_array_index_2056273_comb;
  wire [7:0] p67_array_index_2056274_comb;
  wire [7:0] p67_array_index_2056275_comb;
  wire [7:0] p67_array_index_2056276_comb;
  wire [7:0] p67_res7__868_comb;
  wire [7:0] p67_array_index_2056286_comb;
  wire [7:0] p67_array_index_2056287_comb;
  wire [7:0] p67_array_index_2056288_comb;
  wire [7:0] p67_array_index_2056289_comb;
  wire [7:0] p67_array_index_2056290_comb;
  wire [7:0] p67_res7__870_comb;
  wire [7:0] p67_array_index_2056301_comb;
  wire [7:0] p67_array_index_2056302_comb;
  wire [7:0] p67_array_index_2056303_comb;
  wire [7:0] p67_array_index_2056304_comb;
  wire [7:0] p67_res7__872_comb;
  wire [7:0] p67_array_index_2056314_comb;
  wire [7:0] p67_array_index_2056315_comb;
  wire [7:0] p67_array_index_2056316_comb;
  wire [7:0] p67_array_index_2056317_comb;
  wire [7:0] p67_res7__874_comb;
  wire [7:0] p67_array_index_2056328_comb;
  wire [7:0] p67_array_index_2056329_comb;
  wire [7:0] p67_array_index_2056330_comb;
  wire [7:0] p67_res7__876_comb;
  wire [7:0] p67_array_index_2056340_comb;
  wire [7:0] p67_array_index_2056341_comb;
  wire [7:0] p67_array_index_2056342_comb;
  wire [7:0] p67_res7__878_comb;
  wire [7:0] p67_array_index_2056353_comb;
  wire [7:0] p67_array_index_2056354_comb;
  wire [7:0] p67_res7__880_comb;
  assign p67_array_index_2056272_comb = p66_literal_2043912[p66_res7__864];
  assign p67_array_index_2056273_comb = p66_literal_2043914[p66_array_index_2056130];
  assign p67_array_index_2056274_comb = p66_literal_2043916[p66_array_index_2056131];
  assign p67_array_index_2056275_comb = p66_literal_2043918[p66_array_index_2056132];
  assign p67_array_index_2056276_comb = p66_literal_2043920[p66_array_index_2056133];
  assign p67_res7__868_comb = p66_literal_2043910[p66_res7__866] ^ p67_array_index_2056272_comb ^ p67_array_index_2056273_comb ^ p67_array_index_2056274_comb ^ p67_array_index_2056275_comb ^ p67_array_index_2056276_comb ^ p66_array_index_2056134 ^ p66_literal_2043923[p66_array_index_2056135] ^ p66_array_index_2056152 ^ p66_literal_2043920[p66_array_index_2056137] ^ p66_literal_2043918[p66_array_index_2056154] ^ p66_literal_2043916[p66_array_index_2056139] ^ p66_literal_2043914[p66_array_index_2056140] ^ p66_literal_2043912[p66_array_index_2056141] ^ p66_literal_2043910[p66_array_index_2056142] ^ p66_array_index_2056143;
  assign p67_array_index_2056286_comb = p66_literal_2043912[p66_res7__866];
  assign p67_array_index_2056287_comb = p66_literal_2043914[p66_res7__864];
  assign p67_array_index_2056288_comb = p66_literal_2043916[p66_array_index_2056130];
  assign p67_array_index_2056289_comb = p66_literal_2043918[p66_array_index_2056131];
  assign p67_array_index_2056290_comb = p66_literal_2043920[p66_array_index_2056132];
  assign p67_res7__870_comb = p66_literal_2043910[p67_res7__868_comb] ^ p67_array_index_2056286_comb ^ p67_array_index_2056287_comb ^ p67_array_index_2056288_comb ^ p67_array_index_2056289_comb ^ p67_array_index_2056290_comb ^ p66_array_index_2056133 ^ p66_literal_2043923[p66_array_index_2056134] ^ p66_array_index_2056135 ^ p66_literal_2043920[p66_array_index_2056152] ^ p66_literal_2043918[p66_array_index_2056137] ^ p66_literal_2043916[p66_array_index_2056154] ^ p66_literal_2043914[p66_array_index_2056139] ^ p66_literal_2043912[p66_array_index_2056140] ^ p66_literal_2043910[p66_array_index_2056141] ^ p66_array_index_2056142;
  assign p67_array_index_2056301_comb = p66_literal_2043914[p66_res7__866];
  assign p67_array_index_2056302_comb = p66_literal_2043916[p66_res7__864];
  assign p67_array_index_2056303_comb = p66_literal_2043918[p66_array_index_2056130];
  assign p67_array_index_2056304_comb = p66_literal_2043920[p66_array_index_2056131];
  assign p67_res7__872_comb = p66_literal_2043910[p67_res7__870_comb] ^ p66_literal_2043912[p67_res7__868_comb] ^ p67_array_index_2056301_comb ^ p67_array_index_2056302_comb ^ p67_array_index_2056303_comb ^ p67_array_index_2056304_comb ^ p66_array_index_2056132 ^ p66_literal_2043923[p66_array_index_2056133] ^ p66_array_index_2056134 ^ p66_array_index_2056151 ^ p66_literal_2043918[p66_array_index_2056152] ^ p66_literal_2043916[p66_array_index_2056137] ^ p66_literal_2043914[p66_array_index_2056154] ^ p66_literal_2043912[p66_array_index_2056139] ^ p66_literal_2043910[p66_array_index_2056140] ^ p66_array_index_2056141;
  assign p67_array_index_2056314_comb = p66_literal_2043914[p67_res7__868_comb];
  assign p67_array_index_2056315_comb = p66_literal_2043916[p66_res7__866];
  assign p67_array_index_2056316_comb = p66_literal_2043918[p66_res7__864];
  assign p67_array_index_2056317_comb = p66_literal_2043920[p66_array_index_2056130];
  assign p67_res7__874_comb = p66_literal_2043910[p67_res7__872_comb] ^ p66_literal_2043912[p67_res7__870_comb] ^ p67_array_index_2056314_comb ^ p67_array_index_2056315_comb ^ p67_array_index_2056316_comb ^ p67_array_index_2056317_comb ^ p66_array_index_2056131 ^ p66_literal_2043923[p66_array_index_2056132] ^ p66_array_index_2056133 ^ p66_array_index_2056168 ^ p66_literal_2043918[p66_array_index_2056135] ^ p66_literal_2043916[p66_array_index_2056152] ^ p66_literal_2043914[p66_array_index_2056137] ^ p66_literal_2043912[p66_array_index_2056154] ^ p66_literal_2043910[p66_array_index_2056139] ^ p66_array_index_2056140;
  assign p67_array_index_2056328_comb = p66_literal_2043916[p67_res7__868_comb];
  assign p67_array_index_2056329_comb = p66_literal_2043918[p66_res7__866];
  assign p67_array_index_2056330_comb = p66_literal_2043920[p66_res7__864];
  assign p67_res7__876_comb = p66_literal_2043910[p67_res7__874_comb] ^ p66_literal_2043912[p67_res7__872_comb] ^ p66_literal_2043914[p67_res7__870_comb] ^ p67_array_index_2056328_comb ^ p67_array_index_2056329_comb ^ p67_array_index_2056330_comb ^ p66_array_index_2056130 ^ p66_literal_2043923[p66_array_index_2056131] ^ p66_array_index_2056132 ^ p67_array_index_2056276_comb ^ p66_array_index_2056150 ^ p66_literal_2043916[p66_array_index_2056135] ^ p66_literal_2043914[p66_array_index_2056152] ^ p66_literal_2043912[p66_array_index_2056137] ^ p66_literal_2043910[p66_array_index_2056154] ^ p66_array_index_2056139;
  assign p67_array_index_2056340_comb = p66_literal_2043916[p67_res7__870_comb];
  assign p67_array_index_2056341_comb = p66_literal_2043918[p67_res7__868_comb];
  assign p67_array_index_2056342_comb = p66_literal_2043920[p66_res7__866];
  assign p67_res7__878_comb = p66_literal_2043910[p67_res7__876_comb] ^ p66_literal_2043912[p67_res7__874_comb] ^ p66_literal_2043914[p67_res7__872_comb] ^ p67_array_index_2056340_comb ^ p67_array_index_2056341_comb ^ p67_array_index_2056342_comb ^ p66_res7__864 ^ p66_literal_2043923[p66_array_index_2056130] ^ p66_array_index_2056131 ^ p67_array_index_2056290_comb ^ p66_array_index_2056167 ^ p66_literal_2043916[p66_array_index_2056134] ^ p66_literal_2043914[p66_array_index_2056135] ^ p66_literal_2043912[p66_array_index_2056152] ^ p66_literal_2043910[p66_array_index_2056137] ^ p66_array_index_2056154;
  assign p67_array_index_2056353_comb = p66_literal_2043918[p67_res7__870_comb];
  assign p67_array_index_2056354_comb = p66_literal_2043920[p67_res7__868_comb];
  assign p67_res7__880_comb = p66_literal_2043910[p67_res7__878_comb] ^ p66_literal_2043912[p67_res7__876_comb] ^ p66_literal_2043914[p67_res7__874_comb] ^ p66_literal_2043916[p67_res7__872_comb] ^ p67_array_index_2056353_comb ^ p67_array_index_2056354_comb ^ p66_res7__866 ^ p66_literal_2043923[p66_res7__864] ^ p66_array_index_2056130 ^ p67_array_index_2056304_comb ^ p67_array_index_2056275_comb ^ p66_array_index_2056149 ^ p66_literal_2043914[p66_array_index_2056134] ^ p66_literal_2043912[p66_array_index_2056135] ^ p66_literal_2043910[p66_array_index_2056152] ^ p66_array_index_2056137;

  // Registers for pipe stage 67:
  reg [127:0] p67_encoded;
  reg [127:0] p67_bit_slice_2043893;
  reg [127:0] p67_bit_slice_2044018;
  reg [127:0] p67_k3;
  reg [127:0] p67_k2;
  reg [127:0] p67_k5;
  reg [127:0] p67_k4;
  reg [127:0] p67_k7;
  reg [127:0] p67_k6;
  reg [127:0] p67_xor_2055662;
  reg [127:0] p67_xor_2056114;
  reg [7:0] p67_array_index_2056130;
  reg [7:0] p67_array_index_2056131;
  reg [7:0] p67_array_index_2056132;
  reg [7:0] p67_array_index_2056133;
  reg [7:0] p67_array_index_2056134;
  reg [7:0] p67_array_index_2056135;
  reg [7:0] p67_array_index_2056146;
  reg [7:0] p67_array_index_2056147;
  reg [7:0] p67_array_index_2056148;
  reg [7:0] p67_array_index_2056152;
  reg [7:0] p67_res7__864;
  reg [7:0] p67_array_index_2056163;
  reg [7:0] p67_array_index_2056164;
  reg [7:0] p67_array_index_2056165;
  reg [7:0] p67_array_index_2056166;
  reg [7:0] p67_res7__866;
  reg [7:0] p67_array_index_2056272;
  reg [7:0] p67_array_index_2056273;
  reg [7:0] p67_array_index_2056274;
  reg [7:0] p67_res7__868;
  reg [7:0] p67_array_index_2056286;
  reg [7:0] p67_array_index_2056287;
  reg [7:0] p67_array_index_2056288;
  reg [7:0] p67_array_index_2056289;
  reg [7:0] p67_res7__870;
  reg [7:0] p67_array_index_2056301;
  reg [7:0] p67_array_index_2056302;
  reg [7:0] p67_array_index_2056303;
  reg [7:0] p67_res7__872;
  reg [7:0] p67_array_index_2056314;
  reg [7:0] p67_array_index_2056315;
  reg [7:0] p67_array_index_2056316;
  reg [7:0] p67_array_index_2056317;
  reg [7:0] p67_res7__874;
  reg [7:0] p67_array_index_2056328;
  reg [7:0] p67_array_index_2056329;
  reg [7:0] p67_array_index_2056330;
  reg [7:0] p67_res7__876;
  reg [7:0] p67_array_index_2056340;
  reg [7:0] p67_array_index_2056341;
  reg [7:0] p67_array_index_2056342;
  reg [7:0] p67_res7__878;
  reg [7:0] p67_array_index_2056353;
  reg [7:0] p67_array_index_2056354;
  reg [7:0] p67_res7__880;
  reg [7:0] p68_literal_2043896[256];
  reg [7:0] p68_literal_2043910[256];
  reg [7:0] p68_literal_2043912[256];
  reg [7:0] p68_literal_2043914[256];
  reg [7:0] p68_literal_2043916[256];
  reg [7:0] p68_literal_2043918[256];
  reg [7:0] p68_literal_2043920[256];
  reg [7:0] p68_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p67_encoded <= p66_encoded;
    p67_bit_slice_2043893 <= p66_bit_slice_2043893;
    p67_bit_slice_2044018 <= p66_bit_slice_2044018;
    p67_k3 <= p66_k3;
    p67_k2 <= p66_k2;
    p67_k5 <= p66_k5;
    p67_k4 <= p66_k4;
    p67_k7 <= p66_k7;
    p67_k6 <= p66_k6;
    p67_xor_2055662 <= p66_xor_2055662;
    p67_xor_2056114 <= p66_xor_2056114;
    p67_array_index_2056130 <= p66_array_index_2056130;
    p67_array_index_2056131 <= p66_array_index_2056131;
    p67_array_index_2056132 <= p66_array_index_2056132;
    p67_array_index_2056133 <= p66_array_index_2056133;
    p67_array_index_2056134 <= p66_array_index_2056134;
    p67_array_index_2056135 <= p66_array_index_2056135;
    p67_array_index_2056146 <= p66_array_index_2056146;
    p67_array_index_2056147 <= p66_array_index_2056147;
    p67_array_index_2056148 <= p66_array_index_2056148;
    p67_array_index_2056152 <= p66_array_index_2056152;
    p67_res7__864 <= p66_res7__864;
    p67_array_index_2056163 <= p66_array_index_2056163;
    p67_array_index_2056164 <= p66_array_index_2056164;
    p67_array_index_2056165 <= p66_array_index_2056165;
    p67_array_index_2056166 <= p66_array_index_2056166;
    p67_res7__866 <= p66_res7__866;
    p67_array_index_2056272 <= p67_array_index_2056272_comb;
    p67_array_index_2056273 <= p67_array_index_2056273_comb;
    p67_array_index_2056274 <= p67_array_index_2056274_comb;
    p67_res7__868 <= p67_res7__868_comb;
    p67_array_index_2056286 <= p67_array_index_2056286_comb;
    p67_array_index_2056287 <= p67_array_index_2056287_comb;
    p67_array_index_2056288 <= p67_array_index_2056288_comb;
    p67_array_index_2056289 <= p67_array_index_2056289_comb;
    p67_res7__870 <= p67_res7__870_comb;
    p67_array_index_2056301 <= p67_array_index_2056301_comb;
    p67_array_index_2056302 <= p67_array_index_2056302_comb;
    p67_array_index_2056303 <= p67_array_index_2056303_comb;
    p67_res7__872 <= p67_res7__872_comb;
    p67_array_index_2056314 <= p67_array_index_2056314_comb;
    p67_array_index_2056315 <= p67_array_index_2056315_comb;
    p67_array_index_2056316 <= p67_array_index_2056316_comb;
    p67_array_index_2056317 <= p67_array_index_2056317_comb;
    p67_res7__874 <= p67_res7__874_comb;
    p67_array_index_2056328 <= p67_array_index_2056328_comb;
    p67_array_index_2056329 <= p67_array_index_2056329_comb;
    p67_array_index_2056330 <= p67_array_index_2056330_comb;
    p67_res7__876 <= p67_res7__876_comb;
    p67_array_index_2056340 <= p67_array_index_2056340_comb;
    p67_array_index_2056341 <= p67_array_index_2056341_comb;
    p67_array_index_2056342 <= p67_array_index_2056342_comb;
    p67_res7__878 <= p67_res7__878_comb;
    p67_array_index_2056353 <= p67_array_index_2056353_comb;
    p67_array_index_2056354 <= p67_array_index_2056354_comb;
    p67_res7__880 <= p67_res7__880_comb;
    p68_literal_2043896 <= p67_literal_2043896;
    p68_literal_2043910 <= p67_literal_2043910;
    p68_literal_2043912 <= p67_literal_2043912;
    p68_literal_2043914 <= p67_literal_2043914;
    p68_literal_2043916 <= p67_literal_2043916;
    p68_literal_2043918 <= p67_literal_2043918;
    p68_literal_2043920 <= p67_literal_2043920;
    p68_literal_2043923 <= p67_literal_2043923;
  end

  // ===== Pipe stage 68:
  wire [7:0] p68_array_index_2056492_comb;
  wire [7:0] p68_array_index_2056493_comb;
  wire [7:0] p68_res7__882_comb;
  wire [7:0] p68_array_index_2056504_comb;
  wire [7:0] p68_res7__884_comb;
  wire [7:0] p68_array_index_2056514_comb;
  wire [7:0] p68_res7__886_comb;
  wire [7:0] p68_res7__888_comb;
  wire [7:0] p68_res7__890_comb;
  wire [7:0] p68_res7__892_comb;
  wire [7:0] p68_res7__894_comb;
  wire [127:0] p68_res__27_comb;
  assign p68_array_index_2056492_comb = p67_literal_2043918[p67_res7__872];
  assign p68_array_index_2056493_comb = p67_literal_2043920[p67_res7__870];
  assign p68_res7__882_comb = p67_literal_2043910[p67_res7__880] ^ p67_literal_2043912[p67_res7__878] ^ p67_literal_2043914[p67_res7__876] ^ p67_literal_2043916[p67_res7__874] ^ p68_array_index_2056492_comb ^ p68_array_index_2056493_comb ^ p67_res7__868 ^ p67_literal_2043923[p67_res7__866] ^ p67_res7__864 ^ p67_array_index_2056317 ^ p67_array_index_2056289 ^ p67_array_index_2056166 ^ p67_literal_2043914[p67_array_index_2056133] ^ p67_literal_2043912[p67_array_index_2056134] ^ p67_literal_2043910[p67_array_index_2056135] ^ p67_array_index_2056152;
  assign p68_array_index_2056504_comb = p67_literal_2043920[p67_res7__872];
  assign p68_res7__884_comb = p67_literal_2043910[p68_res7__882_comb] ^ p67_literal_2043912[p67_res7__880] ^ p67_literal_2043914[p67_res7__878] ^ p67_literal_2043916[p67_res7__876] ^ p67_literal_2043918[p67_res7__874] ^ p68_array_index_2056504_comb ^ p67_res7__870 ^ p67_literal_2043923[p67_res7__868] ^ p67_res7__866 ^ p67_array_index_2056330 ^ p67_array_index_2056303 ^ p67_array_index_2056274 ^ p67_array_index_2056148 ^ p67_literal_2043912[p67_array_index_2056133] ^ p67_literal_2043910[p67_array_index_2056134] ^ p67_array_index_2056135;
  assign p68_array_index_2056514_comb = p67_literal_2043920[p67_res7__874];
  assign p68_res7__886_comb = p67_literal_2043910[p68_res7__884_comb] ^ p67_literal_2043912[p68_res7__882_comb] ^ p67_literal_2043914[p67_res7__880] ^ p67_literal_2043916[p67_res7__878] ^ p67_literal_2043918[p67_res7__876] ^ p68_array_index_2056514_comb ^ p67_res7__872 ^ p67_literal_2043923[p67_res7__870] ^ p67_res7__868 ^ p67_array_index_2056342 ^ p67_array_index_2056316 ^ p67_array_index_2056288 ^ p67_array_index_2056165 ^ p67_literal_2043912[p67_array_index_2056132] ^ p67_literal_2043910[p67_array_index_2056133] ^ p67_array_index_2056134;
  assign p68_res7__888_comb = p67_literal_2043910[p68_res7__886_comb] ^ p67_literal_2043912[p68_res7__884_comb] ^ p67_literal_2043914[p68_res7__882_comb] ^ p67_literal_2043916[p67_res7__880] ^ p67_literal_2043918[p67_res7__878] ^ p67_literal_2043920[p67_res7__876] ^ p67_res7__874 ^ p67_literal_2043923[p67_res7__872] ^ p67_res7__870 ^ p67_array_index_2056354 ^ p67_array_index_2056329 ^ p67_array_index_2056302 ^ p67_array_index_2056273 ^ p67_array_index_2056147 ^ p67_literal_2043910[p67_array_index_2056132] ^ p67_array_index_2056133;
  assign p68_res7__890_comb = p67_literal_2043910[p68_res7__888_comb] ^ p67_literal_2043912[p68_res7__886_comb] ^ p67_literal_2043914[p68_res7__884_comb] ^ p67_literal_2043916[p68_res7__882_comb] ^ p67_literal_2043918[p67_res7__880] ^ p67_literal_2043920[p67_res7__878] ^ p67_res7__876 ^ p67_literal_2043923[p67_res7__874] ^ p67_res7__872 ^ p68_array_index_2056493_comb ^ p67_array_index_2056341 ^ p67_array_index_2056315 ^ p67_array_index_2056287 ^ p67_array_index_2056164 ^ p67_literal_2043910[p67_array_index_2056131] ^ p67_array_index_2056132;
  assign p68_res7__892_comb = p67_literal_2043910[p68_res7__890_comb] ^ p67_literal_2043912[p68_res7__888_comb] ^ p67_literal_2043914[p68_res7__886_comb] ^ p67_literal_2043916[p68_res7__884_comb] ^ p67_literal_2043918[p68_res7__882_comb] ^ p67_literal_2043920[p67_res7__880] ^ p67_res7__878 ^ p67_literal_2043923[p67_res7__876] ^ p67_res7__874 ^ p68_array_index_2056504_comb ^ p67_array_index_2056353 ^ p67_array_index_2056328 ^ p67_array_index_2056301 ^ p67_array_index_2056272 ^ p67_array_index_2056146 ^ p67_array_index_2056131;
  assign p68_res7__894_comb = p67_literal_2043910[p68_res7__892_comb] ^ p67_literal_2043912[p68_res7__890_comb] ^ p67_literal_2043914[p68_res7__888_comb] ^ p67_literal_2043916[p68_res7__886_comb] ^ p67_literal_2043918[p68_res7__884_comb] ^ p67_literal_2043920[p68_res7__882_comb] ^ p67_res7__880 ^ p67_literal_2043923[p67_res7__878] ^ p67_res7__876 ^ p68_array_index_2056514_comb ^ p68_array_index_2056492_comb ^ p67_array_index_2056340 ^ p67_array_index_2056314 ^ p67_array_index_2056286 ^ p67_array_index_2056163 ^ p67_array_index_2056130;
  assign p68_res__27_comb = {p68_res7__894_comb, p68_res7__892_comb, p68_res7__890_comb, p68_res7__888_comb, p68_res7__886_comb, p68_res7__884_comb, p68_res7__882_comb, p67_res7__880, p67_res7__878, p67_res7__876, p67_res7__874, p67_res7__872, p67_res7__870, p67_res7__868, p67_res7__866, p67_res7__864};

  // Registers for pipe stage 68:
  reg [127:0] p68_encoded;
  reg [127:0] p68_bit_slice_2043893;
  reg [127:0] p68_bit_slice_2044018;
  reg [127:0] p68_k3;
  reg [127:0] p68_k2;
  reg [127:0] p68_k5;
  reg [127:0] p68_k4;
  reg [127:0] p68_k7;
  reg [127:0] p68_k6;
  reg [127:0] p68_xor_2055662;
  reg [127:0] p68_xor_2056114;
  reg [127:0] p68_res__27;
  reg [7:0] p69_literal_2043896[256];
  reg [7:0] p69_literal_2043910[256];
  reg [7:0] p69_literal_2043912[256];
  reg [7:0] p69_literal_2043914[256];
  reg [7:0] p69_literal_2043916[256];
  reg [7:0] p69_literal_2043918[256];
  reg [7:0] p69_literal_2043920[256];
  reg [7:0] p69_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p68_encoded <= p67_encoded;
    p68_bit_slice_2043893 <= p67_bit_slice_2043893;
    p68_bit_slice_2044018 <= p67_bit_slice_2044018;
    p68_k3 <= p67_k3;
    p68_k2 <= p67_k2;
    p68_k5 <= p67_k5;
    p68_k4 <= p67_k4;
    p68_k7 <= p67_k7;
    p68_k6 <= p67_k6;
    p68_xor_2055662 <= p67_xor_2055662;
    p68_xor_2056114 <= p67_xor_2056114;
    p68_res__27 <= p68_res__27_comb;
    p69_literal_2043896 <= p68_literal_2043896;
    p69_literal_2043910 <= p68_literal_2043910;
    p69_literal_2043912 <= p68_literal_2043912;
    p69_literal_2043914 <= p68_literal_2043914;
    p69_literal_2043916 <= p68_literal_2043916;
    p69_literal_2043918 <= p68_literal_2043918;
    p69_literal_2043920 <= p68_literal_2043920;
    p69_literal_2043923 <= p68_literal_2043923;
  end

  // ===== Pipe stage 69:
  wire [127:0] p69_xor_2056594_comb;
  wire [127:0] p69_addedKey__60_comb;
  wire [7:0] p69_array_index_2056610_comb;
  wire [7:0] p69_array_index_2056611_comb;
  wire [7:0] p69_array_index_2056612_comb;
  wire [7:0] p69_array_index_2056613_comb;
  wire [7:0] p69_array_index_2056614_comb;
  wire [7:0] p69_array_index_2056615_comb;
  wire [7:0] p69_array_index_2056617_comb;
  wire [7:0] p69_array_index_2056619_comb;
  wire [7:0] p69_array_index_2056620_comb;
  wire [7:0] p69_array_index_2056621_comb;
  wire [7:0] p69_array_index_2056622_comb;
  wire [7:0] p69_array_index_2056623_comb;
  wire [7:0] p69_array_index_2056624_comb;
  wire [7:0] p69_array_index_2056626_comb;
  wire [7:0] p69_array_index_2056627_comb;
  wire [7:0] p69_array_index_2056628_comb;
  wire [7:0] p69_array_index_2056629_comb;
  wire [7:0] p69_array_index_2056630_comb;
  wire [7:0] p69_array_index_2056631_comb;
  wire [7:0] p69_array_index_2056632_comb;
  wire [7:0] p69_array_index_2056634_comb;
  wire [7:0] p69_res7__896_comb;
  wire [7:0] p69_array_index_2056643_comb;
  wire [7:0] p69_array_index_2056644_comb;
  wire [7:0] p69_array_index_2056645_comb;
  wire [7:0] p69_array_index_2056646_comb;
  wire [7:0] p69_array_index_2056647_comb;
  wire [7:0] p69_array_index_2056648_comb;
  wire [7:0] p69_res7__898_comb;
  wire [7:0] p69_array_index_2056658_comb;
  wire [7:0] p69_array_index_2056659_comb;
  wire [7:0] p69_array_index_2056660_comb;
  wire [7:0] p69_array_index_2056661_comb;
  wire [7:0] p69_array_index_2056662_comb;
  wire [7:0] p69_res7__900_comb;
  wire [7:0] p69_array_index_2056672_comb;
  wire [7:0] p69_array_index_2056673_comb;
  wire [7:0] p69_array_index_2056674_comb;
  wire [7:0] p69_array_index_2056675_comb;
  wire [7:0] p69_array_index_2056676_comb;
  wire [7:0] p69_res7__902_comb;
  wire [7:0] p69_array_index_2056687_comb;
  wire [7:0] p69_array_index_2056688_comb;
  wire [7:0] p69_array_index_2056689_comb;
  wire [7:0] p69_array_index_2056690_comb;
  wire [7:0] p69_res7__904_comb;
  wire [7:0] p69_array_index_2056700_comb;
  wire [7:0] p69_array_index_2056701_comb;
  wire [7:0] p69_array_index_2056702_comb;
  wire [7:0] p69_array_index_2056703_comb;
  wire [7:0] p69_res7__906_comb;
  assign p69_xor_2056594_comb = p68_res__27 ^ p68_xor_2055662;
  assign p69_addedKey__60_comb = p69_xor_2056594_comb ^ 128'hcc84_3743_f6a4_ab45_de75_2c13_46ec_ff1d;
  assign p69_array_index_2056610_comb = p68_literal_2043896[p69_addedKey__60_comb[127:120]];
  assign p69_array_index_2056611_comb = p68_literal_2043896[p69_addedKey__60_comb[119:112]];
  assign p69_array_index_2056612_comb = p68_literal_2043896[p69_addedKey__60_comb[111:104]];
  assign p69_array_index_2056613_comb = p68_literal_2043896[p69_addedKey__60_comb[103:96]];
  assign p69_array_index_2056614_comb = p68_literal_2043896[p69_addedKey__60_comb[95:88]];
  assign p69_array_index_2056615_comb = p68_literal_2043896[p69_addedKey__60_comb[87:80]];
  assign p69_array_index_2056617_comb = p68_literal_2043896[p69_addedKey__60_comb[71:64]];
  assign p69_array_index_2056619_comb = p68_literal_2043896[p69_addedKey__60_comb[55:48]];
  assign p69_array_index_2056620_comb = p68_literal_2043896[p69_addedKey__60_comb[47:40]];
  assign p69_array_index_2056621_comb = p68_literal_2043896[p69_addedKey__60_comb[39:32]];
  assign p69_array_index_2056622_comb = p68_literal_2043896[p69_addedKey__60_comb[31:24]];
  assign p69_array_index_2056623_comb = p68_literal_2043896[p69_addedKey__60_comb[23:16]];
  assign p69_array_index_2056624_comb = p68_literal_2043896[p69_addedKey__60_comb[15:8]];
  assign p69_array_index_2056626_comb = p68_literal_2043910[p69_array_index_2056610_comb];
  assign p69_array_index_2056627_comb = p68_literal_2043912[p69_array_index_2056611_comb];
  assign p69_array_index_2056628_comb = p68_literal_2043914[p69_array_index_2056612_comb];
  assign p69_array_index_2056629_comb = p68_literal_2043916[p69_array_index_2056613_comb];
  assign p69_array_index_2056630_comb = p68_literal_2043918[p69_array_index_2056614_comb];
  assign p69_array_index_2056631_comb = p68_literal_2043920[p69_array_index_2056615_comb];
  assign p69_array_index_2056632_comb = p68_literal_2043896[p69_addedKey__60_comb[79:72]];
  assign p69_array_index_2056634_comb = p68_literal_2043896[p69_addedKey__60_comb[63:56]];
  assign p69_res7__896_comb = p69_array_index_2056626_comb ^ p69_array_index_2056627_comb ^ p69_array_index_2056628_comb ^ p69_array_index_2056629_comb ^ p69_array_index_2056630_comb ^ p69_array_index_2056631_comb ^ p69_array_index_2056632_comb ^ p68_literal_2043923[p69_array_index_2056617_comb] ^ p69_array_index_2056634_comb ^ p68_literal_2043920[p69_array_index_2056619_comb] ^ p68_literal_2043918[p69_array_index_2056620_comb] ^ p68_literal_2043916[p69_array_index_2056621_comb] ^ p68_literal_2043914[p69_array_index_2056622_comb] ^ p68_literal_2043912[p69_array_index_2056623_comb] ^ p68_literal_2043910[p69_array_index_2056624_comb] ^ p68_literal_2043896[p69_addedKey__60_comb[7:0]];
  assign p69_array_index_2056643_comb = p68_literal_2043910[p69_res7__896_comb];
  assign p69_array_index_2056644_comb = p68_literal_2043912[p69_array_index_2056610_comb];
  assign p69_array_index_2056645_comb = p68_literal_2043914[p69_array_index_2056611_comb];
  assign p69_array_index_2056646_comb = p68_literal_2043916[p69_array_index_2056612_comb];
  assign p69_array_index_2056647_comb = p68_literal_2043918[p69_array_index_2056613_comb];
  assign p69_array_index_2056648_comb = p68_literal_2043920[p69_array_index_2056614_comb];
  assign p69_res7__898_comb = p69_array_index_2056643_comb ^ p69_array_index_2056644_comb ^ p69_array_index_2056645_comb ^ p69_array_index_2056646_comb ^ p69_array_index_2056647_comb ^ p69_array_index_2056648_comb ^ p69_array_index_2056615_comb ^ p68_literal_2043923[p69_array_index_2056632_comb] ^ p69_array_index_2056617_comb ^ p68_literal_2043920[p69_array_index_2056634_comb] ^ p68_literal_2043918[p69_array_index_2056619_comb] ^ p68_literal_2043916[p69_array_index_2056620_comb] ^ p68_literal_2043914[p69_array_index_2056621_comb] ^ p68_literal_2043912[p69_array_index_2056622_comb] ^ p68_literal_2043910[p69_array_index_2056623_comb] ^ p69_array_index_2056624_comb;
  assign p69_array_index_2056658_comb = p68_literal_2043912[p69_res7__896_comb];
  assign p69_array_index_2056659_comb = p68_literal_2043914[p69_array_index_2056610_comb];
  assign p69_array_index_2056660_comb = p68_literal_2043916[p69_array_index_2056611_comb];
  assign p69_array_index_2056661_comb = p68_literal_2043918[p69_array_index_2056612_comb];
  assign p69_array_index_2056662_comb = p68_literal_2043920[p69_array_index_2056613_comb];
  assign p69_res7__900_comb = p68_literal_2043910[p69_res7__898_comb] ^ p69_array_index_2056658_comb ^ p69_array_index_2056659_comb ^ p69_array_index_2056660_comb ^ p69_array_index_2056661_comb ^ p69_array_index_2056662_comb ^ p69_array_index_2056614_comb ^ p68_literal_2043923[p69_array_index_2056615_comb] ^ p69_array_index_2056632_comb ^ p68_literal_2043920[p69_array_index_2056617_comb] ^ p68_literal_2043918[p69_array_index_2056634_comb] ^ p68_literal_2043916[p69_array_index_2056619_comb] ^ p68_literal_2043914[p69_array_index_2056620_comb] ^ p68_literal_2043912[p69_array_index_2056621_comb] ^ p68_literal_2043910[p69_array_index_2056622_comb] ^ p69_array_index_2056623_comb;
  assign p69_array_index_2056672_comb = p68_literal_2043912[p69_res7__898_comb];
  assign p69_array_index_2056673_comb = p68_literal_2043914[p69_res7__896_comb];
  assign p69_array_index_2056674_comb = p68_literal_2043916[p69_array_index_2056610_comb];
  assign p69_array_index_2056675_comb = p68_literal_2043918[p69_array_index_2056611_comb];
  assign p69_array_index_2056676_comb = p68_literal_2043920[p69_array_index_2056612_comb];
  assign p69_res7__902_comb = p68_literal_2043910[p69_res7__900_comb] ^ p69_array_index_2056672_comb ^ p69_array_index_2056673_comb ^ p69_array_index_2056674_comb ^ p69_array_index_2056675_comb ^ p69_array_index_2056676_comb ^ p69_array_index_2056613_comb ^ p68_literal_2043923[p69_array_index_2056614_comb] ^ p69_array_index_2056615_comb ^ p68_literal_2043920[p69_array_index_2056632_comb] ^ p68_literal_2043918[p69_array_index_2056617_comb] ^ p68_literal_2043916[p69_array_index_2056634_comb] ^ p68_literal_2043914[p69_array_index_2056619_comb] ^ p68_literal_2043912[p69_array_index_2056620_comb] ^ p68_literal_2043910[p69_array_index_2056621_comb] ^ p69_array_index_2056622_comb;
  assign p69_array_index_2056687_comb = p68_literal_2043914[p69_res7__898_comb];
  assign p69_array_index_2056688_comb = p68_literal_2043916[p69_res7__896_comb];
  assign p69_array_index_2056689_comb = p68_literal_2043918[p69_array_index_2056610_comb];
  assign p69_array_index_2056690_comb = p68_literal_2043920[p69_array_index_2056611_comb];
  assign p69_res7__904_comb = p68_literal_2043910[p69_res7__902_comb] ^ p68_literal_2043912[p69_res7__900_comb] ^ p69_array_index_2056687_comb ^ p69_array_index_2056688_comb ^ p69_array_index_2056689_comb ^ p69_array_index_2056690_comb ^ p69_array_index_2056612_comb ^ p68_literal_2043923[p69_array_index_2056613_comb] ^ p69_array_index_2056614_comb ^ p69_array_index_2056631_comb ^ p68_literal_2043918[p69_array_index_2056632_comb] ^ p68_literal_2043916[p69_array_index_2056617_comb] ^ p68_literal_2043914[p69_array_index_2056634_comb] ^ p68_literal_2043912[p69_array_index_2056619_comb] ^ p68_literal_2043910[p69_array_index_2056620_comb] ^ p69_array_index_2056621_comb;
  assign p69_array_index_2056700_comb = p68_literal_2043914[p69_res7__900_comb];
  assign p69_array_index_2056701_comb = p68_literal_2043916[p69_res7__898_comb];
  assign p69_array_index_2056702_comb = p68_literal_2043918[p69_res7__896_comb];
  assign p69_array_index_2056703_comb = p68_literal_2043920[p69_array_index_2056610_comb];
  assign p69_res7__906_comb = p68_literal_2043910[p69_res7__904_comb] ^ p68_literal_2043912[p69_res7__902_comb] ^ p69_array_index_2056700_comb ^ p69_array_index_2056701_comb ^ p69_array_index_2056702_comb ^ p69_array_index_2056703_comb ^ p69_array_index_2056611_comb ^ p68_literal_2043923[p69_array_index_2056612_comb] ^ p69_array_index_2056613_comb ^ p69_array_index_2056648_comb ^ p68_literal_2043918[p69_array_index_2056615_comb] ^ p68_literal_2043916[p69_array_index_2056632_comb] ^ p68_literal_2043914[p69_array_index_2056617_comb] ^ p68_literal_2043912[p69_array_index_2056634_comb] ^ p68_literal_2043910[p69_array_index_2056619_comb] ^ p69_array_index_2056620_comb;

  // Registers for pipe stage 69:
  reg [127:0] p69_encoded;
  reg [127:0] p69_bit_slice_2043893;
  reg [127:0] p69_bit_slice_2044018;
  reg [127:0] p69_k3;
  reg [127:0] p69_k2;
  reg [127:0] p69_k5;
  reg [127:0] p69_k4;
  reg [127:0] p69_k7;
  reg [127:0] p69_k6;
  reg [127:0] p69_xor_2056114;
  reg [127:0] p69_xor_2056594;
  reg [7:0] p69_array_index_2056610;
  reg [7:0] p69_array_index_2056611;
  reg [7:0] p69_array_index_2056612;
  reg [7:0] p69_array_index_2056613;
  reg [7:0] p69_array_index_2056614;
  reg [7:0] p69_array_index_2056615;
  reg [7:0] p69_array_index_2056617;
  reg [7:0] p69_array_index_2056619;
  reg [7:0] p69_array_index_2056626;
  reg [7:0] p69_array_index_2056627;
  reg [7:0] p69_array_index_2056628;
  reg [7:0] p69_array_index_2056629;
  reg [7:0] p69_array_index_2056630;
  reg [7:0] p69_array_index_2056632;
  reg [7:0] p69_array_index_2056634;
  reg [7:0] p69_res7__896;
  reg [7:0] p69_array_index_2056643;
  reg [7:0] p69_array_index_2056644;
  reg [7:0] p69_array_index_2056645;
  reg [7:0] p69_array_index_2056646;
  reg [7:0] p69_array_index_2056647;
  reg [7:0] p69_res7__898;
  reg [7:0] p69_array_index_2056658;
  reg [7:0] p69_array_index_2056659;
  reg [7:0] p69_array_index_2056660;
  reg [7:0] p69_array_index_2056661;
  reg [7:0] p69_array_index_2056662;
  reg [7:0] p69_res7__900;
  reg [7:0] p69_array_index_2056672;
  reg [7:0] p69_array_index_2056673;
  reg [7:0] p69_array_index_2056674;
  reg [7:0] p69_array_index_2056675;
  reg [7:0] p69_array_index_2056676;
  reg [7:0] p69_res7__902;
  reg [7:0] p69_array_index_2056687;
  reg [7:0] p69_array_index_2056688;
  reg [7:0] p69_array_index_2056689;
  reg [7:0] p69_array_index_2056690;
  reg [7:0] p69_res7__904;
  reg [7:0] p69_array_index_2056700;
  reg [7:0] p69_array_index_2056701;
  reg [7:0] p69_array_index_2056702;
  reg [7:0] p69_array_index_2056703;
  reg [7:0] p69_res7__906;
  reg [7:0] p70_literal_2043896[256];
  reg [7:0] p70_literal_2043910[256];
  reg [7:0] p70_literal_2043912[256];
  reg [7:0] p70_literal_2043914[256];
  reg [7:0] p70_literal_2043916[256];
  reg [7:0] p70_literal_2043918[256];
  reg [7:0] p70_literal_2043920[256];
  reg [7:0] p70_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p69_encoded <= p68_encoded;
    p69_bit_slice_2043893 <= p68_bit_slice_2043893;
    p69_bit_slice_2044018 <= p68_bit_slice_2044018;
    p69_k3 <= p68_k3;
    p69_k2 <= p68_k2;
    p69_k5 <= p68_k5;
    p69_k4 <= p68_k4;
    p69_k7 <= p68_k7;
    p69_k6 <= p68_k6;
    p69_xor_2056114 <= p68_xor_2056114;
    p69_xor_2056594 <= p69_xor_2056594_comb;
    p69_array_index_2056610 <= p69_array_index_2056610_comb;
    p69_array_index_2056611 <= p69_array_index_2056611_comb;
    p69_array_index_2056612 <= p69_array_index_2056612_comb;
    p69_array_index_2056613 <= p69_array_index_2056613_comb;
    p69_array_index_2056614 <= p69_array_index_2056614_comb;
    p69_array_index_2056615 <= p69_array_index_2056615_comb;
    p69_array_index_2056617 <= p69_array_index_2056617_comb;
    p69_array_index_2056619 <= p69_array_index_2056619_comb;
    p69_array_index_2056626 <= p69_array_index_2056626_comb;
    p69_array_index_2056627 <= p69_array_index_2056627_comb;
    p69_array_index_2056628 <= p69_array_index_2056628_comb;
    p69_array_index_2056629 <= p69_array_index_2056629_comb;
    p69_array_index_2056630 <= p69_array_index_2056630_comb;
    p69_array_index_2056632 <= p69_array_index_2056632_comb;
    p69_array_index_2056634 <= p69_array_index_2056634_comb;
    p69_res7__896 <= p69_res7__896_comb;
    p69_array_index_2056643 <= p69_array_index_2056643_comb;
    p69_array_index_2056644 <= p69_array_index_2056644_comb;
    p69_array_index_2056645 <= p69_array_index_2056645_comb;
    p69_array_index_2056646 <= p69_array_index_2056646_comb;
    p69_array_index_2056647 <= p69_array_index_2056647_comb;
    p69_res7__898 <= p69_res7__898_comb;
    p69_array_index_2056658 <= p69_array_index_2056658_comb;
    p69_array_index_2056659 <= p69_array_index_2056659_comb;
    p69_array_index_2056660 <= p69_array_index_2056660_comb;
    p69_array_index_2056661 <= p69_array_index_2056661_comb;
    p69_array_index_2056662 <= p69_array_index_2056662_comb;
    p69_res7__900 <= p69_res7__900_comb;
    p69_array_index_2056672 <= p69_array_index_2056672_comb;
    p69_array_index_2056673 <= p69_array_index_2056673_comb;
    p69_array_index_2056674 <= p69_array_index_2056674_comb;
    p69_array_index_2056675 <= p69_array_index_2056675_comb;
    p69_array_index_2056676 <= p69_array_index_2056676_comb;
    p69_res7__902 <= p69_res7__902_comb;
    p69_array_index_2056687 <= p69_array_index_2056687_comb;
    p69_array_index_2056688 <= p69_array_index_2056688_comb;
    p69_array_index_2056689 <= p69_array_index_2056689_comb;
    p69_array_index_2056690 <= p69_array_index_2056690_comb;
    p69_res7__904 <= p69_res7__904_comb;
    p69_array_index_2056700 <= p69_array_index_2056700_comb;
    p69_array_index_2056701 <= p69_array_index_2056701_comb;
    p69_array_index_2056702 <= p69_array_index_2056702_comb;
    p69_array_index_2056703 <= p69_array_index_2056703_comb;
    p69_res7__906 <= p69_res7__906_comb;
    p70_literal_2043896 <= p69_literal_2043896;
    p70_literal_2043910 <= p69_literal_2043910;
    p70_literal_2043912 <= p69_literal_2043912;
    p70_literal_2043914 <= p69_literal_2043914;
    p70_literal_2043916 <= p69_literal_2043916;
    p70_literal_2043918 <= p69_literal_2043918;
    p70_literal_2043920 <= p69_literal_2043920;
    p70_literal_2043923 <= p69_literal_2043923;
  end

  // ===== Pipe stage 70:
  wire [7:0] p70_array_index_2056840_comb;
  wire [7:0] p70_array_index_2056841_comb;
  wire [7:0] p70_array_index_2056842_comb;
  wire [7:0] p70_res7__908_comb;
  wire [7:0] p70_array_index_2056852_comb;
  wire [7:0] p70_array_index_2056853_comb;
  wire [7:0] p70_array_index_2056854_comb;
  wire [7:0] p70_res7__910_comb;
  wire [7:0] p70_array_index_2056865_comb;
  wire [7:0] p70_array_index_2056866_comb;
  wire [7:0] p70_res7__912_comb;
  wire [7:0] p70_array_index_2056876_comb;
  wire [7:0] p70_array_index_2056877_comb;
  wire [7:0] p70_res7__914_comb;
  wire [7:0] p70_array_index_2056888_comb;
  wire [7:0] p70_res7__916_comb;
  wire [7:0] p70_array_index_2056898_comb;
  wire [7:0] p70_res7__918_comb;
  wire [7:0] p70_res7__920_comb;
  assign p70_array_index_2056840_comb = p69_literal_2043916[p69_res7__900];
  assign p70_array_index_2056841_comb = p69_literal_2043918[p69_res7__898];
  assign p70_array_index_2056842_comb = p69_literal_2043920[p69_res7__896];
  assign p70_res7__908_comb = p69_literal_2043910[p69_res7__906] ^ p69_literal_2043912[p69_res7__904] ^ p69_literal_2043914[p69_res7__902] ^ p70_array_index_2056840_comb ^ p70_array_index_2056841_comb ^ p70_array_index_2056842_comb ^ p69_array_index_2056610 ^ p69_literal_2043923[p69_array_index_2056611] ^ p69_array_index_2056612 ^ p69_array_index_2056662 ^ p69_array_index_2056630 ^ p69_literal_2043916[p69_array_index_2056615] ^ p69_literal_2043914[p69_array_index_2056632] ^ p69_literal_2043912[p69_array_index_2056617] ^ p69_literal_2043910[p69_array_index_2056634] ^ p69_array_index_2056619;
  assign p70_array_index_2056852_comb = p69_literal_2043916[p69_res7__902];
  assign p70_array_index_2056853_comb = p69_literal_2043918[p69_res7__900];
  assign p70_array_index_2056854_comb = p69_literal_2043920[p69_res7__898];
  assign p70_res7__910_comb = p69_literal_2043910[p70_res7__908_comb] ^ p69_literal_2043912[p69_res7__906] ^ p69_literal_2043914[p69_res7__904] ^ p70_array_index_2056852_comb ^ p70_array_index_2056853_comb ^ p70_array_index_2056854_comb ^ p69_res7__896 ^ p69_literal_2043923[p69_array_index_2056610] ^ p69_array_index_2056611 ^ p69_array_index_2056676 ^ p69_array_index_2056647 ^ p69_literal_2043916[p69_array_index_2056614] ^ p69_literal_2043914[p69_array_index_2056615] ^ p69_literal_2043912[p69_array_index_2056632] ^ p69_literal_2043910[p69_array_index_2056617] ^ p69_array_index_2056634;
  assign p70_array_index_2056865_comb = p69_literal_2043918[p69_res7__902];
  assign p70_array_index_2056866_comb = p69_literal_2043920[p69_res7__900];
  assign p70_res7__912_comb = p69_literal_2043910[p70_res7__910_comb] ^ p69_literal_2043912[p70_res7__908_comb] ^ p69_literal_2043914[p69_res7__906] ^ p69_literal_2043916[p69_res7__904] ^ p70_array_index_2056865_comb ^ p70_array_index_2056866_comb ^ p69_res7__898 ^ p69_literal_2043923[p69_res7__896] ^ p69_array_index_2056610 ^ p69_array_index_2056690 ^ p69_array_index_2056661 ^ p69_array_index_2056629 ^ p69_literal_2043914[p69_array_index_2056614] ^ p69_literal_2043912[p69_array_index_2056615] ^ p69_literal_2043910[p69_array_index_2056632] ^ p69_array_index_2056617;
  assign p70_array_index_2056876_comb = p69_literal_2043918[p69_res7__904];
  assign p70_array_index_2056877_comb = p69_literal_2043920[p69_res7__902];
  assign p70_res7__914_comb = p69_literal_2043910[p70_res7__912_comb] ^ p69_literal_2043912[p70_res7__910_comb] ^ p69_literal_2043914[p70_res7__908_comb] ^ p69_literal_2043916[p69_res7__906] ^ p70_array_index_2056876_comb ^ p70_array_index_2056877_comb ^ p69_res7__900 ^ p69_literal_2043923[p69_res7__898] ^ p69_res7__896 ^ p69_array_index_2056703 ^ p69_array_index_2056675 ^ p69_array_index_2056646 ^ p69_literal_2043914[p69_array_index_2056613] ^ p69_literal_2043912[p69_array_index_2056614] ^ p69_literal_2043910[p69_array_index_2056615] ^ p69_array_index_2056632;
  assign p70_array_index_2056888_comb = p69_literal_2043920[p69_res7__904];
  assign p70_res7__916_comb = p69_literal_2043910[p70_res7__914_comb] ^ p69_literal_2043912[p70_res7__912_comb] ^ p69_literal_2043914[p70_res7__910_comb] ^ p69_literal_2043916[p70_res7__908_comb] ^ p69_literal_2043918[p69_res7__906] ^ p70_array_index_2056888_comb ^ p69_res7__902 ^ p69_literal_2043923[p69_res7__900] ^ p69_res7__898 ^ p70_array_index_2056842_comb ^ p69_array_index_2056689 ^ p69_array_index_2056660 ^ p69_array_index_2056628 ^ p69_literal_2043912[p69_array_index_2056613] ^ p69_literal_2043910[p69_array_index_2056614] ^ p69_array_index_2056615;
  assign p70_array_index_2056898_comb = p69_literal_2043920[p69_res7__906];
  assign p70_res7__918_comb = p69_literal_2043910[p70_res7__916_comb] ^ p69_literal_2043912[p70_res7__914_comb] ^ p69_literal_2043914[p70_res7__912_comb] ^ p69_literal_2043916[p70_res7__910_comb] ^ p69_literal_2043918[p70_res7__908_comb] ^ p70_array_index_2056898_comb ^ p69_res7__904 ^ p69_literal_2043923[p69_res7__902] ^ p69_res7__900 ^ p70_array_index_2056854_comb ^ p69_array_index_2056702 ^ p69_array_index_2056674 ^ p69_array_index_2056645 ^ p69_literal_2043912[p69_array_index_2056612] ^ p69_literal_2043910[p69_array_index_2056613] ^ p69_array_index_2056614;
  assign p70_res7__920_comb = p69_literal_2043910[p70_res7__918_comb] ^ p69_literal_2043912[p70_res7__916_comb] ^ p69_literal_2043914[p70_res7__914_comb] ^ p69_literal_2043916[p70_res7__912_comb] ^ p69_literal_2043918[p70_res7__910_comb] ^ p69_literal_2043920[p70_res7__908_comb] ^ p69_res7__906 ^ p69_literal_2043923[p69_res7__904] ^ p69_res7__902 ^ p70_array_index_2056866_comb ^ p70_array_index_2056841_comb ^ p69_array_index_2056688 ^ p69_array_index_2056659 ^ p69_array_index_2056627 ^ p69_literal_2043910[p69_array_index_2056612] ^ p69_array_index_2056613;

  // Registers for pipe stage 70:
  reg [127:0] p70_encoded;
  reg [127:0] p70_bit_slice_2043893;
  reg [127:0] p70_bit_slice_2044018;
  reg [127:0] p70_k3;
  reg [127:0] p70_k2;
  reg [127:0] p70_k5;
  reg [127:0] p70_k4;
  reg [127:0] p70_k7;
  reg [127:0] p70_k6;
  reg [127:0] p70_xor_2056114;
  reg [127:0] p70_xor_2056594;
  reg [7:0] p70_array_index_2056610;
  reg [7:0] p70_array_index_2056611;
  reg [7:0] p70_array_index_2056612;
  reg [7:0] p70_array_index_2056626;
  reg [7:0] p70_res7__896;
  reg [7:0] p70_array_index_2056643;
  reg [7:0] p70_array_index_2056644;
  reg [7:0] p70_res7__898;
  reg [7:0] p70_array_index_2056658;
  reg [7:0] p70_res7__900;
  reg [7:0] p70_array_index_2056672;
  reg [7:0] p70_array_index_2056673;
  reg [7:0] p70_res7__902;
  reg [7:0] p70_array_index_2056687;
  reg [7:0] p70_res7__904;
  reg [7:0] p70_array_index_2056700;
  reg [7:0] p70_array_index_2056701;
  reg [7:0] p70_res7__906;
  reg [7:0] p70_array_index_2056840;
  reg [7:0] p70_res7__908;
  reg [7:0] p70_array_index_2056852;
  reg [7:0] p70_array_index_2056853;
  reg [7:0] p70_res7__910;
  reg [7:0] p70_array_index_2056865;
  reg [7:0] p70_res7__912;
  reg [7:0] p70_array_index_2056876;
  reg [7:0] p70_array_index_2056877;
  reg [7:0] p70_res7__914;
  reg [7:0] p70_array_index_2056888;
  reg [7:0] p70_res7__916;
  reg [7:0] p70_array_index_2056898;
  reg [7:0] p70_res7__918;
  reg [7:0] p70_res7__920;
  reg [7:0] p71_literal_2043896[256];
  reg [7:0] p71_literal_2043910[256];
  reg [7:0] p71_literal_2043912[256];
  reg [7:0] p71_literal_2043914[256];
  reg [7:0] p71_literal_2043916[256];
  reg [7:0] p71_literal_2043918[256];
  reg [7:0] p71_literal_2043920[256];
  reg [7:0] p71_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p70_encoded <= p69_encoded;
    p70_bit_slice_2043893 <= p69_bit_slice_2043893;
    p70_bit_slice_2044018 <= p69_bit_slice_2044018;
    p70_k3 <= p69_k3;
    p70_k2 <= p69_k2;
    p70_k5 <= p69_k5;
    p70_k4 <= p69_k4;
    p70_k7 <= p69_k7;
    p70_k6 <= p69_k6;
    p70_xor_2056114 <= p69_xor_2056114;
    p70_xor_2056594 <= p69_xor_2056594;
    p70_array_index_2056610 <= p69_array_index_2056610;
    p70_array_index_2056611 <= p69_array_index_2056611;
    p70_array_index_2056612 <= p69_array_index_2056612;
    p70_array_index_2056626 <= p69_array_index_2056626;
    p70_res7__896 <= p69_res7__896;
    p70_array_index_2056643 <= p69_array_index_2056643;
    p70_array_index_2056644 <= p69_array_index_2056644;
    p70_res7__898 <= p69_res7__898;
    p70_array_index_2056658 <= p69_array_index_2056658;
    p70_res7__900 <= p69_res7__900;
    p70_array_index_2056672 <= p69_array_index_2056672;
    p70_array_index_2056673 <= p69_array_index_2056673;
    p70_res7__902 <= p69_res7__902;
    p70_array_index_2056687 <= p69_array_index_2056687;
    p70_res7__904 <= p69_res7__904;
    p70_array_index_2056700 <= p69_array_index_2056700;
    p70_array_index_2056701 <= p69_array_index_2056701;
    p70_res7__906 <= p69_res7__906;
    p70_array_index_2056840 <= p70_array_index_2056840_comb;
    p70_res7__908 <= p70_res7__908_comb;
    p70_array_index_2056852 <= p70_array_index_2056852_comb;
    p70_array_index_2056853 <= p70_array_index_2056853_comb;
    p70_res7__910 <= p70_res7__910_comb;
    p70_array_index_2056865 <= p70_array_index_2056865_comb;
    p70_res7__912 <= p70_res7__912_comb;
    p70_array_index_2056876 <= p70_array_index_2056876_comb;
    p70_array_index_2056877 <= p70_array_index_2056877_comb;
    p70_res7__914 <= p70_res7__914_comb;
    p70_array_index_2056888 <= p70_array_index_2056888_comb;
    p70_res7__916 <= p70_res7__916_comb;
    p70_array_index_2056898 <= p70_array_index_2056898_comb;
    p70_res7__918 <= p70_res7__918_comb;
    p70_res7__920 <= p70_res7__920_comb;
    p71_literal_2043896 <= p70_literal_2043896;
    p71_literal_2043910 <= p70_literal_2043910;
    p71_literal_2043912 <= p70_literal_2043912;
    p71_literal_2043914 <= p70_literal_2043914;
    p71_literal_2043916 <= p70_literal_2043916;
    p71_literal_2043918 <= p70_literal_2043918;
    p71_literal_2043920 <= p70_literal_2043920;
    p71_literal_2043923 <= p70_literal_2043923;
  end

  // ===== Pipe stage 71:
  wire [7:0] p71_res7__922_comb;
  wire [7:0] p71_res7__924_comb;
  wire [7:0] p71_res7__926_comb;
  wire [127:0] p71_res__28_comb;
  wire [127:0] p71_xor_2057042_comb;
  wire [127:0] p71_addedKey__61_comb;
  wire [7:0] p71_array_index_2057058_comb;
  wire [7:0] p71_array_index_2057059_comb;
  wire [7:0] p71_array_index_2057060_comb;
  wire [7:0] p71_array_index_2057061_comb;
  wire [7:0] p71_array_index_2057062_comb;
  wire [7:0] p71_array_index_2057063_comb;
  wire [7:0] p71_array_index_2057065_comb;
  wire [7:0] p71_array_index_2057067_comb;
  wire [7:0] p71_array_index_2057068_comb;
  wire [7:0] p71_array_index_2057069_comb;
  wire [7:0] p71_array_index_2057070_comb;
  wire [7:0] p71_array_index_2057071_comb;
  wire [7:0] p71_array_index_2057072_comb;
  wire [7:0] p71_array_index_2057074_comb;
  wire [7:0] p71_array_index_2057075_comb;
  wire [7:0] p71_array_index_2057076_comb;
  wire [7:0] p71_array_index_2057077_comb;
  wire [7:0] p71_array_index_2057078_comb;
  wire [7:0] p71_array_index_2057079_comb;
  wire [7:0] p71_array_index_2057080_comb;
  wire [7:0] p71_array_index_2057082_comb;
  wire [7:0] p71_res7__928_comb;
  wire [7:0] p71_array_index_2057091_comb;
  wire [7:0] p71_array_index_2057092_comb;
  wire [7:0] p71_array_index_2057093_comb;
  wire [7:0] p71_array_index_2057094_comb;
  wire [7:0] p71_array_index_2057095_comb;
  wire [7:0] p71_array_index_2057096_comb;
  wire [7:0] p71_res7__930_comb;
  wire [7:0] p71_array_index_2057106_comb;
  wire [7:0] p71_array_index_2057107_comb;
  wire [7:0] p71_array_index_2057108_comb;
  wire [7:0] p71_array_index_2057109_comb;
  wire [7:0] p71_array_index_2057110_comb;
  wire [7:0] p71_res7__932_comb;
  assign p71_res7__922_comb = p70_literal_2043910[p70_res7__920] ^ p70_literal_2043912[p70_res7__918] ^ p70_literal_2043914[p70_res7__916] ^ p70_literal_2043916[p70_res7__914] ^ p70_literal_2043918[p70_res7__912] ^ p70_literal_2043920[p70_res7__910] ^ p70_res7__908 ^ p70_literal_2043923[p70_res7__906] ^ p70_res7__904 ^ p70_array_index_2056877 ^ p70_array_index_2056853 ^ p70_array_index_2056701 ^ p70_array_index_2056673 ^ p70_array_index_2056644 ^ p70_literal_2043910[p70_array_index_2056611] ^ p70_array_index_2056612;
  assign p71_res7__924_comb = p70_literal_2043910[p71_res7__922_comb] ^ p70_literal_2043912[p70_res7__920] ^ p70_literal_2043914[p70_res7__918] ^ p70_literal_2043916[p70_res7__916] ^ p70_literal_2043918[p70_res7__914] ^ p70_literal_2043920[p70_res7__912] ^ p70_res7__910 ^ p70_literal_2043923[p70_res7__908] ^ p70_res7__906 ^ p70_array_index_2056888 ^ p70_array_index_2056865 ^ p70_array_index_2056840 ^ p70_array_index_2056687 ^ p70_array_index_2056658 ^ p70_array_index_2056626 ^ p70_array_index_2056611;
  assign p71_res7__926_comb = p70_literal_2043910[p71_res7__924_comb] ^ p70_literal_2043912[p71_res7__922_comb] ^ p70_literal_2043914[p70_res7__920] ^ p70_literal_2043916[p70_res7__918] ^ p70_literal_2043918[p70_res7__916] ^ p70_literal_2043920[p70_res7__914] ^ p70_res7__912 ^ p70_literal_2043923[p70_res7__910] ^ p70_res7__908 ^ p70_array_index_2056898 ^ p70_array_index_2056876 ^ p70_array_index_2056852 ^ p70_array_index_2056700 ^ p70_array_index_2056672 ^ p70_array_index_2056643 ^ p70_array_index_2056610;
  assign p71_res__28_comb = {p71_res7__926_comb, p71_res7__924_comb, p71_res7__922_comb, p70_res7__920, p70_res7__918, p70_res7__916, p70_res7__914, p70_res7__912, p70_res7__910, p70_res7__908, p70_res7__906, p70_res7__904, p70_res7__902, p70_res7__900, p70_res7__898, p70_res7__896};
  assign p71_xor_2057042_comb = p71_res__28_comb ^ p70_xor_2056114;
  assign p71_addedKey__61_comb = p71_xor_2057042_comb ^ 128'h7ea1_add5_427c_254e_391c_2823_e2a3_801e;
  assign p71_array_index_2057058_comb = p70_literal_2043896[p71_addedKey__61_comb[127:120]];
  assign p71_array_index_2057059_comb = p70_literal_2043896[p71_addedKey__61_comb[119:112]];
  assign p71_array_index_2057060_comb = p70_literal_2043896[p71_addedKey__61_comb[111:104]];
  assign p71_array_index_2057061_comb = p70_literal_2043896[p71_addedKey__61_comb[103:96]];
  assign p71_array_index_2057062_comb = p70_literal_2043896[p71_addedKey__61_comb[95:88]];
  assign p71_array_index_2057063_comb = p70_literal_2043896[p71_addedKey__61_comb[87:80]];
  assign p71_array_index_2057065_comb = p70_literal_2043896[p71_addedKey__61_comb[71:64]];
  assign p71_array_index_2057067_comb = p70_literal_2043896[p71_addedKey__61_comb[55:48]];
  assign p71_array_index_2057068_comb = p70_literal_2043896[p71_addedKey__61_comb[47:40]];
  assign p71_array_index_2057069_comb = p70_literal_2043896[p71_addedKey__61_comb[39:32]];
  assign p71_array_index_2057070_comb = p70_literal_2043896[p71_addedKey__61_comb[31:24]];
  assign p71_array_index_2057071_comb = p70_literal_2043896[p71_addedKey__61_comb[23:16]];
  assign p71_array_index_2057072_comb = p70_literal_2043896[p71_addedKey__61_comb[15:8]];
  assign p71_array_index_2057074_comb = p70_literal_2043910[p71_array_index_2057058_comb];
  assign p71_array_index_2057075_comb = p70_literal_2043912[p71_array_index_2057059_comb];
  assign p71_array_index_2057076_comb = p70_literal_2043914[p71_array_index_2057060_comb];
  assign p71_array_index_2057077_comb = p70_literal_2043916[p71_array_index_2057061_comb];
  assign p71_array_index_2057078_comb = p70_literal_2043918[p71_array_index_2057062_comb];
  assign p71_array_index_2057079_comb = p70_literal_2043920[p71_array_index_2057063_comb];
  assign p71_array_index_2057080_comb = p70_literal_2043896[p71_addedKey__61_comb[79:72]];
  assign p71_array_index_2057082_comb = p70_literal_2043896[p71_addedKey__61_comb[63:56]];
  assign p71_res7__928_comb = p71_array_index_2057074_comb ^ p71_array_index_2057075_comb ^ p71_array_index_2057076_comb ^ p71_array_index_2057077_comb ^ p71_array_index_2057078_comb ^ p71_array_index_2057079_comb ^ p71_array_index_2057080_comb ^ p70_literal_2043923[p71_array_index_2057065_comb] ^ p71_array_index_2057082_comb ^ p70_literal_2043920[p71_array_index_2057067_comb] ^ p70_literal_2043918[p71_array_index_2057068_comb] ^ p70_literal_2043916[p71_array_index_2057069_comb] ^ p70_literal_2043914[p71_array_index_2057070_comb] ^ p70_literal_2043912[p71_array_index_2057071_comb] ^ p70_literal_2043910[p71_array_index_2057072_comb] ^ p70_literal_2043896[p71_addedKey__61_comb[7:0]];
  assign p71_array_index_2057091_comb = p70_literal_2043910[p71_res7__928_comb];
  assign p71_array_index_2057092_comb = p70_literal_2043912[p71_array_index_2057058_comb];
  assign p71_array_index_2057093_comb = p70_literal_2043914[p71_array_index_2057059_comb];
  assign p71_array_index_2057094_comb = p70_literal_2043916[p71_array_index_2057060_comb];
  assign p71_array_index_2057095_comb = p70_literal_2043918[p71_array_index_2057061_comb];
  assign p71_array_index_2057096_comb = p70_literal_2043920[p71_array_index_2057062_comb];
  assign p71_res7__930_comb = p71_array_index_2057091_comb ^ p71_array_index_2057092_comb ^ p71_array_index_2057093_comb ^ p71_array_index_2057094_comb ^ p71_array_index_2057095_comb ^ p71_array_index_2057096_comb ^ p71_array_index_2057063_comb ^ p70_literal_2043923[p71_array_index_2057080_comb] ^ p71_array_index_2057065_comb ^ p70_literal_2043920[p71_array_index_2057082_comb] ^ p70_literal_2043918[p71_array_index_2057067_comb] ^ p70_literal_2043916[p71_array_index_2057068_comb] ^ p70_literal_2043914[p71_array_index_2057069_comb] ^ p70_literal_2043912[p71_array_index_2057070_comb] ^ p70_literal_2043910[p71_array_index_2057071_comb] ^ p71_array_index_2057072_comb;
  assign p71_array_index_2057106_comb = p70_literal_2043912[p71_res7__928_comb];
  assign p71_array_index_2057107_comb = p70_literal_2043914[p71_array_index_2057058_comb];
  assign p71_array_index_2057108_comb = p70_literal_2043916[p71_array_index_2057059_comb];
  assign p71_array_index_2057109_comb = p70_literal_2043918[p71_array_index_2057060_comb];
  assign p71_array_index_2057110_comb = p70_literal_2043920[p71_array_index_2057061_comb];
  assign p71_res7__932_comb = p70_literal_2043910[p71_res7__930_comb] ^ p71_array_index_2057106_comb ^ p71_array_index_2057107_comb ^ p71_array_index_2057108_comb ^ p71_array_index_2057109_comb ^ p71_array_index_2057110_comb ^ p71_array_index_2057062_comb ^ p70_literal_2043923[p71_array_index_2057063_comb] ^ p71_array_index_2057080_comb ^ p70_literal_2043920[p71_array_index_2057065_comb] ^ p70_literal_2043918[p71_array_index_2057082_comb] ^ p70_literal_2043916[p71_array_index_2057067_comb] ^ p70_literal_2043914[p71_array_index_2057068_comb] ^ p70_literal_2043912[p71_array_index_2057069_comb] ^ p70_literal_2043910[p71_array_index_2057070_comb] ^ p71_array_index_2057071_comb;

  // Registers for pipe stage 71:
  reg [127:0] p71_encoded;
  reg [127:0] p71_bit_slice_2043893;
  reg [127:0] p71_bit_slice_2044018;
  reg [127:0] p71_k3;
  reg [127:0] p71_k2;
  reg [127:0] p71_k5;
  reg [127:0] p71_k4;
  reg [127:0] p71_k7;
  reg [127:0] p71_k6;
  reg [127:0] p71_xor_2056594;
  reg [127:0] p71_xor_2057042;
  reg [7:0] p71_array_index_2057058;
  reg [7:0] p71_array_index_2057059;
  reg [7:0] p71_array_index_2057060;
  reg [7:0] p71_array_index_2057061;
  reg [7:0] p71_array_index_2057062;
  reg [7:0] p71_array_index_2057063;
  reg [7:0] p71_array_index_2057065;
  reg [7:0] p71_array_index_2057067;
  reg [7:0] p71_array_index_2057068;
  reg [7:0] p71_array_index_2057069;
  reg [7:0] p71_array_index_2057070;
  reg [7:0] p71_array_index_2057074;
  reg [7:0] p71_array_index_2057075;
  reg [7:0] p71_array_index_2057076;
  reg [7:0] p71_array_index_2057077;
  reg [7:0] p71_array_index_2057078;
  reg [7:0] p71_array_index_2057079;
  reg [7:0] p71_array_index_2057080;
  reg [7:0] p71_array_index_2057082;
  reg [7:0] p71_res7__928;
  reg [7:0] p71_array_index_2057091;
  reg [7:0] p71_array_index_2057092;
  reg [7:0] p71_array_index_2057093;
  reg [7:0] p71_array_index_2057094;
  reg [7:0] p71_array_index_2057095;
  reg [7:0] p71_array_index_2057096;
  reg [7:0] p71_res7__930;
  reg [7:0] p71_array_index_2057106;
  reg [7:0] p71_array_index_2057107;
  reg [7:0] p71_array_index_2057108;
  reg [7:0] p71_array_index_2057109;
  reg [7:0] p71_array_index_2057110;
  reg [7:0] p71_res7__932;
  reg [7:0] p72_literal_2043896[256];
  reg [7:0] p72_literal_2043910[256];
  reg [7:0] p72_literal_2043912[256];
  reg [7:0] p72_literal_2043914[256];
  reg [7:0] p72_literal_2043916[256];
  reg [7:0] p72_literal_2043918[256];
  reg [7:0] p72_literal_2043920[256];
  reg [7:0] p72_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p71_encoded <= p70_encoded;
    p71_bit_slice_2043893 <= p70_bit_slice_2043893;
    p71_bit_slice_2044018 <= p70_bit_slice_2044018;
    p71_k3 <= p70_k3;
    p71_k2 <= p70_k2;
    p71_k5 <= p70_k5;
    p71_k4 <= p70_k4;
    p71_k7 <= p70_k7;
    p71_k6 <= p70_k6;
    p71_xor_2056594 <= p70_xor_2056594;
    p71_xor_2057042 <= p71_xor_2057042_comb;
    p71_array_index_2057058 <= p71_array_index_2057058_comb;
    p71_array_index_2057059 <= p71_array_index_2057059_comb;
    p71_array_index_2057060 <= p71_array_index_2057060_comb;
    p71_array_index_2057061 <= p71_array_index_2057061_comb;
    p71_array_index_2057062 <= p71_array_index_2057062_comb;
    p71_array_index_2057063 <= p71_array_index_2057063_comb;
    p71_array_index_2057065 <= p71_array_index_2057065_comb;
    p71_array_index_2057067 <= p71_array_index_2057067_comb;
    p71_array_index_2057068 <= p71_array_index_2057068_comb;
    p71_array_index_2057069 <= p71_array_index_2057069_comb;
    p71_array_index_2057070 <= p71_array_index_2057070_comb;
    p71_array_index_2057074 <= p71_array_index_2057074_comb;
    p71_array_index_2057075 <= p71_array_index_2057075_comb;
    p71_array_index_2057076 <= p71_array_index_2057076_comb;
    p71_array_index_2057077 <= p71_array_index_2057077_comb;
    p71_array_index_2057078 <= p71_array_index_2057078_comb;
    p71_array_index_2057079 <= p71_array_index_2057079_comb;
    p71_array_index_2057080 <= p71_array_index_2057080_comb;
    p71_array_index_2057082 <= p71_array_index_2057082_comb;
    p71_res7__928 <= p71_res7__928_comb;
    p71_array_index_2057091 <= p71_array_index_2057091_comb;
    p71_array_index_2057092 <= p71_array_index_2057092_comb;
    p71_array_index_2057093 <= p71_array_index_2057093_comb;
    p71_array_index_2057094 <= p71_array_index_2057094_comb;
    p71_array_index_2057095 <= p71_array_index_2057095_comb;
    p71_array_index_2057096 <= p71_array_index_2057096_comb;
    p71_res7__930 <= p71_res7__930_comb;
    p71_array_index_2057106 <= p71_array_index_2057106_comb;
    p71_array_index_2057107 <= p71_array_index_2057107_comb;
    p71_array_index_2057108 <= p71_array_index_2057108_comb;
    p71_array_index_2057109 <= p71_array_index_2057109_comb;
    p71_array_index_2057110 <= p71_array_index_2057110_comb;
    p71_res7__932 <= p71_res7__932_comb;
    p72_literal_2043896 <= p71_literal_2043896;
    p72_literal_2043910 <= p71_literal_2043910;
    p72_literal_2043912 <= p71_literal_2043912;
    p72_literal_2043914 <= p71_literal_2043914;
    p72_literal_2043916 <= p71_literal_2043916;
    p72_literal_2043918 <= p71_literal_2043918;
    p72_literal_2043920 <= p71_literal_2043920;
    p72_literal_2043923 <= p71_literal_2043923;
  end

  // ===== Pipe stage 72:
  wire [7:0] p72_array_index_2057224_comb;
  wire [7:0] p72_array_index_2057225_comb;
  wire [7:0] p72_array_index_2057226_comb;
  wire [7:0] p72_array_index_2057227_comb;
  wire [7:0] p72_array_index_2057228_comb;
  wire [7:0] p72_res7__934_comb;
  wire [7:0] p72_array_index_2057239_comb;
  wire [7:0] p72_array_index_2057240_comb;
  wire [7:0] p72_array_index_2057241_comb;
  wire [7:0] p72_array_index_2057242_comb;
  wire [7:0] p72_res7__936_comb;
  wire [7:0] p72_array_index_2057252_comb;
  wire [7:0] p72_array_index_2057253_comb;
  wire [7:0] p72_array_index_2057254_comb;
  wire [7:0] p72_array_index_2057255_comb;
  wire [7:0] p72_res7__938_comb;
  wire [7:0] p72_array_index_2057266_comb;
  wire [7:0] p72_array_index_2057267_comb;
  wire [7:0] p72_array_index_2057268_comb;
  wire [7:0] p72_res7__940_comb;
  wire [7:0] p72_array_index_2057278_comb;
  wire [7:0] p72_array_index_2057279_comb;
  wire [7:0] p72_array_index_2057280_comb;
  wire [7:0] p72_res7__942_comb;
  wire [7:0] p72_array_index_2057291_comb;
  wire [7:0] p72_array_index_2057292_comb;
  wire [7:0] p72_res7__944_comb;
  wire [7:0] p72_array_index_2057302_comb;
  wire [7:0] p72_array_index_2057303_comb;
  wire [7:0] p72_res7__946_comb;
  assign p72_array_index_2057224_comb = p71_literal_2043912[p71_res7__930];
  assign p72_array_index_2057225_comb = p71_literal_2043914[p71_res7__928];
  assign p72_array_index_2057226_comb = p71_literal_2043916[p71_array_index_2057058];
  assign p72_array_index_2057227_comb = p71_literal_2043918[p71_array_index_2057059];
  assign p72_array_index_2057228_comb = p71_literal_2043920[p71_array_index_2057060];
  assign p72_res7__934_comb = p71_literal_2043910[p71_res7__932] ^ p72_array_index_2057224_comb ^ p72_array_index_2057225_comb ^ p72_array_index_2057226_comb ^ p72_array_index_2057227_comb ^ p72_array_index_2057228_comb ^ p71_array_index_2057061 ^ p71_literal_2043923[p71_array_index_2057062] ^ p71_array_index_2057063 ^ p71_literal_2043920[p71_array_index_2057080] ^ p71_literal_2043918[p71_array_index_2057065] ^ p71_literal_2043916[p71_array_index_2057082] ^ p71_literal_2043914[p71_array_index_2057067] ^ p71_literal_2043912[p71_array_index_2057068] ^ p71_literal_2043910[p71_array_index_2057069] ^ p71_array_index_2057070;
  assign p72_array_index_2057239_comb = p71_literal_2043914[p71_res7__930];
  assign p72_array_index_2057240_comb = p71_literal_2043916[p71_res7__928];
  assign p72_array_index_2057241_comb = p71_literal_2043918[p71_array_index_2057058];
  assign p72_array_index_2057242_comb = p71_literal_2043920[p71_array_index_2057059];
  assign p72_res7__936_comb = p71_literal_2043910[p72_res7__934_comb] ^ p71_literal_2043912[p71_res7__932] ^ p72_array_index_2057239_comb ^ p72_array_index_2057240_comb ^ p72_array_index_2057241_comb ^ p72_array_index_2057242_comb ^ p71_array_index_2057060 ^ p71_literal_2043923[p71_array_index_2057061] ^ p71_array_index_2057062 ^ p71_array_index_2057079 ^ p71_literal_2043918[p71_array_index_2057080] ^ p71_literal_2043916[p71_array_index_2057065] ^ p71_literal_2043914[p71_array_index_2057082] ^ p71_literal_2043912[p71_array_index_2057067] ^ p71_literal_2043910[p71_array_index_2057068] ^ p71_array_index_2057069;
  assign p72_array_index_2057252_comb = p71_literal_2043914[p71_res7__932];
  assign p72_array_index_2057253_comb = p71_literal_2043916[p71_res7__930];
  assign p72_array_index_2057254_comb = p71_literal_2043918[p71_res7__928];
  assign p72_array_index_2057255_comb = p71_literal_2043920[p71_array_index_2057058];
  assign p72_res7__938_comb = p71_literal_2043910[p72_res7__936_comb] ^ p71_literal_2043912[p72_res7__934_comb] ^ p72_array_index_2057252_comb ^ p72_array_index_2057253_comb ^ p72_array_index_2057254_comb ^ p72_array_index_2057255_comb ^ p71_array_index_2057059 ^ p71_literal_2043923[p71_array_index_2057060] ^ p71_array_index_2057061 ^ p71_array_index_2057096 ^ p71_literal_2043918[p71_array_index_2057063] ^ p71_literal_2043916[p71_array_index_2057080] ^ p71_literal_2043914[p71_array_index_2057065] ^ p71_literal_2043912[p71_array_index_2057082] ^ p71_literal_2043910[p71_array_index_2057067] ^ p71_array_index_2057068;
  assign p72_array_index_2057266_comb = p71_literal_2043916[p71_res7__932];
  assign p72_array_index_2057267_comb = p71_literal_2043918[p71_res7__930];
  assign p72_array_index_2057268_comb = p71_literal_2043920[p71_res7__928];
  assign p72_res7__940_comb = p71_literal_2043910[p72_res7__938_comb] ^ p71_literal_2043912[p72_res7__936_comb] ^ p71_literal_2043914[p72_res7__934_comb] ^ p72_array_index_2057266_comb ^ p72_array_index_2057267_comb ^ p72_array_index_2057268_comb ^ p71_array_index_2057058 ^ p71_literal_2043923[p71_array_index_2057059] ^ p71_array_index_2057060 ^ p71_array_index_2057110 ^ p71_array_index_2057078 ^ p71_literal_2043916[p71_array_index_2057063] ^ p71_literal_2043914[p71_array_index_2057080] ^ p71_literal_2043912[p71_array_index_2057065] ^ p71_literal_2043910[p71_array_index_2057082] ^ p71_array_index_2057067;
  assign p72_array_index_2057278_comb = p71_literal_2043916[p72_res7__934_comb];
  assign p72_array_index_2057279_comb = p71_literal_2043918[p71_res7__932];
  assign p72_array_index_2057280_comb = p71_literal_2043920[p71_res7__930];
  assign p72_res7__942_comb = p71_literal_2043910[p72_res7__940_comb] ^ p71_literal_2043912[p72_res7__938_comb] ^ p71_literal_2043914[p72_res7__936_comb] ^ p72_array_index_2057278_comb ^ p72_array_index_2057279_comb ^ p72_array_index_2057280_comb ^ p71_res7__928 ^ p71_literal_2043923[p71_array_index_2057058] ^ p71_array_index_2057059 ^ p72_array_index_2057228_comb ^ p71_array_index_2057095 ^ p71_literal_2043916[p71_array_index_2057062] ^ p71_literal_2043914[p71_array_index_2057063] ^ p71_literal_2043912[p71_array_index_2057080] ^ p71_literal_2043910[p71_array_index_2057065] ^ p71_array_index_2057082;
  assign p72_array_index_2057291_comb = p71_literal_2043918[p72_res7__934_comb];
  assign p72_array_index_2057292_comb = p71_literal_2043920[p71_res7__932];
  assign p72_res7__944_comb = p71_literal_2043910[p72_res7__942_comb] ^ p71_literal_2043912[p72_res7__940_comb] ^ p71_literal_2043914[p72_res7__938_comb] ^ p71_literal_2043916[p72_res7__936_comb] ^ p72_array_index_2057291_comb ^ p72_array_index_2057292_comb ^ p71_res7__930 ^ p71_literal_2043923[p71_res7__928] ^ p71_array_index_2057058 ^ p72_array_index_2057242_comb ^ p71_array_index_2057109 ^ p71_array_index_2057077 ^ p71_literal_2043914[p71_array_index_2057062] ^ p71_literal_2043912[p71_array_index_2057063] ^ p71_literal_2043910[p71_array_index_2057080] ^ p71_array_index_2057065;
  assign p72_array_index_2057302_comb = p71_literal_2043918[p72_res7__936_comb];
  assign p72_array_index_2057303_comb = p71_literal_2043920[p72_res7__934_comb];
  assign p72_res7__946_comb = p71_literal_2043910[p72_res7__944_comb] ^ p71_literal_2043912[p72_res7__942_comb] ^ p71_literal_2043914[p72_res7__940_comb] ^ p71_literal_2043916[p72_res7__938_comb] ^ p72_array_index_2057302_comb ^ p72_array_index_2057303_comb ^ p71_res7__932 ^ p71_literal_2043923[p71_res7__930] ^ p71_res7__928 ^ p72_array_index_2057255_comb ^ p72_array_index_2057227_comb ^ p71_array_index_2057094 ^ p71_literal_2043914[p71_array_index_2057061] ^ p71_literal_2043912[p71_array_index_2057062] ^ p71_literal_2043910[p71_array_index_2057063] ^ p71_array_index_2057080;

  // Registers for pipe stage 72:
  reg [127:0] p72_encoded;
  reg [127:0] p72_bit_slice_2043893;
  reg [127:0] p72_bit_slice_2044018;
  reg [127:0] p72_k3;
  reg [127:0] p72_k2;
  reg [127:0] p72_k5;
  reg [127:0] p72_k4;
  reg [127:0] p72_k7;
  reg [127:0] p72_k6;
  reg [127:0] p72_xor_2056594;
  reg [127:0] p72_xor_2057042;
  reg [7:0] p72_array_index_2057058;
  reg [7:0] p72_array_index_2057059;
  reg [7:0] p72_array_index_2057060;
  reg [7:0] p72_array_index_2057061;
  reg [7:0] p72_array_index_2057062;
  reg [7:0] p72_array_index_2057063;
  reg [7:0] p72_array_index_2057074;
  reg [7:0] p72_array_index_2057075;
  reg [7:0] p72_array_index_2057076;
  reg [7:0] p72_res7__928;
  reg [7:0] p72_array_index_2057091;
  reg [7:0] p72_array_index_2057092;
  reg [7:0] p72_array_index_2057093;
  reg [7:0] p72_res7__930;
  reg [7:0] p72_array_index_2057106;
  reg [7:0] p72_array_index_2057107;
  reg [7:0] p72_array_index_2057108;
  reg [7:0] p72_res7__932;
  reg [7:0] p72_array_index_2057224;
  reg [7:0] p72_array_index_2057225;
  reg [7:0] p72_array_index_2057226;
  reg [7:0] p72_res7__934;
  reg [7:0] p72_array_index_2057239;
  reg [7:0] p72_array_index_2057240;
  reg [7:0] p72_array_index_2057241;
  reg [7:0] p72_res7__936;
  reg [7:0] p72_array_index_2057252;
  reg [7:0] p72_array_index_2057253;
  reg [7:0] p72_array_index_2057254;
  reg [7:0] p72_res7__938;
  reg [7:0] p72_array_index_2057266;
  reg [7:0] p72_array_index_2057267;
  reg [7:0] p72_array_index_2057268;
  reg [7:0] p72_res7__940;
  reg [7:0] p72_array_index_2057278;
  reg [7:0] p72_array_index_2057279;
  reg [7:0] p72_array_index_2057280;
  reg [7:0] p72_res7__942;
  reg [7:0] p72_array_index_2057291;
  reg [7:0] p72_array_index_2057292;
  reg [7:0] p72_res7__944;
  reg [7:0] p72_array_index_2057302;
  reg [7:0] p72_array_index_2057303;
  reg [7:0] p72_res7__946;
  reg [7:0] p73_literal_2043896[256];
  reg [7:0] p73_literal_2043910[256];
  reg [7:0] p73_literal_2043912[256];
  reg [7:0] p73_literal_2043914[256];
  reg [7:0] p73_literal_2043916[256];
  reg [7:0] p73_literal_2043918[256];
  reg [7:0] p73_literal_2043920[256];
  reg [7:0] p73_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p72_encoded <= p71_encoded;
    p72_bit_slice_2043893 <= p71_bit_slice_2043893;
    p72_bit_slice_2044018 <= p71_bit_slice_2044018;
    p72_k3 <= p71_k3;
    p72_k2 <= p71_k2;
    p72_k5 <= p71_k5;
    p72_k4 <= p71_k4;
    p72_k7 <= p71_k7;
    p72_k6 <= p71_k6;
    p72_xor_2056594 <= p71_xor_2056594;
    p72_xor_2057042 <= p71_xor_2057042;
    p72_array_index_2057058 <= p71_array_index_2057058;
    p72_array_index_2057059 <= p71_array_index_2057059;
    p72_array_index_2057060 <= p71_array_index_2057060;
    p72_array_index_2057061 <= p71_array_index_2057061;
    p72_array_index_2057062 <= p71_array_index_2057062;
    p72_array_index_2057063 <= p71_array_index_2057063;
    p72_array_index_2057074 <= p71_array_index_2057074;
    p72_array_index_2057075 <= p71_array_index_2057075;
    p72_array_index_2057076 <= p71_array_index_2057076;
    p72_res7__928 <= p71_res7__928;
    p72_array_index_2057091 <= p71_array_index_2057091;
    p72_array_index_2057092 <= p71_array_index_2057092;
    p72_array_index_2057093 <= p71_array_index_2057093;
    p72_res7__930 <= p71_res7__930;
    p72_array_index_2057106 <= p71_array_index_2057106;
    p72_array_index_2057107 <= p71_array_index_2057107;
    p72_array_index_2057108 <= p71_array_index_2057108;
    p72_res7__932 <= p71_res7__932;
    p72_array_index_2057224 <= p72_array_index_2057224_comb;
    p72_array_index_2057225 <= p72_array_index_2057225_comb;
    p72_array_index_2057226 <= p72_array_index_2057226_comb;
    p72_res7__934 <= p72_res7__934_comb;
    p72_array_index_2057239 <= p72_array_index_2057239_comb;
    p72_array_index_2057240 <= p72_array_index_2057240_comb;
    p72_array_index_2057241 <= p72_array_index_2057241_comb;
    p72_res7__936 <= p72_res7__936_comb;
    p72_array_index_2057252 <= p72_array_index_2057252_comb;
    p72_array_index_2057253 <= p72_array_index_2057253_comb;
    p72_array_index_2057254 <= p72_array_index_2057254_comb;
    p72_res7__938 <= p72_res7__938_comb;
    p72_array_index_2057266 <= p72_array_index_2057266_comb;
    p72_array_index_2057267 <= p72_array_index_2057267_comb;
    p72_array_index_2057268 <= p72_array_index_2057268_comb;
    p72_res7__940 <= p72_res7__940_comb;
    p72_array_index_2057278 <= p72_array_index_2057278_comb;
    p72_array_index_2057279 <= p72_array_index_2057279_comb;
    p72_array_index_2057280 <= p72_array_index_2057280_comb;
    p72_res7__942 <= p72_res7__942_comb;
    p72_array_index_2057291 <= p72_array_index_2057291_comb;
    p72_array_index_2057292 <= p72_array_index_2057292_comb;
    p72_res7__944 <= p72_res7__944_comb;
    p72_array_index_2057302 <= p72_array_index_2057302_comb;
    p72_array_index_2057303 <= p72_array_index_2057303_comb;
    p72_res7__946 <= p72_res7__946_comb;
    p73_literal_2043896 <= p72_literal_2043896;
    p73_literal_2043910 <= p72_literal_2043910;
    p73_literal_2043912 <= p72_literal_2043912;
    p73_literal_2043914 <= p72_literal_2043914;
    p73_literal_2043916 <= p72_literal_2043916;
    p73_literal_2043918 <= p72_literal_2043918;
    p73_literal_2043920 <= p72_literal_2043920;
    p73_literal_2043923 <= p72_literal_2043923;
  end

  // ===== Pipe stage 73:
  wire [7:0] p73_array_index_2057440_comb;
  wire [7:0] p73_res7__948_comb;
  wire [7:0] p73_array_index_2057450_comb;
  wire [7:0] p73_res7__950_comb;
  wire [7:0] p73_res7__952_comb;
  wire [7:0] p73_res7__954_comb;
  wire [7:0] p73_res7__956_comb;
  wire [7:0] p73_res7__958_comb;
  wire [127:0] p73_res__29_comb;
  wire [127:0] p73_xor_2057490_comb;
  wire [127:0] p73_addedKey__62_comb;
  wire [7:0] p73_array_index_2057506_comb;
  wire [7:0] p73_array_index_2057507_comb;
  wire [7:0] p73_array_index_2057508_comb;
  wire [7:0] p73_array_index_2057509_comb;
  wire [7:0] p73_array_index_2057510_comb;
  wire [7:0] p73_array_index_2057511_comb;
  wire [7:0] p73_array_index_2057513_comb;
  wire [7:0] p73_array_index_2057515_comb;
  wire [7:0] p73_array_index_2057516_comb;
  wire [7:0] p73_array_index_2057517_comb;
  wire [7:0] p73_array_index_2057518_comb;
  wire [7:0] p73_array_index_2057519_comb;
  wire [7:0] p73_array_index_2057520_comb;
  wire [7:0] p73_array_index_2057522_comb;
  wire [7:0] p73_array_index_2057523_comb;
  wire [7:0] p73_array_index_2057524_comb;
  assign p73_array_index_2057440_comb = p72_literal_2043920[p72_res7__936];
  assign p73_res7__948_comb = p72_literal_2043910[p72_res7__946] ^ p72_literal_2043912[p72_res7__944] ^ p72_literal_2043914[p72_res7__942] ^ p72_literal_2043916[p72_res7__940] ^ p72_literal_2043918[p72_res7__938] ^ p73_array_index_2057440_comb ^ p72_res7__934 ^ p72_literal_2043923[p72_res7__932] ^ p72_res7__930 ^ p72_array_index_2057268 ^ p72_array_index_2057241 ^ p72_array_index_2057108 ^ p72_array_index_2057076 ^ p72_literal_2043912[p72_array_index_2057061] ^ p72_literal_2043910[p72_array_index_2057062] ^ p72_array_index_2057063;
  assign p73_array_index_2057450_comb = p72_literal_2043920[p72_res7__938];
  assign p73_res7__950_comb = p72_literal_2043910[p73_res7__948_comb] ^ p72_literal_2043912[p72_res7__946] ^ p72_literal_2043914[p72_res7__944] ^ p72_literal_2043916[p72_res7__942] ^ p72_literal_2043918[p72_res7__940] ^ p73_array_index_2057450_comb ^ p72_res7__936 ^ p72_literal_2043923[p72_res7__934] ^ p72_res7__932 ^ p72_array_index_2057280 ^ p72_array_index_2057254 ^ p72_array_index_2057226 ^ p72_array_index_2057093 ^ p72_literal_2043912[p72_array_index_2057060] ^ p72_literal_2043910[p72_array_index_2057061] ^ p72_array_index_2057062;
  assign p73_res7__952_comb = p72_literal_2043910[p73_res7__950_comb] ^ p72_literal_2043912[p73_res7__948_comb] ^ p72_literal_2043914[p72_res7__946] ^ p72_literal_2043916[p72_res7__944] ^ p72_literal_2043918[p72_res7__942] ^ p72_literal_2043920[p72_res7__940] ^ p72_res7__938 ^ p72_literal_2043923[p72_res7__936] ^ p72_res7__934 ^ p72_array_index_2057292 ^ p72_array_index_2057267 ^ p72_array_index_2057240 ^ p72_array_index_2057107 ^ p72_array_index_2057075 ^ p72_literal_2043910[p72_array_index_2057060] ^ p72_array_index_2057061;
  assign p73_res7__954_comb = p72_literal_2043910[p73_res7__952_comb] ^ p72_literal_2043912[p73_res7__950_comb] ^ p72_literal_2043914[p73_res7__948_comb] ^ p72_literal_2043916[p72_res7__946] ^ p72_literal_2043918[p72_res7__944] ^ p72_literal_2043920[p72_res7__942] ^ p72_res7__940 ^ p72_literal_2043923[p72_res7__938] ^ p72_res7__936 ^ p72_array_index_2057303 ^ p72_array_index_2057279 ^ p72_array_index_2057253 ^ p72_array_index_2057225 ^ p72_array_index_2057092 ^ p72_literal_2043910[p72_array_index_2057059] ^ p72_array_index_2057060;
  assign p73_res7__956_comb = p72_literal_2043910[p73_res7__954_comb] ^ p72_literal_2043912[p73_res7__952_comb] ^ p72_literal_2043914[p73_res7__950_comb] ^ p72_literal_2043916[p73_res7__948_comb] ^ p72_literal_2043918[p72_res7__946] ^ p72_literal_2043920[p72_res7__944] ^ p72_res7__942 ^ p72_literal_2043923[p72_res7__940] ^ p72_res7__938 ^ p73_array_index_2057440_comb ^ p72_array_index_2057291 ^ p72_array_index_2057266 ^ p72_array_index_2057239 ^ p72_array_index_2057106 ^ p72_array_index_2057074 ^ p72_array_index_2057059;
  assign p73_res7__958_comb = p72_literal_2043910[p73_res7__956_comb] ^ p72_literal_2043912[p73_res7__954_comb] ^ p72_literal_2043914[p73_res7__952_comb] ^ p72_literal_2043916[p73_res7__950_comb] ^ p72_literal_2043918[p73_res7__948_comb] ^ p72_literal_2043920[p72_res7__946] ^ p72_res7__944 ^ p72_literal_2043923[p72_res7__942] ^ p72_res7__940 ^ p73_array_index_2057450_comb ^ p72_array_index_2057302 ^ p72_array_index_2057278 ^ p72_array_index_2057252 ^ p72_array_index_2057224 ^ p72_array_index_2057091 ^ p72_array_index_2057058;
  assign p73_res__29_comb = {p73_res7__958_comb, p73_res7__956_comb, p73_res7__954_comb, p73_res7__952_comb, p73_res7__950_comb, p73_res7__948_comb, p72_res7__946, p72_res7__944, p72_res7__942, p72_res7__940, p72_res7__938, p72_res7__936, p72_res7__934, p72_res7__932, p72_res7__930, p72_res7__928};
  assign p73_xor_2057490_comb = p73_res__29_comb ^ p72_xor_2056594;
  assign p73_addedKey__62_comb = p73_xor_2057490_comb ^ 128'h1003_dba7_2e34_5ff6_643b_9533_3f27_141f;
  assign p73_array_index_2057506_comb = p72_literal_2043896[p73_addedKey__62_comb[127:120]];
  assign p73_array_index_2057507_comb = p72_literal_2043896[p73_addedKey__62_comb[119:112]];
  assign p73_array_index_2057508_comb = p72_literal_2043896[p73_addedKey__62_comb[111:104]];
  assign p73_array_index_2057509_comb = p72_literal_2043896[p73_addedKey__62_comb[103:96]];
  assign p73_array_index_2057510_comb = p72_literal_2043896[p73_addedKey__62_comb[95:88]];
  assign p73_array_index_2057511_comb = p72_literal_2043896[p73_addedKey__62_comb[87:80]];
  assign p73_array_index_2057513_comb = p72_literal_2043896[p73_addedKey__62_comb[71:64]];
  assign p73_array_index_2057515_comb = p72_literal_2043896[p73_addedKey__62_comb[55:48]];
  assign p73_array_index_2057516_comb = p72_literal_2043896[p73_addedKey__62_comb[47:40]];
  assign p73_array_index_2057517_comb = p72_literal_2043896[p73_addedKey__62_comb[39:32]];
  assign p73_array_index_2057518_comb = p72_literal_2043896[p73_addedKey__62_comb[31:24]];
  assign p73_array_index_2057519_comb = p72_literal_2043896[p73_addedKey__62_comb[23:16]];
  assign p73_array_index_2057520_comb = p72_literal_2043896[p73_addedKey__62_comb[15:8]];
  assign p73_array_index_2057522_comb = p72_literal_2043896[p73_addedKey__62_comb[79:72]];
  assign p73_array_index_2057523_comb = p72_literal_2043896[p73_addedKey__62_comb[63:56]];
  assign p73_array_index_2057524_comb = p72_literal_2043896[p73_addedKey__62_comb[7:0]];

  // Registers for pipe stage 73:
  reg [127:0] p73_encoded;
  reg [127:0] p73_bit_slice_2043893;
  reg [127:0] p73_bit_slice_2044018;
  reg [127:0] p73_k3;
  reg [127:0] p73_k2;
  reg [127:0] p73_k5;
  reg [127:0] p73_k4;
  reg [127:0] p73_k7;
  reg [127:0] p73_k6;
  reg [127:0] p73_xor_2057042;
  reg [127:0] p73_xor_2057490;
  reg [7:0] p73_array_index_2057506;
  reg [7:0] p73_array_index_2057507;
  reg [7:0] p73_array_index_2057508;
  reg [7:0] p73_array_index_2057509;
  reg [7:0] p73_array_index_2057510;
  reg [7:0] p73_array_index_2057511;
  reg [7:0] p73_array_index_2057513;
  reg [7:0] p73_array_index_2057515;
  reg [7:0] p73_array_index_2057516;
  reg [7:0] p73_array_index_2057517;
  reg [7:0] p73_array_index_2057518;
  reg [7:0] p73_array_index_2057519;
  reg [7:0] p73_array_index_2057520;
  reg [7:0] p73_array_index_2057522;
  reg [7:0] p73_array_index_2057523;
  reg [7:0] p73_array_index_2057524;
  reg [7:0] p74_literal_2043896[256];
  reg [7:0] p74_literal_2043910[256];
  reg [7:0] p74_literal_2043912[256];
  reg [7:0] p74_literal_2043914[256];
  reg [7:0] p74_literal_2043916[256];
  reg [7:0] p74_literal_2043918[256];
  reg [7:0] p74_literal_2043920[256];
  reg [7:0] p74_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p73_encoded <= p72_encoded;
    p73_bit_slice_2043893 <= p72_bit_slice_2043893;
    p73_bit_slice_2044018 <= p72_bit_slice_2044018;
    p73_k3 <= p72_k3;
    p73_k2 <= p72_k2;
    p73_k5 <= p72_k5;
    p73_k4 <= p72_k4;
    p73_k7 <= p72_k7;
    p73_k6 <= p72_k6;
    p73_xor_2057042 <= p72_xor_2057042;
    p73_xor_2057490 <= p73_xor_2057490_comb;
    p73_array_index_2057506 <= p73_array_index_2057506_comb;
    p73_array_index_2057507 <= p73_array_index_2057507_comb;
    p73_array_index_2057508 <= p73_array_index_2057508_comb;
    p73_array_index_2057509 <= p73_array_index_2057509_comb;
    p73_array_index_2057510 <= p73_array_index_2057510_comb;
    p73_array_index_2057511 <= p73_array_index_2057511_comb;
    p73_array_index_2057513 <= p73_array_index_2057513_comb;
    p73_array_index_2057515 <= p73_array_index_2057515_comb;
    p73_array_index_2057516 <= p73_array_index_2057516_comb;
    p73_array_index_2057517 <= p73_array_index_2057517_comb;
    p73_array_index_2057518 <= p73_array_index_2057518_comb;
    p73_array_index_2057519 <= p73_array_index_2057519_comb;
    p73_array_index_2057520 <= p73_array_index_2057520_comb;
    p73_array_index_2057522 <= p73_array_index_2057522_comb;
    p73_array_index_2057523 <= p73_array_index_2057523_comb;
    p73_array_index_2057524 <= p73_array_index_2057524_comb;
    p74_literal_2043896 <= p73_literal_2043896;
    p74_literal_2043910 <= p73_literal_2043910;
    p74_literal_2043912 <= p73_literal_2043912;
    p74_literal_2043914 <= p73_literal_2043914;
    p74_literal_2043916 <= p73_literal_2043916;
    p74_literal_2043918 <= p73_literal_2043918;
    p74_literal_2043920 <= p73_literal_2043920;
    p74_literal_2043923 <= p73_literal_2043923;
  end

  // ===== Pipe stage 74:
  wire [7:0] p74_array_index_2057595_comb;
  wire [7:0] p74_array_index_2057596_comb;
  wire [7:0] p74_array_index_2057597_comb;
  wire [7:0] p74_array_index_2057598_comb;
  wire [7:0] p74_array_index_2057599_comb;
  wire [7:0] p74_array_index_2057600_comb;
  wire [7:0] p74_res7__960_comb;
  wire [7:0] p74_array_index_2057609_comb;
  wire [7:0] p74_array_index_2057610_comb;
  wire [7:0] p74_array_index_2057611_comb;
  wire [7:0] p74_array_index_2057612_comb;
  wire [7:0] p74_array_index_2057613_comb;
  wire [7:0] p74_array_index_2057614_comb;
  wire [7:0] p74_res7__962_comb;
  wire [7:0] p74_array_index_2057624_comb;
  wire [7:0] p74_array_index_2057625_comb;
  wire [7:0] p74_array_index_2057626_comb;
  wire [7:0] p74_array_index_2057627_comb;
  wire [7:0] p74_array_index_2057628_comb;
  wire [7:0] p74_res7__964_comb;
  wire [7:0] p74_array_index_2057638_comb;
  wire [7:0] p74_array_index_2057639_comb;
  wire [7:0] p74_array_index_2057640_comb;
  wire [7:0] p74_array_index_2057641_comb;
  wire [7:0] p74_array_index_2057642_comb;
  wire [7:0] p74_res7__966_comb;
  wire [7:0] p74_array_index_2057653_comb;
  wire [7:0] p74_array_index_2057654_comb;
  wire [7:0] p74_array_index_2057655_comb;
  wire [7:0] p74_array_index_2057656_comb;
  wire [7:0] p74_res7__968_comb;
  wire [7:0] p74_array_index_2057666_comb;
  wire [7:0] p74_array_index_2057667_comb;
  wire [7:0] p74_array_index_2057668_comb;
  wire [7:0] p74_array_index_2057669_comb;
  wire [7:0] p74_res7__970_comb;
  wire [7:0] p74_array_index_2057680_comb;
  wire [7:0] p74_array_index_2057681_comb;
  wire [7:0] p74_array_index_2057682_comb;
  wire [7:0] p74_res7__972_comb;
  assign p74_array_index_2057595_comb = p73_literal_2043910[p73_array_index_2057506];
  assign p74_array_index_2057596_comb = p73_literal_2043912[p73_array_index_2057507];
  assign p74_array_index_2057597_comb = p73_literal_2043914[p73_array_index_2057508];
  assign p74_array_index_2057598_comb = p73_literal_2043916[p73_array_index_2057509];
  assign p74_array_index_2057599_comb = p73_literal_2043918[p73_array_index_2057510];
  assign p74_array_index_2057600_comb = p73_literal_2043920[p73_array_index_2057511];
  assign p74_res7__960_comb = p74_array_index_2057595_comb ^ p74_array_index_2057596_comb ^ p74_array_index_2057597_comb ^ p74_array_index_2057598_comb ^ p74_array_index_2057599_comb ^ p74_array_index_2057600_comb ^ p73_array_index_2057522 ^ p73_literal_2043923[p73_array_index_2057513] ^ p73_array_index_2057523 ^ p73_literal_2043920[p73_array_index_2057515] ^ p73_literal_2043918[p73_array_index_2057516] ^ p73_literal_2043916[p73_array_index_2057517] ^ p73_literal_2043914[p73_array_index_2057518] ^ p73_literal_2043912[p73_array_index_2057519] ^ p73_literal_2043910[p73_array_index_2057520] ^ p73_array_index_2057524;
  assign p74_array_index_2057609_comb = p73_literal_2043910[p74_res7__960_comb];
  assign p74_array_index_2057610_comb = p73_literal_2043912[p73_array_index_2057506];
  assign p74_array_index_2057611_comb = p73_literal_2043914[p73_array_index_2057507];
  assign p74_array_index_2057612_comb = p73_literal_2043916[p73_array_index_2057508];
  assign p74_array_index_2057613_comb = p73_literal_2043918[p73_array_index_2057509];
  assign p74_array_index_2057614_comb = p73_literal_2043920[p73_array_index_2057510];
  assign p74_res7__962_comb = p74_array_index_2057609_comb ^ p74_array_index_2057610_comb ^ p74_array_index_2057611_comb ^ p74_array_index_2057612_comb ^ p74_array_index_2057613_comb ^ p74_array_index_2057614_comb ^ p73_array_index_2057511 ^ p73_literal_2043923[p73_array_index_2057522] ^ p73_array_index_2057513 ^ p73_literal_2043920[p73_array_index_2057523] ^ p73_literal_2043918[p73_array_index_2057515] ^ p73_literal_2043916[p73_array_index_2057516] ^ p73_literal_2043914[p73_array_index_2057517] ^ p73_literal_2043912[p73_array_index_2057518] ^ p73_literal_2043910[p73_array_index_2057519] ^ p73_array_index_2057520;
  assign p74_array_index_2057624_comb = p73_literal_2043912[p74_res7__960_comb];
  assign p74_array_index_2057625_comb = p73_literal_2043914[p73_array_index_2057506];
  assign p74_array_index_2057626_comb = p73_literal_2043916[p73_array_index_2057507];
  assign p74_array_index_2057627_comb = p73_literal_2043918[p73_array_index_2057508];
  assign p74_array_index_2057628_comb = p73_literal_2043920[p73_array_index_2057509];
  assign p74_res7__964_comb = p73_literal_2043910[p74_res7__962_comb] ^ p74_array_index_2057624_comb ^ p74_array_index_2057625_comb ^ p74_array_index_2057626_comb ^ p74_array_index_2057627_comb ^ p74_array_index_2057628_comb ^ p73_array_index_2057510 ^ p73_literal_2043923[p73_array_index_2057511] ^ p73_array_index_2057522 ^ p73_literal_2043920[p73_array_index_2057513] ^ p73_literal_2043918[p73_array_index_2057523] ^ p73_literal_2043916[p73_array_index_2057515] ^ p73_literal_2043914[p73_array_index_2057516] ^ p73_literal_2043912[p73_array_index_2057517] ^ p73_literal_2043910[p73_array_index_2057518] ^ p73_array_index_2057519;
  assign p74_array_index_2057638_comb = p73_literal_2043912[p74_res7__962_comb];
  assign p74_array_index_2057639_comb = p73_literal_2043914[p74_res7__960_comb];
  assign p74_array_index_2057640_comb = p73_literal_2043916[p73_array_index_2057506];
  assign p74_array_index_2057641_comb = p73_literal_2043918[p73_array_index_2057507];
  assign p74_array_index_2057642_comb = p73_literal_2043920[p73_array_index_2057508];
  assign p74_res7__966_comb = p73_literal_2043910[p74_res7__964_comb] ^ p74_array_index_2057638_comb ^ p74_array_index_2057639_comb ^ p74_array_index_2057640_comb ^ p74_array_index_2057641_comb ^ p74_array_index_2057642_comb ^ p73_array_index_2057509 ^ p73_literal_2043923[p73_array_index_2057510] ^ p73_array_index_2057511 ^ p73_literal_2043920[p73_array_index_2057522] ^ p73_literal_2043918[p73_array_index_2057513] ^ p73_literal_2043916[p73_array_index_2057523] ^ p73_literal_2043914[p73_array_index_2057515] ^ p73_literal_2043912[p73_array_index_2057516] ^ p73_literal_2043910[p73_array_index_2057517] ^ p73_array_index_2057518;
  assign p74_array_index_2057653_comb = p73_literal_2043914[p74_res7__962_comb];
  assign p74_array_index_2057654_comb = p73_literal_2043916[p74_res7__960_comb];
  assign p74_array_index_2057655_comb = p73_literal_2043918[p73_array_index_2057506];
  assign p74_array_index_2057656_comb = p73_literal_2043920[p73_array_index_2057507];
  assign p74_res7__968_comb = p73_literal_2043910[p74_res7__966_comb] ^ p73_literal_2043912[p74_res7__964_comb] ^ p74_array_index_2057653_comb ^ p74_array_index_2057654_comb ^ p74_array_index_2057655_comb ^ p74_array_index_2057656_comb ^ p73_array_index_2057508 ^ p73_literal_2043923[p73_array_index_2057509] ^ p73_array_index_2057510 ^ p74_array_index_2057600_comb ^ p73_literal_2043918[p73_array_index_2057522] ^ p73_literal_2043916[p73_array_index_2057513] ^ p73_literal_2043914[p73_array_index_2057523] ^ p73_literal_2043912[p73_array_index_2057515] ^ p73_literal_2043910[p73_array_index_2057516] ^ p73_array_index_2057517;
  assign p74_array_index_2057666_comb = p73_literal_2043914[p74_res7__964_comb];
  assign p74_array_index_2057667_comb = p73_literal_2043916[p74_res7__962_comb];
  assign p74_array_index_2057668_comb = p73_literal_2043918[p74_res7__960_comb];
  assign p74_array_index_2057669_comb = p73_literal_2043920[p73_array_index_2057506];
  assign p74_res7__970_comb = p73_literal_2043910[p74_res7__968_comb] ^ p73_literal_2043912[p74_res7__966_comb] ^ p74_array_index_2057666_comb ^ p74_array_index_2057667_comb ^ p74_array_index_2057668_comb ^ p74_array_index_2057669_comb ^ p73_array_index_2057507 ^ p73_literal_2043923[p73_array_index_2057508] ^ p73_array_index_2057509 ^ p74_array_index_2057614_comb ^ p73_literal_2043918[p73_array_index_2057511] ^ p73_literal_2043916[p73_array_index_2057522] ^ p73_literal_2043914[p73_array_index_2057513] ^ p73_literal_2043912[p73_array_index_2057523] ^ p73_literal_2043910[p73_array_index_2057515] ^ p73_array_index_2057516;
  assign p74_array_index_2057680_comb = p73_literal_2043916[p74_res7__964_comb];
  assign p74_array_index_2057681_comb = p73_literal_2043918[p74_res7__962_comb];
  assign p74_array_index_2057682_comb = p73_literal_2043920[p74_res7__960_comb];
  assign p74_res7__972_comb = p73_literal_2043910[p74_res7__970_comb] ^ p73_literal_2043912[p74_res7__968_comb] ^ p73_literal_2043914[p74_res7__966_comb] ^ p74_array_index_2057680_comb ^ p74_array_index_2057681_comb ^ p74_array_index_2057682_comb ^ p73_array_index_2057506 ^ p73_literal_2043923[p73_array_index_2057507] ^ p73_array_index_2057508 ^ p74_array_index_2057628_comb ^ p74_array_index_2057599_comb ^ p73_literal_2043916[p73_array_index_2057511] ^ p73_literal_2043914[p73_array_index_2057522] ^ p73_literal_2043912[p73_array_index_2057513] ^ p73_literal_2043910[p73_array_index_2057523] ^ p73_array_index_2057515;

  // Registers for pipe stage 74:
  reg [127:0] p74_encoded;
  reg [127:0] p74_bit_slice_2043893;
  reg [127:0] p74_bit_slice_2044018;
  reg [127:0] p74_k3;
  reg [127:0] p74_k2;
  reg [127:0] p74_k5;
  reg [127:0] p74_k4;
  reg [127:0] p74_k7;
  reg [127:0] p74_k6;
  reg [127:0] p74_xor_2057042;
  reg [127:0] p74_xor_2057490;
  reg [7:0] p74_array_index_2057506;
  reg [7:0] p74_array_index_2057507;
  reg [7:0] p74_array_index_2057508;
  reg [7:0] p74_array_index_2057509;
  reg [7:0] p74_array_index_2057510;
  reg [7:0] p74_array_index_2057511;
  reg [7:0] p74_array_index_2057513;
  reg [7:0] p74_array_index_2057595;
  reg [7:0] p74_array_index_2057596;
  reg [7:0] p74_array_index_2057597;
  reg [7:0] p74_array_index_2057598;
  reg [7:0] p74_array_index_2057522;
  reg [7:0] p74_array_index_2057523;
  reg [7:0] p74_res7__960;
  reg [7:0] p74_array_index_2057609;
  reg [7:0] p74_array_index_2057610;
  reg [7:0] p74_array_index_2057611;
  reg [7:0] p74_array_index_2057612;
  reg [7:0] p74_array_index_2057613;
  reg [7:0] p74_res7__962;
  reg [7:0] p74_array_index_2057624;
  reg [7:0] p74_array_index_2057625;
  reg [7:0] p74_array_index_2057626;
  reg [7:0] p74_array_index_2057627;
  reg [7:0] p74_res7__964;
  reg [7:0] p74_array_index_2057638;
  reg [7:0] p74_array_index_2057639;
  reg [7:0] p74_array_index_2057640;
  reg [7:0] p74_array_index_2057641;
  reg [7:0] p74_array_index_2057642;
  reg [7:0] p74_res7__966;
  reg [7:0] p74_array_index_2057653;
  reg [7:0] p74_array_index_2057654;
  reg [7:0] p74_array_index_2057655;
  reg [7:0] p74_array_index_2057656;
  reg [7:0] p74_res7__968;
  reg [7:0] p74_array_index_2057666;
  reg [7:0] p74_array_index_2057667;
  reg [7:0] p74_array_index_2057668;
  reg [7:0] p74_array_index_2057669;
  reg [7:0] p74_res7__970;
  reg [7:0] p74_array_index_2057680;
  reg [7:0] p74_array_index_2057681;
  reg [7:0] p74_array_index_2057682;
  reg [7:0] p74_res7__972;
  reg [7:0] p75_literal_2043896[256];
  reg [7:0] p75_literal_2043910[256];
  reg [7:0] p75_literal_2043912[256];
  reg [7:0] p75_literal_2043914[256];
  reg [7:0] p75_literal_2043916[256];
  reg [7:0] p75_literal_2043918[256];
  reg [7:0] p75_literal_2043920[256];
  reg [7:0] p75_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p74_encoded <= p73_encoded;
    p74_bit_slice_2043893 <= p73_bit_slice_2043893;
    p74_bit_slice_2044018 <= p73_bit_slice_2044018;
    p74_k3 <= p73_k3;
    p74_k2 <= p73_k2;
    p74_k5 <= p73_k5;
    p74_k4 <= p73_k4;
    p74_k7 <= p73_k7;
    p74_k6 <= p73_k6;
    p74_xor_2057042 <= p73_xor_2057042;
    p74_xor_2057490 <= p73_xor_2057490;
    p74_array_index_2057506 <= p73_array_index_2057506;
    p74_array_index_2057507 <= p73_array_index_2057507;
    p74_array_index_2057508 <= p73_array_index_2057508;
    p74_array_index_2057509 <= p73_array_index_2057509;
    p74_array_index_2057510 <= p73_array_index_2057510;
    p74_array_index_2057511 <= p73_array_index_2057511;
    p74_array_index_2057513 <= p73_array_index_2057513;
    p74_array_index_2057595 <= p74_array_index_2057595_comb;
    p74_array_index_2057596 <= p74_array_index_2057596_comb;
    p74_array_index_2057597 <= p74_array_index_2057597_comb;
    p74_array_index_2057598 <= p74_array_index_2057598_comb;
    p74_array_index_2057522 <= p73_array_index_2057522;
    p74_array_index_2057523 <= p73_array_index_2057523;
    p74_res7__960 <= p74_res7__960_comb;
    p74_array_index_2057609 <= p74_array_index_2057609_comb;
    p74_array_index_2057610 <= p74_array_index_2057610_comb;
    p74_array_index_2057611 <= p74_array_index_2057611_comb;
    p74_array_index_2057612 <= p74_array_index_2057612_comb;
    p74_array_index_2057613 <= p74_array_index_2057613_comb;
    p74_res7__962 <= p74_res7__962_comb;
    p74_array_index_2057624 <= p74_array_index_2057624_comb;
    p74_array_index_2057625 <= p74_array_index_2057625_comb;
    p74_array_index_2057626 <= p74_array_index_2057626_comb;
    p74_array_index_2057627 <= p74_array_index_2057627_comb;
    p74_res7__964 <= p74_res7__964_comb;
    p74_array_index_2057638 <= p74_array_index_2057638_comb;
    p74_array_index_2057639 <= p74_array_index_2057639_comb;
    p74_array_index_2057640 <= p74_array_index_2057640_comb;
    p74_array_index_2057641 <= p74_array_index_2057641_comb;
    p74_array_index_2057642 <= p74_array_index_2057642_comb;
    p74_res7__966 <= p74_res7__966_comb;
    p74_array_index_2057653 <= p74_array_index_2057653_comb;
    p74_array_index_2057654 <= p74_array_index_2057654_comb;
    p74_array_index_2057655 <= p74_array_index_2057655_comb;
    p74_array_index_2057656 <= p74_array_index_2057656_comb;
    p74_res7__968 <= p74_res7__968_comb;
    p74_array_index_2057666 <= p74_array_index_2057666_comb;
    p74_array_index_2057667 <= p74_array_index_2057667_comb;
    p74_array_index_2057668 <= p74_array_index_2057668_comb;
    p74_array_index_2057669 <= p74_array_index_2057669_comb;
    p74_res7__970 <= p74_res7__970_comb;
    p74_array_index_2057680 <= p74_array_index_2057680_comb;
    p74_array_index_2057681 <= p74_array_index_2057681_comb;
    p74_array_index_2057682 <= p74_array_index_2057682_comb;
    p74_res7__972 <= p74_res7__972_comb;
    p75_literal_2043896 <= p74_literal_2043896;
    p75_literal_2043910 <= p74_literal_2043910;
    p75_literal_2043912 <= p74_literal_2043912;
    p75_literal_2043914 <= p74_literal_2043914;
    p75_literal_2043916 <= p74_literal_2043916;
    p75_literal_2043918 <= p74_literal_2043918;
    p75_literal_2043920 <= p74_literal_2043920;
    p75_literal_2043923 <= p74_literal_2043923;
  end

  // ===== Pipe stage 75:
  wire [7:0] p75_array_index_2057820_comb;
  wire [7:0] p75_array_index_2057821_comb;
  wire [7:0] p75_array_index_2057822_comb;
  wire [7:0] p75_res7__974_comb;
  wire [7:0] p75_array_index_2057833_comb;
  wire [7:0] p75_array_index_2057834_comb;
  wire [7:0] p75_res7__976_comb;
  wire [7:0] p75_array_index_2057844_comb;
  wire [7:0] p75_array_index_2057845_comb;
  wire [7:0] p75_res7__978_comb;
  wire [7:0] p75_array_index_2057856_comb;
  wire [7:0] p75_res7__980_comb;
  wire [7:0] p75_array_index_2057866_comb;
  wire [7:0] p75_res7__982_comb;
  wire [7:0] p75_res7__984_comb;
  wire [7:0] p75_res7__986_comb;
  assign p75_array_index_2057820_comb = p74_literal_2043916[p74_res7__966];
  assign p75_array_index_2057821_comb = p74_literal_2043918[p74_res7__964];
  assign p75_array_index_2057822_comb = p74_literal_2043920[p74_res7__962];
  assign p75_res7__974_comb = p74_literal_2043910[p74_res7__972] ^ p74_literal_2043912[p74_res7__970] ^ p74_literal_2043914[p74_res7__968] ^ p75_array_index_2057820_comb ^ p75_array_index_2057821_comb ^ p75_array_index_2057822_comb ^ p74_res7__960 ^ p74_literal_2043923[p74_array_index_2057506] ^ p74_array_index_2057507 ^ p74_array_index_2057642 ^ p74_array_index_2057613 ^ p74_literal_2043916[p74_array_index_2057510] ^ p74_literal_2043914[p74_array_index_2057511] ^ p74_literal_2043912[p74_array_index_2057522] ^ p74_literal_2043910[p74_array_index_2057513] ^ p74_array_index_2057523;
  assign p75_array_index_2057833_comb = p74_literal_2043918[p74_res7__966];
  assign p75_array_index_2057834_comb = p74_literal_2043920[p74_res7__964];
  assign p75_res7__976_comb = p74_literal_2043910[p75_res7__974_comb] ^ p74_literal_2043912[p74_res7__972] ^ p74_literal_2043914[p74_res7__970] ^ p74_literal_2043916[p74_res7__968] ^ p75_array_index_2057833_comb ^ p75_array_index_2057834_comb ^ p74_res7__962 ^ p74_literal_2043923[p74_res7__960] ^ p74_array_index_2057506 ^ p74_array_index_2057656 ^ p74_array_index_2057627 ^ p74_array_index_2057598 ^ p74_literal_2043914[p74_array_index_2057510] ^ p74_literal_2043912[p74_array_index_2057511] ^ p74_literal_2043910[p74_array_index_2057522] ^ p74_array_index_2057513;
  assign p75_array_index_2057844_comb = p74_literal_2043918[p74_res7__968];
  assign p75_array_index_2057845_comb = p74_literal_2043920[p74_res7__966];
  assign p75_res7__978_comb = p74_literal_2043910[p75_res7__976_comb] ^ p74_literal_2043912[p75_res7__974_comb] ^ p74_literal_2043914[p74_res7__972] ^ p74_literal_2043916[p74_res7__970] ^ p75_array_index_2057844_comb ^ p75_array_index_2057845_comb ^ p74_res7__964 ^ p74_literal_2043923[p74_res7__962] ^ p74_res7__960 ^ p74_array_index_2057669 ^ p74_array_index_2057641 ^ p74_array_index_2057612 ^ p74_literal_2043914[p74_array_index_2057509] ^ p74_literal_2043912[p74_array_index_2057510] ^ p74_literal_2043910[p74_array_index_2057511] ^ p74_array_index_2057522;
  assign p75_array_index_2057856_comb = p74_literal_2043920[p74_res7__968];
  assign p75_res7__980_comb = p74_literal_2043910[p75_res7__978_comb] ^ p74_literal_2043912[p75_res7__976_comb] ^ p74_literal_2043914[p75_res7__974_comb] ^ p74_literal_2043916[p74_res7__972] ^ p74_literal_2043918[p74_res7__970] ^ p75_array_index_2057856_comb ^ p74_res7__966 ^ p74_literal_2043923[p74_res7__964] ^ p74_res7__962 ^ p74_array_index_2057682 ^ p74_array_index_2057655 ^ p74_array_index_2057626 ^ p74_array_index_2057597 ^ p74_literal_2043912[p74_array_index_2057509] ^ p74_literal_2043910[p74_array_index_2057510] ^ p74_array_index_2057511;
  assign p75_array_index_2057866_comb = p74_literal_2043920[p74_res7__970];
  assign p75_res7__982_comb = p74_literal_2043910[p75_res7__980_comb] ^ p74_literal_2043912[p75_res7__978_comb] ^ p74_literal_2043914[p75_res7__976_comb] ^ p74_literal_2043916[p75_res7__974_comb] ^ p74_literal_2043918[p74_res7__972] ^ p75_array_index_2057866_comb ^ p74_res7__968 ^ p74_literal_2043923[p74_res7__966] ^ p74_res7__964 ^ p75_array_index_2057822_comb ^ p74_array_index_2057668 ^ p74_array_index_2057640 ^ p74_array_index_2057611 ^ p74_literal_2043912[p74_array_index_2057508] ^ p74_literal_2043910[p74_array_index_2057509] ^ p74_array_index_2057510;
  assign p75_res7__984_comb = p74_literal_2043910[p75_res7__982_comb] ^ p74_literal_2043912[p75_res7__980_comb] ^ p74_literal_2043914[p75_res7__978_comb] ^ p74_literal_2043916[p75_res7__976_comb] ^ p74_literal_2043918[p75_res7__974_comb] ^ p74_literal_2043920[p74_res7__972] ^ p74_res7__970 ^ p74_literal_2043923[p74_res7__968] ^ p74_res7__966 ^ p75_array_index_2057834_comb ^ p74_array_index_2057681 ^ p74_array_index_2057654 ^ p74_array_index_2057625 ^ p74_array_index_2057596 ^ p74_literal_2043910[p74_array_index_2057508] ^ p74_array_index_2057509;
  assign p75_res7__986_comb = p74_literal_2043910[p75_res7__984_comb] ^ p74_literal_2043912[p75_res7__982_comb] ^ p74_literal_2043914[p75_res7__980_comb] ^ p74_literal_2043916[p75_res7__978_comb] ^ p74_literal_2043918[p75_res7__976_comb] ^ p74_literal_2043920[p75_res7__974_comb] ^ p74_res7__972 ^ p74_literal_2043923[p74_res7__970] ^ p74_res7__968 ^ p75_array_index_2057845_comb ^ p75_array_index_2057821_comb ^ p74_array_index_2057667 ^ p74_array_index_2057639 ^ p74_array_index_2057610 ^ p74_literal_2043910[p74_array_index_2057507] ^ p74_array_index_2057508;

  // Registers for pipe stage 75:
  reg [127:0] p75_encoded;
  reg [127:0] p75_bit_slice_2043893;
  reg [127:0] p75_bit_slice_2044018;
  reg [127:0] p75_k3;
  reg [127:0] p75_k2;
  reg [127:0] p75_k5;
  reg [127:0] p75_k4;
  reg [127:0] p75_k7;
  reg [127:0] p75_k6;
  reg [127:0] p75_xor_2057042;
  reg [127:0] p75_xor_2057490;
  reg [7:0] p75_array_index_2057506;
  reg [7:0] p75_array_index_2057507;
  reg [7:0] p75_array_index_2057595;
  reg [7:0] p75_res7__960;
  reg [7:0] p75_array_index_2057609;
  reg [7:0] p75_res7__962;
  reg [7:0] p75_array_index_2057624;
  reg [7:0] p75_res7__964;
  reg [7:0] p75_array_index_2057638;
  reg [7:0] p75_res7__966;
  reg [7:0] p75_array_index_2057653;
  reg [7:0] p75_res7__968;
  reg [7:0] p75_array_index_2057666;
  reg [7:0] p75_res7__970;
  reg [7:0] p75_array_index_2057680;
  reg [7:0] p75_res7__972;
  reg [7:0] p75_array_index_2057820;
  reg [7:0] p75_res7__974;
  reg [7:0] p75_array_index_2057833;
  reg [7:0] p75_res7__976;
  reg [7:0] p75_array_index_2057844;
  reg [7:0] p75_res7__978;
  reg [7:0] p75_array_index_2057856;
  reg [7:0] p75_res7__980;
  reg [7:0] p75_array_index_2057866;
  reg [7:0] p75_res7__982;
  reg [7:0] p75_res7__984;
  reg [7:0] p75_res7__986;
  reg [7:0] p76_literal_2043910[256];
  reg [7:0] p76_literal_2043912[256];
  reg [7:0] p76_literal_2043914[256];
  reg [7:0] p76_literal_2043916[256];
  reg [7:0] p76_literal_2043918[256];
  reg [7:0] p76_literal_2043920[256];
  reg [7:0] p76_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p75_encoded <= p74_encoded;
    p75_bit_slice_2043893 <= p74_bit_slice_2043893;
    p75_bit_slice_2044018 <= p74_bit_slice_2044018;
    p75_k3 <= p74_k3;
    p75_k2 <= p74_k2;
    p75_k5 <= p74_k5;
    p75_k4 <= p74_k4;
    p75_k7 <= p74_k7;
    p75_k6 <= p74_k6;
    p75_xor_2057042 <= p74_xor_2057042;
    p75_xor_2057490 <= p74_xor_2057490;
    p75_array_index_2057506 <= p74_array_index_2057506;
    p75_array_index_2057507 <= p74_array_index_2057507;
    p75_array_index_2057595 <= p74_array_index_2057595;
    p75_res7__960 <= p74_res7__960;
    p75_array_index_2057609 <= p74_array_index_2057609;
    p75_res7__962 <= p74_res7__962;
    p75_array_index_2057624 <= p74_array_index_2057624;
    p75_res7__964 <= p74_res7__964;
    p75_array_index_2057638 <= p74_array_index_2057638;
    p75_res7__966 <= p74_res7__966;
    p75_array_index_2057653 <= p74_array_index_2057653;
    p75_res7__968 <= p74_res7__968;
    p75_array_index_2057666 <= p74_array_index_2057666;
    p75_res7__970 <= p74_res7__970;
    p75_array_index_2057680 <= p74_array_index_2057680;
    p75_res7__972 <= p74_res7__972;
    p75_array_index_2057820 <= p75_array_index_2057820_comb;
    p75_res7__974 <= p75_res7__974_comb;
    p75_array_index_2057833 <= p75_array_index_2057833_comb;
    p75_res7__976 <= p75_res7__976_comb;
    p75_array_index_2057844 <= p75_array_index_2057844_comb;
    p75_res7__978 <= p75_res7__978_comb;
    p75_array_index_2057856 <= p75_array_index_2057856_comb;
    p75_res7__980 <= p75_res7__980_comb;
    p75_array_index_2057866 <= p75_array_index_2057866_comb;
    p75_res7__982 <= p75_res7__982_comb;
    p75_res7__984 <= p75_res7__984_comb;
    p75_res7__986 <= p75_res7__986_comb;
    p76_literal_2043910 <= p75_literal_2043910;
    p76_literal_2043912 <= p75_literal_2043912;
    p76_literal_2043914 <= p75_literal_2043914;
    p76_literal_2043916 <= p75_literal_2043916;
    p76_literal_2043918 <= p75_literal_2043918;
    p76_literal_2043920 <= p75_literal_2043920;
    p76_literal_2043923 <= p75_literal_2043923;
  end

  // ===== Pipe stage 76:
  wire [7:0] p76_res7__988_comb;
  wire [7:0] p76_res7__990_comb;
  wire [127:0] p76_res__30_comb;
  wire [127:0] p76_k9_comb;
  wire [127:0] p76_addedKey__63_comb;
  wire [127:0] p76_xor_2058003_comb;
  wire [7:0] p76_bit_slice_2058020_comb;
  wire [7:0] p76_bit_slice_2058021_comb;
  wire [7:0] p76_bit_slice_2058022_comb;
  wire [7:0] p76_bit_slice_2058023_comb;
  wire [7:0] p76_bit_slice_2058024_comb;
  wire [7:0] p76_bit_slice_2058025_comb;
  wire [7:0] p76_bit_slice_2058026_comb;
  wire [7:0] p76_bit_slice_2058027_comb;
  wire [7:0] p76_bit_slice_2058028_comb;
  wire [7:0] p76_bit_slice_2058029_comb;
  wire [7:0] p76_array_index_2058030_comb;
  wire [7:0] p76_array_index_2058031_comb;
  wire [7:0] p76_array_index_2058032_comb;
  wire [7:0] p76_array_index_2058033_comb;
  wire [7:0] p76_array_index_2058034_comb;
  wire [7:0] p76_array_index_2058035_comb;
  wire [7:0] p76_array_index_2058037_comb;
  wire [7:0] p76_array_index_2058039_comb;
  wire [7:0] p76_array_index_2058040_comb;
  wire [7:0] p76_array_index_2058041_comb;
  wire [7:0] p76_array_index_2058042_comb;
  wire [7:0] p76_array_index_2058043_comb;
  wire [7:0] p76_array_index_2058044_comb;
  wire [7:0] p76_bit_slice_2058052_comb;
  wire [7:0] p76_bit_slice_2058054_comb;
  wire [7:0] p76_array_index_2058055_comb;
  wire [7:0] p76_array_index_2058056_comb;
  wire [7:0] p76_array_index_2058057_comb;
  wire [7:0] p76_array_index_2058058_comb;
  wire [7:0] p76_array_index_2058059_comb;
  wire [7:0] p76_array_index_2058060_comb;
  wire [7:0] p76_array_index_2058062_comb;
  wire [7:0] p76_array_index_2058063_comb;
  wire [7:0] p76_array_index_2058064_comb;
  wire [7:0] p76_array_index_2058065_comb;
  wire [7:0] p76_array_index_2058066_comb;
  wire [7:0] p76_array_index_2058067_comb;
  wire [7:0] p76_array_index_2058068_comb;
  wire [7:0] p76_array_index_2058070_comb;
  wire [7:0] p76_res7__1025_comb;
  wire [7:0] p76_res7__992_comb;
  wire [7:0] p76_array_index_2058087_comb;
  wire [7:0] p76_array_index_2058088_comb;
  wire [7:0] p76_array_index_2058089_comb;
  wire [7:0] p76_array_index_2058090_comb;
  wire [7:0] p76_array_index_2058091_comb;
  wire [7:0] p76_array_index_2058092_comb;
  wire [7:0] p76_array_index_2058093_comb;
  wire [7:0] p76_array_index_2058094_comb;
  wire [7:0] p76_array_index_2058095_comb;
  wire [7:0] p76_array_index_2058096_comb;
  wire [7:0] p76_array_index_2058097_comb;
  wire [7:0] p76_array_index_2058098_comb;
  wire [7:0] p76_res7__1027_comb;
  wire [7:0] p76_res7__994_comb;
  wire [7:0] p76_array_index_2058115_comb;
  wire [7:0] p76_array_index_2058116_comb;
  wire [7:0] p76_array_index_2058117_comb;
  wire [7:0] p76_array_index_2058118_comb;
  wire [7:0] p76_array_index_2058119_comb;
  wire [7:0] p76_array_index_2058122_comb;
  wire [7:0] p76_array_index_2058123_comb;
  wire [7:0] p76_array_index_2058124_comb;
  wire [7:0] p76_array_index_2058125_comb;
  wire [7:0] p76_array_index_2058126_comb;
  wire [7:0] p76_res7__1029_comb;
  wire [7:0] p76_res7__996_comb;
  wire [7:0] p76_array_index_2058143_comb;
  wire [7:0] p76_array_index_2058144_comb;
  wire [7:0] p76_array_index_2058145_comb;
  wire [7:0] p76_array_index_2058146_comb;
  wire [7:0] p76_array_index_2058147_comb;
  wire [7:0] p76_array_index_2058150_comb;
  wire [7:0] p76_array_index_2058151_comb;
  wire [7:0] p76_array_index_2058152_comb;
  wire [7:0] p76_array_index_2058153_comb;
  wire [7:0] p76_array_index_2058154_comb;
  wire [7:0] p76_res7__1031_comb;
  wire [7:0] p76_res7__998_comb;
  wire [7:0] p76_array_index_2058164_comb;
  wire [7:0] p76_array_index_2058165_comb;
  wire [7:0] p76_array_index_2058166_comb;
  wire [7:0] p76_array_index_2058167_comb;
  wire [7:0] p76_array_index_2058168_comb;
  wire [7:0] p76_array_index_2058169_comb;
  wire [7:0] p76_array_index_2058170_comb;
  wire [7:0] p76_array_index_2058171_comb;
  wire [7:0] p76_array_index_2058172_comb;
  wire [7:0] p76_array_index_2058173_comb;
  wire [7:0] p76_array_index_2058174_comb;
  wire [7:0] p76_array_index_2058175_comb;
  assign p76_res7__988_comb = p75_literal_2043910[p75_res7__986] ^ p75_literal_2043912[p75_res7__984] ^ p75_literal_2043914[p75_res7__982] ^ p75_literal_2043916[p75_res7__980] ^ p75_literal_2043918[p75_res7__978] ^ p75_literal_2043920[p75_res7__976] ^ p75_res7__974 ^ p75_literal_2043923[p75_res7__972] ^ p75_res7__970 ^ p75_array_index_2057856 ^ p75_array_index_2057833 ^ p75_array_index_2057680 ^ p75_array_index_2057653 ^ p75_array_index_2057624 ^ p75_array_index_2057595 ^ p75_array_index_2057507;
  assign p76_res7__990_comb = p75_literal_2043910[p76_res7__988_comb] ^ p75_literal_2043912[p75_res7__986] ^ p75_literal_2043914[p75_res7__984] ^ p75_literal_2043916[p75_res7__982] ^ p75_literal_2043918[p75_res7__980] ^ p75_literal_2043920[p75_res7__978] ^ p75_res7__976 ^ p75_literal_2043923[p75_res7__974] ^ p75_res7__972 ^ p75_array_index_2057866 ^ p75_array_index_2057844 ^ p75_array_index_2057820 ^ p75_array_index_2057666 ^ p75_array_index_2057638 ^ p75_array_index_2057609 ^ p75_array_index_2057506;
  assign p76_res__30_comb = {p76_res7__990_comb, p76_res7__988_comb, p75_res7__986, p75_res7__984, p75_res7__982, p75_res7__980, p75_res7__978, p75_res7__976, p75_res7__974, p75_res7__972, p75_res7__970, p75_res7__968, p75_res7__966, p75_res7__964, p75_res7__962, p75_res7__960};
  assign p76_k9_comb = p76_res__30_comb ^ p75_xor_2057042;
  assign p76_addedKey__63_comb = p76_k9_comb ^ 128'h5ea7_d858_1e14_9b61_f16a_c145_9ced_a820;
  assign p76_xor_2058003_comb = p75_encoded ^ p76_k9_comb;
  assign p76_bit_slice_2058020_comb = p76_xor_2058003_comb[95:88];
  assign p76_bit_slice_2058021_comb = p76_xor_2058003_comb[87:80];
  assign p76_bit_slice_2058022_comb = p76_xor_2058003_comb[79:72];
  assign p76_bit_slice_2058023_comb = p76_xor_2058003_comb[63:56];
  assign p76_bit_slice_2058024_comb = p76_xor_2058003_comb[47:40];
  assign p76_bit_slice_2058025_comb = p76_xor_2058003_comb[39:32];
  assign p76_bit_slice_2058026_comb = p76_xor_2058003_comb[31:24];
  assign p76_bit_slice_2058027_comb = p76_xor_2058003_comb[23:16];
  assign p76_bit_slice_2058028_comb = p76_xor_2058003_comb[15:8];
  assign p76_bit_slice_2058029_comb = p76_xor_2058003_comb[7:0];
  assign p76_array_index_2058030_comb = p75_literal_2043896[p76_addedKey__63_comb[127:120]];
  assign p76_array_index_2058031_comb = p75_literal_2043896[p76_addedKey__63_comb[119:112]];
  assign p76_array_index_2058032_comb = p75_literal_2043896[p76_addedKey__63_comb[111:104]];
  assign p76_array_index_2058033_comb = p75_literal_2043896[p76_addedKey__63_comb[103:96]];
  assign p76_array_index_2058034_comb = p75_literal_2043896[p76_addedKey__63_comb[95:88]];
  assign p76_array_index_2058035_comb = p75_literal_2043896[p76_addedKey__63_comb[87:80]];
  assign p76_array_index_2058037_comb = p75_literal_2043896[p76_addedKey__63_comb[71:64]];
  assign p76_array_index_2058039_comb = p75_literal_2043896[p76_addedKey__63_comb[55:48]];
  assign p76_array_index_2058040_comb = p75_literal_2043896[p76_addedKey__63_comb[47:40]];
  assign p76_array_index_2058041_comb = p75_literal_2043896[p76_addedKey__63_comb[39:32]];
  assign p76_array_index_2058042_comb = p75_literal_2043896[p76_addedKey__63_comb[31:24]];
  assign p76_array_index_2058043_comb = p75_literal_2043896[p76_addedKey__63_comb[23:16]];
  assign p76_array_index_2058044_comb = p75_literal_2043896[p76_addedKey__63_comb[15:8]];
  assign p76_bit_slice_2058052_comb = p76_xor_2058003_comb[71:64];
  assign p76_bit_slice_2058054_comb = p76_xor_2058003_comb[55:48];
  assign p76_array_index_2058055_comb = p75_literal_2043920[p76_bit_slice_2058024_comb];
  assign p76_array_index_2058056_comb = p75_literal_2043918[p76_bit_slice_2058025_comb];
  assign p76_array_index_2058057_comb = p75_literal_2043916[p76_bit_slice_2058026_comb];
  assign p76_array_index_2058058_comb = p75_literal_2043914[p76_bit_slice_2058027_comb];
  assign p76_array_index_2058059_comb = p75_literal_2043912[p76_bit_slice_2058028_comb];
  assign p76_array_index_2058060_comb = p75_literal_2043910[p76_bit_slice_2058029_comb];
  assign p76_array_index_2058062_comb = p75_literal_2043910[p76_array_index_2058030_comb];
  assign p76_array_index_2058063_comb = p75_literal_2043912[p76_array_index_2058031_comb];
  assign p76_array_index_2058064_comb = p75_literal_2043914[p76_array_index_2058032_comb];
  assign p76_array_index_2058065_comb = p75_literal_2043916[p76_array_index_2058033_comb];
  assign p76_array_index_2058066_comb = p75_literal_2043918[p76_array_index_2058034_comb];
  assign p76_array_index_2058067_comb = p75_literal_2043920[p76_array_index_2058035_comb];
  assign p76_array_index_2058068_comb = p75_literal_2043896[p76_addedKey__63_comb[79:72]];
  assign p76_array_index_2058070_comb = p75_literal_2043896[p76_addedKey__63_comb[63:56]];
  assign p76_res7__1025_comb = p75_literal_2043910[p76_xor_2058003_comb[119:112]] ^ p75_literal_2043912[p76_xor_2058003_comb[111:104]] ^ p75_literal_2043914[p76_xor_2058003_comb[103:96]] ^ p75_literal_2043916[p76_bit_slice_2058020_comb] ^ p75_literal_2043918[p76_bit_slice_2058021_comb] ^ p75_literal_2043920[p76_bit_slice_2058022_comb] ^ p76_bit_slice_2058052_comb ^ p75_literal_2043923[p76_bit_slice_2058023_comb] ^ p76_bit_slice_2058054_comb ^ p76_array_index_2058055_comb ^ p76_array_index_2058056_comb ^ p76_array_index_2058057_comb ^ p76_array_index_2058058_comb ^ p76_array_index_2058059_comb ^ p76_array_index_2058060_comb ^ p76_xor_2058003_comb[127:120];
  assign p76_res7__992_comb = p76_array_index_2058062_comb ^ p76_array_index_2058063_comb ^ p76_array_index_2058064_comb ^ p76_array_index_2058065_comb ^ p76_array_index_2058066_comb ^ p76_array_index_2058067_comb ^ p76_array_index_2058068_comb ^ p75_literal_2043923[p76_array_index_2058037_comb] ^ p76_array_index_2058070_comb ^ p75_literal_2043920[p76_array_index_2058039_comb] ^ p75_literal_2043918[p76_array_index_2058040_comb] ^ p75_literal_2043916[p76_array_index_2058041_comb] ^ p75_literal_2043914[p76_array_index_2058042_comb] ^ p75_literal_2043912[p76_array_index_2058043_comb] ^ p75_literal_2043910[p76_array_index_2058044_comb] ^ p75_literal_2043896[p76_addedKey__63_comb[7:0]];
  assign p76_array_index_2058087_comb = p75_literal_2043920[p76_bit_slice_2058025_comb];
  assign p76_array_index_2058088_comb = p75_literal_2043918[p76_bit_slice_2058026_comb];
  assign p76_array_index_2058089_comb = p75_literal_2043916[p76_bit_slice_2058027_comb];
  assign p76_array_index_2058090_comb = p75_literal_2043914[p76_bit_slice_2058028_comb];
  assign p76_array_index_2058091_comb = p75_literal_2043912[p76_bit_slice_2058029_comb];
  assign p76_array_index_2058092_comb = p75_literal_2043910[p76_res7__1025_comb];
  assign p76_array_index_2058093_comb = p75_literal_2043910[p76_res7__992_comb];
  assign p76_array_index_2058094_comb = p75_literal_2043912[p76_array_index_2058030_comb];
  assign p76_array_index_2058095_comb = p75_literal_2043914[p76_array_index_2058031_comb];
  assign p76_array_index_2058096_comb = p75_literal_2043916[p76_array_index_2058032_comb];
  assign p76_array_index_2058097_comb = p75_literal_2043918[p76_array_index_2058033_comb];
  assign p76_array_index_2058098_comb = p75_literal_2043920[p76_array_index_2058034_comb];
  assign p76_res7__1027_comb = p75_literal_2043910[p76_xor_2058003_comb[111:104]] ^ p75_literal_2043912[p76_xor_2058003_comb[103:96]] ^ p75_literal_2043914[p76_bit_slice_2058020_comb] ^ p75_literal_2043916[p76_bit_slice_2058021_comb] ^ p75_literal_2043918[p76_bit_slice_2058022_comb] ^ p75_literal_2043920[p76_bit_slice_2058052_comb] ^ p76_bit_slice_2058023_comb ^ p75_literal_2043923[p76_bit_slice_2058054_comb] ^ p76_bit_slice_2058024_comb ^ p76_array_index_2058087_comb ^ p76_array_index_2058088_comb ^ p76_array_index_2058089_comb ^ p76_array_index_2058090_comb ^ p76_array_index_2058091_comb ^ p76_array_index_2058092_comb ^ p76_xor_2058003_comb[119:112];
  assign p76_res7__994_comb = p76_array_index_2058093_comb ^ p76_array_index_2058094_comb ^ p76_array_index_2058095_comb ^ p76_array_index_2058096_comb ^ p76_array_index_2058097_comb ^ p76_array_index_2058098_comb ^ p76_array_index_2058035_comb ^ p75_literal_2043923[p76_array_index_2058068_comb] ^ p76_array_index_2058037_comb ^ p75_literal_2043920[p76_array_index_2058070_comb] ^ p75_literal_2043918[p76_array_index_2058039_comb] ^ p75_literal_2043916[p76_array_index_2058040_comb] ^ p75_literal_2043914[p76_array_index_2058041_comb] ^ p75_literal_2043912[p76_array_index_2058042_comb] ^ p75_literal_2043910[p76_array_index_2058043_comb] ^ p76_array_index_2058044_comb;
  assign p76_array_index_2058115_comb = p75_literal_2043920[p76_bit_slice_2058026_comb];
  assign p76_array_index_2058116_comb = p75_literal_2043918[p76_bit_slice_2058027_comb];
  assign p76_array_index_2058117_comb = p75_literal_2043916[p76_bit_slice_2058028_comb];
  assign p76_array_index_2058118_comb = p75_literal_2043914[p76_bit_slice_2058029_comb];
  assign p76_array_index_2058119_comb = p75_literal_2043912[p76_res7__1025_comb];
  assign p76_array_index_2058122_comb = p75_literal_2043912[p76_res7__992_comb];
  assign p76_array_index_2058123_comb = p75_literal_2043914[p76_array_index_2058030_comb];
  assign p76_array_index_2058124_comb = p75_literal_2043916[p76_array_index_2058031_comb];
  assign p76_array_index_2058125_comb = p75_literal_2043918[p76_array_index_2058032_comb];
  assign p76_array_index_2058126_comb = p75_literal_2043920[p76_array_index_2058033_comb];
  assign p76_res7__1029_comb = p75_literal_2043910[p76_xor_2058003_comb[103:96]] ^ p75_literal_2043912[p76_bit_slice_2058020_comb] ^ p75_literal_2043914[p76_bit_slice_2058021_comb] ^ p75_literal_2043916[p76_bit_slice_2058022_comb] ^ p75_literal_2043918[p76_bit_slice_2058052_comb] ^ p75_literal_2043920[p76_bit_slice_2058023_comb] ^ p76_bit_slice_2058054_comb ^ p75_literal_2043923[p76_bit_slice_2058024_comb] ^ p76_bit_slice_2058025_comb ^ p76_array_index_2058115_comb ^ p76_array_index_2058116_comb ^ p76_array_index_2058117_comb ^ p76_array_index_2058118_comb ^ p76_array_index_2058119_comb ^ p75_literal_2043910[p76_res7__1027_comb] ^ p76_xor_2058003_comb[111:104];
  assign p76_res7__996_comb = p75_literal_2043910[p76_res7__994_comb] ^ p76_array_index_2058122_comb ^ p76_array_index_2058123_comb ^ p76_array_index_2058124_comb ^ p76_array_index_2058125_comb ^ p76_array_index_2058126_comb ^ p76_array_index_2058034_comb ^ p75_literal_2043923[p76_array_index_2058035_comb] ^ p76_array_index_2058068_comb ^ p75_literal_2043920[p76_array_index_2058037_comb] ^ p75_literal_2043918[p76_array_index_2058070_comb] ^ p75_literal_2043916[p76_array_index_2058039_comb] ^ p75_literal_2043914[p76_array_index_2058040_comb] ^ p75_literal_2043912[p76_array_index_2058041_comb] ^ p75_literal_2043910[p76_array_index_2058042_comb] ^ p76_array_index_2058043_comb;
  assign p76_array_index_2058143_comb = p75_literal_2043920[p76_bit_slice_2058027_comb];
  assign p76_array_index_2058144_comb = p75_literal_2043918[p76_bit_slice_2058028_comb];
  assign p76_array_index_2058145_comb = p75_literal_2043916[p76_bit_slice_2058029_comb];
  assign p76_array_index_2058146_comb = p75_literal_2043914[p76_res7__1025_comb];
  assign p76_array_index_2058147_comb = p75_literal_2043912[p76_res7__1027_comb];
  assign p76_array_index_2058150_comb = p75_literal_2043912[p76_res7__994_comb];
  assign p76_array_index_2058151_comb = p75_literal_2043914[p76_res7__992_comb];
  assign p76_array_index_2058152_comb = p75_literal_2043916[p76_array_index_2058030_comb];
  assign p76_array_index_2058153_comb = p75_literal_2043918[p76_array_index_2058031_comb];
  assign p76_array_index_2058154_comb = p75_literal_2043920[p76_array_index_2058032_comb];
  assign p76_res7__1031_comb = p75_literal_2043910[p76_bit_slice_2058020_comb] ^ p75_literal_2043912[p76_bit_slice_2058021_comb] ^ p75_literal_2043914[p76_bit_slice_2058022_comb] ^ p75_literal_2043916[p76_bit_slice_2058052_comb] ^ p75_literal_2043918[p76_bit_slice_2058023_comb] ^ p75_literal_2043920[p76_bit_slice_2058054_comb] ^ p76_bit_slice_2058024_comb ^ p75_literal_2043923[p76_bit_slice_2058025_comb] ^ p76_bit_slice_2058026_comb ^ p76_array_index_2058143_comb ^ p76_array_index_2058144_comb ^ p76_array_index_2058145_comb ^ p76_array_index_2058146_comb ^ p76_array_index_2058147_comb ^ p75_literal_2043910[p76_res7__1029_comb] ^ p76_xor_2058003_comb[103:96];
  assign p76_res7__998_comb = p75_literal_2043910[p76_res7__996_comb] ^ p76_array_index_2058150_comb ^ p76_array_index_2058151_comb ^ p76_array_index_2058152_comb ^ p76_array_index_2058153_comb ^ p76_array_index_2058154_comb ^ p76_array_index_2058033_comb ^ p75_literal_2043923[p76_array_index_2058034_comb] ^ p76_array_index_2058035_comb ^ p75_literal_2043920[p76_array_index_2058068_comb] ^ p75_literal_2043918[p76_array_index_2058037_comb] ^ p75_literal_2043916[p76_array_index_2058070_comb] ^ p75_literal_2043914[p76_array_index_2058039_comb] ^ p75_literal_2043912[p76_array_index_2058040_comb] ^ p75_literal_2043910[p76_array_index_2058041_comb] ^ p76_array_index_2058042_comb;
  assign p76_array_index_2058164_comb = p75_literal_2043910[p76_bit_slice_2058021_comb];
  assign p76_array_index_2058165_comb = p75_literal_2043912[p76_bit_slice_2058022_comb];
  assign p76_array_index_2058166_comb = p75_literal_2043914[p76_bit_slice_2058052_comb];
  assign p76_array_index_2058167_comb = p75_literal_2043916[p76_bit_slice_2058023_comb];
  assign p76_array_index_2058168_comb = p75_literal_2043918[p76_bit_slice_2058054_comb];
  assign p76_array_index_2058169_comb = p75_literal_2043923[p76_bit_slice_2058026_comb];
  assign p76_array_index_2058170_comb = p75_literal_2043920[p76_bit_slice_2058028_comb];
  assign p76_array_index_2058171_comb = p75_literal_2043918[p76_bit_slice_2058029_comb];
  assign p76_array_index_2058172_comb = p75_literal_2043916[p76_res7__1025_comb];
  assign p76_array_index_2058173_comb = p75_literal_2043914[p76_res7__1027_comb];
  assign p76_array_index_2058174_comb = p75_literal_2043912[p76_res7__1029_comb];
  assign p76_array_index_2058175_comb = p75_literal_2043910[p76_res7__1031_comb];

  // Registers for pipe stage 76:
  reg [127:0] p76_bit_slice_2043893;
  reg [127:0] p76_bit_slice_2044018;
  reg [127:0] p76_k3;
  reg [127:0] p76_k2;
  reg [127:0] p76_k5;
  reg [127:0] p76_k4;
  reg [127:0] p76_k7;
  reg [127:0] p76_k6;
  reg [127:0] p76_xor_2057490;
  reg [7:0] p76_bit_slice_2058020;
  reg [7:0] p76_bit_slice_2058021;
  reg [7:0] p76_bit_slice_2058022;
  reg [7:0] p76_bit_slice_2058023;
  reg [7:0] p76_bit_slice_2058024;
  reg [7:0] p76_bit_slice_2058025;
  reg [7:0] p76_bit_slice_2058026;
  reg [7:0] p76_bit_slice_2058027;
  reg [7:0] p76_bit_slice_2058028;
  reg [7:0] p76_bit_slice_2058029;
  reg [7:0] p76_array_index_2058030;
  reg [7:0] p76_array_index_2058031;
  reg [7:0] p76_array_index_2058032;
  reg [7:0] p76_array_index_2058033;
  reg [7:0] p76_array_index_2058034;
  reg [7:0] p76_array_index_2058035;
  reg [7:0] p76_array_index_2058037;
  reg [7:0] p76_array_index_2058039;
  reg [7:0] p76_array_index_2058040;
  reg [7:0] p76_array_index_2058041;
  reg [7:0] p76_bit_slice_2058052;
  reg [7:0] p76_bit_slice_2058054;
  reg [7:0] p76_array_index_2058055;
  reg [7:0] p76_array_index_2058056;
  reg [7:0] p76_array_index_2058057;
  reg [7:0] p76_array_index_2058058;
  reg [7:0] p76_array_index_2058059;
  reg [7:0] p76_array_index_2058060;
  reg [7:0] p76_array_index_2058062;
  reg [7:0] p76_array_index_2058063;
  reg [7:0] p76_array_index_2058064;
  reg [7:0] p76_array_index_2058065;
  reg [7:0] p76_array_index_2058066;
  reg [7:0] p76_array_index_2058067;
  reg [7:0] p76_array_index_2058068;
  reg [7:0] p76_array_index_2058070;
  reg [7:0] p76_res7__1025;
  reg [7:0] p76_res7__992;
  reg [7:0] p76_array_index_2058087;
  reg [7:0] p76_array_index_2058088;
  reg [7:0] p76_array_index_2058089;
  reg [7:0] p76_array_index_2058090;
  reg [7:0] p76_array_index_2058091;
  reg [7:0] p76_array_index_2058092;
  reg [7:0] p76_array_index_2058093;
  reg [7:0] p76_array_index_2058094;
  reg [7:0] p76_array_index_2058095;
  reg [7:0] p76_array_index_2058096;
  reg [7:0] p76_array_index_2058097;
  reg [7:0] p76_array_index_2058098;
  reg [7:0] p76_res7__1027;
  reg [7:0] p76_res7__994;
  reg [7:0] p76_array_index_2058115;
  reg [7:0] p76_array_index_2058116;
  reg [7:0] p76_array_index_2058117;
  reg [7:0] p76_array_index_2058118;
  reg [7:0] p76_array_index_2058119;
  reg [7:0] p76_array_index_2058122;
  reg [7:0] p76_array_index_2058123;
  reg [7:0] p76_array_index_2058124;
  reg [7:0] p76_array_index_2058125;
  reg [7:0] p76_array_index_2058126;
  reg [7:0] p76_res7__1029;
  reg [7:0] p76_res7__996;
  reg [7:0] p76_array_index_2058143;
  reg [7:0] p76_array_index_2058144;
  reg [7:0] p76_array_index_2058145;
  reg [7:0] p76_array_index_2058146;
  reg [7:0] p76_array_index_2058147;
  reg [7:0] p76_array_index_2058150;
  reg [7:0] p76_array_index_2058151;
  reg [7:0] p76_array_index_2058152;
  reg [7:0] p76_array_index_2058153;
  reg [7:0] p76_array_index_2058154;
  reg [7:0] p76_res7__1031;
  reg [7:0] p76_res7__998;
  reg [7:0] p76_array_index_2058164;
  reg [7:0] p76_array_index_2058165;
  reg [7:0] p76_array_index_2058166;
  reg [7:0] p76_array_index_2058167;
  reg [7:0] p76_array_index_2058168;
  reg [7:0] p76_array_index_2058169;
  reg [7:0] p76_array_index_2058170;
  reg [7:0] p76_array_index_2058171;
  reg [7:0] p76_array_index_2058172;
  reg [7:0] p76_array_index_2058173;
  reg [7:0] p76_array_index_2058174;
  reg [7:0] p76_array_index_2058175;
  reg [7:0] p77_literal_2043910[256];
  reg [7:0] p77_literal_2043912[256];
  reg [7:0] p77_literal_2043914[256];
  reg [7:0] p77_literal_2043916[256];
  reg [7:0] p77_literal_2043918[256];
  reg [7:0] p77_literal_2043920[256];
  reg [7:0] p77_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p76_bit_slice_2043893 <= p75_bit_slice_2043893;
    p76_bit_slice_2044018 <= p75_bit_slice_2044018;
    p76_k3 <= p75_k3;
    p76_k2 <= p75_k2;
    p76_k5 <= p75_k5;
    p76_k4 <= p75_k4;
    p76_k7 <= p75_k7;
    p76_k6 <= p75_k6;
    p76_xor_2057490 <= p75_xor_2057490;
    p76_bit_slice_2058020 <= p76_bit_slice_2058020_comb;
    p76_bit_slice_2058021 <= p76_bit_slice_2058021_comb;
    p76_bit_slice_2058022 <= p76_bit_slice_2058022_comb;
    p76_bit_slice_2058023 <= p76_bit_slice_2058023_comb;
    p76_bit_slice_2058024 <= p76_bit_slice_2058024_comb;
    p76_bit_slice_2058025 <= p76_bit_slice_2058025_comb;
    p76_bit_slice_2058026 <= p76_bit_slice_2058026_comb;
    p76_bit_slice_2058027 <= p76_bit_slice_2058027_comb;
    p76_bit_slice_2058028 <= p76_bit_slice_2058028_comb;
    p76_bit_slice_2058029 <= p76_bit_slice_2058029_comb;
    p76_array_index_2058030 <= p76_array_index_2058030_comb;
    p76_array_index_2058031 <= p76_array_index_2058031_comb;
    p76_array_index_2058032 <= p76_array_index_2058032_comb;
    p76_array_index_2058033 <= p76_array_index_2058033_comb;
    p76_array_index_2058034 <= p76_array_index_2058034_comb;
    p76_array_index_2058035 <= p76_array_index_2058035_comb;
    p76_array_index_2058037 <= p76_array_index_2058037_comb;
    p76_array_index_2058039 <= p76_array_index_2058039_comb;
    p76_array_index_2058040 <= p76_array_index_2058040_comb;
    p76_array_index_2058041 <= p76_array_index_2058041_comb;
    p76_bit_slice_2058052 <= p76_bit_slice_2058052_comb;
    p76_bit_slice_2058054 <= p76_bit_slice_2058054_comb;
    p76_array_index_2058055 <= p76_array_index_2058055_comb;
    p76_array_index_2058056 <= p76_array_index_2058056_comb;
    p76_array_index_2058057 <= p76_array_index_2058057_comb;
    p76_array_index_2058058 <= p76_array_index_2058058_comb;
    p76_array_index_2058059 <= p76_array_index_2058059_comb;
    p76_array_index_2058060 <= p76_array_index_2058060_comb;
    p76_array_index_2058062 <= p76_array_index_2058062_comb;
    p76_array_index_2058063 <= p76_array_index_2058063_comb;
    p76_array_index_2058064 <= p76_array_index_2058064_comb;
    p76_array_index_2058065 <= p76_array_index_2058065_comb;
    p76_array_index_2058066 <= p76_array_index_2058066_comb;
    p76_array_index_2058067 <= p76_array_index_2058067_comb;
    p76_array_index_2058068 <= p76_array_index_2058068_comb;
    p76_array_index_2058070 <= p76_array_index_2058070_comb;
    p76_res7__1025 <= p76_res7__1025_comb;
    p76_res7__992 <= p76_res7__992_comb;
    p76_array_index_2058087 <= p76_array_index_2058087_comb;
    p76_array_index_2058088 <= p76_array_index_2058088_comb;
    p76_array_index_2058089 <= p76_array_index_2058089_comb;
    p76_array_index_2058090 <= p76_array_index_2058090_comb;
    p76_array_index_2058091 <= p76_array_index_2058091_comb;
    p76_array_index_2058092 <= p76_array_index_2058092_comb;
    p76_array_index_2058093 <= p76_array_index_2058093_comb;
    p76_array_index_2058094 <= p76_array_index_2058094_comb;
    p76_array_index_2058095 <= p76_array_index_2058095_comb;
    p76_array_index_2058096 <= p76_array_index_2058096_comb;
    p76_array_index_2058097 <= p76_array_index_2058097_comb;
    p76_array_index_2058098 <= p76_array_index_2058098_comb;
    p76_res7__1027 <= p76_res7__1027_comb;
    p76_res7__994 <= p76_res7__994_comb;
    p76_array_index_2058115 <= p76_array_index_2058115_comb;
    p76_array_index_2058116 <= p76_array_index_2058116_comb;
    p76_array_index_2058117 <= p76_array_index_2058117_comb;
    p76_array_index_2058118 <= p76_array_index_2058118_comb;
    p76_array_index_2058119 <= p76_array_index_2058119_comb;
    p76_array_index_2058122 <= p76_array_index_2058122_comb;
    p76_array_index_2058123 <= p76_array_index_2058123_comb;
    p76_array_index_2058124 <= p76_array_index_2058124_comb;
    p76_array_index_2058125 <= p76_array_index_2058125_comb;
    p76_array_index_2058126 <= p76_array_index_2058126_comb;
    p76_res7__1029 <= p76_res7__1029_comb;
    p76_res7__996 <= p76_res7__996_comb;
    p76_array_index_2058143 <= p76_array_index_2058143_comb;
    p76_array_index_2058144 <= p76_array_index_2058144_comb;
    p76_array_index_2058145 <= p76_array_index_2058145_comb;
    p76_array_index_2058146 <= p76_array_index_2058146_comb;
    p76_array_index_2058147 <= p76_array_index_2058147_comb;
    p76_array_index_2058150 <= p76_array_index_2058150_comb;
    p76_array_index_2058151 <= p76_array_index_2058151_comb;
    p76_array_index_2058152 <= p76_array_index_2058152_comb;
    p76_array_index_2058153 <= p76_array_index_2058153_comb;
    p76_array_index_2058154 <= p76_array_index_2058154_comb;
    p76_res7__1031 <= p76_res7__1031_comb;
    p76_res7__998 <= p76_res7__998_comb;
    p76_array_index_2058164 <= p76_array_index_2058164_comb;
    p76_array_index_2058165 <= p76_array_index_2058165_comb;
    p76_array_index_2058166 <= p76_array_index_2058166_comb;
    p76_array_index_2058167 <= p76_array_index_2058167_comb;
    p76_array_index_2058168 <= p76_array_index_2058168_comb;
    p76_array_index_2058169 <= p76_array_index_2058169_comb;
    p76_array_index_2058170 <= p76_array_index_2058170_comb;
    p76_array_index_2058171 <= p76_array_index_2058171_comb;
    p76_array_index_2058172 <= p76_array_index_2058172_comb;
    p76_array_index_2058173 <= p76_array_index_2058173_comb;
    p76_array_index_2058174 <= p76_array_index_2058174_comb;
    p76_array_index_2058175 <= p76_array_index_2058175_comb;
    p77_literal_2043910 <= p76_literal_2043910;
    p77_literal_2043912 <= p76_literal_2043912;
    p77_literal_2043914 <= p76_literal_2043914;
    p77_literal_2043916 <= p76_literal_2043916;
    p77_literal_2043918 <= p76_literal_2043918;
    p77_literal_2043920 <= p76_literal_2043920;
    p77_literal_2043923 <= p76_literal_2043923;
  end

  // ===== Pipe stage 77:
  wire [7:0] p77_array_index_2058386_comb;
  wire [7:0] p77_array_index_2058387_comb;
  wire [7:0] p77_array_index_2058388_comb;
  wire [7:0] p77_array_index_2058389_comb;
  wire [7:0] p77_res7__1033_comb;
  wire [7:0] p77_res7__1000_comb;
  wire [7:0] p77_array_index_2058404_comb;
  wire [7:0] p77_array_index_2058405_comb;
  wire [7:0] p77_array_index_2058406_comb;
  wire [7:0] p77_array_index_2058407_comb;
  wire [7:0] p77_array_index_2058412_comb;
  wire [7:0] p77_array_index_2058413_comb;
  wire [7:0] p77_array_index_2058414_comb;
  wire [7:0] p77_array_index_2058415_comb;
  wire [7:0] p77_res7__1035_comb;
  wire [7:0] p77_res7__1002_comb;
  wire [7:0] p77_array_index_2058429_comb;
  wire [7:0] p77_array_index_2058430_comb;
  wire [7:0] p77_array_index_2058431_comb;
  wire [7:0] p77_array_index_2058438_comb;
  wire [7:0] p77_array_index_2058439_comb;
  wire [7:0] p77_array_index_2058440_comb;
  wire [7:0] p77_res7__1037_comb;
  wire [7:0] p77_res7__1004_comb;
  wire [7:0] p77_array_index_2058453_comb;
  wire [7:0] p77_array_index_2058454_comb;
  wire [7:0] p77_array_index_2058455_comb;
  wire [7:0] p77_array_index_2058462_comb;
  wire [7:0] p77_array_index_2058463_comb;
  wire [7:0] p77_array_index_2058464_comb;
  wire [7:0] p77_res7__1039_comb;
  wire [7:0] p77_res7__1006_comb;
  wire [7:0] p77_array_index_2058476_comb;
  wire [7:0] p77_array_index_2058477_comb;
  wire [7:0] p77_array_index_2058486_comb;
  wire [7:0] p77_array_index_2058487_comb;
  wire [7:0] p77_res7__1041_comb;
  wire [7:0] p77_res7__1008_comb;
  wire [7:0] p77_array_index_2058498_comb;
  wire [7:0] p77_array_index_2058499_comb;
  wire [7:0] p77_array_index_2058508_comb;
  wire [7:0] p77_array_index_2058509_comb;
  wire [7:0] p77_res7__1043_comb;
  wire [7:0] p77_res7__1010_comb;
  wire [7:0] p77_array_index_2058519_comb;
  wire [7:0] p77_array_index_2058530_comb;
  wire [7:0] p77_res7__1045_comb;
  wire [7:0] p77_res7__1012_comb;
  wire [7:0] p77_array_index_2058536_comb;
  wire [7:0] p77_array_index_2058537_comb;
  wire [7:0] p77_array_index_2058538_comb;
  wire [7:0] p77_array_index_2058539_comb;
  wire [7:0] p77_array_index_2058540_comb;
  wire [7:0] p77_array_index_2058541_comb;
  wire [7:0] p77_array_index_2058542_comb;
  wire [7:0] p77_array_index_2058543_comb;
  wire [7:0] p77_array_index_2058544_comb;
  assign p77_array_index_2058386_comb = p76_literal_2043914[p76_res7__994];
  assign p77_array_index_2058387_comb = p76_literal_2043916[p76_res7__992];
  assign p77_array_index_2058388_comb = p76_literal_2043918[p76_array_index_2058030];
  assign p77_array_index_2058389_comb = p76_literal_2043920[p76_array_index_2058031];
  assign p77_res7__1033_comb = p76_array_index_2058164 ^ p76_array_index_2058165 ^ p76_array_index_2058166 ^ p76_array_index_2058167 ^ p76_array_index_2058168 ^ p76_array_index_2058055 ^ p76_bit_slice_2058025 ^ p76_array_index_2058169 ^ p76_bit_slice_2058027 ^ p76_array_index_2058170 ^ p76_array_index_2058171 ^ p76_array_index_2058172 ^ p76_array_index_2058173 ^ p76_array_index_2058174 ^ p76_array_index_2058175 ^ p76_bit_slice_2058020;
  assign p77_res7__1000_comb = p76_literal_2043910[p76_res7__998] ^ p76_literal_2043912[p76_res7__996] ^ p77_array_index_2058386_comb ^ p77_array_index_2058387_comb ^ p77_array_index_2058388_comb ^ p77_array_index_2058389_comb ^ p76_array_index_2058032 ^ p76_literal_2043923[p76_array_index_2058033] ^ p76_array_index_2058034 ^ p76_array_index_2058067 ^ p76_literal_2043918[p76_array_index_2058068] ^ p76_literal_2043916[p76_array_index_2058037] ^ p76_literal_2043914[p76_array_index_2058070] ^ p76_literal_2043912[p76_array_index_2058039] ^ p76_literal_2043910[p76_array_index_2058040] ^ p76_array_index_2058041;
  assign p77_array_index_2058404_comb = p76_literal_2043920[p76_bit_slice_2058029];
  assign p77_array_index_2058405_comb = p76_literal_2043918[p76_res7__1025];
  assign p77_array_index_2058406_comb = p76_literal_2043916[p76_res7__1027];
  assign p77_array_index_2058407_comb = p76_literal_2043914[p76_res7__1029];
  assign p77_array_index_2058412_comb = p76_literal_2043914[p76_res7__996];
  assign p77_array_index_2058413_comb = p76_literal_2043916[p76_res7__994];
  assign p77_array_index_2058414_comb = p76_literal_2043918[p76_res7__992];
  assign p77_array_index_2058415_comb = p76_literal_2043920[p76_array_index_2058030];
  assign p77_res7__1035_comb = p76_literal_2043910[p76_bit_slice_2058022] ^ p76_literal_2043912[p76_bit_slice_2058052] ^ p76_literal_2043914[p76_bit_slice_2058023] ^ p76_literal_2043916[p76_bit_slice_2058054] ^ p76_literal_2043918[p76_bit_slice_2058024] ^ p76_array_index_2058087 ^ p76_bit_slice_2058026 ^ p76_literal_2043923[p76_bit_slice_2058027] ^ p76_bit_slice_2058028 ^ p77_array_index_2058404_comb ^ p77_array_index_2058405_comb ^ p77_array_index_2058406_comb ^ p77_array_index_2058407_comb ^ p76_literal_2043912[p76_res7__1031] ^ p76_literal_2043910[p77_res7__1033_comb] ^ p76_bit_slice_2058021;
  assign p77_res7__1002_comb = p76_literal_2043910[p77_res7__1000_comb] ^ p76_literal_2043912[p76_res7__998] ^ p77_array_index_2058412_comb ^ p77_array_index_2058413_comb ^ p77_array_index_2058414_comb ^ p77_array_index_2058415_comb ^ p76_array_index_2058031 ^ p76_literal_2043923[p76_array_index_2058032] ^ p76_array_index_2058033 ^ p76_array_index_2058098 ^ p76_literal_2043918[p76_array_index_2058035] ^ p76_literal_2043916[p76_array_index_2058068] ^ p76_literal_2043914[p76_array_index_2058037] ^ p76_literal_2043912[p76_array_index_2058070] ^ p76_literal_2043910[p76_array_index_2058039] ^ p76_array_index_2058040;
  assign p77_array_index_2058429_comb = p76_literal_2043920[p76_res7__1025];
  assign p77_array_index_2058430_comb = p76_literal_2043918[p76_res7__1027];
  assign p77_array_index_2058431_comb = p76_literal_2043916[p76_res7__1029];
  assign p77_array_index_2058438_comb = p76_literal_2043916[p76_res7__996];
  assign p77_array_index_2058439_comb = p76_literal_2043918[p76_res7__994];
  assign p77_array_index_2058440_comb = p76_literal_2043920[p76_res7__992];
  assign p77_res7__1037_comb = p76_literal_2043910[p76_bit_slice_2058052] ^ p76_literal_2043912[p76_bit_slice_2058023] ^ p76_literal_2043914[p76_bit_slice_2058054] ^ p76_literal_2043916[p76_bit_slice_2058024] ^ p76_array_index_2058056 ^ p76_array_index_2058115 ^ p76_bit_slice_2058027 ^ p76_literal_2043923[p76_bit_slice_2058028] ^ p76_bit_slice_2058029 ^ p77_array_index_2058429_comb ^ p77_array_index_2058430_comb ^ p77_array_index_2058431_comb ^ p76_literal_2043914[p76_res7__1031] ^ p76_literal_2043912[p77_res7__1033_comb] ^ p76_literal_2043910[p77_res7__1035_comb] ^ p76_bit_slice_2058022;
  assign p77_res7__1004_comb = p76_literal_2043910[p77_res7__1002_comb] ^ p76_literal_2043912[p77_res7__1000_comb] ^ p76_literal_2043914[p76_res7__998] ^ p77_array_index_2058438_comb ^ p77_array_index_2058439_comb ^ p77_array_index_2058440_comb ^ p76_array_index_2058030 ^ p76_literal_2043923[p76_array_index_2058031] ^ p76_array_index_2058032 ^ p76_array_index_2058126 ^ p76_array_index_2058066 ^ p76_literal_2043916[p76_array_index_2058035] ^ p76_literal_2043914[p76_array_index_2058068] ^ p76_literal_2043912[p76_array_index_2058037] ^ p76_literal_2043910[p76_array_index_2058070] ^ p76_array_index_2058039;
  assign p77_array_index_2058453_comb = p76_literal_2043920[p76_res7__1027];
  assign p77_array_index_2058454_comb = p76_literal_2043918[p76_res7__1029];
  assign p77_array_index_2058455_comb = p76_literal_2043916[p76_res7__1031];
  assign p77_array_index_2058462_comb = p76_literal_2043916[p76_res7__998];
  assign p77_array_index_2058463_comb = p76_literal_2043918[p76_res7__996];
  assign p77_array_index_2058464_comb = p76_literal_2043920[p76_res7__994];
  assign p77_res7__1039_comb = p76_literal_2043910[p76_bit_slice_2058023] ^ p76_literal_2043912[p76_bit_slice_2058054] ^ p76_literal_2043914[p76_bit_slice_2058024] ^ p76_literal_2043916[p76_bit_slice_2058025] ^ p76_array_index_2058088 ^ p76_array_index_2058143 ^ p76_bit_slice_2058028 ^ p76_literal_2043923[p76_bit_slice_2058029] ^ p76_res7__1025 ^ p77_array_index_2058453_comb ^ p77_array_index_2058454_comb ^ p77_array_index_2058455_comb ^ p76_literal_2043914[p77_res7__1033_comb] ^ p76_literal_2043912[p77_res7__1035_comb] ^ p76_literal_2043910[p77_res7__1037_comb] ^ p76_bit_slice_2058052;
  assign p77_res7__1006_comb = p76_literal_2043910[p77_res7__1004_comb] ^ p76_literal_2043912[p77_res7__1002_comb] ^ p76_literal_2043914[p77_res7__1000_comb] ^ p77_array_index_2058462_comb ^ p77_array_index_2058463_comb ^ p77_array_index_2058464_comb ^ p76_res7__992 ^ p76_literal_2043923[p76_array_index_2058030] ^ p76_array_index_2058031 ^ p76_array_index_2058154 ^ p76_array_index_2058097 ^ p76_literal_2043916[p76_array_index_2058034] ^ p76_literal_2043914[p76_array_index_2058035] ^ p76_literal_2043912[p76_array_index_2058068] ^ p76_literal_2043910[p76_array_index_2058037] ^ p76_array_index_2058070;
  assign p77_array_index_2058476_comb = p76_literal_2043920[p76_res7__1029];
  assign p77_array_index_2058477_comb = p76_literal_2043918[p76_res7__1031];
  assign p77_array_index_2058486_comb = p76_literal_2043918[p76_res7__998];
  assign p77_array_index_2058487_comb = p76_literal_2043920[p76_res7__996];
  assign p77_res7__1041_comb = p76_literal_2043910[p76_bit_slice_2058054] ^ p76_literal_2043912[p76_bit_slice_2058024] ^ p76_literal_2043914[p76_bit_slice_2058025] ^ p76_array_index_2058057 ^ p76_array_index_2058116 ^ p76_array_index_2058170 ^ p76_bit_slice_2058029 ^ p76_literal_2043923[p76_res7__1025] ^ p76_res7__1027 ^ p77_array_index_2058476_comb ^ p77_array_index_2058477_comb ^ p76_literal_2043916[p77_res7__1033_comb] ^ p76_literal_2043914[p77_res7__1035_comb] ^ p76_literal_2043912[p77_res7__1037_comb] ^ p76_literal_2043910[p77_res7__1039_comb] ^ p76_bit_slice_2058023;
  assign p77_res7__1008_comb = p76_literal_2043910[p77_res7__1006_comb] ^ p76_literal_2043912[p77_res7__1004_comb] ^ p76_literal_2043914[p77_res7__1002_comb] ^ p76_literal_2043916[p77_res7__1000_comb] ^ p77_array_index_2058486_comb ^ p77_array_index_2058487_comb ^ p76_res7__994 ^ p76_literal_2043923[p76_res7__992] ^ p76_array_index_2058030 ^ p77_array_index_2058389_comb ^ p76_array_index_2058125 ^ p76_array_index_2058065 ^ p76_literal_2043914[p76_array_index_2058034] ^ p76_literal_2043912[p76_array_index_2058035] ^ p76_literal_2043910[p76_array_index_2058068] ^ p76_array_index_2058037;
  assign p77_array_index_2058498_comb = p76_literal_2043920[p76_res7__1031];
  assign p77_array_index_2058499_comb = p76_literal_2043918[p77_res7__1033_comb];
  assign p77_array_index_2058508_comb = p76_literal_2043918[p77_res7__1000_comb];
  assign p77_array_index_2058509_comb = p76_literal_2043920[p76_res7__998];
  assign p77_res7__1043_comb = p76_literal_2043910[p76_bit_slice_2058024] ^ p76_literal_2043912[p76_bit_slice_2058025] ^ p76_literal_2043914[p76_bit_slice_2058026] ^ p76_array_index_2058089 ^ p76_array_index_2058144 ^ p77_array_index_2058404_comb ^ p76_res7__1025 ^ p76_literal_2043923[p76_res7__1027] ^ p76_res7__1029 ^ p77_array_index_2058498_comb ^ p77_array_index_2058499_comb ^ p76_literal_2043916[p77_res7__1035_comb] ^ p76_literal_2043914[p77_res7__1037_comb] ^ p76_literal_2043912[p77_res7__1039_comb] ^ p76_literal_2043910[p77_res7__1041_comb] ^ p76_bit_slice_2058054;
  assign p77_res7__1010_comb = p76_literal_2043910[p77_res7__1008_comb] ^ p76_literal_2043912[p77_res7__1006_comb] ^ p76_literal_2043914[p77_res7__1004_comb] ^ p76_literal_2043916[p77_res7__1002_comb] ^ p77_array_index_2058508_comb ^ p77_array_index_2058509_comb ^ p76_res7__996 ^ p76_literal_2043923[p76_res7__994] ^ p76_res7__992 ^ p77_array_index_2058415_comb ^ p76_array_index_2058153 ^ p76_array_index_2058096 ^ p76_literal_2043914[p76_array_index_2058033] ^ p76_literal_2043912[p76_array_index_2058034] ^ p76_literal_2043910[p76_array_index_2058035] ^ p76_array_index_2058068;
  assign p77_array_index_2058519_comb = p76_literal_2043920[p77_res7__1033_comb];
  assign p77_array_index_2058530_comb = p76_literal_2043920[p77_res7__1000_comb];
  assign p77_res7__1045_comb = p76_literal_2043910[p76_bit_slice_2058025] ^ p76_literal_2043912[p76_bit_slice_2058026] ^ p76_array_index_2058058 ^ p76_array_index_2058117 ^ p76_array_index_2058171 ^ p77_array_index_2058429_comb ^ p76_res7__1027 ^ p76_literal_2043923[p76_res7__1029] ^ p76_res7__1031 ^ p77_array_index_2058519_comb ^ p76_literal_2043918[p77_res7__1035_comb] ^ p76_literal_2043916[p77_res7__1037_comb] ^ p76_literal_2043914[p77_res7__1039_comb] ^ p76_literal_2043912[p77_res7__1041_comb] ^ p76_literal_2043910[p77_res7__1043_comb] ^ p76_bit_slice_2058024;
  assign p77_res7__1012_comb = p76_literal_2043910[p77_res7__1010_comb] ^ p76_literal_2043912[p77_res7__1008_comb] ^ p76_literal_2043914[p77_res7__1006_comb] ^ p76_literal_2043916[p77_res7__1004_comb] ^ p76_literal_2043918[p77_res7__1002_comb] ^ p77_array_index_2058530_comb ^ p76_res7__998 ^ p76_literal_2043923[p76_res7__996] ^ p76_res7__994 ^ p77_array_index_2058440_comb ^ p77_array_index_2058388_comb ^ p76_array_index_2058124 ^ p76_array_index_2058064 ^ p76_literal_2043912[p76_array_index_2058033] ^ p76_literal_2043910[p76_array_index_2058034] ^ p76_array_index_2058035;
  assign p77_array_index_2058536_comb = p76_literal_2043910[p76_bit_slice_2058026];
  assign p77_array_index_2058537_comb = p76_literal_2043912[p76_bit_slice_2058027];
  assign p77_array_index_2058538_comb = p76_literal_2043923[p76_res7__1031];
  assign p77_array_index_2058539_comb = p76_literal_2043920[p77_res7__1035_comb];
  assign p77_array_index_2058540_comb = p76_literal_2043918[p77_res7__1037_comb];
  assign p77_array_index_2058541_comb = p76_literal_2043916[p77_res7__1039_comb];
  assign p77_array_index_2058542_comb = p76_literal_2043914[p77_res7__1041_comb];
  assign p77_array_index_2058543_comb = p76_literal_2043912[p77_res7__1043_comb];
  assign p77_array_index_2058544_comb = p76_literal_2043910[p77_res7__1045_comb];

  // Registers for pipe stage 77:
  reg [127:0] p77_bit_slice_2043893;
  reg [127:0] p77_bit_slice_2044018;
  reg [127:0] p77_k3;
  reg [127:0] p77_k2;
  reg [127:0] p77_k5;
  reg [127:0] p77_k4;
  reg [127:0] p77_k7;
  reg [127:0] p77_k6;
  reg [127:0] p77_xor_2057490;
  reg [7:0] p77_bit_slice_2058025;
  reg [7:0] p77_bit_slice_2058026;
  reg [7:0] p77_bit_slice_2058027;
  reg [7:0] p77_bit_slice_2058028;
  reg [7:0] p77_bit_slice_2058029;
  reg [7:0] p77_array_index_2058030;
  reg [7:0] p77_array_index_2058031;
  reg [7:0] p77_array_index_2058032;
  reg [7:0] p77_array_index_2058033;
  reg [7:0] p77_array_index_2058034;
  reg [7:0] p77_array_index_2058059;
  reg [7:0] p77_array_index_2058060;
  reg [7:0] p77_array_index_2058062;
  reg [7:0] p77_array_index_2058063;
  reg [7:0] p77_res7__1025;
  reg [7:0] p77_res7__992;
  reg [7:0] p77_array_index_2058090;
  reg [7:0] p77_array_index_2058091;
  reg [7:0] p77_array_index_2058092;
  reg [7:0] p77_array_index_2058093;
  reg [7:0] p77_array_index_2058094;
  reg [7:0] p77_array_index_2058095;
  reg [7:0] p77_res7__1027;
  reg [7:0] p77_res7__994;
  reg [7:0] p77_array_index_2058118;
  reg [7:0] p77_array_index_2058119;
  reg [7:0] p77_array_index_2058122;
  reg [7:0] p77_array_index_2058123;
  reg [7:0] p77_res7__1029;
  reg [7:0] p77_res7__996;
  reg [7:0] p77_array_index_2058145;
  reg [7:0] p77_array_index_2058146;
  reg [7:0] p77_array_index_2058147;
  reg [7:0] p77_array_index_2058150;
  reg [7:0] p77_array_index_2058151;
  reg [7:0] p77_array_index_2058152;
  reg [7:0] p77_res7__1031;
  reg [7:0] p77_res7__998;
  reg [7:0] p77_array_index_2058172;
  reg [7:0] p77_array_index_2058173;
  reg [7:0] p77_array_index_2058386;
  reg [7:0] p77_array_index_2058387;
  reg [7:0] p77_res7__1033;
  reg [7:0] p77_res7__1000;
  reg [7:0] p77_array_index_2058405;
  reg [7:0] p77_array_index_2058406;
  reg [7:0] p77_array_index_2058407;
  reg [7:0] p77_array_index_2058412;
  reg [7:0] p77_array_index_2058413;
  reg [7:0] p77_array_index_2058414;
  reg [7:0] p77_res7__1035;
  reg [7:0] p77_res7__1002;
  reg [7:0] p77_array_index_2058430;
  reg [7:0] p77_array_index_2058431;
  reg [7:0] p77_array_index_2058438;
  reg [7:0] p77_array_index_2058439;
  reg [7:0] p77_res7__1037;
  reg [7:0] p77_res7__1004;
  reg [7:0] p77_array_index_2058453;
  reg [7:0] p77_array_index_2058454;
  reg [7:0] p77_array_index_2058455;
  reg [7:0] p77_array_index_2058462;
  reg [7:0] p77_array_index_2058463;
  reg [7:0] p77_array_index_2058464;
  reg [7:0] p77_res7__1039;
  reg [7:0] p77_res7__1006;
  reg [7:0] p77_array_index_2058476;
  reg [7:0] p77_array_index_2058477;
  reg [7:0] p77_array_index_2058486;
  reg [7:0] p77_array_index_2058487;
  reg [7:0] p77_res7__1041;
  reg [7:0] p77_res7__1008;
  reg [7:0] p77_array_index_2058498;
  reg [7:0] p77_array_index_2058499;
  reg [7:0] p77_array_index_2058508;
  reg [7:0] p77_array_index_2058509;
  reg [7:0] p77_res7__1043;
  reg [7:0] p77_res7__1010;
  reg [7:0] p77_array_index_2058519;
  reg [7:0] p77_array_index_2058530;
  reg [7:0] p77_res7__1045;
  reg [7:0] p77_res7__1012;
  reg [7:0] p77_array_index_2058536;
  reg [7:0] p77_array_index_2058537;
  reg [7:0] p77_array_index_2058538;
  reg [7:0] p77_array_index_2058539;
  reg [7:0] p77_array_index_2058540;
  reg [7:0] p77_array_index_2058541;
  reg [7:0] p77_array_index_2058542;
  reg [7:0] p77_array_index_2058543;
  reg [7:0] p77_array_index_2058544;
  reg [7:0] p78_literal_2043910[256];
  reg [7:0] p78_literal_2043912[256];
  reg [7:0] p78_literal_2043914[256];
  reg [7:0] p78_literal_2043916[256];
  reg [7:0] p78_literal_2043918[256];
  reg [7:0] p78_literal_2043920[256];
  reg [7:0] p78_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p77_bit_slice_2043893 <= p76_bit_slice_2043893;
    p77_bit_slice_2044018 <= p76_bit_slice_2044018;
    p77_k3 <= p76_k3;
    p77_k2 <= p76_k2;
    p77_k5 <= p76_k5;
    p77_k4 <= p76_k4;
    p77_k7 <= p76_k7;
    p77_k6 <= p76_k6;
    p77_xor_2057490 <= p76_xor_2057490;
    p77_bit_slice_2058025 <= p76_bit_slice_2058025;
    p77_bit_slice_2058026 <= p76_bit_slice_2058026;
    p77_bit_slice_2058027 <= p76_bit_slice_2058027;
    p77_bit_slice_2058028 <= p76_bit_slice_2058028;
    p77_bit_slice_2058029 <= p76_bit_slice_2058029;
    p77_array_index_2058030 <= p76_array_index_2058030;
    p77_array_index_2058031 <= p76_array_index_2058031;
    p77_array_index_2058032 <= p76_array_index_2058032;
    p77_array_index_2058033 <= p76_array_index_2058033;
    p77_array_index_2058034 <= p76_array_index_2058034;
    p77_array_index_2058059 <= p76_array_index_2058059;
    p77_array_index_2058060 <= p76_array_index_2058060;
    p77_array_index_2058062 <= p76_array_index_2058062;
    p77_array_index_2058063 <= p76_array_index_2058063;
    p77_res7__1025 <= p76_res7__1025;
    p77_res7__992 <= p76_res7__992;
    p77_array_index_2058090 <= p76_array_index_2058090;
    p77_array_index_2058091 <= p76_array_index_2058091;
    p77_array_index_2058092 <= p76_array_index_2058092;
    p77_array_index_2058093 <= p76_array_index_2058093;
    p77_array_index_2058094 <= p76_array_index_2058094;
    p77_array_index_2058095 <= p76_array_index_2058095;
    p77_res7__1027 <= p76_res7__1027;
    p77_res7__994 <= p76_res7__994;
    p77_array_index_2058118 <= p76_array_index_2058118;
    p77_array_index_2058119 <= p76_array_index_2058119;
    p77_array_index_2058122 <= p76_array_index_2058122;
    p77_array_index_2058123 <= p76_array_index_2058123;
    p77_res7__1029 <= p76_res7__1029;
    p77_res7__996 <= p76_res7__996;
    p77_array_index_2058145 <= p76_array_index_2058145;
    p77_array_index_2058146 <= p76_array_index_2058146;
    p77_array_index_2058147 <= p76_array_index_2058147;
    p77_array_index_2058150 <= p76_array_index_2058150;
    p77_array_index_2058151 <= p76_array_index_2058151;
    p77_array_index_2058152 <= p76_array_index_2058152;
    p77_res7__1031 <= p76_res7__1031;
    p77_res7__998 <= p76_res7__998;
    p77_array_index_2058172 <= p76_array_index_2058172;
    p77_array_index_2058173 <= p76_array_index_2058173;
    p77_array_index_2058386 <= p77_array_index_2058386_comb;
    p77_array_index_2058387 <= p77_array_index_2058387_comb;
    p77_res7__1033 <= p77_res7__1033_comb;
    p77_res7__1000 <= p77_res7__1000_comb;
    p77_array_index_2058405 <= p77_array_index_2058405_comb;
    p77_array_index_2058406 <= p77_array_index_2058406_comb;
    p77_array_index_2058407 <= p77_array_index_2058407_comb;
    p77_array_index_2058412 <= p77_array_index_2058412_comb;
    p77_array_index_2058413 <= p77_array_index_2058413_comb;
    p77_array_index_2058414 <= p77_array_index_2058414_comb;
    p77_res7__1035 <= p77_res7__1035_comb;
    p77_res7__1002 <= p77_res7__1002_comb;
    p77_array_index_2058430 <= p77_array_index_2058430_comb;
    p77_array_index_2058431 <= p77_array_index_2058431_comb;
    p77_array_index_2058438 <= p77_array_index_2058438_comb;
    p77_array_index_2058439 <= p77_array_index_2058439_comb;
    p77_res7__1037 <= p77_res7__1037_comb;
    p77_res7__1004 <= p77_res7__1004_comb;
    p77_array_index_2058453 <= p77_array_index_2058453_comb;
    p77_array_index_2058454 <= p77_array_index_2058454_comb;
    p77_array_index_2058455 <= p77_array_index_2058455_comb;
    p77_array_index_2058462 <= p77_array_index_2058462_comb;
    p77_array_index_2058463 <= p77_array_index_2058463_comb;
    p77_array_index_2058464 <= p77_array_index_2058464_comb;
    p77_res7__1039 <= p77_res7__1039_comb;
    p77_res7__1006 <= p77_res7__1006_comb;
    p77_array_index_2058476 <= p77_array_index_2058476_comb;
    p77_array_index_2058477 <= p77_array_index_2058477_comb;
    p77_array_index_2058486 <= p77_array_index_2058486_comb;
    p77_array_index_2058487 <= p77_array_index_2058487_comb;
    p77_res7__1041 <= p77_res7__1041_comb;
    p77_res7__1008 <= p77_res7__1008_comb;
    p77_array_index_2058498 <= p77_array_index_2058498_comb;
    p77_array_index_2058499 <= p77_array_index_2058499_comb;
    p77_array_index_2058508 <= p77_array_index_2058508_comb;
    p77_array_index_2058509 <= p77_array_index_2058509_comb;
    p77_res7__1043 <= p77_res7__1043_comb;
    p77_res7__1010 <= p77_res7__1010_comb;
    p77_array_index_2058519 <= p77_array_index_2058519_comb;
    p77_array_index_2058530 <= p77_array_index_2058530_comb;
    p77_res7__1045 <= p77_res7__1045_comb;
    p77_res7__1012 <= p77_res7__1012_comb;
    p77_array_index_2058536 <= p77_array_index_2058536_comb;
    p77_array_index_2058537 <= p77_array_index_2058537_comb;
    p77_array_index_2058538 <= p77_array_index_2058538_comb;
    p77_array_index_2058539 <= p77_array_index_2058539_comb;
    p77_array_index_2058540 <= p77_array_index_2058540_comb;
    p77_array_index_2058541 <= p77_array_index_2058541_comb;
    p77_array_index_2058542 <= p77_array_index_2058542_comb;
    p77_array_index_2058543 <= p77_array_index_2058543_comb;
    p77_array_index_2058544 <= p77_array_index_2058544_comb;
    p78_literal_2043910 <= p77_literal_2043910;
    p78_literal_2043912 <= p77_literal_2043912;
    p78_literal_2043914 <= p77_literal_2043914;
    p78_literal_2043916 <= p77_literal_2043916;
    p78_literal_2043918 <= p77_literal_2043918;
    p78_literal_2043920 <= p77_literal_2043920;
    p78_literal_2043923 <= p77_literal_2043923;
  end

  // ===== Pipe stage 78:
  wire [7:0] p78_array_index_2058764_comb;
  wire [7:0] p78_res7__1047_comb;
  wire [7:0] p78_res7__1014_comb;
  wire [7:0] p78_res7__1049_comb;
  wire [7:0] p78_res7__1016_comb;
  wire [7:0] p78_res7__1051_comb;
  wire [7:0] p78_res7__1018_comb;
  wire [7:0] p78_res7__1053_comb;
  wire [7:0] p78_res7__1020_comb;
  wire [7:0] p78_res7__1055_comb;
  wire [7:0] p78_res7__1022_comb;
  wire [127:0] p78_res__31_comb;
  wire [127:0] p78_permut__32_comb;
  wire [127:0] p78_xor_2058857_comb;
  wire [7:0] p78_bit_slice_2058858_comb;
  wire [7:0] p78_bit_slice_2058859_comb;
  wire [7:0] p78_bit_slice_2058860_comb;
  wire [7:0] p78_bit_slice_2058861_comb;
  wire [7:0] p78_bit_slice_2058862_comb;
  wire [7:0] p78_bit_slice_2058863_comb;
  wire [7:0] p78_bit_slice_2058864_comb;
  wire [7:0] p78_bit_slice_2058865_comb;
  wire [7:0] p78_bit_slice_2058866_comb;
  wire [7:0] p78_bit_slice_2058867_comb;
  wire [7:0] p78_bit_slice_2058868_comb;
  wire [7:0] p78_bit_slice_2058869_comb;
  wire [7:0] p78_bit_slice_2058870_comb;
  wire [7:0] p78_bit_slice_2058877_comb;
  wire [7:0] p78_bit_slice_2058879_comb;
  wire [7:0] p78_array_index_2058880_comb;
  wire [7:0] p78_array_index_2058881_comb;
  wire [7:0] p78_array_index_2058882_comb;
  wire [7:0] p78_array_index_2058883_comb;
  wire [7:0] p78_array_index_2058884_comb;
  wire [7:0] p78_array_index_2058885_comb;
  wire [7:0] p78_res7__1057_comb;
  wire [7:0] p78_array_index_2058888_comb;
  wire [7:0] p78_array_index_2058889_comb;
  wire [7:0] p78_array_index_2058890_comb;
  wire [7:0] p78_array_index_2058891_comb;
  wire [7:0] p78_array_index_2058892_comb;
  wire [7:0] p78_array_index_2058893_comb;
  wire [7:0] p78_array_index_2058894_comb;
  wire [7:0] p78_array_index_2058895_comb;
  wire [7:0] p78_array_index_2058896_comb;
  wire [7:0] p78_array_index_2058897_comb;
  wire [7:0] p78_array_index_2058898_comb;
  wire [7:0] p78_array_index_2058899_comb;
  wire [7:0] p78_array_index_2058900_comb;
  assign p78_array_index_2058764_comb = p77_literal_2043920[p77_res7__1002];
  assign p78_res7__1047_comb = p77_array_index_2058536 ^ p77_array_index_2058537 ^ p77_array_index_2058090 ^ p77_array_index_2058145 ^ p77_array_index_2058405 ^ p77_array_index_2058453 ^ p77_res7__1029 ^ p77_array_index_2058538 ^ p77_res7__1033 ^ p77_array_index_2058539 ^ p77_array_index_2058540 ^ p77_array_index_2058541 ^ p77_array_index_2058542 ^ p77_array_index_2058543 ^ p77_array_index_2058544 ^ p77_bit_slice_2058025;
  assign p78_res7__1014_comb = p77_literal_2043910[p77_res7__1012] ^ p77_literal_2043912[p77_res7__1010] ^ p77_literal_2043914[p77_res7__1008] ^ p77_literal_2043916[p77_res7__1006] ^ p77_literal_2043918[p77_res7__1004] ^ p78_array_index_2058764_comb ^ p77_res7__1000 ^ p77_literal_2043923[p77_res7__998] ^ p77_res7__996 ^ p77_array_index_2058464 ^ p77_array_index_2058414 ^ p77_array_index_2058152 ^ p77_array_index_2058095 ^ p77_literal_2043912[p77_array_index_2058032] ^ p77_literal_2043910[p77_array_index_2058033] ^ p77_array_index_2058034;
  assign p78_res7__1049_comb = p77_literal_2043910[p77_bit_slice_2058027] ^ p77_array_index_2058059 ^ p77_array_index_2058118 ^ p77_array_index_2058172 ^ p77_array_index_2058430 ^ p77_array_index_2058476 ^ p77_res7__1031 ^ p77_literal_2043923[p77_res7__1033] ^ p77_res7__1035 ^ p77_literal_2043920[p77_res7__1037] ^ p77_literal_2043918[p77_res7__1039] ^ p77_literal_2043916[p77_res7__1041] ^ p77_literal_2043914[p77_res7__1043] ^ p77_literal_2043912[p77_res7__1045] ^ p77_literal_2043910[p78_res7__1047_comb] ^ p77_bit_slice_2058026;
  assign p78_res7__1016_comb = p77_literal_2043910[p78_res7__1014_comb] ^ p77_literal_2043912[p77_res7__1012] ^ p77_literal_2043914[p77_res7__1010] ^ p77_literal_2043916[p77_res7__1008] ^ p77_literal_2043918[p77_res7__1006] ^ p77_literal_2043920[p77_res7__1004] ^ p77_res7__1002 ^ p77_literal_2043923[p77_res7__1000] ^ p77_res7__998 ^ p77_array_index_2058487 ^ p77_array_index_2058439 ^ p77_array_index_2058387 ^ p77_array_index_2058123 ^ p77_array_index_2058063 ^ p77_literal_2043910[p77_array_index_2058032] ^ p77_array_index_2058033;
  assign p78_res7__1051_comb = p77_literal_2043910[p77_bit_slice_2058028] ^ p77_array_index_2058091 ^ p77_array_index_2058146 ^ p77_array_index_2058406 ^ p77_array_index_2058454 ^ p77_array_index_2058498 ^ p77_res7__1033 ^ p77_literal_2043923[p77_res7__1035] ^ p77_res7__1037 ^ p77_literal_2043920[p77_res7__1039] ^ p77_literal_2043918[p77_res7__1041] ^ p77_literal_2043916[p77_res7__1043] ^ p77_literal_2043914[p77_res7__1045] ^ p77_literal_2043912[p78_res7__1047_comb] ^ p77_literal_2043910[p78_res7__1049_comb] ^ p77_bit_slice_2058027;
  assign p78_res7__1018_comb = p77_literal_2043910[p78_res7__1016_comb] ^ p77_literal_2043912[p78_res7__1014_comb] ^ p77_literal_2043914[p77_res7__1012] ^ p77_literal_2043916[p77_res7__1010] ^ p77_literal_2043918[p77_res7__1008] ^ p77_literal_2043920[p77_res7__1006] ^ p77_res7__1004 ^ p77_literal_2043923[p77_res7__1002] ^ p77_res7__1000 ^ p77_array_index_2058509 ^ p77_array_index_2058463 ^ p77_array_index_2058413 ^ p77_array_index_2058151 ^ p77_array_index_2058094 ^ p77_literal_2043910[p77_array_index_2058031] ^ p77_array_index_2058032;
  assign p78_res7__1053_comb = p77_array_index_2058060 ^ p77_array_index_2058119 ^ p77_array_index_2058173 ^ p77_array_index_2058431 ^ p77_array_index_2058477 ^ p77_array_index_2058519 ^ p77_res7__1035 ^ p77_literal_2043923[p77_res7__1037] ^ p77_res7__1039 ^ p77_literal_2043920[p77_res7__1041] ^ p77_literal_2043918[p77_res7__1043] ^ p77_literal_2043916[p77_res7__1045] ^ p77_literal_2043914[p78_res7__1047_comb] ^ p77_literal_2043912[p78_res7__1049_comb] ^ p77_literal_2043910[p78_res7__1051_comb] ^ p77_bit_slice_2058028;
  assign p78_res7__1020_comb = p77_literal_2043910[p78_res7__1018_comb] ^ p77_literal_2043912[p78_res7__1016_comb] ^ p77_literal_2043914[p78_res7__1014_comb] ^ p77_literal_2043916[p77_res7__1012] ^ p77_literal_2043918[p77_res7__1010] ^ p77_literal_2043920[p77_res7__1008] ^ p77_res7__1006 ^ p77_literal_2043923[p77_res7__1004] ^ p77_res7__1002 ^ p77_array_index_2058530 ^ p77_array_index_2058486 ^ p77_array_index_2058438 ^ p77_array_index_2058386 ^ p77_array_index_2058122 ^ p77_array_index_2058062 ^ p77_array_index_2058031;
  assign p78_res7__1055_comb = p77_array_index_2058092 ^ p77_array_index_2058147 ^ p77_array_index_2058407 ^ p77_array_index_2058455 ^ p77_array_index_2058499 ^ p77_array_index_2058539 ^ p77_res7__1037 ^ p77_literal_2043923[p77_res7__1039] ^ p77_res7__1041 ^ p77_literal_2043920[p77_res7__1043] ^ p77_literal_2043918[p77_res7__1045] ^ p77_literal_2043916[p78_res7__1047_comb] ^ p77_literal_2043914[p78_res7__1049_comb] ^ p77_literal_2043912[p78_res7__1051_comb] ^ p77_literal_2043910[p78_res7__1053_comb] ^ p77_bit_slice_2058029;
  assign p78_res7__1022_comb = p77_literal_2043910[p78_res7__1020_comb] ^ p77_literal_2043912[p78_res7__1018_comb] ^ p77_literal_2043914[p78_res7__1016_comb] ^ p77_literal_2043916[p78_res7__1014_comb] ^ p77_literal_2043918[p77_res7__1012] ^ p77_literal_2043920[p77_res7__1010] ^ p77_res7__1008 ^ p77_literal_2043923[p77_res7__1006] ^ p77_res7__1004 ^ p78_array_index_2058764_comb ^ p77_array_index_2058508 ^ p77_array_index_2058462 ^ p77_array_index_2058412 ^ p77_array_index_2058150 ^ p77_array_index_2058093 ^ p77_array_index_2058030;
  assign p78_res__31_comb = {p78_res7__1022_comb, p78_res7__1020_comb, p78_res7__1018_comb, p78_res7__1016_comb, p78_res7__1014_comb, p77_res7__1012, p77_res7__1010, p77_res7__1008, p77_res7__1006, p77_res7__1004, p77_res7__1002, p77_res7__1000, p77_res7__998, p77_res7__996, p77_res7__994, p77_res7__992};
  assign p78_permut__32_comb = {literal_2058836[p77_res7__1025], literal_2058836[p77_res7__1027], literal_2058836[p77_res7__1029], literal_2058836[p77_res7__1031], literal_2058836[p77_res7__1033], literal_2058836[p77_res7__1035], literal_2058836[p77_res7__1037], literal_2058836[p77_res7__1039], literal_2058836[p77_res7__1041], literal_2058836[p77_res7__1043], literal_2058836[p77_res7__1045], literal_2058836[p78_res7__1047_comb], literal_2058836[p78_res7__1049_comb], literal_2058836[p78_res7__1051_comb], literal_2058836[p78_res7__1053_comb], literal_2058836[p78_res7__1055_comb]};
  assign p78_xor_2058857_comb = p78_res__31_comb ^ p77_xor_2057490 ^ p78_permut__32_comb;
  assign p78_bit_slice_2058858_comb = p78_xor_2058857_comb[119:112];
  assign p78_bit_slice_2058859_comb = p78_xor_2058857_comb[111:104];
  assign p78_bit_slice_2058860_comb = p78_xor_2058857_comb[103:96];
  assign p78_bit_slice_2058861_comb = p78_xor_2058857_comb[95:88];
  assign p78_bit_slice_2058862_comb = p78_xor_2058857_comb[87:80];
  assign p78_bit_slice_2058863_comb = p78_xor_2058857_comb[79:72];
  assign p78_bit_slice_2058864_comb = p78_xor_2058857_comb[63:56];
  assign p78_bit_slice_2058865_comb = p78_xor_2058857_comb[47:40];
  assign p78_bit_slice_2058866_comb = p78_xor_2058857_comb[39:32];
  assign p78_bit_slice_2058867_comb = p78_xor_2058857_comb[31:24];
  assign p78_bit_slice_2058868_comb = p78_xor_2058857_comb[23:16];
  assign p78_bit_slice_2058869_comb = p78_xor_2058857_comb[15:8];
  assign p78_bit_slice_2058870_comb = p78_xor_2058857_comb[7:0];
  assign p78_bit_slice_2058877_comb = p78_xor_2058857_comb[71:64];
  assign p78_bit_slice_2058879_comb = p78_xor_2058857_comb[55:48];
  assign p78_array_index_2058880_comb = p77_literal_2043920[p78_bit_slice_2058865_comb];
  assign p78_array_index_2058881_comb = p77_literal_2043918[p78_bit_slice_2058866_comb];
  assign p78_array_index_2058882_comb = p77_literal_2043916[p78_bit_slice_2058867_comb];
  assign p78_array_index_2058883_comb = p77_literal_2043914[p78_bit_slice_2058868_comb];
  assign p78_array_index_2058884_comb = p77_literal_2043912[p78_bit_slice_2058869_comb];
  assign p78_array_index_2058885_comb = p77_literal_2043910[p78_bit_slice_2058870_comb];
  assign p78_res7__1057_comb = p77_literal_2043910[p78_bit_slice_2058858_comb] ^ p77_literal_2043912[p78_bit_slice_2058859_comb] ^ p77_literal_2043914[p78_bit_slice_2058860_comb] ^ p77_literal_2043916[p78_bit_slice_2058861_comb] ^ p77_literal_2043918[p78_bit_slice_2058862_comb] ^ p77_literal_2043920[p78_bit_slice_2058863_comb] ^ p78_bit_slice_2058877_comb ^ p77_literal_2043923[p78_bit_slice_2058864_comb] ^ p78_bit_slice_2058879_comb ^ p78_array_index_2058880_comb ^ p78_array_index_2058881_comb ^ p78_array_index_2058882_comb ^ p78_array_index_2058883_comb ^ p78_array_index_2058884_comb ^ p78_array_index_2058885_comb ^ p78_xor_2058857_comb[127:120];
  assign p78_array_index_2058888_comb = p77_literal_2043910[p78_bit_slice_2058859_comb];
  assign p78_array_index_2058889_comb = p77_literal_2043912[p78_bit_slice_2058860_comb];
  assign p78_array_index_2058890_comb = p77_literal_2043914[p78_bit_slice_2058861_comb];
  assign p78_array_index_2058891_comb = p77_literal_2043916[p78_bit_slice_2058862_comb];
  assign p78_array_index_2058892_comb = p77_literal_2043918[p78_bit_slice_2058863_comb];
  assign p78_array_index_2058893_comb = p77_literal_2043920[p78_bit_slice_2058877_comb];
  assign p78_array_index_2058894_comb = p77_literal_2043923[p78_bit_slice_2058879_comb];
  assign p78_array_index_2058895_comb = p77_literal_2043920[p78_bit_slice_2058866_comb];
  assign p78_array_index_2058896_comb = p77_literal_2043918[p78_bit_slice_2058867_comb];
  assign p78_array_index_2058897_comb = p77_literal_2043916[p78_bit_slice_2058868_comb];
  assign p78_array_index_2058898_comb = p77_literal_2043914[p78_bit_slice_2058869_comb];
  assign p78_array_index_2058899_comb = p77_literal_2043912[p78_bit_slice_2058870_comb];
  assign p78_array_index_2058900_comb = p77_literal_2043910[p78_res7__1057_comb];

  // Registers for pipe stage 78:
  reg [127:0] p78_bit_slice_2043893;
  reg [127:0] p78_bit_slice_2044018;
  reg [127:0] p78_k3;
  reg [127:0] p78_k2;
  reg [127:0] p78_k5;
  reg [127:0] p78_k4;
  reg [127:0] p78_k7;
  reg [127:0] p78_k6;
  reg [7:0] p78_bit_slice_2058858;
  reg [7:0] p78_bit_slice_2058859;
  reg [7:0] p78_bit_slice_2058860;
  reg [7:0] p78_bit_slice_2058861;
  reg [7:0] p78_bit_slice_2058862;
  reg [7:0] p78_bit_slice_2058863;
  reg [7:0] p78_bit_slice_2058864;
  reg [7:0] p78_bit_slice_2058865;
  reg [7:0] p78_bit_slice_2058866;
  reg [7:0] p78_bit_slice_2058867;
  reg [7:0] p78_bit_slice_2058868;
  reg [7:0] p78_bit_slice_2058869;
  reg [7:0] p78_bit_slice_2058870;
  reg [7:0] p78_bit_slice_2058877;
  reg [7:0] p78_bit_slice_2058879;
  reg [7:0] p78_array_index_2058880;
  reg [7:0] p78_array_index_2058881;
  reg [7:0] p78_array_index_2058882;
  reg [7:0] p78_array_index_2058883;
  reg [7:0] p78_array_index_2058884;
  reg [7:0] p78_array_index_2058885;
  reg [7:0] p78_res7__1057;
  reg [7:0] p78_array_index_2058888;
  reg [7:0] p78_array_index_2058889;
  reg [7:0] p78_array_index_2058890;
  reg [7:0] p78_array_index_2058891;
  reg [7:0] p78_array_index_2058892;
  reg [7:0] p78_array_index_2058893;
  reg [7:0] p78_array_index_2058894;
  reg [7:0] p78_array_index_2058895;
  reg [7:0] p78_array_index_2058896;
  reg [7:0] p78_array_index_2058897;
  reg [7:0] p78_array_index_2058898;
  reg [7:0] p78_array_index_2058899;
  reg [7:0] p78_array_index_2058900;
  reg [7:0] p79_literal_2043910[256];
  reg [7:0] p79_literal_2043912[256];
  reg [7:0] p79_literal_2043914[256];
  reg [7:0] p79_literal_2043916[256];
  reg [7:0] p79_literal_2043918[256];
  reg [7:0] p79_literal_2043920[256];
  reg [7:0] p79_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p78_bit_slice_2043893 <= p77_bit_slice_2043893;
    p78_bit_slice_2044018 <= p77_bit_slice_2044018;
    p78_k3 <= p77_k3;
    p78_k2 <= p77_k2;
    p78_k5 <= p77_k5;
    p78_k4 <= p77_k4;
    p78_k7 <= p77_k7;
    p78_k6 <= p77_k6;
    p78_bit_slice_2058858 <= p78_bit_slice_2058858_comb;
    p78_bit_slice_2058859 <= p78_bit_slice_2058859_comb;
    p78_bit_slice_2058860 <= p78_bit_slice_2058860_comb;
    p78_bit_slice_2058861 <= p78_bit_slice_2058861_comb;
    p78_bit_slice_2058862 <= p78_bit_slice_2058862_comb;
    p78_bit_slice_2058863 <= p78_bit_slice_2058863_comb;
    p78_bit_slice_2058864 <= p78_bit_slice_2058864_comb;
    p78_bit_slice_2058865 <= p78_bit_slice_2058865_comb;
    p78_bit_slice_2058866 <= p78_bit_slice_2058866_comb;
    p78_bit_slice_2058867 <= p78_bit_slice_2058867_comb;
    p78_bit_slice_2058868 <= p78_bit_slice_2058868_comb;
    p78_bit_slice_2058869 <= p78_bit_slice_2058869_comb;
    p78_bit_slice_2058870 <= p78_bit_slice_2058870_comb;
    p78_bit_slice_2058877 <= p78_bit_slice_2058877_comb;
    p78_bit_slice_2058879 <= p78_bit_slice_2058879_comb;
    p78_array_index_2058880 <= p78_array_index_2058880_comb;
    p78_array_index_2058881 <= p78_array_index_2058881_comb;
    p78_array_index_2058882 <= p78_array_index_2058882_comb;
    p78_array_index_2058883 <= p78_array_index_2058883_comb;
    p78_array_index_2058884 <= p78_array_index_2058884_comb;
    p78_array_index_2058885 <= p78_array_index_2058885_comb;
    p78_res7__1057 <= p78_res7__1057_comb;
    p78_array_index_2058888 <= p78_array_index_2058888_comb;
    p78_array_index_2058889 <= p78_array_index_2058889_comb;
    p78_array_index_2058890 <= p78_array_index_2058890_comb;
    p78_array_index_2058891 <= p78_array_index_2058891_comb;
    p78_array_index_2058892 <= p78_array_index_2058892_comb;
    p78_array_index_2058893 <= p78_array_index_2058893_comb;
    p78_array_index_2058894 <= p78_array_index_2058894_comb;
    p78_array_index_2058895 <= p78_array_index_2058895_comb;
    p78_array_index_2058896 <= p78_array_index_2058896_comb;
    p78_array_index_2058897 <= p78_array_index_2058897_comb;
    p78_array_index_2058898 <= p78_array_index_2058898_comb;
    p78_array_index_2058899 <= p78_array_index_2058899_comb;
    p78_array_index_2058900 <= p78_array_index_2058900_comb;
    p79_literal_2043910 <= p78_literal_2043910;
    p79_literal_2043912 <= p78_literal_2043912;
    p79_literal_2043914 <= p78_literal_2043914;
    p79_literal_2043916 <= p78_literal_2043916;
    p79_literal_2043918 <= p78_literal_2043918;
    p79_literal_2043920 <= p78_literal_2043920;
    p79_literal_2043923 <= p78_literal_2043923;
  end

  // ===== Pipe stage 79:
  wire [7:0] p79_res7__1059_comb;
  wire [7:0] p79_array_index_2059011_comb;
  wire [7:0] p79_array_index_2059012_comb;
  wire [7:0] p79_array_index_2059013_comb;
  wire [7:0] p79_array_index_2059014_comb;
  wire [7:0] p79_array_index_2059015_comb;
  wire [7:0] p79_res7__1061_comb;
  wire [7:0] p79_array_index_2059025_comb;
  wire [7:0] p79_array_index_2059026_comb;
  wire [7:0] p79_array_index_2059027_comb;
  wire [7:0] p79_array_index_2059028_comb;
  wire [7:0] p79_array_index_2059029_comb;
  wire [7:0] p79_res7__1063_comb;
  wire [7:0] p79_array_index_2059038_comb;
  wire [7:0] p79_array_index_2059039_comb;
  wire [7:0] p79_array_index_2059040_comb;
  wire [7:0] p79_array_index_2059041_comb;
  wire [7:0] p79_res7__1065_comb;
  wire [7:0] p79_array_index_2059051_comb;
  wire [7:0] p79_array_index_2059052_comb;
  wire [7:0] p79_array_index_2059053_comb;
  wire [7:0] p79_array_index_2059054_comb;
  wire [7:0] p79_res7__1067_comb;
  wire [7:0] p79_array_index_2059063_comb;
  wire [7:0] p79_array_index_2059064_comb;
  wire [7:0] p79_array_index_2059065_comb;
  wire [7:0] p79_res7__1069_comb;
  wire [7:0] p79_array_index_2059075_comb;
  wire [7:0] p79_array_index_2059076_comb;
  wire [7:0] p79_array_index_2059077_comb;
  wire [7:0] p79_res7__1071_comb;
  wire [7:0] p79_array_index_2059082_comb;
  wire [7:0] p79_array_index_2059083_comb;
  wire [7:0] p79_array_index_2059084_comb;
  wire [7:0] p79_array_index_2059085_comb;
  wire [7:0] p79_array_index_2059086_comb;
  wire [7:0] p79_array_index_2059087_comb;
  wire [7:0] p79_array_index_2059088_comb;
  wire [7:0] p79_array_index_2059089_comb;
  wire [7:0] p79_array_index_2059090_comb;
  wire [7:0] p79_array_index_2059091_comb;
  assign p79_res7__1059_comb = p78_array_index_2058888 ^ p78_array_index_2058889 ^ p78_array_index_2058890 ^ p78_array_index_2058891 ^ p78_array_index_2058892 ^ p78_array_index_2058893 ^ p78_bit_slice_2058864 ^ p78_array_index_2058894 ^ p78_bit_slice_2058865 ^ p78_array_index_2058895 ^ p78_array_index_2058896 ^ p78_array_index_2058897 ^ p78_array_index_2058898 ^ p78_array_index_2058899 ^ p78_array_index_2058900 ^ p78_bit_slice_2058858;
  assign p79_array_index_2059011_comb = p78_literal_2043920[p78_bit_slice_2058867];
  assign p79_array_index_2059012_comb = p78_literal_2043918[p78_bit_slice_2058868];
  assign p79_array_index_2059013_comb = p78_literal_2043916[p78_bit_slice_2058869];
  assign p79_array_index_2059014_comb = p78_literal_2043914[p78_bit_slice_2058870];
  assign p79_array_index_2059015_comb = p78_literal_2043912[p78_res7__1057];
  assign p79_res7__1061_comb = p78_literal_2043910[p78_bit_slice_2058860] ^ p78_literal_2043912[p78_bit_slice_2058861] ^ p78_literal_2043914[p78_bit_slice_2058862] ^ p78_literal_2043916[p78_bit_slice_2058863] ^ p78_literal_2043918[p78_bit_slice_2058877] ^ p78_literal_2043920[p78_bit_slice_2058864] ^ p78_bit_slice_2058879 ^ p78_literal_2043923[p78_bit_slice_2058865] ^ p78_bit_slice_2058866 ^ p79_array_index_2059011_comb ^ p79_array_index_2059012_comb ^ p79_array_index_2059013_comb ^ p79_array_index_2059014_comb ^ p79_array_index_2059015_comb ^ p78_literal_2043910[p79_res7__1059_comb] ^ p78_bit_slice_2058859;
  assign p79_array_index_2059025_comb = p78_literal_2043920[p78_bit_slice_2058868];
  assign p79_array_index_2059026_comb = p78_literal_2043918[p78_bit_slice_2058869];
  assign p79_array_index_2059027_comb = p78_literal_2043916[p78_bit_slice_2058870];
  assign p79_array_index_2059028_comb = p78_literal_2043914[p78_res7__1057];
  assign p79_array_index_2059029_comb = p78_literal_2043912[p79_res7__1059_comb];
  assign p79_res7__1063_comb = p78_literal_2043910[p78_bit_slice_2058861] ^ p78_literal_2043912[p78_bit_slice_2058862] ^ p78_literal_2043914[p78_bit_slice_2058863] ^ p78_literal_2043916[p78_bit_slice_2058877] ^ p78_literal_2043918[p78_bit_slice_2058864] ^ p78_literal_2043920[p78_bit_slice_2058879] ^ p78_bit_slice_2058865 ^ p78_literal_2043923[p78_bit_slice_2058866] ^ p78_bit_slice_2058867 ^ p79_array_index_2059025_comb ^ p79_array_index_2059026_comb ^ p79_array_index_2059027_comb ^ p79_array_index_2059028_comb ^ p79_array_index_2059029_comb ^ p78_literal_2043910[p79_res7__1061_comb] ^ p78_bit_slice_2058860;
  assign p79_array_index_2059038_comb = p78_literal_2043920[p78_bit_slice_2058869];
  assign p79_array_index_2059039_comb = p78_literal_2043918[p78_bit_slice_2058870];
  assign p79_array_index_2059040_comb = p78_literal_2043916[p78_res7__1057];
  assign p79_array_index_2059041_comb = p78_literal_2043914[p79_res7__1059_comb];
  assign p79_res7__1065_comb = p78_literal_2043910[p78_bit_slice_2058862] ^ p78_literal_2043912[p78_bit_slice_2058863] ^ p78_literal_2043914[p78_bit_slice_2058877] ^ p78_literal_2043916[p78_bit_slice_2058864] ^ p78_literal_2043918[p78_bit_slice_2058879] ^ p78_array_index_2058880 ^ p78_bit_slice_2058866 ^ p78_literal_2043923[p78_bit_slice_2058867] ^ p78_bit_slice_2058868 ^ p79_array_index_2059038_comb ^ p79_array_index_2059039_comb ^ p79_array_index_2059040_comb ^ p79_array_index_2059041_comb ^ p78_literal_2043912[p79_res7__1061_comb] ^ p78_literal_2043910[p79_res7__1063_comb] ^ p78_bit_slice_2058861;
  assign p79_array_index_2059051_comb = p78_literal_2043920[p78_bit_slice_2058870];
  assign p79_array_index_2059052_comb = p78_literal_2043918[p78_res7__1057];
  assign p79_array_index_2059053_comb = p78_literal_2043916[p79_res7__1059_comb];
  assign p79_array_index_2059054_comb = p78_literal_2043914[p79_res7__1061_comb];
  assign p79_res7__1067_comb = p78_literal_2043910[p78_bit_slice_2058863] ^ p78_literal_2043912[p78_bit_slice_2058877] ^ p78_literal_2043914[p78_bit_slice_2058864] ^ p78_literal_2043916[p78_bit_slice_2058879] ^ p78_literal_2043918[p78_bit_slice_2058865] ^ p78_array_index_2058895 ^ p78_bit_slice_2058867 ^ p78_literal_2043923[p78_bit_slice_2058868] ^ p78_bit_slice_2058869 ^ p79_array_index_2059051_comb ^ p79_array_index_2059052_comb ^ p79_array_index_2059053_comb ^ p79_array_index_2059054_comb ^ p78_literal_2043912[p79_res7__1063_comb] ^ p78_literal_2043910[p79_res7__1065_comb] ^ p78_bit_slice_2058862;
  assign p79_array_index_2059063_comb = p78_literal_2043920[p78_res7__1057];
  assign p79_array_index_2059064_comb = p78_literal_2043918[p79_res7__1059_comb];
  assign p79_array_index_2059065_comb = p78_literal_2043916[p79_res7__1061_comb];
  assign p79_res7__1069_comb = p78_literal_2043910[p78_bit_slice_2058877] ^ p78_literal_2043912[p78_bit_slice_2058864] ^ p78_literal_2043914[p78_bit_slice_2058879] ^ p78_literal_2043916[p78_bit_slice_2058865] ^ p78_array_index_2058881 ^ p79_array_index_2059011_comb ^ p78_bit_slice_2058868 ^ p78_literal_2043923[p78_bit_slice_2058869] ^ p78_bit_slice_2058870 ^ p79_array_index_2059063_comb ^ p79_array_index_2059064_comb ^ p79_array_index_2059065_comb ^ p78_literal_2043914[p79_res7__1063_comb] ^ p78_literal_2043912[p79_res7__1065_comb] ^ p78_literal_2043910[p79_res7__1067_comb] ^ p78_bit_slice_2058863;
  assign p79_array_index_2059075_comb = p78_literal_2043920[p79_res7__1059_comb];
  assign p79_array_index_2059076_comb = p78_literal_2043918[p79_res7__1061_comb];
  assign p79_array_index_2059077_comb = p78_literal_2043916[p79_res7__1063_comb];
  assign p79_res7__1071_comb = p78_literal_2043910[p78_bit_slice_2058864] ^ p78_literal_2043912[p78_bit_slice_2058879] ^ p78_literal_2043914[p78_bit_slice_2058865] ^ p78_literal_2043916[p78_bit_slice_2058866] ^ p78_array_index_2058896 ^ p79_array_index_2059025_comb ^ p78_bit_slice_2058869 ^ p78_literal_2043923[p78_bit_slice_2058870] ^ p78_res7__1057 ^ p79_array_index_2059075_comb ^ p79_array_index_2059076_comb ^ p79_array_index_2059077_comb ^ p78_literal_2043914[p79_res7__1065_comb] ^ p78_literal_2043912[p79_res7__1067_comb] ^ p78_literal_2043910[p79_res7__1069_comb] ^ p78_bit_slice_2058877;
  assign p79_array_index_2059082_comb = p78_literal_2043910[p78_bit_slice_2058879];
  assign p79_array_index_2059083_comb = p78_literal_2043912[p78_bit_slice_2058865];
  assign p79_array_index_2059084_comb = p78_literal_2043914[p78_bit_slice_2058866];
  assign p79_array_index_2059085_comb = p78_literal_2043923[p78_res7__1057];
  assign p79_array_index_2059086_comb = p78_literal_2043920[p79_res7__1061_comb];
  assign p79_array_index_2059087_comb = p78_literal_2043918[p79_res7__1063_comb];
  assign p79_array_index_2059088_comb = p78_literal_2043916[p79_res7__1065_comb];
  assign p79_array_index_2059089_comb = p78_literal_2043914[p79_res7__1067_comb];
  assign p79_array_index_2059090_comb = p78_literal_2043912[p79_res7__1069_comb];
  assign p79_array_index_2059091_comb = p78_literal_2043910[p79_res7__1071_comb];

  // Registers for pipe stage 79:
  reg [127:0] p79_bit_slice_2043893;
  reg [127:0] p79_bit_slice_2044018;
  reg [127:0] p79_k3;
  reg [127:0] p79_k2;
  reg [127:0] p79_k5;
  reg [127:0] p79_k4;
  reg [127:0] p79_k7;
  reg [127:0] p79_k6;
  reg [7:0] p79_bit_slice_2058864;
  reg [7:0] p79_bit_slice_2058865;
  reg [7:0] p79_bit_slice_2058866;
  reg [7:0] p79_bit_slice_2058867;
  reg [7:0] p79_bit_slice_2058868;
  reg [7:0] p79_bit_slice_2058869;
  reg [7:0] p79_bit_slice_2058870;
  reg [7:0] p79_bit_slice_2058879;
  reg [7:0] p79_array_index_2058882;
  reg [7:0] p79_array_index_2058883;
  reg [7:0] p79_array_index_2058884;
  reg [7:0] p79_array_index_2058885;
  reg [7:0] p79_res7__1057;
  reg [7:0] p79_array_index_2058897;
  reg [7:0] p79_array_index_2058898;
  reg [7:0] p79_array_index_2058899;
  reg [7:0] p79_array_index_2058900;
  reg [7:0] p79_res7__1059;
  reg [7:0] p79_array_index_2059012;
  reg [7:0] p79_array_index_2059013;
  reg [7:0] p79_array_index_2059014;
  reg [7:0] p79_array_index_2059015;
  reg [7:0] p79_res7__1061;
  reg [7:0] p79_array_index_2059026;
  reg [7:0] p79_array_index_2059027;
  reg [7:0] p79_array_index_2059028;
  reg [7:0] p79_array_index_2059029;
  reg [7:0] p79_res7__1063;
  reg [7:0] p79_array_index_2059038;
  reg [7:0] p79_array_index_2059039;
  reg [7:0] p79_array_index_2059040;
  reg [7:0] p79_array_index_2059041;
  reg [7:0] p79_res7__1065;
  reg [7:0] p79_array_index_2059051;
  reg [7:0] p79_array_index_2059052;
  reg [7:0] p79_array_index_2059053;
  reg [7:0] p79_array_index_2059054;
  reg [7:0] p79_res7__1067;
  reg [7:0] p79_array_index_2059063;
  reg [7:0] p79_array_index_2059064;
  reg [7:0] p79_array_index_2059065;
  reg [7:0] p79_res7__1069;
  reg [7:0] p79_array_index_2059075;
  reg [7:0] p79_array_index_2059076;
  reg [7:0] p79_array_index_2059077;
  reg [7:0] p79_res7__1071;
  reg [7:0] p79_array_index_2059082;
  reg [7:0] p79_array_index_2059083;
  reg [7:0] p79_array_index_2059084;
  reg [7:0] p79_array_index_2059085;
  reg [7:0] p79_array_index_2059086;
  reg [7:0] p79_array_index_2059087;
  reg [7:0] p79_array_index_2059088;
  reg [7:0] p79_array_index_2059089;
  reg [7:0] p79_array_index_2059090;
  reg [7:0] p79_array_index_2059091;
  reg [7:0] p80_literal_2043910[256];
  reg [7:0] p80_literal_2043912[256];
  reg [7:0] p80_literal_2043914[256];
  reg [7:0] p80_literal_2043916[256];
  reg [7:0] p80_literal_2043918[256];
  reg [7:0] p80_literal_2043920[256];
  reg [7:0] p80_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p79_bit_slice_2043893 <= p78_bit_slice_2043893;
    p79_bit_slice_2044018 <= p78_bit_slice_2044018;
    p79_k3 <= p78_k3;
    p79_k2 <= p78_k2;
    p79_k5 <= p78_k5;
    p79_k4 <= p78_k4;
    p79_k7 <= p78_k7;
    p79_k6 <= p78_k6;
    p79_bit_slice_2058864 <= p78_bit_slice_2058864;
    p79_bit_slice_2058865 <= p78_bit_slice_2058865;
    p79_bit_slice_2058866 <= p78_bit_slice_2058866;
    p79_bit_slice_2058867 <= p78_bit_slice_2058867;
    p79_bit_slice_2058868 <= p78_bit_slice_2058868;
    p79_bit_slice_2058869 <= p78_bit_slice_2058869;
    p79_bit_slice_2058870 <= p78_bit_slice_2058870;
    p79_bit_slice_2058879 <= p78_bit_slice_2058879;
    p79_array_index_2058882 <= p78_array_index_2058882;
    p79_array_index_2058883 <= p78_array_index_2058883;
    p79_array_index_2058884 <= p78_array_index_2058884;
    p79_array_index_2058885 <= p78_array_index_2058885;
    p79_res7__1057 <= p78_res7__1057;
    p79_array_index_2058897 <= p78_array_index_2058897;
    p79_array_index_2058898 <= p78_array_index_2058898;
    p79_array_index_2058899 <= p78_array_index_2058899;
    p79_array_index_2058900 <= p78_array_index_2058900;
    p79_res7__1059 <= p79_res7__1059_comb;
    p79_array_index_2059012 <= p79_array_index_2059012_comb;
    p79_array_index_2059013 <= p79_array_index_2059013_comb;
    p79_array_index_2059014 <= p79_array_index_2059014_comb;
    p79_array_index_2059015 <= p79_array_index_2059015_comb;
    p79_res7__1061 <= p79_res7__1061_comb;
    p79_array_index_2059026 <= p79_array_index_2059026_comb;
    p79_array_index_2059027 <= p79_array_index_2059027_comb;
    p79_array_index_2059028 <= p79_array_index_2059028_comb;
    p79_array_index_2059029 <= p79_array_index_2059029_comb;
    p79_res7__1063 <= p79_res7__1063_comb;
    p79_array_index_2059038 <= p79_array_index_2059038_comb;
    p79_array_index_2059039 <= p79_array_index_2059039_comb;
    p79_array_index_2059040 <= p79_array_index_2059040_comb;
    p79_array_index_2059041 <= p79_array_index_2059041_comb;
    p79_res7__1065 <= p79_res7__1065_comb;
    p79_array_index_2059051 <= p79_array_index_2059051_comb;
    p79_array_index_2059052 <= p79_array_index_2059052_comb;
    p79_array_index_2059053 <= p79_array_index_2059053_comb;
    p79_array_index_2059054 <= p79_array_index_2059054_comb;
    p79_res7__1067 <= p79_res7__1067_comb;
    p79_array_index_2059063 <= p79_array_index_2059063_comb;
    p79_array_index_2059064 <= p79_array_index_2059064_comb;
    p79_array_index_2059065 <= p79_array_index_2059065_comb;
    p79_res7__1069 <= p79_res7__1069_comb;
    p79_array_index_2059075 <= p79_array_index_2059075_comb;
    p79_array_index_2059076 <= p79_array_index_2059076_comb;
    p79_array_index_2059077 <= p79_array_index_2059077_comb;
    p79_res7__1071 <= p79_res7__1071_comb;
    p79_array_index_2059082 <= p79_array_index_2059082_comb;
    p79_array_index_2059083 <= p79_array_index_2059083_comb;
    p79_array_index_2059084 <= p79_array_index_2059084_comb;
    p79_array_index_2059085 <= p79_array_index_2059085_comb;
    p79_array_index_2059086 <= p79_array_index_2059086_comb;
    p79_array_index_2059087 <= p79_array_index_2059087_comb;
    p79_array_index_2059088 <= p79_array_index_2059088_comb;
    p79_array_index_2059089 <= p79_array_index_2059089_comb;
    p79_array_index_2059090 <= p79_array_index_2059090_comb;
    p79_array_index_2059091 <= p79_array_index_2059091_comb;
    p80_literal_2043910 <= p79_literal_2043910;
    p80_literal_2043912 <= p79_literal_2043912;
    p80_literal_2043914 <= p79_literal_2043914;
    p80_literal_2043916 <= p79_literal_2043916;
    p80_literal_2043918 <= p79_literal_2043918;
    p80_literal_2043920 <= p79_literal_2043920;
    p80_literal_2043923 <= p79_literal_2043923;
  end

  // ===== Pipe stage 80:
  wire [7:0] p80_res7__1073_comb;
  wire [7:0] p80_array_index_2059241_comb;
  wire [7:0] p80_array_index_2059242_comb;
  wire [7:0] p80_res7__1075_comb;
  wire [7:0] p80_array_index_2059251_comb;
  wire [7:0] p80_res7__1077_comb;
  wire [7:0] p80_array_index_2059261_comb;
  wire [7:0] p80_res7__1079_comb;
  wire [7:0] p80_res7__1081_comb;
  wire [7:0] p80_res7__1083_comb;
  wire [7:0] p80_res7__1085_comb;
  wire [7:0] p80_array_index_2059294_comb;
  wire [7:0] p80_array_index_2059295_comb;
  wire [7:0] p80_array_index_2059296_comb;
  wire [7:0] p80_array_index_2059297_comb;
  wire [7:0] p80_array_index_2059298_comb;
  wire [7:0] p80_array_index_2059299_comb;
  wire [7:0] p80_array_index_2059300_comb;
  wire [7:0] p80_array_index_2059301_comb;
  wire [7:0] p80_array_index_2059302_comb;
  wire [7:0] p80_array_index_2059303_comb;
  wire [7:0] p80_array_index_2059304_comb;
  wire [7:0] p80_array_index_2059305_comb;
  wire [7:0] p80_array_index_2059306_comb;
  wire [7:0] p80_array_index_2059307_comb;
  wire [7:0] p80_array_index_2059308_comb;
  wire [7:0] p80_array_index_2059309_comb;
  wire [7:0] p80_array_index_2059310_comb;
  wire [7:0] p80_array_index_2059311_comb;
  wire [7:0] p80_array_index_2059312_comb;
  wire [7:0] p80_array_index_2059313_comb;
  assign p80_res7__1073_comb = p79_array_index_2059082 ^ p79_array_index_2059083 ^ p79_array_index_2059084 ^ p79_array_index_2058882 ^ p79_array_index_2059012 ^ p79_array_index_2059038 ^ p79_bit_slice_2058870 ^ p79_array_index_2059085 ^ p79_res7__1059 ^ p79_array_index_2059086 ^ p79_array_index_2059087 ^ p79_array_index_2059088 ^ p79_array_index_2059089 ^ p79_array_index_2059090 ^ p79_array_index_2059091 ^ p79_bit_slice_2058864;
  assign p80_array_index_2059241_comb = p79_literal_2043920[p79_res7__1063];
  assign p80_array_index_2059242_comb = p79_literal_2043918[p79_res7__1065];
  assign p80_res7__1075_comb = p79_literal_2043910[p79_bit_slice_2058865] ^ p79_literal_2043912[p79_bit_slice_2058866] ^ p79_literal_2043914[p79_bit_slice_2058867] ^ p79_array_index_2058897 ^ p79_array_index_2059026 ^ p79_array_index_2059051 ^ p79_res7__1057 ^ p79_literal_2043923[p79_res7__1059] ^ p79_res7__1061 ^ p80_array_index_2059241_comb ^ p80_array_index_2059242_comb ^ p79_literal_2043916[p79_res7__1067] ^ p79_literal_2043914[p79_res7__1069] ^ p79_literal_2043912[p79_res7__1071] ^ p79_literal_2043910[p80_res7__1073_comb] ^ p79_bit_slice_2058879;
  assign p80_array_index_2059251_comb = p79_literal_2043920[p79_res7__1065];
  assign p80_res7__1077_comb = p79_literal_2043910[p79_bit_slice_2058866] ^ p79_literal_2043912[p79_bit_slice_2058867] ^ p79_array_index_2058883 ^ p79_array_index_2059013 ^ p79_array_index_2059039 ^ p79_array_index_2059063 ^ p79_res7__1059 ^ p79_literal_2043923[p79_res7__1061] ^ p79_res7__1063 ^ p80_array_index_2059251_comb ^ p79_literal_2043918[p79_res7__1067] ^ p79_literal_2043916[p79_res7__1069] ^ p79_literal_2043914[p79_res7__1071] ^ p79_literal_2043912[p80_res7__1073_comb] ^ p79_literal_2043910[p80_res7__1075_comb] ^ p79_bit_slice_2058865;
  assign p80_array_index_2059261_comb = p79_literal_2043920[p79_res7__1067];
  assign p80_res7__1079_comb = p79_literal_2043910[p79_bit_slice_2058867] ^ p79_literal_2043912[p79_bit_slice_2058868] ^ p79_array_index_2058898 ^ p79_array_index_2059027 ^ p79_array_index_2059052 ^ p79_array_index_2059075 ^ p79_res7__1061 ^ p79_literal_2043923[p79_res7__1063] ^ p79_res7__1065 ^ p80_array_index_2059261_comb ^ p79_literal_2043918[p79_res7__1069] ^ p79_literal_2043916[p79_res7__1071] ^ p79_literal_2043914[p80_res7__1073_comb] ^ p79_literal_2043912[p80_res7__1075_comb] ^ p79_literal_2043910[p80_res7__1077_comb] ^ p79_bit_slice_2058866;
  assign p80_res7__1081_comb = p79_literal_2043910[p79_bit_slice_2058868] ^ p79_array_index_2058884 ^ p79_array_index_2059014 ^ p79_array_index_2059040 ^ p79_array_index_2059064 ^ p79_array_index_2059086 ^ p79_res7__1063 ^ p79_literal_2043923[p79_res7__1065] ^ p79_res7__1067 ^ p79_literal_2043920[p79_res7__1069] ^ p79_literal_2043918[p79_res7__1071] ^ p79_literal_2043916[p80_res7__1073_comb] ^ p79_literal_2043914[p80_res7__1075_comb] ^ p79_literal_2043912[p80_res7__1077_comb] ^ p79_literal_2043910[p80_res7__1079_comb] ^ p79_bit_slice_2058867;
  assign p80_res7__1083_comb = p79_literal_2043910[p79_bit_slice_2058869] ^ p79_array_index_2058899 ^ p79_array_index_2059028 ^ p79_array_index_2059053 ^ p79_array_index_2059076 ^ p80_array_index_2059241_comb ^ p79_res7__1065 ^ p79_literal_2043923[p79_res7__1067] ^ p79_res7__1069 ^ p79_literal_2043920[p79_res7__1071] ^ p79_literal_2043918[p80_res7__1073_comb] ^ p79_literal_2043916[p80_res7__1075_comb] ^ p79_literal_2043914[p80_res7__1077_comb] ^ p79_literal_2043912[p80_res7__1079_comb] ^ p79_literal_2043910[p80_res7__1081_comb] ^ p79_bit_slice_2058868;
  assign p80_res7__1085_comb = p79_array_index_2058885 ^ p79_array_index_2059015 ^ p79_array_index_2059041 ^ p79_array_index_2059065 ^ p79_array_index_2059087 ^ p80_array_index_2059251_comb ^ p79_res7__1067 ^ p79_literal_2043923[p79_res7__1069] ^ p79_res7__1071 ^ p79_literal_2043920[p80_res7__1073_comb] ^ p79_literal_2043918[p80_res7__1075_comb] ^ p79_literal_2043916[p80_res7__1077_comb] ^ p79_literal_2043914[p80_res7__1079_comb] ^ p79_literal_2043912[p80_res7__1081_comb] ^ p79_literal_2043910[p80_res7__1083_comb] ^ p79_bit_slice_2058869;
  assign p80_array_index_2059294_comb = p79_literal_2043923[p79_res7__1071];
  assign p80_array_index_2059295_comb = p79_literal_2043920[p80_res7__1075_comb];
  assign p80_array_index_2059296_comb = p79_literal_2043918[p80_res7__1077_comb];
  assign p80_array_index_2059297_comb = p79_literal_2043916[p80_res7__1079_comb];
  assign p80_array_index_2059298_comb = p79_literal_2043914[p80_res7__1081_comb];
  assign p80_array_index_2059299_comb = p79_literal_2043912[p80_res7__1083_comb];
  assign p80_array_index_2059300_comb = p79_literal_2043910[p80_res7__1085_comb];
  assign p80_array_index_2059301_comb = p79_literal_2058836[p79_res7__1057];
  assign p80_array_index_2059302_comb = p79_literal_2058836[p79_res7__1059];
  assign p80_array_index_2059303_comb = p79_literal_2058836[p79_res7__1061];
  assign p80_array_index_2059304_comb = p79_literal_2058836[p79_res7__1063];
  assign p80_array_index_2059305_comb = p79_literal_2058836[p79_res7__1065];
  assign p80_array_index_2059306_comb = p79_literal_2058836[p79_res7__1067];
  assign p80_array_index_2059307_comb = p79_literal_2058836[p79_res7__1071];
  assign p80_array_index_2059308_comb = p79_literal_2058836[p80_res7__1075_comb];
  assign p80_array_index_2059309_comb = p79_literal_2058836[p80_res7__1077_comb];
  assign p80_array_index_2059310_comb = p79_literal_2058836[p80_res7__1079_comb];
  assign p80_array_index_2059311_comb = p79_literal_2058836[p80_res7__1081_comb];
  assign p80_array_index_2059312_comb = p79_literal_2058836[p80_res7__1083_comb];
  assign p80_array_index_2059313_comb = p79_literal_2058836[p80_res7__1085_comb];

  // Registers for pipe stage 80:
  reg [127:0] p80_bit_slice_2043893;
  reg [127:0] p80_bit_slice_2044018;
  reg [127:0] p80_k3;
  reg [127:0] p80_k2;
  reg [127:0] p80_k5;
  reg [127:0] p80_k4;
  reg [127:0] p80_k7;
  reg [127:0] p80_k6;
  reg [7:0] p80_bit_slice_2058870;
  reg [7:0] p80_array_index_2058900;
  reg [7:0] p80_array_index_2059029;
  reg [7:0] p80_array_index_2059054;
  reg [7:0] p80_res7__1069;
  reg [7:0] p80_array_index_2059077;
  reg [7:0] p80_res7__1073;
  reg [7:0] p80_array_index_2059242;
  reg [7:0] p80_array_index_2059261;
  reg [7:0] p80_array_index_2059294;
  reg [7:0] p80_array_index_2059295;
  reg [7:0] p80_array_index_2059296;
  reg [7:0] p80_array_index_2059297;
  reg [7:0] p80_array_index_2059298;
  reg [7:0] p80_array_index_2059299;
  reg [7:0] p80_array_index_2059300;
  reg [7:0] p80_array_index_2059301;
  reg [7:0] p80_array_index_2059302;
  reg [7:0] p80_array_index_2059303;
  reg [7:0] p80_array_index_2059304;
  reg [7:0] p80_array_index_2059305;
  reg [7:0] p80_array_index_2059306;
  reg [7:0] p80_array_index_2059307;
  reg [7:0] p80_array_index_2059308;
  reg [7:0] p80_array_index_2059309;
  reg [7:0] p80_array_index_2059310;
  reg [7:0] p80_array_index_2059311;
  reg [7:0] p80_array_index_2059312;
  reg [7:0] p80_array_index_2059313;
  reg [7:0] p81_literal_2043910[256];
  reg [7:0] p81_literal_2043912[256];
  reg [7:0] p81_literal_2043914[256];
  reg [7:0] p81_literal_2043916[256];
  reg [7:0] p81_literal_2043918[256];
  reg [7:0] p81_literal_2043920[256];
  reg [7:0] p81_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p80_bit_slice_2043893 <= p79_bit_slice_2043893;
    p80_bit_slice_2044018 <= p79_bit_slice_2044018;
    p80_k3 <= p79_k3;
    p80_k2 <= p79_k2;
    p80_k5 <= p79_k5;
    p80_k4 <= p79_k4;
    p80_k7 <= p79_k7;
    p80_k6 <= p79_k6;
    p80_bit_slice_2058870 <= p79_bit_slice_2058870;
    p80_array_index_2058900 <= p79_array_index_2058900;
    p80_array_index_2059029 <= p79_array_index_2059029;
    p80_array_index_2059054 <= p79_array_index_2059054;
    p80_res7__1069 <= p79_res7__1069;
    p80_array_index_2059077 <= p79_array_index_2059077;
    p80_res7__1073 <= p80_res7__1073_comb;
    p80_array_index_2059242 <= p80_array_index_2059242_comb;
    p80_array_index_2059261 <= p80_array_index_2059261_comb;
    p80_array_index_2059294 <= p80_array_index_2059294_comb;
    p80_array_index_2059295 <= p80_array_index_2059295_comb;
    p80_array_index_2059296 <= p80_array_index_2059296_comb;
    p80_array_index_2059297 <= p80_array_index_2059297_comb;
    p80_array_index_2059298 <= p80_array_index_2059298_comb;
    p80_array_index_2059299 <= p80_array_index_2059299_comb;
    p80_array_index_2059300 <= p80_array_index_2059300_comb;
    p80_array_index_2059301 <= p80_array_index_2059301_comb;
    p80_array_index_2059302 <= p80_array_index_2059302_comb;
    p80_array_index_2059303 <= p80_array_index_2059303_comb;
    p80_array_index_2059304 <= p80_array_index_2059304_comb;
    p80_array_index_2059305 <= p80_array_index_2059305_comb;
    p80_array_index_2059306 <= p80_array_index_2059306_comb;
    p80_array_index_2059307 <= p80_array_index_2059307_comb;
    p80_array_index_2059308 <= p80_array_index_2059308_comb;
    p80_array_index_2059309 <= p80_array_index_2059309_comb;
    p80_array_index_2059310 <= p80_array_index_2059310_comb;
    p80_array_index_2059311 <= p80_array_index_2059311_comb;
    p80_array_index_2059312 <= p80_array_index_2059312_comb;
    p80_array_index_2059313 <= p80_array_index_2059313_comb;
    p81_literal_2043910 <= p80_literal_2043910;
    p81_literal_2043912 <= p80_literal_2043912;
    p81_literal_2043914 <= p80_literal_2043914;
    p81_literal_2043916 <= p80_literal_2043916;
    p81_literal_2043918 <= p80_literal_2043918;
    p81_literal_2043920 <= p80_literal_2043920;
    p81_literal_2043923 <= p80_literal_2043923;
  end

  // ===== Pipe stage 81:
  wire [7:0] p81_res7__1087_comb;
  wire [127:0] p81_permut__33_comb;
  wire [127:0] p81_xor_2059409_comb;
  wire [7:0] p81_bit_slice_2059414_comb;
  wire [7:0] p81_bit_slice_2059415_comb;
  wire [7:0] p81_bit_slice_2059416_comb;
  wire [7:0] p81_bit_slice_2059417_comb;
  wire [7:0] p81_bit_slice_2059418_comb;
  wire [7:0] p81_bit_slice_2059419_comb;
  wire [7:0] p81_bit_slice_2059420_comb;
  wire [7:0] p81_bit_slice_2059421_comb;
  wire [7:0] p81_bit_slice_2059422_comb;
  wire [7:0] p81_bit_slice_2059429_comb;
  wire [7:0] p81_bit_slice_2059431_comb;
  wire [7:0] p81_array_index_2059432_comb;
  wire [7:0] p81_array_index_2059433_comb;
  wire [7:0] p81_array_index_2059434_comb;
  wire [7:0] p81_array_index_2059435_comb;
  wire [7:0] p81_array_index_2059436_comb;
  wire [7:0] p81_array_index_2059437_comb;
  wire [7:0] p81_res7__1089_comb;
  wire [7:0] p81_array_index_2059447_comb;
  wire [7:0] p81_array_index_2059448_comb;
  wire [7:0] p81_array_index_2059449_comb;
  wire [7:0] p81_array_index_2059450_comb;
  wire [7:0] p81_array_index_2059451_comb;
  wire [7:0] p81_array_index_2059452_comb;
  wire [7:0] p81_res7__1091_comb;
  wire [7:0] p81_array_index_2059461_comb;
  wire [7:0] p81_array_index_2059462_comb;
  wire [7:0] p81_array_index_2059463_comb;
  wire [7:0] p81_array_index_2059464_comb;
  wire [7:0] p81_array_index_2059465_comb;
  wire [7:0] p81_res7__1093_comb;
  wire [7:0] p81_array_index_2059475_comb;
  wire [7:0] p81_array_index_2059476_comb;
  wire [7:0] p81_array_index_2059477_comb;
  wire [7:0] p81_array_index_2059478_comb;
  wire [7:0] p81_array_index_2059479_comb;
  wire [7:0] p81_res7__1095_comb;
  wire [7:0] p81_array_index_2059488_comb;
  wire [7:0] p81_array_index_2059489_comb;
  wire [7:0] p81_array_index_2059490_comb;
  wire [7:0] p81_array_index_2059491_comb;
  wire [7:0] p81_res7__1097_comb;
  wire [7:0] p81_array_index_2059495_comb;
  wire [7:0] p81_array_index_2059496_comb;
  wire [7:0] p81_array_index_2059497_comb;
  wire [7:0] p81_array_index_2059498_comb;
  wire [7:0] p81_array_index_2059499_comb;
  wire [7:0] p81_array_index_2059500_comb;
  wire [7:0] p81_array_index_2059501_comb;
  wire [7:0] p81_array_index_2059502_comb;
  wire [7:0] p81_array_index_2059503_comb;
  wire [7:0] p81_array_index_2059504_comb;
  wire [7:0] p81_array_index_2059505_comb;
  wire [7:0] p81_array_index_2059506_comb;
  assign p81_res7__1087_comb = p80_array_index_2058900 ^ p80_array_index_2059029 ^ p80_array_index_2059054 ^ p80_array_index_2059077 ^ p80_array_index_2059242 ^ p80_array_index_2059261 ^ p80_res7__1069 ^ p80_array_index_2059294 ^ p80_res7__1073 ^ p80_array_index_2059295 ^ p80_array_index_2059296 ^ p80_array_index_2059297 ^ p80_array_index_2059298 ^ p80_array_index_2059299 ^ p80_array_index_2059300 ^ p80_bit_slice_2058870;
  assign p81_permut__33_comb = {p80_array_index_2059301, p80_array_index_2059302, p80_array_index_2059303, p80_array_index_2059304, p80_array_index_2059305, p80_array_index_2059306, p80_literal_2058836[p80_res7__1069], p80_array_index_2059307, p80_literal_2058836[p80_res7__1073], p80_array_index_2059308, p80_array_index_2059309, p80_array_index_2059310, p80_array_index_2059311, p80_array_index_2059312, p80_array_index_2059313, p80_literal_2058836[p81_res7__1087_comb]};
  assign p81_xor_2059409_comb = p80_k7 ^ p81_permut__33_comb;
  assign p81_bit_slice_2059414_comb = p81_xor_2059409_comb[87:80];
  assign p81_bit_slice_2059415_comb = p81_xor_2059409_comb[79:72];
  assign p81_bit_slice_2059416_comb = p81_xor_2059409_comb[63:56];
  assign p81_bit_slice_2059417_comb = p81_xor_2059409_comb[47:40];
  assign p81_bit_slice_2059418_comb = p81_xor_2059409_comb[39:32];
  assign p81_bit_slice_2059419_comb = p81_xor_2059409_comb[31:24];
  assign p81_bit_slice_2059420_comb = p81_xor_2059409_comb[23:16];
  assign p81_bit_slice_2059421_comb = p81_xor_2059409_comb[15:8];
  assign p81_bit_slice_2059422_comb = p81_xor_2059409_comb[7:0];
  assign p81_bit_slice_2059429_comb = p81_xor_2059409_comb[71:64];
  assign p81_bit_slice_2059431_comb = p81_xor_2059409_comb[55:48];
  assign p81_array_index_2059432_comb = p80_literal_2043920[p81_bit_slice_2059417_comb];
  assign p81_array_index_2059433_comb = p80_literal_2043918[p81_bit_slice_2059418_comb];
  assign p81_array_index_2059434_comb = p80_literal_2043916[p81_bit_slice_2059419_comb];
  assign p81_array_index_2059435_comb = p80_literal_2043914[p81_bit_slice_2059420_comb];
  assign p81_array_index_2059436_comb = p80_literal_2043912[p81_bit_slice_2059421_comb];
  assign p81_array_index_2059437_comb = p80_literal_2043910[p81_bit_slice_2059422_comb];
  assign p81_res7__1089_comb = p80_literal_2043910[p81_xor_2059409_comb[119:112]] ^ p80_literal_2043912[p81_xor_2059409_comb[111:104]] ^ p80_literal_2043914[p81_xor_2059409_comb[103:96]] ^ p80_literal_2043916[p81_xor_2059409_comb[95:88]] ^ p80_literal_2043918[p81_bit_slice_2059414_comb] ^ p80_literal_2043920[p81_bit_slice_2059415_comb] ^ p81_bit_slice_2059429_comb ^ p80_literal_2043923[p81_bit_slice_2059416_comb] ^ p81_bit_slice_2059431_comb ^ p81_array_index_2059432_comb ^ p81_array_index_2059433_comb ^ p81_array_index_2059434_comb ^ p81_array_index_2059435_comb ^ p81_array_index_2059436_comb ^ p81_array_index_2059437_comb ^ p81_xor_2059409_comb[127:120];
  assign p81_array_index_2059447_comb = p80_literal_2043920[p81_bit_slice_2059418_comb];
  assign p81_array_index_2059448_comb = p80_literal_2043918[p81_bit_slice_2059419_comb];
  assign p81_array_index_2059449_comb = p80_literal_2043916[p81_bit_slice_2059420_comb];
  assign p81_array_index_2059450_comb = p80_literal_2043914[p81_bit_slice_2059421_comb];
  assign p81_array_index_2059451_comb = p80_literal_2043912[p81_bit_slice_2059422_comb];
  assign p81_array_index_2059452_comb = p80_literal_2043910[p81_res7__1089_comb];
  assign p81_res7__1091_comb = p80_literal_2043910[p81_xor_2059409_comb[111:104]] ^ p80_literal_2043912[p81_xor_2059409_comb[103:96]] ^ p80_literal_2043914[p81_xor_2059409_comb[95:88]] ^ p80_literal_2043916[p81_bit_slice_2059414_comb] ^ p80_literal_2043918[p81_bit_slice_2059415_comb] ^ p80_literal_2043920[p81_bit_slice_2059429_comb] ^ p81_bit_slice_2059416_comb ^ p80_literal_2043923[p81_bit_slice_2059431_comb] ^ p81_bit_slice_2059417_comb ^ p81_array_index_2059447_comb ^ p81_array_index_2059448_comb ^ p81_array_index_2059449_comb ^ p81_array_index_2059450_comb ^ p81_array_index_2059451_comb ^ p81_array_index_2059452_comb ^ p81_xor_2059409_comb[119:112];
  assign p81_array_index_2059461_comb = p80_literal_2043920[p81_bit_slice_2059419_comb];
  assign p81_array_index_2059462_comb = p80_literal_2043918[p81_bit_slice_2059420_comb];
  assign p81_array_index_2059463_comb = p80_literal_2043916[p81_bit_slice_2059421_comb];
  assign p81_array_index_2059464_comb = p80_literal_2043914[p81_bit_slice_2059422_comb];
  assign p81_array_index_2059465_comb = p80_literal_2043912[p81_res7__1089_comb];
  assign p81_res7__1093_comb = p80_literal_2043910[p81_xor_2059409_comb[103:96]] ^ p80_literal_2043912[p81_xor_2059409_comb[95:88]] ^ p80_literal_2043914[p81_bit_slice_2059414_comb] ^ p80_literal_2043916[p81_bit_slice_2059415_comb] ^ p80_literal_2043918[p81_bit_slice_2059429_comb] ^ p80_literal_2043920[p81_bit_slice_2059416_comb] ^ p81_bit_slice_2059431_comb ^ p80_literal_2043923[p81_bit_slice_2059417_comb] ^ p81_bit_slice_2059418_comb ^ p81_array_index_2059461_comb ^ p81_array_index_2059462_comb ^ p81_array_index_2059463_comb ^ p81_array_index_2059464_comb ^ p81_array_index_2059465_comb ^ p80_literal_2043910[p81_res7__1091_comb] ^ p81_xor_2059409_comb[111:104];
  assign p81_array_index_2059475_comb = p80_literal_2043920[p81_bit_slice_2059420_comb];
  assign p81_array_index_2059476_comb = p80_literal_2043918[p81_bit_slice_2059421_comb];
  assign p81_array_index_2059477_comb = p80_literal_2043916[p81_bit_slice_2059422_comb];
  assign p81_array_index_2059478_comb = p80_literal_2043914[p81_res7__1089_comb];
  assign p81_array_index_2059479_comb = p80_literal_2043912[p81_res7__1091_comb];
  assign p81_res7__1095_comb = p80_literal_2043910[p81_xor_2059409_comb[95:88]] ^ p80_literal_2043912[p81_bit_slice_2059414_comb] ^ p80_literal_2043914[p81_bit_slice_2059415_comb] ^ p80_literal_2043916[p81_bit_slice_2059429_comb] ^ p80_literal_2043918[p81_bit_slice_2059416_comb] ^ p80_literal_2043920[p81_bit_slice_2059431_comb] ^ p81_bit_slice_2059417_comb ^ p80_literal_2043923[p81_bit_slice_2059418_comb] ^ p81_bit_slice_2059419_comb ^ p81_array_index_2059475_comb ^ p81_array_index_2059476_comb ^ p81_array_index_2059477_comb ^ p81_array_index_2059478_comb ^ p81_array_index_2059479_comb ^ p80_literal_2043910[p81_res7__1093_comb] ^ p81_xor_2059409_comb[103:96];
  assign p81_array_index_2059488_comb = p80_literal_2043920[p81_bit_slice_2059421_comb];
  assign p81_array_index_2059489_comb = p80_literal_2043918[p81_bit_slice_2059422_comb];
  assign p81_array_index_2059490_comb = p80_literal_2043916[p81_res7__1089_comb];
  assign p81_array_index_2059491_comb = p80_literal_2043914[p81_res7__1091_comb];
  assign p81_res7__1097_comb = p80_literal_2043910[p81_bit_slice_2059414_comb] ^ p80_literal_2043912[p81_bit_slice_2059415_comb] ^ p80_literal_2043914[p81_bit_slice_2059429_comb] ^ p80_literal_2043916[p81_bit_slice_2059416_comb] ^ p80_literal_2043918[p81_bit_slice_2059431_comb] ^ p81_array_index_2059432_comb ^ p81_bit_slice_2059418_comb ^ p80_literal_2043923[p81_bit_slice_2059419_comb] ^ p81_bit_slice_2059420_comb ^ p81_array_index_2059488_comb ^ p81_array_index_2059489_comb ^ p81_array_index_2059490_comb ^ p81_array_index_2059491_comb ^ p80_literal_2043912[p81_res7__1093_comb] ^ p80_literal_2043910[p81_res7__1095_comb] ^ p81_xor_2059409_comb[95:88];
  assign p81_array_index_2059495_comb = p80_literal_2043910[p81_bit_slice_2059415_comb];
  assign p81_array_index_2059496_comb = p80_literal_2043912[p81_bit_slice_2059429_comb];
  assign p81_array_index_2059497_comb = p80_literal_2043914[p81_bit_slice_2059416_comb];
  assign p81_array_index_2059498_comb = p80_literal_2043916[p81_bit_slice_2059431_comb];
  assign p81_array_index_2059499_comb = p80_literal_2043918[p81_bit_slice_2059417_comb];
  assign p81_array_index_2059500_comb = p80_literal_2043923[p81_bit_slice_2059420_comb];
  assign p81_array_index_2059501_comb = p80_literal_2043920[p81_bit_slice_2059422_comb];
  assign p81_array_index_2059502_comb = p80_literal_2043918[p81_res7__1089_comb];
  assign p81_array_index_2059503_comb = p80_literal_2043916[p81_res7__1091_comb];
  assign p81_array_index_2059504_comb = p80_literal_2043914[p81_res7__1093_comb];
  assign p81_array_index_2059505_comb = p80_literal_2043912[p81_res7__1095_comb];
  assign p81_array_index_2059506_comb = p80_literal_2043910[p81_res7__1097_comb];

  // Registers for pipe stage 81:
  reg [127:0] p81_bit_slice_2043893;
  reg [127:0] p81_bit_slice_2044018;
  reg [127:0] p81_k3;
  reg [127:0] p81_k2;
  reg [127:0] p81_k5;
  reg [127:0] p81_k4;
  reg [127:0] p81_k6;
  reg [7:0] p81_bit_slice_2059414;
  reg [7:0] p81_bit_slice_2059415;
  reg [7:0] p81_bit_slice_2059416;
  reg [7:0] p81_bit_slice_2059417;
  reg [7:0] p81_bit_slice_2059418;
  reg [7:0] p81_bit_slice_2059419;
  reg [7:0] p81_bit_slice_2059420;
  reg [7:0] p81_bit_slice_2059421;
  reg [7:0] p81_bit_slice_2059422;
  reg [7:0] p81_bit_slice_2059429;
  reg [7:0] p81_bit_slice_2059431;
  reg [7:0] p81_array_index_2059433;
  reg [7:0] p81_array_index_2059434;
  reg [7:0] p81_array_index_2059435;
  reg [7:0] p81_array_index_2059436;
  reg [7:0] p81_array_index_2059437;
  reg [7:0] p81_res7__1089;
  reg [7:0] p81_array_index_2059447;
  reg [7:0] p81_array_index_2059448;
  reg [7:0] p81_array_index_2059449;
  reg [7:0] p81_array_index_2059450;
  reg [7:0] p81_array_index_2059451;
  reg [7:0] p81_array_index_2059452;
  reg [7:0] p81_res7__1091;
  reg [7:0] p81_array_index_2059461;
  reg [7:0] p81_array_index_2059462;
  reg [7:0] p81_array_index_2059463;
  reg [7:0] p81_array_index_2059464;
  reg [7:0] p81_array_index_2059465;
  reg [7:0] p81_res7__1093;
  reg [7:0] p81_array_index_2059475;
  reg [7:0] p81_array_index_2059476;
  reg [7:0] p81_array_index_2059477;
  reg [7:0] p81_array_index_2059478;
  reg [7:0] p81_array_index_2059479;
  reg [7:0] p81_res7__1095;
  reg [7:0] p81_array_index_2059488;
  reg [7:0] p81_array_index_2059489;
  reg [7:0] p81_array_index_2059490;
  reg [7:0] p81_array_index_2059491;
  reg [7:0] p81_res7__1097;
  reg [7:0] p81_array_index_2059495;
  reg [7:0] p81_array_index_2059496;
  reg [7:0] p81_array_index_2059497;
  reg [7:0] p81_array_index_2059498;
  reg [7:0] p81_array_index_2059499;
  reg [7:0] p81_array_index_2059500;
  reg [7:0] p81_array_index_2059501;
  reg [7:0] p81_array_index_2059502;
  reg [7:0] p81_array_index_2059503;
  reg [7:0] p81_array_index_2059504;
  reg [7:0] p81_array_index_2059505;
  reg [7:0] p81_array_index_2059506;
  reg [7:0] p82_literal_2043910[256];
  reg [7:0] p82_literal_2043912[256];
  reg [7:0] p82_literal_2043914[256];
  reg [7:0] p82_literal_2043916[256];
  reg [7:0] p82_literal_2043918[256];
  reg [7:0] p82_literal_2043920[256];
  reg [7:0] p82_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p81_bit_slice_2043893 <= p80_bit_slice_2043893;
    p81_bit_slice_2044018 <= p80_bit_slice_2044018;
    p81_k3 <= p80_k3;
    p81_k2 <= p80_k2;
    p81_k5 <= p80_k5;
    p81_k4 <= p80_k4;
    p81_k6 <= p80_k6;
    p81_bit_slice_2059414 <= p81_bit_slice_2059414_comb;
    p81_bit_slice_2059415 <= p81_bit_slice_2059415_comb;
    p81_bit_slice_2059416 <= p81_bit_slice_2059416_comb;
    p81_bit_slice_2059417 <= p81_bit_slice_2059417_comb;
    p81_bit_slice_2059418 <= p81_bit_slice_2059418_comb;
    p81_bit_slice_2059419 <= p81_bit_slice_2059419_comb;
    p81_bit_slice_2059420 <= p81_bit_slice_2059420_comb;
    p81_bit_slice_2059421 <= p81_bit_slice_2059421_comb;
    p81_bit_slice_2059422 <= p81_bit_slice_2059422_comb;
    p81_bit_slice_2059429 <= p81_bit_slice_2059429_comb;
    p81_bit_slice_2059431 <= p81_bit_slice_2059431_comb;
    p81_array_index_2059433 <= p81_array_index_2059433_comb;
    p81_array_index_2059434 <= p81_array_index_2059434_comb;
    p81_array_index_2059435 <= p81_array_index_2059435_comb;
    p81_array_index_2059436 <= p81_array_index_2059436_comb;
    p81_array_index_2059437 <= p81_array_index_2059437_comb;
    p81_res7__1089 <= p81_res7__1089_comb;
    p81_array_index_2059447 <= p81_array_index_2059447_comb;
    p81_array_index_2059448 <= p81_array_index_2059448_comb;
    p81_array_index_2059449 <= p81_array_index_2059449_comb;
    p81_array_index_2059450 <= p81_array_index_2059450_comb;
    p81_array_index_2059451 <= p81_array_index_2059451_comb;
    p81_array_index_2059452 <= p81_array_index_2059452_comb;
    p81_res7__1091 <= p81_res7__1091_comb;
    p81_array_index_2059461 <= p81_array_index_2059461_comb;
    p81_array_index_2059462 <= p81_array_index_2059462_comb;
    p81_array_index_2059463 <= p81_array_index_2059463_comb;
    p81_array_index_2059464 <= p81_array_index_2059464_comb;
    p81_array_index_2059465 <= p81_array_index_2059465_comb;
    p81_res7__1093 <= p81_res7__1093_comb;
    p81_array_index_2059475 <= p81_array_index_2059475_comb;
    p81_array_index_2059476 <= p81_array_index_2059476_comb;
    p81_array_index_2059477 <= p81_array_index_2059477_comb;
    p81_array_index_2059478 <= p81_array_index_2059478_comb;
    p81_array_index_2059479 <= p81_array_index_2059479_comb;
    p81_res7__1095 <= p81_res7__1095_comb;
    p81_array_index_2059488 <= p81_array_index_2059488_comb;
    p81_array_index_2059489 <= p81_array_index_2059489_comb;
    p81_array_index_2059490 <= p81_array_index_2059490_comb;
    p81_array_index_2059491 <= p81_array_index_2059491_comb;
    p81_res7__1097 <= p81_res7__1097_comb;
    p81_array_index_2059495 <= p81_array_index_2059495_comb;
    p81_array_index_2059496 <= p81_array_index_2059496_comb;
    p81_array_index_2059497 <= p81_array_index_2059497_comb;
    p81_array_index_2059498 <= p81_array_index_2059498_comb;
    p81_array_index_2059499 <= p81_array_index_2059499_comb;
    p81_array_index_2059500 <= p81_array_index_2059500_comb;
    p81_array_index_2059501 <= p81_array_index_2059501_comb;
    p81_array_index_2059502 <= p81_array_index_2059502_comb;
    p81_array_index_2059503 <= p81_array_index_2059503_comb;
    p81_array_index_2059504 <= p81_array_index_2059504_comb;
    p81_array_index_2059505 <= p81_array_index_2059505_comb;
    p81_array_index_2059506 <= p81_array_index_2059506_comb;
    p82_literal_2043910 <= p81_literal_2043910;
    p82_literal_2043912 <= p81_literal_2043912;
    p82_literal_2043914 <= p81_literal_2043914;
    p82_literal_2043916 <= p81_literal_2043916;
    p82_literal_2043918 <= p81_literal_2043918;
    p82_literal_2043920 <= p81_literal_2043920;
    p82_literal_2043923 <= p81_literal_2043923;
  end

  // ===== Pipe stage 82:
  wire [7:0] p82_res7__1099_comb;
  wire [7:0] p82_array_index_2059649_comb;
  wire [7:0] p82_array_index_2059650_comb;
  wire [7:0] p82_array_index_2059651_comb;
  wire [7:0] p82_res7__1101_comb;
  wire [7:0] p82_array_index_2059661_comb;
  wire [7:0] p82_array_index_2059662_comb;
  wire [7:0] p82_array_index_2059663_comb;
  wire [7:0] p82_res7__1103_comb;
  wire [7:0] p82_array_index_2059672_comb;
  wire [7:0] p82_array_index_2059673_comb;
  wire [7:0] p82_res7__1105_comb;
  wire [7:0] p82_array_index_2059683_comb;
  wire [7:0] p82_array_index_2059684_comb;
  wire [7:0] p82_res7__1107_comb;
  wire [7:0] p82_array_index_2059693_comb;
  wire [7:0] p82_res7__1109_comb;
  wire [7:0] p82_array_index_2059703_comb;
  wire [7:0] p82_res7__1111_comb;
  wire [7:0] p82_array_index_2059710_comb;
  wire [7:0] p82_array_index_2059711_comb;
  wire [7:0] p82_array_index_2059712_comb;
  wire [7:0] p82_array_index_2059713_comb;
  wire [7:0] p82_array_index_2059714_comb;
  wire [7:0] p82_array_index_2059715_comb;
  wire [7:0] p82_array_index_2059716_comb;
  wire [7:0] p82_array_index_2059717_comb;
  wire [7:0] p82_array_index_2059718_comb;
  wire [7:0] p82_array_index_2059719_comb;
  wire [7:0] p82_array_index_2059720_comb;
  assign p82_res7__1099_comb = p81_array_index_2059495 ^ p81_array_index_2059496 ^ p81_array_index_2059497 ^ p81_array_index_2059498 ^ p81_array_index_2059499 ^ p81_array_index_2059447 ^ p81_bit_slice_2059419 ^ p81_array_index_2059500 ^ p81_bit_slice_2059421 ^ p81_array_index_2059501 ^ p81_array_index_2059502 ^ p81_array_index_2059503 ^ p81_array_index_2059504 ^ p81_array_index_2059505 ^ p81_array_index_2059506 ^ p81_bit_slice_2059414;
  assign p82_array_index_2059649_comb = p81_literal_2043920[p81_res7__1089];
  assign p82_array_index_2059650_comb = p81_literal_2043918[p81_res7__1091];
  assign p82_array_index_2059651_comb = p81_literal_2043916[p81_res7__1093];
  assign p82_res7__1101_comb = p81_literal_2043910[p81_bit_slice_2059429] ^ p81_literal_2043912[p81_bit_slice_2059416] ^ p81_literal_2043914[p81_bit_slice_2059431] ^ p81_literal_2043916[p81_bit_slice_2059417] ^ p81_array_index_2059433 ^ p81_array_index_2059461 ^ p81_bit_slice_2059420 ^ p81_literal_2043923[p81_bit_slice_2059421] ^ p81_bit_slice_2059422 ^ p82_array_index_2059649_comb ^ p82_array_index_2059650_comb ^ p82_array_index_2059651_comb ^ p81_literal_2043914[p81_res7__1095] ^ p81_literal_2043912[p81_res7__1097] ^ p81_literal_2043910[p82_res7__1099_comb] ^ p81_bit_slice_2059415;
  assign p82_array_index_2059661_comb = p81_literal_2043920[p81_res7__1091];
  assign p82_array_index_2059662_comb = p81_literal_2043918[p81_res7__1093];
  assign p82_array_index_2059663_comb = p81_literal_2043916[p81_res7__1095];
  assign p82_res7__1103_comb = p81_literal_2043910[p81_bit_slice_2059416] ^ p81_literal_2043912[p81_bit_slice_2059431] ^ p81_literal_2043914[p81_bit_slice_2059417] ^ p81_literal_2043916[p81_bit_slice_2059418] ^ p81_array_index_2059448 ^ p81_array_index_2059475 ^ p81_bit_slice_2059421 ^ p81_literal_2043923[p81_bit_slice_2059422] ^ p81_res7__1089 ^ p82_array_index_2059661_comb ^ p82_array_index_2059662_comb ^ p82_array_index_2059663_comb ^ p81_literal_2043914[p81_res7__1097] ^ p81_literal_2043912[p82_res7__1099_comb] ^ p81_literal_2043910[p82_res7__1101_comb] ^ p81_bit_slice_2059429;
  assign p82_array_index_2059672_comb = p81_literal_2043920[p81_res7__1093];
  assign p82_array_index_2059673_comb = p81_literal_2043918[p81_res7__1095];
  assign p82_res7__1105_comb = p81_literal_2043910[p81_bit_slice_2059431] ^ p81_literal_2043912[p81_bit_slice_2059417] ^ p81_literal_2043914[p81_bit_slice_2059418] ^ p81_array_index_2059434 ^ p81_array_index_2059462 ^ p81_array_index_2059488 ^ p81_bit_slice_2059422 ^ p81_literal_2043923[p81_res7__1089] ^ p81_res7__1091 ^ p82_array_index_2059672_comb ^ p82_array_index_2059673_comb ^ p81_literal_2043916[p81_res7__1097] ^ p81_literal_2043914[p82_res7__1099_comb] ^ p81_literal_2043912[p82_res7__1101_comb] ^ p81_literal_2043910[p82_res7__1103_comb] ^ p81_bit_slice_2059416;
  assign p82_array_index_2059683_comb = p81_literal_2043920[p81_res7__1095];
  assign p82_array_index_2059684_comb = p81_literal_2043918[p81_res7__1097];
  assign p82_res7__1107_comb = p81_literal_2043910[p81_bit_slice_2059417] ^ p81_literal_2043912[p81_bit_slice_2059418] ^ p81_literal_2043914[p81_bit_slice_2059419] ^ p81_array_index_2059449 ^ p81_array_index_2059476 ^ p81_array_index_2059501 ^ p81_res7__1089 ^ p81_literal_2043923[p81_res7__1091] ^ p81_res7__1093 ^ p82_array_index_2059683_comb ^ p82_array_index_2059684_comb ^ p81_literal_2043916[p82_res7__1099_comb] ^ p81_literal_2043914[p82_res7__1101_comb] ^ p81_literal_2043912[p82_res7__1103_comb] ^ p81_literal_2043910[p82_res7__1105_comb] ^ p81_bit_slice_2059431;
  assign p82_array_index_2059693_comb = p81_literal_2043920[p81_res7__1097];
  assign p82_res7__1109_comb = p81_literal_2043910[p81_bit_slice_2059418] ^ p81_literal_2043912[p81_bit_slice_2059419] ^ p81_array_index_2059435 ^ p81_array_index_2059463 ^ p81_array_index_2059489 ^ p82_array_index_2059649_comb ^ p81_res7__1091 ^ p81_literal_2043923[p81_res7__1093] ^ p81_res7__1095 ^ p82_array_index_2059693_comb ^ p81_literal_2043918[p82_res7__1099_comb] ^ p81_literal_2043916[p82_res7__1101_comb] ^ p81_literal_2043914[p82_res7__1103_comb] ^ p81_literal_2043912[p82_res7__1105_comb] ^ p81_literal_2043910[p82_res7__1107_comb] ^ p81_bit_slice_2059417;
  assign p82_array_index_2059703_comb = p81_literal_2043920[p82_res7__1099_comb];
  assign p82_res7__1111_comb = p81_literal_2043910[p81_bit_slice_2059419] ^ p81_literal_2043912[p81_bit_slice_2059420] ^ p81_array_index_2059450 ^ p81_array_index_2059477 ^ p81_array_index_2059502 ^ p82_array_index_2059661_comb ^ p81_res7__1093 ^ p81_literal_2043923[p81_res7__1095] ^ p81_res7__1097 ^ p82_array_index_2059703_comb ^ p81_literal_2043918[p82_res7__1101_comb] ^ p81_literal_2043916[p82_res7__1103_comb] ^ p81_literal_2043914[p82_res7__1105_comb] ^ p81_literal_2043912[p82_res7__1107_comb] ^ p81_literal_2043910[p82_res7__1109_comb] ^ p81_bit_slice_2059418;
  assign p82_array_index_2059710_comb = p81_literal_2043910[p81_bit_slice_2059420];
  assign p82_array_index_2059711_comb = p81_literal_2043923[p81_res7__1097];
  assign p82_array_index_2059712_comb = p81_literal_2043920[p82_res7__1101_comb];
  assign p82_array_index_2059713_comb = p81_literal_2043918[p82_res7__1103_comb];
  assign p82_array_index_2059714_comb = p81_literal_2043916[p82_res7__1105_comb];
  assign p82_array_index_2059715_comb = p81_literal_2043914[p82_res7__1107_comb];
  assign p82_array_index_2059716_comb = p81_literal_2043912[p82_res7__1109_comb];
  assign p82_array_index_2059717_comb = p81_literal_2043910[p82_res7__1111_comb];
  assign p82_array_index_2059718_comb = p81_literal_2058836[p81_res7__1089];
  assign p82_array_index_2059719_comb = p81_literal_2058836[p81_res7__1091];
  assign p82_array_index_2059720_comb = p81_literal_2058836[p81_res7__1093];

  // Registers for pipe stage 82:
  reg [127:0] p82_bit_slice_2043893;
  reg [127:0] p82_bit_slice_2044018;
  reg [127:0] p82_k3;
  reg [127:0] p82_k2;
  reg [127:0] p82_k5;
  reg [127:0] p82_k4;
  reg [127:0] p82_k6;
  reg [7:0] p82_bit_slice_2059419;
  reg [7:0] p82_bit_slice_2059420;
  reg [7:0] p82_bit_slice_2059421;
  reg [7:0] p82_bit_slice_2059422;
  reg [7:0] p82_array_index_2059436;
  reg [7:0] p82_array_index_2059437;
  reg [7:0] p82_array_index_2059451;
  reg [7:0] p82_array_index_2059452;
  reg [7:0] p82_array_index_2059464;
  reg [7:0] p82_array_index_2059465;
  reg [7:0] p82_array_index_2059478;
  reg [7:0] p82_array_index_2059479;
  reg [7:0] p82_res7__1095;
  reg [7:0] p82_array_index_2059490;
  reg [7:0] p82_array_index_2059491;
  reg [7:0] p82_res7__1097;
  reg [7:0] p82_array_index_2059503;
  reg [7:0] p82_array_index_2059504;
  reg [7:0] p82_res7__1099;
  reg [7:0] p82_array_index_2059650;
  reg [7:0] p82_array_index_2059651;
  reg [7:0] p82_res7__1101;
  reg [7:0] p82_array_index_2059662;
  reg [7:0] p82_array_index_2059663;
  reg [7:0] p82_res7__1103;
  reg [7:0] p82_array_index_2059672;
  reg [7:0] p82_array_index_2059673;
  reg [7:0] p82_res7__1105;
  reg [7:0] p82_array_index_2059683;
  reg [7:0] p82_array_index_2059684;
  reg [7:0] p82_res7__1107;
  reg [7:0] p82_array_index_2059693;
  reg [7:0] p82_res7__1109;
  reg [7:0] p82_array_index_2059703;
  reg [7:0] p82_res7__1111;
  reg [7:0] p82_array_index_2059710;
  reg [7:0] p82_array_index_2059711;
  reg [7:0] p82_array_index_2059712;
  reg [7:0] p82_array_index_2059713;
  reg [7:0] p82_array_index_2059714;
  reg [7:0] p82_array_index_2059715;
  reg [7:0] p82_array_index_2059716;
  reg [7:0] p82_array_index_2059717;
  reg [7:0] p82_array_index_2059718;
  reg [7:0] p82_array_index_2059719;
  reg [7:0] p82_array_index_2059720;
  reg [7:0] p83_literal_2043910[256];
  reg [7:0] p83_literal_2043912[256];
  reg [7:0] p83_literal_2043914[256];
  reg [7:0] p83_literal_2043916[256];
  reg [7:0] p83_literal_2043918[256];
  reg [7:0] p83_literal_2043920[256];
  reg [7:0] p83_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p82_bit_slice_2043893 <= p81_bit_slice_2043893;
    p82_bit_slice_2044018 <= p81_bit_slice_2044018;
    p82_k3 <= p81_k3;
    p82_k2 <= p81_k2;
    p82_k5 <= p81_k5;
    p82_k4 <= p81_k4;
    p82_k6 <= p81_k6;
    p82_bit_slice_2059419 <= p81_bit_slice_2059419;
    p82_bit_slice_2059420 <= p81_bit_slice_2059420;
    p82_bit_slice_2059421 <= p81_bit_slice_2059421;
    p82_bit_slice_2059422 <= p81_bit_slice_2059422;
    p82_array_index_2059436 <= p81_array_index_2059436;
    p82_array_index_2059437 <= p81_array_index_2059437;
    p82_array_index_2059451 <= p81_array_index_2059451;
    p82_array_index_2059452 <= p81_array_index_2059452;
    p82_array_index_2059464 <= p81_array_index_2059464;
    p82_array_index_2059465 <= p81_array_index_2059465;
    p82_array_index_2059478 <= p81_array_index_2059478;
    p82_array_index_2059479 <= p81_array_index_2059479;
    p82_res7__1095 <= p81_res7__1095;
    p82_array_index_2059490 <= p81_array_index_2059490;
    p82_array_index_2059491 <= p81_array_index_2059491;
    p82_res7__1097 <= p81_res7__1097;
    p82_array_index_2059503 <= p81_array_index_2059503;
    p82_array_index_2059504 <= p81_array_index_2059504;
    p82_res7__1099 <= p82_res7__1099_comb;
    p82_array_index_2059650 <= p82_array_index_2059650_comb;
    p82_array_index_2059651 <= p82_array_index_2059651_comb;
    p82_res7__1101 <= p82_res7__1101_comb;
    p82_array_index_2059662 <= p82_array_index_2059662_comb;
    p82_array_index_2059663 <= p82_array_index_2059663_comb;
    p82_res7__1103 <= p82_res7__1103_comb;
    p82_array_index_2059672 <= p82_array_index_2059672_comb;
    p82_array_index_2059673 <= p82_array_index_2059673_comb;
    p82_res7__1105 <= p82_res7__1105_comb;
    p82_array_index_2059683 <= p82_array_index_2059683_comb;
    p82_array_index_2059684 <= p82_array_index_2059684_comb;
    p82_res7__1107 <= p82_res7__1107_comb;
    p82_array_index_2059693 <= p82_array_index_2059693_comb;
    p82_res7__1109 <= p82_res7__1109_comb;
    p82_array_index_2059703 <= p82_array_index_2059703_comb;
    p82_res7__1111 <= p82_res7__1111_comb;
    p82_array_index_2059710 <= p82_array_index_2059710_comb;
    p82_array_index_2059711 <= p82_array_index_2059711_comb;
    p82_array_index_2059712 <= p82_array_index_2059712_comb;
    p82_array_index_2059713 <= p82_array_index_2059713_comb;
    p82_array_index_2059714 <= p82_array_index_2059714_comb;
    p82_array_index_2059715 <= p82_array_index_2059715_comb;
    p82_array_index_2059716 <= p82_array_index_2059716_comb;
    p82_array_index_2059717 <= p82_array_index_2059717_comb;
    p82_array_index_2059718 <= p82_array_index_2059718_comb;
    p82_array_index_2059719 <= p82_array_index_2059719_comb;
    p82_array_index_2059720 <= p82_array_index_2059720_comb;
    p83_literal_2043910 <= p82_literal_2043910;
    p83_literal_2043912 <= p82_literal_2043912;
    p83_literal_2043914 <= p82_literal_2043914;
    p83_literal_2043916 <= p82_literal_2043916;
    p83_literal_2043918 <= p82_literal_2043918;
    p83_literal_2043920 <= p82_literal_2043920;
    p83_literal_2043923 <= p82_literal_2043923;
  end

  // ===== Pipe stage 83:
  wire [7:0] p83_res7__1113_comb;
  wire [7:0] p83_res7__1115_comb;
  wire [7:0] p83_res7__1117_comb;
  wire [7:0] p83_res7__1119_comb;
  wire [127:0] p83_permut__34_comb;
  wire [127:0] p83_xor_2059883_comb;
  wire [7:0] p83_bit_slice_2059885_comb;
  wire [7:0] p83_bit_slice_2059886_comb;
  wire [7:0] p83_bit_slice_2059887_comb;
  wire [7:0] p83_bit_slice_2059888_comb;
  wire [7:0] p83_bit_slice_2059889_comb;
  wire [7:0] p83_bit_slice_2059890_comb;
  wire [7:0] p83_bit_slice_2059891_comb;
  wire [7:0] p83_bit_slice_2059892_comb;
  wire [7:0] p83_bit_slice_2059893_comb;
  wire [7:0] p83_bit_slice_2059894_comb;
  wire [7:0] p83_bit_slice_2059895_comb;
  wire [7:0] p83_bit_slice_2059896_comb;
  wire [7:0] p83_bit_slice_2059903_comb;
  wire [7:0] p83_bit_slice_2059905_comb;
  wire [7:0] p83_array_index_2059906_comb;
  wire [7:0] p83_array_index_2059907_comb;
  wire [7:0] p83_array_index_2059908_comb;
  wire [7:0] p83_array_index_2059909_comb;
  wire [7:0] p83_array_index_2059910_comb;
  wire [7:0] p83_array_index_2059911_comb;
  wire [7:0] p83_res7__1121_comb;
  wire [7:0] p83_array_index_2059921_comb;
  wire [7:0] p83_array_index_2059922_comb;
  wire [7:0] p83_array_index_2059923_comb;
  wire [7:0] p83_array_index_2059924_comb;
  wire [7:0] p83_array_index_2059925_comb;
  wire [7:0] p83_array_index_2059926_comb;
  wire [7:0] p83_res7__1123_comb;
  wire [7:0] p83_array_index_2059928_comb;
  wire [7:0] p83_array_index_2059929_comb;
  wire [7:0] p83_array_index_2059930_comb;
  wire [7:0] p83_array_index_2059931_comb;
  wire [7:0] p83_array_index_2059932_comb;
  wire [7:0] p83_array_index_2059933_comb;
  wire [7:0] p83_array_index_2059934_comb;
  wire [7:0] p83_array_index_2059935_comb;
  wire [7:0] p83_array_index_2059936_comb;
  wire [7:0] p83_array_index_2059937_comb;
  wire [7:0] p83_array_index_2059938_comb;
  wire [7:0] p83_array_index_2059939_comb;
  wire [7:0] p83_array_index_2059940_comb;
  assign p83_res7__1113_comb = p82_array_index_2059710 ^ p82_array_index_2059436 ^ p82_array_index_2059464 ^ p82_array_index_2059490 ^ p82_array_index_2059650 ^ p82_array_index_2059672 ^ p82_res7__1095 ^ p82_array_index_2059711 ^ p82_res7__1099 ^ p82_array_index_2059712 ^ p82_array_index_2059713 ^ p82_array_index_2059714 ^ p82_array_index_2059715 ^ p82_array_index_2059716 ^ p82_array_index_2059717 ^ p82_bit_slice_2059419;
  assign p83_res7__1115_comb = p82_literal_2043910[p82_bit_slice_2059421] ^ p82_array_index_2059451 ^ p82_array_index_2059478 ^ p82_array_index_2059503 ^ p82_array_index_2059662 ^ p82_array_index_2059683 ^ p82_res7__1097 ^ p82_literal_2043923[p82_res7__1099] ^ p82_res7__1101 ^ p82_literal_2043920[p82_res7__1103] ^ p82_literal_2043918[p82_res7__1105] ^ p82_literal_2043916[p82_res7__1107] ^ p82_literal_2043914[p82_res7__1109] ^ p82_literal_2043912[p82_res7__1111] ^ p82_literal_2043910[p83_res7__1113_comb] ^ p82_bit_slice_2059420;
  assign p83_res7__1117_comb = p82_array_index_2059437 ^ p82_array_index_2059465 ^ p82_array_index_2059491 ^ p82_array_index_2059651 ^ p82_array_index_2059673 ^ p82_array_index_2059693 ^ p82_res7__1099 ^ p82_literal_2043923[p82_res7__1101] ^ p82_res7__1103 ^ p82_literal_2043920[p82_res7__1105] ^ p82_literal_2043918[p82_res7__1107] ^ p82_literal_2043916[p82_res7__1109] ^ p82_literal_2043914[p82_res7__1111] ^ p82_literal_2043912[p83_res7__1113_comb] ^ p82_literal_2043910[p83_res7__1115_comb] ^ p82_bit_slice_2059421;
  assign p83_res7__1119_comb = p82_array_index_2059452 ^ p82_array_index_2059479 ^ p82_array_index_2059504 ^ p82_array_index_2059663 ^ p82_array_index_2059684 ^ p82_array_index_2059703 ^ p82_res7__1101 ^ p82_literal_2043923[p82_res7__1103] ^ p82_res7__1105 ^ p82_literal_2043920[p82_res7__1107] ^ p82_literal_2043918[p82_res7__1109] ^ p82_literal_2043916[p82_res7__1111] ^ p82_literal_2043914[p83_res7__1113_comb] ^ p82_literal_2043912[p83_res7__1115_comb] ^ p82_literal_2043910[p83_res7__1117_comb] ^ p82_bit_slice_2059422;
  assign p83_permut__34_comb = {p82_array_index_2059718, p82_array_index_2059719, p82_array_index_2059720, p82_literal_2058836[p82_res7__1095], p82_literal_2058836[p82_res7__1097], p82_literal_2058836[p82_res7__1099], p82_literal_2058836[p82_res7__1101], p82_literal_2058836[p82_res7__1103], p82_literal_2058836[p82_res7__1105], p82_literal_2058836[p82_res7__1107], p82_literal_2058836[p82_res7__1109], p82_literal_2058836[p82_res7__1111], p82_literal_2058836[p83_res7__1113_comb], p82_literal_2058836[p83_res7__1115_comb], p82_literal_2058836[p83_res7__1117_comb], p82_literal_2058836[p83_res7__1119_comb]};
  assign p83_xor_2059883_comb = p82_k6 ^ p83_permut__34_comb;
  assign p83_bit_slice_2059885_comb = p83_xor_2059883_comb[111:104];
  assign p83_bit_slice_2059886_comb = p83_xor_2059883_comb[103:96];
  assign p83_bit_slice_2059887_comb = p83_xor_2059883_comb[95:88];
  assign p83_bit_slice_2059888_comb = p83_xor_2059883_comb[87:80];
  assign p83_bit_slice_2059889_comb = p83_xor_2059883_comb[79:72];
  assign p83_bit_slice_2059890_comb = p83_xor_2059883_comb[63:56];
  assign p83_bit_slice_2059891_comb = p83_xor_2059883_comb[47:40];
  assign p83_bit_slice_2059892_comb = p83_xor_2059883_comb[39:32];
  assign p83_bit_slice_2059893_comb = p83_xor_2059883_comb[31:24];
  assign p83_bit_slice_2059894_comb = p83_xor_2059883_comb[23:16];
  assign p83_bit_slice_2059895_comb = p83_xor_2059883_comb[15:8];
  assign p83_bit_slice_2059896_comb = p83_xor_2059883_comb[7:0];
  assign p83_bit_slice_2059903_comb = p83_xor_2059883_comb[71:64];
  assign p83_bit_slice_2059905_comb = p83_xor_2059883_comb[55:48];
  assign p83_array_index_2059906_comb = p82_literal_2043920[p83_bit_slice_2059891_comb];
  assign p83_array_index_2059907_comb = p82_literal_2043918[p83_bit_slice_2059892_comb];
  assign p83_array_index_2059908_comb = p82_literal_2043916[p83_bit_slice_2059893_comb];
  assign p83_array_index_2059909_comb = p82_literal_2043914[p83_bit_slice_2059894_comb];
  assign p83_array_index_2059910_comb = p82_literal_2043912[p83_bit_slice_2059895_comb];
  assign p83_array_index_2059911_comb = p82_literal_2043910[p83_bit_slice_2059896_comb];
  assign p83_res7__1121_comb = p82_literal_2043910[p83_xor_2059883_comb[119:112]] ^ p82_literal_2043912[p83_bit_slice_2059885_comb] ^ p82_literal_2043914[p83_bit_slice_2059886_comb] ^ p82_literal_2043916[p83_bit_slice_2059887_comb] ^ p82_literal_2043918[p83_bit_slice_2059888_comb] ^ p82_literal_2043920[p83_bit_slice_2059889_comb] ^ p83_bit_slice_2059903_comb ^ p82_literal_2043923[p83_bit_slice_2059890_comb] ^ p83_bit_slice_2059905_comb ^ p83_array_index_2059906_comb ^ p83_array_index_2059907_comb ^ p83_array_index_2059908_comb ^ p83_array_index_2059909_comb ^ p83_array_index_2059910_comb ^ p83_array_index_2059911_comb ^ p83_xor_2059883_comb[127:120];
  assign p83_array_index_2059921_comb = p82_literal_2043920[p83_bit_slice_2059892_comb];
  assign p83_array_index_2059922_comb = p82_literal_2043918[p83_bit_slice_2059893_comb];
  assign p83_array_index_2059923_comb = p82_literal_2043916[p83_bit_slice_2059894_comb];
  assign p83_array_index_2059924_comb = p82_literal_2043914[p83_bit_slice_2059895_comb];
  assign p83_array_index_2059925_comb = p82_literal_2043912[p83_bit_slice_2059896_comb];
  assign p83_array_index_2059926_comb = p82_literal_2043910[p83_res7__1121_comb];
  assign p83_res7__1123_comb = p82_literal_2043910[p83_bit_slice_2059885_comb] ^ p82_literal_2043912[p83_bit_slice_2059886_comb] ^ p82_literal_2043914[p83_bit_slice_2059887_comb] ^ p82_literal_2043916[p83_bit_slice_2059888_comb] ^ p82_literal_2043918[p83_bit_slice_2059889_comb] ^ p82_literal_2043920[p83_bit_slice_2059903_comb] ^ p83_bit_slice_2059890_comb ^ p82_literal_2043923[p83_bit_slice_2059905_comb] ^ p83_bit_slice_2059891_comb ^ p83_array_index_2059921_comb ^ p83_array_index_2059922_comb ^ p83_array_index_2059923_comb ^ p83_array_index_2059924_comb ^ p83_array_index_2059925_comb ^ p83_array_index_2059926_comb ^ p83_xor_2059883_comb[119:112];
  assign p83_array_index_2059928_comb = p82_literal_2043910[p83_bit_slice_2059886_comb];
  assign p83_array_index_2059929_comb = p82_literal_2043912[p83_bit_slice_2059887_comb];
  assign p83_array_index_2059930_comb = p82_literal_2043914[p83_bit_slice_2059888_comb];
  assign p83_array_index_2059931_comb = p82_literal_2043916[p83_bit_slice_2059889_comb];
  assign p83_array_index_2059932_comb = p82_literal_2043918[p83_bit_slice_2059903_comb];
  assign p83_array_index_2059933_comb = p82_literal_2043920[p83_bit_slice_2059890_comb];
  assign p83_array_index_2059934_comb = p82_literal_2043923[p83_bit_slice_2059891_comb];
  assign p83_array_index_2059935_comb = p82_literal_2043920[p83_bit_slice_2059893_comb];
  assign p83_array_index_2059936_comb = p82_literal_2043918[p83_bit_slice_2059894_comb];
  assign p83_array_index_2059937_comb = p82_literal_2043916[p83_bit_slice_2059895_comb];
  assign p83_array_index_2059938_comb = p82_literal_2043914[p83_bit_slice_2059896_comb];
  assign p83_array_index_2059939_comb = p82_literal_2043912[p83_res7__1121_comb];
  assign p83_array_index_2059940_comb = p82_literal_2043910[p83_res7__1123_comb];

  // Registers for pipe stage 83:
  reg [127:0] p83_bit_slice_2043893;
  reg [127:0] p83_bit_slice_2044018;
  reg [127:0] p83_k3;
  reg [127:0] p83_k2;
  reg [127:0] p83_k5;
  reg [127:0] p83_k4;
  reg [7:0] p83_bit_slice_2059885;
  reg [7:0] p83_bit_slice_2059886;
  reg [7:0] p83_bit_slice_2059887;
  reg [7:0] p83_bit_slice_2059888;
  reg [7:0] p83_bit_slice_2059889;
  reg [7:0] p83_bit_slice_2059890;
  reg [7:0] p83_bit_slice_2059891;
  reg [7:0] p83_bit_slice_2059892;
  reg [7:0] p83_bit_slice_2059893;
  reg [7:0] p83_bit_slice_2059894;
  reg [7:0] p83_bit_slice_2059895;
  reg [7:0] p83_bit_slice_2059896;
  reg [7:0] p83_bit_slice_2059903;
  reg [7:0] p83_bit_slice_2059905;
  reg [7:0] p83_array_index_2059906;
  reg [7:0] p83_array_index_2059907;
  reg [7:0] p83_array_index_2059908;
  reg [7:0] p83_array_index_2059909;
  reg [7:0] p83_array_index_2059910;
  reg [7:0] p83_array_index_2059911;
  reg [7:0] p83_res7__1121;
  reg [7:0] p83_array_index_2059921;
  reg [7:0] p83_array_index_2059922;
  reg [7:0] p83_array_index_2059923;
  reg [7:0] p83_array_index_2059924;
  reg [7:0] p83_array_index_2059925;
  reg [7:0] p83_array_index_2059926;
  reg [7:0] p83_res7__1123;
  reg [7:0] p83_array_index_2059928;
  reg [7:0] p83_array_index_2059929;
  reg [7:0] p83_array_index_2059930;
  reg [7:0] p83_array_index_2059931;
  reg [7:0] p83_array_index_2059932;
  reg [7:0] p83_array_index_2059933;
  reg [7:0] p83_array_index_2059934;
  reg [7:0] p83_array_index_2059935;
  reg [7:0] p83_array_index_2059936;
  reg [7:0] p83_array_index_2059937;
  reg [7:0] p83_array_index_2059938;
  reg [7:0] p83_array_index_2059939;
  reg [7:0] p83_array_index_2059940;
  reg [7:0] p84_literal_2043910[256];
  reg [7:0] p84_literal_2043912[256];
  reg [7:0] p84_literal_2043914[256];
  reg [7:0] p84_literal_2043916[256];
  reg [7:0] p84_literal_2043918[256];
  reg [7:0] p84_literal_2043920[256];
  reg [7:0] p84_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p83_bit_slice_2043893 <= p82_bit_slice_2043893;
    p83_bit_slice_2044018 <= p82_bit_slice_2044018;
    p83_k3 <= p82_k3;
    p83_k2 <= p82_k2;
    p83_k5 <= p82_k5;
    p83_k4 <= p82_k4;
    p83_bit_slice_2059885 <= p83_bit_slice_2059885_comb;
    p83_bit_slice_2059886 <= p83_bit_slice_2059886_comb;
    p83_bit_slice_2059887 <= p83_bit_slice_2059887_comb;
    p83_bit_slice_2059888 <= p83_bit_slice_2059888_comb;
    p83_bit_slice_2059889 <= p83_bit_slice_2059889_comb;
    p83_bit_slice_2059890 <= p83_bit_slice_2059890_comb;
    p83_bit_slice_2059891 <= p83_bit_slice_2059891_comb;
    p83_bit_slice_2059892 <= p83_bit_slice_2059892_comb;
    p83_bit_slice_2059893 <= p83_bit_slice_2059893_comb;
    p83_bit_slice_2059894 <= p83_bit_slice_2059894_comb;
    p83_bit_slice_2059895 <= p83_bit_slice_2059895_comb;
    p83_bit_slice_2059896 <= p83_bit_slice_2059896_comb;
    p83_bit_slice_2059903 <= p83_bit_slice_2059903_comb;
    p83_bit_slice_2059905 <= p83_bit_slice_2059905_comb;
    p83_array_index_2059906 <= p83_array_index_2059906_comb;
    p83_array_index_2059907 <= p83_array_index_2059907_comb;
    p83_array_index_2059908 <= p83_array_index_2059908_comb;
    p83_array_index_2059909 <= p83_array_index_2059909_comb;
    p83_array_index_2059910 <= p83_array_index_2059910_comb;
    p83_array_index_2059911 <= p83_array_index_2059911_comb;
    p83_res7__1121 <= p83_res7__1121_comb;
    p83_array_index_2059921 <= p83_array_index_2059921_comb;
    p83_array_index_2059922 <= p83_array_index_2059922_comb;
    p83_array_index_2059923 <= p83_array_index_2059923_comb;
    p83_array_index_2059924 <= p83_array_index_2059924_comb;
    p83_array_index_2059925 <= p83_array_index_2059925_comb;
    p83_array_index_2059926 <= p83_array_index_2059926_comb;
    p83_res7__1123 <= p83_res7__1123_comb;
    p83_array_index_2059928 <= p83_array_index_2059928_comb;
    p83_array_index_2059929 <= p83_array_index_2059929_comb;
    p83_array_index_2059930 <= p83_array_index_2059930_comb;
    p83_array_index_2059931 <= p83_array_index_2059931_comb;
    p83_array_index_2059932 <= p83_array_index_2059932_comb;
    p83_array_index_2059933 <= p83_array_index_2059933_comb;
    p83_array_index_2059934 <= p83_array_index_2059934_comb;
    p83_array_index_2059935 <= p83_array_index_2059935_comb;
    p83_array_index_2059936 <= p83_array_index_2059936_comb;
    p83_array_index_2059937 <= p83_array_index_2059937_comb;
    p83_array_index_2059938 <= p83_array_index_2059938_comb;
    p83_array_index_2059939 <= p83_array_index_2059939_comb;
    p83_array_index_2059940 <= p83_array_index_2059940_comb;
    p84_literal_2043910 <= p83_literal_2043910;
    p84_literal_2043912 <= p83_literal_2043912;
    p84_literal_2043914 <= p83_literal_2043914;
    p84_literal_2043916 <= p83_literal_2043916;
    p84_literal_2043918 <= p83_literal_2043918;
    p84_literal_2043920 <= p83_literal_2043920;
    p84_literal_2043923 <= p83_literal_2043923;
  end

  // ===== Pipe stage 84:
  wire [7:0] p84_res7__1125_comb;
  wire [7:0] p84_array_index_2060059_comb;
  wire [7:0] p84_array_index_2060060_comb;
  wire [7:0] p84_array_index_2060061_comb;
  wire [7:0] p84_array_index_2060062_comb;
  wire [7:0] p84_array_index_2060063_comb;
  wire [7:0] p84_res7__1127_comb;
  wire [7:0] p84_array_index_2060072_comb;
  wire [7:0] p84_array_index_2060073_comb;
  wire [7:0] p84_array_index_2060074_comb;
  wire [7:0] p84_array_index_2060075_comb;
  wire [7:0] p84_res7__1129_comb;
  wire [7:0] p84_array_index_2060085_comb;
  wire [7:0] p84_array_index_2060086_comb;
  wire [7:0] p84_array_index_2060087_comb;
  wire [7:0] p84_array_index_2060088_comb;
  wire [7:0] p84_res7__1131_comb;
  wire [7:0] p84_array_index_2060097_comb;
  wire [7:0] p84_array_index_2060098_comb;
  wire [7:0] p84_array_index_2060099_comb;
  wire [7:0] p84_res7__1133_comb;
  wire [7:0] p84_array_index_2060109_comb;
  wire [7:0] p84_array_index_2060110_comb;
  wire [7:0] p84_array_index_2060111_comb;
  wire [7:0] p84_res7__1135_comb;
  wire [7:0] p84_array_index_2060120_comb;
  wire [7:0] p84_array_index_2060121_comb;
  wire [7:0] p84_res7__1137_comb;
  wire [7:0] p84_array_index_2060127_comb;
  wire [7:0] p84_array_index_2060128_comb;
  wire [7:0] p84_array_index_2060129_comb;
  wire [7:0] p84_array_index_2060130_comb;
  wire [7:0] p84_array_index_2060131_comb;
  wire [7:0] p84_array_index_2060132_comb;
  wire [7:0] p84_array_index_2060133_comb;
  wire [7:0] p84_array_index_2060134_comb;
  wire [7:0] p84_array_index_2060135_comb;
  wire [7:0] p84_array_index_2060136_comb;
  assign p84_res7__1125_comb = p83_array_index_2059928 ^ p83_array_index_2059929 ^ p83_array_index_2059930 ^ p83_array_index_2059931 ^ p83_array_index_2059932 ^ p83_array_index_2059933 ^ p83_bit_slice_2059905 ^ p83_array_index_2059934 ^ p83_bit_slice_2059892 ^ p83_array_index_2059935 ^ p83_array_index_2059936 ^ p83_array_index_2059937 ^ p83_array_index_2059938 ^ p83_array_index_2059939 ^ p83_array_index_2059940 ^ p83_bit_slice_2059885;
  assign p84_array_index_2060059_comb = p83_literal_2043920[p83_bit_slice_2059894];
  assign p84_array_index_2060060_comb = p83_literal_2043918[p83_bit_slice_2059895];
  assign p84_array_index_2060061_comb = p83_literal_2043916[p83_bit_slice_2059896];
  assign p84_array_index_2060062_comb = p83_literal_2043914[p83_res7__1121];
  assign p84_array_index_2060063_comb = p83_literal_2043912[p83_res7__1123];
  assign p84_res7__1127_comb = p83_literal_2043910[p83_bit_slice_2059887] ^ p83_literal_2043912[p83_bit_slice_2059888] ^ p83_literal_2043914[p83_bit_slice_2059889] ^ p83_literal_2043916[p83_bit_slice_2059903] ^ p83_literal_2043918[p83_bit_slice_2059890] ^ p83_literal_2043920[p83_bit_slice_2059905] ^ p83_bit_slice_2059891 ^ p83_literal_2043923[p83_bit_slice_2059892] ^ p83_bit_slice_2059893 ^ p84_array_index_2060059_comb ^ p84_array_index_2060060_comb ^ p84_array_index_2060061_comb ^ p84_array_index_2060062_comb ^ p84_array_index_2060063_comb ^ p83_literal_2043910[p84_res7__1125_comb] ^ p83_bit_slice_2059886;
  assign p84_array_index_2060072_comb = p83_literal_2043920[p83_bit_slice_2059895];
  assign p84_array_index_2060073_comb = p83_literal_2043918[p83_bit_slice_2059896];
  assign p84_array_index_2060074_comb = p83_literal_2043916[p83_res7__1121];
  assign p84_array_index_2060075_comb = p83_literal_2043914[p83_res7__1123];
  assign p84_res7__1129_comb = p83_literal_2043910[p83_bit_slice_2059888] ^ p83_literal_2043912[p83_bit_slice_2059889] ^ p83_literal_2043914[p83_bit_slice_2059903] ^ p83_literal_2043916[p83_bit_slice_2059890] ^ p83_literal_2043918[p83_bit_slice_2059905] ^ p83_array_index_2059906 ^ p83_bit_slice_2059892 ^ p83_literal_2043923[p83_bit_slice_2059893] ^ p83_bit_slice_2059894 ^ p84_array_index_2060072_comb ^ p84_array_index_2060073_comb ^ p84_array_index_2060074_comb ^ p84_array_index_2060075_comb ^ p83_literal_2043912[p84_res7__1125_comb] ^ p83_literal_2043910[p84_res7__1127_comb] ^ p83_bit_slice_2059887;
  assign p84_array_index_2060085_comb = p83_literal_2043920[p83_bit_slice_2059896];
  assign p84_array_index_2060086_comb = p83_literal_2043918[p83_res7__1121];
  assign p84_array_index_2060087_comb = p83_literal_2043916[p83_res7__1123];
  assign p84_array_index_2060088_comb = p83_literal_2043914[p84_res7__1125_comb];
  assign p84_res7__1131_comb = p83_literal_2043910[p83_bit_slice_2059889] ^ p83_literal_2043912[p83_bit_slice_2059903] ^ p83_literal_2043914[p83_bit_slice_2059890] ^ p83_literal_2043916[p83_bit_slice_2059905] ^ p83_literal_2043918[p83_bit_slice_2059891] ^ p83_array_index_2059921 ^ p83_bit_slice_2059893 ^ p83_literal_2043923[p83_bit_slice_2059894] ^ p83_bit_slice_2059895 ^ p84_array_index_2060085_comb ^ p84_array_index_2060086_comb ^ p84_array_index_2060087_comb ^ p84_array_index_2060088_comb ^ p83_literal_2043912[p84_res7__1127_comb] ^ p83_literal_2043910[p84_res7__1129_comb] ^ p83_bit_slice_2059888;
  assign p84_array_index_2060097_comb = p83_literal_2043920[p83_res7__1121];
  assign p84_array_index_2060098_comb = p83_literal_2043918[p83_res7__1123];
  assign p84_array_index_2060099_comb = p83_literal_2043916[p84_res7__1125_comb];
  assign p84_res7__1133_comb = p83_literal_2043910[p83_bit_slice_2059903] ^ p83_literal_2043912[p83_bit_slice_2059890] ^ p83_literal_2043914[p83_bit_slice_2059905] ^ p83_literal_2043916[p83_bit_slice_2059891] ^ p83_array_index_2059907 ^ p83_array_index_2059935 ^ p83_bit_slice_2059894 ^ p83_literal_2043923[p83_bit_slice_2059895] ^ p83_bit_slice_2059896 ^ p84_array_index_2060097_comb ^ p84_array_index_2060098_comb ^ p84_array_index_2060099_comb ^ p83_literal_2043914[p84_res7__1127_comb] ^ p83_literal_2043912[p84_res7__1129_comb] ^ p83_literal_2043910[p84_res7__1131_comb] ^ p83_bit_slice_2059889;
  assign p84_array_index_2060109_comb = p83_literal_2043920[p83_res7__1123];
  assign p84_array_index_2060110_comb = p83_literal_2043918[p84_res7__1125_comb];
  assign p84_array_index_2060111_comb = p83_literal_2043916[p84_res7__1127_comb];
  assign p84_res7__1135_comb = p83_literal_2043910[p83_bit_slice_2059890] ^ p83_literal_2043912[p83_bit_slice_2059905] ^ p83_literal_2043914[p83_bit_slice_2059891] ^ p83_literal_2043916[p83_bit_slice_2059892] ^ p83_array_index_2059922 ^ p84_array_index_2060059_comb ^ p83_bit_slice_2059895 ^ p83_literal_2043923[p83_bit_slice_2059896] ^ p83_res7__1121 ^ p84_array_index_2060109_comb ^ p84_array_index_2060110_comb ^ p84_array_index_2060111_comb ^ p83_literal_2043914[p84_res7__1129_comb] ^ p83_literal_2043912[p84_res7__1131_comb] ^ p83_literal_2043910[p84_res7__1133_comb] ^ p83_bit_slice_2059903;
  assign p84_array_index_2060120_comb = p83_literal_2043920[p84_res7__1125_comb];
  assign p84_array_index_2060121_comb = p83_literal_2043918[p84_res7__1127_comb];
  assign p84_res7__1137_comb = p83_literal_2043910[p83_bit_slice_2059905] ^ p83_literal_2043912[p83_bit_slice_2059891] ^ p83_literal_2043914[p83_bit_slice_2059892] ^ p83_array_index_2059908 ^ p83_array_index_2059936 ^ p84_array_index_2060072_comb ^ p83_bit_slice_2059896 ^ p83_literal_2043923[p83_res7__1121] ^ p83_res7__1123 ^ p84_array_index_2060120_comb ^ p84_array_index_2060121_comb ^ p83_literal_2043916[p84_res7__1129_comb] ^ p83_literal_2043914[p84_res7__1131_comb] ^ p83_literal_2043912[p84_res7__1133_comb] ^ p83_literal_2043910[p84_res7__1135_comb] ^ p83_bit_slice_2059890;
  assign p84_array_index_2060127_comb = p83_literal_2043910[p83_bit_slice_2059891];
  assign p84_array_index_2060128_comb = p83_literal_2043912[p83_bit_slice_2059892];
  assign p84_array_index_2060129_comb = p83_literal_2043914[p83_bit_slice_2059893];
  assign p84_array_index_2060130_comb = p83_literal_2043923[p83_res7__1123];
  assign p84_array_index_2060131_comb = p83_literal_2043920[p84_res7__1127_comb];
  assign p84_array_index_2060132_comb = p83_literal_2043918[p84_res7__1129_comb];
  assign p84_array_index_2060133_comb = p83_literal_2043916[p84_res7__1131_comb];
  assign p84_array_index_2060134_comb = p83_literal_2043914[p84_res7__1133_comb];
  assign p84_array_index_2060135_comb = p83_literal_2043912[p84_res7__1135_comb];
  assign p84_array_index_2060136_comb = p83_literal_2043910[p84_res7__1137_comb];

  // Registers for pipe stage 84:
  reg [127:0] p84_bit_slice_2043893;
  reg [127:0] p84_bit_slice_2044018;
  reg [127:0] p84_k3;
  reg [127:0] p84_k2;
  reg [127:0] p84_k5;
  reg [127:0] p84_k4;
  reg [7:0] p84_bit_slice_2059891;
  reg [7:0] p84_bit_slice_2059892;
  reg [7:0] p84_bit_slice_2059893;
  reg [7:0] p84_bit_slice_2059894;
  reg [7:0] p84_bit_slice_2059895;
  reg [7:0] p84_bit_slice_2059896;
  reg [7:0] p84_bit_slice_2059905;
  reg [7:0] p84_array_index_2059909;
  reg [7:0] p84_array_index_2059910;
  reg [7:0] p84_array_index_2059911;
  reg [7:0] p84_res7__1121;
  reg [7:0] p84_array_index_2059923;
  reg [7:0] p84_array_index_2059924;
  reg [7:0] p84_array_index_2059925;
  reg [7:0] p84_array_index_2059926;
  reg [7:0] p84_res7__1123;
  reg [7:0] p84_array_index_2059937;
  reg [7:0] p84_array_index_2059938;
  reg [7:0] p84_array_index_2059939;
  reg [7:0] p84_res7__1125;
  reg [7:0] p84_array_index_2060060;
  reg [7:0] p84_array_index_2060061;
  reg [7:0] p84_array_index_2060062;
  reg [7:0] p84_array_index_2060063;
  reg [7:0] p84_res7__1127;
  reg [7:0] p84_array_index_2060073;
  reg [7:0] p84_array_index_2060074;
  reg [7:0] p84_array_index_2060075;
  reg [7:0] p84_res7__1129;
  reg [7:0] p84_array_index_2060085;
  reg [7:0] p84_array_index_2060086;
  reg [7:0] p84_array_index_2060087;
  reg [7:0] p84_array_index_2060088;
  reg [7:0] p84_res7__1131;
  reg [7:0] p84_array_index_2060097;
  reg [7:0] p84_array_index_2060098;
  reg [7:0] p84_array_index_2060099;
  reg [7:0] p84_res7__1133;
  reg [7:0] p84_array_index_2060109;
  reg [7:0] p84_array_index_2060110;
  reg [7:0] p84_array_index_2060111;
  reg [7:0] p84_res7__1135;
  reg [7:0] p84_array_index_2060120;
  reg [7:0] p84_array_index_2060121;
  reg [7:0] p84_res7__1137;
  reg [7:0] p84_array_index_2060127;
  reg [7:0] p84_array_index_2060128;
  reg [7:0] p84_array_index_2060129;
  reg [7:0] p84_array_index_2060130;
  reg [7:0] p84_array_index_2060131;
  reg [7:0] p84_array_index_2060132;
  reg [7:0] p84_array_index_2060133;
  reg [7:0] p84_array_index_2060134;
  reg [7:0] p84_array_index_2060135;
  reg [7:0] p84_array_index_2060136;
  reg [7:0] p85_literal_2043910[256];
  reg [7:0] p85_literal_2043912[256];
  reg [7:0] p85_literal_2043914[256];
  reg [7:0] p85_literal_2043916[256];
  reg [7:0] p85_literal_2043918[256];
  reg [7:0] p85_literal_2043920[256];
  reg [7:0] p85_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p84_bit_slice_2043893 <= p83_bit_slice_2043893;
    p84_bit_slice_2044018 <= p83_bit_slice_2044018;
    p84_k3 <= p83_k3;
    p84_k2 <= p83_k2;
    p84_k5 <= p83_k5;
    p84_k4 <= p83_k4;
    p84_bit_slice_2059891 <= p83_bit_slice_2059891;
    p84_bit_slice_2059892 <= p83_bit_slice_2059892;
    p84_bit_slice_2059893 <= p83_bit_slice_2059893;
    p84_bit_slice_2059894 <= p83_bit_slice_2059894;
    p84_bit_slice_2059895 <= p83_bit_slice_2059895;
    p84_bit_slice_2059896 <= p83_bit_slice_2059896;
    p84_bit_slice_2059905 <= p83_bit_slice_2059905;
    p84_array_index_2059909 <= p83_array_index_2059909;
    p84_array_index_2059910 <= p83_array_index_2059910;
    p84_array_index_2059911 <= p83_array_index_2059911;
    p84_res7__1121 <= p83_res7__1121;
    p84_array_index_2059923 <= p83_array_index_2059923;
    p84_array_index_2059924 <= p83_array_index_2059924;
    p84_array_index_2059925 <= p83_array_index_2059925;
    p84_array_index_2059926 <= p83_array_index_2059926;
    p84_res7__1123 <= p83_res7__1123;
    p84_array_index_2059937 <= p83_array_index_2059937;
    p84_array_index_2059938 <= p83_array_index_2059938;
    p84_array_index_2059939 <= p83_array_index_2059939;
    p84_res7__1125 <= p84_res7__1125_comb;
    p84_array_index_2060060 <= p84_array_index_2060060_comb;
    p84_array_index_2060061 <= p84_array_index_2060061_comb;
    p84_array_index_2060062 <= p84_array_index_2060062_comb;
    p84_array_index_2060063 <= p84_array_index_2060063_comb;
    p84_res7__1127 <= p84_res7__1127_comb;
    p84_array_index_2060073 <= p84_array_index_2060073_comb;
    p84_array_index_2060074 <= p84_array_index_2060074_comb;
    p84_array_index_2060075 <= p84_array_index_2060075_comb;
    p84_res7__1129 <= p84_res7__1129_comb;
    p84_array_index_2060085 <= p84_array_index_2060085_comb;
    p84_array_index_2060086 <= p84_array_index_2060086_comb;
    p84_array_index_2060087 <= p84_array_index_2060087_comb;
    p84_array_index_2060088 <= p84_array_index_2060088_comb;
    p84_res7__1131 <= p84_res7__1131_comb;
    p84_array_index_2060097 <= p84_array_index_2060097_comb;
    p84_array_index_2060098 <= p84_array_index_2060098_comb;
    p84_array_index_2060099 <= p84_array_index_2060099_comb;
    p84_res7__1133 <= p84_res7__1133_comb;
    p84_array_index_2060109 <= p84_array_index_2060109_comb;
    p84_array_index_2060110 <= p84_array_index_2060110_comb;
    p84_array_index_2060111 <= p84_array_index_2060111_comb;
    p84_res7__1135 <= p84_res7__1135_comb;
    p84_array_index_2060120 <= p84_array_index_2060120_comb;
    p84_array_index_2060121 <= p84_array_index_2060121_comb;
    p84_res7__1137 <= p84_res7__1137_comb;
    p84_array_index_2060127 <= p84_array_index_2060127_comb;
    p84_array_index_2060128 <= p84_array_index_2060128_comb;
    p84_array_index_2060129 <= p84_array_index_2060129_comb;
    p84_array_index_2060130 <= p84_array_index_2060130_comb;
    p84_array_index_2060131 <= p84_array_index_2060131_comb;
    p84_array_index_2060132 <= p84_array_index_2060132_comb;
    p84_array_index_2060133 <= p84_array_index_2060133_comb;
    p84_array_index_2060134 <= p84_array_index_2060134_comb;
    p84_array_index_2060135 <= p84_array_index_2060135_comb;
    p84_array_index_2060136 <= p84_array_index_2060136_comb;
    p85_literal_2043910 <= p84_literal_2043910;
    p85_literal_2043912 <= p84_literal_2043912;
    p85_literal_2043914 <= p84_literal_2043914;
    p85_literal_2043916 <= p84_literal_2043916;
    p85_literal_2043918 <= p84_literal_2043918;
    p85_literal_2043920 <= p84_literal_2043920;
    p85_literal_2043923 <= p84_literal_2043923;
  end

  // ===== Pipe stage 85:
  wire [7:0] p85_res7__1139_comb;
  wire [7:0] p85_array_index_2060279_comb;
  wire [7:0] p85_res7__1141_comb;
  wire [7:0] p85_array_index_2060289_comb;
  wire [7:0] p85_res7__1143_comb;
  wire [7:0] p85_res7__1145_comb;
  wire [7:0] p85_res7__1147_comb;
  wire [7:0] p85_res7__1149_comb;
  wire [7:0] p85_res7__1151_comb;
  wire [127:0] p85_permut__35_comb;
  assign p85_res7__1139_comb = p84_array_index_2060127 ^ p84_array_index_2060128 ^ p84_array_index_2060129 ^ p84_array_index_2059923 ^ p84_array_index_2060060 ^ p84_array_index_2060085 ^ p84_res7__1121 ^ p84_array_index_2060130 ^ p84_res7__1125 ^ p84_array_index_2060131 ^ p84_array_index_2060132 ^ p84_array_index_2060133 ^ p84_array_index_2060134 ^ p84_array_index_2060135 ^ p84_array_index_2060136 ^ p84_bit_slice_2059905;
  assign p85_array_index_2060279_comb = p84_literal_2043920[p84_res7__1129];
  assign p85_res7__1141_comb = p84_literal_2043910[p84_bit_slice_2059892] ^ p84_literal_2043912[p84_bit_slice_2059893] ^ p84_array_index_2059909 ^ p84_array_index_2059937 ^ p84_array_index_2060073 ^ p84_array_index_2060097 ^ p84_res7__1123 ^ p84_literal_2043923[p84_res7__1125] ^ p84_res7__1127 ^ p85_array_index_2060279_comb ^ p84_literal_2043918[p84_res7__1131] ^ p84_literal_2043916[p84_res7__1133] ^ p84_literal_2043914[p84_res7__1135] ^ p84_literal_2043912[p84_res7__1137] ^ p84_literal_2043910[p85_res7__1139_comb] ^ p84_bit_slice_2059891;
  assign p85_array_index_2060289_comb = p84_literal_2043920[p84_res7__1131];
  assign p85_res7__1143_comb = p84_literal_2043910[p84_bit_slice_2059893] ^ p84_literal_2043912[p84_bit_slice_2059894] ^ p84_array_index_2059924 ^ p84_array_index_2060061 ^ p84_array_index_2060086 ^ p84_array_index_2060109 ^ p84_res7__1125 ^ p84_literal_2043923[p84_res7__1127] ^ p84_res7__1129 ^ p85_array_index_2060289_comb ^ p84_literal_2043918[p84_res7__1133] ^ p84_literal_2043916[p84_res7__1135] ^ p84_literal_2043914[p84_res7__1137] ^ p84_literal_2043912[p85_res7__1139_comb] ^ p84_literal_2043910[p85_res7__1141_comb] ^ p84_bit_slice_2059892;
  assign p85_res7__1145_comb = p84_literal_2043910[p84_bit_slice_2059894] ^ p84_array_index_2059910 ^ p84_array_index_2059938 ^ p84_array_index_2060074 ^ p84_array_index_2060098 ^ p84_array_index_2060120 ^ p84_res7__1127 ^ p84_literal_2043923[p84_res7__1129] ^ p84_res7__1131 ^ p84_literal_2043920[p84_res7__1133] ^ p84_literal_2043918[p84_res7__1135] ^ p84_literal_2043916[p84_res7__1137] ^ p84_literal_2043914[p85_res7__1139_comb] ^ p84_literal_2043912[p85_res7__1141_comb] ^ p84_literal_2043910[p85_res7__1143_comb] ^ p84_bit_slice_2059893;
  assign p85_res7__1147_comb = p84_literal_2043910[p84_bit_slice_2059895] ^ p84_array_index_2059925 ^ p84_array_index_2060062 ^ p84_array_index_2060087 ^ p84_array_index_2060110 ^ p84_array_index_2060131 ^ p84_res7__1129 ^ p84_literal_2043923[p84_res7__1131] ^ p84_res7__1133 ^ p84_literal_2043920[p84_res7__1135] ^ p84_literal_2043918[p84_res7__1137] ^ p84_literal_2043916[p85_res7__1139_comb] ^ p84_literal_2043914[p85_res7__1141_comb] ^ p84_literal_2043912[p85_res7__1143_comb] ^ p84_literal_2043910[p85_res7__1145_comb] ^ p84_bit_slice_2059894;
  assign p85_res7__1149_comb = p84_array_index_2059911 ^ p84_array_index_2059939 ^ p84_array_index_2060075 ^ p84_array_index_2060099 ^ p84_array_index_2060121 ^ p85_array_index_2060279_comb ^ p84_res7__1131 ^ p84_literal_2043923[p84_res7__1133] ^ p84_res7__1135 ^ p84_literal_2043920[p84_res7__1137] ^ p84_literal_2043918[p85_res7__1139_comb] ^ p84_literal_2043916[p85_res7__1141_comb] ^ p84_literal_2043914[p85_res7__1143_comb] ^ p84_literal_2043912[p85_res7__1145_comb] ^ p84_literal_2043910[p85_res7__1147_comb] ^ p84_bit_slice_2059895;
  assign p85_res7__1151_comb = p84_array_index_2059926 ^ p84_array_index_2060063 ^ p84_array_index_2060088 ^ p84_array_index_2060111 ^ p84_array_index_2060132 ^ p85_array_index_2060289_comb ^ p84_res7__1133 ^ p84_literal_2043923[p84_res7__1135] ^ p84_res7__1137 ^ p84_literal_2043920[p85_res7__1139_comb] ^ p84_literal_2043918[p85_res7__1141_comb] ^ p84_literal_2043916[p85_res7__1143_comb] ^ p84_literal_2043914[p85_res7__1145_comb] ^ p84_literal_2043912[p85_res7__1147_comb] ^ p84_literal_2043910[p85_res7__1149_comb] ^ p84_bit_slice_2059896;
  assign p85_permut__35_comb = {p84_literal_2058836[p84_res7__1121], p84_literal_2058836[p84_res7__1123], p84_literal_2058836[p84_res7__1125], p84_literal_2058836[p84_res7__1127], p84_literal_2058836[p84_res7__1129], p84_literal_2058836[p84_res7__1131], p84_literal_2058836[p84_res7__1133], p84_literal_2058836[p84_res7__1135], p84_literal_2058836[p84_res7__1137], p84_literal_2058836[p85_res7__1139_comb], p84_literal_2058836[p85_res7__1141_comb], p84_literal_2058836[p85_res7__1143_comb], p84_literal_2058836[p85_res7__1145_comb], p84_literal_2058836[p85_res7__1147_comb], p84_literal_2058836[p85_res7__1149_comb], p84_literal_2058836[p85_res7__1151_comb]};

  // Registers for pipe stage 85:
  reg [127:0] p85_bit_slice_2043893;
  reg [127:0] p85_bit_slice_2044018;
  reg [127:0] p85_k3;
  reg [127:0] p85_k2;
  reg [127:0] p85_k5;
  reg [127:0] p85_k4;
  reg [127:0] p85_permut__35;
  reg [7:0] p86_literal_2043910[256];
  reg [7:0] p86_literal_2043912[256];
  reg [7:0] p86_literal_2043914[256];
  reg [7:0] p86_literal_2043916[256];
  reg [7:0] p86_literal_2043918[256];
  reg [7:0] p86_literal_2043920[256];
  reg [7:0] p86_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p85_bit_slice_2043893 <= p84_bit_slice_2043893;
    p85_bit_slice_2044018 <= p84_bit_slice_2044018;
    p85_k3 <= p84_k3;
    p85_k2 <= p84_k2;
    p85_k5 <= p84_k5;
    p85_k4 <= p84_k4;
    p85_permut__35 <= p85_permut__35_comb;
    p86_literal_2043910 <= p85_literal_2043910;
    p86_literal_2043912 <= p85_literal_2043912;
    p86_literal_2043914 <= p85_literal_2043914;
    p86_literal_2043916 <= p85_literal_2043916;
    p86_literal_2043918 <= p85_literal_2043918;
    p86_literal_2043920 <= p85_literal_2043920;
    p86_literal_2043923 <= p85_literal_2043923;
  end

  // ===== Pipe stage 86:
  wire [127:0] p86_xor_2060377_comb;
  wire [7:0] p86_bit_slice_2060383_comb;
  wire [7:0] p86_bit_slice_2060384_comb;
  wire [7:0] p86_bit_slice_2060385_comb;
  wire [7:0] p86_bit_slice_2060386_comb;
  wire [7:0] p86_bit_slice_2060387_comb;
  wire [7:0] p86_bit_slice_2060388_comb;
  wire [7:0] p86_bit_slice_2060389_comb;
  wire [7:0] p86_bit_slice_2060390_comb;
  wire [7:0] p86_bit_slice_2060397_comb;
  wire [7:0] p86_bit_slice_2060399_comb;
  wire [7:0] p86_array_index_2060400_comb;
  wire [7:0] p86_array_index_2060401_comb;
  wire [7:0] p86_array_index_2060402_comb;
  wire [7:0] p86_array_index_2060403_comb;
  wire [7:0] p86_array_index_2060404_comb;
  wire [7:0] p86_array_index_2060405_comb;
  wire [7:0] p86_res7__1153_comb;
  wire [7:0] p86_array_index_2060415_comb;
  wire [7:0] p86_array_index_2060416_comb;
  wire [7:0] p86_array_index_2060417_comb;
  wire [7:0] p86_array_index_2060418_comb;
  wire [7:0] p86_array_index_2060419_comb;
  wire [7:0] p86_array_index_2060420_comb;
  wire [7:0] p86_res7__1155_comb;
  wire [7:0] p86_array_index_2060429_comb;
  wire [7:0] p86_array_index_2060430_comb;
  wire [7:0] p86_array_index_2060431_comb;
  wire [7:0] p86_array_index_2060432_comb;
  wire [7:0] p86_array_index_2060433_comb;
  wire [7:0] p86_res7__1157_comb;
  wire [7:0] p86_array_index_2060443_comb;
  wire [7:0] p86_array_index_2060444_comb;
  wire [7:0] p86_array_index_2060445_comb;
  wire [7:0] p86_array_index_2060446_comb;
  wire [7:0] p86_array_index_2060447_comb;
  wire [7:0] p86_res7__1159_comb;
  wire [7:0] p86_array_index_2060456_comb;
  wire [7:0] p86_array_index_2060457_comb;
  wire [7:0] p86_array_index_2060458_comb;
  wire [7:0] p86_array_index_2060459_comb;
  wire [7:0] p86_res7__1161_comb;
  wire [7:0] p86_array_index_2060469_comb;
  wire [7:0] p86_array_index_2060470_comb;
  wire [7:0] p86_array_index_2060471_comb;
  wire [7:0] p86_array_index_2060472_comb;
  wire [7:0] p86_res7__1163_comb;
  wire [7:0] p86_array_index_2060476_comb;
  wire [7:0] p86_array_index_2060477_comb;
  wire [7:0] p86_array_index_2060478_comb;
  wire [7:0] p86_array_index_2060479_comb;
  wire [7:0] p86_array_index_2060480_comb;
  wire [7:0] p86_array_index_2060481_comb;
  wire [7:0] p86_array_index_2060482_comb;
  wire [7:0] p86_array_index_2060483_comb;
  wire [7:0] p86_array_index_2060484_comb;
  wire [7:0] p86_array_index_2060485_comb;
  wire [7:0] p86_array_index_2060486_comb;
  assign p86_xor_2060377_comb = p85_k5 ^ p85_permut__35;
  assign p86_bit_slice_2060383_comb = p86_xor_2060377_comb[79:72];
  assign p86_bit_slice_2060384_comb = p86_xor_2060377_comb[63:56];
  assign p86_bit_slice_2060385_comb = p86_xor_2060377_comb[47:40];
  assign p86_bit_slice_2060386_comb = p86_xor_2060377_comb[39:32];
  assign p86_bit_slice_2060387_comb = p86_xor_2060377_comb[31:24];
  assign p86_bit_slice_2060388_comb = p86_xor_2060377_comb[23:16];
  assign p86_bit_slice_2060389_comb = p86_xor_2060377_comb[15:8];
  assign p86_bit_slice_2060390_comb = p86_xor_2060377_comb[7:0];
  assign p86_bit_slice_2060397_comb = p86_xor_2060377_comb[71:64];
  assign p86_bit_slice_2060399_comb = p86_xor_2060377_comb[55:48];
  assign p86_array_index_2060400_comb = p85_literal_2043920[p86_bit_slice_2060385_comb];
  assign p86_array_index_2060401_comb = p85_literal_2043918[p86_bit_slice_2060386_comb];
  assign p86_array_index_2060402_comb = p85_literal_2043916[p86_bit_slice_2060387_comb];
  assign p86_array_index_2060403_comb = p85_literal_2043914[p86_bit_slice_2060388_comb];
  assign p86_array_index_2060404_comb = p85_literal_2043912[p86_bit_slice_2060389_comb];
  assign p86_array_index_2060405_comb = p85_literal_2043910[p86_bit_slice_2060390_comb];
  assign p86_res7__1153_comb = p85_literal_2043910[p86_xor_2060377_comb[119:112]] ^ p85_literal_2043912[p86_xor_2060377_comb[111:104]] ^ p85_literal_2043914[p86_xor_2060377_comb[103:96]] ^ p85_literal_2043916[p86_xor_2060377_comb[95:88]] ^ p85_literal_2043918[p86_xor_2060377_comb[87:80]] ^ p85_literal_2043920[p86_bit_slice_2060383_comb] ^ p86_bit_slice_2060397_comb ^ p85_literal_2043923[p86_bit_slice_2060384_comb] ^ p86_bit_slice_2060399_comb ^ p86_array_index_2060400_comb ^ p86_array_index_2060401_comb ^ p86_array_index_2060402_comb ^ p86_array_index_2060403_comb ^ p86_array_index_2060404_comb ^ p86_array_index_2060405_comb ^ p86_xor_2060377_comb[127:120];
  assign p86_array_index_2060415_comb = p85_literal_2043920[p86_bit_slice_2060386_comb];
  assign p86_array_index_2060416_comb = p85_literal_2043918[p86_bit_slice_2060387_comb];
  assign p86_array_index_2060417_comb = p85_literal_2043916[p86_bit_slice_2060388_comb];
  assign p86_array_index_2060418_comb = p85_literal_2043914[p86_bit_slice_2060389_comb];
  assign p86_array_index_2060419_comb = p85_literal_2043912[p86_bit_slice_2060390_comb];
  assign p86_array_index_2060420_comb = p85_literal_2043910[p86_res7__1153_comb];
  assign p86_res7__1155_comb = p85_literal_2043910[p86_xor_2060377_comb[111:104]] ^ p85_literal_2043912[p86_xor_2060377_comb[103:96]] ^ p85_literal_2043914[p86_xor_2060377_comb[95:88]] ^ p85_literal_2043916[p86_xor_2060377_comb[87:80]] ^ p85_literal_2043918[p86_bit_slice_2060383_comb] ^ p85_literal_2043920[p86_bit_slice_2060397_comb] ^ p86_bit_slice_2060384_comb ^ p85_literal_2043923[p86_bit_slice_2060399_comb] ^ p86_bit_slice_2060385_comb ^ p86_array_index_2060415_comb ^ p86_array_index_2060416_comb ^ p86_array_index_2060417_comb ^ p86_array_index_2060418_comb ^ p86_array_index_2060419_comb ^ p86_array_index_2060420_comb ^ p86_xor_2060377_comb[119:112];
  assign p86_array_index_2060429_comb = p85_literal_2043920[p86_bit_slice_2060387_comb];
  assign p86_array_index_2060430_comb = p85_literal_2043918[p86_bit_slice_2060388_comb];
  assign p86_array_index_2060431_comb = p85_literal_2043916[p86_bit_slice_2060389_comb];
  assign p86_array_index_2060432_comb = p85_literal_2043914[p86_bit_slice_2060390_comb];
  assign p86_array_index_2060433_comb = p85_literal_2043912[p86_res7__1153_comb];
  assign p86_res7__1157_comb = p85_literal_2043910[p86_xor_2060377_comb[103:96]] ^ p85_literal_2043912[p86_xor_2060377_comb[95:88]] ^ p85_literal_2043914[p86_xor_2060377_comb[87:80]] ^ p85_literal_2043916[p86_bit_slice_2060383_comb] ^ p85_literal_2043918[p86_bit_slice_2060397_comb] ^ p85_literal_2043920[p86_bit_slice_2060384_comb] ^ p86_bit_slice_2060399_comb ^ p85_literal_2043923[p86_bit_slice_2060385_comb] ^ p86_bit_slice_2060386_comb ^ p86_array_index_2060429_comb ^ p86_array_index_2060430_comb ^ p86_array_index_2060431_comb ^ p86_array_index_2060432_comb ^ p86_array_index_2060433_comb ^ p85_literal_2043910[p86_res7__1155_comb] ^ p86_xor_2060377_comb[111:104];
  assign p86_array_index_2060443_comb = p85_literal_2043920[p86_bit_slice_2060388_comb];
  assign p86_array_index_2060444_comb = p85_literal_2043918[p86_bit_slice_2060389_comb];
  assign p86_array_index_2060445_comb = p85_literal_2043916[p86_bit_slice_2060390_comb];
  assign p86_array_index_2060446_comb = p85_literal_2043914[p86_res7__1153_comb];
  assign p86_array_index_2060447_comb = p85_literal_2043912[p86_res7__1155_comb];
  assign p86_res7__1159_comb = p85_literal_2043910[p86_xor_2060377_comb[95:88]] ^ p85_literal_2043912[p86_xor_2060377_comb[87:80]] ^ p85_literal_2043914[p86_bit_slice_2060383_comb] ^ p85_literal_2043916[p86_bit_slice_2060397_comb] ^ p85_literal_2043918[p86_bit_slice_2060384_comb] ^ p85_literal_2043920[p86_bit_slice_2060399_comb] ^ p86_bit_slice_2060385_comb ^ p85_literal_2043923[p86_bit_slice_2060386_comb] ^ p86_bit_slice_2060387_comb ^ p86_array_index_2060443_comb ^ p86_array_index_2060444_comb ^ p86_array_index_2060445_comb ^ p86_array_index_2060446_comb ^ p86_array_index_2060447_comb ^ p85_literal_2043910[p86_res7__1157_comb] ^ p86_xor_2060377_comb[103:96];
  assign p86_array_index_2060456_comb = p85_literal_2043920[p86_bit_slice_2060389_comb];
  assign p86_array_index_2060457_comb = p85_literal_2043918[p86_bit_slice_2060390_comb];
  assign p86_array_index_2060458_comb = p85_literal_2043916[p86_res7__1153_comb];
  assign p86_array_index_2060459_comb = p85_literal_2043914[p86_res7__1155_comb];
  assign p86_res7__1161_comb = p85_literal_2043910[p86_xor_2060377_comb[87:80]] ^ p85_literal_2043912[p86_bit_slice_2060383_comb] ^ p85_literal_2043914[p86_bit_slice_2060397_comb] ^ p85_literal_2043916[p86_bit_slice_2060384_comb] ^ p85_literal_2043918[p86_bit_slice_2060399_comb] ^ p86_array_index_2060400_comb ^ p86_bit_slice_2060386_comb ^ p85_literal_2043923[p86_bit_slice_2060387_comb] ^ p86_bit_slice_2060388_comb ^ p86_array_index_2060456_comb ^ p86_array_index_2060457_comb ^ p86_array_index_2060458_comb ^ p86_array_index_2060459_comb ^ p85_literal_2043912[p86_res7__1157_comb] ^ p85_literal_2043910[p86_res7__1159_comb] ^ p86_xor_2060377_comb[95:88];
  assign p86_array_index_2060469_comb = p85_literal_2043920[p86_bit_slice_2060390_comb];
  assign p86_array_index_2060470_comb = p85_literal_2043918[p86_res7__1153_comb];
  assign p86_array_index_2060471_comb = p85_literal_2043916[p86_res7__1155_comb];
  assign p86_array_index_2060472_comb = p85_literal_2043914[p86_res7__1157_comb];
  assign p86_res7__1163_comb = p85_literal_2043910[p86_bit_slice_2060383_comb] ^ p85_literal_2043912[p86_bit_slice_2060397_comb] ^ p85_literal_2043914[p86_bit_slice_2060384_comb] ^ p85_literal_2043916[p86_bit_slice_2060399_comb] ^ p85_literal_2043918[p86_bit_slice_2060385_comb] ^ p86_array_index_2060415_comb ^ p86_bit_slice_2060387_comb ^ p85_literal_2043923[p86_bit_slice_2060388_comb] ^ p86_bit_slice_2060389_comb ^ p86_array_index_2060469_comb ^ p86_array_index_2060470_comb ^ p86_array_index_2060471_comb ^ p86_array_index_2060472_comb ^ p85_literal_2043912[p86_res7__1159_comb] ^ p85_literal_2043910[p86_res7__1161_comb] ^ p86_xor_2060377_comb[87:80];
  assign p86_array_index_2060476_comb = p85_literal_2043910[p86_bit_slice_2060397_comb];
  assign p86_array_index_2060477_comb = p85_literal_2043912[p86_bit_slice_2060384_comb];
  assign p86_array_index_2060478_comb = p85_literal_2043914[p86_bit_slice_2060399_comb];
  assign p86_array_index_2060479_comb = p85_literal_2043916[p86_bit_slice_2060385_comb];
  assign p86_array_index_2060480_comb = p85_literal_2043923[p86_bit_slice_2060389_comb];
  assign p86_array_index_2060481_comb = p85_literal_2043920[p86_res7__1153_comb];
  assign p86_array_index_2060482_comb = p85_literal_2043918[p86_res7__1155_comb];
  assign p86_array_index_2060483_comb = p85_literal_2043916[p86_res7__1157_comb];
  assign p86_array_index_2060484_comb = p85_literal_2043914[p86_res7__1159_comb];
  assign p86_array_index_2060485_comb = p85_literal_2043912[p86_res7__1161_comb];
  assign p86_array_index_2060486_comb = p85_literal_2043910[p86_res7__1163_comb];

  // Registers for pipe stage 86:
  reg [127:0] p86_bit_slice_2043893;
  reg [127:0] p86_bit_slice_2044018;
  reg [127:0] p86_k3;
  reg [127:0] p86_k2;
  reg [127:0] p86_k4;
  reg [7:0] p86_bit_slice_2060383;
  reg [7:0] p86_bit_slice_2060384;
  reg [7:0] p86_bit_slice_2060385;
  reg [7:0] p86_bit_slice_2060386;
  reg [7:0] p86_bit_slice_2060387;
  reg [7:0] p86_bit_slice_2060388;
  reg [7:0] p86_bit_slice_2060389;
  reg [7:0] p86_bit_slice_2060390;
  reg [7:0] p86_bit_slice_2060397;
  reg [7:0] p86_bit_slice_2060399;
  reg [7:0] p86_array_index_2060401;
  reg [7:0] p86_array_index_2060402;
  reg [7:0] p86_array_index_2060403;
  reg [7:0] p86_array_index_2060404;
  reg [7:0] p86_array_index_2060405;
  reg [7:0] p86_res7__1153;
  reg [7:0] p86_array_index_2060416;
  reg [7:0] p86_array_index_2060417;
  reg [7:0] p86_array_index_2060418;
  reg [7:0] p86_array_index_2060419;
  reg [7:0] p86_array_index_2060420;
  reg [7:0] p86_res7__1155;
  reg [7:0] p86_array_index_2060429;
  reg [7:0] p86_array_index_2060430;
  reg [7:0] p86_array_index_2060431;
  reg [7:0] p86_array_index_2060432;
  reg [7:0] p86_array_index_2060433;
  reg [7:0] p86_res7__1157;
  reg [7:0] p86_array_index_2060443;
  reg [7:0] p86_array_index_2060444;
  reg [7:0] p86_array_index_2060445;
  reg [7:0] p86_array_index_2060446;
  reg [7:0] p86_array_index_2060447;
  reg [7:0] p86_res7__1159;
  reg [7:0] p86_array_index_2060456;
  reg [7:0] p86_array_index_2060457;
  reg [7:0] p86_array_index_2060458;
  reg [7:0] p86_array_index_2060459;
  reg [7:0] p86_res7__1161;
  reg [7:0] p86_array_index_2060469;
  reg [7:0] p86_array_index_2060470;
  reg [7:0] p86_array_index_2060471;
  reg [7:0] p86_array_index_2060472;
  reg [7:0] p86_res7__1163;
  reg [7:0] p86_array_index_2060476;
  reg [7:0] p86_array_index_2060477;
  reg [7:0] p86_array_index_2060478;
  reg [7:0] p86_array_index_2060479;
  reg [7:0] p86_array_index_2060480;
  reg [7:0] p86_array_index_2060481;
  reg [7:0] p86_array_index_2060482;
  reg [7:0] p86_array_index_2060483;
  reg [7:0] p86_array_index_2060484;
  reg [7:0] p86_array_index_2060485;
  reg [7:0] p86_array_index_2060486;
  reg [7:0] p87_literal_2043910[256];
  reg [7:0] p87_literal_2043912[256];
  reg [7:0] p87_literal_2043914[256];
  reg [7:0] p87_literal_2043916[256];
  reg [7:0] p87_literal_2043918[256];
  reg [7:0] p87_literal_2043920[256];
  reg [7:0] p87_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p86_bit_slice_2043893 <= p85_bit_slice_2043893;
    p86_bit_slice_2044018 <= p85_bit_slice_2044018;
    p86_k3 <= p85_k3;
    p86_k2 <= p85_k2;
    p86_k4 <= p85_k4;
    p86_bit_slice_2060383 <= p86_bit_slice_2060383_comb;
    p86_bit_slice_2060384 <= p86_bit_slice_2060384_comb;
    p86_bit_slice_2060385 <= p86_bit_slice_2060385_comb;
    p86_bit_slice_2060386 <= p86_bit_slice_2060386_comb;
    p86_bit_slice_2060387 <= p86_bit_slice_2060387_comb;
    p86_bit_slice_2060388 <= p86_bit_slice_2060388_comb;
    p86_bit_slice_2060389 <= p86_bit_slice_2060389_comb;
    p86_bit_slice_2060390 <= p86_bit_slice_2060390_comb;
    p86_bit_slice_2060397 <= p86_bit_slice_2060397_comb;
    p86_bit_slice_2060399 <= p86_bit_slice_2060399_comb;
    p86_array_index_2060401 <= p86_array_index_2060401_comb;
    p86_array_index_2060402 <= p86_array_index_2060402_comb;
    p86_array_index_2060403 <= p86_array_index_2060403_comb;
    p86_array_index_2060404 <= p86_array_index_2060404_comb;
    p86_array_index_2060405 <= p86_array_index_2060405_comb;
    p86_res7__1153 <= p86_res7__1153_comb;
    p86_array_index_2060416 <= p86_array_index_2060416_comb;
    p86_array_index_2060417 <= p86_array_index_2060417_comb;
    p86_array_index_2060418 <= p86_array_index_2060418_comb;
    p86_array_index_2060419 <= p86_array_index_2060419_comb;
    p86_array_index_2060420 <= p86_array_index_2060420_comb;
    p86_res7__1155 <= p86_res7__1155_comb;
    p86_array_index_2060429 <= p86_array_index_2060429_comb;
    p86_array_index_2060430 <= p86_array_index_2060430_comb;
    p86_array_index_2060431 <= p86_array_index_2060431_comb;
    p86_array_index_2060432 <= p86_array_index_2060432_comb;
    p86_array_index_2060433 <= p86_array_index_2060433_comb;
    p86_res7__1157 <= p86_res7__1157_comb;
    p86_array_index_2060443 <= p86_array_index_2060443_comb;
    p86_array_index_2060444 <= p86_array_index_2060444_comb;
    p86_array_index_2060445 <= p86_array_index_2060445_comb;
    p86_array_index_2060446 <= p86_array_index_2060446_comb;
    p86_array_index_2060447 <= p86_array_index_2060447_comb;
    p86_res7__1159 <= p86_res7__1159_comb;
    p86_array_index_2060456 <= p86_array_index_2060456_comb;
    p86_array_index_2060457 <= p86_array_index_2060457_comb;
    p86_array_index_2060458 <= p86_array_index_2060458_comb;
    p86_array_index_2060459 <= p86_array_index_2060459_comb;
    p86_res7__1161 <= p86_res7__1161_comb;
    p86_array_index_2060469 <= p86_array_index_2060469_comb;
    p86_array_index_2060470 <= p86_array_index_2060470_comb;
    p86_array_index_2060471 <= p86_array_index_2060471_comb;
    p86_array_index_2060472 <= p86_array_index_2060472_comb;
    p86_res7__1163 <= p86_res7__1163_comb;
    p86_array_index_2060476 <= p86_array_index_2060476_comb;
    p86_array_index_2060477 <= p86_array_index_2060477_comb;
    p86_array_index_2060478 <= p86_array_index_2060478_comb;
    p86_array_index_2060479 <= p86_array_index_2060479_comb;
    p86_array_index_2060480 <= p86_array_index_2060480_comb;
    p86_array_index_2060481 <= p86_array_index_2060481_comb;
    p86_array_index_2060482 <= p86_array_index_2060482_comb;
    p86_array_index_2060483 <= p86_array_index_2060483_comb;
    p86_array_index_2060484 <= p86_array_index_2060484_comb;
    p86_array_index_2060485 <= p86_array_index_2060485_comb;
    p86_array_index_2060486 <= p86_array_index_2060486_comb;
    p87_literal_2043910 <= p86_literal_2043910;
    p87_literal_2043912 <= p86_literal_2043912;
    p87_literal_2043914 <= p86_literal_2043914;
    p87_literal_2043916 <= p86_literal_2043916;
    p87_literal_2043918 <= p86_literal_2043918;
    p87_literal_2043920 <= p86_literal_2043920;
    p87_literal_2043923 <= p86_literal_2043923;
  end

  // ===== Pipe stage 87:
  wire [7:0] p87_res7__1165_comb;
  wire [7:0] p87_array_index_2060629_comb;
  wire [7:0] p87_array_index_2060630_comb;
  wire [7:0] p87_array_index_2060631_comb;
  wire [7:0] p87_res7__1167_comb;
  wire [7:0] p87_array_index_2060640_comb;
  wire [7:0] p87_array_index_2060641_comb;
  wire [7:0] p87_res7__1169_comb;
  wire [7:0] p87_array_index_2060651_comb;
  wire [7:0] p87_array_index_2060652_comb;
  wire [7:0] p87_res7__1171_comb;
  wire [7:0] p87_array_index_2060661_comb;
  wire [7:0] p87_res7__1173_comb;
  wire [7:0] p87_array_index_2060671_comb;
  wire [7:0] p87_res7__1175_comb;
  wire [7:0] p87_res7__1177_comb;
  wire [7:0] p87_array_index_2060687_comb;
  wire [7:0] p87_array_index_2060688_comb;
  wire [7:0] p87_array_index_2060689_comb;
  wire [7:0] p87_array_index_2060690_comb;
  wire [7:0] p87_array_index_2060691_comb;
  wire [7:0] p87_array_index_2060692_comb;
  wire [7:0] p87_array_index_2060693_comb;
  wire [7:0] p87_array_index_2060694_comb;
  wire [7:0] p87_array_index_2060695_comb;
  wire [7:0] p87_array_index_2060696_comb;
  wire [7:0] p87_array_index_2060697_comb;
  wire [7:0] p87_array_index_2060698_comb;
  assign p87_res7__1165_comb = p86_array_index_2060476 ^ p86_array_index_2060477 ^ p86_array_index_2060478 ^ p86_array_index_2060479 ^ p86_array_index_2060401 ^ p86_array_index_2060429 ^ p86_bit_slice_2060388 ^ p86_array_index_2060480 ^ p86_bit_slice_2060390 ^ p86_array_index_2060481 ^ p86_array_index_2060482 ^ p86_array_index_2060483 ^ p86_array_index_2060484 ^ p86_array_index_2060485 ^ p86_array_index_2060486 ^ p86_bit_slice_2060383;
  assign p87_array_index_2060629_comb = p86_literal_2043920[p86_res7__1155];
  assign p87_array_index_2060630_comb = p86_literal_2043918[p86_res7__1157];
  assign p87_array_index_2060631_comb = p86_literal_2043916[p86_res7__1159];
  assign p87_res7__1167_comb = p86_literal_2043910[p86_bit_slice_2060384] ^ p86_literal_2043912[p86_bit_slice_2060399] ^ p86_literal_2043914[p86_bit_slice_2060385] ^ p86_literal_2043916[p86_bit_slice_2060386] ^ p86_array_index_2060416 ^ p86_array_index_2060443 ^ p86_bit_slice_2060389 ^ p86_literal_2043923[p86_bit_slice_2060390] ^ p86_res7__1153 ^ p87_array_index_2060629_comb ^ p87_array_index_2060630_comb ^ p87_array_index_2060631_comb ^ p86_literal_2043914[p86_res7__1161] ^ p86_literal_2043912[p86_res7__1163] ^ p86_literal_2043910[p87_res7__1165_comb] ^ p86_bit_slice_2060397;
  assign p87_array_index_2060640_comb = p86_literal_2043920[p86_res7__1157];
  assign p87_array_index_2060641_comb = p86_literal_2043918[p86_res7__1159];
  assign p87_res7__1169_comb = p86_literal_2043910[p86_bit_slice_2060399] ^ p86_literal_2043912[p86_bit_slice_2060385] ^ p86_literal_2043914[p86_bit_slice_2060386] ^ p86_array_index_2060402 ^ p86_array_index_2060430 ^ p86_array_index_2060456 ^ p86_bit_slice_2060390 ^ p86_literal_2043923[p86_res7__1153] ^ p86_res7__1155 ^ p87_array_index_2060640_comb ^ p87_array_index_2060641_comb ^ p86_literal_2043916[p86_res7__1161] ^ p86_literal_2043914[p86_res7__1163] ^ p86_literal_2043912[p87_res7__1165_comb] ^ p86_literal_2043910[p87_res7__1167_comb] ^ p86_bit_slice_2060384;
  assign p87_array_index_2060651_comb = p86_literal_2043920[p86_res7__1159];
  assign p87_array_index_2060652_comb = p86_literal_2043918[p86_res7__1161];
  assign p87_res7__1171_comb = p86_literal_2043910[p86_bit_slice_2060385] ^ p86_literal_2043912[p86_bit_slice_2060386] ^ p86_literal_2043914[p86_bit_slice_2060387] ^ p86_array_index_2060417 ^ p86_array_index_2060444 ^ p86_array_index_2060469 ^ p86_res7__1153 ^ p86_literal_2043923[p86_res7__1155] ^ p86_res7__1157 ^ p87_array_index_2060651_comb ^ p87_array_index_2060652_comb ^ p86_literal_2043916[p86_res7__1163] ^ p86_literal_2043914[p87_res7__1165_comb] ^ p86_literal_2043912[p87_res7__1167_comb] ^ p86_literal_2043910[p87_res7__1169_comb] ^ p86_bit_slice_2060399;
  assign p87_array_index_2060661_comb = p86_literal_2043920[p86_res7__1161];
  assign p87_res7__1173_comb = p86_literal_2043910[p86_bit_slice_2060386] ^ p86_literal_2043912[p86_bit_slice_2060387] ^ p86_array_index_2060403 ^ p86_array_index_2060431 ^ p86_array_index_2060457 ^ p86_array_index_2060481 ^ p86_res7__1155 ^ p86_literal_2043923[p86_res7__1157] ^ p86_res7__1159 ^ p87_array_index_2060661_comb ^ p86_literal_2043918[p86_res7__1163] ^ p86_literal_2043916[p87_res7__1165_comb] ^ p86_literal_2043914[p87_res7__1167_comb] ^ p86_literal_2043912[p87_res7__1169_comb] ^ p86_literal_2043910[p87_res7__1171_comb] ^ p86_bit_slice_2060385;
  assign p87_array_index_2060671_comb = p86_literal_2043920[p86_res7__1163];
  assign p87_res7__1175_comb = p86_literal_2043910[p86_bit_slice_2060387] ^ p86_literal_2043912[p86_bit_slice_2060388] ^ p86_array_index_2060418 ^ p86_array_index_2060445 ^ p86_array_index_2060470 ^ p87_array_index_2060629_comb ^ p86_res7__1157 ^ p86_literal_2043923[p86_res7__1159] ^ p86_res7__1161 ^ p87_array_index_2060671_comb ^ p86_literal_2043918[p87_res7__1165_comb] ^ p86_literal_2043916[p87_res7__1167_comb] ^ p86_literal_2043914[p87_res7__1169_comb] ^ p86_literal_2043912[p87_res7__1171_comb] ^ p86_literal_2043910[p87_res7__1173_comb] ^ p86_bit_slice_2060386;
  assign p87_res7__1177_comb = p86_literal_2043910[p86_bit_slice_2060388] ^ p86_array_index_2060404 ^ p86_array_index_2060432 ^ p86_array_index_2060458 ^ p86_array_index_2060482 ^ p87_array_index_2060640_comb ^ p86_res7__1159 ^ p86_literal_2043923[p86_res7__1161] ^ p86_res7__1163 ^ p86_literal_2043920[p87_res7__1165_comb] ^ p86_literal_2043918[p87_res7__1167_comb] ^ p86_literal_2043916[p87_res7__1169_comb] ^ p86_literal_2043914[p87_res7__1171_comb] ^ p86_literal_2043912[p87_res7__1173_comb] ^ p86_literal_2043910[p87_res7__1175_comb] ^ p86_bit_slice_2060387;
  assign p87_array_index_2060687_comb = p86_literal_2043910[p86_bit_slice_2060389];
  assign p87_array_index_2060688_comb = p86_literal_2043923[p86_res7__1163];
  assign p87_array_index_2060689_comb = p86_literal_2043920[p87_res7__1167_comb];
  assign p87_array_index_2060690_comb = p86_literal_2043918[p87_res7__1169_comb];
  assign p87_array_index_2060691_comb = p86_literal_2043916[p87_res7__1171_comb];
  assign p87_array_index_2060692_comb = p86_literal_2043914[p87_res7__1173_comb];
  assign p87_array_index_2060693_comb = p86_literal_2043912[p87_res7__1175_comb];
  assign p87_array_index_2060694_comb = p86_literal_2043910[p87_res7__1177_comb];
  assign p87_array_index_2060695_comb = p86_literal_2058836[p86_res7__1153];
  assign p87_array_index_2060696_comb = p86_literal_2058836[p86_res7__1155];
  assign p87_array_index_2060697_comb = p86_literal_2058836[p86_res7__1157];
  assign p87_array_index_2060698_comb = p86_literal_2058836[p86_res7__1159];

  // Registers for pipe stage 87:
  reg [127:0] p87_bit_slice_2043893;
  reg [127:0] p87_bit_slice_2044018;
  reg [127:0] p87_k3;
  reg [127:0] p87_k2;
  reg [127:0] p87_k4;
  reg [7:0] p87_bit_slice_2060388;
  reg [7:0] p87_bit_slice_2060389;
  reg [7:0] p87_bit_slice_2060390;
  reg [7:0] p87_array_index_2060405;
  reg [7:0] p87_array_index_2060419;
  reg [7:0] p87_array_index_2060420;
  reg [7:0] p87_array_index_2060433;
  reg [7:0] p87_array_index_2060446;
  reg [7:0] p87_array_index_2060447;
  reg [7:0] p87_array_index_2060459;
  reg [7:0] p87_res7__1161;
  reg [7:0] p87_array_index_2060471;
  reg [7:0] p87_array_index_2060472;
  reg [7:0] p87_res7__1163;
  reg [7:0] p87_array_index_2060483;
  reg [7:0] p87_res7__1165;
  reg [7:0] p87_array_index_2060630;
  reg [7:0] p87_array_index_2060631;
  reg [7:0] p87_res7__1167;
  reg [7:0] p87_array_index_2060641;
  reg [7:0] p87_res7__1169;
  reg [7:0] p87_array_index_2060651;
  reg [7:0] p87_array_index_2060652;
  reg [7:0] p87_res7__1171;
  reg [7:0] p87_array_index_2060661;
  reg [7:0] p87_res7__1173;
  reg [7:0] p87_array_index_2060671;
  reg [7:0] p87_res7__1175;
  reg [7:0] p87_res7__1177;
  reg [7:0] p87_array_index_2060687;
  reg [7:0] p87_array_index_2060688;
  reg [7:0] p87_array_index_2060689;
  reg [7:0] p87_array_index_2060690;
  reg [7:0] p87_array_index_2060691;
  reg [7:0] p87_array_index_2060692;
  reg [7:0] p87_array_index_2060693;
  reg [7:0] p87_array_index_2060694;
  reg [7:0] p87_array_index_2060695;
  reg [7:0] p87_array_index_2060696;
  reg [7:0] p87_array_index_2060697;
  reg [7:0] p87_array_index_2060698;
  reg [7:0] p88_literal_2043910[256];
  reg [7:0] p88_literal_2043912[256];
  reg [7:0] p88_literal_2043914[256];
  reg [7:0] p88_literal_2043916[256];
  reg [7:0] p88_literal_2043918[256];
  reg [7:0] p88_literal_2043920[256];
  reg [7:0] p88_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p87_bit_slice_2043893 <= p86_bit_slice_2043893;
    p87_bit_slice_2044018 <= p86_bit_slice_2044018;
    p87_k3 <= p86_k3;
    p87_k2 <= p86_k2;
    p87_k4 <= p86_k4;
    p87_bit_slice_2060388 <= p86_bit_slice_2060388;
    p87_bit_slice_2060389 <= p86_bit_slice_2060389;
    p87_bit_slice_2060390 <= p86_bit_slice_2060390;
    p87_array_index_2060405 <= p86_array_index_2060405;
    p87_array_index_2060419 <= p86_array_index_2060419;
    p87_array_index_2060420 <= p86_array_index_2060420;
    p87_array_index_2060433 <= p86_array_index_2060433;
    p87_array_index_2060446 <= p86_array_index_2060446;
    p87_array_index_2060447 <= p86_array_index_2060447;
    p87_array_index_2060459 <= p86_array_index_2060459;
    p87_res7__1161 <= p86_res7__1161;
    p87_array_index_2060471 <= p86_array_index_2060471;
    p87_array_index_2060472 <= p86_array_index_2060472;
    p87_res7__1163 <= p86_res7__1163;
    p87_array_index_2060483 <= p86_array_index_2060483;
    p87_res7__1165 <= p87_res7__1165_comb;
    p87_array_index_2060630 <= p87_array_index_2060630_comb;
    p87_array_index_2060631 <= p87_array_index_2060631_comb;
    p87_res7__1167 <= p87_res7__1167_comb;
    p87_array_index_2060641 <= p87_array_index_2060641_comb;
    p87_res7__1169 <= p87_res7__1169_comb;
    p87_array_index_2060651 <= p87_array_index_2060651_comb;
    p87_array_index_2060652 <= p87_array_index_2060652_comb;
    p87_res7__1171 <= p87_res7__1171_comb;
    p87_array_index_2060661 <= p87_array_index_2060661_comb;
    p87_res7__1173 <= p87_res7__1173_comb;
    p87_array_index_2060671 <= p87_array_index_2060671_comb;
    p87_res7__1175 <= p87_res7__1175_comb;
    p87_res7__1177 <= p87_res7__1177_comb;
    p87_array_index_2060687 <= p87_array_index_2060687_comb;
    p87_array_index_2060688 <= p87_array_index_2060688_comb;
    p87_array_index_2060689 <= p87_array_index_2060689_comb;
    p87_array_index_2060690 <= p87_array_index_2060690_comb;
    p87_array_index_2060691 <= p87_array_index_2060691_comb;
    p87_array_index_2060692 <= p87_array_index_2060692_comb;
    p87_array_index_2060693 <= p87_array_index_2060693_comb;
    p87_array_index_2060694 <= p87_array_index_2060694_comb;
    p87_array_index_2060695 <= p87_array_index_2060695_comb;
    p87_array_index_2060696 <= p87_array_index_2060696_comb;
    p87_array_index_2060697 <= p87_array_index_2060697_comb;
    p87_array_index_2060698 <= p87_array_index_2060698_comb;
    p88_literal_2043910 <= p87_literal_2043910;
    p88_literal_2043912 <= p87_literal_2043912;
    p88_literal_2043914 <= p87_literal_2043914;
    p88_literal_2043916 <= p87_literal_2043916;
    p88_literal_2043918 <= p87_literal_2043918;
    p88_literal_2043920 <= p87_literal_2043920;
    p88_literal_2043923 <= p87_literal_2043923;
  end

  // ===== Pipe stage 88:
  wire [7:0] p88_res7__1179_comb;
  wire [7:0] p88_res7__1181_comb;
  wire [7:0] p88_res7__1183_comb;
  wire [127:0] p88_permut__36_comb;
  wire [127:0] p88_xor_2060837_comb;
  wire [7:0] p88_bit_slice_2060840_comb;
  wire [7:0] p88_bit_slice_2060841_comb;
  wire [7:0] p88_bit_slice_2060842_comb;
  wire [7:0] p88_bit_slice_2060843_comb;
  wire [7:0] p88_bit_slice_2060844_comb;
  wire [7:0] p88_bit_slice_2060845_comb;
  wire [7:0] p88_bit_slice_2060846_comb;
  wire [7:0] p88_bit_slice_2060847_comb;
  wire [7:0] p88_bit_slice_2060848_comb;
  wire [7:0] p88_bit_slice_2060849_comb;
  wire [7:0] p88_bit_slice_2060850_comb;
  wire [7:0] p88_bit_slice_2060857_comb;
  wire [7:0] p88_bit_slice_2060859_comb;
  wire [7:0] p88_array_index_2060860_comb;
  wire [7:0] p88_array_index_2060861_comb;
  wire [7:0] p88_array_index_2060862_comb;
  wire [7:0] p88_array_index_2060863_comb;
  wire [7:0] p88_array_index_2060864_comb;
  wire [7:0] p88_array_index_2060865_comb;
  wire [7:0] p88_res7__1185_comb;
  wire [7:0] p88_array_index_2060875_comb;
  wire [7:0] p88_array_index_2060876_comb;
  wire [7:0] p88_array_index_2060877_comb;
  wire [7:0] p88_array_index_2060878_comb;
  wire [7:0] p88_array_index_2060879_comb;
  wire [7:0] p88_array_index_2060880_comb;
  wire [7:0] p88_res7__1187_comb;
  wire [7:0] p88_array_index_2060889_comb;
  wire [7:0] p88_array_index_2060890_comb;
  wire [7:0] p88_array_index_2060891_comb;
  wire [7:0] p88_array_index_2060892_comb;
  wire [7:0] p88_array_index_2060893_comb;
  wire [7:0] p88_res7__1189_comb;
  wire [7:0] p88_array_index_2060896_comb;
  wire [7:0] p88_array_index_2060897_comb;
  wire [7:0] p88_array_index_2060898_comb;
  wire [7:0] p88_array_index_2060899_comb;
  wire [7:0] p88_array_index_2060900_comb;
  wire [7:0] p88_array_index_2060901_comb;
  wire [7:0] p88_array_index_2060902_comb;
  wire [7:0] p88_array_index_2060903_comb;
  wire [7:0] p88_array_index_2060904_comb;
  wire [7:0] p88_array_index_2060905_comb;
  wire [7:0] p88_array_index_2060906_comb;
  wire [7:0] p88_array_index_2060907_comb;
  wire [7:0] p88_array_index_2060908_comb;
  assign p88_res7__1179_comb = p87_array_index_2060687 ^ p87_array_index_2060419 ^ p87_array_index_2060446 ^ p87_array_index_2060471 ^ p87_array_index_2060630 ^ p87_array_index_2060651 ^ p87_res7__1161 ^ p87_array_index_2060688 ^ p87_res7__1165 ^ p87_array_index_2060689 ^ p87_array_index_2060690 ^ p87_array_index_2060691 ^ p87_array_index_2060692 ^ p87_array_index_2060693 ^ p87_array_index_2060694 ^ p87_bit_slice_2060388;
  assign p88_res7__1181_comb = p87_array_index_2060405 ^ p87_array_index_2060433 ^ p87_array_index_2060459 ^ p87_array_index_2060483 ^ p87_array_index_2060641 ^ p87_array_index_2060661 ^ p87_res7__1163 ^ p87_literal_2043923[p87_res7__1165] ^ p87_res7__1167 ^ p87_literal_2043920[p87_res7__1169] ^ p87_literal_2043918[p87_res7__1171] ^ p87_literal_2043916[p87_res7__1173] ^ p87_literal_2043914[p87_res7__1175] ^ p87_literal_2043912[p87_res7__1177] ^ p87_literal_2043910[p88_res7__1179_comb] ^ p87_bit_slice_2060389;
  assign p88_res7__1183_comb = p87_array_index_2060420 ^ p87_array_index_2060447 ^ p87_array_index_2060472 ^ p87_array_index_2060631 ^ p87_array_index_2060652 ^ p87_array_index_2060671 ^ p87_res7__1165 ^ p87_literal_2043923[p87_res7__1167] ^ p87_res7__1169 ^ p87_literal_2043920[p87_res7__1171] ^ p87_literal_2043918[p87_res7__1173] ^ p87_literal_2043916[p87_res7__1175] ^ p87_literal_2043914[p87_res7__1177] ^ p87_literal_2043912[p88_res7__1179_comb] ^ p87_literal_2043910[p88_res7__1181_comb] ^ p87_bit_slice_2060390;
  assign p88_permut__36_comb = {p87_array_index_2060695, p87_array_index_2060696, p87_array_index_2060697, p87_array_index_2060698, p87_literal_2058836[p87_res7__1161], p87_literal_2058836[p87_res7__1163], p87_literal_2058836[p87_res7__1165], p87_literal_2058836[p87_res7__1167], p87_literal_2058836[p87_res7__1169], p87_literal_2058836[p87_res7__1171], p87_literal_2058836[p87_res7__1173], p87_literal_2058836[p87_res7__1175], p87_literal_2058836[p87_res7__1177], p87_literal_2058836[p88_res7__1179_comb], p87_literal_2058836[p88_res7__1181_comb], p87_literal_2058836[p88_res7__1183_comb]};
  assign p88_xor_2060837_comb = p87_k4 ^ p88_permut__36_comb;
  assign p88_bit_slice_2060840_comb = p88_xor_2060837_comb[103:96];
  assign p88_bit_slice_2060841_comb = p88_xor_2060837_comb[95:88];
  assign p88_bit_slice_2060842_comb = p88_xor_2060837_comb[87:80];
  assign p88_bit_slice_2060843_comb = p88_xor_2060837_comb[79:72];
  assign p88_bit_slice_2060844_comb = p88_xor_2060837_comb[63:56];
  assign p88_bit_slice_2060845_comb = p88_xor_2060837_comb[47:40];
  assign p88_bit_slice_2060846_comb = p88_xor_2060837_comb[39:32];
  assign p88_bit_slice_2060847_comb = p88_xor_2060837_comb[31:24];
  assign p88_bit_slice_2060848_comb = p88_xor_2060837_comb[23:16];
  assign p88_bit_slice_2060849_comb = p88_xor_2060837_comb[15:8];
  assign p88_bit_slice_2060850_comb = p88_xor_2060837_comb[7:0];
  assign p88_bit_slice_2060857_comb = p88_xor_2060837_comb[71:64];
  assign p88_bit_slice_2060859_comb = p88_xor_2060837_comb[55:48];
  assign p88_array_index_2060860_comb = p87_literal_2043920[p88_bit_slice_2060845_comb];
  assign p88_array_index_2060861_comb = p87_literal_2043918[p88_bit_slice_2060846_comb];
  assign p88_array_index_2060862_comb = p87_literal_2043916[p88_bit_slice_2060847_comb];
  assign p88_array_index_2060863_comb = p87_literal_2043914[p88_bit_slice_2060848_comb];
  assign p88_array_index_2060864_comb = p87_literal_2043912[p88_bit_slice_2060849_comb];
  assign p88_array_index_2060865_comb = p87_literal_2043910[p88_bit_slice_2060850_comb];
  assign p88_res7__1185_comb = p87_literal_2043910[p88_xor_2060837_comb[119:112]] ^ p87_literal_2043912[p88_xor_2060837_comb[111:104]] ^ p87_literal_2043914[p88_bit_slice_2060840_comb] ^ p87_literal_2043916[p88_bit_slice_2060841_comb] ^ p87_literal_2043918[p88_bit_slice_2060842_comb] ^ p87_literal_2043920[p88_bit_slice_2060843_comb] ^ p88_bit_slice_2060857_comb ^ p87_literal_2043923[p88_bit_slice_2060844_comb] ^ p88_bit_slice_2060859_comb ^ p88_array_index_2060860_comb ^ p88_array_index_2060861_comb ^ p88_array_index_2060862_comb ^ p88_array_index_2060863_comb ^ p88_array_index_2060864_comb ^ p88_array_index_2060865_comb ^ p88_xor_2060837_comb[127:120];
  assign p88_array_index_2060875_comb = p87_literal_2043920[p88_bit_slice_2060846_comb];
  assign p88_array_index_2060876_comb = p87_literal_2043918[p88_bit_slice_2060847_comb];
  assign p88_array_index_2060877_comb = p87_literal_2043916[p88_bit_slice_2060848_comb];
  assign p88_array_index_2060878_comb = p87_literal_2043914[p88_bit_slice_2060849_comb];
  assign p88_array_index_2060879_comb = p87_literal_2043912[p88_bit_slice_2060850_comb];
  assign p88_array_index_2060880_comb = p87_literal_2043910[p88_res7__1185_comb];
  assign p88_res7__1187_comb = p87_literal_2043910[p88_xor_2060837_comb[111:104]] ^ p87_literal_2043912[p88_bit_slice_2060840_comb] ^ p87_literal_2043914[p88_bit_slice_2060841_comb] ^ p87_literal_2043916[p88_bit_slice_2060842_comb] ^ p87_literal_2043918[p88_bit_slice_2060843_comb] ^ p87_literal_2043920[p88_bit_slice_2060857_comb] ^ p88_bit_slice_2060844_comb ^ p87_literal_2043923[p88_bit_slice_2060859_comb] ^ p88_bit_slice_2060845_comb ^ p88_array_index_2060875_comb ^ p88_array_index_2060876_comb ^ p88_array_index_2060877_comb ^ p88_array_index_2060878_comb ^ p88_array_index_2060879_comb ^ p88_array_index_2060880_comb ^ p88_xor_2060837_comb[119:112];
  assign p88_array_index_2060889_comb = p87_literal_2043920[p88_bit_slice_2060847_comb];
  assign p88_array_index_2060890_comb = p87_literal_2043918[p88_bit_slice_2060848_comb];
  assign p88_array_index_2060891_comb = p87_literal_2043916[p88_bit_slice_2060849_comb];
  assign p88_array_index_2060892_comb = p87_literal_2043914[p88_bit_slice_2060850_comb];
  assign p88_array_index_2060893_comb = p87_literal_2043912[p88_res7__1185_comb];
  assign p88_res7__1189_comb = p87_literal_2043910[p88_bit_slice_2060840_comb] ^ p87_literal_2043912[p88_bit_slice_2060841_comb] ^ p87_literal_2043914[p88_bit_slice_2060842_comb] ^ p87_literal_2043916[p88_bit_slice_2060843_comb] ^ p87_literal_2043918[p88_bit_slice_2060857_comb] ^ p87_literal_2043920[p88_bit_slice_2060844_comb] ^ p88_bit_slice_2060859_comb ^ p87_literal_2043923[p88_bit_slice_2060845_comb] ^ p88_bit_slice_2060846_comb ^ p88_array_index_2060889_comb ^ p88_array_index_2060890_comb ^ p88_array_index_2060891_comb ^ p88_array_index_2060892_comb ^ p88_array_index_2060893_comb ^ p87_literal_2043910[p88_res7__1187_comb] ^ p88_xor_2060837_comb[111:104];
  assign p88_array_index_2060896_comb = p87_literal_2043910[p88_bit_slice_2060841_comb];
  assign p88_array_index_2060897_comb = p87_literal_2043912[p88_bit_slice_2060842_comb];
  assign p88_array_index_2060898_comb = p87_literal_2043914[p88_bit_slice_2060843_comb];
  assign p88_array_index_2060899_comb = p87_literal_2043916[p88_bit_slice_2060857_comb];
  assign p88_array_index_2060900_comb = p87_literal_2043918[p88_bit_slice_2060844_comb];
  assign p88_array_index_2060901_comb = p87_literal_2043920[p88_bit_slice_2060859_comb];
  assign p88_array_index_2060902_comb = p87_literal_2043923[p88_bit_slice_2060846_comb];
  assign p88_array_index_2060903_comb = p87_literal_2043920[p88_bit_slice_2060848_comb];
  assign p88_array_index_2060904_comb = p87_literal_2043918[p88_bit_slice_2060849_comb];
  assign p88_array_index_2060905_comb = p87_literal_2043916[p88_bit_slice_2060850_comb];
  assign p88_array_index_2060906_comb = p87_literal_2043914[p88_res7__1185_comb];
  assign p88_array_index_2060907_comb = p87_literal_2043912[p88_res7__1187_comb];
  assign p88_array_index_2060908_comb = p87_literal_2043910[p88_res7__1189_comb];

  // Registers for pipe stage 88:
  reg [127:0] p88_bit_slice_2043893;
  reg [127:0] p88_bit_slice_2044018;
  reg [127:0] p88_k3;
  reg [127:0] p88_k2;
  reg [7:0] p88_bit_slice_2060840;
  reg [7:0] p88_bit_slice_2060841;
  reg [7:0] p88_bit_slice_2060842;
  reg [7:0] p88_bit_slice_2060843;
  reg [7:0] p88_bit_slice_2060844;
  reg [7:0] p88_bit_slice_2060845;
  reg [7:0] p88_bit_slice_2060846;
  reg [7:0] p88_bit_slice_2060847;
  reg [7:0] p88_bit_slice_2060848;
  reg [7:0] p88_bit_slice_2060849;
  reg [7:0] p88_bit_slice_2060850;
  reg [7:0] p88_bit_slice_2060857;
  reg [7:0] p88_bit_slice_2060859;
  reg [7:0] p88_array_index_2060860;
  reg [7:0] p88_array_index_2060861;
  reg [7:0] p88_array_index_2060862;
  reg [7:0] p88_array_index_2060863;
  reg [7:0] p88_array_index_2060864;
  reg [7:0] p88_array_index_2060865;
  reg [7:0] p88_res7__1185;
  reg [7:0] p88_array_index_2060875;
  reg [7:0] p88_array_index_2060876;
  reg [7:0] p88_array_index_2060877;
  reg [7:0] p88_array_index_2060878;
  reg [7:0] p88_array_index_2060879;
  reg [7:0] p88_array_index_2060880;
  reg [7:0] p88_res7__1187;
  reg [7:0] p88_array_index_2060889;
  reg [7:0] p88_array_index_2060890;
  reg [7:0] p88_array_index_2060891;
  reg [7:0] p88_array_index_2060892;
  reg [7:0] p88_array_index_2060893;
  reg [7:0] p88_res7__1189;
  reg [7:0] p88_array_index_2060896;
  reg [7:0] p88_array_index_2060897;
  reg [7:0] p88_array_index_2060898;
  reg [7:0] p88_array_index_2060899;
  reg [7:0] p88_array_index_2060900;
  reg [7:0] p88_array_index_2060901;
  reg [7:0] p88_array_index_2060902;
  reg [7:0] p88_array_index_2060903;
  reg [7:0] p88_array_index_2060904;
  reg [7:0] p88_array_index_2060905;
  reg [7:0] p88_array_index_2060906;
  reg [7:0] p88_array_index_2060907;
  reg [7:0] p88_array_index_2060908;
  reg [7:0] p89_literal_2043910[256];
  reg [7:0] p89_literal_2043912[256];
  reg [7:0] p89_literal_2043914[256];
  reg [7:0] p89_literal_2043916[256];
  reg [7:0] p89_literal_2043918[256];
  reg [7:0] p89_literal_2043920[256];
  reg [7:0] p89_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p88_bit_slice_2043893 <= p87_bit_slice_2043893;
    p88_bit_slice_2044018 <= p87_bit_slice_2044018;
    p88_k3 <= p87_k3;
    p88_k2 <= p87_k2;
    p88_bit_slice_2060840 <= p88_bit_slice_2060840_comb;
    p88_bit_slice_2060841 <= p88_bit_slice_2060841_comb;
    p88_bit_slice_2060842 <= p88_bit_slice_2060842_comb;
    p88_bit_slice_2060843 <= p88_bit_slice_2060843_comb;
    p88_bit_slice_2060844 <= p88_bit_slice_2060844_comb;
    p88_bit_slice_2060845 <= p88_bit_slice_2060845_comb;
    p88_bit_slice_2060846 <= p88_bit_slice_2060846_comb;
    p88_bit_slice_2060847 <= p88_bit_slice_2060847_comb;
    p88_bit_slice_2060848 <= p88_bit_slice_2060848_comb;
    p88_bit_slice_2060849 <= p88_bit_slice_2060849_comb;
    p88_bit_slice_2060850 <= p88_bit_slice_2060850_comb;
    p88_bit_slice_2060857 <= p88_bit_slice_2060857_comb;
    p88_bit_slice_2060859 <= p88_bit_slice_2060859_comb;
    p88_array_index_2060860 <= p88_array_index_2060860_comb;
    p88_array_index_2060861 <= p88_array_index_2060861_comb;
    p88_array_index_2060862 <= p88_array_index_2060862_comb;
    p88_array_index_2060863 <= p88_array_index_2060863_comb;
    p88_array_index_2060864 <= p88_array_index_2060864_comb;
    p88_array_index_2060865 <= p88_array_index_2060865_comb;
    p88_res7__1185 <= p88_res7__1185_comb;
    p88_array_index_2060875 <= p88_array_index_2060875_comb;
    p88_array_index_2060876 <= p88_array_index_2060876_comb;
    p88_array_index_2060877 <= p88_array_index_2060877_comb;
    p88_array_index_2060878 <= p88_array_index_2060878_comb;
    p88_array_index_2060879 <= p88_array_index_2060879_comb;
    p88_array_index_2060880 <= p88_array_index_2060880_comb;
    p88_res7__1187 <= p88_res7__1187_comb;
    p88_array_index_2060889 <= p88_array_index_2060889_comb;
    p88_array_index_2060890 <= p88_array_index_2060890_comb;
    p88_array_index_2060891 <= p88_array_index_2060891_comb;
    p88_array_index_2060892 <= p88_array_index_2060892_comb;
    p88_array_index_2060893 <= p88_array_index_2060893_comb;
    p88_res7__1189 <= p88_res7__1189_comb;
    p88_array_index_2060896 <= p88_array_index_2060896_comb;
    p88_array_index_2060897 <= p88_array_index_2060897_comb;
    p88_array_index_2060898 <= p88_array_index_2060898_comb;
    p88_array_index_2060899 <= p88_array_index_2060899_comb;
    p88_array_index_2060900 <= p88_array_index_2060900_comb;
    p88_array_index_2060901 <= p88_array_index_2060901_comb;
    p88_array_index_2060902 <= p88_array_index_2060902_comb;
    p88_array_index_2060903 <= p88_array_index_2060903_comb;
    p88_array_index_2060904 <= p88_array_index_2060904_comb;
    p88_array_index_2060905 <= p88_array_index_2060905_comb;
    p88_array_index_2060906 <= p88_array_index_2060906_comb;
    p88_array_index_2060907 <= p88_array_index_2060907_comb;
    p88_array_index_2060908 <= p88_array_index_2060908_comb;
    p89_literal_2043910 <= p88_literal_2043910;
    p89_literal_2043912 <= p88_literal_2043912;
    p89_literal_2043914 <= p88_literal_2043914;
    p89_literal_2043916 <= p88_literal_2043916;
    p89_literal_2043918 <= p88_literal_2043918;
    p89_literal_2043920 <= p88_literal_2043920;
    p89_literal_2043923 <= p88_literal_2043923;
  end

  // ===== Pipe stage 89:
  wire [7:0] p89_res7__1191_comb;
  wire [7:0] p89_array_index_2061032_comb;
  wire [7:0] p89_array_index_2061033_comb;
  wire [7:0] p89_array_index_2061034_comb;
  wire [7:0] p89_array_index_2061035_comb;
  wire [7:0] p89_res7__1193_comb;
  wire [7:0] p89_array_index_2061045_comb;
  wire [7:0] p89_array_index_2061046_comb;
  wire [7:0] p89_array_index_2061047_comb;
  wire [7:0] p89_array_index_2061048_comb;
  wire [7:0] p89_res7__1195_comb;
  wire [7:0] p89_array_index_2061057_comb;
  wire [7:0] p89_array_index_2061058_comb;
  wire [7:0] p89_array_index_2061059_comb;
  wire [7:0] p89_res7__1197_comb;
  wire [7:0] p89_array_index_2061069_comb;
  wire [7:0] p89_array_index_2061070_comb;
  wire [7:0] p89_array_index_2061071_comb;
  wire [7:0] p89_res7__1199_comb;
  wire [7:0] p89_array_index_2061080_comb;
  wire [7:0] p89_array_index_2061081_comb;
  wire [7:0] p89_res7__1201_comb;
  wire [7:0] p89_array_index_2061091_comb;
  wire [7:0] p89_array_index_2061092_comb;
  wire [7:0] p89_res7__1203_comb;
  wire [7:0] p89_array_index_2061098_comb;
  wire [7:0] p89_array_index_2061099_comb;
  wire [7:0] p89_array_index_2061100_comb;
  wire [7:0] p89_array_index_2061101_comb;
  wire [7:0] p89_array_index_2061102_comb;
  wire [7:0] p89_array_index_2061103_comb;
  wire [7:0] p89_array_index_2061104_comb;
  wire [7:0] p89_array_index_2061105_comb;
  wire [7:0] p89_array_index_2061106_comb;
  wire [7:0] p89_array_index_2061107_comb;
  assign p89_res7__1191_comb = p88_array_index_2060896 ^ p88_array_index_2060897 ^ p88_array_index_2060898 ^ p88_array_index_2060899 ^ p88_array_index_2060900 ^ p88_array_index_2060901 ^ p88_bit_slice_2060845 ^ p88_array_index_2060902 ^ p88_bit_slice_2060847 ^ p88_array_index_2060903 ^ p88_array_index_2060904 ^ p88_array_index_2060905 ^ p88_array_index_2060906 ^ p88_array_index_2060907 ^ p88_array_index_2060908 ^ p88_bit_slice_2060840;
  assign p89_array_index_2061032_comb = p88_literal_2043920[p88_bit_slice_2060849];
  assign p89_array_index_2061033_comb = p88_literal_2043918[p88_bit_slice_2060850];
  assign p89_array_index_2061034_comb = p88_literal_2043916[p88_res7__1185];
  assign p89_array_index_2061035_comb = p88_literal_2043914[p88_res7__1187];
  assign p89_res7__1193_comb = p88_literal_2043910[p88_bit_slice_2060842] ^ p88_literal_2043912[p88_bit_slice_2060843] ^ p88_literal_2043914[p88_bit_slice_2060857] ^ p88_literal_2043916[p88_bit_slice_2060844] ^ p88_literal_2043918[p88_bit_slice_2060859] ^ p88_array_index_2060860 ^ p88_bit_slice_2060846 ^ p88_literal_2043923[p88_bit_slice_2060847] ^ p88_bit_slice_2060848 ^ p89_array_index_2061032_comb ^ p89_array_index_2061033_comb ^ p89_array_index_2061034_comb ^ p89_array_index_2061035_comb ^ p88_literal_2043912[p88_res7__1189] ^ p88_literal_2043910[p89_res7__1191_comb] ^ p88_bit_slice_2060841;
  assign p89_array_index_2061045_comb = p88_literal_2043920[p88_bit_slice_2060850];
  assign p89_array_index_2061046_comb = p88_literal_2043918[p88_res7__1185];
  assign p89_array_index_2061047_comb = p88_literal_2043916[p88_res7__1187];
  assign p89_array_index_2061048_comb = p88_literal_2043914[p88_res7__1189];
  assign p89_res7__1195_comb = p88_literal_2043910[p88_bit_slice_2060843] ^ p88_literal_2043912[p88_bit_slice_2060857] ^ p88_literal_2043914[p88_bit_slice_2060844] ^ p88_literal_2043916[p88_bit_slice_2060859] ^ p88_literal_2043918[p88_bit_slice_2060845] ^ p88_array_index_2060875 ^ p88_bit_slice_2060847 ^ p88_literal_2043923[p88_bit_slice_2060848] ^ p88_bit_slice_2060849 ^ p89_array_index_2061045_comb ^ p89_array_index_2061046_comb ^ p89_array_index_2061047_comb ^ p89_array_index_2061048_comb ^ p88_literal_2043912[p89_res7__1191_comb] ^ p88_literal_2043910[p89_res7__1193_comb] ^ p88_bit_slice_2060842;
  assign p89_array_index_2061057_comb = p88_literal_2043920[p88_res7__1185];
  assign p89_array_index_2061058_comb = p88_literal_2043918[p88_res7__1187];
  assign p89_array_index_2061059_comb = p88_literal_2043916[p88_res7__1189];
  assign p89_res7__1197_comb = p88_literal_2043910[p88_bit_slice_2060857] ^ p88_literal_2043912[p88_bit_slice_2060844] ^ p88_literal_2043914[p88_bit_slice_2060859] ^ p88_literal_2043916[p88_bit_slice_2060845] ^ p88_array_index_2060861 ^ p88_array_index_2060889 ^ p88_bit_slice_2060848 ^ p88_literal_2043923[p88_bit_slice_2060849] ^ p88_bit_slice_2060850 ^ p89_array_index_2061057_comb ^ p89_array_index_2061058_comb ^ p89_array_index_2061059_comb ^ p88_literal_2043914[p89_res7__1191_comb] ^ p88_literal_2043912[p89_res7__1193_comb] ^ p88_literal_2043910[p89_res7__1195_comb] ^ p88_bit_slice_2060843;
  assign p89_array_index_2061069_comb = p88_literal_2043920[p88_res7__1187];
  assign p89_array_index_2061070_comb = p88_literal_2043918[p88_res7__1189];
  assign p89_array_index_2061071_comb = p88_literal_2043916[p89_res7__1191_comb];
  assign p89_res7__1199_comb = p88_literal_2043910[p88_bit_slice_2060844] ^ p88_literal_2043912[p88_bit_slice_2060859] ^ p88_literal_2043914[p88_bit_slice_2060845] ^ p88_literal_2043916[p88_bit_slice_2060846] ^ p88_array_index_2060876 ^ p88_array_index_2060903 ^ p88_bit_slice_2060849 ^ p88_literal_2043923[p88_bit_slice_2060850] ^ p88_res7__1185 ^ p89_array_index_2061069_comb ^ p89_array_index_2061070_comb ^ p89_array_index_2061071_comb ^ p88_literal_2043914[p89_res7__1193_comb] ^ p88_literal_2043912[p89_res7__1195_comb] ^ p88_literal_2043910[p89_res7__1197_comb] ^ p88_bit_slice_2060857;
  assign p89_array_index_2061080_comb = p88_literal_2043920[p88_res7__1189];
  assign p89_array_index_2061081_comb = p88_literal_2043918[p89_res7__1191_comb];
  assign p89_res7__1201_comb = p88_literal_2043910[p88_bit_slice_2060859] ^ p88_literal_2043912[p88_bit_slice_2060845] ^ p88_literal_2043914[p88_bit_slice_2060846] ^ p88_array_index_2060862 ^ p88_array_index_2060890 ^ p89_array_index_2061032_comb ^ p88_bit_slice_2060850 ^ p88_literal_2043923[p88_res7__1185] ^ p88_res7__1187 ^ p89_array_index_2061080_comb ^ p89_array_index_2061081_comb ^ p88_literal_2043916[p89_res7__1193_comb] ^ p88_literal_2043914[p89_res7__1195_comb] ^ p88_literal_2043912[p89_res7__1197_comb] ^ p88_literal_2043910[p89_res7__1199_comb] ^ p88_bit_slice_2060844;
  assign p89_array_index_2061091_comb = p88_literal_2043920[p89_res7__1191_comb];
  assign p89_array_index_2061092_comb = p88_literal_2043918[p89_res7__1193_comb];
  assign p89_res7__1203_comb = p88_literal_2043910[p88_bit_slice_2060845] ^ p88_literal_2043912[p88_bit_slice_2060846] ^ p88_literal_2043914[p88_bit_slice_2060847] ^ p88_array_index_2060877 ^ p88_array_index_2060904 ^ p89_array_index_2061045_comb ^ p88_res7__1185 ^ p88_literal_2043923[p88_res7__1187] ^ p88_res7__1189 ^ p89_array_index_2061091_comb ^ p89_array_index_2061092_comb ^ p88_literal_2043916[p89_res7__1195_comb] ^ p88_literal_2043914[p89_res7__1197_comb] ^ p88_literal_2043912[p89_res7__1199_comb] ^ p88_literal_2043910[p89_res7__1201_comb] ^ p88_bit_slice_2060859;
  assign p89_array_index_2061098_comb = p88_literal_2043910[p88_bit_slice_2060846];
  assign p89_array_index_2061099_comb = p88_literal_2043912[p88_bit_slice_2060847];
  assign p89_array_index_2061100_comb = p88_literal_2043923[p88_res7__1189];
  assign p89_array_index_2061101_comb = p88_literal_2043920[p89_res7__1193_comb];
  assign p89_array_index_2061102_comb = p88_literal_2043918[p89_res7__1195_comb];
  assign p89_array_index_2061103_comb = p88_literal_2043916[p89_res7__1197_comb];
  assign p89_array_index_2061104_comb = p88_literal_2043914[p89_res7__1199_comb];
  assign p89_array_index_2061105_comb = p88_literal_2043912[p89_res7__1201_comb];
  assign p89_array_index_2061106_comb = p88_literal_2043910[p89_res7__1203_comb];
  assign p89_array_index_2061107_comb = p88_literal_2058836[p88_res7__1185];

  // Registers for pipe stage 89:
  reg [127:0] p89_bit_slice_2043893;
  reg [127:0] p89_bit_slice_2044018;
  reg [127:0] p89_k3;
  reg [127:0] p89_k2;
  reg [7:0] p89_bit_slice_2060845;
  reg [7:0] p89_bit_slice_2060846;
  reg [7:0] p89_bit_slice_2060847;
  reg [7:0] p89_bit_slice_2060848;
  reg [7:0] p89_bit_slice_2060849;
  reg [7:0] p89_bit_slice_2060850;
  reg [7:0] p89_array_index_2060863;
  reg [7:0] p89_array_index_2060864;
  reg [7:0] p89_array_index_2060865;
  reg [7:0] p89_array_index_2060878;
  reg [7:0] p89_array_index_2060879;
  reg [7:0] p89_array_index_2060880;
  reg [7:0] p89_res7__1187;
  reg [7:0] p89_array_index_2060891;
  reg [7:0] p89_array_index_2060892;
  reg [7:0] p89_array_index_2060893;
  reg [7:0] p89_res7__1189;
  reg [7:0] p89_array_index_2060905;
  reg [7:0] p89_array_index_2060906;
  reg [7:0] p89_array_index_2060907;
  reg [7:0] p89_res7__1191;
  reg [7:0] p89_array_index_2061033;
  reg [7:0] p89_array_index_2061034;
  reg [7:0] p89_array_index_2061035;
  reg [7:0] p89_res7__1193;
  reg [7:0] p89_array_index_2061046;
  reg [7:0] p89_array_index_2061047;
  reg [7:0] p89_array_index_2061048;
  reg [7:0] p89_res7__1195;
  reg [7:0] p89_array_index_2061057;
  reg [7:0] p89_array_index_2061058;
  reg [7:0] p89_array_index_2061059;
  reg [7:0] p89_res7__1197;
  reg [7:0] p89_array_index_2061069;
  reg [7:0] p89_array_index_2061070;
  reg [7:0] p89_array_index_2061071;
  reg [7:0] p89_res7__1199;
  reg [7:0] p89_array_index_2061080;
  reg [7:0] p89_array_index_2061081;
  reg [7:0] p89_res7__1201;
  reg [7:0] p89_array_index_2061091;
  reg [7:0] p89_array_index_2061092;
  reg [7:0] p89_res7__1203;
  reg [7:0] p89_array_index_2061098;
  reg [7:0] p89_array_index_2061099;
  reg [7:0] p89_array_index_2061100;
  reg [7:0] p89_array_index_2061101;
  reg [7:0] p89_array_index_2061102;
  reg [7:0] p89_array_index_2061103;
  reg [7:0] p89_array_index_2061104;
  reg [7:0] p89_array_index_2061105;
  reg [7:0] p89_array_index_2061106;
  reg [7:0] p89_array_index_2061107;
  reg [7:0] p90_literal_2043910[256];
  reg [7:0] p90_literal_2043912[256];
  reg [7:0] p90_literal_2043914[256];
  reg [7:0] p90_literal_2043916[256];
  reg [7:0] p90_literal_2043918[256];
  reg [7:0] p90_literal_2043920[256];
  reg [7:0] p90_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p89_bit_slice_2043893 <= p88_bit_slice_2043893;
    p89_bit_slice_2044018 <= p88_bit_slice_2044018;
    p89_k3 <= p88_k3;
    p89_k2 <= p88_k2;
    p89_bit_slice_2060845 <= p88_bit_slice_2060845;
    p89_bit_slice_2060846 <= p88_bit_slice_2060846;
    p89_bit_slice_2060847 <= p88_bit_slice_2060847;
    p89_bit_slice_2060848 <= p88_bit_slice_2060848;
    p89_bit_slice_2060849 <= p88_bit_slice_2060849;
    p89_bit_slice_2060850 <= p88_bit_slice_2060850;
    p89_array_index_2060863 <= p88_array_index_2060863;
    p89_array_index_2060864 <= p88_array_index_2060864;
    p89_array_index_2060865 <= p88_array_index_2060865;
    p89_array_index_2060878 <= p88_array_index_2060878;
    p89_array_index_2060879 <= p88_array_index_2060879;
    p89_array_index_2060880 <= p88_array_index_2060880;
    p89_res7__1187 <= p88_res7__1187;
    p89_array_index_2060891 <= p88_array_index_2060891;
    p89_array_index_2060892 <= p88_array_index_2060892;
    p89_array_index_2060893 <= p88_array_index_2060893;
    p89_res7__1189 <= p88_res7__1189;
    p89_array_index_2060905 <= p88_array_index_2060905;
    p89_array_index_2060906 <= p88_array_index_2060906;
    p89_array_index_2060907 <= p88_array_index_2060907;
    p89_res7__1191 <= p89_res7__1191_comb;
    p89_array_index_2061033 <= p89_array_index_2061033_comb;
    p89_array_index_2061034 <= p89_array_index_2061034_comb;
    p89_array_index_2061035 <= p89_array_index_2061035_comb;
    p89_res7__1193 <= p89_res7__1193_comb;
    p89_array_index_2061046 <= p89_array_index_2061046_comb;
    p89_array_index_2061047 <= p89_array_index_2061047_comb;
    p89_array_index_2061048 <= p89_array_index_2061048_comb;
    p89_res7__1195 <= p89_res7__1195_comb;
    p89_array_index_2061057 <= p89_array_index_2061057_comb;
    p89_array_index_2061058 <= p89_array_index_2061058_comb;
    p89_array_index_2061059 <= p89_array_index_2061059_comb;
    p89_res7__1197 <= p89_res7__1197_comb;
    p89_array_index_2061069 <= p89_array_index_2061069_comb;
    p89_array_index_2061070 <= p89_array_index_2061070_comb;
    p89_array_index_2061071 <= p89_array_index_2061071_comb;
    p89_res7__1199 <= p89_res7__1199_comb;
    p89_array_index_2061080 <= p89_array_index_2061080_comb;
    p89_array_index_2061081 <= p89_array_index_2061081_comb;
    p89_res7__1201 <= p89_res7__1201_comb;
    p89_array_index_2061091 <= p89_array_index_2061091_comb;
    p89_array_index_2061092 <= p89_array_index_2061092_comb;
    p89_res7__1203 <= p89_res7__1203_comb;
    p89_array_index_2061098 <= p89_array_index_2061098_comb;
    p89_array_index_2061099 <= p89_array_index_2061099_comb;
    p89_array_index_2061100 <= p89_array_index_2061100_comb;
    p89_array_index_2061101 <= p89_array_index_2061101_comb;
    p89_array_index_2061102 <= p89_array_index_2061102_comb;
    p89_array_index_2061103 <= p89_array_index_2061103_comb;
    p89_array_index_2061104 <= p89_array_index_2061104_comb;
    p89_array_index_2061105 <= p89_array_index_2061105_comb;
    p89_array_index_2061106 <= p89_array_index_2061106_comb;
    p89_array_index_2061107 <= p89_array_index_2061107_comb;
    p90_literal_2043910 <= p89_literal_2043910;
    p90_literal_2043912 <= p89_literal_2043912;
    p90_literal_2043914 <= p89_literal_2043914;
    p90_literal_2043916 <= p89_literal_2043916;
    p90_literal_2043918 <= p89_literal_2043918;
    p90_literal_2043920 <= p89_literal_2043920;
    p90_literal_2043923 <= p89_literal_2043923;
  end

  // ===== Pipe stage 90:
  wire [7:0] p90_res7__1205_comb;
  wire [7:0] p90_array_index_2061242_comb;
  wire [7:0] p90_res7__1207_comb;
  wire [7:0] p90_res7__1209_comb;
  wire [7:0] p90_res7__1211_comb;
  wire [7:0] p90_res7__1213_comb;
  wire [7:0] p90_res7__1215_comb;
  wire [127:0] p90_permut__37_comb;
  wire [127:0] p90_xor_2061299_comb;
  wire [7:0] p90_bit_slice_2061300_comb;
  wire [7:0] p90_bit_slice_2061301_comb;
  wire [7:0] p90_bit_slice_2061302_comb;
  wire [7:0] p90_bit_slice_2061303_comb;
  wire [7:0] p90_bit_slice_2061304_comb;
  wire [7:0] p90_bit_slice_2061305_comb;
  wire [7:0] p90_bit_slice_2061306_comb;
  wire [7:0] p90_bit_slice_2061307_comb;
  wire [7:0] p90_bit_slice_2061308_comb;
  wire [7:0] p90_bit_slice_2061309_comb;
  wire [7:0] p90_bit_slice_2061310_comb;
  wire [7:0] p90_bit_slice_2061311_comb;
  wire [7:0] p90_bit_slice_2061312_comb;
  wire [7:0] p90_array_index_2061313_comb;
  wire [7:0] p90_array_index_2061314_comb;
  wire [7:0] p90_array_index_2061315_comb;
  wire [7:0] p90_array_index_2061316_comb;
  wire [7:0] p90_array_index_2061317_comb;
  wire [7:0] p90_array_index_2061318_comb;
  wire [7:0] p90_bit_slice_2061319_comb;
  wire [7:0] p90_array_index_2061320_comb;
  wire [7:0] p90_bit_slice_2061321_comb;
  wire [7:0] p90_array_index_2061322_comb;
  wire [7:0] p90_array_index_2061323_comb;
  wire [7:0] p90_array_index_2061324_comb;
  wire [7:0] p90_array_index_2061325_comb;
  wire [7:0] p90_array_index_2061326_comb;
  wire [7:0] p90_array_index_2061327_comb;
  wire [7:0] p90_bit_slice_2061328_comb;
  assign p90_res7__1205_comb = p89_array_index_2061098 ^ p89_array_index_2061099 ^ p89_array_index_2060863 ^ p89_array_index_2060891 ^ p89_array_index_2061033 ^ p89_array_index_2061057 ^ p89_res7__1187 ^ p89_array_index_2061100 ^ p89_res7__1191 ^ p89_array_index_2061101 ^ p89_array_index_2061102 ^ p89_array_index_2061103 ^ p89_array_index_2061104 ^ p89_array_index_2061105 ^ p89_array_index_2061106 ^ p89_bit_slice_2060845;
  assign p90_array_index_2061242_comb = p89_literal_2043920[p89_res7__1195];
  assign p90_res7__1207_comb = p89_literal_2043910[p89_bit_slice_2060847] ^ p89_literal_2043912[p89_bit_slice_2060848] ^ p89_array_index_2060878 ^ p89_array_index_2060905 ^ p89_array_index_2061046 ^ p89_array_index_2061069 ^ p89_res7__1189 ^ p89_literal_2043923[p89_res7__1191] ^ p89_res7__1193 ^ p90_array_index_2061242_comb ^ p89_literal_2043918[p89_res7__1197] ^ p89_literal_2043916[p89_res7__1199] ^ p89_literal_2043914[p89_res7__1201] ^ p89_literal_2043912[p89_res7__1203] ^ p89_literal_2043910[p90_res7__1205_comb] ^ p89_bit_slice_2060846;
  assign p90_res7__1209_comb = p89_literal_2043910[p89_bit_slice_2060848] ^ p89_array_index_2060864 ^ p89_array_index_2060892 ^ p89_array_index_2061034 ^ p89_array_index_2061058 ^ p89_array_index_2061080 ^ p89_res7__1191 ^ p89_literal_2043923[p89_res7__1193] ^ p89_res7__1195 ^ p89_literal_2043920[p89_res7__1197] ^ p89_literal_2043918[p89_res7__1199] ^ p89_literal_2043916[p89_res7__1201] ^ p89_literal_2043914[p89_res7__1203] ^ p89_literal_2043912[p90_res7__1205_comb] ^ p89_literal_2043910[p90_res7__1207_comb] ^ p89_bit_slice_2060847;
  assign p90_res7__1211_comb = p89_literal_2043910[p89_bit_slice_2060849] ^ p89_array_index_2060879 ^ p89_array_index_2060906 ^ p89_array_index_2061047 ^ p89_array_index_2061070 ^ p89_array_index_2061091 ^ p89_res7__1193 ^ p89_literal_2043923[p89_res7__1195] ^ p89_res7__1197 ^ p89_literal_2043920[p89_res7__1199] ^ p89_literal_2043918[p89_res7__1201] ^ p89_literal_2043916[p89_res7__1203] ^ p89_literal_2043914[p90_res7__1205_comb] ^ p89_literal_2043912[p90_res7__1207_comb] ^ p89_literal_2043910[p90_res7__1209_comb] ^ p89_bit_slice_2060848;
  assign p90_res7__1213_comb = p89_array_index_2060865 ^ p89_array_index_2060893 ^ p89_array_index_2061035 ^ p89_array_index_2061059 ^ p89_array_index_2061081 ^ p89_array_index_2061101 ^ p89_res7__1195 ^ p89_literal_2043923[p89_res7__1197] ^ p89_res7__1199 ^ p89_literal_2043920[p89_res7__1201] ^ p89_literal_2043918[p89_res7__1203] ^ p89_literal_2043916[p90_res7__1205_comb] ^ p89_literal_2043914[p90_res7__1207_comb] ^ p89_literal_2043912[p90_res7__1209_comb] ^ p89_literal_2043910[p90_res7__1211_comb] ^ p89_bit_slice_2060849;
  assign p90_res7__1215_comb = p89_array_index_2060880 ^ p89_array_index_2060907 ^ p89_array_index_2061048 ^ p89_array_index_2061071 ^ p89_array_index_2061092 ^ p90_array_index_2061242_comb ^ p89_res7__1197 ^ p89_literal_2043923[p89_res7__1199] ^ p89_res7__1201 ^ p89_literal_2043920[p89_res7__1203] ^ p89_literal_2043918[p90_res7__1205_comb] ^ p89_literal_2043916[p90_res7__1207_comb] ^ p89_literal_2043914[p90_res7__1209_comb] ^ p89_literal_2043912[p90_res7__1211_comb] ^ p89_literal_2043910[p90_res7__1213_comb] ^ p89_bit_slice_2060850;
  assign p90_permut__37_comb = {p89_array_index_2061107, p89_literal_2058836[p89_res7__1187], p89_literal_2058836[p89_res7__1189], p89_literal_2058836[p89_res7__1191], p89_literal_2058836[p89_res7__1193], p89_literal_2058836[p89_res7__1195], p89_literal_2058836[p89_res7__1197], p89_literal_2058836[p89_res7__1199], p89_literal_2058836[p89_res7__1201], p89_literal_2058836[p89_res7__1203], p89_literal_2058836[p90_res7__1205_comb], p89_literal_2058836[p90_res7__1207_comb], p89_literal_2058836[p90_res7__1209_comb], p89_literal_2058836[p90_res7__1211_comb], p89_literal_2058836[p90_res7__1213_comb], p89_literal_2058836[p90_res7__1215_comb]};
  assign p90_xor_2061299_comb = p89_k3 ^ p90_permut__37_comb;
  assign p90_bit_slice_2061300_comb = p90_xor_2061299_comb[119:112];
  assign p90_bit_slice_2061301_comb = p90_xor_2061299_comb[111:104];
  assign p90_bit_slice_2061302_comb = p90_xor_2061299_comb[103:96];
  assign p90_bit_slice_2061303_comb = p90_xor_2061299_comb[95:88];
  assign p90_bit_slice_2061304_comb = p90_xor_2061299_comb[87:80];
  assign p90_bit_slice_2061305_comb = p90_xor_2061299_comb[79:72];
  assign p90_bit_slice_2061306_comb = p90_xor_2061299_comb[63:56];
  assign p90_bit_slice_2061307_comb = p90_xor_2061299_comb[47:40];
  assign p90_bit_slice_2061308_comb = p90_xor_2061299_comb[39:32];
  assign p90_bit_slice_2061309_comb = p90_xor_2061299_comb[31:24];
  assign p90_bit_slice_2061310_comb = p90_xor_2061299_comb[23:16];
  assign p90_bit_slice_2061311_comb = p90_xor_2061299_comb[15:8];
  assign p90_bit_slice_2061312_comb = p90_xor_2061299_comb[7:0];
  assign p90_array_index_2061313_comb = p89_literal_2043910[p90_bit_slice_2061300_comb];
  assign p90_array_index_2061314_comb = p89_literal_2043912[p90_bit_slice_2061301_comb];
  assign p90_array_index_2061315_comb = p89_literal_2043914[p90_bit_slice_2061302_comb];
  assign p90_array_index_2061316_comb = p89_literal_2043916[p90_bit_slice_2061303_comb];
  assign p90_array_index_2061317_comb = p89_literal_2043918[p90_bit_slice_2061304_comb];
  assign p90_array_index_2061318_comb = p89_literal_2043920[p90_bit_slice_2061305_comb];
  assign p90_bit_slice_2061319_comb = p90_xor_2061299_comb[71:64];
  assign p90_array_index_2061320_comb = p89_literal_2043923[p90_bit_slice_2061306_comb];
  assign p90_bit_slice_2061321_comb = p90_xor_2061299_comb[55:48];
  assign p90_array_index_2061322_comb = p89_literal_2043920[p90_bit_slice_2061307_comb];
  assign p90_array_index_2061323_comb = p89_literal_2043918[p90_bit_slice_2061308_comb];
  assign p90_array_index_2061324_comb = p89_literal_2043916[p90_bit_slice_2061309_comb];
  assign p90_array_index_2061325_comb = p89_literal_2043914[p90_bit_slice_2061310_comb];
  assign p90_array_index_2061326_comb = p89_literal_2043912[p90_bit_slice_2061311_comb];
  assign p90_array_index_2061327_comb = p89_literal_2043910[p90_bit_slice_2061312_comb];
  assign p90_bit_slice_2061328_comb = p90_xor_2061299_comb[127:120];

  // Registers for pipe stage 90:
  reg [127:0] p90_bit_slice_2043893;
  reg [127:0] p90_bit_slice_2044018;
  reg [127:0] p90_k2;
  reg [7:0] p90_bit_slice_2061300;
  reg [7:0] p90_bit_slice_2061301;
  reg [7:0] p90_bit_slice_2061302;
  reg [7:0] p90_bit_slice_2061303;
  reg [7:0] p90_bit_slice_2061304;
  reg [7:0] p90_bit_slice_2061305;
  reg [7:0] p90_bit_slice_2061306;
  reg [7:0] p90_bit_slice_2061307;
  reg [7:0] p90_bit_slice_2061308;
  reg [7:0] p90_bit_slice_2061309;
  reg [7:0] p90_bit_slice_2061310;
  reg [7:0] p90_bit_slice_2061311;
  reg [7:0] p90_bit_slice_2061312;
  reg [7:0] p90_array_index_2061313;
  reg [7:0] p90_array_index_2061314;
  reg [7:0] p90_array_index_2061315;
  reg [7:0] p90_array_index_2061316;
  reg [7:0] p90_array_index_2061317;
  reg [7:0] p90_array_index_2061318;
  reg [7:0] p90_bit_slice_2061319;
  reg [7:0] p90_array_index_2061320;
  reg [7:0] p90_bit_slice_2061321;
  reg [7:0] p90_array_index_2061322;
  reg [7:0] p90_array_index_2061323;
  reg [7:0] p90_array_index_2061324;
  reg [7:0] p90_array_index_2061325;
  reg [7:0] p90_array_index_2061326;
  reg [7:0] p90_array_index_2061327;
  reg [7:0] p90_bit_slice_2061328;
  reg [7:0] p91_literal_2043910[256];
  reg [7:0] p91_literal_2043912[256];
  reg [7:0] p91_literal_2043914[256];
  reg [7:0] p91_literal_2043916[256];
  reg [7:0] p91_literal_2043918[256];
  reg [7:0] p91_literal_2043920[256];
  reg [7:0] p91_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p90_bit_slice_2043893 <= p89_bit_slice_2043893;
    p90_bit_slice_2044018 <= p89_bit_slice_2044018;
    p90_k2 <= p89_k2;
    p90_bit_slice_2061300 <= p90_bit_slice_2061300_comb;
    p90_bit_slice_2061301 <= p90_bit_slice_2061301_comb;
    p90_bit_slice_2061302 <= p90_bit_slice_2061302_comb;
    p90_bit_slice_2061303 <= p90_bit_slice_2061303_comb;
    p90_bit_slice_2061304 <= p90_bit_slice_2061304_comb;
    p90_bit_slice_2061305 <= p90_bit_slice_2061305_comb;
    p90_bit_slice_2061306 <= p90_bit_slice_2061306_comb;
    p90_bit_slice_2061307 <= p90_bit_slice_2061307_comb;
    p90_bit_slice_2061308 <= p90_bit_slice_2061308_comb;
    p90_bit_slice_2061309 <= p90_bit_slice_2061309_comb;
    p90_bit_slice_2061310 <= p90_bit_slice_2061310_comb;
    p90_bit_slice_2061311 <= p90_bit_slice_2061311_comb;
    p90_bit_slice_2061312 <= p90_bit_slice_2061312_comb;
    p90_array_index_2061313 <= p90_array_index_2061313_comb;
    p90_array_index_2061314 <= p90_array_index_2061314_comb;
    p90_array_index_2061315 <= p90_array_index_2061315_comb;
    p90_array_index_2061316 <= p90_array_index_2061316_comb;
    p90_array_index_2061317 <= p90_array_index_2061317_comb;
    p90_array_index_2061318 <= p90_array_index_2061318_comb;
    p90_bit_slice_2061319 <= p90_bit_slice_2061319_comb;
    p90_array_index_2061320 <= p90_array_index_2061320_comb;
    p90_bit_slice_2061321 <= p90_bit_slice_2061321_comb;
    p90_array_index_2061322 <= p90_array_index_2061322_comb;
    p90_array_index_2061323 <= p90_array_index_2061323_comb;
    p90_array_index_2061324 <= p90_array_index_2061324_comb;
    p90_array_index_2061325 <= p90_array_index_2061325_comb;
    p90_array_index_2061326 <= p90_array_index_2061326_comb;
    p90_array_index_2061327 <= p90_array_index_2061327_comb;
    p90_bit_slice_2061328 <= p90_bit_slice_2061328_comb;
    p91_literal_2043910 <= p90_literal_2043910;
    p91_literal_2043912 <= p90_literal_2043912;
    p91_literal_2043914 <= p90_literal_2043914;
    p91_literal_2043916 <= p90_literal_2043916;
    p91_literal_2043918 <= p90_literal_2043918;
    p91_literal_2043920 <= p90_literal_2043920;
    p91_literal_2043923 <= p90_literal_2043923;
  end

  // ===== Pipe stage 91:
  wire [7:0] p91_res7__1217_comb;
  wire [7:0] p91_array_index_2061417_comb;
  wire [7:0] p91_array_index_2061418_comb;
  wire [7:0] p91_array_index_2061419_comb;
  wire [7:0] p91_array_index_2061420_comb;
  wire [7:0] p91_array_index_2061421_comb;
  wire [7:0] p91_array_index_2061422_comb;
  wire [7:0] p91_res7__1219_comb;
  wire [7:0] p91_array_index_2061431_comb;
  wire [7:0] p91_array_index_2061432_comb;
  wire [7:0] p91_array_index_2061433_comb;
  wire [7:0] p91_array_index_2061434_comb;
  wire [7:0] p91_array_index_2061435_comb;
  wire [7:0] p91_res7__1221_comb;
  wire [7:0] p91_array_index_2061445_comb;
  wire [7:0] p91_array_index_2061446_comb;
  wire [7:0] p91_array_index_2061447_comb;
  wire [7:0] p91_array_index_2061448_comb;
  wire [7:0] p91_array_index_2061449_comb;
  wire [7:0] p91_res7__1223_comb;
  wire [7:0] p91_array_index_2061458_comb;
  wire [7:0] p91_array_index_2061459_comb;
  wire [7:0] p91_array_index_2061460_comb;
  wire [7:0] p91_array_index_2061461_comb;
  wire [7:0] p91_res7__1225_comb;
  wire [7:0] p91_array_index_2061471_comb;
  wire [7:0] p91_array_index_2061472_comb;
  wire [7:0] p91_array_index_2061473_comb;
  wire [7:0] p91_array_index_2061474_comb;
  wire [7:0] p91_res7__1227_comb;
  wire [7:0] p91_array_index_2061483_comb;
  wire [7:0] p91_array_index_2061484_comb;
  wire [7:0] p91_array_index_2061485_comb;
  wire [7:0] p91_res7__1229_comb;
  wire [7:0] p91_array_index_2061490_comb;
  wire [7:0] p91_array_index_2061491_comb;
  wire [7:0] p91_array_index_2061492_comb;
  wire [7:0] p91_array_index_2061493_comb;
  wire [7:0] p91_array_index_2061494_comb;
  wire [7:0] p91_array_index_2061495_comb;
  wire [7:0] p91_array_index_2061496_comb;
  wire [7:0] p91_array_index_2061497_comb;
  wire [7:0] p91_array_index_2061498_comb;
  wire [7:0] p91_array_index_2061499_comb;
  wire [7:0] p91_array_index_2061500_comb;
  assign p91_res7__1217_comb = p90_array_index_2061313 ^ p90_array_index_2061314 ^ p90_array_index_2061315 ^ p90_array_index_2061316 ^ p90_array_index_2061317 ^ p90_array_index_2061318 ^ p90_bit_slice_2061319 ^ p90_array_index_2061320 ^ p90_bit_slice_2061321 ^ p90_array_index_2061322 ^ p90_array_index_2061323 ^ p90_array_index_2061324 ^ p90_array_index_2061325 ^ p90_array_index_2061326 ^ p90_array_index_2061327 ^ p90_bit_slice_2061328;
  assign p91_array_index_2061417_comb = p90_literal_2043920[p90_bit_slice_2061308];
  assign p91_array_index_2061418_comb = p90_literal_2043918[p90_bit_slice_2061309];
  assign p91_array_index_2061419_comb = p90_literal_2043916[p90_bit_slice_2061310];
  assign p91_array_index_2061420_comb = p90_literal_2043914[p90_bit_slice_2061311];
  assign p91_array_index_2061421_comb = p90_literal_2043912[p90_bit_slice_2061312];
  assign p91_array_index_2061422_comb = p90_literal_2043910[p91_res7__1217_comb];
  assign p91_res7__1219_comb = p90_literal_2043910[p90_bit_slice_2061301] ^ p90_literal_2043912[p90_bit_slice_2061302] ^ p90_literal_2043914[p90_bit_slice_2061303] ^ p90_literal_2043916[p90_bit_slice_2061304] ^ p90_literal_2043918[p90_bit_slice_2061305] ^ p90_literal_2043920[p90_bit_slice_2061319] ^ p90_bit_slice_2061306 ^ p90_literal_2043923[p90_bit_slice_2061321] ^ p90_bit_slice_2061307 ^ p91_array_index_2061417_comb ^ p91_array_index_2061418_comb ^ p91_array_index_2061419_comb ^ p91_array_index_2061420_comb ^ p91_array_index_2061421_comb ^ p91_array_index_2061422_comb ^ p90_bit_slice_2061300;
  assign p91_array_index_2061431_comb = p90_literal_2043920[p90_bit_slice_2061309];
  assign p91_array_index_2061432_comb = p90_literal_2043918[p90_bit_slice_2061310];
  assign p91_array_index_2061433_comb = p90_literal_2043916[p90_bit_slice_2061311];
  assign p91_array_index_2061434_comb = p90_literal_2043914[p90_bit_slice_2061312];
  assign p91_array_index_2061435_comb = p90_literal_2043912[p91_res7__1217_comb];
  assign p91_res7__1221_comb = p90_literal_2043910[p90_bit_slice_2061302] ^ p90_literal_2043912[p90_bit_slice_2061303] ^ p90_literal_2043914[p90_bit_slice_2061304] ^ p90_literal_2043916[p90_bit_slice_2061305] ^ p90_literal_2043918[p90_bit_slice_2061319] ^ p90_literal_2043920[p90_bit_slice_2061306] ^ p90_bit_slice_2061321 ^ p90_literal_2043923[p90_bit_slice_2061307] ^ p90_bit_slice_2061308 ^ p91_array_index_2061431_comb ^ p91_array_index_2061432_comb ^ p91_array_index_2061433_comb ^ p91_array_index_2061434_comb ^ p91_array_index_2061435_comb ^ p90_literal_2043910[p91_res7__1219_comb] ^ p90_bit_slice_2061301;
  assign p91_array_index_2061445_comb = p90_literal_2043920[p90_bit_slice_2061310];
  assign p91_array_index_2061446_comb = p90_literal_2043918[p90_bit_slice_2061311];
  assign p91_array_index_2061447_comb = p90_literal_2043916[p90_bit_slice_2061312];
  assign p91_array_index_2061448_comb = p90_literal_2043914[p91_res7__1217_comb];
  assign p91_array_index_2061449_comb = p90_literal_2043912[p91_res7__1219_comb];
  assign p91_res7__1223_comb = p90_literal_2043910[p90_bit_slice_2061303] ^ p90_literal_2043912[p90_bit_slice_2061304] ^ p90_literal_2043914[p90_bit_slice_2061305] ^ p90_literal_2043916[p90_bit_slice_2061319] ^ p90_literal_2043918[p90_bit_slice_2061306] ^ p90_literal_2043920[p90_bit_slice_2061321] ^ p90_bit_slice_2061307 ^ p90_literal_2043923[p90_bit_slice_2061308] ^ p90_bit_slice_2061309 ^ p91_array_index_2061445_comb ^ p91_array_index_2061446_comb ^ p91_array_index_2061447_comb ^ p91_array_index_2061448_comb ^ p91_array_index_2061449_comb ^ p90_literal_2043910[p91_res7__1221_comb] ^ p90_bit_slice_2061302;
  assign p91_array_index_2061458_comb = p90_literal_2043920[p90_bit_slice_2061311];
  assign p91_array_index_2061459_comb = p90_literal_2043918[p90_bit_slice_2061312];
  assign p91_array_index_2061460_comb = p90_literal_2043916[p91_res7__1217_comb];
  assign p91_array_index_2061461_comb = p90_literal_2043914[p91_res7__1219_comb];
  assign p91_res7__1225_comb = p90_literal_2043910[p90_bit_slice_2061304] ^ p90_literal_2043912[p90_bit_slice_2061305] ^ p90_literal_2043914[p90_bit_slice_2061319] ^ p90_literal_2043916[p90_bit_slice_2061306] ^ p90_literal_2043918[p90_bit_slice_2061321] ^ p90_array_index_2061322 ^ p90_bit_slice_2061308 ^ p90_literal_2043923[p90_bit_slice_2061309] ^ p90_bit_slice_2061310 ^ p91_array_index_2061458_comb ^ p91_array_index_2061459_comb ^ p91_array_index_2061460_comb ^ p91_array_index_2061461_comb ^ p90_literal_2043912[p91_res7__1221_comb] ^ p90_literal_2043910[p91_res7__1223_comb] ^ p90_bit_slice_2061303;
  assign p91_array_index_2061471_comb = p90_literal_2043920[p90_bit_slice_2061312];
  assign p91_array_index_2061472_comb = p90_literal_2043918[p91_res7__1217_comb];
  assign p91_array_index_2061473_comb = p90_literal_2043916[p91_res7__1219_comb];
  assign p91_array_index_2061474_comb = p90_literal_2043914[p91_res7__1221_comb];
  assign p91_res7__1227_comb = p90_literal_2043910[p90_bit_slice_2061305] ^ p90_literal_2043912[p90_bit_slice_2061319] ^ p90_literal_2043914[p90_bit_slice_2061306] ^ p90_literal_2043916[p90_bit_slice_2061321] ^ p90_literal_2043918[p90_bit_slice_2061307] ^ p91_array_index_2061417_comb ^ p90_bit_slice_2061309 ^ p90_literal_2043923[p90_bit_slice_2061310] ^ p90_bit_slice_2061311 ^ p91_array_index_2061471_comb ^ p91_array_index_2061472_comb ^ p91_array_index_2061473_comb ^ p91_array_index_2061474_comb ^ p90_literal_2043912[p91_res7__1223_comb] ^ p90_literal_2043910[p91_res7__1225_comb] ^ p90_bit_slice_2061304;
  assign p91_array_index_2061483_comb = p90_literal_2043920[p91_res7__1217_comb];
  assign p91_array_index_2061484_comb = p90_literal_2043918[p91_res7__1219_comb];
  assign p91_array_index_2061485_comb = p90_literal_2043916[p91_res7__1221_comb];
  assign p91_res7__1229_comb = p90_literal_2043910[p90_bit_slice_2061319] ^ p90_literal_2043912[p90_bit_slice_2061306] ^ p90_literal_2043914[p90_bit_slice_2061321] ^ p90_literal_2043916[p90_bit_slice_2061307] ^ p90_array_index_2061323 ^ p91_array_index_2061431_comb ^ p90_bit_slice_2061310 ^ p90_literal_2043923[p90_bit_slice_2061311] ^ p90_bit_slice_2061312 ^ p91_array_index_2061483_comb ^ p91_array_index_2061484_comb ^ p91_array_index_2061485_comb ^ p90_literal_2043914[p91_res7__1223_comb] ^ p90_literal_2043912[p91_res7__1225_comb] ^ p90_literal_2043910[p91_res7__1227_comb] ^ p90_bit_slice_2061305;
  assign p91_array_index_2061490_comb = p90_literal_2043910[p90_bit_slice_2061306];
  assign p91_array_index_2061491_comb = p90_literal_2043912[p90_bit_slice_2061321];
  assign p91_array_index_2061492_comb = p90_literal_2043914[p90_bit_slice_2061307];
  assign p91_array_index_2061493_comb = p90_literal_2043916[p90_bit_slice_2061308];
  assign p91_array_index_2061494_comb = p90_literal_2043923[p90_bit_slice_2061312];
  assign p91_array_index_2061495_comb = p90_literal_2043920[p91_res7__1219_comb];
  assign p91_array_index_2061496_comb = p90_literal_2043918[p91_res7__1221_comb];
  assign p91_array_index_2061497_comb = p90_literal_2043916[p91_res7__1223_comb];
  assign p91_array_index_2061498_comb = p90_literal_2043914[p91_res7__1225_comb];
  assign p91_array_index_2061499_comb = p90_literal_2043912[p91_res7__1227_comb];
  assign p91_array_index_2061500_comb = p90_literal_2043910[p91_res7__1229_comb];

  // Registers for pipe stage 91:
  reg [127:0] p91_bit_slice_2043893;
  reg [127:0] p91_bit_slice_2044018;
  reg [127:0] p91_k2;
  reg [7:0] p91_bit_slice_2061306;
  reg [7:0] p91_bit_slice_2061307;
  reg [7:0] p91_bit_slice_2061308;
  reg [7:0] p91_bit_slice_2061309;
  reg [7:0] p91_bit_slice_2061310;
  reg [7:0] p91_bit_slice_2061311;
  reg [7:0] p91_bit_slice_2061312;
  reg [7:0] p91_bit_slice_2061319;
  reg [7:0] p91_bit_slice_2061321;
  reg [7:0] p91_array_index_2061324;
  reg [7:0] p91_array_index_2061325;
  reg [7:0] p91_array_index_2061326;
  reg [7:0] p91_array_index_2061327;
  reg [7:0] p91_res7__1217;
  reg [7:0] p91_array_index_2061418;
  reg [7:0] p91_array_index_2061419;
  reg [7:0] p91_array_index_2061420;
  reg [7:0] p91_array_index_2061421;
  reg [7:0] p91_array_index_2061422;
  reg [7:0] p91_res7__1219;
  reg [7:0] p91_array_index_2061432;
  reg [7:0] p91_array_index_2061433;
  reg [7:0] p91_array_index_2061434;
  reg [7:0] p91_array_index_2061435;
  reg [7:0] p91_res7__1221;
  reg [7:0] p91_array_index_2061445;
  reg [7:0] p91_array_index_2061446;
  reg [7:0] p91_array_index_2061447;
  reg [7:0] p91_array_index_2061448;
  reg [7:0] p91_array_index_2061449;
  reg [7:0] p91_res7__1223;
  reg [7:0] p91_array_index_2061458;
  reg [7:0] p91_array_index_2061459;
  reg [7:0] p91_array_index_2061460;
  reg [7:0] p91_array_index_2061461;
  reg [7:0] p91_res7__1225;
  reg [7:0] p91_array_index_2061471;
  reg [7:0] p91_array_index_2061472;
  reg [7:0] p91_array_index_2061473;
  reg [7:0] p91_array_index_2061474;
  reg [7:0] p91_res7__1227;
  reg [7:0] p91_array_index_2061483;
  reg [7:0] p91_array_index_2061484;
  reg [7:0] p91_array_index_2061485;
  reg [7:0] p91_res7__1229;
  reg [7:0] p91_array_index_2061490;
  reg [7:0] p91_array_index_2061491;
  reg [7:0] p91_array_index_2061492;
  reg [7:0] p91_array_index_2061493;
  reg [7:0] p91_array_index_2061494;
  reg [7:0] p91_array_index_2061495;
  reg [7:0] p91_array_index_2061496;
  reg [7:0] p91_array_index_2061497;
  reg [7:0] p91_array_index_2061498;
  reg [7:0] p91_array_index_2061499;
  reg [7:0] p91_array_index_2061500;
  reg [7:0] p92_literal_2043910[256];
  reg [7:0] p92_literal_2043912[256];
  reg [7:0] p92_literal_2043914[256];
  reg [7:0] p92_literal_2043916[256];
  reg [7:0] p92_literal_2043918[256];
  reg [7:0] p92_literal_2043920[256];
  reg [7:0] p92_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p91_bit_slice_2043893 <= p90_bit_slice_2043893;
    p91_bit_slice_2044018 <= p90_bit_slice_2044018;
    p91_k2 <= p90_k2;
    p91_bit_slice_2061306 <= p90_bit_slice_2061306;
    p91_bit_slice_2061307 <= p90_bit_slice_2061307;
    p91_bit_slice_2061308 <= p90_bit_slice_2061308;
    p91_bit_slice_2061309 <= p90_bit_slice_2061309;
    p91_bit_slice_2061310 <= p90_bit_slice_2061310;
    p91_bit_slice_2061311 <= p90_bit_slice_2061311;
    p91_bit_slice_2061312 <= p90_bit_slice_2061312;
    p91_bit_slice_2061319 <= p90_bit_slice_2061319;
    p91_bit_slice_2061321 <= p90_bit_slice_2061321;
    p91_array_index_2061324 <= p90_array_index_2061324;
    p91_array_index_2061325 <= p90_array_index_2061325;
    p91_array_index_2061326 <= p90_array_index_2061326;
    p91_array_index_2061327 <= p90_array_index_2061327;
    p91_res7__1217 <= p91_res7__1217_comb;
    p91_array_index_2061418 <= p91_array_index_2061418_comb;
    p91_array_index_2061419 <= p91_array_index_2061419_comb;
    p91_array_index_2061420 <= p91_array_index_2061420_comb;
    p91_array_index_2061421 <= p91_array_index_2061421_comb;
    p91_array_index_2061422 <= p91_array_index_2061422_comb;
    p91_res7__1219 <= p91_res7__1219_comb;
    p91_array_index_2061432 <= p91_array_index_2061432_comb;
    p91_array_index_2061433 <= p91_array_index_2061433_comb;
    p91_array_index_2061434 <= p91_array_index_2061434_comb;
    p91_array_index_2061435 <= p91_array_index_2061435_comb;
    p91_res7__1221 <= p91_res7__1221_comb;
    p91_array_index_2061445 <= p91_array_index_2061445_comb;
    p91_array_index_2061446 <= p91_array_index_2061446_comb;
    p91_array_index_2061447 <= p91_array_index_2061447_comb;
    p91_array_index_2061448 <= p91_array_index_2061448_comb;
    p91_array_index_2061449 <= p91_array_index_2061449_comb;
    p91_res7__1223 <= p91_res7__1223_comb;
    p91_array_index_2061458 <= p91_array_index_2061458_comb;
    p91_array_index_2061459 <= p91_array_index_2061459_comb;
    p91_array_index_2061460 <= p91_array_index_2061460_comb;
    p91_array_index_2061461 <= p91_array_index_2061461_comb;
    p91_res7__1225 <= p91_res7__1225_comb;
    p91_array_index_2061471 <= p91_array_index_2061471_comb;
    p91_array_index_2061472 <= p91_array_index_2061472_comb;
    p91_array_index_2061473 <= p91_array_index_2061473_comb;
    p91_array_index_2061474 <= p91_array_index_2061474_comb;
    p91_res7__1227 <= p91_res7__1227_comb;
    p91_array_index_2061483 <= p91_array_index_2061483_comb;
    p91_array_index_2061484 <= p91_array_index_2061484_comb;
    p91_array_index_2061485 <= p91_array_index_2061485_comb;
    p91_res7__1229 <= p91_res7__1229_comb;
    p91_array_index_2061490 <= p91_array_index_2061490_comb;
    p91_array_index_2061491 <= p91_array_index_2061491_comb;
    p91_array_index_2061492 <= p91_array_index_2061492_comb;
    p91_array_index_2061493 <= p91_array_index_2061493_comb;
    p91_array_index_2061494 <= p91_array_index_2061494_comb;
    p91_array_index_2061495 <= p91_array_index_2061495_comb;
    p91_array_index_2061496 <= p91_array_index_2061496_comb;
    p91_array_index_2061497 <= p91_array_index_2061497_comb;
    p91_array_index_2061498 <= p91_array_index_2061498_comb;
    p91_array_index_2061499 <= p91_array_index_2061499_comb;
    p91_array_index_2061500 <= p91_array_index_2061500_comb;
    p92_literal_2043910 <= p91_literal_2043910;
    p92_literal_2043912 <= p91_literal_2043912;
    p92_literal_2043914 <= p91_literal_2043914;
    p92_literal_2043916 <= p91_literal_2043916;
    p92_literal_2043918 <= p91_literal_2043918;
    p92_literal_2043920 <= p91_literal_2043920;
    p92_literal_2043923 <= p91_literal_2043923;
  end

  // ===== Pipe stage 92:
  wire [7:0] p92_res7__1231_comb;
  wire [7:0] p92_array_index_2061640_comb;
  wire [7:0] p92_array_index_2061641_comb;
  wire [7:0] p92_res7__1233_comb;
  wire [7:0] p92_array_index_2061651_comb;
  wire [7:0] p92_array_index_2061652_comb;
  wire [7:0] p92_res7__1235_comb;
  wire [7:0] p92_array_index_2061661_comb;
  wire [7:0] p92_res7__1237_comb;
  wire [7:0] p92_array_index_2061671_comb;
  wire [7:0] p92_res7__1239_comb;
  wire [7:0] p92_res7__1241_comb;
  wire [7:0] p92_res7__1243_comb;
  wire [7:0] p92_array_index_2061696_comb;
  wire [7:0] p92_array_index_2061697_comb;
  wire [7:0] p92_array_index_2061698_comb;
  wire [7:0] p92_array_index_2061699_comb;
  wire [7:0] p92_array_index_2061700_comb;
  wire [7:0] p92_array_index_2061701_comb;
  wire [7:0] p92_array_index_2061702_comb;
  wire [7:0] p92_array_index_2061703_comb;
  wire [7:0] p92_array_index_2061704_comb;
  wire [7:0] p92_array_index_2061705_comb;
  wire [7:0] p92_array_index_2061706_comb;
  wire [7:0] p92_array_index_2061707_comb;
  assign p92_res7__1231_comb = p91_array_index_2061490 ^ p91_array_index_2061491 ^ p91_array_index_2061492 ^ p91_array_index_2061493 ^ p91_array_index_2061418 ^ p91_array_index_2061445 ^ p91_bit_slice_2061311 ^ p91_array_index_2061494 ^ p91_res7__1217 ^ p91_array_index_2061495 ^ p91_array_index_2061496 ^ p91_array_index_2061497 ^ p91_array_index_2061498 ^ p91_array_index_2061499 ^ p91_array_index_2061500 ^ p91_bit_slice_2061319;
  assign p92_array_index_2061640_comb = p91_literal_2043920[p91_res7__1221];
  assign p92_array_index_2061641_comb = p91_literal_2043918[p91_res7__1223];
  assign p92_res7__1233_comb = p91_literal_2043910[p91_bit_slice_2061321] ^ p91_literal_2043912[p91_bit_slice_2061307] ^ p91_literal_2043914[p91_bit_slice_2061308] ^ p91_array_index_2061324 ^ p91_array_index_2061432 ^ p91_array_index_2061458 ^ p91_bit_slice_2061312 ^ p91_literal_2043923[p91_res7__1217] ^ p91_res7__1219 ^ p92_array_index_2061640_comb ^ p92_array_index_2061641_comb ^ p91_literal_2043916[p91_res7__1225] ^ p91_literal_2043914[p91_res7__1227] ^ p91_literal_2043912[p91_res7__1229] ^ p91_literal_2043910[p92_res7__1231_comb] ^ p91_bit_slice_2061306;
  assign p92_array_index_2061651_comb = p91_literal_2043920[p91_res7__1223];
  assign p92_array_index_2061652_comb = p91_literal_2043918[p91_res7__1225];
  assign p92_res7__1235_comb = p91_literal_2043910[p91_bit_slice_2061307] ^ p91_literal_2043912[p91_bit_slice_2061308] ^ p91_literal_2043914[p91_bit_slice_2061309] ^ p91_array_index_2061419 ^ p91_array_index_2061446 ^ p91_array_index_2061471 ^ p91_res7__1217 ^ p91_literal_2043923[p91_res7__1219] ^ p91_res7__1221 ^ p92_array_index_2061651_comb ^ p92_array_index_2061652_comb ^ p91_literal_2043916[p91_res7__1227] ^ p91_literal_2043914[p91_res7__1229] ^ p91_literal_2043912[p92_res7__1231_comb] ^ p91_literal_2043910[p92_res7__1233_comb] ^ p91_bit_slice_2061321;
  assign p92_array_index_2061661_comb = p91_literal_2043920[p91_res7__1225];
  assign p92_res7__1237_comb = p91_literal_2043910[p91_bit_slice_2061308] ^ p91_literal_2043912[p91_bit_slice_2061309] ^ p91_array_index_2061325 ^ p91_array_index_2061433 ^ p91_array_index_2061459 ^ p91_array_index_2061483 ^ p91_res7__1219 ^ p91_literal_2043923[p91_res7__1221] ^ p91_res7__1223 ^ p92_array_index_2061661_comb ^ p91_literal_2043918[p91_res7__1227] ^ p91_literal_2043916[p91_res7__1229] ^ p91_literal_2043914[p92_res7__1231_comb] ^ p91_literal_2043912[p92_res7__1233_comb] ^ p91_literal_2043910[p92_res7__1235_comb] ^ p91_bit_slice_2061307;
  assign p92_array_index_2061671_comb = p91_literal_2043920[p91_res7__1227];
  assign p92_res7__1239_comb = p91_literal_2043910[p91_bit_slice_2061309] ^ p91_literal_2043912[p91_bit_slice_2061310] ^ p91_array_index_2061420 ^ p91_array_index_2061447 ^ p91_array_index_2061472 ^ p91_array_index_2061495 ^ p91_res7__1221 ^ p91_literal_2043923[p91_res7__1223] ^ p91_res7__1225 ^ p92_array_index_2061671_comb ^ p91_literal_2043918[p91_res7__1229] ^ p91_literal_2043916[p92_res7__1231_comb] ^ p91_literal_2043914[p92_res7__1233_comb] ^ p91_literal_2043912[p92_res7__1235_comb] ^ p91_literal_2043910[p92_res7__1237_comb] ^ p91_bit_slice_2061308;
  assign p92_res7__1241_comb = p91_literal_2043910[p91_bit_slice_2061310] ^ p91_array_index_2061326 ^ p91_array_index_2061434 ^ p91_array_index_2061460 ^ p91_array_index_2061484 ^ p92_array_index_2061640_comb ^ p91_res7__1223 ^ p91_literal_2043923[p91_res7__1225] ^ p91_res7__1227 ^ p91_literal_2043920[p91_res7__1229] ^ p91_literal_2043918[p92_res7__1231_comb] ^ p91_literal_2043916[p92_res7__1233_comb] ^ p91_literal_2043914[p92_res7__1235_comb] ^ p91_literal_2043912[p92_res7__1237_comb] ^ p91_literal_2043910[p92_res7__1239_comb] ^ p91_bit_slice_2061309;
  assign p92_res7__1243_comb = p91_literal_2043910[p91_bit_slice_2061311] ^ p91_array_index_2061421 ^ p91_array_index_2061448 ^ p91_array_index_2061473 ^ p91_array_index_2061496 ^ p92_array_index_2061651_comb ^ p91_res7__1225 ^ p91_literal_2043923[p91_res7__1227] ^ p91_res7__1229 ^ p91_literal_2043920[p92_res7__1231_comb] ^ p91_literal_2043918[p92_res7__1233_comb] ^ p91_literal_2043916[p92_res7__1235_comb] ^ p91_literal_2043914[p92_res7__1237_comb] ^ p91_literal_2043912[p92_res7__1239_comb] ^ p91_literal_2043910[p92_res7__1241_comb] ^ p91_bit_slice_2061310;
  assign p92_array_index_2061696_comb = p91_literal_2043923[p91_res7__1229];
  assign p92_array_index_2061697_comb = p91_literal_2043920[p92_res7__1233_comb];
  assign p92_array_index_2061698_comb = p91_literal_2043918[p92_res7__1235_comb];
  assign p92_array_index_2061699_comb = p91_literal_2043916[p92_res7__1237_comb];
  assign p92_array_index_2061700_comb = p91_literal_2043914[p92_res7__1239_comb];
  assign p92_array_index_2061701_comb = p91_literal_2043912[p92_res7__1241_comb];
  assign p92_array_index_2061702_comb = p91_literal_2043910[p92_res7__1243_comb];
  assign p92_array_index_2061703_comb = p91_literal_2058836[p91_res7__1217];
  assign p92_array_index_2061704_comb = p91_literal_2058836[p91_res7__1219];
  assign p92_array_index_2061705_comb = p91_literal_2058836[p91_res7__1221];
  assign p92_array_index_2061706_comb = p91_literal_2058836[p91_res7__1223];
  assign p92_array_index_2061707_comb = p91_literal_2058836[p91_res7__1225];

  // Registers for pipe stage 92:
  reg [127:0] p92_bit_slice_2043893;
  reg [127:0] p92_bit_slice_2044018;
  reg [127:0] p92_k2;
  reg [7:0] p92_bit_slice_2061311;
  reg [7:0] p92_bit_slice_2061312;
  reg [7:0] p92_array_index_2061327;
  reg [7:0] p92_array_index_2061422;
  reg [7:0] p92_array_index_2061435;
  reg [7:0] p92_array_index_2061449;
  reg [7:0] p92_array_index_2061461;
  reg [7:0] p92_array_index_2061474;
  reg [7:0] p92_res7__1227;
  reg [7:0] p92_array_index_2061485;
  reg [7:0] p92_res7__1229;
  reg [7:0] p92_array_index_2061497;
  reg [7:0] p92_res7__1231;
  reg [7:0] p92_array_index_2061641;
  reg [7:0] p92_res7__1233;
  reg [7:0] p92_array_index_2061652;
  reg [7:0] p92_res7__1235;
  reg [7:0] p92_array_index_2061661;
  reg [7:0] p92_res7__1237;
  reg [7:0] p92_array_index_2061671;
  reg [7:0] p92_res7__1239;
  reg [7:0] p92_res7__1241;
  reg [7:0] p92_res7__1243;
  reg [7:0] p92_array_index_2061696;
  reg [7:0] p92_array_index_2061697;
  reg [7:0] p92_array_index_2061698;
  reg [7:0] p92_array_index_2061699;
  reg [7:0] p92_array_index_2061700;
  reg [7:0] p92_array_index_2061701;
  reg [7:0] p92_array_index_2061702;
  reg [7:0] p92_array_index_2061703;
  reg [7:0] p92_array_index_2061704;
  reg [7:0] p92_array_index_2061705;
  reg [7:0] p92_array_index_2061706;
  reg [7:0] p92_array_index_2061707;
  reg [7:0] p93_literal_2043910[256];
  reg [7:0] p93_literal_2043912[256];
  reg [7:0] p93_literal_2043914[256];
  reg [7:0] p93_literal_2043916[256];
  reg [7:0] p93_literal_2043918[256];
  reg [7:0] p93_literal_2043920[256];
  reg [7:0] p93_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p92_bit_slice_2043893 <= p91_bit_slice_2043893;
    p92_bit_slice_2044018 <= p91_bit_slice_2044018;
    p92_k2 <= p91_k2;
    p92_bit_slice_2061311 <= p91_bit_slice_2061311;
    p92_bit_slice_2061312 <= p91_bit_slice_2061312;
    p92_array_index_2061327 <= p91_array_index_2061327;
    p92_array_index_2061422 <= p91_array_index_2061422;
    p92_array_index_2061435 <= p91_array_index_2061435;
    p92_array_index_2061449 <= p91_array_index_2061449;
    p92_array_index_2061461 <= p91_array_index_2061461;
    p92_array_index_2061474 <= p91_array_index_2061474;
    p92_res7__1227 <= p91_res7__1227;
    p92_array_index_2061485 <= p91_array_index_2061485;
    p92_res7__1229 <= p91_res7__1229;
    p92_array_index_2061497 <= p91_array_index_2061497;
    p92_res7__1231 <= p92_res7__1231_comb;
    p92_array_index_2061641 <= p92_array_index_2061641_comb;
    p92_res7__1233 <= p92_res7__1233_comb;
    p92_array_index_2061652 <= p92_array_index_2061652_comb;
    p92_res7__1235 <= p92_res7__1235_comb;
    p92_array_index_2061661 <= p92_array_index_2061661_comb;
    p92_res7__1237 <= p92_res7__1237_comb;
    p92_array_index_2061671 <= p92_array_index_2061671_comb;
    p92_res7__1239 <= p92_res7__1239_comb;
    p92_res7__1241 <= p92_res7__1241_comb;
    p92_res7__1243 <= p92_res7__1243_comb;
    p92_array_index_2061696 <= p92_array_index_2061696_comb;
    p92_array_index_2061697 <= p92_array_index_2061697_comb;
    p92_array_index_2061698 <= p92_array_index_2061698_comb;
    p92_array_index_2061699 <= p92_array_index_2061699_comb;
    p92_array_index_2061700 <= p92_array_index_2061700_comb;
    p92_array_index_2061701 <= p92_array_index_2061701_comb;
    p92_array_index_2061702 <= p92_array_index_2061702_comb;
    p92_array_index_2061703 <= p92_array_index_2061703_comb;
    p92_array_index_2061704 <= p92_array_index_2061704_comb;
    p92_array_index_2061705 <= p92_array_index_2061705_comb;
    p92_array_index_2061706 <= p92_array_index_2061706_comb;
    p92_array_index_2061707 <= p92_array_index_2061707_comb;
    p93_literal_2043910 <= p92_literal_2043910;
    p93_literal_2043912 <= p92_literal_2043912;
    p93_literal_2043914 <= p92_literal_2043914;
    p93_literal_2043916 <= p92_literal_2043916;
    p93_literal_2043918 <= p92_literal_2043918;
    p93_literal_2043920 <= p92_literal_2043920;
    p93_literal_2043923 <= p92_literal_2043923;
  end

  // ===== Pipe stage 93:
  wire [7:0] p93_res7__1245_comb;
  wire [7:0] p93_res7__1247_comb;
  wire [127:0] p93_permut__38_comb;
  wire [127:0] p93_xor_2061821_comb;
  wire [7:0] p93_bit_slice_2061825_comb;
  wire [7:0] p93_bit_slice_2061826_comb;
  wire [7:0] p93_bit_slice_2061827_comb;
  wire [7:0] p93_bit_slice_2061828_comb;
  wire [7:0] p93_bit_slice_2061829_comb;
  wire [7:0] p93_bit_slice_2061830_comb;
  wire [7:0] p93_bit_slice_2061831_comb;
  wire [7:0] p93_bit_slice_2061832_comb;
  wire [7:0] p93_bit_slice_2061833_comb;
  wire [7:0] p93_bit_slice_2061834_comb;
  wire [7:0] p93_bit_slice_2061841_comb;
  wire [7:0] p93_bit_slice_2061843_comb;
  wire [7:0] p93_array_index_2061844_comb;
  wire [7:0] p93_array_index_2061845_comb;
  wire [7:0] p93_array_index_2061846_comb;
  wire [7:0] p93_array_index_2061847_comb;
  wire [7:0] p93_array_index_2061848_comb;
  wire [7:0] p93_array_index_2061849_comb;
  wire [7:0] p93_res7__1249_comb;
  wire [7:0] p93_array_index_2061859_comb;
  wire [7:0] p93_array_index_2061860_comb;
  wire [7:0] p93_array_index_2061861_comb;
  wire [7:0] p93_array_index_2061862_comb;
  wire [7:0] p93_array_index_2061863_comb;
  wire [7:0] p93_array_index_2061864_comb;
  wire [7:0] p93_res7__1251_comb;
  wire [7:0] p93_array_index_2061873_comb;
  wire [7:0] p93_array_index_2061874_comb;
  wire [7:0] p93_array_index_2061875_comb;
  wire [7:0] p93_array_index_2061876_comb;
  wire [7:0] p93_array_index_2061877_comb;
  wire [7:0] p93_res7__1253_comb;
  wire [7:0] p93_array_index_2061887_comb;
  wire [7:0] p93_array_index_2061888_comb;
  wire [7:0] p93_array_index_2061889_comb;
  wire [7:0] p93_array_index_2061890_comb;
  wire [7:0] p93_array_index_2061891_comb;
  wire [7:0] p93_res7__1255_comb;
  wire [7:0] p93_array_index_2061894_comb;
  wire [7:0] p93_array_index_2061895_comb;
  wire [7:0] p93_array_index_2061896_comb;
  wire [7:0] p93_array_index_2061897_comb;
  wire [7:0] p93_array_index_2061898_comb;
  wire [7:0] p93_array_index_2061899_comb;
  wire [7:0] p93_array_index_2061900_comb;
  wire [7:0] p93_array_index_2061901_comb;
  wire [7:0] p93_array_index_2061902_comb;
  wire [7:0] p93_array_index_2061903_comb;
  wire [7:0] p93_array_index_2061904_comb;
  wire [7:0] p93_array_index_2061905_comb;
  assign p93_res7__1245_comb = p92_array_index_2061327 ^ p92_array_index_2061435 ^ p92_array_index_2061461 ^ p92_array_index_2061485 ^ p92_array_index_2061641 ^ p92_array_index_2061661 ^ p92_res7__1227 ^ p92_array_index_2061696 ^ p92_res7__1231 ^ p92_array_index_2061697 ^ p92_array_index_2061698 ^ p92_array_index_2061699 ^ p92_array_index_2061700 ^ p92_array_index_2061701 ^ p92_array_index_2061702 ^ p92_bit_slice_2061311;
  assign p93_res7__1247_comb = p92_array_index_2061422 ^ p92_array_index_2061449 ^ p92_array_index_2061474 ^ p92_array_index_2061497 ^ p92_array_index_2061652 ^ p92_array_index_2061671 ^ p92_res7__1229 ^ p92_literal_2043923[p92_res7__1231] ^ p92_res7__1233 ^ p92_literal_2043920[p92_res7__1235] ^ p92_literal_2043918[p92_res7__1237] ^ p92_literal_2043916[p92_res7__1239] ^ p92_literal_2043914[p92_res7__1241] ^ p92_literal_2043912[p92_res7__1243] ^ p92_literal_2043910[p93_res7__1245_comb] ^ p92_bit_slice_2061312;
  assign p93_permut__38_comb = {p92_array_index_2061703, p92_array_index_2061704, p92_array_index_2061705, p92_array_index_2061706, p92_array_index_2061707, p92_literal_2058836[p92_res7__1227], p92_literal_2058836[p92_res7__1229], p92_literal_2058836[p92_res7__1231], p92_literal_2058836[p92_res7__1233], p92_literal_2058836[p92_res7__1235], p92_literal_2058836[p92_res7__1237], p92_literal_2058836[p92_res7__1239], p92_literal_2058836[p92_res7__1241], p92_literal_2058836[p92_res7__1243], p92_literal_2058836[p93_res7__1245_comb], p92_literal_2058836[p93_res7__1247_comb]};
  assign p93_xor_2061821_comb = p92_k2 ^ p93_permut__38_comb;
  assign p93_bit_slice_2061825_comb = p93_xor_2061821_comb[95:88];
  assign p93_bit_slice_2061826_comb = p93_xor_2061821_comb[87:80];
  assign p93_bit_slice_2061827_comb = p93_xor_2061821_comb[79:72];
  assign p93_bit_slice_2061828_comb = p93_xor_2061821_comb[63:56];
  assign p93_bit_slice_2061829_comb = p93_xor_2061821_comb[47:40];
  assign p93_bit_slice_2061830_comb = p93_xor_2061821_comb[39:32];
  assign p93_bit_slice_2061831_comb = p93_xor_2061821_comb[31:24];
  assign p93_bit_slice_2061832_comb = p93_xor_2061821_comb[23:16];
  assign p93_bit_slice_2061833_comb = p93_xor_2061821_comb[15:8];
  assign p93_bit_slice_2061834_comb = p93_xor_2061821_comb[7:0];
  assign p93_bit_slice_2061841_comb = p93_xor_2061821_comb[71:64];
  assign p93_bit_slice_2061843_comb = p93_xor_2061821_comb[55:48];
  assign p93_array_index_2061844_comb = p92_literal_2043920[p93_bit_slice_2061829_comb];
  assign p93_array_index_2061845_comb = p92_literal_2043918[p93_bit_slice_2061830_comb];
  assign p93_array_index_2061846_comb = p92_literal_2043916[p93_bit_slice_2061831_comb];
  assign p93_array_index_2061847_comb = p92_literal_2043914[p93_bit_slice_2061832_comb];
  assign p93_array_index_2061848_comb = p92_literal_2043912[p93_bit_slice_2061833_comb];
  assign p93_array_index_2061849_comb = p92_literal_2043910[p93_bit_slice_2061834_comb];
  assign p93_res7__1249_comb = p92_literal_2043910[p93_xor_2061821_comb[119:112]] ^ p92_literal_2043912[p93_xor_2061821_comb[111:104]] ^ p92_literal_2043914[p93_xor_2061821_comb[103:96]] ^ p92_literal_2043916[p93_bit_slice_2061825_comb] ^ p92_literal_2043918[p93_bit_slice_2061826_comb] ^ p92_literal_2043920[p93_bit_slice_2061827_comb] ^ p93_bit_slice_2061841_comb ^ p92_literal_2043923[p93_bit_slice_2061828_comb] ^ p93_bit_slice_2061843_comb ^ p93_array_index_2061844_comb ^ p93_array_index_2061845_comb ^ p93_array_index_2061846_comb ^ p93_array_index_2061847_comb ^ p93_array_index_2061848_comb ^ p93_array_index_2061849_comb ^ p93_xor_2061821_comb[127:120];
  assign p93_array_index_2061859_comb = p92_literal_2043920[p93_bit_slice_2061830_comb];
  assign p93_array_index_2061860_comb = p92_literal_2043918[p93_bit_slice_2061831_comb];
  assign p93_array_index_2061861_comb = p92_literal_2043916[p93_bit_slice_2061832_comb];
  assign p93_array_index_2061862_comb = p92_literal_2043914[p93_bit_slice_2061833_comb];
  assign p93_array_index_2061863_comb = p92_literal_2043912[p93_bit_slice_2061834_comb];
  assign p93_array_index_2061864_comb = p92_literal_2043910[p93_res7__1249_comb];
  assign p93_res7__1251_comb = p92_literal_2043910[p93_xor_2061821_comb[111:104]] ^ p92_literal_2043912[p93_xor_2061821_comb[103:96]] ^ p92_literal_2043914[p93_bit_slice_2061825_comb] ^ p92_literal_2043916[p93_bit_slice_2061826_comb] ^ p92_literal_2043918[p93_bit_slice_2061827_comb] ^ p92_literal_2043920[p93_bit_slice_2061841_comb] ^ p93_bit_slice_2061828_comb ^ p92_literal_2043923[p93_bit_slice_2061843_comb] ^ p93_bit_slice_2061829_comb ^ p93_array_index_2061859_comb ^ p93_array_index_2061860_comb ^ p93_array_index_2061861_comb ^ p93_array_index_2061862_comb ^ p93_array_index_2061863_comb ^ p93_array_index_2061864_comb ^ p93_xor_2061821_comb[119:112];
  assign p93_array_index_2061873_comb = p92_literal_2043920[p93_bit_slice_2061831_comb];
  assign p93_array_index_2061874_comb = p92_literal_2043918[p93_bit_slice_2061832_comb];
  assign p93_array_index_2061875_comb = p92_literal_2043916[p93_bit_slice_2061833_comb];
  assign p93_array_index_2061876_comb = p92_literal_2043914[p93_bit_slice_2061834_comb];
  assign p93_array_index_2061877_comb = p92_literal_2043912[p93_res7__1249_comb];
  assign p93_res7__1253_comb = p92_literal_2043910[p93_xor_2061821_comb[103:96]] ^ p92_literal_2043912[p93_bit_slice_2061825_comb] ^ p92_literal_2043914[p93_bit_slice_2061826_comb] ^ p92_literal_2043916[p93_bit_slice_2061827_comb] ^ p92_literal_2043918[p93_bit_slice_2061841_comb] ^ p92_literal_2043920[p93_bit_slice_2061828_comb] ^ p93_bit_slice_2061843_comb ^ p92_literal_2043923[p93_bit_slice_2061829_comb] ^ p93_bit_slice_2061830_comb ^ p93_array_index_2061873_comb ^ p93_array_index_2061874_comb ^ p93_array_index_2061875_comb ^ p93_array_index_2061876_comb ^ p93_array_index_2061877_comb ^ p92_literal_2043910[p93_res7__1251_comb] ^ p93_xor_2061821_comb[111:104];
  assign p93_array_index_2061887_comb = p92_literal_2043920[p93_bit_slice_2061832_comb];
  assign p93_array_index_2061888_comb = p92_literal_2043918[p93_bit_slice_2061833_comb];
  assign p93_array_index_2061889_comb = p92_literal_2043916[p93_bit_slice_2061834_comb];
  assign p93_array_index_2061890_comb = p92_literal_2043914[p93_res7__1249_comb];
  assign p93_array_index_2061891_comb = p92_literal_2043912[p93_res7__1251_comb];
  assign p93_res7__1255_comb = p92_literal_2043910[p93_bit_slice_2061825_comb] ^ p92_literal_2043912[p93_bit_slice_2061826_comb] ^ p92_literal_2043914[p93_bit_slice_2061827_comb] ^ p92_literal_2043916[p93_bit_slice_2061841_comb] ^ p92_literal_2043918[p93_bit_slice_2061828_comb] ^ p92_literal_2043920[p93_bit_slice_2061843_comb] ^ p93_bit_slice_2061829_comb ^ p92_literal_2043923[p93_bit_slice_2061830_comb] ^ p93_bit_slice_2061831_comb ^ p93_array_index_2061887_comb ^ p93_array_index_2061888_comb ^ p93_array_index_2061889_comb ^ p93_array_index_2061890_comb ^ p93_array_index_2061891_comb ^ p92_literal_2043910[p93_res7__1253_comb] ^ p93_xor_2061821_comb[103:96];
  assign p93_array_index_2061894_comb = p92_literal_2043910[p93_bit_slice_2061826_comb];
  assign p93_array_index_2061895_comb = p92_literal_2043912[p93_bit_slice_2061827_comb];
  assign p93_array_index_2061896_comb = p92_literal_2043914[p93_bit_slice_2061841_comb];
  assign p93_array_index_2061897_comb = p92_literal_2043916[p93_bit_slice_2061828_comb];
  assign p93_array_index_2061898_comb = p92_literal_2043918[p93_bit_slice_2061843_comb];
  assign p93_array_index_2061899_comb = p92_literal_2043923[p93_bit_slice_2061831_comb];
  assign p93_array_index_2061900_comb = p92_literal_2043920[p93_bit_slice_2061833_comb];
  assign p93_array_index_2061901_comb = p92_literal_2043918[p93_bit_slice_2061834_comb];
  assign p93_array_index_2061902_comb = p92_literal_2043916[p93_res7__1249_comb];
  assign p93_array_index_2061903_comb = p92_literal_2043914[p93_res7__1251_comb];
  assign p93_array_index_2061904_comb = p92_literal_2043912[p93_res7__1253_comb];
  assign p93_array_index_2061905_comb = p92_literal_2043910[p93_res7__1255_comb];

  // Registers for pipe stage 93:
  reg [127:0] p93_bit_slice_2043893;
  reg [127:0] p93_bit_slice_2044018;
  reg [7:0] p93_bit_slice_2061825;
  reg [7:0] p93_bit_slice_2061826;
  reg [7:0] p93_bit_slice_2061827;
  reg [7:0] p93_bit_slice_2061828;
  reg [7:0] p93_bit_slice_2061829;
  reg [7:0] p93_bit_slice_2061830;
  reg [7:0] p93_bit_slice_2061831;
  reg [7:0] p93_bit_slice_2061832;
  reg [7:0] p93_bit_slice_2061833;
  reg [7:0] p93_bit_slice_2061834;
  reg [7:0] p93_bit_slice_2061841;
  reg [7:0] p93_bit_slice_2061843;
  reg [7:0] p93_array_index_2061844;
  reg [7:0] p93_array_index_2061845;
  reg [7:0] p93_array_index_2061846;
  reg [7:0] p93_array_index_2061847;
  reg [7:0] p93_array_index_2061848;
  reg [7:0] p93_array_index_2061849;
  reg [7:0] p93_res7__1249;
  reg [7:0] p93_array_index_2061859;
  reg [7:0] p93_array_index_2061860;
  reg [7:0] p93_array_index_2061861;
  reg [7:0] p93_array_index_2061862;
  reg [7:0] p93_array_index_2061863;
  reg [7:0] p93_array_index_2061864;
  reg [7:0] p93_res7__1251;
  reg [7:0] p93_array_index_2061873;
  reg [7:0] p93_array_index_2061874;
  reg [7:0] p93_array_index_2061875;
  reg [7:0] p93_array_index_2061876;
  reg [7:0] p93_array_index_2061877;
  reg [7:0] p93_res7__1253;
  reg [7:0] p93_array_index_2061887;
  reg [7:0] p93_array_index_2061888;
  reg [7:0] p93_array_index_2061889;
  reg [7:0] p93_array_index_2061890;
  reg [7:0] p93_array_index_2061891;
  reg [7:0] p93_res7__1255;
  reg [7:0] p93_array_index_2061894;
  reg [7:0] p93_array_index_2061895;
  reg [7:0] p93_array_index_2061896;
  reg [7:0] p93_array_index_2061897;
  reg [7:0] p93_array_index_2061898;
  reg [7:0] p93_array_index_2061899;
  reg [7:0] p93_array_index_2061900;
  reg [7:0] p93_array_index_2061901;
  reg [7:0] p93_array_index_2061902;
  reg [7:0] p93_array_index_2061903;
  reg [7:0] p93_array_index_2061904;
  reg [7:0] p93_array_index_2061905;
  reg [7:0] p94_literal_2043910[256];
  reg [7:0] p94_literal_2043912[256];
  reg [7:0] p94_literal_2043914[256];
  reg [7:0] p94_literal_2043916[256];
  reg [7:0] p94_literal_2043918[256];
  reg [7:0] p94_literal_2043920[256];
  reg [7:0] p94_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p93_bit_slice_2043893 <= p92_bit_slice_2043893;
    p93_bit_slice_2044018 <= p92_bit_slice_2044018;
    p93_bit_slice_2061825 <= p93_bit_slice_2061825_comb;
    p93_bit_slice_2061826 <= p93_bit_slice_2061826_comb;
    p93_bit_slice_2061827 <= p93_bit_slice_2061827_comb;
    p93_bit_slice_2061828 <= p93_bit_slice_2061828_comb;
    p93_bit_slice_2061829 <= p93_bit_slice_2061829_comb;
    p93_bit_slice_2061830 <= p93_bit_slice_2061830_comb;
    p93_bit_slice_2061831 <= p93_bit_slice_2061831_comb;
    p93_bit_slice_2061832 <= p93_bit_slice_2061832_comb;
    p93_bit_slice_2061833 <= p93_bit_slice_2061833_comb;
    p93_bit_slice_2061834 <= p93_bit_slice_2061834_comb;
    p93_bit_slice_2061841 <= p93_bit_slice_2061841_comb;
    p93_bit_slice_2061843 <= p93_bit_slice_2061843_comb;
    p93_array_index_2061844 <= p93_array_index_2061844_comb;
    p93_array_index_2061845 <= p93_array_index_2061845_comb;
    p93_array_index_2061846 <= p93_array_index_2061846_comb;
    p93_array_index_2061847 <= p93_array_index_2061847_comb;
    p93_array_index_2061848 <= p93_array_index_2061848_comb;
    p93_array_index_2061849 <= p93_array_index_2061849_comb;
    p93_res7__1249 <= p93_res7__1249_comb;
    p93_array_index_2061859 <= p93_array_index_2061859_comb;
    p93_array_index_2061860 <= p93_array_index_2061860_comb;
    p93_array_index_2061861 <= p93_array_index_2061861_comb;
    p93_array_index_2061862 <= p93_array_index_2061862_comb;
    p93_array_index_2061863 <= p93_array_index_2061863_comb;
    p93_array_index_2061864 <= p93_array_index_2061864_comb;
    p93_res7__1251 <= p93_res7__1251_comb;
    p93_array_index_2061873 <= p93_array_index_2061873_comb;
    p93_array_index_2061874 <= p93_array_index_2061874_comb;
    p93_array_index_2061875 <= p93_array_index_2061875_comb;
    p93_array_index_2061876 <= p93_array_index_2061876_comb;
    p93_array_index_2061877 <= p93_array_index_2061877_comb;
    p93_res7__1253 <= p93_res7__1253_comb;
    p93_array_index_2061887 <= p93_array_index_2061887_comb;
    p93_array_index_2061888 <= p93_array_index_2061888_comb;
    p93_array_index_2061889 <= p93_array_index_2061889_comb;
    p93_array_index_2061890 <= p93_array_index_2061890_comb;
    p93_array_index_2061891 <= p93_array_index_2061891_comb;
    p93_res7__1255 <= p93_res7__1255_comb;
    p93_array_index_2061894 <= p93_array_index_2061894_comb;
    p93_array_index_2061895 <= p93_array_index_2061895_comb;
    p93_array_index_2061896 <= p93_array_index_2061896_comb;
    p93_array_index_2061897 <= p93_array_index_2061897_comb;
    p93_array_index_2061898 <= p93_array_index_2061898_comb;
    p93_array_index_2061899 <= p93_array_index_2061899_comb;
    p93_array_index_2061900 <= p93_array_index_2061900_comb;
    p93_array_index_2061901 <= p93_array_index_2061901_comb;
    p93_array_index_2061902 <= p93_array_index_2061902_comb;
    p93_array_index_2061903 <= p93_array_index_2061903_comb;
    p93_array_index_2061904 <= p93_array_index_2061904_comb;
    p93_array_index_2061905 <= p93_array_index_2061905_comb;
    p94_literal_2043910 <= p93_literal_2043910;
    p94_literal_2043912 <= p93_literal_2043912;
    p94_literal_2043914 <= p93_literal_2043914;
    p94_literal_2043916 <= p93_literal_2043916;
    p94_literal_2043918 <= p93_literal_2043918;
    p94_literal_2043920 <= p93_literal_2043920;
    p94_literal_2043923 <= p93_literal_2043923;
  end

  // ===== Pipe stage 94:
  wire [7:0] p94_res7__1257_comb;
  wire [7:0] p94_array_index_2062033_comb;
  wire [7:0] p94_array_index_2062034_comb;
  wire [7:0] p94_array_index_2062035_comb;
  wire [7:0] p94_array_index_2062036_comb;
  wire [7:0] p94_res7__1259_comb;
  wire [7:0] p94_array_index_2062045_comb;
  wire [7:0] p94_array_index_2062046_comb;
  wire [7:0] p94_array_index_2062047_comb;
  wire [7:0] p94_res7__1261_comb;
  wire [7:0] p94_array_index_2062057_comb;
  wire [7:0] p94_array_index_2062058_comb;
  wire [7:0] p94_array_index_2062059_comb;
  wire [7:0] p94_res7__1263_comb;
  wire [7:0] p94_array_index_2062068_comb;
  wire [7:0] p94_array_index_2062069_comb;
  wire [7:0] p94_res7__1265_comb;
  wire [7:0] p94_array_index_2062079_comb;
  wire [7:0] p94_array_index_2062080_comb;
  wire [7:0] p94_res7__1267_comb;
  wire [7:0] p94_array_index_2062089_comb;
  wire [7:0] p94_res7__1269_comb;
  wire [7:0] p94_array_index_2062096_comb;
  wire [7:0] p94_array_index_2062097_comb;
  wire [7:0] p94_array_index_2062098_comb;
  wire [7:0] p94_array_index_2062099_comb;
  wire [7:0] p94_array_index_2062100_comb;
  wire [7:0] p94_array_index_2062101_comb;
  wire [7:0] p94_array_index_2062102_comb;
  wire [7:0] p94_array_index_2062103_comb;
  wire [7:0] p94_array_index_2062104_comb;
  wire [7:0] p94_array_index_2062105_comb;
  wire [7:0] p94_array_index_2062106_comb;
  assign p94_res7__1257_comb = p93_array_index_2061894 ^ p93_array_index_2061895 ^ p93_array_index_2061896 ^ p93_array_index_2061897 ^ p93_array_index_2061898 ^ p93_array_index_2061844 ^ p93_bit_slice_2061830 ^ p93_array_index_2061899 ^ p93_bit_slice_2061832 ^ p93_array_index_2061900 ^ p93_array_index_2061901 ^ p93_array_index_2061902 ^ p93_array_index_2061903 ^ p93_array_index_2061904 ^ p93_array_index_2061905 ^ p93_bit_slice_2061825;
  assign p94_array_index_2062033_comb = p93_literal_2043920[p93_bit_slice_2061834];
  assign p94_array_index_2062034_comb = p93_literal_2043918[p93_res7__1249];
  assign p94_array_index_2062035_comb = p93_literal_2043916[p93_res7__1251];
  assign p94_array_index_2062036_comb = p93_literal_2043914[p93_res7__1253];
  assign p94_res7__1259_comb = p93_literal_2043910[p93_bit_slice_2061827] ^ p93_literal_2043912[p93_bit_slice_2061841] ^ p93_literal_2043914[p93_bit_slice_2061828] ^ p93_literal_2043916[p93_bit_slice_2061843] ^ p93_literal_2043918[p93_bit_slice_2061829] ^ p93_array_index_2061859 ^ p93_bit_slice_2061831 ^ p93_literal_2043923[p93_bit_slice_2061832] ^ p93_bit_slice_2061833 ^ p94_array_index_2062033_comb ^ p94_array_index_2062034_comb ^ p94_array_index_2062035_comb ^ p94_array_index_2062036_comb ^ p93_literal_2043912[p93_res7__1255] ^ p93_literal_2043910[p94_res7__1257_comb] ^ p93_bit_slice_2061826;
  assign p94_array_index_2062045_comb = p93_literal_2043920[p93_res7__1249];
  assign p94_array_index_2062046_comb = p93_literal_2043918[p93_res7__1251];
  assign p94_array_index_2062047_comb = p93_literal_2043916[p93_res7__1253];
  assign p94_res7__1261_comb = p93_literal_2043910[p93_bit_slice_2061841] ^ p93_literal_2043912[p93_bit_slice_2061828] ^ p93_literal_2043914[p93_bit_slice_2061843] ^ p93_literal_2043916[p93_bit_slice_2061829] ^ p93_array_index_2061845 ^ p93_array_index_2061873 ^ p93_bit_slice_2061832 ^ p93_literal_2043923[p93_bit_slice_2061833] ^ p93_bit_slice_2061834 ^ p94_array_index_2062045_comb ^ p94_array_index_2062046_comb ^ p94_array_index_2062047_comb ^ p93_literal_2043914[p93_res7__1255] ^ p93_literal_2043912[p94_res7__1257_comb] ^ p93_literal_2043910[p94_res7__1259_comb] ^ p93_bit_slice_2061827;
  assign p94_array_index_2062057_comb = p93_literal_2043920[p93_res7__1251];
  assign p94_array_index_2062058_comb = p93_literal_2043918[p93_res7__1253];
  assign p94_array_index_2062059_comb = p93_literal_2043916[p93_res7__1255];
  assign p94_res7__1263_comb = p93_literal_2043910[p93_bit_slice_2061828] ^ p93_literal_2043912[p93_bit_slice_2061843] ^ p93_literal_2043914[p93_bit_slice_2061829] ^ p93_literal_2043916[p93_bit_slice_2061830] ^ p93_array_index_2061860 ^ p93_array_index_2061887 ^ p93_bit_slice_2061833 ^ p93_literal_2043923[p93_bit_slice_2061834] ^ p93_res7__1249 ^ p94_array_index_2062057_comb ^ p94_array_index_2062058_comb ^ p94_array_index_2062059_comb ^ p93_literal_2043914[p94_res7__1257_comb] ^ p93_literal_2043912[p94_res7__1259_comb] ^ p93_literal_2043910[p94_res7__1261_comb] ^ p93_bit_slice_2061841;
  assign p94_array_index_2062068_comb = p93_literal_2043920[p93_res7__1253];
  assign p94_array_index_2062069_comb = p93_literal_2043918[p93_res7__1255];
  assign p94_res7__1265_comb = p93_literal_2043910[p93_bit_slice_2061843] ^ p93_literal_2043912[p93_bit_slice_2061829] ^ p93_literal_2043914[p93_bit_slice_2061830] ^ p93_array_index_2061846 ^ p93_array_index_2061874 ^ p93_array_index_2061900 ^ p93_bit_slice_2061834 ^ p93_literal_2043923[p93_res7__1249] ^ p93_res7__1251 ^ p94_array_index_2062068_comb ^ p94_array_index_2062069_comb ^ p93_literal_2043916[p94_res7__1257_comb] ^ p93_literal_2043914[p94_res7__1259_comb] ^ p93_literal_2043912[p94_res7__1261_comb] ^ p93_literal_2043910[p94_res7__1263_comb] ^ p93_bit_slice_2061828;
  assign p94_array_index_2062079_comb = p93_literal_2043920[p93_res7__1255];
  assign p94_array_index_2062080_comb = p93_literal_2043918[p94_res7__1257_comb];
  assign p94_res7__1267_comb = p93_literal_2043910[p93_bit_slice_2061829] ^ p93_literal_2043912[p93_bit_slice_2061830] ^ p93_literal_2043914[p93_bit_slice_2061831] ^ p93_array_index_2061861 ^ p93_array_index_2061888 ^ p94_array_index_2062033_comb ^ p93_res7__1249 ^ p93_literal_2043923[p93_res7__1251] ^ p93_res7__1253 ^ p94_array_index_2062079_comb ^ p94_array_index_2062080_comb ^ p93_literal_2043916[p94_res7__1259_comb] ^ p93_literal_2043914[p94_res7__1261_comb] ^ p93_literal_2043912[p94_res7__1263_comb] ^ p93_literal_2043910[p94_res7__1265_comb] ^ p93_bit_slice_2061843;
  assign p94_array_index_2062089_comb = p93_literal_2043920[p94_res7__1257_comb];
  assign p94_res7__1269_comb = p93_literal_2043910[p93_bit_slice_2061830] ^ p93_literal_2043912[p93_bit_slice_2061831] ^ p93_array_index_2061847 ^ p93_array_index_2061875 ^ p93_array_index_2061901 ^ p94_array_index_2062045_comb ^ p93_res7__1251 ^ p93_literal_2043923[p93_res7__1253] ^ p93_res7__1255 ^ p94_array_index_2062089_comb ^ p93_literal_2043918[p94_res7__1259_comb] ^ p93_literal_2043916[p94_res7__1261_comb] ^ p93_literal_2043914[p94_res7__1263_comb] ^ p93_literal_2043912[p94_res7__1265_comb] ^ p93_literal_2043910[p94_res7__1267_comb] ^ p93_bit_slice_2061829;
  assign p94_array_index_2062096_comb = p93_literal_2043910[p93_bit_slice_2061831];
  assign p94_array_index_2062097_comb = p93_literal_2043912[p93_bit_slice_2061832];
  assign p94_array_index_2062098_comb = p93_literal_2043923[p93_res7__1255];
  assign p94_array_index_2062099_comb = p93_literal_2043920[p94_res7__1259_comb];
  assign p94_array_index_2062100_comb = p93_literal_2043918[p94_res7__1261_comb];
  assign p94_array_index_2062101_comb = p93_literal_2043916[p94_res7__1263_comb];
  assign p94_array_index_2062102_comb = p93_literal_2043914[p94_res7__1265_comb];
  assign p94_array_index_2062103_comb = p93_literal_2043912[p94_res7__1267_comb];
  assign p94_array_index_2062104_comb = p93_literal_2043910[p94_res7__1269_comb];
  assign p94_array_index_2062105_comb = p93_literal_2058836[p93_res7__1249];
  assign p94_array_index_2062106_comb = p93_literal_2058836[p93_res7__1251];

  // Registers for pipe stage 94:
  reg [127:0] p94_bit_slice_2043893;
  reg [127:0] p94_bit_slice_2044018;
  reg [7:0] p94_bit_slice_2061830;
  reg [7:0] p94_bit_slice_2061831;
  reg [7:0] p94_bit_slice_2061832;
  reg [7:0] p94_bit_slice_2061833;
  reg [7:0] p94_bit_slice_2061834;
  reg [7:0] p94_array_index_2061848;
  reg [7:0] p94_array_index_2061849;
  reg [7:0] p94_array_index_2061862;
  reg [7:0] p94_array_index_2061863;
  reg [7:0] p94_array_index_2061864;
  reg [7:0] p94_array_index_2061876;
  reg [7:0] p94_array_index_2061877;
  reg [7:0] p94_res7__1253;
  reg [7:0] p94_array_index_2061889;
  reg [7:0] p94_array_index_2061890;
  reg [7:0] p94_array_index_2061891;
  reg [7:0] p94_res7__1255;
  reg [7:0] p94_array_index_2061902;
  reg [7:0] p94_array_index_2061903;
  reg [7:0] p94_res7__1257;
  reg [7:0] p94_array_index_2062034;
  reg [7:0] p94_array_index_2062035;
  reg [7:0] p94_array_index_2062036;
  reg [7:0] p94_res7__1259;
  reg [7:0] p94_array_index_2062046;
  reg [7:0] p94_array_index_2062047;
  reg [7:0] p94_res7__1261;
  reg [7:0] p94_array_index_2062057;
  reg [7:0] p94_array_index_2062058;
  reg [7:0] p94_array_index_2062059;
  reg [7:0] p94_res7__1263;
  reg [7:0] p94_array_index_2062068;
  reg [7:0] p94_array_index_2062069;
  reg [7:0] p94_res7__1265;
  reg [7:0] p94_array_index_2062079;
  reg [7:0] p94_array_index_2062080;
  reg [7:0] p94_res7__1267;
  reg [7:0] p94_array_index_2062089;
  reg [7:0] p94_res7__1269;
  reg [7:0] p94_array_index_2062096;
  reg [7:0] p94_array_index_2062097;
  reg [7:0] p94_array_index_2062098;
  reg [7:0] p94_array_index_2062099;
  reg [7:0] p94_array_index_2062100;
  reg [7:0] p94_array_index_2062101;
  reg [7:0] p94_array_index_2062102;
  reg [7:0] p94_array_index_2062103;
  reg [7:0] p94_array_index_2062104;
  reg [7:0] p94_array_index_2062105;
  reg [7:0] p94_array_index_2062106;
  reg [7:0] p95_literal_2043910[256];
  reg [7:0] p95_literal_2043912[256];
  reg [7:0] p95_literal_2043914[256];
  reg [7:0] p95_literal_2043916[256];
  reg [7:0] p95_literal_2043918[256];
  reg [7:0] p95_literal_2043920[256];
  reg [7:0] p95_literal_2043923[256];
  always_ff @ (posedge clk) begin
    p94_bit_slice_2043893 <= p93_bit_slice_2043893;
    p94_bit_slice_2044018 <= p93_bit_slice_2044018;
    p94_bit_slice_2061830 <= p93_bit_slice_2061830;
    p94_bit_slice_2061831 <= p93_bit_slice_2061831;
    p94_bit_slice_2061832 <= p93_bit_slice_2061832;
    p94_bit_slice_2061833 <= p93_bit_slice_2061833;
    p94_bit_slice_2061834 <= p93_bit_slice_2061834;
    p94_array_index_2061848 <= p93_array_index_2061848;
    p94_array_index_2061849 <= p93_array_index_2061849;
    p94_array_index_2061862 <= p93_array_index_2061862;
    p94_array_index_2061863 <= p93_array_index_2061863;
    p94_array_index_2061864 <= p93_array_index_2061864;
    p94_array_index_2061876 <= p93_array_index_2061876;
    p94_array_index_2061877 <= p93_array_index_2061877;
    p94_res7__1253 <= p93_res7__1253;
    p94_array_index_2061889 <= p93_array_index_2061889;
    p94_array_index_2061890 <= p93_array_index_2061890;
    p94_array_index_2061891 <= p93_array_index_2061891;
    p94_res7__1255 <= p93_res7__1255;
    p94_array_index_2061902 <= p93_array_index_2061902;
    p94_array_index_2061903 <= p93_array_index_2061903;
    p94_res7__1257 <= p94_res7__1257_comb;
    p94_array_index_2062034 <= p94_array_index_2062034_comb;
    p94_array_index_2062035 <= p94_array_index_2062035_comb;
    p94_array_index_2062036 <= p94_array_index_2062036_comb;
    p94_res7__1259 <= p94_res7__1259_comb;
    p94_array_index_2062046 <= p94_array_index_2062046_comb;
    p94_array_index_2062047 <= p94_array_index_2062047_comb;
    p94_res7__1261 <= p94_res7__1261_comb;
    p94_array_index_2062057 <= p94_array_index_2062057_comb;
    p94_array_index_2062058 <= p94_array_index_2062058_comb;
    p94_array_index_2062059 <= p94_array_index_2062059_comb;
    p94_res7__1263 <= p94_res7__1263_comb;
    p94_array_index_2062068 <= p94_array_index_2062068_comb;
    p94_array_index_2062069 <= p94_array_index_2062069_comb;
    p94_res7__1265 <= p94_res7__1265_comb;
    p94_array_index_2062079 <= p94_array_index_2062079_comb;
    p94_array_index_2062080 <= p94_array_index_2062080_comb;
    p94_res7__1267 <= p94_res7__1267_comb;
    p94_array_index_2062089 <= p94_array_index_2062089_comb;
    p94_res7__1269 <= p94_res7__1269_comb;
    p94_array_index_2062096 <= p94_array_index_2062096_comb;
    p94_array_index_2062097 <= p94_array_index_2062097_comb;
    p94_array_index_2062098 <= p94_array_index_2062098_comb;
    p94_array_index_2062099 <= p94_array_index_2062099_comb;
    p94_array_index_2062100 <= p94_array_index_2062100_comb;
    p94_array_index_2062101 <= p94_array_index_2062101_comb;
    p94_array_index_2062102 <= p94_array_index_2062102_comb;
    p94_array_index_2062103 <= p94_array_index_2062103_comb;
    p94_array_index_2062104 <= p94_array_index_2062104_comb;
    p94_array_index_2062105 <= p94_array_index_2062105_comb;
    p94_array_index_2062106 <= p94_array_index_2062106_comb;
    p95_literal_2043910 <= p94_literal_2043910;
    p95_literal_2043912 <= p94_literal_2043912;
    p95_literal_2043914 <= p94_literal_2043914;
    p95_literal_2043916 <= p94_literal_2043916;
    p95_literal_2043918 <= p94_literal_2043918;
    p95_literal_2043920 <= p94_literal_2043920;
    p95_literal_2043923 <= p94_literal_2043923;
  end

  // ===== Pipe stage 95:
  wire [7:0] p95_res7__1271_comb;
  wire [7:0] p95_res7__1273_comb;
  wire [7:0] p95_res7__1275_comb;
  wire [7:0] p95_res7__1277_comb;
  wire [7:0] p95_res7__1279_comb;
  wire [127:0] p95_permut__39_comb;
  wire [127:0] p95_xor_2062277_comb;
  wire [7:0] p95_bit_slice_2062278_comb;
  wire [7:0] p95_bit_slice_2062279_comb;
  wire [7:0] p95_bit_slice_2062280_comb;
  wire [7:0] p95_bit_slice_2062281_comb;
  wire [7:0] p95_bit_slice_2062282_comb;
  wire [7:0] p95_bit_slice_2062283_comb;
  wire [7:0] p95_bit_slice_2062284_comb;
  wire [7:0] p95_bit_slice_2062285_comb;
  wire [7:0] p95_bit_slice_2062286_comb;
  wire [7:0] p95_bit_slice_2062287_comb;
  wire [7:0] p95_bit_slice_2062288_comb;
  wire [7:0] p95_bit_slice_2062289_comb;
  wire [7:0] p95_bit_slice_2062290_comb;
  wire [7:0] p95_bit_slice_2062297_comb;
  wire [7:0] p95_bit_slice_2062299_comb;
  wire [7:0] p95_array_index_2062300_comb;
  wire [7:0] p95_array_index_2062301_comb;
  wire [7:0] p95_array_index_2062302_comb;
  wire [7:0] p95_array_index_2062303_comb;
  wire [7:0] p95_array_index_2062304_comb;
  wire [7:0] p95_array_index_2062305_comb;
  wire [7:0] p95_res7__1281_comb;
  wire [7:0] p95_array_index_2062308_comb;
  wire [7:0] p95_array_index_2062309_comb;
  wire [7:0] p95_array_index_2062310_comb;
  wire [7:0] p95_array_index_2062311_comb;
  wire [7:0] p95_array_index_2062312_comb;
  wire [7:0] p95_array_index_2062313_comb;
  wire [7:0] p95_array_index_2062314_comb;
  wire [7:0] p95_array_index_2062315_comb;
  wire [7:0] p95_array_index_2062316_comb;
  wire [7:0] p95_array_index_2062317_comb;
  wire [7:0] p95_array_index_2062318_comb;
  wire [7:0] p95_array_index_2062319_comb;
  wire [7:0] p95_array_index_2062320_comb;
  assign p95_res7__1271_comb = p94_array_index_2062096 ^ p94_array_index_2062097 ^ p94_array_index_2061862 ^ p94_array_index_2061889 ^ p94_array_index_2062034 ^ p94_array_index_2062057 ^ p94_res7__1253 ^ p94_array_index_2062098 ^ p94_res7__1257 ^ p94_array_index_2062099 ^ p94_array_index_2062100 ^ p94_array_index_2062101 ^ p94_array_index_2062102 ^ p94_array_index_2062103 ^ p94_array_index_2062104 ^ p94_bit_slice_2061830;
  assign p95_res7__1273_comb = p94_literal_2043910[p94_bit_slice_2061832] ^ p94_array_index_2061848 ^ p94_array_index_2061876 ^ p94_array_index_2061902 ^ p94_array_index_2062046 ^ p94_array_index_2062068 ^ p94_res7__1255 ^ p94_literal_2043923[p94_res7__1257] ^ p94_res7__1259 ^ p94_literal_2043920[p94_res7__1261] ^ p94_literal_2043918[p94_res7__1263] ^ p94_literal_2043916[p94_res7__1265] ^ p94_literal_2043914[p94_res7__1267] ^ p94_literal_2043912[p94_res7__1269] ^ p94_literal_2043910[p95_res7__1271_comb] ^ p94_bit_slice_2061831;
  assign p95_res7__1275_comb = p94_literal_2043910[p94_bit_slice_2061833] ^ p94_array_index_2061863 ^ p94_array_index_2061890 ^ p94_array_index_2062035 ^ p94_array_index_2062058 ^ p94_array_index_2062079 ^ p94_res7__1257 ^ p94_literal_2043923[p94_res7__1259] ^ p94_res7__1261 ^ p94_literal_2043920[p94_res7__1263] ^ p94_literal_2043918[p94_res7__1265] ^ p94_literal_2043916[p94_res7__1267] ^ p94_literal_2043914[p94_res7__1269] ^ p94_literal_2043912[p95_res7__1271_comb] ^ p94_literal_2043910[p95_res7__1273_comb] ^ p94_bit_slice_2061832;
  assign p95_res7__1277_comb = p94_array_index_2061849 ^ p94_array_index_2061877 ^ p94_array_index_2061903 ^ p94_array_index_2062047 ^ p94_array_index_2062069 ^ p94_array_index_2062089 ^ p94_res7__1259 ^ p94_literal_2043923[p94_res7__1261] ^ p94_res7__1263 ^ p94_literal_2043920[p94_res7__1265] ^ p94_literal_2043918[p94_res7__1267] ^ p94_literal_2043916[p94_res7__1269] ^ p94_literal_2043914[p95_res7__1271_comb] ^ p94_literal_2043912[p95_res7__1273_comb] ^ p94_literal_2043910[p95_res7__1275_comb] ^ p94_bit_slice_2061833;
  assign p95_res7__1279_comb = p94_array_index_2061864 ^ p94_array_index_2061891 ^ p94_array_index_2062036 ^ p94_array_index_2062059 ^ p94_array_index_2062080 ^ p94_array_index_2062099 ^ p94_res7__1261 ^ p94_literal_2043923[p94_res7__1263] ^ p94_res7__1265 ^ p94_literal_2043920[p94_res7__1267] ^ p94_literal_2043918[p94_res7__1269] ^ p94_literal_2043916[p95_res7__1271_comb] ^ p94_literal_2043914[p95_res7__1273_comb] ^ p94_literal_2043912[p95_res7__1275_comb] ^ p94_literal_2043910[p95_res7__1277_comb] ^ p94_bit_slice_2061834;
  assign p95_permut__39_comb = {p94_array_index_2062105, p94_array_index_2062106, p94_literal_2058836[p94_res7__1253], p94_literal_2058836[p94_res7__1255], p94_literal_2058836[p94_res7__1257], p94_literal_2058836[p94_res7__1259], p94_literal_2058836[p94_res7__1261], p94_literal_2058836[p94_res7__1263], p94_literal_2058836[p94_res7__1265], p94_literal_2058836[p94_res7__1267], p94_literal_2058836[p94_res7__1269], p94_literal_2058836[p95_res7__1271_comb], p94_literal_2058836[p95_res7__1273_comb], p94_literal_2058836[p95_res7__1275_comb], p94_literal_2058836[p95_res7__1277_comb], p94_literal_2058836[p95_res7__1279_comb]};
  assign p95_xor_2062277_comb = p94_bit_slice_2044018 ^ p95_permut__39_comb;
  assign p95_bit_slice_2062278_comb = p95_xor_2062277_comb[119:112];
  assign p95_bit_slice_2062279_comb = p95_xor_2062277_comb[111:104];
  assign p95_bit_slice_2062280_comb = p95_xor_2062277_comb[103:96];
  assign p95_bit_slice_2062281_comb = p95_xor_2062277_comb[95:88];
  assign p95_bit_slice_2062282_comb = p95_xor_2062277_comb[87:80];
  assign p95_bit_slice_2062283_comb = p95_xor_2062277_comb[79:72];
  assign p95_bit_slice_2062284_comb = p95_xor_2062277_comb[63:56];
  assign p95_bit_slice_2062285_comb = p95_xor_2062277_comb[47:40];
  assign p95_bit_slice_2062286_comb = p95_xor_2062277_comb[39:32];
  assign p95_bit_slice_2062287_comb = p95_xor_2062277_comb[31:24];
  assign p95_bit_slice_2062288_comb = p95_xor_2062277_comb[23:16];
  assign p95_bit_slice_2062289_comb = p95_xor_2062277_comb[15:8];
  assign p95_bit_slice_2062290_comb = p95_xor_2062277_comb[7:0];
  assign p95_bit_slice_2062297_comb = p95_xor_2062277_comb[71:64];
  assign p95_bit_slice_2062299_comb = p95_xor_2062277_comb[55:48];
  assign p95_array_index_2062300_comb = p94_literal_2043920[p95_bit_slice_2062285_comb];
  assign p95_array_index_2062301_comb = p94_literal_2043918[p95_bit_slice_2062286_comb];
  assign p95_array_index_2062302_comb = p94_literal_2043916[p95_bit_slice_2062287_comb];
  assign p95_array_index_2062303_comb = p94_literal_2043914[p95_bit_slice_2062288_comb];
  assign p95_array_index_2062304_comb = p94_literal_2043912[p95_bit_slice_2062289_comb];
  assign p95_array_index_2062305_comb = p94_literal_2043910[p95_bit_slice_2062290_comb];
  assign p95_res7__1281_comb = p94_literal_2043910[p95_bit_slice_2062278_comb] ^ p94_literal_2043912[p95_bit_slice_2062279_comb] ^ p94_literal_2043914[p95_bit_slice_2062280_comb] ^ p94_literal_2043916[p95_bit_slice_2062281_comb] ^ p94_literal_2043918[p95_bit_slice_2062282_comb] ^ p94_literal_2043920[p95_bit_slice_2062283_comb] ^ p95_bit_slice_2062297_comb ^ p94_literal_2043923[p95_bit_slice_2062284_comb] ^ p95_bit_slice_2062299_comb ^ p95_array_index_2062300_comb ^ p95_array_index_2062301_comb ^ p95_array_index_2062302_comb ^ p95_array_index_2062303_comb ^ p95_array_index_2062304_comb ^ p95_array_index_2062305_comb ^ p95_xor_2062277_comb[127:120];
  assign p95_array_index_2062308_comb = p94_literal_2043910[p95_bit_slice_2062279_comb];
  assign p95_array_index_2062309_comb = p94_literal_2043912[p95_bit_slice_2062280_comb];
  assign p95_array_index_2062310_comb = p94_literal_2043914[p95_bit_slice_2062281_comb];
  assign p95_array_index_2062311_comb = p94_literal_2043916[p95_bit_slice_2062282_comb];
  assign p95_array_index_2062312_comb = p94_literal_2043918[p95_bit_slice_2062283_comb];
  assign p95_array_index_2062313_comb = p94_literal_2043920[p95_bit_slice_2062297_comb];
  assign p95_array_index_2062314_comb = p94_literal_2043923[p95_bit_slice_2062299_comb];
  assign p95_array_index_2062315_comb = p94_literal_2043920[p95_bit_slice_2062286_comb];
  assign p95_array_index_2062316_comb = p94_literal_2043918[p95_bit_slice_2062287_comb];
  assign p95_array_index_2062317_comb = p94_literal_2043916[p95_bit_slice_2062288_comb];
  assign p95_array_index_2062318_comb = p94_literal_2043914[p95_bit_slice_2062289_comb];
  assign p95_array_index_2062319_comb = p94_literal_2043912[p95_bit_slice_2062290_comb];
  assign p95_array_index_2062320_comb = p94_literal_2043910[p95_res7__1281_comb];

  // Registers for pipe stage 95:
  reg [127:0] p95_bit_slice_2043893;
  reg [7:0] p95_bit_slice_2062278;
  reg [7:0] p95_bit_slice_2062279;
  reg [7:0] p95_bit_slice_2062280;
  reg [7:0] p95_bit_slice_2062281;
  reg [7:0] p95_bit_slice_2062282;
  reg [7:0] p95_bit_slice_2062283;
  reg [7:0] p95_bit_slice_2062284;
  reg [7:0] p95_bit_slice_2062285;
  reg [7:0] p95_bit_slice_2062286;
  reg [7:0] p95_bit_slice_2062287;
  reg [7:0] p95_bit_slice_2062288;
  reg [7:0] p95_bit_slice_2062289;
  reg [7:0] p95_bit_slice_2062290;
  reg [7:0] p95_bit_slice_2062297;
  reg [7:0] p95_bit_slice_2062299;
  reg [7:0] p95_array_index_2062300;
  reg [7:0] p95_array_index_2062301;
  reg [7:0] p95_array_index_2062302;
  reg [7:0] p95_array_index_2062303;
  reg [7:0] p95_array_index_2062304;
  reg [7:0] p95_array_index_2062305;
  reg [7:0] p95_res7__1281;
  reg [7:0] p95_array_index_2062308;
  reg [7:0] p95_array_index_2062309;
  reg [7:0] p95_array_index_2062310;
  reg [7:0] p95_array_index_2062311;
  reg [7:0] p95_array_index_2062312;
  reg [7:0] p95_array_index_2062313;
  reg [7:0] p95_array_index_2062314;
  reg [7:0] p95_array_index_2062315;
  reg [7:0] p95_array_index_2062316;
  reg [7:0] p95_array_index_2062317;
  reg [7:0] p95_array_index_2062318;
  reg [7:0] p95_array_index_2062319;
  reg [7:0] p95_array_index_2062320;
  reg [7:0] p96_literal_2043910[256];
  reg [7:0] p96_literal_2043912[256];
  reg [7:0] p96_literal_2043914[256];
  reg [7:0] p96_literal_2043916[256];
  reg [7:0] p96_literal_2043918[256];
  reg [7:0] p96_literal_2043920[256];
  always_ff @ (posedge clk) begin
    p95_bit_slice_2043893 <= p94_bit_slice_2043893;
    p95_bit_slice_2062278 <= p95_bit_slice_2062278_comb;
    p95_bit_slice_2062279 <= p95_bit_slice_2062279_comb;
    p95_bit_slice_2062280 <= p95_bit_slice_2062280_comb;
    p95_bit_slice_2062281 <= p95_bit_slice_2062281_comb;
    p95_bit_slice_2062282 <= p95_bit_slice_2062282_comb;
    p95_bit_slice_2062283 <= p95_bit_slice_2062283_comb;
    p95_bit_slice_2062284 <= p95_bit_slice_2062284_comb;
    p95_bit_slice_2062285 <= p95_bit_slice_2062285_comb;
    p95_bit_slice_2062286 <= p95_bit_slice_2062286_comb;
    p95_bit_slice_2062287 <= p95_bit_slice_2062287_comb;
    p95_bit_slice_2062288 <= p95_bit_slice_2062288_comb;
    p95_bit_slice_2062289 <= p95_bit_slice_2062289_comb;
    p95_bit_slice_2062290 <= p95_bit_slice_2062290_comb;
    p95_bit_slice_2062297 <= p95_bit_slice_2062297_comb;
    p95_bit_slice_2062299 <= p95_bit_slice_2062299_comb;
    p95_array_index_2062300 <= p95_array_index_2062300_comb;
    p95_array_index_2062301 <= p95_array_index_2062301_comb;
    p95_array_index_2062302 <= p95_array_index_2062302_comb;
    p95_array_index_2062303 <= p95_array_index_2062303_comb;
    p95_array_index_2062304 <= p95_array_index_2062304_comb;
    p95_array_index_2062305 <= p95_array_index_2062305_comb;
    p95_res7__1281 <= p95_res7__1281_comb;
    p95_array_index_2062308 <= p95_array_index_2062308_comb;
    p95_array_index_2062309 <= p95_array_index_2062309_comb;
    p95_array_index_2062310 <= p95_array_index_2062310_comb;
    p95_array_index_2062311 <= p95_array_index_2062311_comb;
    p95_array_index_2062312 <= p95_array_index_2062312_comb;
    p95_array_index_2062313 <= p95_array_index_2062313_comb;
    p95_array_index_2062314 <= p95_array_index_2062314_comb;
    p95_array_index_2062315 <= p95_array_index_2062315_comb;
    p95_array_index_2062316 <= p95_array_index_2062316_comb;
    p95_array_index_2062317 <= p95_array_index_2062317_comb;
    p95_array_index_2062318 <= p95_array_index_2062318_comb;
    p95_array_index_2062319 <= p95_array_index_2062319_comb;
    p95_array_index_2062320 <= p95_array_index_2062320_comb;
    p96_literal_2043910 <= p95_literal_2043910;
    p96_literal_2043912 <= p95_literal_2043912;
    p96_literal_2043914 <= p95_literal_2043914;
    p96_literal_2043916 <= p95_literal_2043916;
    p96_literal_2043918 <= p95_literal_2043918;
    p96_literal_2043920 <= p95_literal_2043920;
  end

  // ===== Pipe stage 96:
  wire [7:0] p96_res7__1283_comb;
  wire [7:0] p96_array_index_2062417_comb;
  wire [7:0] p96_array_index_2062418_comb;
  wire [7:0] p96_array_index_2062419_comb;
  wire [7:0] p96_array_index_2062420_comb;
  wire [7:0] p96_array_index_2062421_comb;
  wire [7:0] p96_res7__1285_comb;
  wire [7:0] p96_array_index_2062431_comb;
  wire [7:0] p96_array_index_2062432_comb;
  wire [7:0] p96_array_index_2062433_comb;
  wire [7:0] p96_array_index_2062434_comb;
  wire [7:0] p96_array_index_2062435_comb;
  wire [7:0] p96_res7__1287_comb;
  wire [7:0] p96_array_index_2062444_comb;
  wire [7:0] p96_array_index_2062445_comb;
  wire [7:0] p96_array_index_2062446_comb;
  wire [7:0] p96_array_index_2062447_comb;
  wire [7:0] p96_res7__1289_comb;
  wire [7:0] p96_array_index_2062457_comb;
  wire [7:0] p96_array_index_2062458_comb;
  wire [7:0] p96_array_index_2062459_comb;
  wire [7:0] p96_array_index_2062460_comb;
  wire [7:0] p96_res7__1291_comb;
  wire [7:0] p96_array_index_2062469_comb;
  wire [7:0] p96_array_index_2062470_comb;
  wire [7:0] p96_array_index_2062471_comb;
  wire [7:0] p96_res7__1293_comb;
  wire [7:0] p96_array_index_2062481_comb;
  wire [7:0] p96_array_index_2062482_comb;
  wire [7:0] p96_array_index_2062483_comb;
  wire [7:0] p96_res7__1295_comb;
  wire [7:0] p96_array_index_2062488_comb;
  wire [7:0] p96_array_index_2062489_comb;
  wire [7:0] p96_array_index_2062490_comb;
  wire [7:0] p96_array_index_2062491_comb;
  wire [7:0] p96_array_index_2062492_comb;
  wire [7:0] p96_array_index_2062493_comb;
  wire [7:0] p96_array_index_2062494_comb;
  wire [7:0] p96_array_index_2062495_comb;
  wire [7:0] p96_array_index_2062496_comb;
  wire [7:0] p96_array_index_2062497_comb;
  wire [7:0] p96_array_index_2062498_comb;
  wire [7:0] p96_array_index_2062499_comb;
  wire [7:0] p96_array_index_2062500_comb;
  wire [7:0] p96_array_index_2062501_comb;
  wire [7:0] p96_array_index_2062502_comb;
  wire [7:0] p96_array_index_2062503_comb;
  wire [7:0] p96_array_index_2062504_comb;
  assign p96_res7__1283_comb = p95_array_index_2062308 ^ p95_array_index_2062309 ^ p95_array_index_2062310 ^ p95_array_index_2062311 ^ p95_array_index_2062312 ^ p95_array_index_2062313 ^ p95_bit_slice_2062284 ^ p95_array_index_2062314 ^ p95_bit_slice_2062285 ^ p95_array_index_2062315 ^ p95_array_index_2062316 ^ p95_array_index_2062317 ^ p95_array_index_2062318 ^ p95_array_index_2062319 ^ p95_array_index_2062320 ^ p95_bit_slice_2062278;
  assign p96_array_index_2062417_comb = p95_literal_2043920[p95_bit_slice_2062287];
  assign p96_array_index_2062418_comb = p95_literal_2043918[p95_bit_slice_2062288];
  assign p96_array_index_2062419_comb = p95_literal_2043916[p95_bit_slice_2062289];
  assign p96_array_index_2062420_comb = p95_literal_2043914[p95_bit_slice_2062290];
  assign p96_array_index_2062421_comb = p95_literal_2043912[p95_res7__1281];
  assign p96_res7__1285_comb = p95_literal_2043910[p95_bit_slice_2062280] ^ p95_literal_2043912[p95_bit_slice_2062281] ^ p95_literal_2043914[p95_bit_slice_2062282] ^ p95_literal_2043916[p95_bit_slice_2062283] ^ p95_literal_2043918[p95_bit_slice_2062297] ^ p95_literal_2043920[p95_bit_slice_2062284] ^ p95_bit_slice_2062299 ^ p95_literal_2043923[p95_bit_slice_2062285] ^ p95_bit_slice_2062286 ^ p96_array_index_2062417_comb ^ p96_array_index_2062418_comb ^ p96_array_index_2062419_comb ^ p96_array_index_2062420_comb ^ p96_array_index_2062421_comb ^ p95_literal_2043910[p96_res7__1283_comb] ^ p95_bit_slice_2062279;
  assign p96_array_index_2062431_comb = p95_literal_2043920[p95_bit_slice_2062288];
  assign p96_array_index_2062432_comb = p95_literal_2043918[p95_bit_slice_2062289];
  assign p96_array_index_2062433_comb = p95_literal_2043916[p95_bit_slice_2062290];
  assign p96_array_index_2062434_comb = p95_literal_2043914[p95_res7__1281];
  assign p96_array_index_2062435_comb = p95_literal_2043912[p96_res7__1283_comb];
  assign p96_res7__1287_comb = p95_literal_2043910[p95_bit_slice_2062281] ^ p95_literal_2043912[p95_bit_slice_2062282] ^ p95_literal_2043914[p95_bit_slice_2062283] ^ p95_literal_2043916[p95_bit_slice_2062297] ^ p95_literal_2043918[p95_bit_slice_2062284] ^ p95_literal_2043920[p95_bit_slice_2062299] ^ p95_bit_slice_2062285 ^ p95_literal_2043923[p95_bit_slice_2062286] ^ p95_bit_slice_2062287 ^ p96_array_index_2062431_comb ^ p96_array_index_2062432_comb ^ p96_array_index_2062433_comb ^ p96_array_index_2062434_comb ^ p96_array_index_2062435_comb ^ p95_literal_2043910[p96_res7__1285_comb] ^ p95_bit_slice_2062280;
  assign p96_array_index_2062444_comb = p95_literal_2043920[p95_bit_slice_2062289];
  assign p96_array_index_2062445_comb = p95_literal_2043918[p95_bit_slice_2062290];
  assign p96_array_index_2062446_comb = p95_literal_2043916[p95_res7__1281];
  assign p96_array_index_2062447_comb = p95_literal_2043914[p96_res7__1283_comb];
  assign p96_res7__1289_comb = p95_literal_2043910[p95_bit_slice_2062282] ^ p95_literal_2043912[p95_bit_slice_2062283] ^ p95_literal_2043914[p95_bit_slice_2062297] ^ p95_literal_2043916[p95_bit_slice_2062284] ^ p95_literal_2043918[p95_bit_slice_2062299] ^ p95_array_index_2062300 ^ p95_bit_slice_2062286 ^ p95_literal_2043923[p95_bit_slice_2062287] ^ p95_bit_slice_2062288 ^ p96_array_index_2062444_comb ^ p96_array_index_2062445_comb ^ p96_array_index_2062446_comb ^ p96_array_index_2062447_comb ^ p95_literal_2043912[p96_res7__1285_comb] ^ p95_literal_2043910[p96_res7__1287_comb] ^ p95_bit_slice_2062281;
  assign p96_array_index_2062457_comb = p95_literal_2043920[p95_bit_slice_2062290];
  assign p96_array_index_2062458_comb = p95_literal_2043918[p95_res7__1281];
  assign p96_array_index_2062459_comb = p95_literal_2043916[p96_res7__1283_comb];
  assign p96_array_index_2062460_comb = p95_literal_2043914[p96_res7__1285_comb];
  assign p96_res7__1291_comb = p95_literal_2043910[p95_bit_slice_2062283] ^ p95_literal_2043912[p95_bit_slice_2062297] ^ p95_literal_2043914[p95_bit_slice_2062284] ^ p95_literal_2043916[p95_bit_slice_2062299] ^ p95_literal_2043918[p95_bit_slice_2062285] ^ p95_array_index_2062315 ^ p95_bit_slice_2062287 ^ p95_literal_2043923[p95_bit_slice_2062288] ^ p95_bit_slice_2062289 ^ p96_array_index_2062457_comb ^ p96_array_index_2062458_comb ^ p96_array_index_2062459_comb ^ p96_array_index_2062460_comb ^ p95_literal_2043912[p96_res7__1287_comb] ^ p95_literal_2043910[p96_res7__1289_comb] ^ p95_bit_slice_2062282;
  assign p96_array_index_2062469_comb = p95_literal_2043920[p95_res7__1281];
  assign p96_array_index_2062470_comb = p95_literal_2043918[p96_res7__1283_comb];
  assign p96_array_index_2062471_comb = p95_literal_2043916[p96_res7__1285_comb];
  assign p96_res7__1293_comb = p95_literal_2043910[p95_bit_slice_2062297] ^ p95_literal_2043912[p95_bit_slice_2062284] ^ p95_literal_2043914[p95_bit_slice_2062299] ^ p95_literal_2043916[p95_bit_slice_2062285] ^ p95_array_index_2062301 ^ p96_array_index_2062417_comb ^ p95_bit_slice_2062288 ^ p95_literal_2043923[p95_bit_slice_2062289] ^ p95_bit_slice_2062290 ^ p96_array_index_2062469_comb ^ p96_array_index_2062470_comb ^ p96_array_index_2062471_comb ^ p95_literal_2043914[p96_res7__1287_comb] ^ p95_literal_2043912[p96_res7__1289_comb] ^ p95_literal_2043910[p96_res7__1291_comb] ^ p95_bit_slice_2062283;
  assign p96_array_index_2062481_comb = p95_literal_2043920[p96_res7__1283_comb];
  assign p96_array_index_2062482_comb = p95_literal_2043918[p96_res7__1285_comb];
  assign p96_array_index_2062483_comb = p95_literal_2043916[p96_res7__1287_comb];
  assign p96_res7__1295_comb = p95_literal_2043910[p95_bit_slice_2062284] ^ p95_literal_2043912[p95_bit_slice_2062299] ^ p95_literal_2043914[p95_bit_slice_2062285] ^ p95_literal_2043916[p95_bit_slice_2062286] ^ p95_array_index_2062316 ^ p96_array_index_2062431_comb ^ p95_bit_slice_2062289 ^ p95_literal_2043923[p95_bit_slice_2062290] ^ p95_res7__1281 ^ p96_array_index_2062481_comb ^ p96_array_index_2062482_comb ^ p96_array_index_2062483_comb ^ p95_literal_2043914[p96_res7__1289_comb] ^ p95_literal_2043912[p96_res7__1291_comb] ^ p95_literal_2043910[p96_res7__1293_comb] ^ p95_bit_slice_2062297;
  assign p96_array_index_2062488_comb = p95_literal_2043910[p95_bit_slice_2062299];
  assign p96_array_index_2062489_comb = p95_literal_2043912[p95_bit_slice_2062285];
  assign p96_array_index_2062490_comb = p95_literal_2043914[p95_bit_slice_2062286];
  assign p96_array_index_2062491_comb = p95_literal_2043923[p95_res7__1281];
  assign p96_array_index_2062492_comb = p95_literal_2043920[p96_res7__1285_comb];
  assign p96_array_index_2062493_comb = p95_literal_2043918[p96_res7__1287_comb];
  assign p96_array_index_2062494_comb = p95_literal_2043916[p96_res7__1289_comb];
  assign p96_array_index_2062495_comb = p95_literal_2043914[p96_res7__1291_comb];
  assign p96_array_index_2062496_comb = p95_literal_2043912[p96_res7__1293_comb];
  assign p96_array_index_2062497_comb = p95_literal_2043910[p96_res7__1295_comb];
  assign p96_array_index_2062498_comb = p95_literal_2043923[p96_res7__1283_comb];
  assign p96_array_index_2062499_comb = p95_literal_2043923[p96_res7__1285_comb];
  assign p96_array_index_2062500_comb = p95_literal_2043923[p96_res7__1287_comb];
  assign p96_array_index_2062501_comb = p95_literal_2043923[p96_res7__1289_comb];
  assign p96_array_index_2062502_comb = p95_literal_2043923[p96_res7__1291_comb];
  assign p96_array_index_2062503_comb = p95_literal_2043923[p96_res7__1293_comb];
  assign p96_array_index_2062504_comb = p95_literal_2043923[p96_res7__1295_comb];

  // Registers for pipe stage 96:
  reg [127:0] p96_bit_slice_2043893;
  reg [7:0] p96_bit_slice_2062284;
  reg [7:0] p96_bit_slice_2062285;
  reg [7:0] p96_bit_slice_2062286;
  reg [7:0] p96_bit_slice_2062287;
  reg [7:0] p96_bit_slice_2062288;
  reg [7:0] p96_bit_slice_2062289;
  reg [7:0] p96_bit_slice_2062290;
  reg [7:0] p96_bit_slice_2062299;
  reg [7:0] p96_array_index_2062302;
  reg [7:0] p96_array_index_2062303;
  reg [7:0] p96_array_index_2062304;
  reg [7:0] p96_array_index_2062305;
  reg [7:0] p96_res7__1281;
  reg [7:0] p96_array_index_2062317;
  reg [7:0] p96_array_index_2062318;
  reg [7:0] p96_array_index_2062319;
  reg [7:0] p96_array_index_2062320;
  reg [7:0] p96_res7__1283;
  reg [7:0] p96_array_index_2062418;
  reg [7:0] p96_array_index_2062419;
  reg [7:0] p96_array_index_2062420;
  reg [7:0] p96_array_index_2062421;
  reg [7:0] p96_res7__1285;
  reg [7:0] p96_array_index_2062432;
  reg [7:0] p96_array_index_2062433;
  reg [7:0] p96_array_index_2062434;
  reg [7:0] p96_array_index_2062435;
  reg [7:0] p96_res7__1287;
  reg [7:0] p96_array_index_2062444;
  reg [7:0] p96_array_index_2062445;
  reg [7:0] p96_array_index_2062446;
  reg [7:0] p96_array_index_2062447;
  reg [7:0] p96_res7__1289;
  reg [7:0] p96_array_index_2062457;
  reg [7:0] p96_array_index_2062458;
  reg [7:0] p96_array_index_2062459;
  reg [7:0] p96_array_index_2062460;
  reg [7:0] p96_res7__1291;
  reg [7:0] p96_array_index_2062469;
  reg [7:0] p96_array_index_2062470;
  reg [7:0] p96_array_index_2062471;
  reg [7:0] p96_res7__1293;
  reg [7:0] p96_array_index_2062481;
  reg [7:0] p96_array_index_2062482;
  reg [7:0] p96_array_index_2062483;
  reg [7:0] p96_res7__1295;
  reg [7:0] p96_array_index_2062488;
  reg [7:0] p96_array_index_2062489;
  reg [7:0] p96_array_index_2062490;
  reg [7:0] p96_array_index_2062491;
  reg [7:0] p96_array_index_2062492;
  reg [7:0] p96_array_index_2062493;
  reg [7:0] p96_array_index_2062494;
  reg [7:0] p96_array_index_2062495;
  reg [7:0] p96_array_index_2062496;
  reg [7:0] p96_array_index_2062497;
  reg [7:0] p96_array_index_2062498;
  reg [7:0] p96_array_index_2062499;
  reg [7:0] p96_array_index_2062500;
  reg [7:0] p96_array_index_2062501;
  reg [7:0] p96_array_index_2062502;
  reg [7:0] p96_array_index_2062503;
  reg [7:0] p96_array_index_2062504;
  always_ff @ (posedge clk) begin
    p96_bit_slice_2043893 <= p95_bit_slice_2043893;
    p96_bit_slice_2062284 <= p95_bit_slice_2062284;
    p96_bit_slice_2062285 <= p95_bit_slice_2062285;
    p96_bit_slice_2062286 <= p95_bit_slice_2062286;
    p96_bit_slice_2062287 <= p95_bit_slice_2062287;
    p96_bit_slice_2062288 <= p95_bit_slice_2062288;
    p96_bit_slice_2062289 <= p95_bit_slice_2062289;
    p96_bit_slice_2062290 <= p95_bit_slice_2062290;
    p96_bit_slice_2062299 <= p95_bit_slice_2062299;
    p96_array_index_2062302 <= p95_array_index_2062302;
    p96_array_index_2062303 <= p95_array_index_2062303;
    p96_array_index_2062304 <= p95_array_index_2062304;
    p96_array_index_2062305 <= p95_array_index_2062305;
    p96_res7__1281 <= p95_res7__1281;
    p96_array_index_2062317 <= p95_array_index_2062317;
    p96_array_index_2062318 <= p95_array_index_2062318;
    p96_array_index_2062319 <= p95_array_index_2062319;
    p96_array_index_2062320 <= p95_array_index_2062320;
    p96_res7__1283 <= p96_res7__1283_comb;
    p96_array_index_2062418 <= p96_array_index_2062418_comb;
    p96_array_index_2062419 <= p96_array_index_2062419_comb;
    p96_array_index_2062420 <= p96_array_index_2062420_comb;
    p96_array_index_2062421 <= p96_array_index_2062421_comb;
    p96_res7__1285 <= p96_res7__1285_comb;
    p96_array_index_2062432 <= p96_array_index_2062432_comb;
    p96_array_index_2062433 <= p96_array_index_2062433_comb;
    p96_array_index_2062434 <= p96_array_index_2062434_comb;
    p96_array_index_2062435 <= p96_array_index_2062435_comb;
    p96_res7__1287 <= p96_res7__1287_comb;
    p96_array_index_2062444 <= p96_array_index_2062444_comb;
    p96_array_index_2062445 <= p96_array_index_2062445_comb;
    p96_array_index_2062446 <= p96_array_index_2062446_comb;
    p96_array_index_2062447 <= p96_array_index_2062447_comb;
    p96_res7__1289 <= p96_res7__1289_comb;
    p96_array_index_2062457 <= p96_array_index_2062457_comb;
    p96_array_index_2062458 <= p96_array_index_2062458_comb;
    p96_array_index_2062459 <= p96_array_index_2062459_comb;
    p96_array_index_2062460 <= p96_array_index_2062460_comb;
    p96_res7__1291 <= p96_res7__1291_comb;
    p96_array_index_2062469 <= p96_array_index_2062469_comb;
    p96_array_index_2062470 <= p96_array_index_2062470_comb;
    p96_array_index_2062471 <= p96_array_index_2062471_comb;
    p96_res7__1293 <= p96_res7__1293_comb;
    p96_array_index_2062481 <= p96_array_index_2062481_comb;
    p96_array_index_2062482 <= p96_array_index_2062482_comb;
    p96_array_index_2062483 <= p96_array_index_2062483_comb;
    p96_res7__1295 <= p96_res7__1295_comb;
    p96_array_index_2062488 <= p96_array_index_2062488_comb;
    p96_array_index_2062489 <= p96_array_index_2062489_comb;
    p96_array_index_2062490 <= p96_array_index_2062490_comb;
    p96_array_index_2062491 <= p96_array_index_2062491_comb;
    p96_array_index_2062492 <= p96_array_index_2062492_comb;
    p96_array_index_2062493 <= p96_array_index_2062493_comb;
    p96_array_index_2062494 <= p96_array_index_2062494_comb;
    p96_array_index_2062495 <= p96_array_index_2062495_comb;
    p96_array_index_2062496 <= p96_array_index_2062496_comb;
    p96_array_index_2062497 <= p96_array_index_2062497_comb;
    p96_array_index_2062498 <= p96_array_index_2062498_comb;
    p96_array_index_2062499 <= p96_array_index_2062499_comb;
    p96_array_index_2062500 <= p96_array_index_2062500_comb;
    p96_array_index_2062501 <= p96_array_index_2062501_comb;
    p96_array_index_2062502 <= p96_array_index_2062502_comb;
    p96_array_index_2062503 <= p96_array_index_2062503_comb;
    p96_array_index_2062504 <= p96_array_index_2062504_comb;
  end

  // ===== Pipe stage 97:
  wire [7:0] p97_res7__1297_comb;
  wire [7:0] p97_array_index_2062651_comb;
  wire [7:0] p97_array_index_2062652_comb;
  wire [7:0] p97_res7__1299_comb;
  wire [7:0] p97_array_index_2062660_comb;
  wire [7:0] p97_res7__1301_comb;
  wire [7:0] p97_array_index_2062669_comb;
  wire [7:0] p97_res7__1303_comb;
  wire [7:0] p97_res7__1305_comb;
  wire [7:0] p97_res7__1307_comb;
  wire [7:0] p97_res7__1309_comb;
  wire [7:0] p97_array_index_2062699_comb;
  wire [7:0] p97_array_index_2062700_comb;
  wire [7:0] p97_array_index_2062701_comb;
  wire [7:0] p97_array_index_2062702_comb;
  wire [7:0] p97_array_index_2062703_comb;
  wire [7:0] p97_array_index_2062704_comb;
  wire [7:0] p97_array_index_2062705_comb;
  wire [7:0] p97_array_index_2062706_comb;
  wire [7:0] p97_array_index_2062707_comb;
  wire [7:0] p97_array_index_2062708_comb;
  wire [7:0] p97_array_index_2062709_comb;
  wire [7:0] p97_array_index_2062710_comb;
  wire [7:0] p97_array_index_2062711_comb;
  wire [7:0] p97_array_index_2062712_comb;
  wire [7:0] p97_array_index_2062713_comb;
  wire [7:0] p97_array_index_2062714_comb;
  wire [7:0] p97_array_index_2062715_comb;
  wire [7:0] p97_array_index_2062716_comb;
  wire [7:0] p97_array_index_2062717_comb;
  assign p97_res7__1297_comb = p96_array_index_2062488 ^ p96_array_index_2062489 ^ p96_array_index_2062490 ^ p96_array_index_2062302 ^ p96_array_index_2062418 ^ p96_array_index_2062444 ^ p96_bit_slice_2062290 ^ p96_array_index_2062491 ^ p96_res7__1283 ^ p96_array_index_2062492 ^ p96_array_index_2062493 ^ p96_array_index_2062494 ^ p96_array_index_2062495 ^ p96_array_index_2062496 ^ p96_array_index_2062497 ^ p96_bit_slice_2062284;
  assign p97_array_index_2062651_comb = p96_literal_2043920[p96_res7__1287];
  assign p97_array_index_2062652_comb = p96_literal_2043918[p96_res7__1289];
  assign p97_res7__1299_comb = p96_literal_2043910[p96_bit_slice_2062285] ^ p96_literal_2043912[p96_bit_slice_2062286] ^ p96_literal_2043914[p96_bit_slice_2062287] ^ p96_array_index_2062317 ^ p96_array_index_2062432 ^ p96_array_index_2062457 ^ p96_res7__1281 ^ p96_array_index_2062498 ^ p96_res7__1285 ^ p97_array_index_2062651_comb ^ p97_array_index_2062652_comb ^ p96_literal_2043916[p96_res7__1291] ^ p96_literal_2043914[p96_res7__1293] ^ p96_literal_2043912[p96_res7__1295] ^ p96_literal_2043910[p97_res7__1297_comb] ^ p96_bit_slice_2062299;
  assign p97_array_index_2062660_comb = p96_literal_2043920[p96_res7__1289];
  assign p97_res7__1301_comb = p96_literal_2043910[p96_bit_slice_2062286] ^ p96_literal_2043912[p96_bit_slice_2062287] ^ p96_array_index_2062303 ^ p96_array_index_2062419 ^ p96_array_index_2062445 ^ p96_array_index_2062469 ^ p96_res7__1283 ^ p96_array_index_2062499 ^ p96_res7__1287 ^ p97_array_index_2062660_comb ^ p96_literal_2043918[p96_res7__1291] ^ p96_literal_2043916[p96_res7__1293] ^ p96_literal_2043914[p96_res7__1295] ^ p96_literal_2043912[p97_res7__1297_comb] ^ p96_literal_2043910[p97_res7__1299_comb] ^ p96_bit_slice_2062285;
  assign p97_array_index_2062669_comb = p96_literal_2043920[p96_res7__1291];
  assign p97_res7__1303_comb = p96_literal_2043910[p96_bit_slice_2062287] ^ p96_literal_2043912[p96_bit_slice_2062288] ^ p96_array_index_2062318 ^ p96_array_index_2062433 ^ p96_array_index_2062458 ^ p96_array_index_2062481 ^ p96_res7__1285 ^ p96_array_index_2062500 ^ p96_res7__1289 ^ p97_array_index_2062669_comb ^ p96_literal_2043918[p96_res7__1293] ^ p96_literal_2043916[p96_res7__1295] ^ p96_literal_2043914[p97_res7__1297_comb] ^ p96_literal_2043912[p97_res7__1299_comb] ^ p96_literal_2043910[p97_res7__1301_comb] ^ p96_bit_slice_2062286;
  assign p97_res7__1305_comb = p96_literal_2043910[p96_bit_slice_2062288] ^ p96_array_index_2062304 ^ p96_array_index_2062420 ^ p96_array_index_2062446 ^ p96_array_index_2062470 ^ p96_array_index_2062492 ^ p96_res7__1287 ^ p96_array_index_2062501 ^ p96_res7__1291 ^ p96_literal_2043920[p96_res7__1293] ^ p96_literal_2043918[p96_res7__1295] ^ p96_literal_2043916[p97_res7__1297_comb] ^ p96_literal_2043914[p97_res7__1299_comb] ^ p96_literal_2043912[p97_res7__1301_comb] ^ p96_literal_2043910[p97_res7__1303_comb] ^ p96_bit_slice_2062287;
  assign p97_res7__1307_comb = p96_literal_2043910[p96_bit_slice_2062289] ^ p96_array_index_2062319 ^ p96_array_index_2062434 ^ p96_array_index_2062459 ^ p96_array_index_2062482 ^ p97_array_index_2062651_comb ^ p96_res7__1289 ^ p96_array_index_2062502 ^ p96_res7__1293 ^ p96_literal_2043920[p96_res7__1295] ^ p96_literal_2043918[p97_res7__1297_comb] ^ p96_literal_2043916[p97_res7__1299_comb] ^ p96_literal_2043914[p97_res7__1301_comb] ^ p96_literal_2043912[p97_res7__1303_comb] ^ p96_literal_2043910[p97_res7__1305_comb] ^ p96_bit_slice_2062288;
  assign p97_res7__1309_comb = p96_array_index_2062305 ^ p96_array_index_2062421 ^ p96_array_index_2062447 ^ p96_array_index_2062471 ^ p96_array_index_2062493 ^ p97_array_index_2062660_comb ^ p96_res7__1291 ^ p96_array_index_2062503 ^ p96_res7__1295 ^ p96_literal_2043920[p97_res7__1297_comb] ^ p96_literal_2043918[p97_res7__1299_comb] ^ p96_literal_2043916[p97_res7__1301_comb] ^ p96_literal_2043914[p97_res7__1303_comb] ^ p96_literal_2043912[p97_res7__1305_comb] ^ p96_literal_2043910[p97_res7__1307_comb] ^ p96_bit_slice_2062289;
  assign p97_array_index_2062699_comb = p96_literal_2043920[p97_res7__1299_comb];
  assign p97_array_index_2062700_comb = p96_literal_2043918[p97_res7__1301_comb];
  assign p97_array_index_2062701_comb = p96_literal_2043916[p97_res7__1303_comb];
  assign p97_array_index_2062702_comb = p96_literal_2043914[p97_res7__1305_comb];
  assign p97_array_index_2062703_comb = p96_literal_2043912[p97_res7__1307_comb];
  assign p97_array_index_2062704_comb = p96_literal_2043910[p97_res7__1309_comb];
  assign p97_array_index_2062705_comb = p96_literal_2058836[p96_res7__1281];
  assign p97_array_index_2062706_comb = p96_literal_2058836[p96_res7__1283];
  assign p97_array_index_2062707_comb = p96_literal_2058836[p96_res7__1285];
  assign p97_array_index_2062708_comb = p96_literal_2058836[p96_res7__1287];
  assign p97_array_index_2062709_comb = p96_literal_2058836[p96_res7__1289];
  assign p97_array_index_2062710_comb = p96_literal_2058836[p96_res7__1291];
  assign p97_array_index_2062711_comb = p96_literal_2058836[p96_res7__1295];
  assign p97_array_index_2062712_comb = p96_literal_2058836[p97_res7__1299_comb];
  assign p97_array_index_2062713_comb = p96_literal_2058836[p97_res7__1301_comb];
  assign p97_array_index_2062714_comb = p96_literal_2058836[p97_res7__1303_comb];
  assign p97_array_index_2062715_comb = p96_literal_2058836[p97_res7__1305_comb];
  assign p97_array_index_2062716_comb = p96_literal_2058836[p97_res7__1307_comb];
  assign p97_array_index_2062717_comb = p96_literal_2058836[p97_res7__1309_comb];

  // Registers for pipe stage 97:
  reg [127:0] p97_bit_slice_2043893;
  reg [7:0] p97_bit_slice_2062290;
  reg [7:0] p97_array_index_2062320;
  reg [7:0] p97_array_index_2062435;
  reg [7:0] p97_array_index_2062460;
  reg [7:0] p97_res7__1293;
  reg [7:0] p97_array_index_2062483;
  reg [7:0] p97_res7__1297;
  reg [7:0] p97_array_index_2062652;
  reg [7:0] p97_array_index_2062669;
  reg [7:0] p97_array_index_2062504;
  reg [7:0] p97_array_index_2062699;
  reg [7:0] p97_array_index_2062700;
  reg [7:0] p97_array_index_2062701;
  reg [7:0] p97_array_index_2062702;
  reg [7:0] p97_array_index_2062703;
  reg [7:0] p97_array_index_2062704;
  reg [7:0] p97_array_index_2062705;
  reg [7:0] p97_array_index_2062706;
  reg [7:0] p97_array_index_2062707;
  reg [7:0] p97_array_index_2062708;
  reg [7:0] p97_array_index_2062709;
  reg [7:0] p97_array_index_2062710;
  reg [7:0] p97_array_index_2062711;
  reg [7:0] p97_array_index_2062712;
  reg [7:0] p97_array_index_2062713;
  reg [7:0] p97_array_index_2062714;
  reg [7:0] p97_array_index_2062715;
  reg [7:0] p97_array_index_2062716;
  reg [7:0] p97_array_index_2062717;
  always_ff @ (posedge clk) begin
    p97_bit_slice_2043893 <= p96_bit_slice_2043893;
    p97_bit_slice_2062290 <= p96_bit_slice_2062290;
    p97_array_index_2062320 <= p96_array_index_2062320;
    p97_array_index_2062435 <= p96_array_index_2062435;
    p97_array_index_2062460 <= p96_array_index_2062460;
    p97_res7__1293 <= p96_res7__1293;
    p97_array_index_2062483 <= p96_array_index_2062483;
    p97_res7__1297 <= p97_res7__1297_comb;
    p97_array_index_2062652 <= p97_array_index_2062652_comb;
    p97_array_index_2062669 <= p97_array_index_2062669_comb;
    p97_array_index_2062504 <= p96_array_index_2062504;
    p97_array_index_2062699 <= p97_array_index_2062699_comb;
    p97_array_index_2062700 <= p97_array_index_2062700_comb;
    p97_array_index_2062701 <= p97_array_index_2062701_comb;
    p97_array_index_2062702 <= p97_array_index_2062702_comb;
    p97_array_index_2062703 <= p97_array_index_2062703_comb;
    p97_array_index_2062704 <= p97_array_index_2062704_comb;
    p97_array_index_2062705 <= p97_array_index_2062705_comb;
    p97_array_index_2062706 <= p97_array_index_2062706_comb;
    p97_array_index_2062707 <= p97_array_index_2062707_comb;
    p97_array_index_2062708 <= p97_array_index_2062708_comb;
    p97_array_index_2062709 <= p97_array_index_2062709_comb;
    p97_array_index_2062710 <= p97_array_index_2062710_comb;
    p97_array_index_2062711 <= p97_array_index_2062711_comb;
    p97_array_index_2062712 <= p97_array_index_2062712_comb;
    p97_array_index_2062713 <= p97_array_index_2062713_comb;
    p97_array_index_2062714 <= p97_array_index_2062714_comb;
    p97_array_index_2062715 <= p97_array_index_2062715_comb;
    p97_array_index_2062716 <= p97_array_index_2062716_comb;
    p97_array_index_2062717 <= p97_array_index_2062717_comb;
  end

  // ===== Pipe stage 98:
  wire [7:0] p98_res7__1311_comb;
  wire [127:0] p98_permut__40_comb;
  assign p98_res7__1311_comb = p97_array_index_2062320 ^ p97_array_index_2062435 ^ p97_array_index_2062460 ^ p97_array_index_2062483 ^ p97_array_index_2062652 ^ p97_array_index_2062669 ^ p97_res7__1293 ^ p97_array_index_2062504 ^ p97_res7__1297 ^ p97_array_index_2062699 ^ p97_array_index_2062700 ^ p97_array_index_2062701 ^ p97_array_index_2062702 ^ p97_array_index_2062703 ^ p97_array_index_2062704 ^ p97_bit_slice_2062290;
  assign p98_permut__40_comb = {p97_array_index_2062705, p97_array_index_2062706, p97_array_index_2062707, p97_array_index_2062708, p97_array_index_2062709, p97_array_index_2062710, p97_literal_2058836[p97_res7__1293], p97_array_index_2062711, p97_literal_2058836[p97_res7__1297], p97_array_index_2062712, p97_array_index_2062713, p97_array_index_2062714, p97_array_index_2062715, p97_array_index_2062716, p97_array_index_2062717, p97_literal_2058836[p98_res7__1311_comb]};

  // Registers for pipe stage 98:
  reg [127:0] p98_bit_slice_2043893;
  reg [127:0] p98_permut__40;
  always_ff @ (posedge clk) begin
    p98_bit_slice_2043893 <= p97_bit_slice_2043893;
    p98_permut__40 <= p98_permut__40_comb;
  end

  // ===== Pipe stage 99:
  wire [127:0] p99_newValue_comb;
  assign p99_newValue_comb = p98_bit_slice_2043893 ^ p98_permut__40;

  // Registers for pipe stage 99:
  reg [127:0] p99_newValue;
  always_ff @ (posedge clk) begin
    p99_newValue <= p99_newValue_comb;
  end
  assign out = p99_newValue;
endmodule
