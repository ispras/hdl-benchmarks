// IWLS benchmark module "MultiplierA_16" printed on Wed May 29 22:12:32 2002
module MultiplierA_16(\1 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \13 , \14 , \15 , \16 , \17 , \18 , \36 );
input
  \1 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ,
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ;
output
  \36 ;
reg
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ,
  \34 ,
  \2 ;
wire
  \[40] ,
  \[26] ,
  \[41] ,
  \[27] ,
  \[42] ,
  \[28] ,
  \[43] ,
  \[29] ,
  \[44] ,
  \[45] ,
  \[60] ,
  \[46] ,
  \86 ,
  \87 ,
  \88 ,
  \89 ,
  \[61] ,
  \90 ,
  \91 ,
  \92 ,
  \93 ,
  \94 ,
  \[47] ,
  \95 ,
  \96 ,
  \97 ,
  \98 ,
  \99 ,
  \[62] ,
  \[48] ,
  \[30] ,
  \[31] ,
  \[17] ,
  \[32] ,
  \[18] ,
  \[33] ,
  \[19] ,
  \[34] ,
  \[35] ,
  \[36] ,
  \[37] ,
  \[38] ,
  \100 ,
  \101 ,
  \102 ,
  \107 ,
  \[39] ,
  \113 ,
  \115 ,
  \117 ,
  \119 ,
  \[20] ,
  \121 ,
  \123 ,
  \125 ,
  \127 ,
  \129 ,
  \[21] ,
  \131 ,
  \133 ,
  \135 ,
  \137 ,
  \[22] ,
  \140 ,
  \[23] ,
  \[24] ,
  \[25] ;
assign
  \[40]  = \121  | \26 ,
  \[26]  = \96 ,
  \[41]  = \123  | \27 ,
  \36  = \87 ,
  \[27]  = \97 ,
  \[42]  = \125  | \28 ,
  \[28]  = \98 ,
  \[43]  = \127  | \29 ,
  \[29]  = \99 ,
  \[44]  = \129  | \30 ,
  \[45]  = \131  | \31 ,
  \[60]  = ~\87  & \20 ,
  \[46]  = \133  | \32 ,
  \86  = (\[62]  & \137 ) | (\[35]  & \34 ),
  \87  = (~\[48]  & ~\20 ) | (\[48]  & \20 ),
  \88  = (\[60]  & (\21  & \4 )) | ((\[33]  & ~\113 ) | (~\113  & \21 )),
  \89  = (~\115  & (\5  & \1 )) | ((\113  & (\22  & \5 )) | (\[36]  & ~\115 )),
  \[61]  = \16  & \1 ,
  \90  = (~\117  & (\6  & \1 )) | ((\115  & (\23  & \6 )) | (\[37]  & ~\117 )),
  \91  = (~\119  & (\7  & \1 )) | ((\117  & (\24  & \7 )) | (\[38]  & ~\119 )),
  \92  = (~\121  & (\8  & \1 )) | ((\119  & (\25  & \8 )) | (\[39]  & ~\121 )),
  \93  = (~\123  & (\9  & \1 )) | ((\121  & (\26  & \9 )) | (\[40]  & ~\123 )),
  \94  = (~\125  & (\10  & \1 )) | ((\123  & (\27  & \10 )) | (\[41]  & ~\125 )),
  \[47]  = ~\18  | ~\1 ,
  \95  = (~\127  & (\11  & \1 )) | ((\125  & (\28  & \11 )) | (\[42]  & ~\127 )),
  \96  = (~\129  & (\12  & \1 )) | ((\127  & (\29  & \12 )) | (\[43]  & ~\129 )),
  \97  = (~\131  & (\13  & \1 )) | ((\129  & (\30  & \13 )) | (\[44]  & ~\131 )),
  \98  = (~\133  & (\14  & \1 )) | ((\131  & (\31  & \14 )) | (\[45]  & ~\133 )),
  \99  = (~\135  & (\15  & \1 )) | ((\133  & (\32  & \15 )) | (\[46]  & ~\135 )),
  \[62]  = \17  & \1 ,
  \[48]  = ~\3  | ~\1 ,
  \[30]  = \100 ,
  \[31]  = \101 ,
  \[17]  = \107 ,
  \[32]  = \102 ,
  \[18]  = \88 ,
  \[33]  = (\4  & \1 ) | \[60] ,
  \[19]  = \89 ,
  \[34]  = \[61]  | \135 ,
  \[35]  = \[62]  | \137 ,
  \[36]  = \113  | \22 ,
  \[37]  = \115  | \23 ,
  \[38]  = \117  | \24 ,
  \100  = (\[61]  & (\135  & \33 )) | ((\[34]  & ~\137 ) | (~\137  & \33 )),
  \101  = (\[62]  & (\137  & \34 )) | ((\[35]  & ~\86 ) | (~\86  & \34 )),
  \102  = (~\140  & \2 ) | (\140  & ~\2 ),
  \107  = (~\[47]  & ~\140 ) | (\140  & \2 ),
  \[39]  = \119  | \25 ,
  \113  = (\[60]  & \4 ) | (\[33]  & \21 ),
  \115  = (\[36]  & (\5  & \1 )) | (\113  & \22 ),
  \117  = (\[37]  & (\6  & \1 )) | (\115  & \23 ),
  \119  = (\[38]  & (\7  & \1 )) | (\117  & \24 ),
  \[20]  = \90 ,
  \121  = (\[39]  & (\8  & \1 )) | (\119  & \25 ),
  \123  = (\[40]  & (\9  & \1 )) | (\121  & \26 ),
  \125  = (\[41]  & (\10  & \1 )) | (\123  & \27 ),
  \127  = (\[42]  & (\11  & \1 )) | (\125  & \28 ),
  \129  = (\[43]  & (\12  & \1 )) | (\127  & \29 ),
  \[21]  = \91 ,
  \131  = (\[44]  & (\13  & \1 )) | (\129  & \30 ),
  \133  = (\[45]  & (\14  & \1 )) | (\131  & \31 ),
  \135  = (\[46]  & (\15  & \1 )) | (\133  & \32 ),
  \137  = (\[61]  & \135 ) | (\[34]  & \33 ),
  \[22]  = \92 ,
  \140  = (~\[47]  & ~\86 ) | (\[47]  & \86 ),
  \[23]  = \93 ,
  \[24]  = \94 ,
  \[25]  = \95 ;
always begin
  \20  = \[18] ;
  \21  = \[19] ;
  \22  = \[20] ;
  \23  = \[21] ;
  \24  = \[22] ;
  \25  = \[23] ;
  \26  = \[24] ;
  \27  = \[25] ;
  \28  = \[26] ;
  \29  = \[27] ;
  \30  = \[28] ;
  \31  = \[29] ;
  \32  = \[30] ;
  \33  = \[31] ;
  \34  = \[32] ;
  \2  = \[17] ;
end
initial begin
  \20  = 0;
  \21  = 0;
  \22  = 0;
  \23  = 0;
  \24  = 0;
  \25  = 0;
  \26  = 0;
  \27  = 0;
  \28  = 0;
  \29  = 0;
  \30  = 0;
  \31  = 0;
  \32  = 0;
  \33  = 0;
  \34  = 0;
  \2  = 0;
end
endmodule

