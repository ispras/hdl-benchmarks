//NOTE: no-implementation module stub

module NAND4X1 (
    input wire A,
    input wire B,
    input wire C,
    input wire D,
    output wire Y
);

endmodule

module INVX1 (
    input wire A,
    output wire Y
);

endmodule

module DFFSRX1 (
    input wire RN,
    input wire SN,
    input wire CK,
    input wire D,
    output wire Q,
    output wire QN
);

endmodule

module OAI21X1 (
    input wire A0,
    input wire A1,
    input wire B0,
    output wire Y
);

endmodule

module AOI22X1 (
    input wire A0,
    input wire A1,
    input wire B0,
    input wire B1,
    output wire Y
);

endmodule

module NAND3X1 (
    input wire A,
    input wire B,
    input wire C,
    output wire Y
);

endmodule

module NAND2X1 (
    input wire A,
    input wire B,
    output wire Y
);

endmodule

module AOI21X1 (
    input wire A0,
    input wire A1,
    input wire B0,
    output wire Y
);

endmodule

module OR2X1 (
    input wire A,
    input wire B,
    output wire Y
);

endmodule

module INVX2 (
    input wire A,
    output wire Y
);

endmodule

module OAI22X1 (
    input wire A0,
    input wire A1,
    input wire B0,
    input wire B1,
    output wire Y
);

endmodule

module NOR2X1 (
    input wire A,
    input wire B,
    output wire Y
);

endmodule

module NAND2X2 (
    input wire A,
    input wire B,
    output wire Y
);

endmodule

module AND2X1 (
    input wire A,
    input wire B,
    output wire Y
);

endmodule

module CLKBUFX3 (
    input wire A,
    output wire Y
);

endmodule

module MX2X1 (
    input wire A,
    input wire B,
    input wire S0,
    output wire Y
);

endmodule

module CLKBUFX1 (
    input wire A,
    output wire Y
);

endmodule

module INVX4 (
    input wire A,
    output wire Y
);

endmodule

module CLKBUFX2 (
    input wire A,
    output wire Y
);

endmodule

module INVX8 (
    input wire A,
    output wire Y
);

endmodule

module BUFX3 (
    input wire A,
    output wire Y
);

endmodule

module XOR2X1 (
    input wire A,
    input wire B,
    output wire Y
);

endmodule

module OR4X1 (
    input wire A,
    input wire B,
    input wire C,
    input wire D,
    output wire Y
);

endmodule

module ADDHX1 (
    input wire A,
    input wire B,
    output wire CO,
    output wire S
);

endmodule

module NOR3X1 (
    input wire A,
    input wire B,
    input wire C,
    output wire Y
);

endmodule

module OAI33X1 (
    input wire A0,
    input wire A1,
    input wire A2,
    input wire B0,
    input wire B1,
    input wire B2,
    output wire Y
);

endmodule

module BUFX1 (
    input wire A,
    output wire Y
);

endmodule

module SDFFSRX1 (
    input wire RN,
    input wire SN,
    input wire CK,
    input wire D,
    input wire SE,
    input wire SI,
    output wire Q,
    output wire QN
);

endmodule
