module sub_2_6_1(a, b, c);
  input [1:0] a;
  input [5:0] b;
  output c;
  assign c = a - b;
endmodule
