// IWLS benchmark module "i5" printed on Wed May 29 17:26:46 2002
module i5(\V4(0) , \V2(1) , \V4(1) , \V2(0) , \V28(1) , \V16(2) , \V28(2) , \V16(3) , \V28(3) , \V28(5) , \V16(6) , \V28(6) , \V16(7) , \V28(7) , \V28(9) , \V16(10) , \V28(10) , \V16(11) , \V28(11) , \V28(13) , \V16(14) , \V28(14) , \V16(15) , \V28(15) , \V16(1) , \V16(5) , \V16(9) , \V16(13) , \V52(1) , \V40(2) , \V52(2) , \V40(3) , \V52(3) , \V52(5) , \V40(6) , \V52(6) , \V40(7) , \V52(7) , \V52(9) , \V40(10) , \V52(10) , \V40(11) , \V52(11) , \V52(13) , \V40(14) , \V52(14) , \V40(15) , \V52(15) , \V40(1) , \V40(5) , \V40(9) , \V40(13) , \V76(1) , \V64(2) , \V76(2) , \V64(3) , \V76(3) , \V76(5) , \V64(6) , \V76(6) , \V64(7) , \V76(7) , \V76(9) , \V64(10) , \V76(10) , \V64(11) , \V76(11) , \V76(13) , \V64(14) , \V76(14) , \V64(15) , \V76(15) , \V64(1) , \V64(5) , \V64(9) , \V64(13) , \V100(1) , \V88(2) , \V100(2) , \V88(3) , \V100(3) , \V100(5) , \V88(6) , \V100(6) , \V88(7) , \V100(7) , \V100(9) , \V88(10) , \V100(10) , \V88(11) , \V100(11) , \V100(13) , \V88(14) , \V100(14) , \V88(15) , \V133(0) , \V100(15) , \V88(1) , \V88(5) , \V88(9) , \V88(13) , \V106(1) , \V103(2) , \V106(2) , \V103(3) , \V106(3) , \V112(1) , \V109(2) , \V112(2) , \V109(3) , \V112(3) , \V118(1) , \V115(2) , \V118(2) , \V115(3) , \V118(3) , \V124(1) , \V121(2) , \V124(2) , \V121(3) , \V124(3) , \V103(1) , \V109(1) , \V115(1) , \V121(1) , \V132(0) , \V128(1) , \V132(1) , \V128(2) , \V132(2) , \V128(3) , \V132(3) , \V128(0) , \V135(0) , \V135(1) , \V151(1) , \V151(2) , \V151(3) , \V151(5) , \V151(6) , \V151(7) , \V151(9) , \V151(10) , \V151(11) , \V151(13) , \V151(14) , \V151(15) , \V167(1) , \V167(2) , \V167(3) , \V167(5) , \V167(6) , \V167(7) , \V167(9) , \V167(10) , \V167(11) , \V167(13) , \V167(14) , \V167(15) , \V183(1) , \V183(2) , \V183(3) , \V183(5) , \V183(6) , \V183(7) , \V183(9) , \V183(10) , \V183(11) , \V183(13) , \V183(14) , \V183(15) , \V199(1) , \V199(2) , \V199(3) , \V199(5) , \V199(6) , \V199(7) , \V199(9) , \V199(10) , \V199(11) , \V199(13) , \V199(14) , \V199(15) , \V151(4) , \V151(8) , \V151(12) , \V167(4) , \V167(8) , \V167(12) , \V183(4) , \V183(8) , \V183(12) , \V199(4) , \V199(8) , \V199(12) , \V151(0) , \V167(0) , \V183(0) , \V199(0) );
input
  \V124(2) ,
  \V40(3) ,
  \V88(11) ,
  \V40(5) ,
  \V88(10) ,
  \V40(6) ,
  \V40(7) ,
  \V124(1) ,
  \V40(9) ,
  \V112(3) ,
  \V112(2) ,
  \V112(1) ,
  \V40(13) ,
  \V40(15) ,
  \V40(14) ,
  \V100(3) ,
  \V100(2) ,
  \V100(5) ,
  \V40(11) ,
  \V40(10) ,
  \V128(3) ,
  \V100(1) ,
  \V128(2) ,
  \V115(3) ,
  \V115(2) ,
  \V128(1) ,
  \V100(7) ,
  \V128(0) ,
  \V76(13) ,
  \V100(6) ,
  \V100(9) ,
  \V76(15) ,
  \V115(1) ,
  \V76(14) ,
  \V76(11) ,
  \V103(3) ,
  \V76(10) ,
  \V103(2) ,
  \V103(1) ,
  \V2(0) ,
  \V2(1) ,
  \V118(3) ,
  \V118(2) ,
  \V118(1) ,
  \V106(3) ,
  \V4(0) ,
  \V106(2) ,
  \V100(11) ,
  \V4(1) ,
  \V100(10) ,
  \V100(13) ,
  \V100(15) ,
  \V106(1) ,
  \V100(14) ,
  \V28(13) ,
  \V28(15) ,
  \V28(14) ,
  \V64(13) ,
  \V28(11) ,
  \V64(15) ,
  \V28(10) ,
  \V64(14) ,
  \V64(11) ,
  \V64(10) ,
  \V109(3) ,
  \V109(2) ,
  \V109(1) ,
  \V88(1) ,
  \V88(2) ,
  \V88(3) ,
  \V88(5) ,
  \V88(6) ,
  \V132(3) ,
  \V88(7) ,
  \V132(2) ,
  \V88(9) ,
  \V76(1) ,
  \V76(2) ,
  \V132(1) ,
  \V28(1) ,
  \V76(3) ,
  \V132(0) ,
  \V28(2) ,
  \V28(3) ,
  \V76(5) ,
  \V76(6) ,
  \V28(5) ,
  \V76(7) ,
  \V28(6) ,
  \V16(13) ,
  \V28(7) ,
  \V76(9) ,
  \V133(0) ,
  \V16(15) ,
  \V28(9) ,
  \V64(1) ,
  \V16(14) ,
  \V64(2) ,
  \V52(13) ,
  \V121(3) ,
  \V16(1) ,
  \V64(3) ,
  \V121(2) ,
  \V16(2) ,
  \V16(11) ,
  \V52(15) ,
  \V16(3) ,
  \V64(5) ,
  \V16(10) ,
  \V52(14) ,
  \V64(6) ,
  \V16(5) ,
  \V64(7) ,
  \V16(6) ,
  \V52(11) ,
  \V121(1) ,
  \V16(7) ,
  \V64(9) ,
  \V52(10) ,
  \V16(9) ,
  \V52(1) ,
  \V52(2) ,
  \V52(3) ,
  \V52(5) ,
  \V52(6) ,
  \V52(7) ,
  \V88(13) ,
  \V52(9) ,
  \V88(15) ,
  \V40(1) ,
  \V88(14) ,
  \V124(3) ,
  \V40(2) ;
output
  \V199(1) ,
  \V199(0) ,
  \V199(7) ,
  \V199(6) ,
  \V199(9) ,
  \V199(8) ,
  \V151(3) ,
  \V151(2) ,
  \V151(5) ,
  \V151(4) ,
  \V151(1) ,
  \V151(0) ,
  \V151(7) ,
  \V151(6) ,
  \V151(9) ,
  \V151(8) ,
  \V167(3) ,
  \V167(2) ,
  \V167(5) ,
  \V167(4) ,
  \V167(1) ,
  \V167(0) ,
  \V199(11) ,
  \V167(7) ,
  \V199(10) ,
  \V167(6) ,
  \V199(13) ,
  \V183(11) ,
  \V167(9) ,
  \V199(12) ,
  \V183(10) ,
  \V167(8) ,
  \V199(15) ,
  \V183(13) ,
  \V199(14) ,
  \V183(12) ,
  \V183(15) ,
  \V183(14) ,
  \V167(11) ,
  \V167(10) ,
  \V167(13) ,
  \V151(11) ,
  \V167(12) ,
  \V151(10) ,
  \V167(15) ,
  \V151(13) ,
  \V167(14) ,
  \V151(12) ,
  \V151(15) ,
  \V151(14) ,
  \V183(3) ,
  \V183(2) ,
  \V183(5) ,
  \V183(4) ,
  \V183(1) ,
  \V183(0) ,
  \V135(1) ,
  \V135(0) ,
  \V183(7) ,
  \V183(6) ,
  \V183(9) ,
  \V183(8) ,
  \V199(3) ,
  \V199(2) ,
  \V199(5) ,
  \V199(4) ;
wire
  \[60] ,
  \[61] ,
  \[62] ,
  \[63] ,
  \[64] ,
  \[65] ,
  \[0] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \[5] ,
  \[6] ,
  \[7] ,
  \[8] ,
  \[9] ,
  V200,
  V201,
  V202,
  V203,
  V204,
  V205,
  V206,
  V207,
  V208,
  V209,
  V210,
  V211,
  V212,
  V213,
  V214,
  V215,
  V216,
  V217,
  V218,
  V219,
  V220,
  V221,
  V222,
  V223,
  V224,
  V225,
  V226,
  V227,
  V228,
  V229,
  V230,
  V231,
  V232,
  V233,
  V234,
  V235,
  V236,
  V237,
  V238,
  V239,
  V240,
  V241,
  V242,
  V243,
  V244,
  V245,
  V246,
  V247,
  V248,
  V249,
  V250,
  V251,
  V252,
  V253,
  V254,
  V255,
  V256,
  V257,
  V258,
  V259,
  V260,
  V261,
  V262,
  V263,
  V264,
  V265,
  V266,
  V267,
  V268,
  V269,
  V270,
  V271,
  V272,
  V273,
  V274,
  V275,
  V276,
  V277,
  V278,
  V279,
  V280,
  V281,
  V282,
  V283,
  V284,
  V285,
  V286,
  V287,
  V288,
  V289,
  V290,
  V291,
  V292,
  V293,
  V294,
  V295,
  V296,
  V297,
  V298,
  V299,
  V300,
  V301,
  V302,
  V303,
  V304,
  V305,
  V306,
  V307,
  V308,
  V309,
  V310,
  V311,
  V312,
  V313,
  V314,
  V315,
  V316,
  V317,
  V318,
  V319,
  V320,
  V321,
  V322,
  V323,
  V324,
  V325,
  V326,
  V327,
  V328,
  V329,
  \[10] ,
  V330,
  V331,
  V332,
  \[11] ,
  \[12] ,
  \[13] ,
  \[14] ,
  \[15] ,
  \[16] ,
  \[17] ,
  \[18] ,
  \[19] ,
  \[20] ,
  \[21] ,
  \[22] ,
  \[23] ,
  \[24] ,
  \[25] ,
  \[26] ,
  \[27] ,
  \[28] ,
  \[29] ,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \[36] ,
  \[37] ,
  \[38] ,
  \[39] ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ,
  \[59] ;
assign
  \[60]  = V320 | (\V121(2)  | V321),
  \[61]  = \V121(3)  | V322,
  \[62]  = V325 | (V323 | (\V128(0)  | (V324 | V326))),
  \V199(1)  = \[38] ,
  \[63]  = V328 | (\V128(1)  | (V327 | V329)),
  \V199(0)  = \[65] ,
  \[64]  = V330 | (\V128(2)  | V331),
  \[65]  = \V128(3)  | V332,
  \V199(7)  = \[43] ,
  \V199(6)  = \[42] ,
  \V199(9)  = \[44] ,
  \V199(8)  = \[60] ,
  \[0]  = V200 | (\V2(0)  | V201),
  \[1]  = \V2(1)  | V202,
  \[2]  = V204 | (\V16(1)  | (V203 | V205)),
  \[3]  = V206 | (\V16(2)  | V207),
  \[4]  = \V16(3)  | V208,
  \[5]  = V210 | (\V16(5)  | (V209 | V211)),
  \[6]  = V212 | (\V16(6)  | V213),
  \[7]  = \V16(7)  | V214,
  \[8]  = V216 | (\V16(9)  | (V215 | V217)),
  \[9]  = V218 | (\V16(10)  | V219),
  V200 = \V2(1)  & \V4(0) ,
  V201 = \V4(1)  & (\V4(0)  & \[62] ),
  V202 = \V4(1)  & \[62] ,
  V203 = \V16(2)  & \V28(1) ,
  V204 = \V28(1)  & (\V16(3)  & \V28(2) ),
  V205 = \V28(3)  & (\V28(1)  & (\V28(2)  & \[50] )),
  V206 = \V16(3)  & \V28(2) ,
  V207 = \V28(3)  & (\V28(2)  & \[50] ),
  V208 = \V28(3)  & \[50] ,
  V209 = \V16(6)  & \V28(5) ,
  V210 = \V28(5)  & (\V16(7)  & \V28(6) ),
  V211 = \V28(7)  & (\V28(5)  & (\V28(6)  & \[51] )),
  V212 = \V16(7)  & \V28(6) ,
  V213 = \V28(7)  & (\V28(6)  & \[51] ),
  V214 = \V28(7)  & \[51] ,
  V215 = \V16(10)  & \V28(9) ,
  V216 = \V28(9)  & (\V16(11)  & \V28(10) ),
  V217 = \V28(11)  & (\V28(9)  & (\V28(10)  & \[52] )),
  V218 = \V16(11)  & \V28(10) ,
  V219 = \V28(11)  & (\V28(10)  & \[52] ),
  V220 = \V28(11)  & \[52] ,
  V221 = \V16(14)  & \V28(13) ,
  V222 = \V28(13)  & (\V16(15)  & \V28(14) ),
  V223 = \V28(15)  & (\V28(13)  & (\V28(14)  & \[63] )),
  V224 = \V16(15)  & \V28(14) ,
  V225 = \V28(15)  & (\V28(14)  & \[63] ),
  V226 = \V28(15)  & \[63] ,
  V227 = \V40(2)  & \V52(1) ,
  V228 = \V52(1)  & (\V40(3)  & \V52(2) ),
  V229 = \V52(3)  & (\V52(1)  & (\V52(2)  & \[53] )),
  V230 = \V40(3)  & \V52(2) ,
  V231 = \V52(3)  & (\V52(2)  & \[53] ),
  V232 = \V52(3)  & \[53] ,
  V233 = \V40(6)  & \V52(5) ,
  V234 = \V52(5)  & (\V40(7)  & \V52(6) ),
  V235 = \V52(7)  & (\V52(5)  & (\V52(6)  & \[54] )),
  V236 = \V40(7)  & \V52(6) ,
  V237 = \V52(7)  & (\V52(6)  & \[54] ),
  V238 = \V52(7)  & \[54] ,
  V239 = \V40(10)  & \V52(9) ,
  V240 = \V52(9)  & (\V40(11)  & \V52(10) ),
  V241 = \V52(11)  & (\V52(9)  & (\V52(10)  & \[55] )),
  V242 = \V40(11)  & \V52(10) ,
  V243 = \V52(11)  & (\V52(10)  & \[55] ),
  V244 = \V52(11)  & \[55] ,
  V245 = \V40(14)  & \V52(13) ,
  V246 = \V52(13)  & (\V40(15)  & \V52(14) ),
  V247 = \V52(15)  & (\V52(13)  & (\V52(14)  & \[64] )),
  V248 = \V40(15)  & \V52(14) ,
  V249 = \V52(15)  & (\V52(14)  & \[64] ),
  V250 = \V52(15)  & \[64] ,
  V251 = \V64(2)  & \V76(1) ,
  V252 = \V76(1)  & (\V64(3)  & \V76(2) ),
  V253 = \V76(3)  & (\V76(1)  & (\V76(2)  & \[56] )),
  V254 = \V64(3)  & \V76(2) ,
  V255 = \V76(3)  & (\V76(2)  & \[56] ),
  V256 = \V76(3)  & \[56] ,
  V257 = \V64(6)  & \V76(5) ,
  V258 = \V76(5)  & (\V64(7)  & \V76(6) ),
  V259 = \V76(7)  & (\V76(5)  & (\V76(6)  & \[57] )),
  V260 = \V64(7)  & \V76(6) ,
  V261 = \V76(7)  & (\V76(6)  & \[57] ),
  V262 = \V76(7)  & \[57] ,
  V263 = \V64(10)  & \V76(9) ,
  V264 = \V76(9)  & (\V64(11)  & \V76(10) ),
  V265 = \V76(11)  & (\V76(9)  & (\V76(10)  & \[58] )),
  V266 = \V64(11)  & \V76(10) ,
  V267 = \V76(11)  & (\V76(10)  & \[58] ),
  V268 = \V76(11)  & \[58] ,
  V269 = \V64(14)  & \V76(13) ,
  V270 = \V76(13)  & (\V64(15)  & \V76(14) ),
  V271 = \V76(15)  & (\V76(13)  & (\V76(14)  & \[65] )),
  V272 = \V64(15)  & \V76(14) ,
  V273 = \V76(15)  & (\V76(14)  & \[65] ),
  V274 = \V76(15)  & \[65] ,
  V275 = \V88(2)  & \V100(1) ,
  V276 = \V100(1)  & (\V88(3)  & \V100(2) ),
  V277 = \V100(3)  & (\V100(1)  & (\V100(2)  & \[59] )),
  V278 = \V88(3)  & \V100(2) ,
  V279 = \V100(3)  & (\V100(2)  & \[59] ),
  V280 = \V100(3)  & \[59] ,
  V281 = \V88(6)  & \V100(5) ,
  V282 = \V100(5)  & (\V88(7)  & \V100(6) ),
  V283 = \V100(7)  & (\V100(5)  & (\V100(6)  & \[60] )),
  V284 = \V88(7)  & \V100(6) ,
  V285 = \V100(7)  & (\V100(6)  & \[60] ),
  V286 = \V100(7)  & \[60] ,
  V287 = \V88(10)  & \V100(9) ,
  V288 = \V100(9)  & (\V88(11)  & \V100(10) ),
  V289 = \V100(11)  & (\V100(9)  & (\V100(10)  & \[61] )),
  V290 = \V88(11)  & \V100(10) ,
  V291 = \V100(11)  & (\V100(10)  & \[61] ),
  V292 = \V100(11)  & \[61] ,
  V293 = \V88(14)  & \V100(13) ,
  V294 = \V100(13)  & (\V88(15)  & \V100(14) ),
  V295 = \V100(15)  & (\V100(13)  & (\V100(14)  & \V133(0) )),
  V296 = \V88(15)  & \V100(14) ,
  V297 = \V100(15)  & (\V100(14)  & \V133(0) ),
  V298 = \V100(15)  & \V133(0) ,
  V299 = \V103(2)  & \V106(1) ,
  \V151(3)  = \[4] ,
  \V151(2)  = \[3] ,
  \V151(5)  = \[5] ,
  \V151(4)  = \[50] ,
  V300 = \V106(1)  & (\V103(3)  & \V106(2) ),
  V301 = \V106(3)  & (\V106(1)  & (\V106(2)  & \[63] )),
  V302 = \V103(3)  & \V106(2) ,
  V303 = \V106(3)  & (\V106(2)  & \[63] ),
  V304 = \V106(3)  & \[63] ,
  V305 = \V109(2)  & \V112(1) ,
  V306 = \V112(1)  & (\V109(3)  & \V112(2) ),
  V307 = \V112(3)  & (\V112(1)  & (\V112(2)  & \[64] )),
  V308 = \V109(3)  & \V112(2) ,
  V309 = \V112(3)  & (\V112(2)  & \[64] ),
  \V151(1)  = \[2] ,
  V310 = \V112(3)  & \[64] ,
  V311 = \V115(2)  & \V118(1) ,
  V312 = \V118(1)  & (\V115(3)  & \V118(2) ),
  V313 = \V118(3)  & (\V118(1)  & (\V118(2)  & \[65] )),
  V314 = \V115(3)  & \V118(2) ,
  V315 = \V118(3)  & (\V118(2)  & \[65] ),
  V316 = \V118(3)  & \[65] ,
  V317 = \V121(2)  & \V124(1) ,
  V318 = \V124(1)  & (\V121(3)  & \V124(2) ),
  V319 = \V124(3)  & (\V124(1)  & (\V124(2)  & \V133(0) )),
  \V151(0)  = \[62] ,
  V320 = \V121(3)  & \V124(2) ,
  V321 = \V124(3)  & (\V124(2)  & \V133(0) ),
  V322 = \V124(3)  & \V133(0) ,
  V323 = \V128(1)  & \V132(0) ,
  V324 = \V132(0)  & (\V128(2)  & \V132(1) ),
  V325 = \V132(1)  & (\V128(3)  & (\V132(0)  & \V132(2) )),
  V326 = \V132(3)  & (\V132(1)  & (\V132(0)  & (\V132(2)  & \V133(0) ))),
  V327 = \V128(2)  & \V132(1) ,
  V328 = \V132(1)  & (\V128(3)  & \V132(2) ),
  V329 = \V132(3)  & (\V132(1)  & (\V132(2)  & \V133(0) )),
  \[10]  = \V16(11)  | V220,
  V330 = \V128(3)  & \V132(2) ,
  V331 = \V132(3)  & (\V132(2)  & \V133(0) ),
  V332 = \V132(3)  & \V133(0) ,
  \[11]  = V222 | (\V16(13)  | (V221 | V223)),
  \[12]  = V224 | (\V16(14)  | V225),
  \[13]  = \V16(15)  | V226,
  \[14]  = V228 | (\V40(1)  | (V227 | V229)),
  \V151(7)  = \[7] ,
  \[15]  = V230 | (\V40(2)  | V231),
  \V151(6)  = \[6] ,
  \[16]  = \V40(3)  | V232,
  \V151(9)  = \[8] ,
  \[17]  = V234 | (\V40(5)  | (V233 | V235)),
  \V151(8)  = \[51] ,
  \V167(3)  = \[16] ,
  \[18]  = V236 | (\V40(6)  | V237),
  \V167(2)  = \[15] ,
  \[19]  = \V40(7)  | V238,
  \V167(5)  = \[17] ,
  \V167(4)  = \[53] ,
  \V167(1)  = \[14] ,
  \V167(0)  = \[63] ,
  \[20]  = V240 | (\V40(9)  | (V239 | V241)),
  \[21]  = V242 | (\V40(10)  | V243),
  \[22]  = \V40(11)  | V244,
  \V199(11)  = \[46] ,
  \[23]  = V246 | (\V40(13)  | (V245 | V247)),
  \V167(7)  = \[19] ,
  \V199(10)  = \[45] ,
  \[24]  = V248 | (\V40(14)  | V249),
  \V167(6)  = \[18] ,
  \V199(13)  = \[47] ,
  \[25]  = \V40(15)  | V250,
  \V183(11)  = \[34] ,
  \V167(9)  = \[20] ,
  \V199(12)  = \[61] ,
  \[26]  = V252 | (\V64(1)  | (V251 | V253)),
  \V183(10)  = \[33] ,
  \V167(8)  = \[54] ,
  \V199(15)  = \[49] ,
  \[27]  = V254 | (\V64(2)  | V255),
  \V183(13)  = \[35] ,
  \V199(14)  = \[48] ,
  \[28]  = \V64(3)  | V256,
  \V183(12)  = \[58] ,
  \[29]  = V258 | (\V64(5)  | (V257 | V259)),
  \V183(15)  = \[37] ,
  \V183(14)  = \[36] ,
  \[30]  = V260 | (\V64(6)  | V261),
  \[31]  = \V64(7)  | V262,
  \[32]  = V264 | (\V64(9)  | (V263 | V265)),
  \[33]  = V266 | (\V64(10)  | V267),
  \[34]  = \V64(11)  | V268,
  \V167(11)  = \[22] ,
  \[35]  = V270 | (\V64(13)  | (V269 | V271)),
  \V167(10)  = \[21] ,
  \[36]  = V272 | (\V64(14)  | V273),
  \V167(13)  = \[23] ,
  \V151(11)  = \[10] ,
  \[37]  = \V64(15)  | V274,
  \V167(12)  = \[55] ,
  \V151(10)  = \[9] ,
  \[38]  = V276 | (\V88(1)  | (V275 | V277)),
  \V167(15)  = \[25] ,
  \V151(13)  = \[11] ,
  \[39]  = V278 | (\V88(2)  | V279),
  \V167(14)  = \[24] ,
  \V151(12)  = \[52] ,
  \V151(15)  = \[13] ,
  \V151(14)  = \[12] ,
  \[40]  = \V88(3)  | V280,
  \[41]  = V282 | (\V88(5)  | (V281 | V283)),
  \[42]  = V284 | (\V88(6)  | V285),
  \[43]  = \V88(7)  | V286,
  \[44]  = V288 | (\V88(9)  | (V287 | V289)),
  \[45]  = V290 | (\V88(10)  | V291),
  \[46]  = \V88(11)  | V292,
  \[47]  = V294 | (\V88(13)  | (V293 | V295)),
  \[48]  = V296 | (\V88(14)  | V297),
  \[49]  = \V88(15)  | V298,
  \V183(3)  = \[28] ,
  \V183(2)  = \[27] ,
  \V183(5)  = \[29] ,
  \[50]  = V300 | (\V103(1)  | (V299 | V301)),
  \V183(4)  = \[56] ,
  \[51]  = V302 | (\V103(2)  | V303),
  \[52]  = \V103(3)  | V304,
  \[53]  = V306 | (\V109(1)  | (V305 | V307)),
  \V183(1)  = \[26] ,
  \[54]  = V308 | (\V109(2)  | V309),
  \V183(0)  = \[64] ,
  \[55]  = \V109(3)  | V310,
  \V135(1)  = \[1] ,
  \[56]  = V312 | (\V115(1)  | (V311 | V313)),
  \V135(0)  = \[0] ,
  \[57]  = V314 | (\V115(2)  | V315),
  \[58]  = \V115(3)  | V316,
  \[59]  = V318 | (\V121(1)  | (V317 | V319)),
  \V183(7)  = \[31] ,
  \V183(6)  = \[30] ,
  \V183(9)  = \[32] ,
  \V183(8)  = \[57] ,
  \V199(3)  = \[40] ,
  \V199(2)  = \[39] ,
  \V199(5)  = \[41] ,
  \V199(4)  = \[59] ;
endmodule

