// IWLS benchmark module "i9" printed on Wed May 29 17:27:10 2002
module i9(\V9(3) , \V9(1) , \V9(2) , \V9(10) , \V9(0) , \V9(5) , \V9(6) , \V9(7) , \V9(8) , \V56(31) , \V56(30) , \V56(29) , \V56(28) , \V56(27) , \V56(26) , \V56(25) , \V56(24) , \V56(23) , \V56(22) , \V56(21) , \V56(20) , \V56(19) , \V56(18) , \V56(17) , \V56(16) , \V56(15) , \V56(14) , \V56(13) , \V56(12) , \V56(11) , \V56(10) , \V56(9) , \V56(8) , \V56(7) , \V56(6) , \V56(5) , \V56(4) , \V56(3) , \V56(2) , \V56(1) , \V56(0) , \V88(11) , \V88(10) , \V88(9) , \V88(8) , \V88(7) , \V88(6) , \V88(5) , \V88(4) , \V88(3) , \V88(2) , \V88(1) , \V24(14) , \V24(13) , \V24(12) , \V24(11) , \V24(10) , \V24(9) , \V24(8) , \V24(7) , \V24(6) , \V24(5) , \V24(4) , \V24(3) , \V24(2) , \V24(1) , \V24(0) , \V88(31) , \V88(30) , \V88(29) , \V88(28) , \V88(27) , \V88(26) , \V88(25) , \V88(24) , \V88(23) , \V88(22) , \V88(21) , \V88(20) , \V88(19) , \V88(18) , \V88(17) , \V88(16) , \V88(15) , \V88(14) , \V88(13) , \V88(12) , \V88(0) , \V119(30) , \V119(29) , \V119(28) , \V119(27) , \V119(26) , \V119(25) , \V119(24) , \V119(23) , \V119(22) , \V119(21) , \V119(20) , \V119(19) , \V119(18) , \V119(17) , \V119(16) , \V119(15) , \V119(14) , \V119(13) , \V119(12) , \V119(11) , \V119(10) , \V119(9) , \V119(8) , \V119(7) , \V119(6) , \V119(5) , \V119(4) , \V119(3) , \V119(2) , \V119(1) , \V119(0) , \V151(15) , \V151(14) , \V151(13) , \V151(12) , \V151(11) , \V151(10) , \V151(9) , \V151(8) , \V151(7) , \V151(6) , \V151(5) , \V151(4) , \V151(3) , \V151(2) , \V151(1) , \V151(0) , \V151(31) , \V151(30) , \V151(29) , \V151(28) , \V151(27) , \V151(26) , \V151(25) , \V151(24) , \V151(23) , \V151(22) , \V151(21) , \V151(20) , \V151(19) , \V151(18) , \V151(17) , \V151(16) );
input
  \V88(21) ,
  \V88(20) ,
  \V88(27) ,
  \V9(0) ,
  \V88(0) ,
  \V88(26) ,
  \V9(1) ,
  \V88(1) ,
  \V88(29) ,
  \V9(2) ,
  \V88(2) ,
  \V88(28) ,
  \V9(3) ,
  \V88(3) ,
  \V88(4) ,
  \V9(5) ,
  \V88(5) ,
  \V9(6) ,
  \V88(6) ,
  \V56(13) ,
  \V9(7) ,
  \V88(7) ,
  \V56(12) ,
  \V9(8) ,
  \V9(10) ,
  \V88(8) ,
  \V56(15) ,
  \V88(9) ,
  \V88(31) ,
  \V56(14) ,
  \V88(30) ,
  \V56(11) ,
  \V56(10) ,
  \V56(17) ,
  \V56(0) ,
  \V56(16) ,
  \V56(1) ,
  \V56(19) ,
  \V56(2) ,
  \V56(18) ,
  \V56(3) ,
  \V56(23) ,
  \V56(4) ,
  \V56(22) ,
  \V56(5) ,
  \V56(25) ,
  \V56(6) ,
  \V56(24) ,
  \V56(7) ,
  \V56(8) ,
  \V56(9) ,
  \V56(21) ,
  \V56(20) ,
  \V56(27) ,
  \V56(26) ,
  \V56(29) ,
  \V56(28) ,
  \V24(0) ,
  \V88(13) ,
  \V24(1) ,
  \V88(12) ,
  \V24(2) ,
  \V88(15) ,
  \V24(3) ,
  \V24(13) ,
  \V88(14) ,
  \V24(4) ,
  \V24(12) ,
  \V24(5) ,
  \V56(31) ,
  \V24(6) ,
  \V24(14) ,
  \V88(11) ,
  \V56(30) ,
  \V24(7) ,
  \V88(10) ,
  \V24(8) ,
  \V24(9) ,
  \V24(11) ,
  \V24(10) ,
  \V88(17) ,
  \V88(16) ,
  \V88(19) ,
  \V88(18) ,
  \V88(23) ,
  \V88(22) ,
  \V88(25) ,
  \V88(24) ;
output
  \V119(21) ,
  \V151(16) ,
  \V119(20) ,
  \V151(19) ,
  \V119(23) ,
  \V151(18) ,
  \V119(22) ,
  \V119(25) ,
  \V119(24) ,
  \V119(17) ,
  \V119(16) ,
  \V119(3) ,
  \V119(19) ,
  \V119(2) ,
  \V119(18) ,
  \V151(11) ,
  \V119(5) ,
  \V151(10) ,
  \V119(4) ,
  \V151(13) ,
  \V151(12) ,
  \V151(15) ,
  \V119(1) ,
  \V151(14) ,
  \V119(0) ,
  \V119(11) ,
  \V119(10) ,
  \V119(13) ,
  \V119(12) ,
  \V119(7) ,
  \V119(15) ,
  \V119(6) ,
  \V119(14) ,
  \V119(9) ,
  \V119(8) ,
  \V151(3) ,
  \V151(2) ,
  \V151(5) ,
  \V151(4) ,
  \V151(1) ,
  \V151(0) ,
  \V151(7) ,
  \V151(6) ,
  \V151(9) ,
  \V151(8) ,
  \V151(31) ,
  \V151(30) ,
  \V119(30) ,
  \V151(27) ,
  \V151(26) ,
  \V151(29) ,
  \V151(28) ,
  \V119(27) ,
  \V119(26) ,
  \V119(29) ,
  \V119(28) ,
  \V151(21) ,
  \V151(20) ,
  \V151(23) ,
  \V151(22) ,
  \V151(25) ,
  \V151(24) ,
  \V151(17) ;
wire
  \[59] ,
  \[15] ,
  \[16] ,
  \[17] ,
  \[18] ,
  \[19] ,
  \[60] ,
  \[61] ,
  \[62] ,
  \[0] ,
  \[63] ,
  \[1] ,
  \[64] ,
  \[20] ,
  \[2] ,
  \[65] ,
  \[21] ,
  \[3] ,
  \[66] ,
  \[22] ,
  \[4] ,
  \[67] ,
  \[23] ,
  \[5] ,
  \[68] ,
  \[24] ,
  \[6] ,
  \[69] ,
  \[25] ,
  \[7] ,
  \[26] ,
  \[8] ,
  \[27] ,
  \[9] ,
  \[28] ,
  \[29] ,
  \[71] ,
  V207,
  \[72] ,
  \[73] ,
  \[74] ,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \[36] ,
  \[37] ,
  \[38] ,
  \[39] ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \V174(2) ,
  \V174(1) ,
  \[50] ,
  \V174(0) ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[10] ,
  \[55] ,
  \[11] ,
  \[56] ,
  \[12] ,
  \[57] ,
  \[13] ,
  \[58] ,
  \[14] ;
assign
  \[59]  = (\[65]  & \V88(4) ) | ((\[64]  & \V88(19) ) | ((V207 & \V88(11) ) | \[74] )),
  \[15]  = (\[67]  & \V56(1) ) | ((~\[66]  & \V56(16) ) | ((\[63]  & \V56(5) ) | ((V207 & \V56(8) ) | ~\V174(0) ))),
  \V119(21)  = \[9] ,
  \V151(16)  = \[62] ,
  \[16]  = (\[67]  & \V24(14) ) | ((~\[66]  & \V56(15) ) | ((\[63]  & \V56(4) ) | ((V207 & \V56(7) ) | ~\V174(0) ))),
  \V119(20)  = \[10] ,
  \V151(19)  = \[59] ,
  \[17]  = (\[67]  & \V24(13) ) | ((~\[66]  & \V56(14) ) | ((\[63]  & \V56(3) ) | ((V207 & \V56(6) ) | ~\V174(0) ))),
  \V119(23)  = \[7] ,
  \V151(18)  = \[60] ,
  \[18]  = (\[67]  & \V24(12) ) | ((~\[66]  & \V56(13) ) | ((\[63]  & \V56(2) ) | ((V207 & \V56(5) ) | ~\V174(0) ))),
  \V119(22)  = \[8] ,
  \[19]  = (\[67]  & \V24(11) ) | ((~\[66]  & \V56(12) ) | ((\[63]  & \V56(1) ) | ((V207 & \V56(4) ) | ~\V174(0) ))),
  \V119(25)  = \[5] ,
  \V119(24)  = \[6] ,
  \V119(17)  = \[13] ,
  \[60]  = (\[65]  & \V88(3) ) | ((\[64]  & \V88(18) ) | ((\[63]  & \V88(7) ) | ((V207 & \V88(10) ) | ~\V174(0) ))),
  \V119(16)  = \[14] ,
  \[61]  = (\[65]  & \V88(2) ) | ((\[64]  & \V88(17) ) | ((\[63]  & \V88(6) ) | ((V207 & \V88(9) ) | ~\V174(0) ))),
  \V119(3)  = \[27] ,
  \V119(19)  = \[11] ,
  \[62]  = (\[65]  & \V88(1) ) | ((\[64]  & \V88(16) ) | ((\[63]  & \V88(5) ) | ((V207 & \V88(8) ) | ~\V174(0) ))),
  \V119(2)  = \[28] ,
  \[0]  = (\[67]  & \V56(16) ) | ((~\[66]  & \V56(31) ) | ((\[63]  & \V56(20) ) | ((V207 & \V56(23) ) | ~\V174(0) ))),
  \V119(18)  = \[12] ,
  \V151(11)  = \[35] ,
  \[63]  = ~\V174(2)  & \V174(1) ,
  \V119(5)  = \[25] ,
  \[1]  = (\[67]  & \V56(15) ) | ((~\[66]  & \V56(30) ) | ((\[63]  & \V56(19) ) | ((V207 & \V56(22) ) | ~\V174(0) ))),
  \V151(10)  = \[36] ,
  \[64]  = ~V207 & ~\V174(1) ,
  \V119(4)  = \[26] ,
  \[20]  = (\[67]  & \V24(10) ) | ((~\[66]  & \V56(11) ) | ((V207 & \V56(3) ) | \[71] )),
  \[2]  = (\[67]  & \V56(14) ) | ((~\[66]  & \V56(29) ) | ((\[63]  & \V56(18) ) | ((V207 & \V56(21) ) | ~\V174(0) ))),
  \V151(13)  = \[33] ,
  \[65]  = ~V207 & \V174(2) ,
  \[21]  = (\[67]  & \V24(9) ) | ((~\[66]  & \V56(10) ) | ((V207 & \V56(2) ) | \[72] )),
  \[3]  = (\[67]  & \V56(13) ) | ((~\[66]  & \V56(28) ) | ((\[63]  & \V56(17) ) | ((V207 & \V56(20) ) | ~\V174(0) ))),
  \V151(12)  = \[34] ,
  \[66]  = \V174(2)  | \V174(1) ,
  \[22]  = (\[67]  & \V24(8) ) | ((~\[66]  & \V56(9) ) | ((V207 & \V56(1) ) | \[73] )),
  \[4]  = (\[67]  & \V56(12) ) | ((~\[66]  & \V56(27) ) | ((\[63]  & \V56(16) ) | ((V207 & \V56(19) ) | ~\V174(0) ))),
  \V151(15)  = \[31] ,
  \[67]  = \V174(2)  & \V174(1) ,
  \V119(1)  = \[29] ,
  \[23]  = (\[67]  & \V24(7) ) | ((~\[66]  & \V56(8) ) | ((V207 & \V56(0) ) | \[74] )),
  \[5]  = (\[67]  & \V56(11) ) | ((~\[66]  & \V56(26) ) | ((\[63]  & \V56(15) ) | ((V207 & \V56(18) ) | ~\V174(0) ))),
  \V151(14)  = \[32] ,
  \[68]  = V207 | ~\V174(0) ,
  \V119(0)  = \[30] ,
  \[24]  = (\[63]  & \V88(7) ) | ((\V174(2)  & \V24(6) ) | ((~\V174(1)  & \V56(7) ) | \[68] )),
  \[6]  = (\[67]  & \V56(10) ) | ((~\[66]  & \V56(25) ) | ((\[63]  & \V56(14) ) | ((V207 & \V56(17) ) | ~\V174(0) ))),
  \[69]  = \V9(7)  | \V9(10) ,
  \[25]  = (\[63]  & \V88(6) ) | ((\V174(2)  & \V24(5) ) | ((~\V174(1)  & \V56(6) ) | \[68] )),
  \[7]  = (\[67]  & \V56(9) ) | ((~\[66]  & \V56(24) ) | ((\[63]  & \V56(13) ) | ((V207 & \V56(16) ) | ~\V174(0) ))),
  \V119(11)  = \[19] ,
  \[26]  = (\[63]  & \V88(5) ) | ((\V174(2)  & \V24(4) ) | ((~\V174(1)  & \V56(5) ) | \[68] )),
  \[8]  = (\[67]  & \V56(8) ) | ((~\[66]  & \V56(23) ) | ((\[63]  & \V56(12) ) | ((V207 & \V56(15) ) | ~\V174(0) ))),
  \V119(10)  = \[20] ,
  \[27]  = (\[63]  & \V88(4) ) | ((\V174(2)  & \V24(3) ) | ((~\V174(1)  & \V56(4) ) | \[68] )),
  \[9]  = (\[67]  & \V56(7) ) | ((~\[66]  & \V56(22) ) | ((\[63]  & \V56(11) ) | ((V207 & \V56(14) ) | ~\V174(0) ))),
  \V119(13)  = \[17] ,
  \[28]  = (\[63]  & \V88(3) ) | ((\V174(2)  & \V24(2) ) | ((~\V174(1)  & \V56(3) ) | \[68] )),
  \V119(12)  = \[18] ,
  \V119(7)  = \[23] ,
  \[29]  = (\[63]  & \V88(2) ) | ((\V174(2)  & \V24(1) ) | ((~\V174(1)  & \V56(2) ) | \[68] )),
  \V119(15)  = \[15] ,
  \V119(6)  = \[24] ,
  \V119(14)  = \[16] ,
  \V119(9)  = \[21] ,
  \V119(8)  = \[22] ,
  \[71]  = (\[63]  & \V88(11) ) | ~\V174(0) ,
  V207 = \V174(2)  & ~\V174(1) ,
  \V151(3)  = \[43] ,
  \[72]  = (\[63]  & \V88(10) ) | ~\V174(0) ,
  \V151(2)  = \[44] ,
  \[73]  = (\[63]  & \V88(9) ) | ~\V174(0) ,
  \V151(5)  = \[41] ,
  \[74]  = (\[63]  & \V88(8) ) | ~\V174(0) ,
  \[30]  = (\[63]  & \V88(1) ) | ((\V174(2)  & \V24(0) ) | ((~\V174(1)  & \V56(1) ) | \[68] )),
  \V151(4)  = \[42] ,
  \[31]  = (\[65]  & \V88(0) ) | ((\[64]  & \V88(15) ) | ((\[63]  & \V88(4) ) | ((V207 & \V88(7) ) | ~\V174(0) ))),
  \[32]  = (\[65]  & \V56(31) ) | ((\[64]  & \V88(14) ) | ((\[63]  & \V88(3) ) | ((V207 & \V88(6) ) | ~\V174(0) ))),
  \[33]  = (\[65]  & \V56(30) ) | ((\[64]  & \V88(13) ) | ((\[63]  & \V88(2) ) | ((V207 & \V88(5) ) | ~\V174(0) ))),
  \V151(1)  = \[45] ,
  \[34]  = (\[65]  & \V56(29) ) | ((\[64]  & \V88(12) ) | ((\[63]  & \V88(1) ) | ((V207 & \V88(4) ) | ~\V174(0) ))),
  \V151(0)  = \[46] ,
  \[35]  = (\[65]  & \V56(28) ) | ((\[64]  & \V88(11) ) | ((\[63]  & \V88(0) ) | ((V207 & \V88(3) ) | ~\V174(0) ))),
  \[36]  = (\[65]  & \V56(27) ) | ((\[64]  & \V88(10) ) | ((\[63]  & \V56(31) ) | ((V207 & \V88(2) ) | ~\V174(0) ))),
  \[37]  = (\[65]  & \V56(26) ) | ((\[64]  & \V88(9) ) | ((\[63]  & \V56(30) ) | ((V207 & \V88(1) ) | ~\V174(0) ))),
  \[38]  = (\[65]  & \V56(25) ) | ((\[64]  & \V88(8) ) | ((\[63]  & \V56(29) ) | ((V207 & \V88(0) ) | ~\V174(0) ))),
  \[39]  = (\[65]  & \V56(24) ) | ((\[64]  & \V88(7) ) | ((\[63]  & \V56(28) ) | ((V207 & \V56(31) ) | ~\V174(0) ))),
  \V151(7)  = \[39] ,
  \V151(6)  = \[40] ,
  \V151(9)  = \[37] ,
  \V151(8)  = \[38] ,
  \V151(31)  = \[47] ,
  \V151(30)  = \[48] ,
  \[40]  = (\[65]  & \V56(23) ) | ((\[64]  & \V88(6) ) | ((\[63]  & \V56(27) ) | ((V207 & \V56(30) ) | ~\V174(0) ))),
  \[41]  = (\[65]  & \V56(22) ) | ((\[64]  & \V88(5) ) | ((\[63]  & \V56(26) ) | ((V207 & \V56(29) ) | ~\V174(0) ))),
  \[42]  = (\[65]  & \V56(21) ) | ((\[64]  & \V88(4) ) | ((\[63]  & \V56(25) ) | ((V207 & \V56(28) ) | ~\V174(0) ))),
  \[43]  = (\[65]  & \V56(20) ) | ((\[64]  & \V88(3) ) | ((\[63]  & \V56(24) ) | ((V207 & \V56(27) ) | ~\V174(0) ))),
  \[44]  = (\[65]  & \V56(19) ) | ((\[64]  & \V88(2) ) | ((\[63]  & \V56(23) ) | ((V207 & \V56(26) ) | ~\V174(0) ))),
  \[45]  = (\[65]  & \V56(18) ) | ((\[64]  & \V88(1) ) | ((\[63]  & \V56(22) ) | ((V207 & \V56(25) ) | ~\V174(0) ))),
  \[46]  = (\[65]  & \V56(17) ) | ((\[64]  & \V88(0) ) | ((\[63]  & \V56(21) ) | ((V207 & \V56(24) ) | ~\V174(0) ))),
  \V119(30)  = \[0] ,
  \[47]  = (\[65]  & \V88(16) ) | ((\[64]  & \V88(31) ) | ((\[63]  & \V88(20) ) | ((V207 & \V88(23) ) | ~\V174(0) ))),
  \[48]  = (\[65]  & \V88(15) ) | ((\[64]  & \V88(30) ) | ((\[63]  & \V88(19) ) | ((V207 & \V88(22) ) | ~\V174(0) ))),
  \V151(27)  = \[51] ,
  \[49]  = (\[65]  & \V88(14) ) | ((\[64]  & \V88(29) ) | ((\[63]  & \V88(18) ) | ((V207 & \V88(21) ) | ~\V174(0) ))),
  \V151(26)  = \[52] ,
  \V174(2)  = (~\V9(6)  & (~\V9(5)  & (~\V9(10)  & ~\V9(2) ))) | ((\[69]  & (~\V9(2)  & ~\V9(1) )) | ((\V9(8)  & (~\V9(10)  & \V9(1) )) | ((\V9(7)  & (~\V9(0)  & ~\V9(10) )) | (~\V9(5)  & (~\V9(0)  & ~\V9(10) ))))),
  \V151(29)  = \[49] ,
  \V151(28)  = \[50] ,
  \V174(1)  = (~\V9(6)  & (~\V9(5)  & (\V9(0)  & (~\V9(10)  & ~\V9(1) )))) | ((\V9(8)  & (~\V9(10)  & (\V9(2)  & ~\V9(1) ))) | ((~\V9(6)  & (~\V9(5)  & (~\V9(2)  & ~\V9(1) ))) | ((~\V9(10)  & (\V9(2)  & (\V9(1)  & ~\V9(3) ))) | (\[69]  & (~\V9(2)  & ~\V9(1) ))))),
  \V119(27)  = \[3] ,
  \[50]  = (\[65]  & \V88(13) ) | ((\[64]  & \V88(28) ) | ((\[63]  & \V88(17) ) | ((V207 & \V88(20) ) | ~\V174(0) ))),
  \V174(0)  = (\V9(2)  & \V9(1) ) | (\[66]  | \V9(10) ),
  \V119(26)  = \[4] ,
  \[51]  = (\[65]  & \V88(12) ) | ((\[64]  & \V88(27) ) | ((\[63]  & \V88(16) ) | ((V207 & \V88(19) ) | ~\V174(0) ))),
  \V119(29)  = \[1] ,
  \[52]  = (\[65]  & \V88(11) ) | ((\[64]  & \V88(26) ) | ((\[63]  & \V88(15) ) | ((V207 & \V88(18) ) | ~\V174(0) ))),
  \V119(28)  = \[2] ,
  \V151(21)  = \[57] ,
  \[53]  = (\[65]  & \V88(10) ) | ((\[64]  & \V88(25) ) | ((\[63]  & \V88(14) ) | ((V207 & \V88(17) ) | ~\V174(0) ))),
  \V151(20)  = \[58] ,
  \[54]  = (\[65]  & \V88(9) ) | ((\[64]  & \V88(24) ) | ((\[63]  & \V88(13) ) | ((V207 & \V88(16) ) | ~\V174(0) ))),
  \[10]  = (\[67]  & \V56(6) ) | ((~\[66]  & \V56(21) ) | ((\[63]  & \V56(10) ) | ((V207 & \V56(13) ) | ~\V174(0) ))),
  \V151(23)  = \[55] ,
  \[55]  = (\[65]  & \V88(8) ) | ((\[64]  & \V88(23) ) | ((\[63]  & \V88(12) ) | ((V207 & \V88(15) ) | ~\V174(0) ))),
  \[11]  = (\[67]  & \V56(5) ) | ((~\[66]  & \V56(20) ) | ((\[63]  & \V56(9) ) | ((V207 & \V56(12) ) | ~\V174(0) ))),
  \V151(22)  = \[56] ,
  \[56]  = (\[65]  & \V88(7) ) | ((\[64]  & \V88(22) ) | ((V207 & \V88(14) ) | \[71] )),
  \[12]  = (\[67]  & \V56(4) ) | ((~\[66]  & \V56(19) ) | ((\[63]  & \V56(8) ) | ((V207 & \V56(11) ) | ~\V174(0) ))),
  \V151(25)  = \[53] ,
  \[57]  = (\[65]  & \V88(6) ) | ((\[64]  & \V88(21) ) | ((V207 & \V88(13) ) | \[72] )),
  \[13]  = (\[67]  & \V56(3) ) | ((~\[66]  & \V56(18) ) | ((\[63]  & \V56(7) ) | ((V207 & \V56(10) ) | ~\V174(0) ))),
  \V151(24)  = \[54] ,
  \[58]  = (\[65]  & \V88(5) ) | ((\[64]  & \V88(20) ) | ((V207 & \V88(12) ) | \[73] )),
  \[14]  = (\[67]  & \V56(2) ) | ((~\[66]  & \V56(17) ) | ((\[63]  & \V56(6) ) | ((V207 & \V56(9) ) | ~\V174(0) ))),
  \V151(17)  = \[61] ;
endmodule

