// IWLS benchmark module "MultiplierA_32" printed on Wed May 29 22:12:35 2002
module MultiplierA_32(\1 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \13 , \14 , \15 , \16 , \17 , \18 , \19 , \20 , \21 , \22 , \23 , \24 , \25 , \26 , \27 , \28 , \29 , \30 , \31 , \32 , \33 , \34 , \68 );
input
  \1 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ,
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ,
  \19 ,
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ,
  \34 ;
output
  \68 ;
reg
  \2 ,
  \36 ,
  \37 ,
  \38 ,
  \39 ,
  \40 ,
  \41 ,
  \42 ,
  \43 ,
  \44 ,
  \45 ,
  \46 ,
  \47 ,
  \48 ,
  \49 ,
  \50 ,
  \51 ,
  \52 ,
  \53 ,
  \54 ,
  \55 ,
  \56 ,
  \57 ,
  \58 ,
  \59 ,
  \60 ,
  \61 ,
  \62 ,
  \63 ,
  \64 ,
  \65 ,
  \66 ;
wire
  \[59] ,
  \[60] ,
  \[61] ,
  \[62] ,
  \[63] ,
  \[64] ,
  \[65] ,
  \[66] ,
  \[67] ,
  \[68] ,
  \[69] ,
  \166 ,
  \167 ,
  \168 ,
  \[70] ,
  \169 ,
  \170 ,
  \171 ,
  \172 ,
  \173 ,
  \174 ,
  \175 ,
  \176 ,
  \177 ,
  \178 ,
  \[71] ,
  \179 ,
  \180 ,
  \181 ,
  \182 ,
  \183 ,
  \184 ,
  \185 ,
  \186 ,
  \187 ,
  \188 ,
  \[72] ,
  \189 ,
  \190 ,
  \191 ,
  \192 ,
  \193 ,
  \194 ,
  \195 ,
  \196 ,
  \197 ,
  \198 ,
  \[73] ,
  \[74] ,
  \[75] ,
  \[76] ,
  \[77] ,
  \[33] ,
  \[78] ,
  \[34] ,
  \[79] ,
  \[35] ,
  \203 ,
  \209 ,
  \[36] ,
  \211 ,
  \213 ,
  \215 ,
  \217 ,
  \219 ,
  \[37] ,
  \221 ,
  \223 ,
  \225 ,
  \227 ,
  \229 ,
  \[38] ,
  \231 ,
  \233 ,
  \235 ,
  \237 ,
  \239 ,
  \[39] ,
  \241 ,
  \243 ,
  \245 ,
  \247 ,
  \249 ,
  \251 ,
  \253 ,
  \255 ,
  \257 ,
  \259 ,
  \261 ,
  \263 ,
  \265 ,
  \268 ,
  \[80] ,
  \[81] ,
  \[82] ,
  \[83] ,
  \[84] ,
  \[40] ,
  \[85] ,
  \[41] ,
  \[86] ,
  \[42] ,
  \[87] ,
  \[43] ,
  \[88] ,
  \[44] ,
  \[89] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \[90] ,
  \[91] ,
  \[92] ,
  \[93] ,
  \[94] ,
  \[50] ,
  \[124] ,
  \[95] ,
  \[51] ,
  \[125] ,
  \[96] ,
  \[52] ,
  \[126] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ;
assign
  \[59]  = \193 ,
  \[60]  = \194 ,
  \[61]  = \195 ,
  \[62]  = \196 ,
  \[63]  = \197 ,
  \[64]  = \198 ,
  \[65]  = (\4  & \1 ) | \[124] ,
  \[66]  = \[125]  | \263 ,
  \[67]  = \[126]  | \265 ,
  \[68]  = \209  | \38 ,
  \[69]  = \211  | \39 ,
  \166  = (\[126]  & \265 ) | (\[67]  & \66 ),
  \167  = (~\[96]  & ~\36 ) | (\[96]  & \36 ),
  \168  = (\[124]  & (\37  & \4 )) | ((\[65]  & ~\209 ) | (~\209  & \37 )),
  \[70]  = \213  | \40 ,
  \169  = (~\211  & (\5  & \1 )) | ((\209  & (\38  & \5 )) | (\[68]  & ~\211 )),
  \170  = (~\213  & (\6  & \1 )) | ((\211  & (\39  & \6 )) | (\[69]  & ~\213 )),
  \171  = (~\215  & (\7  & \1 )) | ((\213  & (\40  & \7 )) | (\[70]  & ~\215 )),
  \172  = (~\217  & (\8  & \1 )) | ((\215  & (\41  & \8 )) | (\[71]  & ~\217 )),
  \173  = (~\219  & (\9  & \1 )) | ((\217  & (\42  & \9 )) | (\[72]  & ~\219 )),
  \174  = (~\221  & (\10  & \1 )) | ((\219  & (\43  & \10 )) | (\[73]  & ~\221 )),
  \175  = (~\223  & (\11  & \1 )) | ((\221  & (\44  & \11 )) | (\[74]  & ~\223 )),
  \176  = (~\225  & (\12  & \1 )) | ((\223  & (\45  & \12 )) | (\[75]  & ~\225 )),
  \177  = (~\227  & (\13  & \1 )) | ((\225  & (\46  & \13 )) | (\[76]  & ~\227 )),
  \178  = (~\229  & (\14  & \1 )) | ((\227  & (\47  & \14 )) | (\[77]  & ~\229 )),
  \[71]  = \215  | \41 ,
  \179  = (~\231  & (\15  & \1 )) | ((\229  & (\48  & \15 )) | (\[78]  & ~\231 )),
  \180  = (~\233  & (\16  & \1 )) | ((\231  & (\49  & \16 )) | (\[79]  & ~\233 )),
  \181  = (~\235  & (\17  & \1 )) | ((\233  & (\50  & \17 )) | (\[80]  & ~\235 )),
  \182  = (~\237  & (\18  & \1 )) | ((\235  & (\51  & \18 )) | (\[81]  & ~\237 )),
  \183  = (~\239  & (\19  & \1 )) | ((\237  & (\52  & \19 )) | (\[82]  & ~\239 )),
  \184  = (~\241  & (\20  & \1 )) | ((\239  & (\53  & \20 )) | (\[83]  & ~\241 )),
  \185  = (~\243  & (\21  & \1 )) | ((\241  & (\54  & \21 )) | (\[84]  & ~\243 )),
  \186  = (~\245  & (\22  & \1 )) | ((\243  & (\55  & \22 )) | (\[85]  & ~\245 )),
  \187  = (~\247  & (\23  & \1 )) | ((\245  & (\56  & \23 )) | (\[86]  & ~\247 )),
  \188  = (~\249  & (\24  & \1 )) | ((\247  & (\57  & \24 )) | (\[87]  & ~\249 )),
  \[72]  = \217  | \42 ,
  \189  = (~\251  & (\25  & \1 )) | ((\249  & (\58  & \25 )) | (\[88]  & ~\251 )),
  \190  = (~\253  & (\26  & \1 )) | ((\251  & (\59  & \26 )) | (\[89]  & ~\253 )),
  \191  = (~\255  & (\27  & \1 )) | ((\253  & (\60  & \27 )) | (\[90]  & ~\255 )),
  \192  = (~\257  & (\28  & \1 )) | ((\255  & (\61  & \28 )) | (\[91]  & ~\257 )),
  \193  = (~\259  & (\29  & \1 )) | ((\257  & (\62  & \29 )) | (\[92]  & ~\259 )),
  \194  = (~\261  & (\30  & \1 )) | ((\259  & (\63  & \30 )) | (\[93]  & ~\261 )),
  \195  = (~\263  & (\31  & \1 )) | ((\261  & (\64  & \31 )) | (\[94]  & ~\263 )),
  \196  = (\[125]  & (\263  & \65 )) | ((\[66]  & ~\265 ) | (~\265  & \65 )),
  \197  = (\[126]  & (\265  & \66 )) | ((\[67]  & ~\166 ) | (~\166  & \66 )),
  \198  = (~\268  & \2 ) | (\268  & ~\2 ),
  \[73]  = \219  | \43 ,
  \[74]  = \221  | \44 ,
  \[75]  = \223  | \45 ,
  \[76]  = \225  | \46 ,
  \[77]  = \227  | \47 ,
  \[33]  = \203 ,
  \[78]  = \229  | \48 ,
  \[34]  = \168 ,
  \[79]  = \231  | \49 ,
  \[35]  = \169 ,
  \203  = (~\[95]  & ~\268 ) | (\268  & \2 ),
  \209  = (\[124]  & \4 ) | (\[65]  & \37 ),
  \[36]  = \170 ,
  \211  = (\[68]  & (\5  & \1 )) | (\209  & \38 ),
  \213  = (\[69]  & (\6  & \1 )) | (\211  & \39 ),
  \215  = (\[70]  & (\7  & \1 )) | (\213  & \40 ),
  \217  = (\[71]  & (\8  & \1 )) | (\215  & \41 ),
  \219  = (\[72]  & (\9  & \1 )) | (\217  & \42 ),
  \[37]  = \171 ,
  \221  = (\[73]  & (\10  & \1 )) | (\219  & \43 ),
  \223  = (\[74]  & (\11  & \1 )) | (\221  & \44 ),
  \225  = (\[75]  & (\12  & \1 )) | (\223  & \45 ),
  \227  = (\[76]  & (\13  & \1 )) | (\225  & \46 ),
  \229  = (\[77]  & (\14  & \1 )) | (\227  & \47 ),
  \[38]  = \172 ,
  \231  = (\[78]  & (\15  & \1 )) | (\229  & \48 ),
  \233  = (\[79]  & (\16  & \1 )) | (\231  & \49 ),
  \235  = (\[80]  & (\17  & \1 )) | (\233  & \50 ),
  \237  = (\[81]  & (\18  & \1 )) | (\235  & \51 ),
  \239  = (\[82]  & (\19  & \1 )) | (\237  & \52 ),
  \[39]  = \173 ,
  \241  = (\[83]  & (\20  & \1 )) | (\239  & \53 ),
  \243  = (\[84]  & (\21  & \1 )) | (\241  & \54 ),
  \245  = (\[85]  & (\22  & \1 )) | (\243  & \55 ),
  \247  = (\[86]  & (\23  & \1 )) | (\245  & \56 ),
  \249  = (\[87]  & (\24  & \1 )) | (\247  & \57 ),
  \251  = (\[88]  & (\25  & \1 )) | (\249  & \58 ),
  \253  = (\[89]  & (\26  & \1 )) | (\251  & \59 ),
  \255  = (\[90]  & (\27  & \1 )) | (\253  & \60 ),
  \257  = (\[91]  & (\28  & \1 )) | (\255  & \61 ),
  \259  = (\[92]  & (\29  & \1 )) | (\257  & \62 ),
  \261  = (\[93]  & (\30  & \1 )) | (\259  & \63 ),
  \263  = (\[94]  & (\31  & \1 )) | (\261  & \64 ),
  \265  = (\[125]  & \263 ) | (\[66]  & \65 ),
  \268  = (~\[95]  & ~\166 ) | (\[95]  & \166 ),
  \[80]  = \233  | \50 ,
  \[81]  = \235  | \51 ,
  \[82]  = \237  | \52 ,
  \[83]  = \239  | \53 ,
  \[84]  = \241  | \54 ,
  \[40]  = \174 ,
  \[85]  = \243  | \55 ,
  \[41]  = \175 ,
  \[86]  = \245  | \56 ,
  \[42]  = \176 ,
  \[87]  = \247  | \57 ,
  \[43]  = \177 ,
  \[88]  = \249  | \58 ,
  \[44]  = \178 ,
  \[89]  = \251  | \59 ,
  \[45]  = \179 ,
  \[46]  = \180 ,
  \[47]  = \181 ,
  \[48]  = \182 ,
  \[49]  = \183 ,
  \[90]  = \253  | \60 ,
  \[91]  = \255  | \61 ,
  \[92]  = \257  | \62 ,
  \68  = \167 ,
  \[93]  = \259  | \63 ,
  \[94]  = \261  | \64 ,
  \[50]  = \184 ,
  \[124]  = ~\167  & \36 ,
  \[95]  = ~\34  | ~\1 ,
  \[51]  = \185 ,
  \[125]  = \32  & \1 ,
  \[96]  = ~\3  | ~\1 ,
  \[52]  = \186 ,
  \[126]  = \33  & \1 ,
  \[53]  = \187 ,
  \[54]  = \188 ,
  \[55]  = \189 ,
  \[56]  = \190 ,
  \[57]  = \191 ,
  \[58]  = \192 ;
always begin
  \2  = \[33] ;
  \36  = \[34] ;
  \37  = \[35] ;
  \38  = \[36] ;
  \39  = \[37] ;
  \40  = \[38] ;
  \41  = \[39] ;
  \42  = \[40] ;
  \43  = \[41] ;
  \44  = \[42] ;
  \45  = \[43] ;
  \46  = \[44] ;
  \47  = \[45] ;
  \48  = \[46] ;
  \49  = \[47] ;
  \50  = \[48] ;
  \51  = \[49] ;
  \52  = \[50] ;
  \53  = \[51] ;
  \54  = \[52] ;
  \55  = \[53] ;
  \56  = \[54] ;
  \57  = \[55] ;
  \58  = \[56] ;
  \59  = \[57] ;
  \60  = \[58] ;
  \61  = \[59] ;
  \62  = \[60] ;
  \63  = \[61] ;
  \64  = \[62] ;
  \65  = \[63] ;
  \66  = \[64] ;
end
initial begin
  \2  = 0;
  \36  = 0;
  \37  = 0;
  \38  = 0;
  \39  = 0;
  \40  = 0;
  \41  = 0;
  \42  = 0;
  \43  = 0;
  \44  = 0;
  \45  = 0;
  \46  = 0;
  \47  = 0;
  \48  = 0;
  \49  = 0;
  \50  = 0;
  \51  = 0;
  \52  = 0;
  \53  = 0;
  \54  = 0;
  \55  = 0;
  \56  = 0;
  \57  = 0;
  \58  = 0;
  \59  = 0;
  \60  = 0;
  \61  = 0;
  \62  = 0;
  \63  = 0;
  \64  = 0;
  \65  = 0;
  \66  = 0;
end
endmodule

