module soft_module(clk, d, ena, adata, clrn, q);
  input clk;
  input d;
  input ena;
  input clrn;
  output adata;
  output q;
endmodule
