// IWLS benchmark module "Min_Max9_4" printed on Wed May 29 22:12:22 2002
module Min_Max9_4(\1 , \2 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \40 , \41 , \42 , \43 , \44 , \45 , \46 , \47 , \48 );
input
  \1 ,
  \2 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ;
output
  \40 ,
  \41 ,
  \42 ,
  \43 ,
  \44 ,
  \45 ,
  \46 ,
  \47 ,
  \48 ;
reg
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ,
  \19 ,
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ,
  \34 ,
  \35 ,
  \36 ,
  \37 ,
  \38 ,
  \39 ;
wire
  \49 ,
  \50 ,
  \51 ,
  \52 ,
  \53 ,
  \54 ,
  \55 ,
  \56 ,
  \57 ,
  \58 ,
  \59 ,
  \60 ,
  \61 ,
  \62 ,
  \63 ,
  \64 ,
  \65 ,
  \66 ,
  \67 ,
  \68 ,
  \69 ,
  \70 ,
  \71 ,
  \72 ,
  \73 ,
  \74 ,
  \75 ,
  \76 ,
  \77 ,
  \78 ,
  \79 ,
  \80 ,
  \81 ,
  \82 ,
  \83 ,
  \84 ,
  \85 ,
  \86 ,
  \87 ,
  \88 ,
  \89 ,
  \90 ,
  \91 ,
  \92 ,
  \93 ,
  \94 ,
  \95 ,
  \96 ,
  \97 ,
  \98 ,
  \99 ,
  \100 ,
  \101 ,
  \102 ,
  \103 ,
  \104 ,
  \105 ,
  \106 ,
  \107 ,
  \108 ,
  \109 ,
  \110 ,
  \111 ,
  \112 ,
  \113 ,
  \114 ,
  \115 ,
  \116 ,
  \117 ,
  \118 ,
  \119 ,
  \120 ,
  \121 ,
  \122 ,
  \123 ,
  \124 ,
  \125 ,
  \126 ,
  \127 ,
  \128 ,
  \129 ,
  \130 ,
  \131 ,
  \132 ,
  \133 ,
  \134 ,
  \135 ,
  \136 ,
  \137 ,
  \138 ,
  \139 ,
  \140 ,
  \141 ,
  \142 ,
  \143 ,
  \144 ,
  \145 ,
  \146 ,
  \147 ,
  \148 ,
  \149 ,
  \150 ,
  \151 ,
  \152 ,
  \153 ,
  \154 ,
  \155 ,
  \156 ,
  \157 ,
  \158 ,
  \159 ,
  \160 ,
  \161 ,
  \162 ,
  \163 ,
  \164 ,
  \165 ,
  \166 ,
  \167 ,
  \168 ,
  \169 ,
  \170 ,
  \171 ,
  \172 ,
  \173 ,
  \174 ,
  \175 ,
  \176 ,
  \177 ,
  \178 ,
  \179 ,
  \180 ,
  \181 ,
  \182 ,
  \183 ,
  \184 ,
  \185 ,
  \186 ,
  \187 ,
  \188 ,
  \189 ,
  \190 ,
  \191 ,
  \192 ,
  \193 ,
  \194 ,
  \195 ,
  \196 ,
  \197 ,
  \198 ,
  \199 ,
  \200 ,
  \201 ,
  \202 ,
  \203 ,
  \204 ,
  \205 ,
  \206 ,
  \207 ,
  \208 ,
  \209 ,
  \210 ,
  \211 ,
  \212 ,
  \213 ,
  \214 ,
  \215 ,
  \216 ,
  \217 ,
  \218 ,
  \219 ,
  \220 ,
  \221 ,
  \222 ,
  \223 ,
  \224 ,
  \225 ,
  \226 ,
  \227 ,
  \228 ,
  \229 ,
  \230 ,
  \231 ,
  \232 ,
  \233 ,
  \234 ,
  \235 ,
  \236 ,
  \237 ,
  \238 ,
  \239 ,
  \240 ,
  \241 ,
  \242 ,
  \243 ,
  \244 ,
  \245 ,
  \246 ,
  \247 ,
  \248 ,
  \249 ,
  \250 ,
  \251 ,
  \252 ,
  \253 ,
  \254 ,
  \255 ,
  \256 ,
  \257 ,
  \258 ,
  \259 ,
  \260 ,
  \261 ,
  \262 ,
  \263 ,
  \264 ,
  \265 ,
  \266 ,
  \267 ,
  \268 ,
  \269 ,
  \270 ,
  \271 ,
  \272 ,
  \273 ,
  \274 ,
  \275 ,
  \276 ,
  \277 ,
  \278 ,
  \279 ,
  \280 ,
  \281 ,
  \282 ,
  \283 ,
  \284 ,
  \285 ,
  \286 ,
  \287 ,
  \288 ,
  \289 ,
  \290 ,
  \291 ,
  \292 ,
  \293 ,
  \294 ,
  \295 ,
  \296 ,
  \297 ,
  \298 ,
  \299 ,
  \300 ,
  \301 ,
  \302 ,
  \303 ,
  \304 ,
  \305 ,
  \306 ,
  \307 ,
  \308 ,
  \309 ,
  \310 ,
  \311 ,
  \312 ,
  \313 ,
  \314 ,
  \315 ,
  \316 ,
  \317 ,
  \318 ,
  \319 ,
  \320 ,
  \321 ,
  \322 ,
  \323 ,
  \324 ,
  \325 ,
  \326 ,
  \327 ,
  \328 ,
  \329 ,
  \330 ,
  \331 ,
  \332 ,
  \333 ,
  \334 ,
  \335 ,
  \336 ,
  \337 ,
  \338 ,
  \339 ,
  \340 ,
  \341 ,
  \342 ,
  \343 ,
  \344 ,
  \345 ,
  \346 ,
  \347 ,
  \348 ,
  \349 ,
  \350 ,
  \351 ,
  \352 ,
  \353 ,
  \354 ,
  \355 ,
  \356 ,
  \357 ,
  \358 ,
  \359 ,
  \360 ,
  \361 ,
  \362 ,
  \363 ,
  \364 ,
  \365 ,
  \366 ,
  \367 ,
  \368 ,
  \369 ,
  \370 ,
  \371 ,
  \372 ,
  \373 ,
  \374 ,
  \375 ,
  \376 ,
  \377 ,
  \378 ,
  \379 ,
  \380 ,
  \381 ,
  \382 ,
  \383 ,
  \384 ,
  \385 ,
  \386 ,
  \387 ,
  \388 ,
  \389 ,
  \390 ,
  \391 ,
  \392 ,
  \393 ,
  \394 ,
  \395 ,
  \396 ,
  \397 ,
  \398 ,
  \399 ,
  \400 ,
  \401 ,
  \402 ,
  \403 ,
  \404 ,
  \405 ,
  \406 ,
  \407 ,
  \408 ,
  \409 ,
  \410 ,
  \411 ,
  \412 ,
  \413 ,
  \414 ,
  \415 ,
  \416 ,
  \417 ,
  \418 ,
  \419 ,
  \420 ,
  \421 ,
  \422 ,
  \423 ,
  \424 ,
  \425 ,
  \426 ,
  \427 ,
  \428 ,
  \429 ,
  \430 ,
  \431 ,
  \432 ,
  \433 ,
  \434 ,
  \435 ,
  \436 ,
  \437 ,
  \438 ,
  \439 ,
  \440 ,
  \441 ,
  \442 ,
  \443 ,
  \444 ,
  \445 ,
  \446 ,
  \447 ,
  \448 ,
  \449 ,
  \450 ,
  \451 ,
  \452 ,
  \453 ,
  \454 ,
  \455 ,
  \456 ,
  \457 ,
  \458 ,
  \459 ,
  \460 ,
  \461 ,
  \462 ,
  \463 ,
  \464 ,
  \465 ,
  \466 ,
  \467 ,
  \468 ,
  \469 ,
  \470 ,
  \471 ,
  \472 ,
  \473 ,
  \474 ,
  \475 ,
  \476 ,
  \477 ,
  \478 ,
  \479 ,
  \480 ,
  \481 ,
  \482 ,
  \483 ,
  \484 ,
  \485 ,
  \486 ,
  \487 ,
  \488 ,
  \489 ,
  \490 ,
  \491 ,
  \492 ,
  \493 ,
  \494 ,
  \495 ,
  \496 ,
  \497 ,
  \498 ,
  \499 ,
  \500 ,
  \501 ,
  \502 ,
  \503 ,
  \504 ,
  \505 ,
  \506 ,
  \507 ,
  \508 ,
  \509 ,
  \[27] ,
  \510 ,
  \511 ,
  \512 ,
  \513 ,
  \514 ,
  \515 ,
  \516 ,
  \517 ,
  \518 ,
  \519 ,
  \[28] ,
  \520 ,
  \521 ,
  \522 ,
  \523 ,
  \524 ,
  \525 ,
  \526 ,
  \527 ,
  \528 ,
  \529 ,
  \[29] ,
  \530 ,
  \531 ,
  \532 ,
  \533 ,
  \534 ,
  \535 ,
  \536 ,
  \537 ,
  \538 ,
  \539 ,
  \540 ,
  \541 ,
  \542 ,
  \543 ,
  \544 ,
  \545 ,
  \546 ,
  \547 ,
  \548 ,
  \549 ,
  \550 ,
  \551 ,
  \552 ,
  \553 ,
  \554 ,
  \555 ,
  \556 ,
  \557 ,
  \558 ,
  \559 ,
  \560 ,
  \561 ,
  \562 ,
  \563 ,
  \564 ,
  \565 ,
  \566 ,
  \567 ,
  \568 ,
  \569 ,
  \570 ,
  \571 ,
  \572 ,
  \573 ,
  \574 ,
  \575 ,
  \576 ,
  \577 ,
  \578 ,
  \579 ,
  \580 ,
  \581 ,
  \582 ,
  \583 ,
  \584 ,
  \585 ,
  \586 ,
  \587 ,
  \588 ,
  \589 ,
  \590 ,
  \591 ,
  \592 ,
  \593 ,
  \594 ,
  \595 ,
  \596 ,
  \597 ,
  \598 ,
  \599 ,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \[36] ,
  \600 ,
  \601 ,
  \602 ,
  \603 ,
  \604 ,
  \605 ,
  \606 ,
  \607 ,
  \608 ,
  \609 ,
  \[37] ,
  \610 ,
  \611 ,
  \612 ,
  \613 ,
  \614 ,
  \615 ,
  \616 ,
  \617 ,
  \618 ,
  \619 ,
  \[38] ,
  \620 ,
  \621 ,
  \622 ,
  \623 ,
  \624 ,
  \625 ,
  \626 ,
  \627 ,
  \628 ,
  \629 ,
  \[39] ,
  \630 ,
  \631 ,
  \632 ,
  \633 ,
  \634 ,
  \635 ,
  \636 ,
  \637 ,
  \638 ,
  \639 ,
  \640 ,
  \641 ,
  \642 ,
  \643 ,
  \644 ,
  \645 ,
  \646 ,
  \647 ,
  \648 ,
  \649 ,
  \650 ,
  \651 ,
  \652 ,
  \653 ,
  \654 ,
  \655 ,
  \656 ,
  \657 ,
  \658 ,
  \659 ,
  \660 ,
  \661 ,
  \662 ,
  \663 ,
  \664 ,
  \665 ,
  \666 ,
  \667 ,
  \668 ,
  \669 ,
  \670 ,
  \671 ,
  \672 ,
  \673 ,
  \674 ,
  \675 ,
  \676 ,
  \677 ,
  \678 ,
  \679 ,
  \680 ,
  \681 ,
  \682 ,
  \683 ,
  \684 ,
  \685 ,
  \686 ,
  \687 ,
  \688 ,
  \689 ,
  \690 ,
  \691 ,
  \692 ,
  \693 ,
  \694 ,
  \695 ,
  \696 ,
  \697 ,
  \698 ,
  \699 ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \700 ,
  \701 ,
  \702 ,
  \703 ,
  \704 ,
  \705 ,
  \706 ,
  \707 ,
  \708 ,
  \709 ,
  \[47] ,
  \710 ,
  \711 ,
  \712 ,
  \713 ,
  \714 ,
  \715 ,
  \716 ,
  \717 ,
  \718 ,
  \719 ,
  \[48] ,
  \720 ,
  \721 ,
  \722 ,
  \723 ,
  \724 ,
  \725 ,
  \726 ,
  \727 ,
  \728 ,
  \729 ,
  \[49] ,
  \730 ,
  \731 ,
  \732 ,
  \733 ,
  \734 ,
  \735 ,
  \736 ,
  \737 ,
  \738 ,
  \739 ,
  \740 ,
  \741 ,
  \742 ,
  \743 ,
  \744 ,
  \745 ,
  \746 ,
  \747 ,
  \748 ,
  \749 ,
  \750 ,
  \751 ,
  \752 ,
  \753 ,
  \754 ,
  \755 ,
  \756 ,
  \757 ,
  \758 ,
  \759 ,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ,
  \[59] ,
  \[60] ,
  \[61] ,
  \[62] ;
assign
  \40  = \[27] ,
  \41  = \[28] ,
  \42  = \[29] ,
  \43  = \[30] ,
  \44  = \[31] ,
  \45  = \[32] ,
  \46  = \[33] ,
  \47  = \[34] ,
  \48  = \[35] ,
  \49  = \427  | \426 ,
  \50  = \432  | \431 ,
  \51  = \437  | \436 ,
  \52  = \442  | \441 ,
  \53  = \447  | \446 ,
  \54  = \452  | \451 ,
  \55  = \457  | \456 ,
  \56  = \462  | \461 ,
  \57  = \467  | \466 ,
  \58  = \475  | \474 ,
  \59  = \483  | \482 ,
  \60  = \491  | \490 ,
  \61  = \499  | \498 ,
  \62  = \507  | \506 ,
  \63  = \515  | \514 ,
  \64  = \523  | \522 ,
  \65  = \531  | \530 ,
  \66  = \539  | \538 ,
  \67  = \547  | \546 ,
  \68  = \555  | \554 ,
  \69  = \563  | \562 ,
  \70  = \571  | \570 ,
  \71  = \579  | \578 ,
  \72  = \587  | \586 ,
  \73  = \595  | \594 ,
  \74  = \603  | \602 ,
  \75  = \611  | \610 ,
  \76  = ~\77 ,
  \77  = \1 ,
  \78  = ~\79 ,
  \79  = ~\2 ,
  \80  = ~\81 ,
  \81  = \3 ,
  \82  = ~\83 ,
  \83  = (~\12  & \39 ) | (\12  & ~\39 ),
  \84  = ~\85 ,
  \85  = (~\11  & \38 ) | (\11  & ~\38 ),
  \86  = ~\87 ,
  \87  = (~\10  & \37 ) | (\10  & ~\37 ),
  \88  = ~\89 ,
  \89  = (~\9  & \36 ) | (\9  & ~\36 ),
  \90  = ~\91 ,
  \91  = (~\8  & \35 ) | (\8  & ~\35 ),
  \92  = ~\93 ,
  \93  = (~\7  & \34 ) | (\7  & ~\34 ),
  \94  = ~\95 ,
  \95  = (~\6  & \33 ) | (\6  & ~\33 ),
  \96  = ~\97 ,
  \97  = (~\5  & \32 ) | (\5  & ~\32 ),
  \98  = ~\99 ,
  \99  = (~\4  & \31 ) | (\4  & ~\31 ),
  \100  = ~\101 ,
  \101  = \322 ,
  \102  = ~\103 ,
  \103  = (~\12  & \30 ) | (\12  & ~\30 ),
  \104  = ~\105 ,
  \105  = (~\11  & \29 ) | (\11  & ~\29 ),
  \106  = ~\107 ,
  \107  = (~\10  & \28 ) | (\10  & ~\28 ),
  \108  = ~\109 ,
  \109  = (~\9  & \27 ) | (\9  & ~\27 ),
  \110  = ~\111 ,
  \111  = (~\8  & \26 ) | (\8  & ~\26 ),
  \112  = ~\113 ,
  \113  = (~\7  & \25 ) | (\7  & ~\25 ),
  \114  = ~\115 ,
  \115  = (~\6  & \24 ) | (\6  & ~\24 ),
  \116  = ~\117 ,
  \117  = (~\5  & \23 ) | (\5  & ~\23 ),
  \118  = ~\119 ,
  \119  = (~\4  & \22 ) | (\4  & ~\22 ),
  \120  = ~\121 ,
  \121  = ~\323 ,
  \122  = 0,
  \123  = 0,
  \124  = 0,
  \125  = 0,
  \126  = 0,
  \127  = 0,
  \128  = 0,
  \129  = 0,
  \130  = 0,
  \131  = 0,
  \132  = 0,
  \133  = 0,
  \134  = 0,
  \135  = 0,
  \136  = 0,
  \137  = 0,
  \138  = 0,
  \139  = 0,
  \140  = \4 ,
  \141  = \5 ,
  \142  = \6 ,
  \143  = \7 ,
  \144  = \8 ,
  \145  = \9 ,
  \146  = \10 ,
  \147  = \11 ,
  \148  = \12 ,
  \149  = \13 ,
  \150  = \14 ,
  \151  = \15 ,
  \152  = \16 ,
  \153  = \17 ,
  \154  = \18 ,
  \155  = \19 ,
  \156  = \20 ,
  \157  = \21 ,
  \158  = 0,
  \159  = 0,
  \160  = 0,
  \161  = 0,
  \162  = 0,
  \163  = 0,
  \164  = 0,
  \165  = 0,
  \166  = 0,
  \167  = 0,
  \168  = 0,
  \169  = 0,
  \170  = 0,
  \171  = 0,
  \172  = 0,
  \173  = 0,
  \174  = 0,
  \175  = 0,
  \176  = 1,
  \177  = 1,
  \178  = 1,
  \179  = 1,
  \180  = 1,
  \181  = 1,
  \182  = 1,
  \183  = 1,
  \184  = 1,
  \185  = \4 ,
  \186  = \5 ,
  \187  = \6 ,
  \188  = \7 ,
  \189  = \8 ,
  \190  = \9 ,
  \191  = \10 ,
  \192  = \11 ,
  \193  = \12 ,
  \194  = 1,
  \195  = 1,
  \196  = 1,
  \197  = 1,
  \198  = 1,
  \199  = 1,
  \200  = 1,
  \201  = 1,
  \202  = 1,
  \203  = 0,
  \204  = 0,
  \205  = 0,
  \206  = 0,
  \207  = 0,
  \208  = 0,
  \209  = 0,
  \210  = 0,
  \211  = 0,
  \212  = \13 ,
  \213  = \14 ,
  \214  = \15 ,
  \215  = \16 ,
  \216  = \17 ,
  \217  = \18 ,
  \218  = \19 ,
  \219  = \20 ,
  \220  = \21 ,
  \221  = \12 ,
  \222  = 1,
  \223  = 1,
  \224  = 1,
  \225  = 1,
  \226  = 1,
  \227  = 1,
  \228  = 1,
  \229  = 1,
  \230  = 1,
  \231  = \11 ,
  \232  = \10 ,
  \233  = \9 ,
  \234  = \8 ,
  \235  = \7 ,
  \236  = \6 ,
  \237  = \5 ,
  \238  = 0,
  \239  = \4 ,
  \240  = \31 ,
  \241  = \32 ,
  \242  = \33 ,
  \243  = \34 ,
  \244  = \35 ,
  \245  = \36 ,
  \246  = \37 ,
  \247  = \38 ,
  \248  = \39 ,
  \249  = \4 ,
  \250  = \5 ,
  \251  = \6 ,
  \252  = \7 ,
  \253  = \8 ,
  \254  = \9 ,
  \255  = \10 ,
  \256  = \11 ,
  \257  = \12 ,
  \258  = \12 ,
  \259  = \11 ,
  \260  = \10 ,
  \261  = \9 ,
  \262  = \8 ,
  \263  = \7 ,
  \264  = \6 ,
  \265  = \5 ,
  \266  = 0,
  \267  = \4 ,
  \268  = \22 ,
  \269  = \23 ,
  \270  = \24 ,
  \271  = \25 ,
  \272  = \26 ,
  \273  = \27 ,
  \274  = \28 ,
  \275  = \29 ,
  \276  = \30 ,
  \277  = \4 ,
  \278  = \5 ,
  \279  = \6 ,
  \280  = \7 ,
  \281  = \8 ,
  \282  = \9 ,
  \283  = \10 ,
  \284  = \11 ,
  \285  = \12 ,
  \286  = (\350  & \349 ) | ((\350  & \348 ) | (\349  & \348 )),
  \287  = (~\329  & (~\328  & \327 )) | ((~\329  & (\328  & ~\327 )) | ((\329  & (~\328  & ~\327 )) | (\329  & (\328  & \327 )))),
  \288  = (~\332  & (~\331  & \330 )) | ((~\332  & (\331  & ~\330 )) | ((\332  & (~\331  & ~\330 )) | (\332  & (\331  & \330 )))),
  \289  = (~\335  & (~\334  & \333 )) | ((~\335  & (\334  & ~\333 )) | ((\335  & (~\334  & ~\333 )) | (\335  & (\334  & \333 )))),
  \290  = (~\338  & (~\337  & \336 )) | ((~\338  & (\337  & ~\336 )) | ((\338  & (~\337  & ~\336 )) | (\338  & (\337  & \336 )))),
  \291  = (~\341  & (~\340  & \339 )) | ((~\341  & (\340  & ~\339 )) | ((\341  & (~\340  & ~\339 )) | (\341  & (\340  & \339 )))),
  \292  = (~\344  & (~\343  & \342 )) | ((~\344  & (\343  & ~\342 )) | ((\344  & (~\343  & ~\342 )) | (\344  & (\343  & \342 )))),
  \293  = (~\347  & (~\346  & \345 )) | ((~\347  & (\346  & ~\345 )) | ((\347  & (~\346  & ~\345 )) | (\347  & (\346  & \345 )))),
  \294  = (~\350  & (~\349  & \348 )) | ((~\350  & (\349  & ~\348 )) | ((\350  & (~\349  & ~\348 )) | (\350  & (\349  & \348 )))),
  \295  = \286 ,
  \296  = \287 ,
  \297  = \288 ,
  \298  = \289 ,
  \299  = \290 ,
  \300  = \291 ,
  \301  = \292 ,
  \302  = \293 ,
  \303  = \294 ,
  \304  = \325 ,
  \305  = \328 ,
  \306  = \331 ,
  \307  = \334 ,
  \308  = \337 ,
  \309  = \340 ,
  \310  = \343 ,
  \311  = \346 ,
  \312  = \349 ,
  \313  = \326 ,
  \314  = \329 ,
  \315  = \332 ,
  \316  = \335 ,
  \317  = \338 ,
  \318  = \341 ,
  \319  = \344 ,
  \320  = \347 ,
  \321  = \350 ,
  \322  = \759  & \757 ,
  \323  = \730  & \728 ,
  \324  = 0,
  \325  = \701  & \699 ,
  \326  = \696  & \694 ,
  \327  = (\326  & \325 ) | ((\326  & \324 ) | (\325  & \324 )),
  \328  = \691  & \689 ,
  \329  = \686  & \684 ,
  \330  = (\329  & \328 ) | ((\329  & \327 ) | (\328  & \327 )),
  \331  = \681  & \679 ,
  \332  = \676  & \674 ,
  \333  = (\332  & \331 ) | ((\332  & \330 ) | (\331  & \330 )),
  \334  = \671  & \669 ,
  \335  = \666  & \664 ,
  \336  = (\335  & \334 ) | ((\335  & \333 ) | (\334  & \333 )),
  \337  = \661  & \659 ,
  \338  = \656  & \654 ,
  \339  = (\338  & \337 ) | ((\338  & \336 ) | (\337  & \336 )),
  \340  = \651  & \649 ,
  \341  = \646  & \644 ,
  \342  = (\341  & \340 ) | ((\341  & \339 ) | (\340  & \339 )),
  \343  = \641  & \639 ,
  \344  = \636  & \634 ,
  \345  = (\344  & \343 ) | ((\344  & \342 ) | (\343  & \342 )),
  \346  = \631  & \629 ,
  \347  = \626  & \624 ,
  \348  = (\347  & \346 ) | ((\347  & \345 ) | (\346  & \345 )),
  \349  = \621  & \619 ,
  \350  = \616  & \614 ,
  \351  = \296  & \80 ,
  \352  = \185  & \81 ,
  \353  = \352  | \351 ,
  \354  = \353  & \78 ,
  \355  = \149  & \79 ,
  \356  = \355  | \354 ,
  \357  = \356  & \76 ,
  \358  = \122  & \77 ,
  \359  = \297  & \80 ,
  \360  = \186  & \81 ,
  \361  = \360  | \359 ,
  \362  = \361  & \78 ,
  \363  = \150  & \79 ,
  \364  = \363  | \362 ,
  \365  = \364  & \76 ,
  \366  = \123  & \77 ,
  \367  = \298  & \80 ,
  \368  = \187  & \81 ,
  \369  = \368  | \367 ,
  \370  = \369  & \78 ,
  \371  = \151  & \79 ,
  \372  = \371  | \370 ,
  \373  = \372  & \76 ,
  \374  = \124  & \77 ,
  \375  = \299  & \80 ,
  \376  = \188  & \81 ,
  \377  = \376  | \375 ,
  \378  = \377  & \78 ,
  \379  = \152  & \79 ,
  \380  = \379  | \378 ,
  \381  = \380  & \76 ,
  \382  = \125  & \77 ,
  \383  = \300  & \80 ,
  \384  = \189  & \81 ,
  \385  = \384  | \383 ,
  \386  = \385  & \78 ,
  \387  = \153  & \79 ,
  \388  = \387  | \386 ,
  \389  = \388  & \76 ,
  \390  = \126  & \77 ,
  \391  = \301  & \80 ,
  \392  = \190  & \81 ,
  \393  = \392  | \391 ,
  \394  = \393  & \78 ,
  \395  = \154  & \79 ,
  \396  = \395  | \394 ,
  \397  = \396  & \76 ,
  \398  = \127  & \77 ,
  \399  = \302  & \80 ,
  \400  = \191  & \81 ,
  \401  = \400  | \399 ,
  \402  = \401  & \78 ,
  \403  = \155  & \79 ,
  \404  = \403  | \402 ,
  \405  = \404  & \76 ,
  \406  = \128  & \77 ,
  \407  = \303  & \80 ,
  \408  = \192  & \81 ,
  \409  = \408  | \407 ,
  \410  = \409  & \78 ,
  \411  = \156  & \79 ,
  \412  = \411  | \410 ,
  \413  = \412  & \76 ,
  \414  = \129  & \77 ,
  \415  = \295  & \80 ,
  \416  = \193  & \81 ,
  \417  = \416  | \415 ,
  \418  = \417  & \78 ,
  \419  = \157  & \79 ,
  \420  = \419  | \418 ,
  \421  = \420  & \76 ,
  \422  = \130  & \77 ,
  \423  = \140  & \78 ,
  \424  = \212  & \79 ,
  \425  = \424  | \423 ,
  \426  = \425  & \76 ,
  \427  = \131  & \77 ,
  \428  = \141  & \78 ,
  \429  = \213  & \79 ,
  \430  = \429  | \428 ,
  \431  = \430  & \76 ,
  \432  = \132  & \77 ,
  \433  = \142  & \78 ,
  \434  = \214  & \79 ,
  \435  = \434  | \433 ,
  \436  = \435  & \76 ,
  \437  = \133  & \77 ,
  \438  = \143  & \78 ,
  \439  = \215  & \79 ,
  \440  = \439  | \438 ,
  \441  = \440  & \76 ,
  \442  = \134  & \77 ,
  \443  = \144  & \78 ,
  \444  = \216  & \79 ,
  \445  = \444  | \443 ,
  \446  = \445  & \76 ,
  \447  = \135  & \77 ,
  \448  = \145  & \78 ,
  \449  = \217  & \79 ,
  \450  = \449  | \448 ,
  \451  = \450  & \76 ,
  \452  = \136  & \77 ,
  \453  = \146  & \78 ,
  \454  = \218  & \79 ,
  \455  = \454  | \453 ,
  \456  = \455  & \76 ,
  \457  = \137  & \77 ,
  \458  = \147  & \78 ,
  \459  = \219  & \79 ,
  \460  = \459  | \458 ,
  \461  = \460  & \76 ,
  \462  = \138  & \77 ,
  \463  = \148  & \78 ,
  \464  = \220  & \79 ,
  \465  = \464  | \463 ,
  \466  = \465  & \76 ,
  \467  = \139  & \77 ,
  \468  = \313  & \80 ,
  \469  = \222  & \81 ,
  \470  = \469  | \468 ,
  \471  = \470  & \78 ,
  \472  = \194  & \79 ,
  \473  = \472  | \471 ,
  \474  = \473  & \76 ,
  \475  = \176  & \77 ,
  \476  = \314  & \80 ,
  \477  = \223  & \81 ,
  \478  = \477  | \476 ,
  \479  = \478  & \78 ,
  \480  = \195  & \79 ,
  \481  = \480  | \479 ,
  \482  = \481  & \76 ,
  \483  = \177  & \77 ,
  \484  = \315  & \80 ,
  \485  = \224  & \81 ,
  \486  = \485  | \484 ,
  \487  = \486  & \78 ,
  \488  = \196  & \79 ,
  \489  = \488  | \487 ,
  \490  = \489  & \76 ,
  \491  = \178  & \77 ,
  \492  = \316  & \80 ,
  \493  = \225  & \81 ,
  \494  = \493  | \492 ,
  \495  = \494  & \78 ,
  \496  = \197  & \79 ,
  \497  = \496  | \495 ,
  \498  = \497  & \76 ,
  \499  = \179  & \77 ,
  \500  = \317  & \80 ,
  \501  = \226  & \81 ,
  \502  = \501  | \500 ,
  \503  = \502  & \78 ,
  \504  = \198  & \79 ,
  \505  = \504  | \503 ,
  \506  = \505  & \76 ,
  \507  = \180  & \77 ,
  \508  = \318  & \80 ,
  \509  = \227  & \81 ,
  \[27]  = \358  | \357 ,
  \510  = \509  | \508 ,
  \511  = \510  & \78 ,
  \512  = \199  & \79 ,
  \513  = \512  | \511 ,
  \514  = \513  & \76 ,
  \515  = \181  & \77 ,
  \516  = \319  & \80 ,
  \517  = \228  & \81 ,
  \518  = \517  | \516 ,
  \519  = \518  & \78 ,
  \[28]  = \366  | \365 ,
  \520  = \200  & \79 ,
  \521  = \520  | \519 ,
  \522  = \521  & \76 ,
  \523  = \182  & \77 ,
  \524  = \320  & \80 ,
  \525  = \229  & \81 ,
  \526  = \525  | \524 ,
  \527  = \526  & \78 ,
  \528  = \201  & \79 ,
  \529  = \528  | \527 ,
  \[29]  = \374  | \373 ,
  \530  = \529  & \76 ,
  \531  = \183  & \77 ,
  \532  = \321  & \80 ,
  \533  = \230  & \81 ,
  \534  = \533  | \532 ,
  \535  = \534  & \78 ,
  \536  = \202  & \79 ,
  \537  = \536  | \535 ,
  \538  = \537  & \76 ,
  \539  = \184  & \77 ,
  \540  = \304  & \80 ,
  \541  = \203  & \81 ,
  \542  = \541  | \540 ,
  \543  = \542  & \78 ,
  \544  = \167  & \79 ,
  \545  = \544  | \543 ,
  \546  = \545  & \76 ,
  \547  = \158  & \77 ,
  \548  = \305  & \80 ,
  \549  = \204  & \81 ,
  \550  = \549  | \548 ,
  \551  = \550  & \78 ,
  \552  = \168  & \79 ,
  \553  = \552  | \551 ,
  \554  = \553  & \76 ,
  \555  = \159  & \77 ,
  \556  = \306  & \80 ,
  \557  = \205  & \81 ,
  \558  = \557  | \556 ,
  \559  = \558  & \78 ,
  \560  = \169  & \79 ,
  \561  = \560  | \559 ,
  \562  = \561  & \76 ,
  \563  = \160  & \77 ,
  \564  = \307  & \80 ,
  \565  = \206  & \81 ,
  \566  = \565  | \564 ,
  \567  = \566  & \78 ,
  \568  = \170  & \79 ,
  \569  = \568  | \567 ,
  \570  = \569  & \76 ,
  \571  = \161  & \77 ,
  \572  = \308  & \80 ,
  \573  = \207  & \81 ,
  \574  = \573  | \572 ,
  \575  = \574  & \78 ,
  \576  = \171  & \79 ,
  \577  = \576  | \575 ,
  \578  = \577  & \76 ,
  \579  = \162  & \77 ,
  \580  = \309  & \80 ,
  \581  = \208  & \81 ,
  \582  = \581  | \580 ,
  \583  = \582  & \78 ,
  \584  = \172  & \79 ,
  \585  = \584  | \583 ,
  \586  = \585  & \76 ,
  \587  = \163  & \77 ,
  \588  = \310  & \80 ,
  \589  = \209  & \81 ,
  \590  = \589  | \588 ,
  \591  = \590  & \78 ,
  \592  = \173  & \79 ,
  \593  = \592  | \591 ,
  \594  = \593  & \76 ,
  \595  = \164  & \77 ,
  \596  = \311  & \80 ,
  \597  = \210  & \81 ,
  \598  = \597  | \596 ,
  \599  = \598  & \78 ,
  \[30]  = \382  | \381 ,
  \[31]  = \390  | \389 ,
  \[32]  = \398  | \397 ,
  \[33]  = \406  | \405 ,
  \[34]  = \414  | \413 ,
  \[35]  = \422  | \421 ,
  \[36]  = \49 ,
  \600  = \174  & \79 ,
  \601  = \600  | \599 ,
  \602  = \601  & \76 ,
  \603  = \165  & \77 ,
  \604  = \312  & \80 ,
  \605  = \211  & \81 ,
  \606  = \605  | \604 ,
  \607  = \606  & \78 ,
  \608  = \175  & \79 ,
  \609  = \608  | \607 ,
  \[37]  = \50 ,
  \610  = \609  & \76 ,
  \611  = \166  & \77 ,
  \612  = \276  & \120 ,
  \613  = \285  & \121 ,
  \614  = \613  | \612 ,
  \615  = \80  & \78 ,
  \616  = \615  & \76 ,
  \617  = \248  & \100 ,
  \618  = \257  & \101 ,
  \619  = \618  | \617 ,
  \[38]  = \51 ,
  \620  = \80  & \78 ,
  \621  = \620  & \76 ,
  \622  = \275  & \120 ,
  \623  = \284  & \121 ,
  \624  = \623  | \622 ,
  \625  = \80  & \78 ,
  \626  = \625  & \76 ,
  \627  = \247  & \100 ,
  \628  = \256  & \101 ,
  \629  = \628  | \627 ,
  \[39]  = \52 ,
  \630  = \80  & \78 ,
  \631  = \630  & \76 ,
  \632  = \274  & \120 ,
  \633  = \283  & \121 ,
  \634  = \633  | \632 ,
  \635  = \80  & \78 ,
  \636  = \635  & \76 ,
  \637  = \246  & \100 ,
  \638  = \255  & \101 ,
  \639  = \638  | \637 ,
  \640  = \80  & \78 ,
  \641  = \640  & \76 ,
  \642  = \273  & \120 ,
  \643  = \282  & \121 ,
  \644  = \643  | \642 ,
  \645  = \80  & \78 ,
  \646  = \645  & \76 ,
  \647  = \245  & \100 ,
  \648  = \254  & \101 ,
  \649  = \648  | \647 ,
  \650  = \80  & \78 ,
  \651  = \650  & \76 ,
  \652  = \272  & \120 ,
  \653  = \281  & \121 ,
  \654  = \653  | \652 ,
  \655  = \80  & \78 ,
  \656  = \655  & \76 ,
  \657  = \244  & \100 ,
  \658  = \253  & \101 ,
  \659  = \658  | \657 ,
  \660  = \80  & \78 ,
  \661  = \660  & \76 ,
  \662  = \271  & \120 ,
  \663  = \280  & \121 ,
  \664  = \663  | \662 ,
  \665  = \80  & \78 ,
  \666  = \665  & \76 ,
  \667  = \243  & \100 ,
  \668  = \252  & \101 ,
  \669  = \668  | \667 ,
  \670  = \80  & \78 ,
  \671  = \670  & \76 ,
  \672  = \270  & \120 ,
  \673  = \279  & \121 ,
  \674  = \673  | \672 ,
  \675  = \80  & \78 ,
  \676  = \675  & \76 ,
  \677  = \242  & \100 ,
  \678  = \251  & \101 ,
  \679  = \678  | \677 ,
  \680  = \80  & \78 ,
  \681  = \680  & \76 ,
  \682  = \269  & \120 ,
  \683  = \278  & \121 ,
  \684  = \683  | \682 ,
  \685  = \80  & \78 ,
  \686  = \685  & \76 ,
  \687  = \241  & \100 ,
  \688  = \250  & \101 ,
  \689  = \688  | \687 ,
  \690  = \80  & \78 ,
  \691  = \690  & \76 ,
  \692  = \268  & \120 ,
  \693  = \277  & \121 ,
  \694  = \693  | \692 ,
  \695  = \80  & \78 ,
  \696  = \695  & \76 ,
  \697  = \240  & \100 ,
  \698  = \249  & \101 ,
  \699  = \698  | \697 ,
  \[40]  = \53 ,
  \[41]  = \54 ,
  \[42]  = \55 ,
  \[43]  = \56 ,
  \[44]  = \57 ,
  \[45]  = \58 ,
  \[46]  = \59 ,
  \700  = \80  & \78 ,
  \701  = \700  & \76 ,
  \702  = \266  & \118 ,
  \703  = \267  & \119 ,
  \704  = \703  | \702 ,
  \705  = \704  & \116 ,
  \706  = \265  & \117 ,
  \707  = \706  | \705 ,
  \708  = \707  & \114 ,
  \709  = \264  & \115 ,
  \[47]  = \60 ,
  \710  = \709  | \708 ,
  \711  = \710  & \112 ,
  \712  = \263  & \113 ,
  \713  = \712  | \711 ,
  \714  = \713  & \110 ,
  \715  = \262  & \111 ,
  \716  = \715  | \714 ,
  \717  = \716  & \108 ,
  \718  = \261  & \109 ,
  \719  = \718  | \717 ,
  \[48]  = \61 ,
  \720  = \719  & \106 ,
  \721  = \260  & \107 ,
  \722  = \721  | \720 ,
  \723  = \722  & \104 ,
  \724  = \259  & \105 ,
  \725  = \724  | \723 ,
  \726  = \725  & \102 ,
  \727  = \258  & \103 ,
  \728  = \727  | \726 ,
  \729  = \80  & \78 ,
  \[49]  = \62 ,
  \730  = \729  & \76 ,
  \731  = \238  & \98 ,
  \732  = \239  & \99 ,
  \733  = \732  | \731 ,
  \734  = \733  & \96 ,
  \735  = \237  & \97 ,
  \736  = \735  | \734 ,
  \737  = \736  & \94 ,
  \738  = \236  & \95 ,
  \739  = \738  | \737 ,
  \740  = \739  & \92 ,
  \741  = \235  & \93 ,
  \742  = \741  | \740 ,
  \743  = \742  & \90 ,
  \744  = \234  & \91 ,
  \745  = \744  | \743 ,
  \746  = \745  & \88 ,
  \747  = \233  & \89 ,
  \748  = \747  | \746 ,
  \749  = \748  & \86 ,
  \750  = \232  & \87 ,
  \751  = \750  | \749 ,
  \752  = \751  & \84 ,
  \753  = \231  & \85 ,
  \754  = \753  | \752 ,
  \755  = \754  & \82 ,
  \756  = \221  & \83 ,
  \757  = \756  | \755 ,
  \758  = \80  & \78 ,
  \759  = \758  & \76 ,
  \[50]  = \63 ,
  \[51]  = \64 ,
  \[52]  = \65 ,
  \[53]  = \66 ,
  \[54]  = \67 ,
  \[55]  = \68 ,
  \[56]  = \69 ,
  \[57]  = \70 ,
  \[58]  = \71 ,
  \[59]  = \72 ,
  \[60]  = \73 ,
  \[61]  = \74 ,
  \[62]  = \75 ;
always begin
  \13  = \[36] ;
  \14  = \[37] ;
  \15  = \[38] ;
  \16  = \[39] ;
  \17  = \[40] ;
  \18  = \[41] ;
  \19  = \[42] ;
  \20  = \[43] ;
  \21  = \[44] ;
  \22  = \[45] ;
  \23  = \[46] ;
  \24  = \[47] ;
  \25  = \[48] ;
  \26  = \[49] ;
  \27  = \[50] ;
  \28  = \[51] ;
  \29  = \[52] ;
  \30  = \[53] ;
  \31  = \[54] ;
  \32  = \[55] ;
  \33  = \[56] ;
  \34  = \[57] ;
  \35  = \[58] ;
  \36  = \[59] ;
  \37  = \[60] ;
  \38  = \[61] ;
  \39  = \[62] ;
end
initial begin
  \22  = 1;
  \23  = 1;
  \24  = 1;
  \25  = 1;
  \26  = 1;
  \27  = 1;
  \28  = 1;
  \29  = 1;
  \30  = 1;
  \31  = 0;
  \32  = 0;
  \33  = 0;
  \34  = 0;
  \35  = 0;
  \36  = 0;
  \37  = 0;
  \38  = 0;
  \39  = 0;
end
endmodule

