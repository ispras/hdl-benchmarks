// IWLS benchmark module "DES" printed on Wed May 29 16:32:30 2002
module DES(\data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , \data_in<1> , \data_in<0> , \reset<0> , \encrypt<0> , \load_key<0> , \inreg<55> , \inreg<54> , \inreg<53> , \inreg<52> , \inreg<51> , \inreg<50> , \inreg<49> , \inreg<48> , \inreg<47> , \inreg<46> , \inreg<45> , \inreg<44> , \inreg<43> , \inreg<42> , \inreg<41> , \inreg<40> , \inreg<39> , \inreg<38> , \inreg<37> , \inreg<36> , \inreg<35> , \inreg<34> , \inreg<33> , \inreg<32> , \inreg<31> , \inreg<30> , \inreg<29> , \inreg<28> , \inreg<27> , \inreg<26> , \inreg<25> , \inreg<24> , \inreg<23> , \inreg<22> , \inreg<21> , \inreg<20> , \inreg<19> , \inreg<18> , \inreg<17> , \inreg<16> , \inreg<15> , \inreg<14> , \inreg<13> , \inreg<12> , \inreg<11> , \inreg<10> , \inreg<9> , \inreg<8> , \inreg<7> , \inreg<6> , \inreg<5> , \inreg<4> , \inreg<3> , \inreg<2> , \inreg<1> , \inreg<0> , \outreg<63> , \outreg<62> , \outreg<61> , \outreg<60> , \outreg<59> , \outreg<58> , \outreg<57> , \outreg<56> , \outreg<55> , \outreg<54> , \outreg<53> , \outreg<52> , \outreg<51> , \outreg<50> , \outreg<49> , \outreg<48> , \outreg<47> , \outreg<46> , \outreg<45> , \outreg<44> , \outreg<43> , \outreg<42> , \outreg<41> , \outreg<40> , \outreg<39> , \outreg<38> , \outreg<37> , \outreg<36> , \outreg<35> , \outreg<34> , \outreg<33> , \outreg<32> , \outreg<31> , \outreg<30> , \outreg<29> , \outreg<28> , \outreg<27> , \outreg<26> , \outreg<25> , \outreg<24> , \outreg<23> , \outreg<22> , \outreg<21> , \outreg<20> , \outreg<19> , \outreg<18> , \outreg<17> , \outreg<16> , \outreg<15> , \outreg<14> , \outreg<13> , \outreg<12> , \outreg<11> , \outreg<10> , \outreg<9> , \outreg<8> , \outreg<7> , \outreg<6> , \outreg<5> , \outreg<4> , \outreg<3> , \outreg<2> , \outreg<1> , \outreg<0> , \data<63> , \data<62> , \data<61> , \data<60> , \data<59> , \data<58> , \data<57> , \data<56> , \data<55> , \data<54> , \data<53> , \data<52> , \data<51> , \data<50> , \data<49> , \data<48> , \data<47> , \data<46> , \data<45> , \data<44> , \data<43> , \data<42> , \data<41> , \data<40> , \data<39> , \data<38> , \data<37> , \data<36> , \data<35> , \data<34> , \data<33> , \data<32> , \data<31> , \data<30> , \data<29> , \data<28> , \data<27> , \data<26> , \data<25> , \data<24> , \data<23> , \data<22> , \data<21> , \data<20> , \data<19> , \data<18> , \data<17> , \data<16> , \data<15> , \data<14> , \data<13> , \data<12> , \data<11> , \data<10> , \data<9> , \data<8> , \data<7> , \data<6> , \data<5> , \data<4> , \data<3> , \data<2> , \data<1> , \data<0> , \count<3> , \count<2> , \count<1> , \count<0> , \C<27> , \C<26> , \C<25> , \C<24> , \C<23> , \C<22> , \C<21> , \C<20> , \C<19> , \C<18> , \C<17> , \C<16> , \C<15> , \C<14> , \C<13> , \C<12> , \C<11> , \C<10> , \C<9> , \C<8> , \C<7> , \C<6> , \C<5> , \C<4> , \C<3> , \C<2> , \C<1> , \C<0> , \D<27> , \D<26> , \D<25> , \D<24> , \D<23> , \D<22> , \D<21> , \D<20> , \D<19> , \D<18> , \D<17> , \D<16> , \D<15> , \D<14> , \D<13> , \D<12> , \D<11> , \D<10> , \D<9> , \D<8> , \D<7> , \D<6> , \D<5> , \D<4> , \D<3> , \D<2> , \D<1> , \D<0> , \encrypt_mode<0> , \inreg_new<55> , \inreg_new<54> , \inreg_new<53> , \inreg_new<52> , \inreg_new<51> , \inreg_new<50> , \inreg_new<49> , \inreg_new<48> , \inreg_new<47> , \inreg_new<46> , \inreg_new<45> , \inreg_new<44> , \inreg_new<43> , \inreg_new<42> , \inreg_new<41> , \inreg_new<40> , \inreg_new<39> , \inreg_new<38> , \inreg_new<37> , \inreg_new<36> , \inreg_new<35> , \inreg_new<34> , \inreg_new<33> , \inreg_new<32> , \inreg_new<31> , \inreg_new<30> , \inreg_new<29> , \inreg_new<28> , \inreg_new<27> , \inreg_new<26> , \inreg_new<25> , \inreg_new<24> , \inreg_new<23> , \inreg_new<22> , \inreg_new<21> , \inreg_new<20> , \inreg_new<19> , \inreg_new<18> , \inreg_new<17> , \inreg_new<16> , \inreg_new<15> , \inreg_new<14> , \inreg_new<13> , \inreg_new<12> , \inreg_new<11> , \inreg_new<10> , \inreg_new<9> , \inreg_new<8> , \inreg_new<7> , \inreg_new<6> , \inreg_new<5> , \inreg_new<4> , \inreg_new<3> , \inreg_new<2> , \inreg_new<1> , \inreg_new<0> , \outreg_new<63> , \outreg_new<62> , \outreg_new<61> , \outreg_new<60> , \outreg_new<59> , \outreg_new<58> , \outreg_new<57> , \outreg_new<56> , \outreg_new<55> , \outreg_new<54> , \outreg_new<53> , \outreg_new<52> , \outreg_new<51> , \outreg_new<50> , \outreg_new<49> , \outreg_new<48> , \outreg_new<47> , \outreg_new<46> , \outreg_new<45> , \outreg_new<44> , \outreg_new<43> , \outreg_new<42> , \outreg_new<41> , \outreg_new<40> , \outreg_new<39> , \outreg_new<38> , \outreg_new<37> , \outreg_new<36> , \outreg_new<35> , \outreg_new<34> , \outreg_new<33> , \outreg_new<32> , \outreg_new<31> , \outreg_new<30> , \outreg_new<29> , \outreg_new<28> , \outreg_new<27> , \outreg_new<26> , \outreg_new<25> , \outreg_new<24> , \outreg_new<23> , \outreg_new<22> , \outreg_new<21> , \outreg_new<20> , \outreg_new<19> , \outreg_new<18> , \outreg_new<17> , \outreg_new<16> , \outreg_new<15> , \outreg_new<14> , \outreg_new<13> , \outreg_new<12> , \outreg_new<11> , \outreg_new<10> , \outreg_new<9> , \outreg_new<8> , \outreg_new<7> , \outreg_new<6> , \outreg_new<5> , \outreg_new<4> , \outreg_new<3> , \outreg_new<2> , \outreg_new<1> , \outreg_new<0> , \data_new<63> , \data_new<62> , \data_new<61> , \data_new<60> , \data_new<59> , \data_new<58> , \data_new<57> , \data_new<56> , \data_new<55> , \data_new<54> , \data_new<53> , \data_new<52> , \data_new<51> , \data_new<50> , \data_new<49> , \data_new<48> , \data_new<47> , \data_new<46> , \data_new<45> , \data_new<44> , \data_new<43> , \data_new<42> , \data_new<41> , \data_new<40> , \data_new<39> , \data_new<38> , \data_new<37> , \data_new<36> , \data_new<35> , \data_new<34> , \data_new<33> , \data_new<32> , \data_new<31> , \data_new<30> , \data_new<29> , \data_new<28> , \data_new<27> , \data_new<26> , \data_new<25> , \data_new<24> , \data_new<23> , \data_new<22> , \data_new<21> , \data_new<20> , \data_new<19> , \data_new<18> , \data_new<17> , \data_new<16> , \data_new<15> , \data_new<14> , \data_new<13> , \data_new<12> , \data_new<11> , \data_new<10> , \data_new<9> , \data_new<8> , \data_new<7> , \data_new<6> , \data_new<5> , \data_new<4> , \data_new<3> , \data_new<2> , \data_new<1> , \data_new<0> , \count_new<3> , \count_new<2> , \count_new<1> , \count_new<0> , \C_new<27> , \C_new<26> , \C_new<25> , \C_new<24> , \C_new<23> , \C_new<22> , \C_new<21> , \C_new<20> , \C_new<19> , \C_new<18> , \C_new<17> , \C_new<16> , \C_new<15> , \C_new<14> , \C_new<13> , \C_new<12> , \C_new<11> , \C_new<10> , \C_new<9> , \C_new<8> , \C_new<7> , \C_new<6> , \C_new<5> , \C_new<4> , \C_new<3> , \C_new<2> , \C_new<1> , \C_new<0> , \D_new<27> , \D_new<26> , \D_new<25> , \D_new<24> , \D_new<23> , \D_new<22> , \D_new<21> , \D_new<20> , \D_new<19> , \D_new<18> , \D_new<17> , \D_new<16> , \D_new<15> , \D_new<14> , \D_new<13> , \D_new<12> , \D_new<11> , \D_new<10> , \D_new<9> , \D_new<8> , \D_new<7> , \D_new<6> , \D_new<5> , \D_new<4> , \D_new<3> , \D_new<2> , \D_new<1> , \D_new<0> , \encrypt_mode_new<0> );
input
  \data<63> ,
  \data<61> ,
  \data<62> ,
  \reset<0> ,
  \outreg<58> ,
  \inreg<0> ,
  \outreg<57> ,
  \inreg<1> ,
  \outreg<56> ,
  \inreg<2> ,
  \outreg<55> ,
  \inreg<3> ,
  \inreg<4> ,
  \inreg<5> ,
  \inreg<6> ,
  \outreg<59> ,
  \inreg<7> ,
  \outreg<50> ,
  \inreg<8> ,
  \inreg<9> ,
  \outreg<54> ,
  \outreg<53> ,
  \outreg<52> ,
  \outreg<51> ,
  \load_key<0> ,
  \outreg<60> ,
  \outreg<63> ,
  \outreg<62> ,
  \outreg<61> ,
  \D<0> ,
  \D<1> ,
  \D<2> ,
  \D<3> ,
  \D<4> ,
  \D<5> ,
  \D<6> ,
  \C<10> ,
  \D<7> ,
  \C<11> ,
  \D<8> ,
  \C<12> ,
  \D<9> ,
  \C<13> ,
  \C<14> ,
  \C<15> ,
  \C<16> ,
  \C<17> ,
  \C<18> ,
  \C<19> ,
  \outreg<18> ,
  \outreg<17> ,
  \outreg<16> ,
  \outreg<15> ,
  \C<20> ,
  \outreg<19> ,
  \C<21> ,
  \outreg<10> ,
  \C<22> ,
  \C<23> ,
  \C<24> ,
  \C<25> ,
  \outreg<14> ,
  \C<26> ,
  \outreg<13> ,
  \C<27> ,
  \outreg<12> ,
  \outreg<11> ,
  \outreg<28> ,
  \outreg<27> ,
  \outreg<26> ,
  \outreg<25> ,
  \outreg<29> ,
  \outreg<20> ,
  \data<3> ,
  \data<4> ,
  \data<1> ,
  \outreg<24> ,
  \data<2> ,
  \outreg<23> ,
  \outreg<22> ,
  \data<0> ,
  \outreg<21> ,
  \outreg<38> ,
  \outreg<37> ,
  \outreg<36> ,
  \outreg<35> ,
  \data<9> ,
  \data<7> ,
  \data<8> ,
  \outreg<39> ,
  \data<5> ,
  \outreg<30> ,
  \data<6> ,
  \outreg<34> ,
  \outreg<33> ,
  \outreg<32> ,
  \outreg<31> ,
  \outreg<48> ,
  \outreg<47> ,
  \outreg<46> ,
  \outreg<45> ,
  \outreg<49> ,
  \outreg<40> ,
  \outreg<44> ,
  \outreg<43> ,
  \outreg<42> ,
  \outreg<41> ,
  \D<10> ,
  \D<11> ,
  \D<12> ,
  \D<13> ,
  \D<14> ,
  \D<15> ,
  \D<16> ,
  \D<17> ,
  \D<18> ,
  \D<19> ,
  \D<20> ,
  \D<21> ,
  \data_in<7> ,
  \D<22> ,
  \D<23> ,
  \data_in<5> ,
  \D<24> ,
  \data_in<6> ,
  \D<25> ,
  \D<26> ,
  \D<27> ,
  \data_in<0> ,
  \data_in<3> ,
  \data_in<4> ,
  \data_in<1> ,
  \data_in<2> ,
  \data<37> ,
  \data<38> ,
  \data<35> ,
  \data<36> ,
  \data<39> ,
  \data<30> ,
  \data<33> ,
  \data<34> ,
  \data<31> ,
  \data<32> ,
  \data<47> ,
  \data<48> ,
  \data<45> ,
  \data<46> ,
  \data<49> ,
  \data<40> ,
  \data<43> ,
  \data<44> ,
  \data<41> ,
  \data<42> ,
  \data<17> ,
  \data<18> ,
  \data<15> ,
  \count<0> ,
  \data<16> ,
  \count<3> ,
  \data<19> ,
  \count<1> ,
  \count<2> ,
  \data<10> ,
  \data<13> ,
  \data<14> ,
  \data<11> ,
  \data<12> ,
  \data<27> ,
  \data<28> ,
  \data<25> ,
  \data<26> ,
  \data<29> ,
  \data<20> ,
  \data<23> ,
  \data<24> ,
  \data<21> ,
  \data<22> ,
  \C<0> ,
  \C<1> ,
  \C<2> ,
  \C<3> ,
  \C<4> ,
  \C<5> ,
  \C<6> ,
  \C<7> ,
  \C<8> ,
  \C<9> ,
  \inreg<12> ,
  \inreg<11> ,
  \inreg<14> ,
  \inreg<13> ,
  \inreg<10> ,
  \inreg<19> ,
  \inreg<16> ,
  \inreg<15> ,
  \inreg<18> ,
  \inreg<17> ,
  \inreg<22> ,
  \inreg<21> ,
  \inreg<24> ,
  \inreg<23> ,
  \inreg<20> ,
  \inreg<29> ,
  \inreg<26> ,
  \inreg<25> ,
  \outreg<9> ,
  \inreg<28> ,
  \inreg<27> ,
  \inreg<32> ,
  \inreg<31> ,
  \outreg<5> ,
  \inreg<34> ,
  \outreg<6> ,
  \inreg<33> ,
  \outreg<7> ,
  \outreg<8> ,
  \outreg<1> ,
  \inreg<30> ,
  \outreg<2> ,
  \outreg<3> ,
  \outreg<4> ,
  \inreg<39> ,
  \inreg<36> ,
  \outreg<0> ,
  \inreg<35> ,
  \inreg<38> ,
  \inreg<37> ,
  \inreg<42> ,
  \inreg<41> ,
  \inreg<44> ,
  \inreg<43> ,
  \inreg<40> ,
  \inreg<49> ,
  \inreg<46> ,
  \inreg<45> ,
  \encrypt_mode<0> ,
  \inreg<48> ,
  \inreg<47> ,
  \inreg<52> ,
  \inreg<51> ,
  \inreg<54> ,
  \inreg<53> ,
  \inreg<50> ,
  \inreg<55> ,
  \data<57> ,
  \data<58> ,
  \data<55> ,
  \data<56> ,
  \encrypt<0> ,
  \data<59> ,
  \data<50> ,
  \data<53> ,
  \data<54> ,
  \data<51> ,
  \data<52> ,
  \data<60> ;
output
  \data_new<25> ,
  \inreg_new<45> ,
  \data_new<26> ,
  \data_new<13> ,
  \data_new<14> ,
  \data_new<11> ,
  \inreg_new<49> ,
  \data_new<12> ,
  \inreg_new<30> ,
  \outreg_new<11> ,
  \count_new<0> ,
  \outreg_new<12> ,
  \data_new<10> ,
  \outreg_new<13> ,
  \outreg_new<14> ,
  \inreg_new<34> ,
  \count_new<3> ,
  \inreg_new<33> ,
  \inreg_new<32> ,
  \count_new<1> ,
  \data_new<19> ,
  \inreg_new<31> ,
  \count_new<2> ,
  \outreg_new<10> ,
  \inreg_new<38> ,
  \outreg_new<19> ,
  \data_new<17> ,
  \inreg_new<37> ,
  \data_new<18> ,
  \inreg_new<36> ,
  \data_new<15> ,
  \inreg_new<35> ,
  \data_new<16> ,
  \outreg_new<15> ,
  \outreg_new<16> ,
  \outreg_new<17> ,
  \inreg_new<39> ,
  \outreg_new<18> ,
  \outreg_new<21> ,
  \outreg_new<22> ,
  \outreg_new<23> ,
  \outreg_new<24> ,
  \outreg_new<20> ,
  \outreg_new<29> ,
  \outreg_new<25> ,
  \outreg_new<26> ,
  \outreg_new<27> ,
  \outreg_new<28> ,
  \outreg_new<31> ,
  \outreg_new<32> ,
  \outreg_new<33> ,
  \outreg_new<34> ,
  \outreg_new<30> ,
  \outreg_new<39> ,
  \outreg_new<35> ,
  \outreg_new<36> ,
  \outreg_new<37> ,
  \outreg_new<38> ,
  \outreg_new<41> ,
  \outreg_new<42> ,
  \outreg_new<43> ,
  \outreg_new<44> ,
  \outreg_new<40> ,
  \outreg_new<49> ,
  \outreg_new<45> ,
  \outreg_new<46> ,
  \outreg_new<47> ,
  \outreg_new<48> ,
  \C_new<23> ,
  \C_new<24> ,
  \C_new<21> ,
  \C_new<22> ,
  \C_new<20> ,
  \data_new<4> ,
  \data_new<3> ,
  \C_new<27> ,
  \data_new<2> ,
  \data_new<1> ,
  \C_new<25> ,
  \data_new<0> ,
  \C_new<26> ,
  \C_new<13> ,
  \C_new<14> ,
  \C_new<11> ,
  \C_new<12> ,
  \C_new<10> ,
  \data_new<9> ,
  \data_new<8> ,
  \data_new<7> ,
  \data_new<6> ,
  \data_new<5> ,
  \C_new<19> ,
  \C_new<17> ,
  \C_new<18> ,
  \C_new<15> ,
  \C_new<16> ,
  \D_new<13> ,
  \D_new<14> ,
  \D_new<11> ,
  \D_new<12> ,
  \D_new<10> ,
  \data_new<63> ,
  \data_new<61> ,
  \data_new<62> ,
  \D_new<19> ,
  \data_new<60> ,
  \D_new<17> ,
  \D_new<18> ,
  \D_new<15> ,
  \D_new<16> ,
  \D_new<23> ,
  \D_new<24> ,
  \D_new<21> ,
  \D_new<22> ,
  \D_new<20> ,
  \data_new<53> ,
  \data_new<54> ,
  \data_new<51> ,
  \data_new<52> ,
  \data_new<50> ,
  \D_new<27> ,
  \D_new<25> ,
  \D_new<26> ,
  \data_new<59> ,
  \data_new<57> ,
  \data_new<58> ,
  \data_new<55> ,
  \data_new<56> ,
  \D_new<7> ,
  \C_new<6> ,
  \D_new<8> ,
  \C_new<5> ,
  \D_new<5> ,
  \C_new<8> ,
  \D_new<6> ,
  \C_new<7> ,
  \C_new<9> ,
  \D_new<9> ,
  \D_new<0> ,
  \C_new<0> ,
  \D_new<3> ,
  \C_new<2> ,
  \D_new<4> ,
  \C_new<1> ,
  \D_new<1> ,
  \C_new<4> ,
  \D_new<2> ,
  \C_new<3> ,
  \inreg_new<50> ,
  \inreg_new<9> ,
  \inreg_new<54> ,
  \inreg_new<53> ,
  \inreg_new<52> ,
  \inreg_new<6> ,
  \inreg_new<51> ,
  \inreg_new<5> ,
  \inreg_new<8> ,
  \inreg_new<7> ,
  \inreg_new<2> ,
  \inreg_new<55> ,
  \inreg_new<1> ,
  \inreg_new<4> ,
  \inreg_new<3> ,
  \inreg_new<0> ,
  \encrypt_mode_new<0> ,
  \outreg_new<9> ,
  \outreg_new<51> ,
  \outreg_new<52> ,
  \outreg_new<53> ,
  \outreg_new<5> ,
  \outreg_new<54> ,
  \outreg_new<6> ,
  \outreg_new<7> ,
  \outreg_new<8> ,
  \outreg_new<1> ,
  \outreg_new<50> ,
  \outreg_new<2> ,
  \outreg_new<59> ,
  \outreg_new<3> ,
  \outreg_new<4> ,
  \outreg_new<55> ,
  \data_new<43> ,
  \outreg_new<56> ,
  \data_new<44> ,
  \outreg_new<0> ,
  \outreg_new<57> ,
  \data_new<41> ,
  \outreg_new<58> ,
  \data_new<42> ,
  \inreg_new<20> ,
  \outreg_new<61> ,
  \outreg_new<62> ,
  \data_new<40> ,
  \outreg_new<63> ,
  \inreg_new<24> ,
  \inreg_new<23> ,
  \inreg_new<22> ,
  \data_new<49> ,
  \inreg_new<21> ,
  \outreg_new<60> ,
  \inreg_new<28> ,
  \data_new<47> ,
  \inreg_new<27> ,
  \data_new<48> ,
  \inreg_new<26> ,
  \data_new<45> ,
  \inreg_new<25> ,
  \data_new<46> ,
  \data_new<33> ,
  \data_new<34> ,
  \data_new<31> ,
  \inreg_new<29> ,
  \data_new<32> ,
  \inreg_new<10> ,
  \data_new<30> ,
  \inreg_new<14> ,
  \inreg_new<13> ,
  \inreg_new<12> ,
  \data_new<39> ,
  \inreg_new<11> ,
  \inreg_new<18> ,
  \data_new<37> ,
  \inreg_new<17> ,
  \data_new<38> ,
  \inreg_new<16> ,
  \data_new<35> ,
  \inreg_new<15> ,
  \data_new<36> ,
  \data_new<23> ,
  \data_new<24> ,
  \data_new<21> ,
  \inreg_new<19> ,
  \data_new<22> ,
  \inreg_new<40> ,
  \data_new<20> ,
  \inreg_new<44> ,
  \inreg_new<43> ,
  \inreg_new<42> ,
  \data_new<29> ,
  \inreg_new<41> ,
  \inreg_new<48> ,
  \data_new<27> ,
  \inreg_new<47> ,
  \data_new<28> ,
  \inreg_new<46> ;
wire
  \$$COND258<0>226.1 ,
  \$$COND348<0>376.1 ,
  \$$COND327<0>376.1 ,
  \$$COND216<0>226.1 ,
  \$$COND516<0>526.1 ,
  \$$COND235<0>226.1 ,
  \$$COND365<0>376.1 ,
  \$$COND180<0>151.1 ,
  \$$COND6<0>1.1 ,
  \[189] ,
  \$$COND391<0>451.1 ,
  \$$COND460<0>526.1 ,
  \$$COND56<0>1.1 ,
  \[190] ,
  \[191] ,
  \[192] ,
  \[193] ,
  \main_1/preS<28>0.1 ,
  \[194] ,
  \[195] ,
  \main_1/S7_1/$S7<3>526.1 ,
  \[196] ,
  \$$COND289<0>301.1 ,
  \main_1/preS<11>0.1 ,
  \[197] ,
  \[198] ,
  \$$COND403<0>451.1 ,
  \$$COND424<0>451.1 ,
  \$$COND349<0>376.1 ,
  \$$COND328<0>376.1 ,
  \$$COND517<0>526.1 ,
  \[199] ,
  \$$COND319<0>301.1 ,
  \$$COND521<0>601.1 ,
  \main_1/preS<7>0.1 ,
  \$$COND461<0>526.1 ,
  \$$COND480<0>526.1 ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \main_1/S2_1/$S2<1>151.1 ,
  \[5] ,
  \[6] ,
  \[7] ,
  \$$COND269<0>301.1 ,
  \[8] ,
  \[9] ,
  \$$COND402<0>451.1 ,
  \$$COND444<0>451.1 ,
  \$$COND329<0>376.1 ,
  \$$COND218<0>226.1 ,
  \$$COND518<0>526.1 ,
  \$$COND388<0>376.1 ,
  \$$COND237<0>226.1 ,
  \$$COND310<0>301.1 ,
  \main_1/preS<24>0.1 ,
  \main_1/S0_1/$S0<2>1.1 ,
  \$$COND481<0>526.1 ,
  \main_1/S3_1/$S3<3>226.1 ,
  \main_1/S4_1/$S4<2>301.1 ,
  \$$COND44<0>1.1 ,
  \main_1/S1_1/$S1<3>76.1 ,
  \$$COND34<0>1.1 ,
  \$$COND24<0>1.1 ,
  \main_1/preS<36>0.1 ,
  \$$COND401<0>451.1 ,
  \$$COND238<0>226.1 ,
  \$$COND368<0>376.1 ,
  \$$COND195<0>226.1 ,
  \$$COND96<0>76.1 ,
  \$$COND463<0>526.1 ,
  \$$COND482<0>526.1 ,
  \$$COND95<0>76.1 ,
  \$$COND98<0>76.1 ,
  \main_1/preS<20>0.1 ,
  \$$COND99<0>76.1 ,
  \$$COND45<0>1.1 ,
  \main_1/preS<2>0.1 ,
  \$$COND25<0>1.1 ,
  \$$COND15<0>1.1 ,
  \main_1/preS<32>0.1 ,
  \$$COND421<0>451.1 ,
  \$$COND92<0>76.1 ,
  \$$COND142<0>151.1 ,
  \$$COND163<0>151.1 ,
  \$$COND239<0>226.1 ,
  \$$COND196<0>226.1 ,
  \$$COND94<0>76.1 ,
  \$$COND93<0>76.1 ,
  \$$COND5<0>1.1 ,
  \$$COND464<0>526.1 ,
  \$$COND55<0>1.1 ,
  \main_1/S5_1/$S5<0>376.1 ,
  \$$COND417<0>451.1 ,
  \$$COND438<0>451.1 ,
  \$$COND141<0>151.1 ,
  \$$COND162<0>151.1 ,
  \$$COND183<0>151.1 ,
  \$$COND197<0>226.1 ,
  \main_1/preS<45>0.1 ,
  \$$COND105<0>76.1 ,
  \$$COND76<0>76.1 ,
  \$$COND108<0>76.1 ,
  \$$COND465<0>526.1 ,
  \$$COND484<0>526.1 ,
  \$$COND107<0>76.1 ,
  \$$COND77<0>76.1 ,
  \$$COND109<0>76.1 ,
  \$$COND79<0>76.1 ,
  \$$COND100<0>76.1 ,
  \$$COND284<0>301.1 ,
  \$$COND70<0>76.1 ,
  \$$COND101<0>76.1 ,
  \$$COND416<0>451.1 ,
  \$$COND137<0>151.1 ,
  \$$COND308<0>301.1 ,
  \$$COND158<0>151.1 ,
  \$$COND182<0>151.1 ,
  \$$COND71<0>76.1 ,
  \$$COND198<0>226.1 ,
  \$$COND103<0>76.1 ,
  \$$COND74<0>76.1 ,
  \$$COND73<0>76.1 ,
  \$$COND115<0>76.1 ,
  \main_1/preS<18>0.1 ,
  \$$COND118<0>76.1 ,
  \$$COND466<0>526.1 ,
  \$$COND485<0>526.1 ,
  \$$COND85<0>76.1 ,
  \$$COND117<0>76.1 ,
  \$$COND88<0>76.1 ,
  \main_1/preS<41>0.1 ,
  \$$COND89<0>76.1 ,
  \main_1/S4_1/$S4<1>301.1 ,
  \$$COND43<0>1.1 ,
  \main_1/S6_1/$S6<0>451.1 ,
  \$$COND110<0>76.1 ,
  \$$COND13<0>1.1 ,
  \$$COND80<0>76.1 ,
  \$$COND264<0>301.1 ,
  \$$COND112<0>76.1 ,
  \$$COND415<0>451.1 ,
  \$$COND436<0>451.1 ,
  \$$COND136<0>151.1 ,
  \$$COND82<0>76.1 ,
  \$$COND307<0>301.1 ,
  \$$COND157<0>151.1 ,
  \$$COND313<0>301.1 ,
  \$$COND81<0>76.1 ,
  \$$COND113<0>76.1 ,
  \$$COND84<0>76.1 ,
  \$$COND126<0>76.1 ,
  \$$COND128<0>76.1 ,
  \$$COND467<0>526.1 ,
  \$$COND127<0>76.1 ,
  \$$COND63<0>1.1 ,
  \[200] ,
  \$$COND53<0>1.1 ,
  \[201] ,
  \[202] ,
  \main_1/preS<14>0.1 ,
  \[203] ,
  \[204] ,
  \[205] ,
  \[206] ,
  \$$COND282<0>301.1 ,
  \$$COND122<0>76.1 ,
  \main_1/preS<6>0.1 ,
  \[207] ,
  \$$COND121<0>76.1 ,
  \[208] ,
  \$$COND331<0>376.1 ,
  \$$COND435<0>451.1 ,
  \$$COND135<0>151.1 ,
  \$$COND156<0>151.1 ,
  \$$COND177<0>151.1 ,
  \$$COND124<0>76.1 ,
  \[209] ,
  \$$COND123<0>76.1 ,
  \$$COND487<0>526.1 ,
  \$$COND65<0>76.1 ,
  \$$COND68<0>76.1 ,
  \$$COND8<0>1.1 ,
  \[210] ,
  \[211] ,
  \$$COND69<0>76.1 ,
  \[212] ,
  \[213] ,
  \[214] ,
  \main_1/preS<27>0.1 ,
  \[215] ,
  \[216] ,
  \$$COND281<0>301.1 ,
  \[217] ,
  \main_1/S0_1/$S0<3>1.1 ,
  \[218] ,
  \main_1/preS<10>0.1 ,
  \$$COND220<0>226.1 ,
  \$$COND305<0>301.1 ,
  \$$COND370<0>376.1 ,
  \$$COND176<0>151.1 ,
  \[219] ,
  \$$COND311<0>301.1 ,
  \main_1/preS<39>0.1 ,
  \$$COND469<0>526.1 ,
  \$$COND488<0>526.1 ,
  \[220] ,
  \[221] ,
  \[222] ,
  \[223] ,
  \[224] ,
  \[225] ,
  \[226] ,
  \$$COND261<0>301.1 ,
  \[227] ,
  \[228] ,
  \$$COND371<0>376.1 ,
  \$$COND175<0>151.1 ,
  \[229] ,
  \main_1/S2_1/$S2<3>151.1 ,
  \main_1/preS<23>0.1 ,
  \main_1/S5_1/$S5<2>376.1 ,
  \[230] ,
  \[231] ,
  \[232] ,
  \main_1/preS<35>0.1 ,
  \[233] ,
  \[234] ,
  \[235] ,
  \$$COND42<0>1.1 ,
  \[236] ,
  \$$COND277<0>301.1 ,
  \[237] ,
  \$$COND22<0>1.1 ,
  \[238] ,
  \$$COND419<0>451.1 ,
  \$$COND334<0>376.1 ,
  \$$COND12<0>1.1 ,
  \$$COND222<0>226.1 ,
  \$$COND372<0>376.1 ,
  \$$COND351<0>376.1 ,
  \[239] ,
  \$$COND0<0>1.1 ,
  \[240] ,
  \[241] ,
  \[242] ,
  \[243] ,
  \$$COND62<0>1.1 ,
  \[244] ,
  \[245] ,
  \main_1/preS<1>0.1 ,
  \$$COND276<0>301.1 ,
  \$$COND335<0>376.1 ,
  \$$COND439<0>451.1 ,
  \$$COND139<0>151.1 ,
  \main_1/preS<31>0.1 ,
  \$$COND352<0>376.1 ,
  \$$COND200<0>226.1 ,
  \$$COND500<0>526.1 ,
  \main_1/S6_1/$S6<2>451.1 ,
  \$$COND275<0>301.1 ,
  \$$COND298<0>301.1 ,
  \$$COND430<0>451.1 ,
  \$$COND130<0>151.1 ,
  \$$COND224<0>226.1 ,
  \$$COND374<0>376.1 ,
  \$$COND159<0>151.1 ,
  \$$COND243<0>226.1 ,
  \$$COND201<0>226.1 ,
  \$$COND501<0>526.1 ,
  \main_1/preS<44>0.1 ,
  \main_1/S7_1/$S7<0>526.1 ,
  \main_1/S1_1/$S1<1>76.1 ,
  \$$COND297<0>301.1 ,
  \$$COND337<0>376.1 ,
  \$$COND225<0>226.1 ,
  \$$COND300<0>301.1 ,
  \$$COND450<0>451.1 ,
  \$$COND150<0>151.1 ,
  \$$COND244<0>226.1 ,
  \$$COND354<0>376.1 ,
  \$$COND179<0>151.1 ,
  \$$COND202<0>226.1 ,
  \main_1/preS<17>0.1 ,
  \main_1/S5_1/$S5<1>376.1 ,
  \main_1/preS<40>0.1 ,
  \main_1/preS<9>0.1 ,
  \$$COND296<0>301.1 ,
  \main_1/S3_1/$S3<0>226.1 ,
  \$$COND338<0>376.1 ,
  \main_1/S4_1/$S4<3>301.1 ,
  \$$COND226<0>226.1 ,
  \$$COND376<0>376.1 ,
  \$$COND355<0>376.1 ,
  \$$COND170<0>151.1 ,
  \$$COND41<0>1.1 ,
  \$$COND11<0>1.1 ,
  \$$COND491<0>526.1 ,
  \$$COND520<0>0.1 ,
  \main_1/S0_1/$S0<0>1.1 ,
  \main_1/preS<13>0.1 ,
  \$$COND295<0>301.1 ,
  \$$COND414<0>451.1 ,
  \$$COND339<0>376.1 ,
  \main_1/preS<5>0.1 ,
  \$$COND227<0>226.1 ,
  \$$COND377<0>376.1 ,
  \$$COND246<0>226.1 ,
  \$$COND190<0>151.1 ,
  \$$COND398<0>451.1 ,
  \$$COND492<0>526.1 ,
  \main_1/S6_1/$S6<1>451.1 ,
  \main_1/S1_1/$S1<0>76.1 ,
  \$$COND279<0>301.1 ,
  \main_1/preS<26>0.1 ,
  \$$COND413<0>451.1 ,
  \$$COND134<0>151.1 ,
  \$$COND228<0>226.1 ,
  \$$COND378<0>376.1 ,
  \$$COND247<0>226.1 ,
  \$$COND357<0>376.1 ,
  \$$COND320<0>301.1 ,
  \$$COND505<0>526.1 ,
  \$$COND397<0>451.1 ,
  \$$COND493<0>526.1 ,
  \$$COND470<0>526.1 ,
  \main_1/preS<38>0.1 ,
  \$$COND49<0>1.1 ,
  \$$COND39<0>1.1 ,
  \$$COND270<0>301.1 ,
  \$$COND29<0>1.1 ,
  \$$COND133<0>151.1 ,
  \$$COND229<0>226.1 ,
  \$$COND304<0>301.1 ,
  \$$COND379<0>376.1 ,
  \$$COND358<0>376.1 ,
  \$$COND206<0>226.1 ,
  \$$COND506<0>526.1 ,
  \main_1/preS<22>0.1 ,
  \generate_key_1/freeze<0>605.1 ,
  \$$COND59<0>1.1 ,
  \main_1/preS<34>0.1 ,
  \$$COND408<0>451.1 ,
  \$$COND411<0>451.1 ,
  \$$COND432<0>451.1 ,
  \$$COND132<0>151.1 ,
  \$$COND303<0>301.1 ,
  \$$COND453<0>451.1 ,
  \$$COND153<0>151.1 ,
  \$$COND249<0>226.1 ,
  \$$COND359<0>376.1 ,
  \$$COND174<0>151.1 ,
  \$$COND207<0>226.1 ,
  \main_1/S1_1/$S1<2>76.1 ,
  \main_1/S7_1/$S7<2>526.1 ,
  \$$COND40<0>1.1 ,
  \$$COND472<0>526.1 ,
  \$$COND30<0>1.1 ,
  \$$COND20<0>1.1 ,
  \$$COND10<0>1.1 ,
  \$$COND2<0>1.1 ,
  \main_1/preS<47>0.1 ,
  \main_1/preS<4>0.1 ,
  \$$COND428<0>451.1 ,
  \$$COND431<0>451.1 ,
  \$$COND302<0>301.1 ,
  \$$COND452<0>451.1 ,
  \$$COND152<0>151.1 ,
  \$$COND173<0>151.1 ,
  \$$COND208<0>226.1 ,
  \$$COND508<0>526.1 ,
  \main_1/preS<30>0.1 ,
  \$$COND60<0>1.1 ,
  \$$COND496<0>526.1 ,
  \$$COND473<0>526.1 ,
  \main_1/S3_1/$S3<2>226.1 ,
  \[10] ,
  \$$COND406<0>451.1 ,
  \[11] ,
  \$$COND427<0>451.1 ,
  \$$COND301<0>301.1 ,
  \$$COND193<0>151.1 ,
  \[12] ,
  \[13] ,
  \$$COND9<0>1.1 ,
  \[14] ,
  \[15] ,
  \$$COND497<0>526.1 ,
  \main_1/preS<43>0.1 ,
  \$$COND455<0>526.1 ,
  \[16] ,
  \main_1/preS<0>0.1 ,
  \[17] ,
  \[18] ,
  \[19] ,
  \$$COND274<0>301.1 ,
  \[20] ,
  \$$COND48<0>1.1 ,
  \[21] ,
  \$$COND426<0>451.1 ,
  \$$COND447<0>451.1 ,
  \$$COND147<0>151.1 ,
  \$$COND168<0>151.1 ,
  \[22] ,
  \$$COND323<0>301.1 ,
  \$$COND28<0>1.1 ,
  \[23] ,
  \$$COND18<0>1.1 ,
  \[24] ,
  \[25] ,
  \$$COND498<0>526.1 ,
  \[26] ,
  \$$COND475<0>526.1 ,
  \[27] ,
  \[28] ,
  \main_1/preS<16>0.1 ,
  \[100] ,
  \[29] ,
  \[101] ,
  \[102] ,
  \[103] ,
  \[104] ,
  \main_1/S2_1/$S2<0>151.1 ,
  \[105] ,
  \[106] ,
  \[107] ,
  \$$COND58<0>1.1 ,
  \[30] ,
  \main_1/S5_1/$S5<3>376.1 ,
  \[108] ,
  \[31] ,
  \$$COND425<0>451.1 ,
  \$$COND340<0>376.1 ,
  \$$COND446<0>451.1 ,
  \$$COND146<0>151.1 ,
  \$$COND167<0>151.1 ,
  \$$COND188<0>151.1 ,
  \[109] ,
  \$$COND191<0>151.1 ,
  \[32] ,
  \$$COND322<0>301.1 ,
  \[33] ,
  \$$COND399<0>451.1 ,
  \[34] ,
  \[35] ,
  \$$COND499<0>526.1 ,
  \[36] ,
  \$$COND476<0>526.1 ,
  \[37] ,
  \main_1/S7_1/$S7<1>526.1 ,
  \[38] ,
  \[110] ,
  \[39] ,
  \[111] ,
  \main_1/preS<29>0.1 ,
  \[112] ,
  \[113] ,
  \[114] ,
  \[115] ,
  \main_1/preS<12>0.1 ,
  \[116] ,
  \$$COND272<0>301.1 ,
  \[117] ,
  \[40] ,
  \[118] ,
  \[41] ,
  \$$COND251<0>226.1 ,
  \$$COND341<0>376.1 ,
  \$$COND445<0>451.1 ,
  \$$COND187<0>151.1 ,
  \[119] ,
  \[42] ,
  \main_1/preS<8>0.1 ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \$$COND477<0>526.1 ,
  \[47] ,
  \[48] ,
  \[120] ,
  \[49] ,
  \[121] ,
  \[122] ,
  \[123] ,
  \[124] ,
  \[125] ,
  \[126] ,
  \$$COND288<0>301.1 ,
  \main_1/S3_1/$S3<1>226.1 ,
  \$$COND271<0>301.1 ,
  \[127] ,
  \[50] ,
  \main_1/preS<25>0.1 ,
  \[128] ,
  \[51] ,
  \$$COND342<0>376.1 ,
  \$$COND210<0>226.1 ,
  \$$COND510<0>526.1 ,
  \$$COND380<0>376.1 ,
  \$$COND165<0>151.1 ,
  \main_1/S6_1/$S6<3>451.1 ,
  \[129] ,
  \[52] ,
  \[53] ,
  \main_1/S0_1/$S0<1>1.1 ,
  \[54] ,
  \[55] ,
  \$$COND459<0>526.1 ,
  \[56] ,
  \[57] ,
  \[58] ,
  \main_1/preS<37>0.1 ,
  \[130] ,
  \[59] ,
  \[131] ,
  \[132] ,
  \[133] ,
  \[134] ,
  \[135] ,
  \[136] ,
  \$$COND287<0>301.1 ,
  \[137] ,
  \[60] ,
  \[138] ,
  \$$COND409<0>451.1 ,
  \[61] ,
  \$$COND253<0>226.1 ,
  \$$COND211<0>226.1 ,
  \$$COND511<0>526.1 ,
  \$$COND381<0>376.1 ,
  \$$COND360<0>376.1 ,
  \$$COND185<0>151.1 ,
  \[139] ,
  \[62] ,
  \$$COND317<0>301.1 ,
  \[63] ,
  \[64] ,
  \[65] ,
  \$$COND37<0>1.1 ,
  \[66] ,
  \$$COND479<0>526.1 ,
  \$$COND27<0>1.1 ,
  \[67] ,
  \main_1/preS<21>0.1 ,
  \$$COND17<0>1.1 ,
  \[68] ,
  \[140] ,
  \[69] ,
  \[141] ,
  \generate_key_1/shift_by_one<0>605.1 ,
  \[142] ,
  \[143] ,
  \[144] ,
  \[145] ,
  \main_1/preS<33>0.1 ,
  \[146] ,
  \$$COND286<0>301.1 ,
  \$$COND267<0>301.1 ,
  \[147] ,
  \[70] ,
  \[148] ,
  \$$COND400<0>451.1 ,
  \[71] ,
  \$$COND254<0>226.1 ,
  \$$COND429<0>451.1 ,
  \$$COND512<0>526.1 ,
  \$$COND382<0>376.1 ,
  \$$COND231<0>226.1 ,
  \[149] ,
  \[72] ,
  \$$COND316<0>301.1 ,
  \[73] ,
  \$$COND57<0>1.1 ,
  \[74] ,
  \[75] ,
  \[76] ,
  \[77] ,
  \[78] ,
  \[150] ,
  \[79] ,
  \[151] ,
  \[152] ,
  \main_1/S4_1/$S4<0>301.1 ,
  \[153] ,
  \[154] ,
  \[155] ,
  \[156] ,
  \$$COND266<0>301.1 ,
  \$$COND291<0>301.1 ,
  \[157] ,
  \[80] ,
  \main_1/preS<46>0.1 ,
  \[158] ,
  \[81] ,
  \$$COND255<0>226.1 ,
  \$$COND345<0>376.1 ,
  \$$COND449<0>451.1 ,
  \$$COND149<0>151.1 ,
  \$$COND213<0>226.1 ,
  \$$COND513<0>526.1 ,
  \$$COND232<0>226.1 ,
  \main_1/preS<3>0.1 ,
  \[159] ,
  \[82] ,
  \$$COND315<0>301.1 ,
  \[83] ,
  \$$COND394<0>451.1 ,
  \[84] ,
  \[85] ,
  \[86] ,
  \[87] ,
  \[88] ,
  \[160] ,
  \main_1/S2_1/$S2<2>151.1 ,
  \[89] ,
  \[161] ,
  \[162] ,
  \[163] ,
  \[164] ,
  \[165] ,
  \[166] ,
  \$$COND265<0>301.1 ,
  \[167] ,
  \[90] ,
  \[168] ,
  \[91] ,
  \$$COND256<0>226.1 ,
  \$$COND346<0>376.1 ,
  \$$COND140<0>151.1 ,
  \$$COND440<0>451.1 ,
  \$$COND325<0>376.1 ,
  \$$COND214<0>226.1 ,
  \$$COND384<0>376.1 ,
  \$$COND233<0>226.1 ,
  \$$COND363<0>376.1 ,
  \[169] ,
  \[92] ,
  \[93] ,
  \$$COND393<0>451.1 ,
  \main_1/preS<19>0.1 ,
  \[94] ,
  \[95] ,
  \[96] ,
  \[97] ,
  \main_1/preS<42>0.1 ,
  \[98] ,
  \[170] ,
  \[99] ,
  \[171] ,
  \[172] ,
  \[173] ,
  \[174] ,
  \[175] ,
  \[176] ,
  \[177] ,
  \[178] ,
  \$$COND347<0>376.1 ,
  \$$COND215<0>226.1 ,
  \$$COND515<0>526.1 ,
  \$$COND385<0>376.1 ,
  \$$COND160<0>151.1 ,
  \$$COND234<0>226.1 ,
  \$$COND364<0>376.1 ,
  \$$COND189<0>151.1 ,
  \[179] ,
  \$$COND46<0>1.1 ,
  \$$COND36<0>1.1 ,
  \[180] ,
  \main_1/preS<15>0.1 ,
  \$$COND26<0>1.1 ,
  \[181] ,
  \[182] ,
  \[183] ,
  \[184] ,
  \[185] ,
  \[186] ,
  \[187] ,
  \[188] ,
  \$$COND404<0>451.1 ;
assign
  \$$COND258<0>226.1  = \main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND348<0>376.1  = \main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \data_new<25>  = \[159] ,
  \$$COND327<0>376.1  = ~\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \$$COND216<0>226.1  = \main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND516<0>526.1  = \main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \inreg_new<45>  = \[11] ,
  \$$COND235<0>226.1  = ~\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND365<0>376.1  = ~\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND180<0>151.1  = \main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \$$COND6<0>1.1  = ~\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \[189]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<25>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<1>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<26>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<0>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<48>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<27>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<27>  & ~\$$COND521<0>601.1 )))))))),
  \data_new<26>  = \[158] ,
  \data_new<13>  = \[171] ,
  \$$COND391<0>451.1  = ~\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \data_new<14>  = \[170] ,
  \data_new<11>  = \[173] ,
  \$$COND460<0>526.1  = ~\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \inreg_new<49>  = \[7] ,
  \data_new<12>  = \[172] ,
  \inreg_new<30>  = \[26] ,
  \$$COND56<0>1.1  = \main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \outreg_new<11>  = \[109] ,
  \count_new<0>  = \[188] ,
  \outreg_new<12>  = \[108] ,
  \data_new<10>  = \[174] ,
  \[190]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<24>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<0>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<25>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<27>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<35>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<27>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<26>  & ~\$$COND521<0>601.1 )))))))),
  \outreg_new<13>  = \[107] ,
  \[191]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<23>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<27>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<24>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<26>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<43>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<35>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<25>  & ~\$$COND521<0>601.1 )))))))),
  \outreg_new<14>  = \[106] ,
  \inreg_new<34>  = \[22] ,
  \[192]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<22>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<26>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<23>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<25>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<51>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<43>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<24>  & ~\$$COND521<0>601.1 )))))))),
  \count_new<3>  = \[185] ,
  \inreg_new<33>  = \[23] ,
  \[193]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<21>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<25>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<22>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<24>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<51>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<23>  & ~\$$COND521<0>601.1 ))) | (~\reset<0>  & (~\encrypt<0>  & (\data_in<2>  & \$$COND521<0>601.1 )))))))),
  \main_1/preS<28>0.1  = (~\data<51>  & \D<18> ) | (\data<51>  & ~\D<18> ),
  \inreg_new<32>  = \[24] ,
  \[194]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<20>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<24>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<21>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<23>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<2>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<22>  & ~\$$COND521<0>601.1 ))) | (~\reset<0>  & (\encrypt<0>  & (\data_in<2>  & \$$COND521<0>601.1 )))))))),
  \count_new<1>  = \[187] ,
  \data_new<19>  = \[165] ,
  \inreg_new<31>  = \[25] ,
  \[195]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<19>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<23>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<20>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<22>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<2>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<10>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<21>  & ~\$$COND521<0>601.1 )))))))),
  \count_new<2>  = \[186] ,
  \outreg_new<10>  = \[110] ,
  \main_1/S7_1/$S7<3>526.1  = (~\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 ))))) | ((~\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & \main_1/preS<42>0.1 ))))) | ((\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/preS<42>0.1 ))))) | ((\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 ))))) | (\$$COND518<0>526.1  | (\$$COND513<0>526.1  | (\$$COND512<0>526.1  | (\$$COND511<0>526.1  | (\$$COND510<0>526.1  | (\$$COND508<0>526.1  | (\$$COND505<0>526.1  | (\$$COND499<0>526.1  | (\$$COND498<0>526.1  | (\$$COND497<0>526.1  | (\$$COND493<0>526.1  | (\$$COND492<0>526.1  | (\$$COND491<0>526.1  | (\$$COND488<0>526.1  | (\$$COND485<0>526.1  | (\$$COND484<0>526.1  | (\$$COND482<0>526.1  | (\$$COND479<0>526.1  | (\$$COND475<0>526.1  | (\$$COND473<0>526.1  | (\$$COND472<0>526.1  | (\$$COND469<0>526.1  | (\$$COND466<0>526.1  | (\$$COND464<0>526.1  | (\$$COND463<0>526.1  | (\$$COND461<0>526.1  | (\$$COND460<0>526.1  | \$$COND455<0>526.1 )))))))))))))))))))))))))))))),
  \inreg_new<38>  = \[18] ,
  \[196]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<18>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<22>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<19>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<21>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<18>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<10>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<20>  & ~\$$COND521<0>601.1 )))))))),
  \$$COND289<0>301.1  = \main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \outreg_new<19>  = \[101] ,
  \data_new<17>  = \[167] ,
  \inreg_new<37>  = \[19] ,
  \main_1/preS<11>0.1  = (~\data<40>  & \C<9> ) | (\data<40>  & ~\C<9> ),
  \[197]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<17>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<21>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<18>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<20>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<26>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<18>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<19>  & ~\$$COND521<0>601.1 )))))))),
  \data_new<18>  = \[166] ,
  \inreg_new<36>  = \[20] ,
  \[198]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<16>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<20>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<17>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<19>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<34>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<26>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<18>  & ~\$$COND521<0>601.1 )))))))),
  \$$COND403<0>451.1  = ~\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \$$COND424<0>451.1  = ~\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND349<0>376.1  = \main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \data_new<15>  = \[169] ,
  \$$COND328<0>376.1  = ~\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \$$COND517<0>526.1  = \main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \inreg_new<35>  = \[21] ,
  \[199]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<15>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<19>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<16>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<18>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<42>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<34>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<17>  & ~\$$COND521<0>601.1 )))))))),
  \$$COND319<0>301.1  = \main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \data_new<16>  = \[168] ,
  \outreg_new<15>  = \[105] ,
  \$$COND521<0>601.1  = \load_key<0>  & (\count<3>  & (\count<2>  & (\count<1>  & \count<0> ))),
  \outreg_new<16>  = \[104] ,
  \main_1/preS<7>0.1  = (~\data<36>  & \C<27> ) | (\data<36>  & ~\C<27> ),
  \outreg_new<17>  = \[103] ,
  \$$COND461<0>526.1  = ~\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \inreg_new<39>  = \[17] ,
  \$$COND480<0>526.1  = \main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \outreg_new<18>  = \[102] ,
  \outreg_new<21>  = \[99] ,
  \outreg_new<22>  = \[98] ,
  \[1]  = (\inreg<55>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<47>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \outreg_new<23>  = \[97] ,
  \[2]  = (\inreg<54>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<46>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \outreg_new<24>  = \[96] ,
  \[3]  = (\inreg<53>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<45>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[4]  = (\inreg<52>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<44>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \main_1/S2_1/$S2<1>151.1  = (~\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & \main_1/preS<12>0.1 ))))) | ((~\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 ))))) | ((\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 ))))) | ((\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & \main_1/preS<12>0.1 ))))) | (\$$COND190<0>151.1  | (\$$COND189<0>151.1  | (\$$COND188<0>151.1  | (\$$COND187<0>151.1  | (\$$COND185<0>151.1  | (\$$COND182<0>151.1  | (\$$COND179<0>151.1  | (\$$COND177<0>151.1  | (\$$COND176<0>151.1  | (\$$COND175<0>151.1  | (\$$COND170<0>151.1  | (\$$COND168<0>151.1  | (\$$COND167<0>151.1  | (\$$COND163<0>151.1  | (\$$COND160<0>151.1  | (\$$COND159<0>151.1  | (\$$COND157<0>151.1  | (\$$COND153<0>151.1  | (\$$COND152<0>151.1  | (\$$COND150<0>151.1  | (\$$COND147<0>151.1  | (\$$COND142<0>151.1  | (\$$COND141<0>151.1  | (\$$COND136<0>151.1  | (\$$COND135<0>151.1  | (\$$COND134<0>151.1  | (\$$COND133<0>151.1  | \$$COND130<0>151.1 )))))))))))))))))))))))))))))),
  \[5]  = (\inreg<51>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<43>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[6]  = (\inreg<50>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<42>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \outreg_new<20>  = \[100] ,
  \[7]  = (\inreg<49>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<41>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \outreg_new<29>  = \[91] ,
  \$$COND269<0>301.1  = ~\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \[8]  = (\inreg<48>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<40>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[9]  = (\inreg<47>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<39>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND402<0>451.1  = ~\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \$$COND444<0>451.1  = \main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND329<0>376.1  = ~\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \$$COND218<0>226.1  = \main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND518<0>526.1  = \main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \$$COND388<0>376.1  = \main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND237<0>226.1  = ~\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND310<0>301.1  = \main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \main_1/preS<24>0.1  = (~\data<47>  & \D<12> ) | (\data<47>  & ~\D<12> ),
  \outreg_new<25>  = \[95] ,
  \outreg_new<26>  = \[94] ,
  \main_1/S0_1/$S0<2>1.1  = (~\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & \main_1/preS<0>0.1 ))))) | ((~\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 ))))) | ((\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & \main_1/preS<0>0.1 ))))) | ((\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 ))))) | (\$$COND63<0>1.1  | (\$$COND62<0>1.1  | (\$$COND5<0>1.1  | (\$$COND59<0>1.1  | (\$$COND56<0>1.1  | (\$$COND55<0>1.1  | (\$$COND49<0>1.1  | (\$$COND48<0>1.1  | (\$$COND46<0>1.1  | (\$$COND43<0>1.1  | (\$$COND41<0>1.1  | (\$$COND40<0>1.1  | (\$$COND37<0>1.1  | (\$$COND36<0>1.1  | (\$$COND34<0>1.1  | (\$$COND2<0>1.1  | (\$$COND29<0>1.1  | (\$$COND26<0>1.1  | (\$$COND25<0>1.1  | (\$$COND22<0>1.1  | (\$$COND20<0>1.1  | (\$$COND18<0>1.1  | (\$$COND17<0>1.1  | (\$$COND15<0>1.1  | (\$$COND12<0>1.1  | (\$$COND11<0>1.1  | (\$$COND10<0>1.1  | \$$COND0<0>1.1 )))))))))))))))))))))))))))))),
  \outreg_new<27>  = \[93] ,
  \$$COND481<0>526.1  = \main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \main_1/S3_1/$S3<3>226.1  = (~\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 ))))) | ((~\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & \main_1/preS<18>0.1 ))))) | ((\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 ))))) | ((\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & \main_1/preS<18>0.1 ))))) | (\$$COND258<0>226.1  | (\$$COND255<0>226.1  | (\$$COND254<0>226.1  | (\$$COND251<0>226.1  | (\$$COND249<0>226.1  | (\$$COND247<0>226.1  | (\$$COND244<0>226.1  | (\$$COND238<0>226.1  | (\$$COND235<0>226.1  | (\$$COND234<0>226.1  | (\$$COND232<0>226.1  | (\$$COND231<0>226.1  | (\$$COND229<0>226.1  | (\$$COND227<0>226.1  | (\$$COND226<0>226.1  | (\$$COND225<0>226.1  | (\$$COND224<0>226.1  | (\$$COND222<0>226.1  | (\$$COND216<0>226.1  | (\$$COND213<0>226.1  | (\$$COND211<0>226.1  | (\$$COND210<0>226.1  | (\$$COND208<0>226.1  | (\$$COND207<0>226.1  | (\$$COND202<0>226.1  | (\$$COND201<0>226.1  | (\$$COND197<0>226.1  | \$$COND196<0>226.1 )))))))))))))))))))))))))))))),
  \outreg_new<28>  = \[92] ,
  \main_1/S4_1/$S4<2>301.1  = (~\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & \main_1/preS<24>0.1 ))))) | ((~\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 ))))) | ((\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 ))))) | ((\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & \main_1/preS<24>0.1 ))))) | (\$$COND322<0>301.1  | (\$$COND317<0>301.1  | (\$$COND316<0>301.1  | (\$$COND315<0>301.1  | (\$$COND313<0>301.1  | (\$$COND311<0>301.1  | (\$$COND310<0>301.1  | (\$$COND307<0>301.1  | (\$$COND304<0>301.1  | (\$$COND303<0>301.1  | (\$$COND302<0>301.1  | (\$$COND300<0>301.1  | (\$$COND298<0>301.1  | (\$$COND297<0>301.1  | (\$$COND291<0>301.1  | (\$$COND286<0>301.1  | (\$$COND284<0>301.1  | (\$$COND282<0>301.1  | (\$$COND281<0>301.1  | (\$$COND279<0>301.1  | (\$$COND276<0>301.1  | (\$$COND274<0>301.1  | (\$$COND272<0>301.1  | (\$$COND271<0>301.1  | (\$$COND269<0>301.1  | (\$$COND267<0>301.1  | (\$$COND264<0>301.1  | \$$COND261<0>301.1 )))))))))))))))))))))))))))))),
  \outreg_new<31>  = \[89] ,
  \$$COND44<0>1.1  = ~\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \main_1/S1_1/$S1<3>76.1  = (~\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & \main_1/preS<10>0.1 ))))) | ((~\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & \main_1/preS<10>0.1 ))))) | ((\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 ))))) | ((\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 ))))) | (\$$COND98<0>76.1  | (\$$COND95<0>76.1  | (\$$COND94<0>76.1  | (\$$COND92<0>76.1  | (\$$COND89<0>76.1  | (\$$COND88<0>76.1  | (\$$COND85<0>76.1  | (\$$COND82<0>76.1  | (\$$COND80<0>76.1  | (\$$COND77<0>76.1  | (\$$COND76<0>76.1  | (\$$COND73<0>76.1  | (\$$COND70<0>76.1  | (\$$COND68<0>76.1  | (\$$COND65<0>76.1  | (\$$COND128<0>76.1  | (\$$COND127<0>76.1  | (\$$COND124<0>76.1  | (\$$COND121<0>76.1  | (\$$COND118<0>76.1  | (\$$COND115<0>76.1  | (\$$COND113<0>76.1  | (\$$COND112<0>76.1  | (\$$COND109<0>76.1  | (\$$COND107<0>76.1  | (\$$COND103<0>76.1  | (\$$COND101<0>76.1  | \$$COND100<0>76.1 )))))))))))))))))))))))))))))),
  \outreg_new<32>  = \[88] ,
  \$$COND34<0>1.1  = ~\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \outreg_new<33>  = \[87] ,
  \$$COND24<0>1.1  = \main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \main_1/preS<36>0.1  = (~\data<55>  & \D<15> ) | (\data<55>  & ~\D<15> ),
  \outreg_new<34>  = \[86] ,
  \outreg_new<30>  = \[90] ,
  \outreg_new<39>  = \[81] ,
  \$$COND401<0>451.1  = ~\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \$$COND238<0>226.1  = ~\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND368<0>376.1  = ~\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND195<0>226.1  = ~\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \outreg_new<35>  = \[85] ,
  \outreg_new<36>  = \[84] ,
  \$$COND96<0>76.1  = \main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \outreg_new<37>  = \[83] ,
  \$$COND463<0>526.1  = ~\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \$$COND482<0>526.1  = \main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \$$COND95<0>76.1  = \main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \outreg_new<38>  = \[82] ,
  \$$COND98<0>76.1  = ~\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \outreg_new<41>  = \[79] ,
  \outreg_new<42>  = \[78] ,
  \main_1/preS<20>0.1  = (~\data<45>  & \C<26> ) | (\data<45>  & ~\C<26> ),
  \outreg_new<43>  = \[77] ,
  \$$COND99<0>76.1  = \main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \outreg_new<44>  = \[76] ,
  \$$COND45<0>1.1  = ~\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \main_1/preS<2>0.1  = (~\data<33>  & \C<10> ) | (\data<33>  & ~\C<10> ),
  \$$COND25<0>1.1  = \main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \outreg_new<40>  = \[80] ,
  \$$COND15<0>1.1  = ~\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \outreg_new<49>  = \[71] ,
  \main_1/preS<32>0.1  = (~\data<53>  & \D<22> ) | (\data<53>  & ~\D<22> ),
  \$$COND421<0>451.1  = \main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \$$COND92<0>76.1  = \main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \$$COND142<0>151.1  = ~\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND163<0>151.1  = ~\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \$$COND239<0>226.1  = ~\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND196<0>226.1  = ~\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND94<0>76.1  = ~\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \outreg_new<45>  = \[75] ,
  \$$COND93<0>76.1  = ~\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \outreg_new<46>  = \[74] ,
  \$$COND5<0>1.1  = ~\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \outreg_new<47>  = \[73] ,
  \$$COND464<0>526.1  = ~\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \outreg_new<48>  = \[72] ,
  \$$COND55<0>1.1  = \main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \main_1/S5_1/$S5<0>376.1  = (~\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & \main_1/preS<30>0.1 ))))) | ((~\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 ))))) | ((\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & \main_1/preS<30>0.1 ))))) | ((\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 ))))) | (\$$COND388<0>376.1  | (\$$COND384<0>376.1  | (\$$COND381<0>376.1  | (\$$COND379<0>376.1  | (\$$COND378<0>376.1  | (\$$COND377<0>376.1  | (\$$COND374<0>376.1  | (\$$COND371<0>376.1  | (\$$COND370<0>376.1  | (\$$COND365<0>376.1  | (\$$COND364<0>376.1  | (\$$COND360<0>376.1  | (\$$COND359<0>376.1  | (\$$COND357<0>376.1  | (\$$COND355<0>376.1  | (\$$COND354<0>376.1  | (\$$COND351<0>376.1  | (\$$COND348<0>376.1  | (\$$COND347<0>376.1  | (\$$COND345<0>376.1  | (\$$COND342<0>376.1  | (\$$COND340<0>376.1  | (\$$COND339<0>376.1  | (\$$COND338<0>376.1  | (\$$COND335<0>376.1  | (\$$COND334<0>376.1  | (\$$COND329<0>376.1  | \$$COND328<0>376.1 )))))))))))))))))))))))))))))),
  \$$COND417<0>451.1  = \main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \$$COND438<0>451.1  = \main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND141<0>151.1  = ~\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND162<0>151.1  = ~\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \$$COND183<0>151.1  = \main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \$$COND197<0>226.1  = ~\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \main_1/preS<45>0.1  = (~\data<62>  & \D<7> ) | (\data<62>  & ~\D<7> ),
  \$$COND105<0>76.1  = ~\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \$$COND76<0>76.1  = \main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \$$COND108<0>76.1  = \main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \$$COND465<0>526.1  = ~\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \$$COND484<0>526.1  = \main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \$$COND107<0>76.1  = \main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \$$COND77<0>76.1  = ~\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \$$COND109<0>76.1  = ~\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \$$COND79<0>76.1  = \main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \$$COND100<0>76.1  = \main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \$$COND284<0>301.1  = \main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \$$COND70<0>76.1  = ~\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \$$COND101<0>76.1  = ~\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \$$COND416<0>451.1  = \main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \$$COND137<0>151.1  = ~\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND308<0>301.1  = \main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \$$COND158<0>151.1  = \main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND182<0>151.1  = \main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \$$COND71<0>76.1  = \main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \$$COND198<0>226.1  = ~\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND103<0>76.1  = \main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \$$COND74<0>76.1  = ~\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \$$COND73<0>76.1  = ~\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \$$COND115<0>76.1  = \main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \main_1/preS<18>0.1  = (~\data<43>  & \C<15> ) | (\data<43>  & ~\C<15> ),
  \$$COND118<0>76.1  = ~\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \$$COND466<0>526.1  = ~\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \$$COND485<0>526.1  = \main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \$$COND85<0>76.1  = ~\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \$$COND117<0>76.1  = ~\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \$$COND88<0>76.1  = \main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \main_1/preS<41>0.1  = (~\data<60>  & \D<24> ) | (\data<60>  & ~\D<24> ),
  \$$COND89<0>76.1  = ~\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \main_1/S4_1/$S4<1>301.1  = (~\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 ))))) | ((~\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & \main_1/preS<24>0.1 ))))) | ((\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 ))))) | ((\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & \main_1/preS<24>0.1 ))))) | (\$$COND323<0>301.1  | (\$$COND320<0>301.1  | (\$$COND317<0>301.1  | (\$$COND316<0>301.1  | (\$$COND313<0>301.1  | (\$$COND311<0>301.1  | (\$$COND308<0>301.1  | (\$$COND307<0>301.1  | (\$$COND305<0>301.1  | (\$$COND304<0>301.1  | (\$$COND300<0>301.1  | (\$$COND298<0>301.1  | (\$$COND296<0>301.1  | (\$$COND295<0>301.1  | (\$$COND291<0>301.1  | (\$$COND288<0>301.1  | (\$$COND287<0>301.1  | (\$$COND286<0>301.1  | (\$$COND281<0>301.1  | (\$$COND277<0>301.1  | (\$$COND276<0>301.1  | (\$$COND274<0>301.1  | (\$$COND271<0>301.1  | (\$$COND270<0>301.1  | (\$$COND267<0>301.1  | (\$$COND266<0>301.1  | (\$$COND265<0>301.1  | \$$COND264<0>301.1 )))))))))))))))))))))))))))))),
  \$$COND43<0>1.1  = ~\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \main_1/S6_1/$S6<0>451.1  = (~\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & \main_1/preS<36>0.1 ))))) | ((~\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 ))))) | ((\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & \main_1/preS<36>0.1 ))))) | ((\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 ))))) | (\$$COND452<0>451.1  | (\$$COND449<0>451.1  | (\$$COND447<0>451.1  | (\$$COND446<0>451.1  | (\$$COND445<0>451.1  | (\$$COND440<0>451.1  | (\$$COND439<0>451.1  | (\$$COND436<0>451.1  | (\$$COND435<0>451.1  | (\$$COND431<0>451.1  | (\$$COND428<0>451.1  | (\$$COND427<0>451.1  | (\$$COND425<0>451.1  | (\$$COND424<0>451.1  | (\$$COND419<0>451.1  | (\$$COND416<0>451.1  | (\$$COND415<0>451.1  | (\$$COND411<0>451.1  | (\$$COND409<0>451.1  | (\$$COND408<0>451.1  | (\$$COND406<0>451.1  | (\$$COND402<0>451.1  | (\$$COND401<0>451.1  | (\$$COND400<0>451.1  | (\$$COND398<0>451.1  | (\$$COND397<0>451.1  | (\$$COND394<0>451.1  | \$$COND391<0>451.1 )))))))))))))))))))))))))))))),
  \$$COND110<0>76.1  = ~\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \$$COND13<0>1.1  = ~\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \$$COND80<0>76.1  = \main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \$$COND264<0>301.1  = ~\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \$$COND112<0>76.1  = \main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \$$COND415<0>451.1  = \main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \$$COND436<0>451.1  = ~\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND136<0>151.1  = ~\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND82<0>76.1  = ~\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \$$COND307<0>301.1  = ~\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \$$COND157<0>151.1  = \main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND313<0>301.1  = \main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \$$COND81<0>76.1  = ~\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \$$COND113<0>76.1  = ~\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \$$COND84<0>76.1  = \main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \$$COND126<0>76.1  = ~\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \$$COND128<0>76.1  = \main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \$$COND467<0>526.1  = ~\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \$$COND127<0>76.1  = \main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \$$COND63<0>1.1  = \main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \[200]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<14>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<18>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<15>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<17>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<50>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<42>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<16>  & ~\$$COND521<0>601.1 )))))))),
  \$$COND53<0>1.1  = \main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \[201]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<13>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<17>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<14>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<16>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<50>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<15>  & ~\$$COND521<0>601.1 ))) | (~\reset<0>  & (~\encrypt<0>  & (\data_in<1>  & \$$COND521<0>601.1 )))))))),
  \[202]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<12>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<16>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<13>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<15>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<1>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<14>  & ~\$$COND521<0>601.1 ))) | (~\reset<0>  & (\encrypt<0>  & (\data_in<1>  & \$$COND521<0>601.1 )))))))),
  \main_1/preS<14>0.1  = (~\data<41>  & \C<11> ) | (\data<41>  & ~\C<11> ),
  \[203]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<11>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<15>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<12>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<14>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<9>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<1>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<13>  & ~\$$COND521<0>601.1 )))))))),
  \[204]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<10>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<14>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<11>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<13>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<9>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<17>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<12>  & ~\$$COND521<0>601.1 )))))))),
  \[205]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<9>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<13>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<10>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<12>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<25>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<17>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<11>  & ~\$$COND521<0>601.1 )))))))),
  \[206]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<8>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<12>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<9>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<11>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<33>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<25>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<10>  & ~\$$COND521<0>601.1 )))))))),
  \$$COND282<0>301.1  = \main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \$$COND122<0>76.1  = ~\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \main_1/preS<6>0.1  = (~\data<35>  & \C<2> ) | (\data<35>  & ~\C<2> ),
  \[207]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<7>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<11>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<8>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<10>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<41>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<33>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<9>  & ~\$$COND521<0>601.1 )))))))),
  \$$COND121<0>76.1  = ~\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \[208]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<6>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<10>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<7>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<9>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<49>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<41>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<8>  & ~\$$COND521<0>601.1 )))))))),
  \$$COND331<0>376.1  = ~\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \$$COND435<0>451.1  = ~\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND135<0>151.1  = ~\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND156<0>151.1  = \main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND177<0>151.1  = ~\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \$$COND124<0>76.1  = \main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \[209]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<5>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<9>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<6>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<8>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<49>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<7>  & ~\$$COND521<0>601.1 ))) | (~\reset<0>  & (~\encrypt<0>  & (\data_in<0>  & \$$COND521<0>601.1 )))))))),
  \$$COND123<0>76.1  = \main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \$$COND487<0>526.1  = ~\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \$$COND65<0>76.1  = ~\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \$$COND68<0>76.1  = \main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & \main_1/preS<10>0.1 )))),
  \$$COND8<0>1.1  = ~\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \[210]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<4>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<8>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<5>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<7>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<0>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<6>  & ~\$$COND521<0>601.1 ))) | (~\reset<0>  & (\encrypt<0>  & (\data_in<0>  & \$$COND521<0>601.1 )))))))),
  \[211]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<3>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<7>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<4>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<6>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<8>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<0>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<5>  & ~\$$COND521<0>601.1 )))))))),
  \$$COND69<0>76.1  = ~\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 )))),
  \[212]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<2>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<6>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<3>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<5>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<8>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<16>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<4>  & ~\$$COND521<0>601.1 )))))))),
  \[213]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<1>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<5>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<2>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<4>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<24>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<16>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<3>  & ~\$$COND521<0>601.1 )))))))),
  \[214]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<0>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<4>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<1>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<3>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<32>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<24>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<2>  & ~\$$COND521<0>601.1 )))))))),
  \main_1/preS<27>0.1  = (~\data<50>  & \D<8> ) | (\data<50>  & ~\D<8> ),
  \[215]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<27>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<3>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<0>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<2>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<40>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<32>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<1>  & ~\$$COND521<0>601.1 )))))))),
  \C_new<23>  = \[193] ,
  \[216]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<26>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<2>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\C<27>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\C<1>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<48>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<40>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\C<0>  & ~\$$COND521<0>601.1 )))))))),
  \C_new<24>  = \[192] ,
  \$$COND281<0>301.1  = \main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \[217]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<25>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<1>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<26>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<0>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<54>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<27>  & ~\$$COND521<0>601.1 ))) | (~\reset<0>  & (~\encrypt<0>  & (\data_in<3>  & \$$COND521<0>601.1 )))))))),
  \C_new<21>  = \[195] ,
  \main_1/S0_1/$S0<3>1.1  = (~\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & \main_1/preS<0>0.1 ))))) | ((~\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 ))))) | ((\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & \main_1/preS<0>0.1 ))))) | ((\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 ))))) | (\$$COND9<0>1.1  | (\$$COND6<0>1.1  | (\$$COND63<0>1.1  | (\$$COND60<0>1.1  | (\$$COND5<0>1.1  | (\$$COND59<0>1.1  | (\$$COND57<0>1.1  | (\$$COND53<0>1.1  | (\$$COND49<0>1.1  | (\$$COND48<0>1.1  | (\$$COND45<0>1.1  | (\$$COND42<0>1.1  | (\$$COND41<0>1.1  | (\$$COND40<0>1.1  | (\$$COND39<0>1.1  | (\$$COND36<0>1.1  | (\$$COND34<0>1.1  | (\$$COND2<0>1.1  | (\$$COND28<0>1.1  | (\$$COND27<0>1.1  | (\$$COND26<0>1.1  | (\$$COND24<0>1.1  | (\$$COND22<0>1.1  | (\$$COND20<0>1.1  | (\$$COND17<0>1.1  | (\$$COND13<0>1.1  | (\$$COND11<0>1.1  | \$$COND0<0>1.1 )))))))))))))))))))))))))))))),
  \[218]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<24>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<0>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<25>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<27>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<3>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<26>  & ~\$$COND521<0>601.1 ))) | (~\reset<0>  & (\encrypt<0>  & (\data_in<3>  & \$$COND521<0>601.1 )))))))),
  \C_new<22>  = \[194] ,
  \main_1/preS<10>0.1  = (~\data<39>  & \C<20> ) | (\data<39>  & ~\C<20> ),
  \$$COND220<0>226.1  = \main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND305<0>301.1  = ~\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \$$COND370<0>376.1  = ~\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND176<0>151.1  = ~\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \[219]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<23>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<27>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<24>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<26>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<3>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<11>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<25>  & ~\$$COND521<0>601.1 )))))))),
  \$$COND311<0>301.1  = \main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \C_new<20>  = \[196] ,
  \main_1/preS<39>0.1  = (~\data<58>  & \D<27> ) | (\data<58>  & ~\D<27> ),
  \$$COND469<0>526.1  = ~\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \$$COND488<0>526.1  = ~\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \data_new<4>  = \[180] ,
  \[220]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<22>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<26>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<23>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<25>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<19>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<11>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<24>  & ~\$$COND521<0>601.1 )))))))),
  \data_new<3>  = \[181] ,
  \[221]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<21>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<25>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<22>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<24>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<19>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<23>  & ~\$$COND521<0>601.1 ))) | (~\reset<0>  & (~\encrypt<0>  & (\data_in<4>  & \$$COND521<0>601.1 )))))))),
  \C_new<27>  = \[189] ,
  \data_new<2>  = \[182] ,
  \[222]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<20>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<24>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<21>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<23>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<4>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<22>  & ~\$$COND521<0>601.1 ))) | (~\reset<0>  & (\encrypt<0>  & (\data_in<4>  & \$$COND521<0>601.1 )))))))),
  \data_new<1>  = \[183] ,
  \[223]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<19>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<23>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<20>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<22>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<4>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<12>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<21>  & ~\$$COND521<0>601.1 )))))))),
  \C_new<25>  = \[191] ,
  \data_new<0>  = \[184] ,
  \[224]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<18>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<22>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<19>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<21>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<20>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<12>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<20>  & ~\$$COND521<0>601.1 )))))))),
  \C_new<26>  = \[190] ,
  \[225]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<17>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<21>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<18>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<20>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<28>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<20>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<19>  & ~\$$COND521<0>601.1 )))))))),
  \C_new<13>  = \[203] ,
  \[226]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<16>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<20>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<17>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<19>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<36>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<28>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<18>  & ~\$$COND521<0>601.1 )))))))),
  \C_new<14>  = \[202] ,
  \$$COND261<0>301.1  = ~\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \[227]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<15>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<19>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<16>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<18>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<44>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<36>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<17>  & ~\$$COND521<0>601.1 )))))))),
  \C_new<11>  = \[205] ,
  \[228]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<14>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<18>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<15>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<17>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<52>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<44>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<16>  & ~\$$COND521<0>601.1 )))))))),
  \C_new<12>  = \[204] ,
  \$$COND371<0>376.1  = ~\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND175<0>151.1  = ~\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \[229]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<13>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<17>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<14>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<16>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<52>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<15>  & ~\$$COND521<0>601.1 ))) | (~\reset<0>  & (~\encrypt<0>  & (\data_in<5>  & \$$COND521<0>601.1 )))))))),
  \C_new<10>  = \[206] ,
  \data_new<9>  = \[175] ,
  \main_1/S2_1/$S2<3>151.1  = (~\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & \main_1/preS<12>0.1 ))))) | ((~\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 ))))) | ((\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & \main_1/preS<12>0.1 ))))) | ((\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 ))))) | (\$$COND193<0>151.1  | (\$$COND190<0>151.1  | (\$$COND188<0>151.1  | (\$$COND187<0>151.1  | (\$$COND183<0>151.1  | (\$$COND180<0>151.1  | (\$$COND179<0>151.1  | (\$$COND176<0>151.1  | (\$$COND175<0>151.1  | (\$$COND173<0>151.1  | (\$$COND170<0>151.1  | (\$$COND167<0>151.1  | (\$$COND165<0>151.1  | (\$$COND162<0>151.1  | (\$$COND160<0>151.1  | (\$$COND159<0>151.1  | (\$$COND158<0>151.1  | (\$$COND157<0>151.1  | (\$$COND153<0>151.1  | (\$$COND149<0>151.1  | (\$$COND146<0>151.1  | (\$$COND142<0>151.1  | (\$$COND140<0>151.1  | (\$$COND139<0>151.1  | (\$$COND136<0>151.1  | (\$$COND133<0>151.1  | (\$$COND132<0>151.1  | \$$COND130<0>151.1 )))))))))))))))))))))))))))))),
  \main_1/preS<23>0.1  = (~\data<48>  & \C<1> ) | (\data<48>  & ~\C<1> ),
  \data_new<8>  = \[176] ,
  \data_new<7>  = \[177] ,
  \main_1/S5_1/$S5<2>376.1  = (~\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & \main_1/preS<30>0.1 ))))) | ((~\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 ))))) | ((\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & \main_1/preS<30>0.1 ))))) | ((\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 ))))) | (\$$COND388<0>376.1  | (\$$COND385<0>376.1  | (\$$COND384<0>376.1  | (\$$COND382<0>376.1  | (\$$COND379<0>376.1  | (\$$COND378<0>376.1  | (\$$COND376<0>376.1  | (\$$COND372<0>376.1  | (\$$COND370<0>376.1  | (\$$COND365<0>376.1  | (\$$COND363<0>376.1  | (\$$COND360<0>376.1  | (\$$COND359<0>376.1  | (\$$COND358<0>376.1  | (\$$COND352<0>376.1  | (\$$COND351<0>376.1  | (\$$COND349<0>376.1  | (\$$COND348<0>376.1  | (\$$COND346<0>376.1  | (\$$COND345<0>376.1  | (\$$COND342<0>376.1  | (\$$COND339<0>376.1  | (\$$COND338<0>376.1  | (\$$COND337<0>376.1  | (\$$COND334<0>376.1  | (\$$COND331<0>376.1  | (\$$COND328<0>376.1  | \$$COND325<0>376.1 )))))))))))))))))))))))))))))),
  \data_new<6>  = \[178] ,
  \data_new<5>  = \[179] ,
  \C_new<19>  = \[197] ,
  \[230]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<12>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<16>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<13>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<15>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<5>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<14>  & ~\$$COND521<0>601.1 ))) | (~\reset<0>  & (\encrypt<0>  & (\data_in<5>  & \$$COND521<0>601.1 )))))))),
  \[231]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<11>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<15>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<12>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<14>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<5>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<13>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<13>  & ~\$$COND521<0>601.1 )))))))),
  \C_new<17>  = \[199] ,
  \[232]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<10>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<14>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<11>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<13>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<21>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<13>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<12>  & ~\$$COND521<0>601.1 )))))))),
  \C_new<18>  = \[198] ,
  \main_1/preS<35>0.1  = (~\data<56>  & \D<19> ) | (\data<56>  & ~\D<19> ),
  \[233]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<9>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<13>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<10>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<12>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<29>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<21>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<11>  & ~\$$COND521<0>601.1 )))))))),
  \C_new<15>  = \[201] ,
  \[234]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<8>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<12>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<9>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<11>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<37>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<29>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<10>  & ~\$$COND521<0>601.1 )))))))),
  \C_new<16>  = \[200] ,
  \[235]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<7>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<11>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<8>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<10>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<45>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<37>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<9>  & ~\$$COND521<0>601.1 )))))))),
  \D_new<13>  = \[231] ,
  \$$COND42<0>1.1  = ~\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \[236]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<6>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<10>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<7>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<9>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<53>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<45>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<8>  & ~\$$COND521<0>601.1 )))))))),
  \D_new<14>  = \[230] ,
  \$$COND277<0>301.1  = \main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \[237]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<5>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<9>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<6>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<8>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<53>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<7>  & ~\$$COND521<0>601.1 ))) | (~\reset<0>  & (~\encrypt<0>  & (\data_in<6>  & \$$COND521<0>601.1 )))))))),
  \D_new<11>  = \[233] ,
  \$$COND22<0>1.1  = \main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \[238]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<4>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<8>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<5>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<7>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<6>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<6>  & ~\$$COND521<0>601.1 ))) | (~\reset<0>  & (\encrypt<0>  & (\data_in<6>  & \$$COND521<0>601.1 )))))))),
  \$$COND419<0>451.1  = \main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \$$COND334<0>376.1  = ~\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \D_new<12>  = \[232] ,
  \$$COND12<0>1.1  = ~\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \$$COND222<0>226.1  = \main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND372<0>376.1  = ~\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND351<0>376.1  = \main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \[239]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<3>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<7>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<4>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<6>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<6>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<14>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<5>  & ~\$$COND521<0>601.1 )))))))),
  \D_new<10>  = \[234] ,
  \data_new<63>  = \[121] ,
  \$$COND0<0>1.1  = ~\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \data_new<61>  = \[123] ,
  \data_new<62>  = \[122] ,
  \D_new<19>  = \[225] ,
  \data_new<60>  = \[124] ,
  \[240]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<2>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<6>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<3>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<5>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<22>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<14>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<4>  & ~\$$COND521<0>601.1 )))))))),
  \[241]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<1>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<5>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<2>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<4>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<30>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<22>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<3>  & ~\$$COND521<0>601.1 )))))))),
  \D_new<17>  = \[227] ,
  \[242]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<0>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<4>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<1>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<3>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<38>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<30>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<2>  & ~\$$COND521<0>601.1 )))))))),
  \D_new<18>  = \[226] ,
  \[243]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<27>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<3>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<0>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<2>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<46>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<38>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<1>  & ~\$$COND521<0>601.1 )))))))),
  \D_new<15>  = \[229] ,
  \$$COND62<0>1.1  = \main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \[244]  = (~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<26>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (~\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<2>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (~\encrypt_mode<0>  & (\D<27>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\generate_key_1/shift_by_one<0>605.1  & (~\generate_key_1/freeze<0>605.1  & (\encrypt_mode<0>  & (\D<1>  & ~\$$COND521<0>601.1 ))))) | ((~\reset<0>  & (\inreg<54>  & (~\encrypt<0>  & \$$COND521<0>601.1 ))) | ((~\reset<0>  & (\inreg<46>  & (\encrypt<0>  & \$$COND521<0>601.1 ))) | (~\reset<0>  & (\generate_key_1/freeze<0>605.1  & (\D<0>  & ~\$$COND521<0>601.1 )))))))),
  \D_new<16>  = \[228] ,
  \[245]  = (\count<3>  & (\count<2>  & (\count<1>  & (\count<0>  & \encrypt<0> )))) | ((~\count<3>  & \encrypt_mode<0> ) | ((~\count<2>  & \encrypt_mode<0> ) | ((~\count<1>  & \encrypt_mode<0> ) | (~\count<0>  & \encrypt_mode<0> )))),
  \D_new<23>  = \[221] ,
  \main_1/preS<1>0.1  = (~\data<32>  & \C<16> ) | (\data<32>  & ~\C<16> ),
  \D_new<24>  = \[220] ,
  \$$COND276<0>301.1  = \main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \D_new<21>  = \[223] ,
  \$$COND335<0>376.1  = ~\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \D_new<22>  = \[222] ,
  \$$COND439<0>451.1  = \main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND139<0>151.1  = ~\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \main_1/preS<31>0.1  = (~\data<52>  & \D<11> ) | (\data<52>  & ~\D<11> ),
  \$$COND352<0>376.1  = \main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \$$COND200<0>226.1  = ~\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND500<0>526.1  = ~\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \D_new<20>  = \[224] ,
  \data_new<53>  = \[131] ,
  \data_new<54>  = \[130] ,
  \data_new<51>  = \[133] ,
  \data_new<52>  = \[132] ,
  \main_1/S6_1/$S6<2>451.1  = (~\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 ))))) | ((~\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & \main_1/preS<36>0.1 ))))) | ((\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 ))))) | ((\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & \main_1/preS<36>0.1 ))))) | (\$$COND453<0>451.1  | (\$$COND450<0>451.1  | (\$$COND449<0>451.1  | (\$$COND447<0>451.1  | (\$$COND445<0>451.1  | (\$$COND440<0>451.1  | (\$$COND438<0>451.1  | (\$$COND435<0>451.1  | (\$$COND432<0>451.1  | (\$$COND431<0>451.1  | (\$$COND429<0>451.1  | (\$$COND428<0>451.1  | (\$$COND426<0>451.1  | (\$$COND425<0>451.1  | (\$$COND421<0>451.1  | (\$$COND419<0>451.1  | (\$$COND417<0>451.1  | (\$$COND416<0>451.1  | (\$$COND414<0>451.1  | (\$$COND409<0>451.1  | (\$$COND406<0>451.1  | (\$$COND404<0>451.1  | (\$$COND402<0>451.1  | (\$$COND401<0>451.1  | (\$$COND399<0>451.1  | (\$$COND397<0>451.1  | (\$$COND394<0>451.1  | \$$COND393<0>451.1 )))))))))))))))))))))))))))))),
  \data_new<50>  = \[134] ,
  \D_new<27>  = \[217] ,
  \D_new<25>  = \[219] ,
  \D_new<26>  = \[218] ,
  \data_new<59>  = \[125] ,
  \$$COND275<0>301.1  = ~\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \data_new<57>  = \[127] ,
  \$$COND298<0>301.1  = ~\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \data_new<58>  = \[126] ,
  \$$COND430<0>451.1  = ~\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND130<0>151.1  = ~\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \data_new<55>  = \[129] ,
  \$$COND224<0>226.1  = \main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND374<0>376.1  = \main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND159<0>151.1  = \main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND243<0>226.1  = \main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND201<0>226.1  = ~\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND501<0>526.1  = ~\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \data_new<56>  = \[128] ,
  \main_1/preS<44>0.1  = (~\data<61>  & \D<21> ) | (\data<61>  & ~\D<21> ),
  \main_1/S7_1/$S7<0>526.1  = (~\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/preS<42>0.1 ))))) | ((~\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 ))))) | ((\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 ))))) | ((\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/preS<42>0.1 ))))) | (\$$COND518<0>526.1  | (\$$COND516<0>526.1  | (\$$COND515<0>526.1  | (\$$COND513<0>526.1  | (\$$COND511<0>526.1  | (\$$COND510<0>526.1  | (\$$COND506<0>526.1  | (\$$COND501<0>526.1  | (\$$COND500<0>526.1  | (\$$COND499<0>526.1  | (\$$COND498<0>526.1  | (\$$COND491<0>526.1  | (\$$COND488<0>526.1  | (\$$COND487<0>526.1  | (\$$COND485<0>526.1  | (\$$COND482<0>526.1  | (\$$COND480<0>526.1  | (\$$COND477<0>526.1  | (\$$COND476<0>526.1  | (\$$COND473<0>526.1  | (\$$COND472<0>526.1  | (\$$COND470<0>526.1  | (\$$COND467<0>526.1  | (\$$COND465<0>526.1  | (\$$COND464<0>526.1  | (\$$COND461<0>526.1  | (\$$COND460<0>526.1  | \$$COND455<0>526.1 )))))))))))))))))))))))))))))),
  \main_1/S1_1/$S1<1>76.1  = (~\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & \main_1/preS<10>0.1 ))))) | ((\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 ))))) | ((\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & \main_1/preS<10>0.1 ))))) | ((\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 ))))) | (\$$COND99<0>76.1  | (\$$COND98<0>76.1  | (\$$COND95<0>76.1  | (\$$COND93<0>76.1  | (\$$COND92<0>76.1  | (\$$COND88<0>76.1  | (\$$COND85<0>76.1  | (\$$COND84<0>76.1  | (\$$COND81<0>76.1  | (\$$COND80<0>76.1  | (\$$COND74<0>76.1  | (\$$COND71<0>76.1  | (\$$COND70<0>76.1  | (\$$COND69<0>76.1  | (\$$COND68<0>76.1  | (\$$COND65<0>76.1  | (\$$COND127<0>76.1  | (\$$COND123<0>76.1  | (\$$COND122<0>76.1  | (\$$COND121<0>76.1  | (\$$COND118<0>76.1  | (\$$COND117<0>76.1  | (\$$COND115<0>76.1  | (\$$COND112<0>76.1  | (\$$COND110<0>76.1  | (\$$COND108<0>76.1  | (\$$COND101<0>76.1  | \$$COND100<0>76.1 )))))))))))))))))))))))))))))),
  \$$COND297<0>301.1  = ~\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \$$COND337<0>376.1  = ~\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \$$COND225<0>226.1  = \main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND300<0>301.1  = ~\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \$$COND450<0>451.1  = \main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND150<0>151.1  = \main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND244<0>226.1  = \main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND354<0>376.1  = \main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \$$COND179<0>151.1  = \main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \$$COND202<0>226.1  = ~\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \main_1/preS<17>0.1  = (~\data<44>  & \C<7> ) | (\data<44>  & ~\C<7> ),
  \main_1/S5_1/$S5<1>376.1  = (~\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & \main_1/preS<30>0.1 ))))) | ((~\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 ))))) | ((\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & \main_1/preS<30>0.1 ))))) | ((\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 ))))) | (\$$COND385<0>376.1  | (\$$COND384<0>376.1  | (\$$COND382<0>376.1  | (\$$COND381<0>376.1  | (\$$COND380<0>376.1  | (\$$COND379<0>376.1  | (\$$COND374<0>376.1  | (\$$COND372<0>376.1  | (\$$COND371<0>376.1  | (\$$COND368<0>376.1  | (\$$COND365<0>376.1  | (\$$COND364<0>376.1  | (\$$COND359<0>376.1  | (\$$COND358<0>376.1  | (\$$COND355<0>376.1  | (\$$COND354<0>376.1  | (\$$COND352<0>376.1  | (\$$COND349<0>376.1  | (\$$COND345<0>376.1  | (\$$COND342<0>376.1  | (\$$COND341<0>376.1  | (\$$COND340<0>376.1  | (\$$COND338<0>376.1  | (\$$COND337<0>376.1  | (\$$COND335<0>376.1  | (\$$COND331<0>376.1  | (\$$COND328<0>376.1  | \$$COND327<0>376.1 )))))))))))))))))))))))))))))),
  \main_1/preS<40>0.1  = (~\data<59>  & \D<5> ) | (\data<59>  & ~\D<5> ),
  \main_1/preS<9>0.1  = (~\data<38>  & \C<5> ) | (\data<38>  & ~\C<5> ),
  \$$COND296<0>301.1  = ~\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \main_1/S3_1/$S3<0>226.1  = (~\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 ))))) | ((~\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & \main_1/preS<18>0.1 ))))) | ((\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 ))))) | ((\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & \main_1/preS<18>0.1 ))))) | (\$$COND256<0>226.1  | (\$$COND254<0>226.1  | (\$$COND253<0>226.1  | (\$$COND251<0>226.1  | (\$$COND249<0>226.1  | (\$$COND244<0>226.1  | (\$$COND243<0>226.1  | (\$$COND239<0>226.1  | (\$$COND237<0>226.1  | (\$$COND235<0>226.1  | (\$$COND234<0>226.1  | (\$$COND233<0>226.1  | (\$$COND232<0>226.1  | (\$$COND229<0>226.1  | (\$$COND226<0>226.1  | (\$$COND220<0>226.1  | (\$$COND218<0>226.1  | (\$$COND216<0>226.1  | (\$$COND214<0>226.1  | (\$$COND213<0>226.1  | (\$$COND211<0>226.1  | (\$$COND210<0>226.1  | (\$$COND207<0>226.1  | (\$$COND206<0>226.1  | (\$$COND201<0>226.1  | (\$$COND198<0>226.1  | (\$$COND196<0>226.1  | \$$COND195<0>226.1 )))))))))))))))))))))))))))))),
  \$$COND338<0>376.1  = ~\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \main_1/S4_1/$S4<3>301.1  = (~\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 ))))) | ((~\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & \main_1/preS<24>0.1 ))))) | ((\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 ))))) | ((\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & \main_1/preS<24>0.1 ))))) | (\$$COND320<0>301.1  | (\$$COND319<0>301.1  | (\$$COND317<0>301.1  | (\$$COND315<0>301.1  | (\$$COND313<0>301.1  | (\$$COND310<0>301.1  | (\$$COND308<0>301.1  | (\$$COND307<0>301.1  | (\$$COND302<0>301.1  | (\$$COND301<0>301.1  | (\$$COND300<0>301.1  | (\$$COND297<0>301.1  | (\$$COND296<0>301.1  | (\$$COND295<0>301.1  | (\$$COND289<0>301.1  | (\$$COND287<0>301.1  | (\$$COND286<0>301.1  | (\$$COND282<0>301.1  | (\$$COND279<0>301.1  | (\$$COND277<0>301.1  | (\$$COND276<0>301.1  | (\$$COND275<0>301.1  | (\$$COND274<0>301.1  | (\$$COND272<0>301.1  | (\$$COND271<0>301.1  | (\$$COND266<0>301.1  | (\$$COND265<0>301.1  | \$$COND261<0>301.1 )))))))))))))))))))))))))))))),
  \$$COND226<0>226.1  = \main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND376<0>376.1  = \main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND355<0>376.1  = \main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \$$COND170<0>151.1  = ~\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \$$COND41<0>1.1  = ~\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \$$COND11<0>1.1  = ~\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \$$COND491<0>526.1  = ~\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \$$COND520<0>0.1  = \count<3>  & (\count<2>  & (\count<1>  & \count<0> )),
  \main_1/S0_1/$S0<0>1.1  = (~\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & \main_1/preS<0>0.1 ))))) | ((~\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 ))))) | ((\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & \main_1/preS<0>0.1 ))))) | ((\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 ))))) | (\$$COND8<0>1.1  | (\$$COND6<0>1.1  | (\$$COND63<0>1.1  | (\$$COND5<0>1.1  | (\$$COND58<0>1.1  | (\$$COND57<0>1.1  | (\$$COND56<0>1.1  | (\$$COND55<0>1.1  | (\$$COND53<0>1.1  | (\$$COND48<0>1.1  | (\$$COND46<0>1.1  | (\$$COND44<0>1.1  | (\$$COND43<0>1.1  | (\$$COND42<0>1.1  | (\$$COND40<0>1.1  | (\$$COND39<0>1.1  | (\$$COND36<0>1.1  | (\$$COND30<0>1.1  | (\$$COND2<0>1.1  | (\$$COND29<0>1.1  | (\$$COND28<0>1.1  | (\$$COND27<0>1.1  | (\$$COND22<0>1.1  | (\$$COND18<0>1.1  | (\$$COND17<0>1.1  | (\$$COND15<0>1.1  | (\$$COND13<0>1.1  | \$$COND12<0>1.1 )))))))))))))))))))))))))))))),
  \main_1/preS<13>0.1  = (~\data<40>  & \C<18> ) | (\data<40>  & ~\C<18> ),
  \$$COND295<0>301.1  = ~\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \$$COND414<0>451.1  = \main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \$$COND339<0>376.1  = ~\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \main_1/preS<5>0.1  = (~\data<36>  & \C<4> ) | (\data<36>  & ~\C<4> ),
  \$$COND227<0>226.1  = ~\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND377<0>376.1  = \main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND246<0>226.1  = \main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND190<0>151.1  = \main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \$$COND398<0>451.1  = ~\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \$$COND492<0>526.1  = ~\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \main_1/S6_1/$S6<1>451.1  = (~\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 ))))) | ((~\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & \main_1/preS<36>0.1 ))))) | ((\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 ))))) | ((\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & \main_1/preS<36>0.1 ))))) | (\$$COND452<0>451.1  | (\$$COND450<0>451.1  | (\$$COND449<0>451.1  | (\$$COND445<0>451.1  | (\$$COND444<0>451.1  | (\$$COND439<0>451.1  | (\$$COND438<0>451.1  | (\$$COND432<0>451.1  | (\$$COND431<0>451.1  | (\$$COND430<0>451.1  | (\$$COND429<0>451.1  | (\$$COND428<0>451.1  | (\$$COND427<0>451.1  | (\$$COND424<0>451.1  | (\$$COND421<0>451.1  | (\$$COND419<0>451.1  | (\$$COND415<0>451.1  | (\$$COND414<0>451.1  | (\$$COND413<0>451.1  | (\$$COND409<0>451.1  | (\$$COND408<0>451.1  | (\$$COND404<0>451.1  | (\$$COND403<0>451.1  | (\$$COND401<0>451.1  | (\$$COND398<0>451.1  | (\$$COND394<0>451.1  | (\$$COND393<0>451.1  | \$$COND391<0>451.1 )))))))))))))))))))))))))))))),
  \main_1/S1_1/$S1<0>76.1  = (~\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & \main_1/preS<10>0.1 ))))) | ((\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & \main_1/preS<10>0.1 ))))) | ((\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 ))))) | ((\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & \main_1/preS<10>0.1 ))))) | (\$$COND99<0>76.1  | (\$$COND96<0>76.1  | (\$$COND95<0>76.1  | (\$$COND94<0>76.1  | (\$$COND85<0>76.1  | (\$$COND84<0>76.1  | (\$$COND82<0>76.1  | (\$$COND81<0>76.1  | (\$$COND79<0>76.1  | (\$$COND76<0>76.1  | (\$$COND74<0>76.1  | (\$$COND73<0>76.1  | (\$$COND71<0>76.1  | (\$$COND70<0>76.1  | (\$$COND65<0>76.1  | (\$$COND128<0>76.1  | (\$$COND126<0>76.1  | (\$$COND123<0>76.1  | (\$$COND121<0>76.1  | (\$$COND118<0>76.1  | (\$$COND117<0>76.1  | (\$$COND113<0>76.1  | (\$$COND112<0>76.1  | (\$$COND110<0>76.1  | (\$$COND109<0>76.1  | (\$$COND105<0>76.1  | (\$$COND103<0>76.1  | \$$COND100<0>76.1 )))))))))))))))))))))))))))))),
  \$$COND279<0>301.1  = \main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \main_1/preS<26>0.1  = (~\data<49>  & \D<2> ) | (\data<49>  & ~\D<2> ),
  \$$COND413<0>451.1  = \main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \$$COND134<0>151.1  = ~\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND228<0>226.1  = ~\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND378<0>376.1  = \main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND247<0>226.1  = \main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND357<0>376.1  = ~\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND320<0>301.1  = \main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \$$COND505<0>526.1  = \main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \$$COND397<0>451.1  = ~\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \D_new<7>  = \[237] ,
  \C_new<6>  = \[210] ,
  \D_new<8>  = \[236] ,
  \C_new<5>  = \[211] ,
  \$$COND493<0>526.1  = ~\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \D_new<5>  = \[239] ,
  \C_new<8>  = \[208] ,
  \$$COND470<0>526.1  = ~\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \main_1/preS<38>0.1  = (~\data<57>  & \D<10> ) | (\data<57>  & ~\D<10> ),
  \D_new<6>  = \[238] ,
  \C_new<7>  = \[209] ,
  \C_new<9>  = \[207] ,
  \D_new<9>  = \[235] ,
  \D_new<0>  = \[244] ,
  \$$COND49<0>1.1  = \main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \C_new<0>  = \[216] ,
  \$$COND39<0>1.1  = ~\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \$$COND270<0>301.1  = ~\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \$$COND29<0>1.1  = \main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \D_new<3>  = \[241] ,
  \C_new<2>  = \[214] ,
  \D_new<4>  = \[240] ,
  \C_new<1>  = \[215] ,
  \$$COND133<0>151.1  = ~\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND229<0>226.1  = ~\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND304<0>301.1  = ~\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \$$COND379<0>376.1  = \main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND358<0>376.1  = ~\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \D_new<1>  = \[243] ,
  \C_new<4>  = \[212] ,
  \$$COND206<0>226.1  = ~\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND506<0>526.1  = \main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \D_new<2>  = \[242] ,
  \C_new<3>  = \[213] ,
  \main_1/preS<22>0.1  = (~\data<47>  & \C<12> ) | (\data<47>  & ~\C<12> ),
  \generate_key_1/freeze<0>605.1  = (~\encrypt_mode<0>  & (\encrypt<0>  & (\count<3>  & (\count<2>  & (\count<1>  & \count<0> ))))) | (\encrypt_mode<0>  & (~\encrypt<0>  & (\count<3>  & (\count<2>  & (\count<1>  & \count<0> ))))),
  \$$COND59<0>1.1  = \main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \main_1/preS<34>0.1  = (~\data<55>  & \D<4> ) | (\data<55>  & ~\D<4> ),
  \$$COND408<0>451.1  = \main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \$$COND411<0>451.1  = \main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \$$COND432<0>451.1  = ~\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND132<0>151.1  = ~\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND303<0>301.1  = ~\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \$$COND453<0>451.1  = \main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND153<0>151.1  = \main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND249<0>226.1  = \main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND359<0>376.1  = ~\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND174<0>151.1  = ~\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \$$COND207<0>226.1  = ~\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \main_1/S1_1/$S1<2>76.1  = (~\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & \main_1/preS<10>0.1 ))))) | ((\main_1/preS<9>0.1  & (~\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 ))))) | ((\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (~\main_1/preS<6>0.1  & (~\main_1/preS<11>0.1  & \main_1/preS<10>0.1 ))))) | ((\main_1/preS<9>0.1  & (\main_1/preS<8>0.1  & (~\main_1/preS<7>0.1  & (\main_1/preS<6>0.1  & (\main_1/preS<11>0.1  & ~\main_1/preS<10>0.1 ))))) | (\$$COND99<0>76.1  | (\$$COND98<0>76.1  | (\$$COND96<0>76.1  | (\$$COND93<0>76.1  | (\$$COND89<0>76.1  | (\$$COND88<0>76.1  | (\$$COND85<0>76.1  | (\$$COND84<0>76.1  | (\$$COND82<0>76.1  | (\$$COND79<0>76.1  | (\$$COND77<0>76.1  | (\$$COND76<0>76.1  | (\$$COND74<0>76.1  | (\$$COND69<0>76.1  | (\$$COND68<0>76.1  | (\$$COND65<0>76.1  | (\$$COND127<0>76.1  | (\$$COND126<0>76.1  | (\$$COND124<0>76.1  | (\$$COND123<0>76.1  | (\$$COND122<0>76.1  | (\$$COND118<0>76.1  | (\$$COND113<0>76.1  | (\$$COND112<0>76.1  | (\$$COND108<0>76.1  | (\$$COND107<0>76.1  | (\$$COND105<0>76.1  | \$$COND103<0>76.1 )))))))))))))))))))))))))))))),
  \main_1/S7_1/$S7<2>526.1  = (~\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/preS<42>0.1 ))))) | ((~\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 ))))) | ((\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/preS<42>0.1 ))))) | ((\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 ))))) | (\$$COND517<0>526.1  | (\$$COND516<0>526.1  | (\$$COND512<0>526.1  | (\$$COND511<0>526.1  | (\$$COND510<0>526.1  | (\$$COND506<0>526.1  | (\$$COND505<0>526.1  | (\$$COND501<0>526.1  | (\$$COND499<0>526.1  | (\$$COND498<0>526.1  | (\$$COND496<0>526.1  | (\$$COND493<0>526.1  | (\$$COND492<0>526.1  | (\$$COND487<0>526.1  | (\$$COND484<0>526.1  | (\$$COND481<0>526.1  | (\$$COND480<0>526.1  | (\$$COND479<0>526.1  | (\$$COND477<0>526.1  | (\$$COND473<0>526.1  | (\$$COND472<0>526.1  | (\$$COND470<0>526.1  | (\$$COND469<0>526.1  | (\$$COND467<0>526.1  | (\$$COND466<0>526.1  | (\$$COND460<0>526.1  | (\$$COND459<0>526.1  | \$$COND455<0>526.1 )))))))))))))))))))))))))))))),
  \$$COND40<0>1.1  = ~\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \$$COND472<0>526.1  = \main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \$$COND30<0>1.1  = \main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \$$COND20<0>1.1  = \main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \$$COND10<0>1.1  = ~\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \$$COND2<0>1.1  = ~\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \main_1/preS<47>0.1  = (~\data<32>  & \D<3> ) | (\data<32>  & ~\D<3> ),
  \main_1/preS<4>0.1  = (~\data<35>  & \C<0> ) | (\data<35>  & ~\C<0> ),
  \$$COND428<0>451.1  = ~\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND431<0>451.1  = ~\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND302<0>301.1  = ~\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \$$COND452<0>451.1  = \main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND152<0>151.1  = \main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND173<0>151.1  = ~\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \$$COND208<0>226.1  = ~\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND508<0>526.1  = \main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \main_1/preS<30>0.1  = (~\data<51>  & \D<1> ) | (\data<51>  & ~\D<1> ),
  \$$COND60<0>1.1  = \main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \$$COND496<0>526.1  = ~\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \$$COND473<0>526.1  = \main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \main_1/S3_1/$S3<2>226.1  = (~\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 ))))) | ((~\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & \main_1/preS<18>0.1 ))))) | ((\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 ))))) | ((\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & \main_1/preS<18>0.1 ))))) | (\$$COND258<0>226.1  | (\$$COND256<0>226.1  | (\$$COND255<0>226.1  | (\$$COND253<0>226.1  | (\$$COND249<0>226.1  | (\$$COND246<0>226.1  | (\$$COND244<0>226.1  | (\$$COND239<0>226.1  | (\$$COND238<0>226.1  | (\$$COND235<0>226.1  | (\$$COND234<0>226.1  | (\$$COND233<0>226.1  | (\$$COND231<0>226.1  | (\$$COND228<0>226.1  | (\$$COND225<0>226.1  | (\$$COND222<0>226.1  | (\$$COND220<0>226.1  | (\$$COND216<0>226.1  | (\$$COND215<0>226.1  | (\$$COND214<0>226.1  | (\$$COND211<0>226.1  | (\$$COND210<0>226.1  | (\$$COND208<0>226.1  | (\$$COND206<0>226.1  | (\$$COND200<0>226.1  | (\$$COND197<0>226.1  | (\$$COND196<0>226.1  | \$$COND195<0>226.1 )))))))))))))))))))))))))))))),
  \[10]  = (\inreg<46>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<38>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND406<0>451.1  = \main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \[11]  = (\inreg<45>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<37>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND427<0>451.1  = ~\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND301<0>301.1  = ~\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \$$COND193<0>151.1  = \main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \[12]  = (\inreg<44>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<36>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[13]  = (\inreg<43>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<35>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND9<0>1.1  = ~\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \[14]  = (\inreg<42>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<34>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[15]  = (\inreg<41>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<33>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND497<0>526.1  = ~\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \main_1/preS<43>0.1  = (~\data<60>  & \D<13> ) | (\data<60>  & ~\D<13> ),
  \$$COND455<0>526.1  = ~\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \[16]  = (\inreg<40>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<32>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \main_1/preS<0>0.1  = (~\data<63>  & \C<13> ) | (\data<63>  & ~\C<13> ),
  \[17]  = (\inreg<39>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<31>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[18]  = (\inreg<38>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<30>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[19]  = (\inreg<37>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<29>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND274<0>301.1  = ~\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \[20]  = (\inreg<36>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<28>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND48<0>1.1  = \main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \[21]  = (\inreg<35>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<27>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND426<0>451.1  = ~\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND447<0>451.1  = \main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND147<0>151.1  = \main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND168<0>151.1  = ~\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \[22]  = (\inreg<34>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<26>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND323<0>301.1  = \main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \$$COND28<0>1.1  = \main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \[23]  = (\inreg<33>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<25>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND18<0>1.1  = \main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \[24]  = (\inreg<32>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<24>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[25]  = (\inreg<31>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<23>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND498<0>526.1  = ~\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \[26]  = (\inreg<30>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<22>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND475<0>526.1  = \main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \[27]  = (\inreg<29>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<21>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[28]  = (\inreg<28>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<20>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \main_1/preS<16>0.1  = (~\data<43>  & \C<25> ) | (\data<43>  & ~\C<25> ),
  \[100]  = (\outreg<28>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<20>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<53>  & \$$COND520<0>0.1 )),
  \[29]  = (\inreg<27>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<19>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[101]  = (~\main_1/S4_1/$S4<2>301.1  & (\data<13>  & \$$COND520<0>0.1 )) | ((\main_1/S4_1/$S4<2>301.1  & (~\data<13>  & \$$COND520<0>0.1 )) | ((\outreg<27>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<19>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \[102]  = (\outreg<26>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<18>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<45>  & \$$COND520<0>0.1 )),
  \[103]  = (~\main_1/S2_1/$S2<0>151.1  & (\data<5>  & \$$COND520<0>0.1 )) | ((\main_1/S2_1/$S2<0>151.1  & (~\data<5>  & \$$COND520<0>0.1 )) | ((\outreg<25>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<17>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \[104]  = (\outreg<24>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<16>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<37>  & \$$COND520<0>0.1 )),
  \main_1/S2_1/$S2<0>151.1  = (~\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 ))))) | ((~\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & \main_1/preS<12>0.1 ))))) | ((\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & \main_1/preS<12>0.1 ))))) | ((\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 ))))) | (\$$COND191<0>151.1  | (\$$COND190<0>151.1  | (\$$COND189<0>151.1  | (\$$COND187<0>151.1  | (\$$COND185<0>151.1  | (\$$COND183<0>151.1  | (\$$COND180<0>151.1  | (\$$COND177<0>151.1  | (\$$COND174<0>151.1  | (\$$COND170<0>151.1  | (\$$COND168<0>151.1  | (\$$COND167<0>151.1  | (\$$COND165<0>151.1  | (\$$COND162<0>151.1  | (\$$COND160<0>151.1  | (\$$COND159<0>151.1  | (\$$COND156<0>151.1  | (\$$COND150<0>151.1  | (\$$COND149<0>151.1  | (\$$COND147<0>151.1  | (\$$COND146<0>151.1  | (\$$COND142<0>151.1  | (\$$COND141<0>151.1  | (\$$COND139<0>151.1  | (\$$COND137<0>151.1  | (\$$COND136<0>151.1  | (\$$COND135<0>151.1  | \$$COND132<0>151.1 )))))))))))))))))))))))))))))),
  \[105]  = (~\main_1/S0_1/$S0<0>1.1  & (\data<30>  & \$$COND520<0>0.1 )) | ((\main_1/S0_1/$S0<0>1.1  & (~\data<30>  & \$$COND520<0>0.1 )) | ((\outreg<23>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<15>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \[106]  = (\outreg<22>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<14>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<62>  & \$$COND520<0>0.1 )),
  \[107]  = (~\main_1/S0_1/$S0<1>1.1  & (\data<22>  & \$$COND520<0>0.1 )) | ((\main_1/S0_1/$S0<1>1.1  & (~\data<22>  & \$$COND520<0>0.1 )) | ((\outreg<21>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<13>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \$$COND58<0>1.1  = \main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \[30]  = (\inreg<26>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<18>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \main_1/S5_1/$S5<3>376.1  = (~\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & \main_1/preS<30>0.1 ))))) | ((~\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 ))))) | ((\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & \main_1/preS<30>0.1 ))))) | ((\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 ))))) | (\$$COND388<0>376.1  | (\$$COND382<0>376.1  | (\$$COND381<0>376.1  | (\$$COND380<0>376.1  | (\$$COND379<0>376.1  | (\$$COND377<0>376.1  | (\$$COND376<0>376.1  | (\$$COND371<0>376.1  | (\$$COND370<0>376.1  | (\$$COND368<0>376.1  | (\$$COND363<0>376.1  | (\$$COND359<0>376.1  | (\$$COND358<0>376.1  | (\$$COND357<0>376.1  | (\$$COND354<0>376.1  | (\$$COND352<0>376.1  | (\$$COND351<0>376.1  | (\$$COND347<0>376.1  | (\$$COND346<0>376.1  | (\$$COND342<0>376.1  | (\$$COND341<0>376.1  | (\$$COND340<0>376.1  | (\$$COND337<0>376.1  | (\$$COND334<0>376.1  | (\$$COND329<0>376.1  | (\$$COND328<0>376.1  | (\$$COND327<0>376.1  | \$$COND325<0>376.1 )))))))))))))))))))))))))))))),
  \[108]  = (\outreg<20>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<12>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<54>  & \$$COND520<0>0.1 )),
  \[31]  = (\inreg<25>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<17>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND425<0>451.1  = ~\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND340<0>376.1  = ~\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \$$COND446<0>451.1  = \main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND146<0>151.1  = \main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND167<0>151.1  = ~\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \$$COND188<0>151.1  = \main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \[109]  = (~\main_1/S7_1/$S7<1>526.1  & (\data<14>  & \$$COND520<0>0.1 )) | ((\main_1/S7_1/$S7<1>526.1  & (~\data<14>  & \$$COND520<0>0.1 )) | ((\outreg<19>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<11>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \$$COND191<0>151.1  = \main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \[32]  = (\inreg<24>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<16>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND322<0>301.1  = \main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \[33]  = (\inreg<23>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<15>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND399<0>451.1  = ~\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \[34]  = (\inreg<22>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<14>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[35]  = (\inreg<21>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<13>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND499<0>526.1  = ~\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \[36]  = (\inreg<20>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<12>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND476<0>526.1  = \main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \[37]  = (\inreg<19>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<11>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \main_1/S7_1/$S7<1>526.1  = (~\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 ))))) | ((~\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/preS<42>0.1 ))))) | ((\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/preS<42>0.1 ))))) | ((\main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 ))))) | (\$$COND518<0>526.1  | (\$$COND517<0>526.1  | (\$$COND515<0>526.1  | (\$$COND511<0>526.1  | (\$$COND508<0>526.1  | (\$$COND506<0>526.1  | (\$$COND505<0>526.1  | (\$$COND500<0>526.1  | (\$$COND499<0>526.1  | (\$$COND497<0>526.1  | (\$$COND496<0>526.1  | (\$$COND493<0>526.1  | (\$$COND488<0>526.1  | (\$$COND487<0>526.1  | (\$$COND484<0>526.1  | (\$$COND482<0>526.1  | (\$$COND481<0>526.1  | (\$$COND477<0>526.1  | (\$$COND476<0>526.1  | (\$$COND475<0>526.1  | (\$$COND472<0>526.1  | (\$$COND470<0>526.1  | (\$$COND466<0>526.1  | (\$$COND465<0>526.1  | (\$$COND463<0>526.1  | (\$$COND461<0>526.1  | (\$$COND460<0>526.1  | \$$COND459<0>526.1 )))))))))))))))))))))))))))))),
  \[38]  = (\inreg<18>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<10>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[110]  = (\outreg<18>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<10>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<46>  & \$$COND520<0>0.1 )),
  \[39]  = (\inreg<9>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<17>  & (~\count<0>  & ~\$$COND520<0>0.1 )),
  \[111]  = (~\main_1/S6_1/$S6<0>451.1  & (\data<6>  & \$$COND520<0>0.1 )) | ((\main_1/S6_1/$S6<0>451.1  & (~\data<6>  & \$$COND520<0>0.1 )) | ((\outreg<9>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<17>  & (\count<0>  & ~\$$COND520<0>0.1 )))),
  \main_1/preS<29>0.1  = (~\data<52>  & \D<26> ) | (\data<52>  & ~\D<26> ),
  \[112]  = (\outreg<8>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<16>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\data<38>  & \$$COND520<0>0.1 )),
  \[113]  = (~\main_1/S6_1/$S6<3>451.1  & (\data<31>  & \$$COND520<0>0.1 )) | ((\main_1/S6_1/$S6<3>451.1  & (~\data<31>  & \$$COND520<0>0.1 )) | ((\outreg<7>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<15>  & (\count<0>  & ~\$$COND520<0>0.1 )))),
  \[114]  = (\outreg<6>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<14>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\data<63>  & \$$COND520<0>0.1 )),
  \[115]  = (~\main_1/S2_1/$S2<3>151.1  & (\data<23>  & \$$COND520<0>0.1 )) | ((\main_1/S2_1/$S2<3>151.1  & (~\data<23>  & \$$COND520<0>0.1 )) | ((\outreg<5>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<13>  & (\count<0>  & ~\$$COND520<0>0.1 )))),
  \main_1/preS<12>0.1  = (~\data<39>  & \C<22> ) | (\data<39>  & ~\C<22> ),
  \[116]  = (\outreg<4>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<12>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\data<55>  & \$$COND520<0>0.1 )),
  \$$COND272<0>301.1  = ~\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \[117]  = (~\main_1/S2_1/$S2<2>151.1  & (\data<15>  & \$$COND520<0>0.1 )) | ((\main_1/S2_1/$S2<2>151.1  & (~\data<15>  & \$$COND520<0>0.1 )) | ((\outreg<3>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<11>  & (\count<0>  & ~\$$COND520<0>0.1 )))),
  \[40]  = (\inreg<8>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<16>  & (~\count<0>  & ~\$$COND520<0>0.1 )),
  \[118]  = (\outreg<2>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<10>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\data<47>  & \$$COND520<0>0.1 )),
  \[41]  = (\inreg<7>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<15>  & (~\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND251<0>226.1  = \main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND341<0>376.1  = \main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \$$COND445<0>451.1  = \main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND187<0>151.1  = \main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \[119]  = (~\main_1/S4_1/$S4<3>301.1  & (\data<7>  & \$$COND520<0>0.1 )) | ((\main_1/S4_1/$S4<3>301.1  & (~\data<7>  & \$$COND520<0>0.1 )) | ((\outreg<9>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<1>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \[42]  = (\inreg<6>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<14>  & (~\count<0>  & ~\$$COND520<0>0.1 )),
  \main_1/preS<8>0.1  = (~\data<37>  & \C<14> ) | (\data<37>  & ~\C<14> ),
  \[43]  = (\inreg<5>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<13>  & (~\count<0>  & ~\$$COND520<0>0.1 )),
  \[44]  = (\inreg<4>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<12>  & (~\count<0>  & ~\$$COND520<0>0.1 )),
  \[45]  = (\inreg<3>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<11>  & (~\count<0>  & ~\$$COND520<0>0.1 )),
  \[46]  = (\inreg<2>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<10>  & (~\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND477<0>526.1  = \main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \[47]  = (\inreg<9>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<1>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[48]  = (\inreg<8>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\inreg<0>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[120]  = (\outreg<8>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<0>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<39>  & \$$COND520<0>0.1 )),
  \[49]  = (\inreg<7>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data_in<7>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[121]  = (~\main_1/S6_1/$S6<3>451.1  & (\data<31>  & ~\$$COND520<0>0.1 )) | ((\main_1/S6_1/$S6<3>451.1  & (~\data<31>  & ~\$$COND520<0>0.1 )) | (\data_in<6>  & \$$COND520<0>0.1 )),
  \[122]  = (~\main_1/S0_1/$S0<0>1.1  & (\data<30>  & ~\$$COND520<0>0.1 )) | ((\main_1/S0_1/$S0<0>1.1  & (~\data<30>  & ~\$$COND520<0>0.1 )) | (\inreg<6>  & \$$COND520<0>0.1 )),
  \[123]  = (~\main_1/S2_1/$S2<1>151.1  & (\data<29>  & ~\$$COND520<0>0.1 )) | ((\main_1/S2_1/$S2<1>151.1  & (~\data<29>  & ~\$$COND520<0>0.1 )) | (\inreg<14>  & \$$COND520<0>0.1 )),
  \[124]  = (~\main_1/S5_1/$S5<2>376.1  & (\data<28>  & ~\$$COND520<0>0.1 )) | ((\main_1/S5_1/$S5<2>376.1  & (~\data<28>  & ~\$$COND520<0>0.1 )) | (\inreg<22>  & \$$COND520<0>0.1 )),
  \[125]  = (~\main_1/S1_1/$S1<2>76.1  & (\data<27>  & ~\$$COND520<0>0.1 )) | ((\main_1/S1_1/$S1<2>76.1  & (~\data<27>  & ~\$$COND520<0>0.1 )) | (\inreg<30>  & \$$COND520<0>0.1 )),
  \[126]  = (~\main_1/S7_1/$S7<2>526.1  & (\data<26>  & ~\$$COND520<0>0.1 )) | ((\main_1/S7_1/$S7<2>526.1  & (~\data<26>  & ~\$$COND520<0>0.1 )) | (\inreg<38>  & \$$COND520<0>0.1 )),
  \$$COND288<0>301.1  = \main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \main_1/S3_1/$S3<1>226.1  = (~\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 ))))) | ((~\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & \main_1/preS<18>0.1 ))))) | ((\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 ))))) | ((\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & \main_1/preS<18>0.1 ))))) | (\$$COND258<0>226.1  | (\$$COND256<0>226.1  | (\$$COND254<0>226.1  | (\$$COND247<0>226.1  | (\$$COND246<0>226.1  | (\$$COND244<0>226.1  | (\$$COND243<0>226.1  | (\$$COND238<0>226.1  | (\$$COND237<0>226.1  | (\$$COND235<0>226.1  | (\$$COND233<0>226.1  | (\$$COND232<0>226.1  | (\$$COND228<0>226.1  | (\$$COND227<0>226.1  | (\$$COND225<0>226.1  | (\$$COND224<0>226.1  | (\$$COND220<0>226.1  | (\$$COND218<0>226.1  | (\$$COND216<0>226.1  | (\$$COND215<0>226.1  | (\$$COND213<0>226.1  | (\$$COND210<0>226.1  | (\$$COND207<0>226.1  | (\$$COND202<0>226.1  | (\$$COND200<0>226.1  | (\$$COND198<0>226.1  | (\$$COND197<0>226.1  | \$$COND195<0>226.1 )))))))))))))))))))))))))))))),
  \$$COND271<0>301.1  = ~\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \[127]  = (~\main_1/S3_1/$S3<3>226.1  & (\data<25>  & ~\$$COND520<0>0.1 )) | ((\main_1/S3_1/$S3<3>226.1  & (~\data<25>  & ~\$$COND520<0>0.1 )) | (\inreg<46>  & \$$COND520<0>0.1 )),
  \[50]  = (\inreg<6>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data_in<6>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \main_1/preS<25>0.1  = (~\data<48>  & \D<23> ) | (\data<48>  & ~\D<23> ),
  \[128]  = (~\main_1/S4_1/$S4<1>301.1  & (\data<24>  & ~\$$COND520<0>0.1 )) | ((\main_1/S4_1/$S4<1>301.1  & (~\data<24>  & ~\$$COND520<0>0.1 )) | (\inreg<54>  & \$$COND520<0>0.1 )),
  \[51]  = (\inreg<5>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data_in<5>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND342<0>376.1  = \main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \$$COND210<0>226.1  = ~\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND510<0>526.1  = \main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \$$COND380<0>376.1  = \main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND165<0>151.1  = ~\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \main_1/S6_1/$S6<3>451.1  = (~\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 ))))) | ((~\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & \main_1/preS<36>0.1 ))))) | ((\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 ))))) | ((\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & \main_1/preS<36>0.1 ))))) | (\$$COND453<0>451.1  | (\$$COND450<0>451.1  | (\$$COND449<0>451.1  | (\$$COND446<0>451.1  | (\$$COND444<0>451.1  | (\$$COND440<0>451.1  | (\$$COND439<0>451.1  | (\$$COND436<0>451.1  | (\$$COND431<0>451.1  | (\$$COND430<0>451.1  | (\$$COND429<0>451.1  | (\$$COND426<0>451.1  | (\$$COND425<0>451.1  | (\$$COND424<0>451.1  | (\$$COND419<0>451.1  | (\$$COND417<0>451.1  | (\$$COND414<0>451.1  | (\$$COND413<0>451.1  | (\$$COND411<0>451.1  | (\$$COND408<0>451.1  | (\$$COND406<0>451.1  | (\$$COND403<0>451.1  | (\$$COND400<0>451.1  | (\$$COND399<0>451.1  | (\$$COND397<0>451.1  | (\$$COND394<0>451.1  | (\$$COND393<0>451.1  | \$$COND391<0>451.1 )))))))))))))))))))))))))))))),
  \[129]  = (~\main_1/S2_1/$S2<3>151.1  & (\data<23>  & ~\$$COND520<0>0.1 )) | ((\main_1/S2_1/$S2<3>151.1  & (~\data<23>  & ~\$$COND520<0>0.1 )) | (\data_in<4>  & \$$COND520<0>0.1 )),
  \[52]  = (\inreg<4>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data_in<4>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[53]  = (\inreg<3>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data_in<3>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \main_1/S0_1/$S0<1>1.1  = (~\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 ))))) | ((~\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & \main_1/preS<0>0.1 ))))) | ((\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 ))))) | ((\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & \main_1/preS<0>0.1 ))))) | (\$$COND9<0>1.1  | (\$$COND8<0>1.1  | (\$$COND6<0>1.1  | (\$$COND62<0>1.1  | (\$$COND60<0>1.1  | (\$$COND5<0>1.1  | (\$$COND59<0>1.1  | (\$$COND58<0>1.1  | (\$$COND57<0>1.1  | (\$$COND55<0>1.1  | (\$$COND48<0>1.1  | (\$$COND45<0>1.1  | (\$$COND44<0>1.1  | (\$$COND43<0>1.1  | (\$$COND40<0>1.1  | (\$$COND39<0>1.1  | (\$$COND37<0>1.1  | (\$$COND34<0>1.1  | (\$$COND30<0>1.1  | (\$$COND27<0>1.1  | (\$$COND25<0>1.1  | (\$$COND24<0>1.1  | (\$$COND20<0>1.1  | (\$$COND18<0>1.1  | (\$$COND17<0>1.1  | (\$$COND15<0>1.1  | (\$$COND10<0>1.1  | \$$COND0<0>1.1 )))))))))))))))))))))))))))))),
  \[54]  = (\inreg<2>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data_in<2>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \[55]  = (\inreg<1>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data_in<1>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \$$COND459<0>526.1  = ~\main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (~\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \[56]  = (\inreg<0>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data_in<0>  & (\count<0>  & ~\$$COND520<0>0.1 )),
  \inreg_new<50>  = \[6] ,
  \[57]  = (~\main_1/S4_1/$S4<1>301.1  & (\data<24>  & \$$COND520<0>0.1 )) | ((\main_1/S4_1/$S4<1>301.1  & (~\data<24>  & \$$COND520<0>0.1 )) | (\outreg<63>  & (~\count<0>  & ~\$$COND520<0>0.1 ))),
  \[58]  = (\outreg<62>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<56>  & \$$COND520<0>0.1 ),
  \main_1/preS<37>0.1  = (~\data<56>  & \D<20> ) | (\data<56>  & ~\D<20> ),
  \[130]  = (~\main_1/S0_1/$S0<1>1.1  & (\data<22>  & ~\$$COND520<0>0.1 )) | ((\main_1/S0_1/$S0<1>1.1  & (~\data<22>  & ~\$$COND520<0>0.1 )) | (\inreg<4>  & \$$COND520<0>0.1 )),
  \[59]  = (~\main_1/S0_1/$S0<2>1.1  & (\data<16>  & \$$COND520<0>0.1 )) | ((\main_1/S0_1/$S0<2>1.1  & (~\data<16>  & \$$COND520<0>0.1 )) | (\outreg<61>  & (~\count<0>  & ~\$$COND520<0>0.1 ))),
  \inreg_new<9>  = \[47] ,
  \[131]  = (~\main_1/S6_1/$S6<1>451.1  & (\data<21>  & ~\$$COND520<0>0.1 )) | ((\main_1/S6_1/$S6<1>451.1  & (~\data<21>  & ~\$$COND520<0>0.1 )) | (\inreg<12>  & \$$COND520<0>0.1 )),
  \inreg_new<54>  = \[2] ,
  \[132]  = (~\main_1/S7_1/$S7<0>526.1  & (\data<20>  & ~\$$COND520<0>0.1 )) | ((\main_1/S7_1/$S7<0>526.1  & (~\data<20>  & ~\$$COND520<0>0.1 )) | (\inreg<20>  & \$$COND520<0>0.1 )),
  \inreg_new<53>  = \[3] ,
  \[133]  = (~\main_1/S3_1/$S3<2>226.1  & (\data<19>  & ~\$$COND520<0>0.1 )) | ((\main_1/S3_1/$S3<2>226.1  & (~\data<19>  & ~\$$COND520<0>0.1 )) | (\inreg<28>  & \$$COND520<0>0.1 )),
  \inreg_new<52>  = \[4] ,
  \inreg_new<6>  = \[50] ,
  \[134]  = (~\main_1/S5_1/$S5<0>376.1  & (\data<18>  & ~\$$COND520<0>0.1 )) | ((\main_1/S5_1/$S5<0>376.1  & (~\data<18>  & ~\$$COND520<0>0.1 )) | (\inreg<36>  & \$$COND520<0>0.1 )),
  \inreg_new<51>  = \[5] ,
  \inreg_new<5>  = \[51] ,
  \[135]  = (~\main_1/S1_1/$S1<0>76.1  & (\data<17>  & ~\$$COND520<0>0.1 )) | ((\main_1/S1_1/$S1<0>76.1  & (~\data<17>  & ~\$$COND520<0>0.1 )) | (\inreg<44>  & \$$COND520<0>0.1 )),
  \inreg_new<8>  = \[48] ,
  \[136]  = (~\main_1/S0_1/$S0<2>1.1  & (\data<16>  & ~\$$COND520<0>0.1 )) | ((\main_1/S0_1/$S0<2>1.1  & (~\data<16>  & ~\$$COND520<0>0.1 )) | (\inreg<52>  & \$$COND520<0>0.1 )),
  \$$COND287<0>301.1  = \main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \inreg_new<7>  = \[49] ,
  \[137]  = (~\main_1/S2_1/$S2<2>151.1  & (\data<15>  & ~\$$COND520<0>0.1 )) | ((\main_1/S2_1/$S2<2>151.1  & (~\data<15>  & ~\$$COND520<0>0.1 )) | (\data_in<2>  & \$$COND520<0>0.1 )),
  \[60]  = (\outreg<60>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<48>  & \$$COND520<0>0.1 ),
  \inreg_new<2>  = \[54] ,
  \[138]  = (~\main_1/S7_1/$S7<1>526.1  & (\data<14>  & ~\$$COND520<0>0.1 )) | ((\main_1/S7_1/$S7<1>526.1  & (~\data<14>  & ~\$$COND520<0>0.1 )) | (\inreg<2>  & \$$COND520<0>0.1 )),
  \$$COND409<0>451.1  = \main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \[61]  = (~\main_1/S0_1/$S0<3>1.1  & (\data<8>  & \$$COND520<0>0.1 )) | ((\main_1/S0_1/$S0<3>1.1  & (~\data<8>  & \$$COND520<0>0.1 )) | (\outreg<59>  & (~\count<0>  & ~\$$COND520<0>0.1 ))),
  \$$COND253<0>226.1  = \main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND211<0>226.1  = \main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND511<0>526.1  = \main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \$$COND381<0>376.1  = \main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \inreg_new<55>  = \[1] ,
  \$$COND360<0>376.1  = ~\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND185<0>151.1  = \main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \inreg_new<1>  = \[55] ,
  \[139]  = (~\main_1/S4_1/$S4<2>301.1  & (\data<13>  & ~\$$COND520<0>0.1 )) | ((\main_1/S4_1/$S4<2>301.1  & (~\data<13>  & ~\$$COND520<0>0.1 )) | (\inreg<10>  & \$$COND520<0>0.1 )),
  \[62]  = (\outreg<58>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<40>  & \$$COND520<0>0.1 ),
  \$$COND317<0>301.1  = \main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \inreg_new<4>  = \[52] ,
  \[63]  = (~\main_1/S3_1/$S3<0>226.1  & (\data<0>  & \$$COND520<0>0.1 )) | ((\main_1/S3_1/$S3<0>226.1  & (~\data<0>  & \$$COND520<0>0.1 )) | (\outreg<57>  & (~\count<0>  & ~\$$COND520<0>0.1 ))),
  \inreg_new<3>  = \[53] ,
  \[64]  = (\outreg<56>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<32>  & \$$COND520<0>0.1 ),
  \[65]  = (~\main_1/S3_1/$S3<3>226.1  & (\data<25>  & \$$COND520<0>0.1 )) | ((\main_1/S3_1/$S3<3>226.1  & (~\data<25>  & \$$COND520<0>0.1 )) | ((\outreg<63>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<55>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \$$COND37<0>1.1  = ~\main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \[66]  = (\outreg<62>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<54>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<57>  & \$$COND520<0>0.1 )),
  \$$COND479<0>526.1  = \main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & ~\main_1/preS<42>0.1 )))),
  \$$COND27<0>1.1  = \main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \inreg_new<0>  = \[56] ,
  \[67]  = (~\main_1/S1_1/$S1<0>76.1  & (\data<17>  & \$$COND520<0>0.1 )) | ((\main_1/S1_1/$S1<0>76.1  & (~\data<17>  & \$$COND520<0>0.1 )) | ((\outreg<61>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<53>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \main_1/preS<21>0.1  = (~\data<46>  & \C<19> ) | (\data<46>  & ~\C<19> ),
  \$$COND17<0>1.1  = \main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \[68]  = (\outreg<60>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<52>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<49>  & \$$COND520<0>0.1 )),
  \[140]  = (~\main_1/S1_1/$S1<3>76.1  & (\data<12>  & ~\$$COND520<0>0.1 )) | ((\main_1/S1_1/$S1<3>76.1  & (~\data<12>  & ~\$$COND520<0>0.1 )) | (\inreg<18>  & \$$COND520<0>0.1 )),
  \[69]  = (~\main_1/S3_1/$S3<1>226.1  & (\data<9>  & \$$COND520<0>0.1 )) | ((\main_1/S3_1/$S3<1>226.1  & (~\data<9>  & \$$COND520<0>0.1 )) | ((\outreg<59>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<51>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \[141]  = (~\main_1/S6_1/$S6<2>451.1  & (\data<11>  & ~\$$COND520<0>0.1 )) | ((\main_1/S6_1/$S6<2>451.1  & (~\data<11>  & ~\$$COND520<0>0.1 )) | (\inreg<26>  & \$$COND520<0>0.1 )),
  \generate_key_1/shift_by_one<0>605.1  = (~\count<3>  & (~\count<2>  & (~\count<1>  & ~\count<0> ))) | ((~\count<3>  & (\count<2>  & (\count<1>  & \count<0> ))) | ((\count<3>  & (\count<2>  & (\count<1>  & ~\count<0> ))) | (\count<3>  & (\count<2>  & (\count<1>  & \count<0> ))))),
  \[142]  = (~\main_1/S5_1/$S5<1>376.1  & (\data<10>  & ~\$$COND520<0>0.1 )) | ((\main_1/S5_1/$S5<1>376.1  & (~\data<10>  & ~\$$COND520<0>0.1 )) | (\inreg<34>  & \$$COND520<0>0.1 )),
  \[143]  = (~\main_1/S3_1/$S3<1>226.1  & (\data<9>  & ~\$$COND520<0>0.1 )) | ((\main_1/S3_1/$S3<1>226.1  & (~\data<9>  & ~\$$COND520<0>0.1 )) | (\inreg<42>  & \$$COND520<0>0.1 )),
  \[144]  = (~\main_1/S0_1/$S0<3>1.1  & (\data<8>  & ~\$$COND520<0>0.1 )) | ((\main_1/S0_1/$S0<3>1.1  & (~\data<8>  & ~\$$COND520<0>0.1 )) | (\inreg<50>  & \$$COND520<0>0.1 )),
  \[145]  = (~\main_1/S4_1/$S4<3>301.1  & (\data<7>  & ~\$$COND520<0>0.1 )) | ((\main_1/S4_1/$S4<3>301.1  & (~\data<7>  & ~\$$COND520<0>0.1 )) | (\data_in<0>  & \$$COND520<0>0.1 )),
  \main_1/preS<33>0.1  = (~\data<54>  & \D<16> ) | (\data<54>  & ~\D<16> ),
  \[146]  = (~\main_1/S6_1/$S6<0>451.1  & (\data<6>  & ~\$$COND520<0>0.1 )) | ((\main_1/S6_1/$S6<0>451.1  & (~\data<6>  & ~\$$COND520<0>0.1 )) | (\inreg<0>  & \$$COND520<0>0.1 )),
  \$$COND286<0>301.1  = \main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \$$COND267<0>301.1  = ~\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \[147]  = (~\main_1/S2_1/$S2<0>151.1  & (\data<5>  & ~\$$COND520<0>0.1 )) | ((\main_1/S2_1/$S2<0>151.1  & (~\data<5>  & ~\$$COND520<0>0.1 )) | (\inreg<8>  & \$$COND520<0>0.1 )),
  \[70]  = (\outreg<58>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<50>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<41>  & \$$COND520<0>0.1 )),
  \[148]  = (~\main_1/S7_1/$S7<3>526.1  & (\data<4>  & ~\$$COND520<0>0.1 )) | ((\main_1/S7_1/$S7<3>526.1  & (~\data<4>  & ~\$$COND520<0>0.1 )) | (\inreg<16>  & \$$COND520<0>0.1 )),
  \$$COND400<0>451.1  = ~\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \[71]  = (~\main_1/S1_1/$S1<1>76.1  & (\data<1>  & \$$COND520<0>0.1 )) | ((\main_1/S1_1/$S1<1>76.1  & (~\data<1>  & \$$COND520<0>0.1 )) | ((\outreg<57>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<49>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \$$COND254<0>226.1  = \main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND429<0>451.1  = ~\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND512<0>526.1  = \main_1/preS<47>0.1  & (\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \$$COND382<0>376.1  = \main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \encrypt_mode_new<0>  = \[245] ,
  \$$COND231<0>226.1  = ~\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \[149]  = (~\main_1/S5_1/$S5<3>376.1  & (\data<3>  & ~\$$COND520<0>0.1 )) | ((\main_1/S5_1/$S5<3>376.1  & (~\data<3>  & ~\$$COND520<0>0.1 )) | (\inreg<24>  & \$$COND520<0>0.1 )),
  \[72]  = (\outreg<56>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<48>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<33>  & \$$COND520<0>0.1 )),
  \$$COND316<0>301.1  = \main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \[73]  = (~\main_1/S7_1/$S7<2>526.1  & (\data<26>  & \$$COND520<0>0.1 )) | ((\main_1/S7_1/$S7<2>526.1  & (~\data<26>  & \$$COND520<0>0.1 )) | ((\outreg<55>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<47>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \$$COND57<0>1.1  = \main_1/preS<5>0.1  & (\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \[74]  = (\outreg<54>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<46>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<58>  & \$$COND520<0>0.1 )),
  \[75]  = (~\main_1/S5_1/$S5<0>376.1  & (\data<18>  & \$$COND520<0>0.1 )) | ((\main_1/S5_1/$S5<0>376.1  & (~\data<18>  & \$$COND520<0>0.1 )) | ((\outreg<53>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<45>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \outreg_new<9>  = \[111] ,
  \[76]  = (\outreg<52>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<44>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<50>  & \$$COND520<0>0.1 )),
  \[77]  = (~\main_1/S5_1/$S5<1>376.1  & (\data<10>  & \$$COND520<0>0.1 )) | ((\main_1/S5_1/$S5<1>376.1  & (~\data<10>  & \$$COND520<0>0.1 )) | ((\outreg<51>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<43>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \outreg_new<51>  = \[69] ,
  \[78]  = (\outreg<50>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<42>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<42>  & \$$COND520<0>0.1 )),
  \outreg_new<52>  = \[68] ,
  \[150]  = (~\main_1/S4_1/$S4<0>301.1  & (\data<2>  & ~\$$COND520<0>0.1 )) | ((\main_1/S4_1/$S4<0>301.1  & (~\data<2>  & ~\$$COND520<0>0.1 )) | (\inreg<32>  & \$$COND520<0>0.1 )),
  \[79]  = (~\main_1/S4_1/$S4<0>301.1  & (\data<2>  & \$$COND520<0>0.1 )) | ((\main_1/S4_1/$S4<0>301.1  & (~\data<2>  & \$$COND520<0>0.1 )) | ((\outreg<49>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<41>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \outreg_new<53>  = \[67] ,
  \outreg_new<5>  = \[115] ,
  \[151]  = (~\main_1/S1_1/$S1<1>76.1  & (\data<1>  & ~\$$COND520<0>0.1 )) | ((\main_1/S1_1/$S1<1>76.1  & (~\data<1>  & ~\$$COND520<0>0.1 )) | (\inreg<40>  & \$$COND520<0>0.1 )),
  \outreg_new<54>  = \[66] ,
  \outreg_new<6>  = \[114] ,
  \[152]  = (~\main_1/S3_1/$S3<0>226.1  & (\data<0>  & ~\$$COND520<0>0.1 )) | ((\main_1/S3_1/$S3<0>226.1  & (~\data<0>  & ~\$$COND520<0>0.1 )) | (\inreg<48>  & \$$COND520<0>0.1 )),
  \outreg_new<7>  = \[113] ,
  \main_1/S4_1/$S4<0>301.1  = (~\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & \main_1/preS<24>0.1 ))))) | ((~\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (~\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 ))))) | ((\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & \main_1/preS<24>0.1 ))))) | ((\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 ))))) | (\$$COND323<0>301.1  | (\$$COND322<0>301.1  | (\$$COND319<0>301.1  | (\$$COND317<0>301.1  | (\$$COND315<0>301.1  | (\$$COND311<0>301.1  | (\$$COND308<0>301.1  | (\$$COND305<0>301.1  | (\$$COND303<0>301.1  | (\$$COND301<0>301.1  | (\$$COND300<0>301.1  | (\$$COND298<0>301.1  | (\$$COND297<0>301.1  | (\$$COND295<0>301.1  | (\$$COND289<0>301.1  | (\$$COND288<0>301.1  | (\$$COND286<0>301.1  | (\$$COND284<0>301.1  | (\$$COND282<0>301.1  | (\$$COND281<0>301.1  | (\$$COND277<0>301.1  | (\$$COND275<0>301.1  | (\$$COND272<0>301.1  | (\$$COND271<0>301.1  | (\$$COND270<0>301.1  | (\$$COND269<0>301.1  | (\$$COND266<0>301.1  | \$$COND264<0>301.1 )))))))))))))))))))))))))))))),
  \[153]  = (\data_in<7>  & \$$COND520<0>0.1 ) | (\data<63>  & ~\$$COND520<0>0.1 ),
  \outreg_new<8>  = \[112] ,
  \[154]  = (\inreg<7>  & \$$COND520<0>0.1 ) | (\data<62>  & ~\$$COND520<0>0.1 ),
  \outreg_new<1>  = \[119] ,
  \[155]  = (\inreg<15>  & \$$COND520<0>0.1 ) | (\data<61>  & ~\$$COND520<0>0.1 ),
  \outreg_new<50>  = \[70] ,
  \outreg_new<2>  = \[118] ,
  \[156]  = (\inreg<23>  & \$$COND520<0>0.1 ) | (\data<60>  & ~\$$COND520<0>0.1 ),
  \outreg_new<59>  = \[61] ,
  \$$COND266<0>301.1  = ~\main_1/preS<29>0.1  & (~\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \outreg_new<3>  = \[117] ,
  \$$COND291<0>301.1  = \main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \[157]  = (\inreg<31>  & \$$COND520<0>0.1 ) | (\data<59>  & ~\$$COND520<0>0.1 ),
  \[80]  = (\outreg<48>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<40>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<34>  & \$$COND520<0>0.1 )),
  \outreg_new<4>  = \[116] ,
  \main_1/preS<46>0.1  = (~\data<63>  & \D<0> ) | (\data<63>  & ~\D<0> ),
  \[158]  = (\inreg<39>  & \$$COND520<0>0.1 ) | (\data<58>  & ~\$$COND520<0>0.1 ),
  \[81]  = (~\main_1/S1_1/$S1<2>76.1  & (\data<27>  & \$$COND520<0>0.1 )) | ((\main_1/S1_1/$S1<2>76.1  & (~\data<27>  & \$$COND520<0>0.1 )) | ((\outreg<47>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<39>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \$$COND255<0>226.1  = \main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND345<0>376.1  = \main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \$$COND449<0>451.1  = \main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND149<0>151.1  = \main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND213<0>226.1  = \main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND513<0>526.1  = \main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (\main_1/preS<45>0.1  & (~\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \$$COND232<0>226.1  = ~\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \main_1/preS<3>0.1  = (~\data<34>  & \C<23> ) | (\data<34>  & ~\C<23> ),
  \[159]  = (\inreg<47>  & \$$COND520<0>0.1 ) | (\data<57>  & ~\$$COND520<0>0.1 ),
  \[82]  = (\outreg<46>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<38>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<59>  & \$$COND520<0>0.1 )),
  \$$COND315<0>301.1  = \main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & \main_1/preS<24>0.1 )))),
  \[83]  = (~\main_1/S3_1/$S3<2>226.1  & (\data<19>  & \$$COND520<0>0.1 )) | ((\main_1/S3_1/$S3<2>226.1  & (~\data<19>  & \$$COND520<0>0.1 )) | ((\outreg<45>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<37>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \outreg_new<55>  = \[65] ,
  \data_new<43>  = \[141] ,
  \$$COND394<0>451.1  = ~\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (~\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \[84]  = (\outreg<44>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<36>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<51>  & \$$COND520<0>0.1 )),
  \outreg_new<56>  = \[64] ,
  \data_new<44>  = \[140] ,
  \outreg_new<0>  = \[120] ,
  \[85]  = (~\main_1/S6_1/$S6<2>451.1  & (\data<11>  & \$$COND520<0>0.1 )) | ((\main_1/S6_1/$S6<2>451.1  & (~\data<11>  & \$$COND520<0>0.1 )) | ((\outreg<43>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<35>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \outreg_new<57>  = \[63] ,
  \data_new<41>  = \[143] ,
  \[86]  = (\outreg<42>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<34>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<43>  & \$$COND520<0>0.1 )),
  \outreg_new<58>  = \[62] ,
  \data_new<42>  = \[142] ,
  \inreg_new<20>  = \[36] ,
  \[87]  = (~\main_1/S5_1/$S5<3>376.1  & (\data<3>  & \$$COND520<0>0.1 )) | ((\main_1/S5_1/$S5<3>376.1  & (~\data<3>  & \$$COND520<0>0.1 )) | ((\outreg<41>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<33>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \outreg_new<61>  = \[59] ,
  \[88]  = (\outreg<40>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<32>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<35>  & \$$COND520<0>0.1 )),
  \outreg_new<62>  = \[58] ,
  \data_new<40>  = \[144] ,
  \[160]  = (\inreg<55>  & \$$COND520<0>0.1 ) | (\data<56>  & ~\$$COND520<0>0.1 ),
  \main_1/S2_1/$S2<2>151.1  = (~\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & \main_1/preS<12>0.1 ))))) | ((~\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 ))))) | ((\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & \main_1/preS<12>0.1 ))))) | ((\main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (~\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (~\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 ))))) | (\$$COND193<0>151.1  | (\$$COND191<0>151.1  | (\$$COND188<0>151.1  | (\$$COND187<0>151.1  | (\$$COND185<0>151.1  | (\$$COND182<0>151.1  | (\$$COND180<0>151.1  | (\$$COND177<0>151.1  | (\$$COND176<0>151.1  | (\$$COND174<0>151.1  | (\$$COND173<0>151.1  | (\$$COND167<0>151.1  | (\$$COND163<0>151.1  | (\$$COND162<0>151.1  | (\$$COND160<0>151.1  | (\$$COND158<0>151.1  | (\$$COND157<0>151.1  | (\$$COND156<0>151.1  | (\$$COND152<0>151.1  | (\$$COND147<0>151.1  | (\$$COND146<0>151.1  | (\$$COND141<0>151.1  | (\$$COND140<0>151.1  | (\$$COND139<0>151.1  | (\$$COND137<0>151.1  | (\$$COND136<0>151.1  | (\$$COND134<0>151.1  | \$$COND133<0>151.1 )))))))))))))))))))))))))))))),
  \[89]  = (~\main_1/S5_1/$S5<2>376.1  & (\data<28>  & \$$COND520<0>0.1 )) | ((\main_1/S5_1/$S5<2>376.1  & (~\data<28>  & \$$COND520<0>0.1 )) | ((\outreg<39>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<31>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \outreg_new<63>  = \[57] ,
  \[161]  = (\data_in<5>  & \$$COND520<0>0.1 ) | (\data<55>  & ~\$$COND520<0>0.1 ),
  \inreg_new<24>  = \[32] ,
  \[162]  = (\inreg<5>  & \$$COND520<0>0.1 ) | (\data<54>  & ~\$$COND520<0>0.1 ),
  \inreg_new<23>  = \[33] ,
  \[163]  = (\inreg<13>  & \$$COND520<0>0.1 ) | (\data<53>  & ~\$$COND520<0>0.1 ),
  \inreg_new<22>  = \[34] ,
  \[164]  = (\inreg<21>  & \$$COND520<0>0.1 ) | (\data<52>  & ~\$$COND520<0>0.1 ),
  \data_new<49>  = \[135] ,
  \inreg_new<21>  = \[35] ,
  \[165]  = (\inreg<29>  & \$$COND520<0>0.1 ) | (\data<51>  & ~\$$COND520<0>0.1 ),
  \outreg_new<60>  = \[60] ,
  \inreg_new<28>  = \[28] ,
  \[166]  = (\inreg<37>  & \$$COND520<0>0.1 ) | (\data<50>  & ~\$$COND520<0>0.1 ),
  \$$COND265<0>301.1  = ~\main_1/preS<29>0.1  & (\main_1/preS<28>0.1  & (~\main_1/preS<27>0.1  & (\main_1/preS<26>0.1  & (~\main_1/preS<25>0.1  & ~\main_1/preS<24>0.1 )))),
  \data_new<47>  = \[137] ,
  \inreg_new<27>  = \[29] ,
  \[167]  = (\inreg<45>  & \$$COND520<0>0.1 ) | (\data<49>  & ~\$$COND520<0>0.1 ),
  \[90]  = (\outreg<38>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<30>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<60>  & \$$COND520<0>0.1 )),
  \data_new<48>  = \[136] ,
  \inreg_new<26>  = \[30] ,
  \[168]  = (\inreg<53>  & \$$COND520<0>0.1 ) | (\data<48>  & ~\$$COND520<0>0.1 ),
  \[91]  = (~\main_1/S7_1/$S7<0>526.1  & (\data<20>  & \$$COND520<0>0.1 )) | ((\main_1/S7_1/$S7<0>526.1  & (~\data<20>  & \$$COND520<0>0.1 )) | ((\outreg<37>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<29>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \$$COND256<0>226.1  = \main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND346<0>376.1  = \main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \data_new<45>  = \[139] ,
  \$$COND140<0>151.1  = ~\main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \$$COND440<0>451.1  = \main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & \main_1/preS<36>0.1 )))),
  \$$COND325<0>376.1  = ~\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \$$COND214<0>226.1  = \main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (~\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND384<0>376.1  = \main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (~\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \inreg_new<25>  = \[31] ,
  \$$COND233<0>226.1  = ~\main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND363<0>376.1  = ~\main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \[169]  = (\data_in<3>  & \$$COND520<0>0.1 ) | (\data<47>  & ~\$$COND520<0>0.1 ),
  \[92]  = (\outreg<36>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<28>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<52>  & \$$COND520<0>0.1 )),
  \data_new<46>  = \[138] ,
  \[93]  = (~\main_1/S1_1/$S1<3>76.1  & (\data<12>  & \$$COND520<0>0.1 )) | ((\main_1/S1_1/$S1<3>76.1  & (~\data<12>  & \$$COND520<0>0.1 )) | ((\outreg<35>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<27>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \data_new<33>  = \[151] ,
  \$$COND393<0>451.1  = ~\main_1/preS<41>0.1  & (\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (~\main_1/preS<38>0.1  & (~\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 )))),
  \main_1/preS<19>0.1  = (~\data<44>  & \C<6> ) | (\data<44>  & ~\C<6> ),
  \[94]  = (\outreg<34>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<26>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<44>  & \$$COND520<0>0.1 )),
  \data_new<34>  = \[150] ,
  \[95]  = (~\main_1/S7_1/$S7<3>526.1  & (\data<4>  & \$$COND520<0>0.1 )) | ((\main_1/S7_1/$S7<3>526.1  & (~\data<4>  & \$$COND520<0>0.1 )) | ((\outreg<33>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<25>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \data_new<31>  = \[153] ,
  \inreg_new<29>  = \[27] ,
  \[96]  = (\outreg<32>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<24>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<36>  & \$$COND520<0>0.1 )),
  \data_new<32>  = \[152] ,
  \inreg_new<10>  = \[46] ,
  \[97]  = (~\main_1/S2_1/$S2<1>151.1  & (\data<29>  & \$$COND520<0>0.1 )) | ((\main_1/S2_1/$S2<1>151.1  & (~\data<29>  & \$$COND520<0>0.1 )) | ((\outreg<31>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<23>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \main_1/preS<42>0.1  = (~\data<59>  & \D<17> ) | (\data<59>  & ~\D<17> ),
  \[98]  = (\outreg<30>  & (\count<0>  & ~\$$COND520<0>0.1 )) | ((\outreg<22>  & (~\count<0>  & ~\$$COND520<0>0.1 )) | (\data<61>  & \$$COND520<0>0.1 )),
  \data_new<30>  = \[154] ,
  \[170]  = (\inreg<3>  & \$$COND520<0>0.1 ) | (\data<46>  & ~\$$COND520<0>0.1 ),
  \[99]  = (~\main_1/S6_1/$S6<1>451.1  & (\data<21>  & \$$COND520<0>0.1 )) | ((\main_1/S6_1/$S6<1>451.1  & (~\data<21>  & \$$COND520<0>0.1 )) | ((\outreg<29>  & (\count<0>  & ~\$$COND520<0>0.1 )) | (\outreg<21>  & (~\count<0>  & ~\$$COND520<0>0.1 )))),
  \[171]  = (\inreg<11>  & \$$COND520<0>0.1 ) | (\data<45>  & ~\$$COND520<0>0.1 ),
  \inreg_new<14>  = \[42] ,
  \[172]  = (\inreg<19>  & \$$COND520<0>0.1 ) | (\data<44>  & ~\$$COND520<0>0.1 ),
  \inreg_new<13>  = \[43] ,
  \[173]  = (\inreg<27>  & \$$COND520<0>0.1 ) | (\data<43>  & ~\$$COND520<0>0.1 ),
  \inreg_new<12>  = \[44] ,
  \[174]  = (\inreg<35>  & \$$COND520<0>0.1 ) | (\data<42>  & ~\$$COND520<0>0.1 ),
  \data_new<39>  = \[145] ,
  \inreg_new<11>  = \[45] ,
  \[175]  = (\inreg<43>  & \$$COND520<0>0.1 ) | (\data<41>  & ~\$$COND520<0>0.1 ),
  \inreg_new<18>  = \[38] ,
  \[176]  = (\inreg<51>  & \$$COND520<0>0.1 ) | (\data<40>  & ~\$$COND520<0>0.1 ),
  \data_new<37>  = \[147] ,
  \inreg_new<17>  = \[39] ,
  \[177]  = (\data_in<1>  & \$$COND520<0>0.1 ) | (\data<39>  & ~\$$COND520<0>0.1 ),
  \data_new<38>  = \[146] ,
  \inreg_new<16>  = \[40] ,
  \[178]  = (\inreg<1>  & \$$COND520<0>0.1 ) | (\data<38>  & ~\$$COND520<0>0.1 ),
  \$$COND347<0>376.1  = \main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & ~\main_1/preS<30>0.1 )))),
  \data_new<35>  = \[149] ,
  \$$COND215<0>226.1  = \main_1/preS<23>0.1  & (~\main_1/preS<22>0.1  & (~\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & ~\main_1/preS<18>0.1 )))),
  \$$COND515<0>526.1  = \main_1/preS<47>0.1  & (~\main_1/preS<46>0.1  & (~\main_1/preS<45>0.1  & (\main_1/preS<44>0.1  & (\main_1/preS<43>0.1  & \main_1/preS<42>0.1 )))),
  \$$COND385<0>376.1  = \main_1/preS<35>0.1  & (~\main_1/preS<34>0.1  & (~\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND160<0>151.1  = \main_1/preS<17>0.1  & (~\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & ~\main_1/preS<12>0.1 )))),
  \inreg_new<15>  = \[41] ,
  \$$COND234<0>226.1  = ~\main_1/preS<23>0.1  & (\main_1/preS<22>0.1  & (\main_1/preS<21>0.1  & (\main_1/preS<20>0.1  & (~\main_1/preS<19>0.1  & \main_1/preS<18>0.1 )))),
  \$$COND364<0>376.1  = ~\main_1/preS<35>0.1  & (\main_1/preS<34>0.1  & (\main_1/preS<33>0.1  & (\main_1/preS<32>0.1  & (~\main_1/preS<31>0.1  & \main_1/preS<30>0.1 )))),
  \$$COND189<0>151.1  = \main_1/preS<17>0.1  & (\main_1/preS<16>0.1  & (\main_1/preS<15>0.1  & (~\main_1/preS<14>0.1  & (\main_1/preS<13>0.1  & \main_1/preS<12>0.1 )))),
  \[179]  = (\inreg<9>  & \$$COND520<0>0.1 ) | (\data<37>  & ~\$$COND520<0>0.1 ),
  \data_new<36>  = \[148] ,
  \data_new<23>  = \[161] ,
  \data_new<24>  = \[160] ,
  \data_new<21>  = \[163] ,
  \inreg_new<19>  = \[37] ,
  \data_new<22>  = \[162] ,
  \inreg_new<40>  = \[16] ,
  \$$COND46<0>1.1  = ~\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \data_new<20>  = \[164] ,
  \$$COND36<0>1.1  = ~\main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (~\main_1/preS<3>0.1  & (\main_1/preS<2>0.1  & (~\main_1/preS<1>0.1  & \main_1/preS<0>0.1 )))),
  \[180]  = (\inreg<17>  & \$$COND520<0>0.1 ) | (\data<36>  & ~\$$COND520<0>0.1 ),
  \main_1/preS<15>0.1  = (~\data<42>  & \C<3> ) | (\data<42>  & ~\C<3> ),
  \$$COND26<0>1.1  = \main_1/preS<5>0.1  & (~\main_1/preS<4>0.1  & (\main_1/preS<3>0.1  & (~\main_1/preS<2>0.1  & (\main_1/preS<1>0.1  & ~\main_1/preS<0>0.1 )))),
  \[181]  = (\inreg<25>  & \$$COND520<0>0.1 ) | (\data<35>  & ~\$$COND520<0>0.1 ),
  \inreg_new<44>  = \[12] ,
  \[182]  = (\inreg<33>  & \$$COND520<0>0.1 ) | (\data<34>  & ~\$$COND520<0>0.1 ),
  \inreg_new<43>  = \[13] ,
  \[183]  = (\inreg<41>  & \$$COND520<0>0.1 ) | (\data<33>  & ~\$$COND520<0>0.1 ),
  \inreg_new<42>  = \[14] ,
  \[184]  = (\inreg<49>  & \$$COND520<0>0.1 ) | (\data<32>  & ~\$$COND520<0>0.1 ),
  \data_new<29>  = \[155] ,
  \inreg_new<41>  = \[15] ,
  \[185]  = (\count<1>  & (\count<0>  & (\count<2>  & (~\count<3>  & (~\reset<0>  & ~\$$COND521<0>601.1 ))))) | ((~\count<1>  & (\count<3>  & (~\reset<0>  & ~\$$COND521<0>601.1 ))) | ((~\count<0>  & (\count<3>  & (~\reset<0>  & ~\$$COND521<0>601.1 ))) | (~\count<2>  & (\count<3>  & (~\reset<0>  & ~\$$COND521<0>601.1 ))))),
  \inreg_new<48>  = \[8] ,
  \[186]  = (\count<1>  & (\count<0>  & (~\count<2>  & (~\reset<0>  & ~\$$COND521<0>601.1 )))) | ((~\count<1>  & (\count<2>  & (~\reset<0>  & ~\$$COND521<0>601.1 ))) | (~\count<0>  & (\count<2>  & (~\reset<0>  & ~\$$COND521<0>601.1 )))),
  \data_new<27>  = \[157] ,
  \inreg_new<47>  = \[9] ,
  \[187]  = (~\count<1>  & (\count<0>  & (~\reset<0>  & ~\$$COND521<0>601.1 ))) | (\count<1>  & (~\count<0>  & (~\reset<0>  & ~\$$COND521<0>601.1 ))),
  \data_new<28>  = \[156] ,
  \inreg_new<46>  = \[10] ,
  \[188]  = ~\count<0>  & (~\reset<0>  & ~\$$COND521<0>601.1 ),
  \$$COND404<0>451.1  = ~\main_1/preS<41>0.1  & (~\main_1/preS<40>0.1  & (\main_1/preS<39>0.1  & (\main_1/preS<38>0.1  & (\main_1/preS<37>0.1  & ~\main_1/preS<36>0.1 ))));
endmodule

