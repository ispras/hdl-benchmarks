// IWLS benchmark module "frg2" printed on Wed May 29 16:34:07 2002
module frg2(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5, s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, f8, g8, h8, i8, j8, k8, l8, m8, n8, o8, p8, q8, r8, s8, t8, u8, v8, w8, x8, y8, z8, a9, b9, c9, d9, e9, f9, g9, h9, i9, j9, k9, l9, m9, n9, o9, p9, q9, r9, s9, t9, u9, v9, w9);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  a1,
  a2,
  a3,
  a4,
  b0,
  b1,
  b2,
  b3,
  b4,
  c0,
  c1,
  c2,
  c3,
  c4,
  d0,
  d1,
  d2,
  d3,
  d4,
  e0,
  e1,
  e2,
  e3,
  e4,
  f0,
  f1,
  f2,
  f3,
  f4,
  g0,
  g1,
  g2,
  g3,
  g4,
  h0,
  h1,
  h2,
  h3,
  h4,
  i0,
  i1,
  i2,
  i3,
  i4,
  j0,
  j1,
  j2,
  j3,
  j4,
  k0,
  k1,
  k2,
  k3,
  k4,
  l0,
  l1,
  l2,
  l3,
  l4,
  m0,
  m1,
  m2,
  m3,
  m4,
  n0,
  n1,
  n2,
  n3,
  n4,
  o0,
  o1,
  o2,
  o3,
  p0,
  p1,
  p2,
  p3,
  q0,
  q1,
  q2,
  q3,
  r1,
  r2,
  r3,
  s0,
  s1,
  s2,
  s3,
  t0,
  t1,
  t2,
  t3,
  u0,
  u1,
  u2,
  u3,
  v0,
  v1,
  v2,
  v3,
  w0,
  w1,
  w2,
  w3,
  x0,
  x1,
  x2,
  x3,
  y0,
  y1,
  y2,
  y3,
  z0,
  z1,
  z2,
  z3;
output
  a5,
  a6,
  a7,
  a8,
  a9,
  b5,
  b6,
  b7,
  b8,
  b9,
  c5,
  c6,
  c7,
  c8,
  c9,
  d5,
  d6,
  d7,
  d8,
  d9,
  e5,
  e6,
  e7,
  e8,
  e9,
  f5,
  f6,
  f7,
  f8,
  f9,
  g5,
  g6,
  g7,
  g8,
  g9,
  h5,
  h6,
  h7,
  h8,
  h9,
  i5,
  i6,
  i7,
  i8,
  i9,
  j5,
  j6,
  j7,
  j8,
  j9,
  k5,
  k6,
  k7,
  k8,
  k9,
  l5,
  l6,
  l7,
  l8,
  l9,
  m5,
  m6,
  m7,
  m8,
  m9,
  n5,
  n6,
  n7,
  n8,
  n9,
  o4,
  o5,
  o6,
  o7,
  o8,
  o9,
  p4,
  p5,
  p6,
  p7,
  p8,
  p9,
  q4,
  q5,
  q6,
  q7,
  q8,
  q9,
  r4,
  r5,
  r6,
  r7,
  r8,
  r9,
  s4,
  s5,
  s6,
  s7,
  s8,
  s9,
  t4,
  t5,
  t6,
  t7,
  t8,
  t9,
  u4,
  u5,
  u6,
  u7,
  u8,
  u9,
  v4,
  v5,
  v6,
  v7,
  v8,
  v9,
  w4,
  w5,
  w6,
  w7,
  w8,
  w9,
  x4,
  x5,
  x6,
  x7,
  x8,
  y4,
  y5,
  y6,
  y7,
  y8,
  z4,
  z5,
  z6,
  z7,
  z8;
wire
  \[77] ,
  \[78] ,
  \[79] ,
  h16,
  h18,
  h19,
  h21,
  h22,
  h23,
  h24,
  h25,
  h27,
  h28,
  h30,
  h31,
  h33,
  h34,
  h35,
  \[80] ,
  \[81] ,
  \[82] ,
  \[83] ,
  \[84] ,
  x15,
  x16,
  x17,
  x18,
  \[85] ,
  x20,
  x21,
  x24,
  x25,
  x26,
  x28,
  x29,
  \[86] ,
  x30,
  x32,
  x33,
  x34,
  \[87] ,
  \[88] ,
  \[89] ,
  i17,
  i18,
  i20,
  i21,
  i23,
  i24,
  i25,
  i26,
  i28,
  i29,
  i31,
  i32,
  i33,
  i34,
  i35,
  \[90] ,
  \[91] ,
  \[92] ,
  \[93] ,
  \[94] ,
  y15,
  y17,
  y19,
  \[95] ,
  y21,
  y23,
  y24,
  y26,
  y27,
  y29,
  \[96] ,
  y31,
  y32,
  y33,
  \[97] ,
  \[100] ,
  \[98] ,
  \[101] ,
  \[99] ,
  \[102] ,
  j15,
  j16,
  j17,
  j19,
  j21,
  j23,
  \[103] ,
  j25,
  j26,
  j27,
  j28,
  j29,
  j30,
  j31,
  j32,
  j33,
  \[104] ,
  j35,
  \[105] ,
  \[106] ,
  \[107] ,
  \[108] ,
  \[0] ,
  \[109] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  z15,
  z18,
  z20,
  z21,
  z22,
  z23,
  z24,
  z25,
  z27,
  z29,
  z31,
  z33,
  \[7] ,
  \[110] ,
  \[8] ,
  \[111] ,
  \[9] ,
  \[112] ,
  k15,
  k18,
  k20,
  k21,
  \[113] ,
  k24,
  k25,
  k27,
  k28,
  k29,
  k30,
  k31,
  k32,
  k33,
  \[114] ,
  k34,
  k35,
  \[115] ,
  \[116] ,
  \[117] ,
  \[118] ,
  \[119] ,
  \[120] ,
  \[121] ,
  \[122] ,
  l15,
  l16,
  l17,
  l19,
  l20,
  l21,
  l22,
  \[123] ,
  l24,
  l25,
  l26,
  l28,
  l29,
  l30,
  l31,
  l32,
  l33,
  \[124] ,
  l34,
  l35,
  \[125] ,
  \[126] ,
  \[127] ,
  \[128] ,
  \[129] ,
  \[130] ,
  \[131] ,
  \[132] ,
  m15,
  m16,
  m18,
  m19,
  m22,
  \[133] ,
  m24,
  m25,
  m26,
  m27,
  m28,
  m29,
  m30,
  m31,
  m32,
  m33,
  \[134] ,
  m34,
  m35,
  \[135] ,
  \[136] ,
  \[137] ,
  \[138] ,
  n17,
  n18,
  n20,
  n22,
  n23,
  n25,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n33,
  n34,
  n35,
  o15,
  o17,
  o19,
  o22,
  o23,
  o24,
  o25,
  o26,
  o29,
  o30,
  o31,
  o32,
  o33,
  o34,
  o35,
  p16,
  p18,
  p20,
  p23,
  p24,
  p25,
  p26,
  p27,
  p28,
  p29,
  p30,
  p31,
  p32,
  p33,
  p34,
  p35,
  a17,
  a18,
  a20,
  a21,
  a22,
  a23,
  a24,
  a25,
  a26,
  a27,
  a29,
  a30,
  a32,
  a33,
  a34,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[14] ,
  q17,
  q19,
  \[15] ,
  q20,
  q21,
  q23,
  q24,
  q25,
  q27,
  q28,
  q29,
  \[16] ,
  q30,
  q31,
  q32,
  q33,
  q34,
  q35,
  \[17] ,
  \[18] ,
  \[19] ,
  b16,
  b17,
  b19,
  b20,
  b23,
  b25,
  b27,
  b28,
  b29,
  b30,
  b31,
  b32,
  b33,
  b34,
  b35,
  \[20] ,
  \[21] ,
  \[22] ,
  \[23] ,
  r16,
  r18,
  r19,
  \[25] ,
  r21,
  r23,
  r25,
  r26,
  r28,
  r29,
  \[26] ,
  r30,
  r31,
  r32,
  r33,
  r34,
  r35,
  \[27] ,
  \[28] ,
  \[29] ,
  c16,
  c18,
  c19,
  c21,
  c23,
  c24,
  c25,
  c26,
  c28,
  c30,
  c31,
  c32,
  c33,
  c34,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  s16,
  s17,
  s18,
  \[35] ,
  s20,
  s21,
  s22,
  s23,
  s24,
  s25,
  s26,
  s27,
  s28,
  \[36] ,
  s31,
  s32,
  s33,
  s34,
  \[37] ,
  \[38] ,
  \[39] ,
  d16,
  d17,
  d18,
  d20,
  d24,
  d25,
  d26,
  d27,
  d29,
  d30,
  d31,
  d32,
  d33,
  d34,
  d35,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  t15,
  t17,
  t19,
  \[45] ,
  t21,
  t22,
  t23,
  t24,
  t25,
  t27,
  t29,
  \[46] ,
  t30,
  t31,
  t32,
  t33,
  t34,
  \[47] ,
  \[48] ,
  \[49] ,
  e17,
  e19,
  e21,
  e22,
  e24,
  e25,
  e27,
  e28,
  e29,
  e30,
  e31,
  e32,
  e33,
  e34,
  e35,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  u16,
  u18,
  \[55] ,
  u20,
  u22,
  u23,
  u24,
  u26,
  u28,
  u29,
  \[56] ,
  u30,
  u31,
  u32,
  u33,
  \[57] ,
  \[58] ,
  \[59] ,
  f16,
  f18,
  f20,
  f21,
  f22,
  f25,
  f26,
  f28,
  f29,
  f30,
  f31,
  f32,
  f34,
  f35,
  \[60] ,
  \[61] ,
  \[62] ,
  \[63] ,
  \[64] ,
  v16,
  v17,
  v19,
  \[65] ,
  v20,
  v22,
  v26,
  v27,
  v28,
  v29,
  \[66] ,
  v30,
  v31,
  v33,
  v34,
  \[67] ,
  \[68] ,
  \[69] ,
  g15,
  g16,
  g17,
  g19,
  g20,
  g22,
  g23,
  g24,
  g25,
  g26,
  g27,
  g29,
  g30,
  g34,
  g35,
  \[70] ,
  \[71] ,
  \[72] ,
  \[73] ,
  \[74] ,
  w15,
  w16,
  w18,
  w19,
  \[75] ,
  w23,
  w24,
  w25,
  w27,
  w28,
  w29,
  \[76] ,
  w30,
  w31,
  w32,
  w33,
  w34;
assign
  \[77]  = (~f20 & (~u16 & ~s16)) | ((~f20 & (~u16 & ~d20)) | ((~f20 & (~u16 & a17)) | ((~f20 & (~n0 & ~s16)) | ((~f20 & (~n0 & ~d20)) | ((~f20 & (~n0 & a17)) | ((~f20 & (e2 & ~s16)) | ((~f20 & (e2 & ~d20)) | (~f20 & (e2 & a17))))))))),
  \[78]  = (~k20 & (~u16 & ~s16)) | ((~k20 & (~u16 & ~i20)) | ((~k20 & (~u16 & a17)) | ((~k20 & (~n0 & ~s16)) | ((~k20 & (~n0 & ~i20)) | ((~k20 & (~n0 & a17)) | ((~k20 & (f2 & ~s16)) | ((~k20 & (f2 & ~i20)) | (~k20 & (f2 & a17))))))))),
  \[79]  = (~p20 & (~u16 & ~s16)) | ((~p20 & (~u16 & ~n20)) | ((~p20 & (~u16 & a17)) | ((~p20 & (~n0 & ~s16)) | ((~p20 & (~n0 & ~n20)) | ((~p20 & (~n0 & a17)) | ((~p20 & (g2 & ~s16)) | ((~p20 & (g2 & ~n20)) | (~p20 & (g2 & a17))))))))),
  h16 = (t15 & (~e1 & ~n0)) | k1,
  h18 = (~w16 & (~t15 & ~u1)) | ~i18,
  h19 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & s))),
  h21 = (~k21 & (~j21 & ~a17)) | ((~i21 & (~s16 & ~m0)) | ~l21),
  h22 = (t15 & (~n0 & ~m0)) | ((l4 & ~a17) | n2),
  h23 = (p & (~l0 & k0)) | ((h & l0) | (h & ~k0)),
  h24 = w2 & l4,
  h25 = (k1 & l1) | (~i25 | ~k4),
  h27 = q0 | ~n3,
  h28 = ~o0 | q0,
  h30 = ~a4 & (~b4 & l4),
  h31 = ~m31 & (l25 & ~j25),
  h33 = (~l3 & ~d3) | ((~l3 & l0) | (~d3 & ~l0)),
  h34 = (~i4 & f1) | (i4 & ~f1),
  h35 = (~j35 & (a1 & z0)) | ((~j35 & (a1 & ~j1)) | ((~j35 & (z0 & ~k1)) | ((~j35 & (~k1 & ~j1)) | (~j35 & ~i35)))),
  \[80]  = (~u20 & (~u16 & ~s16)) | ((~u20 & (~u16 & ~s20)) | ((~u20 & (~u16 & a17)) | ((~u20 & (~n0 & ~s16)) | ((~u20 & (~n0 & ~s20)) | ((~u20 & (~n0 & a17)) | ((~u20 & (h2 & ~s16)) | ((~u20 & (h2 & ~s20)) | (~u20 & (h2 & a17))))))))),
  \[81]  = (~z20 & (~u16 & ~s16)) | ((~z20 & (~u16 & ~x20)) | ((~z20 & (~u16 & a17)) | ((~z20 & (~n0 & ~s16)) | ((~z20 & (~n0 & ~x20)) | ((~z20 & (~n0 & a17)) | ((~z20 & (i2 & ~s16)) | ((~z20 & (i2 & ~x20)) | (~z20 & (i2 & a17))))))))),
  \[82]  = (~e21 & (~u16 & ~s16)) | ((~e21 & (~u16 & ~c21)) | ((~e21 & (~u16 & a17)) | ((~e21 & (~n0 & ~s16)) | ((~e21 & (~n0 & ~c21)) | ((~e21 & (~n0 & a17)) | ((~e21 & (j2 & ~s16)) | ((~e21 & (j2 & ~c21)) | (~e21 & (j2 & a17))))))))),
  \[83]  = ~h21 & (o0 & ~q0),
  \[84]  = ~q21 & (o0 & ~q0),
  x15 = n0 | (e1 | ~t15),
  x16 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & j0))),
  x17 = (~w16 & (~t15 & ~s1)) | ~y17,
  x18 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & q))),
  \[85]  = ~x21 & (o0 & ~q0),
  x20 = ~j2 & l4,
  x21 = (~k21 & (~z21 & ~a17)) | ((~y21 & (~s16 & ~m0)) | ~a22),
  x24 = ~o0 | (q0 | ~t15),
  x25 = q0 | ~b3,
  x26 = j25 | (~l3 | ~k4),
  x28 = ~v0 | (j1 | ~k1),
  x29 = ~h30 | (~g30 | ~o0),
  \[86]  = ~e22 & (o0 & ~q0),
  x30 = l25 & (~j25 & k4),
  x32 = (~j25 & (~l1 & ~k1)) | (~j25 & ~j1),
  x33 = (~i3 & (~l0 & ~k0)) | ((~i3 & (l0 & k0)) | ~m0),
  x34 = (~l1 & (~k1 & ~j1)) | ((~l1 & (~k1 & z0)) | ((~l1 & (a1 & ~j1)) | ((~l1 & (a1 & z0)) | ((b1 & (~k1 & ~j1)) | ((b1 & (~k1 & z0)) | ((b1 & (a1 & ~j1)) | (b1 & (a1 & z0)))))))),
  \[87]  = ~l22 & (o0 & ~q0),
  \[88]  = ~s22 & (o0 & ~q0),
  \[89]  = ~z22 & (o0 & ~q0),
  i17 = (~w16 & (~t15 & ~p1)) | ~j17,
  i18 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & m0))),
  i20 = ~g2 & l4,
  i21 = (i & (~l0 & k0)) | ((a & l0) | (a & ~k0)),
  i23 = s2 | ~l4,
  i24 = (~t23 & (v2 & ~l4)) | (~s23 & (~r23 & l)),
  i25 = (~k25 & (~j25 & ~j1)) | (~k25 & (~j25 & ~l1)),
  i26 = j25 | (~g3 | ~k4),
  i28 = ~l25 | (j25 | ~k4),
  i29 = ~m29 & (~a17 & ~x3),
  i31 = ~j31 & (~g1 & ~q0),
  i32 = (n1 & i4) | ~j32,
  i33 = (~l3 & ~d3) | ((~l3 & ~l0) | (~d3 & l0)),
  i34 = ~g34 | (~y3 | ~z3),
  i35 = ~n35 | (~e4 | ~f4),
  \[90]  = ~g23 & (o0 & ~q0),
  \[91]  = ~n23 & (o0 & ~q0),
  \[92]  = ~y23 & (o0 & ~q0),
  \[93]  = ~c24 & (o0 & ~q0),
  \[94]  = ~g24 & (o0 & ~q0),
  y15 = ~z15 | (~o0 | q0),
  y17 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & e0))),
  y19 = ~e2 & l4,
  \[95]  = ~k24 & (o0 & ~q0),
  y21 = (k & (~l0 & k0)) | ((c & l0) | (c & ~k0)),
  y23 = (~a24 & (~z23 & ~a17)) | ((~a24 & (~z23 & ~t2)) | ((~a24 & (a17 & ~t2)) | (~a24 & ~p23))),
  y24 = q0 | ~z2,
  y26 = q0 | ~k3,
  y27 = j25 | (~u3 | ~k4),
  y29 = q0 | (a17 | x3),
  \[96]  = ~o24 & (o0 & ~q0),
  y31 = ~f32 | (~e32 | ~d32),
  y32 = ~j4 & (k4 & n4),
  y33 = (~j3 & (~l0 & ~k0)) | ((~j3 & (l0 & k0)) | ~m0),
  \[97]  = ~s24 & (o0 & ~q0),
  \[100]  = (~e25 & (~x25 & o0)) | (~c25 & (~w25 & ~a25)),
  \[98]  = (~z24 & (~y24 & o0)) | (~s23 & (~x24 & ~w24)),
  \[101]  = (~e25 & (~a26 & o0)) | (~c25 & (~z25 & ~a25)),
  \[99]  = (~e25 & (~d25 & o0)) | (~c25 & (~b25 & ~a25)),
  \[102]  = (~e25 & (~d26 & o0)) | (~c25 & (~c26 & ~a25)),
  j15 = ~o0 | (q0 | c1),
  j16 = ~m16 | (n0 | c1),
  j17 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & h0))),
  j19 = ~b2 & l4,
  j21 = l2 | ~l4,
  j23 = (t15 & (~n0 & ~m0)) | ((l4 & ~a17) | r2),
  \[103]  = (~e25 & (~g26 & o0)) | (~c25 & (~f26 & ~a25)),
  j25 = ~r35 & ~h4,
  j26 = q0 | ~f3,
  j27 = j25 | (~p3 | ~k4),
  j28 = (~s28 & ~q25) | ((~s28 & ~r28) | ((~s28 & ~s0) | ((h1 & ~q25) | ((h1 & ~r28) | (h1 & ~s0))))),
  j29 = (~k29 & (~q0 & n0)) | (~k29 & (~q0 & ~t15)),
  j30 = ~r30 | (~q30 | ~o0),
  j31 = (~l31 & (~k31 & l25)) | (~n0 & t15),
  j32 = o0 & (~q0 & ~a17),
  j33 = ~m0 & ~t3,
  \[104]  = (~e25 & (~j26 & o0)) | (~c25 & (~i26 & ~a25)),
  j35 = (~k35 & (l1 & ~b1)) | ((~k35 & ~i35) | (~k35 & ~n4)),
  \[105]  = (~e25 & (~m26 & o0)) | (~c25 & (~l26 & ~a25)),
  \[106]  = (~e25 & (~p26 & o0)) | (~c25 & (~o26 & ~a25)),
  \[107]  = (~e25 & (~s26 & o0)) | (~c25 & (~r26 & ~a25)),
  \[108]  = (~e25 & (~v26 & o0)) | (~c25 & (~u26 & ~a25)),
  \[0]  = ~g1,
  \[109]  = (~e25 & (~y26 & o0)) | (~c25 & (~x26 & ~a25)),
  \[1]  = (~j33 & (~i33 & ~h33)) | ((~j33 & (~i33 & k0)) | ((~j33 & (~h33 & ~k0)) | (~j33 & ~m0))),
  \[2]  = (~m33 & (~l33 & ~k33)) | ((~m33 & (~l33 & k0)) | ((~m33 & (~k33 & ~k0)) | (~m33 & ~m0))),
  \[3]  = (~p33 & (~o33 & ~n33)) | ((~p33 & (~o33 & k0)) | ((~p33 & (~n33 & ~k0)) | (~p33 & ~m0))),
  \[4]  = (~s33 & (~r33 & ~q33)) | ((~s33 & (~r33 & k0)) | ((~s33 & (~q33 & ~k0)) | (~s33 & ~m0))),
  z15 = (t15 & (~e1 & ~n0)) | i1,
  z18 = ~z1 & l4,
  z20 = (~w16 & (~t15 & ~i2)) | ~a21,
  z21 = n2 | ~l4,
  z22 = (~k21 & (~b23 & ~a17)) | ((~a23 & (~s16 & ~m0)) | ~c23),
  z23 = u2 & l4,
  z24 = (~s23 & (~s16 & ~m0)) | (~a17 & l4),
  z25 = j25 | (~d3 | ~k4),
  z27 = q0 | ~t3,
  z29 = ~n0 & t15,
  z31 = q0 | (g1 | ~h4),
  z33 = (~k3 & (~l0 & ~k0)) | ((~k3 & (l0 & k0)) | ~m0),
  \[7]  = (~t33 & (~l0 & ~k0)) | ((~t33 & (l0 & k0)) | (~t33 & m3)),
  \[110]  = (~e25 & (~b27 & o0)) | (~c25 & (~a27 & ~a25)),
  \[8]  = (~u33 & (~l0 & ~k0)) | ((~u33 & (l0 & k0)) | (~u33 & n3)),
  \[111]  = (~e25 & (~e27 & o0)) | (~c25 & (~d27 & ~a25)),
  \[9]  = (~v33 & (~l0 & ~k0)) | ((~v33 & (l0 & k0)) | (~v33 & o3)),
  \[112]  = (~e25 & (~h27 & o0)) | (~c25 & (~g27 & ~a25)),
  k15 = d1 | (e1 | ~t15),
  k18 = ~w1 & l4,
  k20 = (~w16 & (~t15 & ~f2)) | ~l20,
  k21 = ~m0 & (~n0 & t15),
  \[113]  = (~e25 & (~k27 & o0)) | (~c25 & (~j27 & ~a25)),
  k24 = (~m24 & (~l24 & ~a17)) | ((~m24 & (~l24 & ~w2)) | ((~m24 & (a17 & ~w2)) | (~m24 & ~p23))),
  k25 = (j1 & k1) | (~m25 | ~l25),
  k27 = q0 | ~o3,
  k28 = q0 | ~w3,
  k29 = ~l29 & (~z3 & l4),
  k30 = q0 | ~c4,
  k31 = j25 | d4,
  k32 = ~y32 | (~o0 | q0),
  k33 = (~k3 & ~c3) | ((~k3 & l0) | (~c3 & ~l0)),
  \[114]  = (~e25 & (~n27 & o0)) | (~c25 & (~m27 & ~a25)),
  k34 = h1 & (m1 & ~k4),
  k35 = ~l35 & (~g4 & ~h4),
  \[115]  = (~e25 & (~q27 & o0)) | (~c25 & (~p27 & ~a25)),
  \[116]  = (~e25 & (~t27 & o0)) | (~c25 & (~s27 & ~a25)),
  \[117]  = (~e25 & (~w27 & o0)) | (~c25 & (~v27 & ~a25)),
  \[118]  = (~e25 & (~z27 & o0)) | (~c25 & (~y27 & ~a25)),
  \[119]  = (~e25 & (~c28 & o0)) | (~c25 & (~b28 & ~a25)),
  \[120]  = (~e25 & (~f28 & o0)) | (~c25 & (~e28 & ~a25)),
  \[121]  = (~l28 & (~k28 & o0)) | (~j28 & (~i28 & ~h28)),
  \[122]  = (~a29 & (~a17 & l4)) | (~a29 & x3),
  l15 = q0 | (g1 | ~h1),
  l16 = (t15 & (~e1 & ~n0)) | (~o0 | q0),
  l17 = ~r1 & l4,
  l19 = (~w16 & (~t15 & ~a2)) | ~m19,
  l20 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & y))),
  l21 = (t15 & (~n0 & ~m0)) | ((l4 & ~a17) | k2),
  l22 = (~k21 & (~n22 & ~a17)) | ((~m22 & (~s16 & ~m0)) | ~o22),
  \[123]  = (~d29 & y3) | (~e29 | ~o0),
  l24 = x2 & l4,
  l25 = (~y0 & i1) | ((~x0 & h1) | ~x34),
  l26 = j25 | (~h3 | ~k4),
  l28 = (~m28 & (~g25 & ~f25)) | ((~m28 & (~g25 & ~h1)) | ((~m28 & (~i1 & ~f25)) | (~m28 & (~i1 & ~h1)))),
  l29 = a17 | (x3 | ~y3),
  l30 = (~p30 & (~o30 & ~a17)) | (~n0 & t15),
  l31 = ~e4 | (f4 | ~k4),
  l32 = ~l25 | (j25 | g1),
  l33 = (~k3 & ~c3) | ((~k3 & ~l0) | (~c3 & l0)),
  \[124]  = (~i29 & z3) | (~j29 | ~o0),
  l34 = i1 & (m1 & ~k4),
  l35 = ~m35 | (g1 | ~d4),
  \[125]  = ~n29 & (o0 & ~q0),
  \[126]  = (~b30 & (~a30 & o0)) | ((~z29 & (~y29 & ~x29)) | ~c30),
  \[127]  = (~l30 & (~k30 & o0)) | ((~z29 & (~y29 & ~j30)) | ~m30),
  \[128]  = (~v30 & (o0 & ~n0)) | (~u30 & (~t30 & o0)),
  \[129]  = (~b31 & e4) | (~c31 | ~o0),
  \[130]  = (~h31 & f4) | (~i31 | ~o0),
  \[131]  = (~q31 & (~p31 & o0)) | ((~z29 & (~o31 & ~n31)) | ~r31),
  \[132]  = (~a32 & (~z31 & o0)) | ((~z29 & (~a25 & ~y31)) | ~c30),
  m15 = ~o15 & (~n0 & t15),
  m16 = ~d1 & t15,
  m18 = (~w16 & (~t15 & ~v1)) | ~n18,
  m19 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & t))),
  m22 = (m & (~l0 & k0)) | ((e & l0) | (e & ~k0)),
  \[133]  = (~i32 & (l4 & n1)) | (~i32 & (l4 & i4)),
  m24 = (~t23 & (w2 & ~l4)) | (~s23 & (~r23 & m)),
  m25 = ~n25 | (k1 | l1),
  m26 = q0 | ~g3,
  m27 = j25 | (~q3 | ~k4),
  m28 = ~n28 | (j25 | ~k4),
  m29 = ~y3 | ~l4,
  m30 = ~n30 | (q0 | ~t15),
  m31 = d4 | (~e4 | ~k4),
  m32 = q0 | (g1 | ~j4),
  m33 = ~m0 & ~s3,
  \[134]  = (~n32 & (~m32 & o0)) | (~j28 & (~l32 & ~k32)),
  m34 = j1 & (m1 & ~k4),
  m35 = e4 & f4,
  \[135]  = ~a33 & (~b4 & ~c4),
  \[136]  = ~c33 & m1,
  \[137]  = (~e33 & ~d33) | (~e33 & ~g15),
  \[138]  = ~a25 & k4,
  n17 = (~w16 & (~t15 & ~q1)) | ~o17,
  n18 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & k0))),
  n20 = ~h2 & l4,
  n22 = p2 | ~l4,
  n23 = (~q23 & (~o23 & ~a17)) | ((~q23 & (~o23 & ~s2)) | ((~q23 & (a17 & ~s2)) | (~q23 & ~p23))),
  n25 = ~h1 & (~i1 & ~j1),
  n27 = q0 | ~p3,
  n28 = (~p28 & (l25 & ~k1)) | (~p28 & (l25 & ~l1)),
  n29 = (~r29 & (~q29 & ~s16)) | ((~r29 & (~q29 & ~p29)) | ((~r29 & (~q29 & ~o29)) | ((~r29 & (~n0 & ~s16)) | ((~r29 & (~n0 & ~p29)) | ((~r29 & (~n0 & ~o29)) | ((~r29 & (~a4 & ~s16)) | ((~r29 & (~a4 & ~p29)) | (~r29 & (~a4 & ~o29))))))))),
  a5 = \[12] ,
  n30 = ~m0 & (~n0 & o0),
  a6 = \[38] ,
  n31 = ~w31 | (~v31 | ~o0),
  a7 = \[64] ,
  n32 = (~r32 & (~q32 & ~p32)) | ((~r32 & (~q32 & ~o32)) | ((~r32 & (~q32 & h1)) | ((~r32 & (~p32 & ~h1)) | (~r32 & (~o32 & ~h1))))),
  a8 = \[90] ,
  n33 = (~j3 & ~b3) | ((~j3 & l0) | (~b3 & ~l0)),
  a9 = \[116] ,
  n34 = k1 & (m1 & ~k4),
  n35 = ~g4 & ~h4,
  b5 = \[13] ,
  b6 = \[39] ,
  b7 = \[65] ,
  b8 = \[91] ,
  b9 = \[117] ,
  c5 = \[14] ,
  c6 = \[40] ,
  c7 = \[66] ,
  c8 = \[92] ,
  c9 = \[118] ,
  d5 = \[15] ,
  d6 = \[41] ,
  d7 = \[67] ,
  d8 = \[93] ,
  d9 = \[119] ,
  e5 = \[16] ,
  e6 = \[42] ,
  e7 = \[68] ,
  e8 = \[94] ,
  e9 = \[120] ,
  f5 = \[17] ,
  f6 = \[43] ,
  f7 = \[69] ,
  f8 = \[95] ,
  f9 = \[121] ,
  g5 = \[18] ,
  g6 = \[44] ,
  g7 = \[70] ,
  g8 = \[96] ,
  g9 = \[122] ,
  h5 = \[19] ,
  h6 = \[45] ,
  h7 = \[71] ,
  h8 = \[97] ,
  h9 = \[123] ,
  i5 = \[20] ,
  i6 = \[46] ,
  i7 = \[72] ,
  i8 = \[98] ,
  i9 = \[124] ,
  j5 = \[21] ,
  j6 = \[47] ,
  j7 = \[73] ,
  j8 = \[99] ,
  j9 = \[125] ,
  k5 = \[22] ,
  k6 = \[48] ,
  k7 = \[74] ,
  k8 = \[100] ,
  k9 = \[126] ,
  l5 = \[23] ,
  l6 = \[49] ,
  l7 = \[75] ,
  l8 = \[101] ,
  l9 = \[127] ,
  m5 = m4,
  m6 = k4,
  m7 = \[76] ,
  m8 = \[102] ,
  m9 = \[128] ,
  n5 = \[25] ,
  n6 = \[51] ,
  n7 = \[77] ,
  n8 = \[103] ,
  n9 = \[129] ,
  o4 = \[0] ,
  o5 = \[26] ,
  o6 = \[52] ,
  o7 = \[78] ,
  o8 = \[104] ,
  o9 = \[130] ,
  o15 = (c1 & e1) | (e1 & d1),
  o17 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & g0))),
  o19 = ~c2 & l4,
  p4 = \[1] ,
  p5 = \[27] ,
  p6 = \[53] ,
  p7 = \[79] ,
  o22 = (t15 & (~n0 & ~m0)) | ((l4 & ~a17) | o2),
  p8 = \[105] ,
  o23 = t2 & l4,
  p9 = \[131] ,
  o24 = (~q24 & (~p24 & ~a17)) | ((~q24 & (~p24 & ~x2)) | ((~q24 & (a17 & ~x2)) | (~q24 & ~p23))),
  o25 = ~k1 & ~l1,
  o26 = j25 | (~i3 | ~k4),
  o29 = ~a17 & (~x3 & y3),
  q4 = \[2] ,
  q5 = \[28] ,
  o30 = x3 | (~y3 | ~z3),
  q6 = \[54] ,
  o31 = q0 | (~l25 | j25),
  q7 = \[80] ,
  o32 = ~i1 & ~j1,
  q8 = \[106] ,
  o33 = (~j3 & ~b3) | ((~j3 & ~l0) | (~b3 & l0)),
  q9 = \[132] ,
  o34 = l1 & (m1 & ~k4),
  o35 = g4 | h4,
  r4 = \[3] ,
  r5 = \[29] ,
  r6 = \[55] ,
  r7 = \[81] ,
  r8 = \[107] ,
  r9 = \[133] ,
  s4 = \[4] ,
  s5 = \[30] ,
  s6 = \[56] ,
  s7 = \[82] ,
  s8 = \[108] ,
  s9 = \[134] ,
  t4 = u3,
  t5 = \[31] ,
  t6 = \[57] ,
  t7 = \[83] ,
  t8 = \[109] ,
  t9 = \[135] ,
  u4 = v3,
  u5 = \[32] ,
  u6 = \[58] ,
  u7 = \[84] ,
  u8 = \[110] ,
  u9 = \[136] ,
  v4 = \[7] ,
  v5 = \[33] ,
  v6 = \[59] ,
  v7 = \[85] ,
  v8 = \[111] ,
  v9 = \[137] ,
  w4 = \[8] ,
  w5 = \[34] ,
  w6 = \[60] ,
  w7 = \[86] ,
  w8 = \[112] ,
  w9 = \[138] ,
  x4 = \[9] ,
  x5 = \[35] ,
  x6 = \[61] ,
  x7 = \[87] ,
  x8 = \[113] ,
  y4 = \[10] ,
  y5 = \[36] ,
  y6 = \[62] ,
  y7 = \[88] ,
  y8 = \[114] ,
  z4 = \[11] ,
  z5 = \[37] ,
  z6 = \[63] ,
  z7 = \[89] ,
  z8 = \[115] ,
  p16 = (m1 & ~g15) | (~o0 | q0),
  p18 = ~x1 & l4,
  p20 = (~w16 & (~t15 & ~g2)) | ~q20,
  p23 = ~w23 | (m0 | n0),
  p24 = y2 & l4,
  p25 = ~t25 & (~i1 & ~j1),
  p26 = q0 | ~h3,
  p27 = j25 | (~r3 | ~k4),
  p28 = (~g25 & (~h1 & ~i1)) | ~q28,
  p29 = z3 & (~a4 & l4),
  p30 = a4 | (b4 | ~l4),
  p31 = q0 | (g1 | ~g4),
  p32 = (~l1 & ~k1) | ((~l1 & ~v0) | (~k1 & ~w0)),
  p33 = ~m0 & ~r3,
  p34 = h1 & l4,
  p35 = h1 | (i1 | j1),
  a17 = ~q35 & (~b4 & ~c4),
  a18 = ~u1 & l4,
  a20 = (~w16 & (~t15 & ~d2)) | ~b20,
  a21 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & b0))),
  a22 = (t15 & (~n0 & ~m0)) | ((l4 & ~a17) | m2),
  a23 = (o & (~l0 & k0)) | ((g & l0) | (g & ~k0)),
  a24 = (~t23 & (t2 & ~l4)) | (~s23 & (~r23 & j)),
  a25 = ~o0 | (q0 | ~l25),
  a26 = q0 | ~c3,
  a27 = j25 | (~m3 | ~k4),
  a29 = (~a17 & (x3 & l4)) | ~b29,
  a30 = q0 | ~b4,
  a32 = (~c32 & (~b32 & l25)) | (~n0 & t15),
  a33 = ~q30 | (~b33 | ~o0),
  a34 = (~l3 & (~l0 & ~k0)) | ((~l3 & (l0 & k0)) | ~m0),
  \[10]  = (~w33 & (~l0 & ~k0)) | ((~w33 & (l0 & k0)) | (~w33 & p3)),
  \[11]  = (~x33 & (~l0 & ~k0)) | ((~x33 & (l0 & k0)) | (~x33 & q3)),
  \[12]  = (~y33 & (~l0 & ~k0)) | ((~y33 & (l0 & k0)) | (~y33 & r3)),
  \[13]  = (~z33 & (~l0 & ~k0)) | ((~z33 & (l0 & k0)) | (~z33 & s3)),
  \[14]  = (~a34 & (~l0 & ~k0)) | ((~a34 & (l0 & k0)) | (~a34 & t3)),
  q17 = ~s1 & l4,
  q19 = (~w16 & (~t15 & ~b2)) | ~r19,
  \[15]  = m0 & m3,
  q20 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & z))),
  q21 = (~k21 & (~s21 & ~a17)) | ((~r21 & (~s16 & ~m0)) | ~t21),
  q23 = (~t23 & (s2 & ~l4)) | (~s23 & (~r23 & i)),
  q24 = (~t23 & (x2 & ~l4)) | (~s23 & (~r23 & n)),
  q25 = ~j1 & (~k1 & ~l1),
  q27 = q0 | ~q3,
  q28 = (~l1 & ~k1) | ~j1,
  q29 = ~w29 | (a17 | x3),
  \[16]  = m0 & n3,
  q30 = y3 & (z3 & ~a4),
  q31 = (~u31 & (~k31 & l25)) | (~n0 & t15),
  q32 = ~q25 | (~s0 | i1),
  q33 = (~i3 & ~a3) | ((~i3 & l0) | (~a3 & ~l0)),
  q34 = i1 & l4,
  q35 = ~w34 | (x3 | ~y3),
  \[17]  = m0 & o3,
  \[18]  = m0 & p3,
  \[19]  = m0 & q3,
  b16 = (~e1 & ~d1) | ((~e1 & c1) | (~d1 & ~c1)),
  b17 = ~p1 & l4,
  b19 = (~w16 & (~t15 & ~y1)) | ~c19,
  b20 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & w))),
  b23 = r2 | ~l4,
  b25 = j25 | (~b3 | ~k4),
  b27 = q0 | ~l3,
  b28 = j25 | (~v3 | ~k4),
  b29 = (~q0 & (o0 & ~t15)) | (~q0 & (o0 & n0)),
  b30 = (~f30 & (~e30 & ~a17)) | (~n0 & t15),
  b31 = ~f31 & (l25 & ~j25),
  b32 = j25 | (d4 | ~e4),
  b33 = ~q0 & m1,
  b34 = ~n0 & (h1 & ~k4),
  b35 = (~d35 & (z0 & y0)) | ((~d35 & (z0 & ~i1)) | ((~d35 & (~j1 & y0)) | (~d35 & (~j1 & ~i1)))),
  \[20]  = m0 & r3,
  \[21]  = m0 & s3,
  \[22]  = m0 & t3,
  \[23]  = g1 & ~j4,
  r16 = ~o1 & l4,
  r18 = (~w16 & (~t15 & ~w1)) | ~s18,
  r19 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & u))),
  \[25]  = ~b34,
  r21 = (j & (~l0 & k0)) | ((b & l0) | (b & ~k0)),
  r23 = m0 | (n0 | ~t15),
  r25 = (~s25 & ~q25) | ((~s25 & h1) | (~s25 & i1)),
  r26 = j25 | (~j3 | ~k4),
  r28 = h1 & ~i1,
  r29 = (~t29 & (~s23 & t15)) | ((~t29 & (~s23 & a4)) | ((~t29 & (~t15 & a4)) | ((~t29 & (t15 & m0)) | (~t29 & (a4 & m0))))),
  \[26]  = ~c34,
  r30 = ~b4 & (~c4 & l4),
  r31 = ~s31 | (q0 | ~t15),
  r32 = (~s32 & (~u0 & ~h1)) | ((~t32 & i1) | ~u32),
  r33 = (~i3 & ~a3) | ((~i3 & ~l0) | (~a3 & l0)),
  r34 = j1 & l4,
  r35 = ~e4 | (~f4 | g4),
  \[27]  = ~d34,
  \[28]  = ~e34,
  \[29]  = ~f34,
  c16 = ~d16 | (~o0 | q0),
  c18 = (~w16 & (~t15 & ~t1)) | ~d18,
  c19 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & r))),
  c21 = ~k2 & l4,
  c23 = (t15 & (~n0 & ~m0)) | ((l4 & ~a17) | q2),
  c24 = (~e24 & (~d24 & ~a17)) | ((~e24 & (~d24 & ~u2)) | ((~e24 & (a17 & ~u2)) | (~e24 & ~p23))),
  c25 = (~q25 & i1) | ((~p25 & h1) | ~r25),
  c26 = j25 | (~e3 | ~k4),
  c28 = q0 | ~u3,
  c30 = ~d30 | (q0 | ~t15),
  c31 = ~d31 & (~g1 & ~q0),
  c32 = ~f4 | (g4 | ~k4),
  c33 = ~o0 | (q0 | a17),
  c34 = ~n0 & (i1 & ~k4),
  \[30]  = (~i34 & ~h34) | ((~i34 & ~g34) | ((~i34 & ~g30) | ((n1 & ~h34) | ((n1 & ~g34) | (n1 & ~g30))))),
  \[31]  = (~i34 & ~h34) | ((~i34 & ~g34) | ((~i34 & ~g30) | ((n1 & ~h34) | ((n1 & ~g34) | (n1 & ~g30))))),
  \[32]  = (~i34 & ~h34) | ((~i34 & ~g34) | ((~i34 & ~g30) | ((n1 & ~h34) | ((n1 & ~g34) | (n1 & ~g30))))),
  \[33]  = (~i34 & ~h34) | ((~i34 & ~g34) | ((~i34 & ~g30) | ((n1 & ~h34) | ((n1 & ~g34) | (n1 & ~g30))))),
  \[34]  = (~i34 & ~h34) | ((~i34 & ~g34) | ((~i34 & ~g30) | ((n1 & ~h34) | ((n1 & ~g34) | (n1 & ~g30))))),
  s16 = n0 | ~t15,
  s17 = (~w16 & (~t15 & ~r1)) | ~t17,
  s18 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & l0))),
  \[35]  = ~k34,
  s20 = ~i2 & l4,
  s21 = m2 | ~l4,
  s22 = (~k21 & (~u22 & ~a17)) | ((~t22 & (~s16 & ~m0)) | ~v22),
  s23 = (~l0 & k0) | (l0 & ~k0),
  s24 = (~u24 & (~t24 & ~a17)) | ((~u24 & (~t24 & ~y2)) | ((~u24 & (a17 & ~y2)) | (~u24 & ~p23))),
  s25 = (l1 & k1) | ((l1 & j1) | (k1 & j1)),
  s26 = q0 | ~i3,
  s27 = j25 | (~s3 | ~k4),
  s28 = (t0 & (~g25 & i1)) | (~u28 & ~i1),
  \[36]  = ~l34,
  s31 = ~t31 & o0,
  s32 = i1 | (k1 | l1),
  s33 = ~m0 & ~q3,
  s34 = k1 & l4,
  \[37]  = ~m34,
  \[38]  = ~n34,
  \[39]  = ~o34,
  d16 = (t15 & (~e1 & ~n0)) | j1,
  d17 = (~w16 & (~t15 & ~o1)) | ~e17,
  d18 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & d0))),
  d20 = ~f2 & l4,
  d24 = v2 & l4,
  d25 = q0 | ~a3,
  d26 = q0 | ~d3,
  d27 = j25 | (~n3 | ~k4),
  d29 = ~a17 & (~x3 & l4),
  d30 = m0 & (~n0 & o0),
  d31 = (~e31 & (l25 & ~j25)) | (~n0 & t15),
  d32 = ~j25 & ~g1,
  d33 = (~x0 & h1) | (~b35 | ~n4),
  d34 = ~n0 & (j1 & ~k4),
  d35 = (~b1 & l1) | ((~a1 & k1) | ~e35),
  \[40]  = ~p34,
  \[41]  = ~q34,
  \[42]  = ~r34,
  \[43]  = ~s34,
  \[44]  = ~t34,
  t15 = ~p35 & (~k1 & ~l1),
  t17 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & f0))),
  t19 = ~d2 & l4,
  \[45]  = ~h1,
  t21 = (t15 & (~n0 & ~m0)) | ((l4 & ~a17) | l2),
  t22 = (n & (~l0 & k0)) | ((f & l0) | (f & ~k0)),
  t23 = ~u23 & (~m0 & ~n0),
  t24 = z2 & l4,
  t25 = k1 | l1,
  t27 = q0 | ~r3,
  t29 = (~v29 & (~u29 & ~t15)) | (n0 & t15),
  \[46]  = ~i1,
  t30 = q0 | g1,
  t31 = (m0 & (~l0 & k0)) | ((m0 & (l0 & ~k0)) | n0),
  t32 = ~t25 & (t0 & ~j1),
  t33 = (~e3 & (~l0 & ~k0)) | ((~e3 & (l0 & k0)) | ~m0),
  t34 = l1 & l4,
  \[47]  = ~j1,
  \[48]  = ~k1,
  \[49]  = ~l1,
  e17 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & i0))),
  e19 = ~a2 & l4,
  e21 = (~w16 & (~t15 & ~j2)) | ~f21,
  e22 = (~k21 & (~g22 & ~a17)) | ((~f22 & (~s16 & ~m0)) | ~h22),
  e24 = (~t23 & (u2 & ~l4)) | (~s23 & (~r23 & k)),
  e25 = (~h25 & (~g25 & ~f25)) | ((~h25 & (~g25 & ~h1)) | ((~h25 & (~i1 & ~f25)) | (~h25 & (~i1 & ~h1)))),
  e27 = q0 | ~m3,
  e28 = j25 | (~w3 | ~k4),
  e29 = (~f29 & (~q0 & n0)) | (~f29 & (~q0 & ~t15)),
  e30 = x3 | ~y3,
  e31 = d4 | (e4 | ~k4),
  e32 = ~d4 & (e4 & f4),
  e33 = (d33 & ~l25) | (~o0 | q0),
  e34 = ~n0 & (k1 & ~k4),
  e35 = ~f35 | h4,
  \[51]  = (~i4 & ~f1) | (i4 & f1),
  \[52]  = ~v34 & (~b4 & ~c4),
  \[53]  = o0 & (~q0 & ~g15),
  \[54]  = (~m15 & (~l15 & o0)) | (~k15 & (~j15 & ~n0)),
  u16 = a17 | ~l4,
  u18 = ~y1 & l4,
  \[55]  = (~y15 & (~x15 & ~w15)) | ((~y15 & (~x15 & n0)) | ((~y15 & (~x15 & ~t15)) | ((~y15 & (~g1 & ~w15)) | ((~y15 & (~g1 & n0)) | (~y15 & (~g1 & ~t15)))))),
  u20 = (~w16 & (~t15 & ~h2)) | ~v20,
  u22 = q2 | ~l4,
  u23 = (~l0 & k0) | ((l0 & ~k0) | ~t15),
  u24 = (~t23 & (y2 & ~l4)) | (~s23 & (~r23 & o)),
  u26 = j25 | (~k3 | ~k4),
  u28 = (~w28 & (~v28 & ~o25)) | ((~w28 & (~v28 & ~j1)) | ((~w28 & (~v28 & ~u0)) | ((~w28 & (~o25 & j1)) | ((~w28 & (~o25 & ~w0)) | ((~w28 & (~j1 & ~w0)) | ((~w28 & (j1 & ~u0)) | (~w28 & (~w0 & ~u0)))))))),
  u29 = a17 | x3,
  \[56]  = (~c16 & (~x15 & ~b16)) | ((~c16 & (~x15 & n0)) | ((~c16 & (~x15 & ~t15)) | ((~c16 & (~g1 & ~b16)) | ((~c16 & (~g1 & n0)) | (~c16 & (~g1 & ~t15)))))),
  u30 = (~w30 & (l25 & ~j25)) | (~x30 & ~d4),
  u31 = ~e4 | (~f4 | ~k4),
  u32 = ~w32 & (k4 & n4),
  u33 = (~f3 & (~l0 & ~k0)) | ((~f3 & (l0 & k0)) | ~m0),
  \[57]  = (~g16 & (~x15 & ~f16)) | ((~g16 & (~x15 & n0)) | ((~g16 & (~x15 & ~t15)) | ((~g16 & (~g1 & ~f16)) | ((~g16 & (~g1 & n0)) | (~g16 & (~g1 & ~t15)))))),
  \[58]  = (~l16 & (l1 & ~g1)) | (~l16 & ~j16),
  \[59]  = (~p16 & (p0 & ~n0)) | (~p16 & m1),
  f16 = (~e1 & ~d1) | ((~e1 & ~c1) | (~d1 & ~c1)),
  f18 = ~v1 & l4,
  f20 = (~w16 & (~t15 & ~e2)) | ~g20,
  f21 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & c0))),
  f22 = (l & (~l0 & k0)) | ((d & l0) | (d & ~k0)),
  f25 = ~o25 | (i1 | j1),
  f26 = j25 | (~f3 | ~k4),
  f28 = q0 | ~v3,
  f29 = ~g29 & l4,
  f30 = ~z3 | (a4 | ~l4),
  f31 = d4 | ~k4,
  f32 = ~g4 & (~h4 & k4),
  f34 = ~n0 & (l1 & ~k4),
  f35 = e4 & (f4 & ~g4),
  \[60]  = (~v16 & (~u16 & ~s16)) | ((~v16 & (~u16 & ~r16)) | ((~v16 & (~u16 & a17)) | ((~v16 & (~n0 & ~s16)) | ((~v16 & (~n0 & ~r16)) | ((~v16 & (~n0 & a17)) | ((~v16 & (n1 & ~s16)) | ((~v16 & (n1 & ~r16)) | (~v16 & (n1 & a17))))))))),
  \[61]  = (~d17 & (~u16 & ~s16)) | ((~d17 & (~u16 & ~b17)) | ((~d17 & (~u16 & a17)) | ((~d17 & (~n0 & ~s16)) | ((~d17 & (~n0 & ~b17)) | ((~d17 & (~n0 & a17)) | ((~d17 & (o1 & ~s16)) | ((~d17 & (o1 & ~b17)) | (~d17 & (o1 & a17))))))))),
  \[62]  = (~i17 & (~u16 & ~s16)) | ((~i17 & (~u16 & ~g17)) | ((~i17 & (~u16 & a17)) | ((~i17 & (~n0 & ~s16)) | ((~i17 & (~n0 & ~g17)) | ((~i17 & (~n0 & a17)) | ((~i17 & (p1 & ~s16)) | ((~i17 & (p1 & ~g17)) | (~i17 & (p1 & a17))))))))),
  \[63]  = (~n17 & (~u16 & ~s16)) | ((~n17 & (~u16 & ~l17)) | ((~n17 & (~u16 & a17)) | ((~n17 & (~n0 & ~s16)) | ((~n17 & (~n0 & ~l17)) | ((~n17 & (~n0 & a17)) | ((~n17 & (q1 & ~s16)) | ((~n17 & (q1 & ~l17)) | (~n17 & (q1 & a17))))))))),
  \[64]  = (~s17 & (~u16 & ~s16)) | ((~s17 & (~u16 & ~q17)) | ((~s17 & (~u16 & a17)) | ((~s17 & (~n0 & ~s16)) | ((~s17 & (~n0 & ~q17)) | ((~s17 & (~n0 & a17)) | ((~s17 & (r1 & ~s16)) | ((~s17 & (r1 & ~q17)) | (~s17 & (r1 & a17))))))))),
  v16 = (~w16 & (~t15 & ~n1)) | ~x16,
  v17 = ~t1 & l4,
  v19 = (~w16 & (~t15 & ~c2)) | ~w19,
  \[65]  = (~x17 & (~u16 & ~s16)) | ((~x17 & (~u16 & ~v17)) | ((~x17 & (~u16 & a17)) | ((~x17 & (~n0 & ~s16)) | ((~x17 & (~n0 & ~v17)) | ((~x17 & (~n0 & a17)) | ((~x17 & (s1 & ~s16)) | ((~x17 & (s1 & ~v17)) | (~x17 & (s1 & a17))))))))),
  v20 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & a0))),
  v22 = (t15 & (~n0 & ~m0)) | ((l4 & ~a17) | p2),
  v26 = q0 | ~j3,
  v27 = j25 | (~t3 | ~k4),
  v28 = ~k1 & l1,
  v29 = ~y3 | (~z3 | ~l4),
  \[66]  = (~c18 & (~u16 & ~s16)) | ((~c18 & (~u16 & ~a18)) | ((~c18 & (~u16 & a17)) | ((~c18 & (~n0 & ~s16)) | ((~c18 & (~n0 & ~a18)) | ((~c18 & (~n0 & a17)) | ((~c18 & (t1 & ~s16)) | ((~c18 & (t1 & ~a18)) | (~c18 & (t1 & a17))))))))),
  v30 = q0 | ~t15,
  v31 = ~g1 & (~d4 & e4),
  v33 = (~g3 & (~l0 & ~k0)) | ((~g3 & (l0 & k0)) | ~m0),
  v34 = ~w34 | (~x3 | ~y3),
  \[67]  = (~h18 & (~u16 & ~s16)) | ((~h18 & (~u16 & ~f18)) | ((~h18 & (~u16 & a17)) | ((~h18 & (~n0 & ~s16)) | ((~h18 & (~n0 & ~f18)) | ((~h18 & (~n0 & a17)) | ((~h18 & (u1 & ~s16)) | ((~h18 & (u1 & ~f18)) | (~h18 & (u1 & a17))))))))),
  \[68]  = (~m18 & (~u16 & ~s16)) | ((~m18 & (~u16 & ~k18)) | ((~m18 & (~u16 & a17)) | ((~m18 & (~n0 & ~s16)) | ((~m18 & (~n0 & ~k18)) | ((~m18 & (~n0 & a17)) | ((~m18 & (v1 & ~s16)) | ((~m18 & (v1 & ~k18)) | (~m18 & (v1 & a17))))))))),
  \[69]  = (~r18 & (~u16 & ~s16)) | ((~r18 & (~u16 & ~p18)) | ((~r18 & (~u16 & a17)) | ((~r18 & (~n0 & ~s16)) | ((~r18 & (~n0 & ~p18)) | ((~r18 & (~n0 & a17)) | ((~r18 & (w1 & ~s16)) | ((~r18 & (w1 & ~p18)) | (~r18 & (w1 & a17))))))))),
  g15 = (~g35 & (i1 & ~y0)) | ((~g35 & (h1 & ~x0)) | ~h35),
  g16 = ~h16 | (~o0 | q0),
  g17 = ~q1 & l4,
  g19 = (~w16 & (~t15 & ~z1)) | ~h19,
  g20 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & \x ))),
  g22 = o2 | ~l4,
  g23 = (~k21 & (~i23 & ~a17)) | ((~h23 & (~s16 & ~m0)) | ~j23),
  g24 = (~i24 & (~h24 & ~a17)) | ((~i24 & (~h24 & ~v2)) | ((~i24 & (a17 & ~v2)) | (~i24 & ~p23))),
  g25 = j1 | (k1 | l1),
  g26 = q0 | ~e3,
  g27 = j25 | (~o3 | ~k4),
  g29 = a17 | (x3 | y3),
  g30 = y3 & z3,
  g34 = ~a4 & (~b4 & ~c4),
  g35 = ~o35 & (e4 & f4),
  \[70]  = (~w18 & (~u16 & ~s16)) | ((~w18 & (~u16 & ~u18)) | ((~w18 & (~u16 & a17)) | ((~w18 & (~n0 & ~s16)) | ((~w18 & (~n0 & ~u18)) | ((~w18 & (~n0 & a17)) | ((~w18 & (x1 & ~s16)) | ((~w18 & (x1 & ~u18)) | (~w18 & (x1 & a17))))))))),
  \[71]  = (~b19 & (~u16 & ~s16)) | ((~b19 & (~u16 & ~z18)) | ((~b19 & (~u16 & a17)) | ((~b19 & (~n0 & ~s16)) | ((~b19 & (~n0 & ~z18)) | ((~b19 & (~n0 & a17)) | ((~b19 & (y1 & ~s16)) | ((~b19 & (y1 & ~z18)) | (~b19 & (y1 & a17))))))))),
  \[72]  = (~g19 & (~u16 & ~s16)) | ((~g19 & (~u16 & ~e19)) | ((~g19 & (~u16 & a17)) | ((~g19 & (~n0 & ~s16)) | ((~g19 & (~n0 & ~e19)) | ((~g19 & (~n0 & a17)) | ((~g19 & (z1 & ~s16)) | ((~g19 & (z1 & ~e19)) | (~g19 & (z1 & a17))))))))),
  \[73]  = (~l19 & (~u16 & ~s16)) | ((~l19 & (~u16 & ~j19)) | ((~l19 & (~u16 & a17)) | ((~l19 & (~n0 & ~s16)) | ((~l19 & (~n0 & ~j19)) | ((~l19 & (~n0 & a17)) | ((~l19 & (a2 & ~s16)) | ((~l19 & (a2 & ~j19)) | (~l19 & (a2 & a17))))))))),
  \[74]  = (~q19 & (~u16 & ~s16)) | ((~q19 & (~u16 & ~o19)) | ((~q19 & (~u16 & a17)) | ((~q19 & (~n0 & ~s16)) | ((~q19 & (~n0 & ~o19)) | ((~q19 & (~n0 & a17)) | ((~q19 & (b2 & ~s16)) | ((~q19 & (b2 & ~o19)) | (~q19 & (b2 & a17))))))))),
  w15 = (~e1 & d1) | ((~e1 & ~c1) | (~d1 & ~c1)),
  w16 = ~a17 & l4,
  w18 = (~w16 & (~t15 & ~x1)) | ~x18,
  w19 = (~q0 & (o0 & ~t15)) | ((~q0 & (o0 & n0)) | (~q0 & (o0 & v))),
  \[75]  = (~v19 & (~u16 & ~s16)) | ((~v19 & (~u16 & ~t19)) | ((~v19 & (~u16 & a17)) | ((~v19 & (~n0 & ~s16)) | ((~v19 & (~n0 & ~t19)) | ((~v19 & (~n0 & a17)) | ((~v19 & (c2 & ~s16)) | ((~v19 & (c2 & ~t19)) | (~v19 & (c2 & a17))))))))),
  w23 = (t15 & (~l0 & ~k0)) | (t15 & (l0 & k0)),
  w24 = ~p | (m0 | n0),
  w25 = j25 | (~c3 | ~k4),
  w27 = q0 | ~s3,
  w28 = ~x28 & ~l1,
  w29 = y3 & (z3 & l4),
  \[76]  = (~a20 & (~u16 & ~s16)) | ((~a20 & (~u16 & ~y19)) | ((~a20 & (~u16 & a17)) | ((~a20 & (~n0 & ~s16)) | ((~a20 & (~n0 & ~y19)) | ((~a20 & (~n0 & a17)) | ((~a20 & (d2 & ~s16)) | ((~a20 & (d2 & ~y19)) | (~a20 & (d2 & a17))))))))),
  w30 = ~d4 | ~k4,
  w31 = f4 & (~g4 & k4),
  w32 = (k1 & l1) | (~x32 | ~l25),
  w33 = (~h3 & (~l0 & ~k0)) | ((~h3 & (l0 & k0)) | ~m0),
  w34 = z3 & ~a4;
endmodule

