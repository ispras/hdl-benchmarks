module reduce_or_1s(a, b);
  input signed a;
  output signed b;
  assign b = |a;
endmodule
