// IWLS benchmark module "i7" printed on Wed May 29 17:26:49 2002
module i7(\V199(1) , \V32(27) , \V199(0) , \V32(26) , \V32(25) , \V32(24) , \V32(23) , \V32(22) , \V32(21) , \V32(20) , \V32(19) , \V32(18) , \V32(17) , \V32(16) , \V32(15) , \V32(14) , \V32(13) , \V32(12) , \V32(11) , \V32(10) , \V32(9) , \V32(8) , \V32(7) , \V32(6) , \V32(5) , \V32(4) , \V32(3) , \V32(2) , \V32(1) , \V32(0) , \V96(27) , \V96(26) , \V96(25) , \V96(24) , \V96(23) , \V96(22) , \V96(21) , \V96(20) , \V96(19) , \V96(18) , \V96(17) , \V96(16) , \V96(15) , \V96(14) , \V96(13) , \V96(12) , \V96(11) , \V96(10) , \V96(9) , \V96(8) , \V96(7) , \V96(6) , \V96(5) , \V96(4) , \V96(3) , \V96(2) , \V96(1) , \V96(0) , \V64(27) , \V64(26) , \V64(25) , \V64(24) , \V64(23) , \V64(22) , \V64(21) , \V64(20) , \V64(19) , \V64(18) , \V64(17) , \V64(16) , \V64(15) , \V64(14) , \V64(13) , \V64(12) , \V64(11) , \V64(10) , \V64(9) , \V64(8) , \V64(7) , \V64(6) , \V64(5) , \V64(4) , \V64(3) , \V64(2) , \V64(1) , \V64(0) , \V128(27) , \V199(4) , \V128(26) , \V128(25) , \V128(24) , \V128(23) , \V128(22) , \V128(21) , \V128(20) , \V128(19) , \V128(18) , \V128(17) , \V128(16) , \V128(15) , \V128(14) , \V128(13) , \V128(12) , \V128(11) , \V128(10) , \V128(9) , \V128(8) , \V128(7) , \V128(6) , \V128(5) , \V128(4) , \V128(3) , \V128(2) , \V128(1) , \V128(0) , \V32(31) , \V32(30) , \V32(29) , \V32(28) , \V192(27) , \V192(26) , \V192(25) , \V192(24) , \V192(23) , \V192(22) , \V192(21) , \V192(20) , \V192(19) , \V192(18) , \V192(17) , \V192(16) , \V192(15) , \V192(14) , \V192(13) , \V192(12) , \V192(11) , \V192(10) , \V192(9) , \V192(8) , \V192(7) , \V192(6) , \V192(5) , \V192(4) , \V192(3) , \V192(2) , \V192(1) , \V192(0) , \V96(31) , \V96(30) , \V96(29) , \V96(28) , \V160(27) , \V160(26) , \V160(25) , \V160(24) , \V160(23) , \V160(22) , \V160(21) , \V160(20) , \V160(19) , \V160(18) , \V160(17) , \V160(16) , \V160(15) , \V160(14) , \V160(13) , \V160(12) , \V160(11) , \V160(10) , \V160(9) , \V160(8) , \V160(7) , \V160(6) , \V160(5) , \V160(4) , \V160(3) , \V160(2) , \V160(1) , \V160(0) , \V64(31) , \V64(30) , \V64(29) , \V64(28) , \V128(31) , \V199(3) , \V128(30) , \V128(29) , \V128(28) , \V195(0) , \V194(1) , \V194(0) , \V192(31) , \V192(30) , \V192(29) , \V192(28) , \V160(31) , \V160(30) , \V160(29) , \V160(28) , \V227(27) , \V227(26) , \V227(25) , \V227(24) , \V227(23) , \V227(22) , \V227(21) , \V227(20) , \V227(19) , \V227(18) , \V227(17) , \V227(16) , \V227(15) , \V227(14) , \V227(13) , \V227(12) , \V227(11) , \V227(10) , \V227(9) , \V227(8) , \V227(7) , \V227(6) , \V227(5) , \V227(4) , \V227(3) , \V227(2) , \V227(1) , \V227(0) , \V259(31) , \V259(30) , \V259(29) , \V259(28) , \V259(27) , \V259(26) , \V259(25) , \V259(24) , \V259(23) , \V259(22) , \V259(21) , \V259(20) , \V259(19) , \V259(18) , \V259(17) , \V259(16) , \V259(15) , \V259(14) , \V259(13) , \V259(12) , \V259(11) , \V259(10) , \V259(9) , \V259(8) , \V259(7) , \V259(6) , \V259(5) , \V259(4) , \V259(3) , \V259(2) , \V259(1) , \V259(0) , \V266(6) , \V266(5) , \V266(4) , \V266(3) , \V266(2) , \V266(1) , \V266(0) );
input
  \V160(21) ,
  \V160(20) ,
  \V160(23) ,
  \V160(22) ,
  \V128(27) ,
  \V160(25) ,
  \V128(26) ,
  \V160(24) ,
  \V128(29) ,
  \V160(17) ,
  \V128(28) ,
  \V160(16) ,
  \V160(19) ,
  \V160(18) ,
  \V96(0) ,
  \V96(1) ,
  \V64(13) ,
  \V96(2) ,
  \V64(12) ,
  \V96(3) ,
  \V64(15) ,
  \V128(21) ,
  \V96(4) ,
  \V64(14) ,
  \V128(20) ,
  \V96(5) ,
  \V128(23) ,
  \V160(11) ,
  \V96(6) ,
  \V128(22) ,
  \V160(10) ,
  \V96(7) ,
  \V64(11) ,
  \V128(25) ,
  \V160(13) ,
  \V96(8) ,
  \V64(10) ,
  \V128(24) ,
  \V192(3) ,
  \V160(12) ,
  \V96(9) ,
  \V128(17) ,
  \V192(2) ,
  \V160(15) ,
  \V128(16) ,
  \V192(5) ,
  \V160(14) ,
  \V128(19) ,
  \V192(4) ,
  \V128(18) ,
  \V64(17) ,
  \V64(16) ,
  \V192(1) ,
  \V64(19) ,
  \V192(0) ,
  \V64(18) ,
  \V64(23) ,
  \V64(22) ,
  \V64(25) ,
  \V128(11) ,
  \V64(24) ,
  \V128(10) ,
  \V192(7) ,
  \V128(13) ,
  \V192(6) ,
  \V128(12) ,
  \V192(9) ,
  \V64(21) ,
  \V128(15) ,
  \V192(8) ,
  \V64(20) ,
  \V128(14) ,
  \V64(27) ,
  \V64(26) ,
  \V64(29) ,
  \V64(28) ,
  \V194(1) ,
  \V160(31) ,
  \V194(0) ,
  \V160(30) ,
  \V64(31) ,
  \V64(30) ,
  \V128(3) ,
  \V128(2) ,
  \V128(5) ,
  \V195(0) ,
  \V128(4) ,
  \V128(31) ,
  \V128(30) ,
  \V128(1) ,
  \V128(0) ,
  \V128(7) ,
  \V128(6) ,
  \V128(9) ,
  \V128(8) ,
  \V199(3) ,
  \V199(4) ,
  \V199(1) ,
  \V199(0) ,
  \V32(0) ,
  \V32(1) ,
  \V32(2) ,
  \V32(3) ,
  \V32(13) ,
  \V32(4) ,
  \V32(12) ,
  \V32(5) ,
  \V32(15) ,
  \V32(6) ,
  \V32(14) ,
  \V32(7) ,
  \V32(8) ,
  \V32(9) ,
  \V32(11) ,
  \V32(10) ,
  \V192(27) ,
  \V192(26) ,
  \V192(29) ,
  \V192(28) ,
  \V32(17) ,
  \V32(16) ,
  \V32(19) ,
  \V32(18) ,
  \V32(23) ,
  \V32(22) ,
  \V192(21) ,
  \V32(25) ,
  \V192(20) ,
  \V32(24) ,
  \V192(23) ,
  \V192(22) ,
  \V192(25) ,
  \V32(21) ,
  \V192(24) ,
  \V32(20) ,
  \V192(17) ,
  \V192(16) ,
  \V192(19) ,
  \V192(18) ,
  \V32(27) ,
  \V96(13) ,
  \V32(26) ,
  \V96(12) ,
  \V32(29) ,
  \V96(15) ,
  \V32(28) ,
  \V96(14) ,
  \V192(11) ,
  \V192(10) ,
  \V96(11) ,
  \V192(13) ,
  \V96(10) ,
  \V192(12) ,
  \V192(15) ,
  \V32(31) ,
  \V192(14) ,
  \V32(30) ,
  \V96(17) ,
  \V96(16) ,
  \V96(19) ,
  \V96(18) ,
  \V96(23) ,
  \V96(22) ,
  \V96(25) ,
  \V96(24) ,
  \V96(21) ,
  \V96(20) ,
  \V96(27) ,
  \V96(26) ,
  \V96(29) ,
  \V96(28) ,
  \V192(31) ,
  \V64(0) ,
  \V192(30) ,
  \V96(31) ,
  \V64(1) ,
  \V96(30) ,
  \V64(2) ,
  \V64(3) ,
  \V64(4) ,
  \V64(5) ,
  \V64(6) ,
  \V64(7) ,
  \V64(8) ,
  \V160(3) ,
  \V64(9) ,
  \V160(2) ,
  \V160(5) ,
  \V160(4) ,
  \V160(1) ,
  \V160(0) ,
  \V160(7) ,
  \V160(6) ,
  \V160(9) ,
  \V160(8) ,
  \V160(27) ,
  \V160(26) ,
  \V160(29) ,
  \V160(28) ;
output
  \V259(27) ,
  \V259(26) ,
  \V259(29) ,
  \V259(28) ,
  \V259(21) ,
  \V259(20) ,
  \V259(23) ,
  \V259(22) ,
  \V259(25) ,
  \V259(24) ,
  \V259(17) ,
  \V259(16) ,
  \V259(19) ,
  \V259(18) ,
  \V259(11) ,
  \V259(10) ,
  \V259(13) ,
  \V259(12) ,
  \V259(15) ,
  \V259(14) ,
  \V259(3) ,
  \V259(2) ,
  \V259(5) ,
  \V259(4) ,
  \V259(1) ,
  \V259(0) ,
  \V259(7) ,
  \V259(6) ,
  \V259(9) ,
  \V259(8) ,
  \V259(31) ,
  \V259(30) ,
  \V227(27) ,
  \V227(26) ,
  \V227(21) ,
  \V227(20) ,
  \V227(23) ,
  \V227(22) ,
  \V227(25) ,
  \V227(24) ,
  \V227(17) ,
  \V227(16) ,
  \V227(19) ,
  \V227(18) ,
  \V227(11) ,
  \V227(10) ,
  \V227(13) ,
  \V227(12) ,
  \V227(15) ,
  \V227(14) ,
  \V266(3) ,
  \V266(2) ,
  \V266(5) ,
  \V266(4) ,
  \V266(1) ,
  \V266(0) ,
  \V266(6) ,
  \V227(3) ,
  \V227(2) ,
  \V227(5) ,
  \V227(4) ,
  \V227(1) ,
  \V227(0) ,
  \V227(7) ,
  \V227(6) ,
  \V227(9) ,
  \V227(8) ;
wire
  \V594(1) ,
  \V594(0) ,
  \V596(1) ,
  \V596(0) ,
  \[0] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \[5] ,
  \[6] ,
  \[7] ,
  \[8] ,
  \[9] ,
  V267,
  V268,
  V269,
  V270,
  V271,
  V272,
  V273,
  V274,
  V275,
  V276,
  V277,
  V278,
  V279,
  V280,
  V281,
  V282,
  V283,
  V284,
  V285,
  V286,
  V287,
  V288,
  V289,
  V290,
  V291,
  V292,
  V293,
  V294,
  V295,
  V296,
  V297,
  V298,
  V299,
  \V538(27) ,
  \V538(26) ,
  V300,
  V301,
  V302,
  V303,
  V304,
  V305,
  V306,
  V307,
  V308,
  V309,
  V310,
  V311,
  V312,
  V313,
  V314,
  V315,
  V316,
  V317,
  V318,
  V319,
  V320,
  V321,
  V322,
  V323,
  V324,
  V325,
  V326,
  V327,
  V328,
  V329,
  V330,
  V331,
  V332,
  V333,
  V334,
  V335,
  V336,
  V337,
  V338,
  V339,
  V340,
  V341,
  V342,
  V343,
  V344,
  V345,
  V346,
  V347,
  V348,
  \V538(21) ,
  V349,
  V350,
  V351,
  V352,
  \V538(20) ,
  \V538(23) ,
  \V538(22) ,
  V381,
  V382,
  V383,
  V384,
  V385,
  V386,
  V387,
  V388,
  \V538(25) ,
  V389,
  V390,
  V391,
  V392,
  V393,
  V394,
  V395,
  V396,
  V397,
  V398,
  \V538(24) ,
  V399,
  \V538(17) ,
  \V538(16) ,
  \V538(19) ,
  \V538(18) ,
  V400,
  V401,
  V402,
  V403,
  V404,
  V405,
  V406,
  V407,
  V408,
  V409,
  V410,
  V411,
  V412,
  V413,
  V414,
  V415,
  V416,
  V417,
  V418,
  V419,
  V420,
  V421,
  V422,
  V423,
  V424,
  V425,
  V426,
  V427,
  V428,
  V429,
  V430,
  V431,
  V432,
  V433,
  V434,
  V435,
  V436,
  V437,
  V438,
  V439,
  V440,
  V441,
  V442,
  V443,
  V444,
  V445,
  V446,
  V447,
  V448,
  \V538(11) ,
  V449,
  V450,
  V451,
  V452,
  V453,
  V454,
  V455,
  V456,
  V457,
  V458,
  \V538(10) ,
  V459,
  V460,
  V461,
  V462,
  V463,
  V464,
  V465,
  V466,
  V467,
  V468,
  \V538(13) ,
  V469,
  V470,
  V471,
  V472,
  V473,
  V474,
  V475,
  V476,
  V477,
  V478,
  \V538(12) ,
  V479,
  V480,
  V481,
  V482,
  V483,
  V484,
  V485,
  V486,
  V487,
  V488,
  \V538(15) ,
  V489,
  V490,
  V491,
  V492,
  V493,
  V494,
  V495,
  V496,
  V497,
  V498,
  \V538(14) ,
  V499,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[14] ,
  \[15] ,
  V500,
  V501,
  V502,
  V503,
  V504,
  V505,
  V506,
  \[16] ,
  \[17] ,
  \[18] ,
  V539,
  \[19] ,
  V540,
  V541,
  V542,
  V543,
  V544,
  V545,
  V546,
  V547,
  V548,
  V549,
  V550,
  V551,
  V552,
  V553,
  V554,
  V555,
  V556,
  V557,
  V558,
  V559,
  V560,
  V561,
  V562,
  V563,
  V564,
  V565,
  V566,
  V567,
  V568,
  V569,
  V570,
  V571,
  V572,
  V573,
  V574,
  V575,
  V576,
  V577,
  V578,
  V579,
  V580,
  V581,
  V582,
  V583,
  V584,
  V585,
  V586,
  V587,
  V588,
  V589,
  V590,
  V597,
  V598,
  V599,
  \[20] ,
  \[21] ,
  \[22] ,
  \[23] ,
  \[24] ,
  \[25] ,
  V600,
  V601,
  \V380(3) ,
  V602,
  V603,
  V604,
  V605,
  \[26] ,
  \V380(2) ,
  \[27] ,
  \V380(5) ,
  \[28] ,
  \V380(4) ,
  \[29] ,
  \V380(1) ,
  \V380(0) ,
  \[30] ,
  \[31] ,
  \V380(7) ,
  \[32] ,
  \V380(6) ,
  \[33] ,
  \V380(9) ,
  \[34] ,
  \V380(8) ,
  \[35] ,
  \V380(27) ,
  \[36] ,
  \V380(26) ,
  \[37] ,
  \[38] ,
  \[39] ,
  \V380(21) ,
  \V538(3) ,
  \[40] ,
  \V380(20) ,
  \V538(2) ,
  \[41] ,
  \V380(23) ,
  \V538(5) ,
  \[42] ,
  \V380(22) ,
  \V538(4) ,
  \[43] ,
  \V380(25) ,
  \[44] ,
  \V380(24) ,
  \[45] ,
  \V380(17) ,
  \V538(1) ,
  \[46] ,
  \V380(16) ,
  \V538(0) ,
  \[47] ,
  \V380(19) ,
  \[48] ,
  \V380(18) ,
  \[49] ,
  \V538(7) ,
  \V538(6) ,
  \V538(9) ,
  \V538(8) ,
  \V380(11) ,
  \[50] ,
  \V380(10) ,
  \[51] ,
  \V380(13) ,
  \[52] ,
  \V380(12) ,
  \[53] ,
  \V380(15) ,
  \[54] ,
  \V380(14) ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ,
  \[59] ,
  \[60] ,
  \[61] ,
  \[62] ,
  \[63] ,
  \[64] ,
  \[65] ,
  \[66] ,
  \V510(3) ,
  \V510(2) ,
  \V510(1) ,
  \V510(0) ,
  \V594(3) ,
  \V594(2) ;
assign
  \V594(1)  = ~\V192(29) ,
  \V594(0)  = ~\V192(28) ,
  \V259(27)  = \[32] ,
  \V259(26)  = \[33] ,
  \V259(29)  = \[30] ,
  \V259(28)  = \[31] ,
  \V259(21)  = \[38] ,
  \V259(20)  = \[39] ,
  \V259(23)  = \[36] ,
  \V259(22)  = \[37] ,
  \V259(25)  = \[34] ,
  \V596(1)  = ~\V194(1) ,
  \V259(24)  = \[35] ,
  \V596(0)  = ~\V194(0) ,
  \V259(17)  = \[42] ,
  \V259(16)  = \[43] ,
  \V259(19)  = \[40] ,
  \V259(18)  = \[41] ,
  \V259(11)  = \[48] ,
  \V259(10)  = \[49] ,
  \V259(13)  = \[46] ,
  \V259(12)  = \[47] ,
  \V259(15)  = \[44] ,
  \V259(14)  = \[45] ,
  \[0]  = V381 | (V325 | (V297 | V268)),
  \[1]  = V382 | (V326 | (V298 | V269)),
  \[2]  = V383 | (V327 | (V299 | V270)),
  \[3]  = V384 | (V328 | (V300 | V271)),
  \[4]  = V385 | (V329 | (V301 | V272)),
  \V259(3)  = \[56] ,
  \[5]  = V386 | (V330 | (V302 | V273)),
  \V259(2)  = \[57] ,
  \[6]  = V387 | (V331 | (V303 | V274)),
  \V259(5)  = \[54] ,
  \[7]  = V388 | (V332 | (V304 | V275)),
  \V259(4)  = \[55] ,
  \[8]  = V389 | (V333 | (V305 | V276)),
  \[9]  = V390 | (V334 | (V306 | V277)),
  \V259(1)  = \[58] ,
  \V259(0)  = \[59] ,
  \V259(7)  = \[52] ,
  \V259(6)  = \[53] ,
  \V259(9)  = \[50] ,
  \V259(8)  = \[51] ,
  \V259(31)  = \[28] ,
  \V259(30)  = \[29] ,
  V267 = ~\V199(1) ,
  V268 = \V199(0)  & (V267 & \V32(27) ),
  V269 = \V199(0)  & (V267 & \V32(26) ),
  V270 = \V199(0)  & (V267 & \V32(25) ),
  V271 = \V199(0)  & (V267 & \V32(24) ),
  V272 = \V199(0)  & (V267 & \V32(23) ),
  V273 = \V199(0)  & (V267 & \V32(22) ),
  V274 = \V199(0)  & (V267 & \V32(21) ),
  V275 = \V199(0)  & (V267 & \V32(20) ),
  V276 = \V199(0)  & (V267 & \V32(19) ),
  V277 = \V199(0)  & (V267 & \V32(18) ),
  V278 = \V199(0)  & (V267 & \V32(17) ),
  V279 = \V199(0)  & (V267 & \V32(16) ),
  V280 = \V199(0)  & (V267 & \V32(15) ),
  V281 = \V199(0)  & (V267 & \V32(14) ),
  V282 = \V199(0)  & (V267 & \V32(13) ),
  V283 = \V199(0)  & (V267 & \V32(12) ),
  V284 = \V199(0)  & (V267 & \V32(11) ),
  V285 = \V199(0)  & (V267 & \V32(10) ),
  V286 = \V199(0)  & (V267 & \V32(9) ),
  V287 = \V199(0)  & (V267 & \V32(8) ),
  V288 = \V199(0)  & (V267 & \V32(7) ),
  V289 = \V199(0)  & (V267 & \V32(6) ),
  V290 = \V199(0)  & (V267 & \V32(5) ),
  V291 = \V199(0)  & (V267 & \V32(4) ),
  V292 = \V199(0)  & (V267 & \V32(3) ),
  V293 = \V199(0)  & (V267 & \V32(2) ),
  V294 = \V199(0)  & (V267 & \V32(1) ),
  V295 = \V199(0)  & (V267 & \V32(0) ),
  V296 = ~\V199(0) ,
  V297 = V296 & (V267 & \V96(27) ),
  V298 = V296 & (V267 & \V96(26) ),
  V299 = V296 & (V267 & \V96(25) ),
  \V538(27)  = ~\V192(27) ,
  \V538(26)  = ~\V192(26) ,
  V300 = V296 & (V267 & \V96(24) ),
  V301 = V296 & (V267 & \V96(23) ),
  V302 = V296 & (V267 & \V96(22) ),
  V303 = V296 & (V267 & \V96(21) ),
  V304 = V296 & (V267 & \V96(20) ),
  V305 = V296 & (V267 & \V96(19) ),
  V306 = V296 & (V267 & \V96(18) ),
  V307 = V296 & (V267 & \V96(17) ),
  V308 = V296 & (V267 & \V96(16) ),
  V309 = V296 & (V267 & \V96(15) ),
  V310 = V296 & (V267 & \V96(14) ),
  V311 = V296 & (V267 & \V96(13) ),
  V312 = V296 & (V267 & \V96(12) ),
  V313 = V296 & (V267 & \V96(11) ),
  V314 = V296 & (V267 & \V96(10) ),
  V315 = V296 & (V267 & \V96(9) ),
  V316 = V296 & (V267 & \V96(8) ),
  V317 = V296 & (V267 & \V96(7) ),
  V318 = V296 & (V267 & \V96(6) ),
  V319 = V296 & (V267 & \V96(5) ),
  \V227(27)  = \[0] ,
  V320 = V296 & (V267 & \V96(4) ),
  V321 = V296 & (V267 & \V96(3) ),
  V322 = V296 & (V267 & \V96(2) ),
  V323 = V296 & (V267 & \V96(1) ),
  V324 = V296 & (V267 & \V96(0) ),
  V325 = \V199(0)  & (\V199(1)  & \V64(27) ),
  V326 = \V199(0)  & (\V199(1)  & \V64(26) ),
  V327 = \V199(0)  & (\V199(1)  & \V64(25) ),
  V328 = \V199(0)  & (\V199(1)  & \V64(24) ),
  V329 = \V199(0)  & (\V199(1)  & \V64(23) ),
  \V227(26)  = \[1] ,
  V330 = \V199(0)  & (\V199(1)  & \V64(22) ),
  V331 = \V199(0)  & (\V199(1)  & \V64(21) ),
  V332 = \V199(0)  & (\V199(1)  & \V64(20) ),
  V333 = \V199(0)  & (\V199(1)  & \V64(19) ),
  V334 = \V199(0)  & (\V199(1)  & \V64(18) ),
  V335 = \V199(0)  & (\V199(1)  & \V64(17) ),
  V336 = \V199(0)  & (\V199(1)  & \V64(16) ),
  V337 = \V199(0)  & (\V199(1)  & \V64(15) ),
  V338 = \V199(0)  & (\V199(1)  & \V64(14) ),
  V339 = \V199(0)  & (\V199(1)  & \V64(13) ),
  V340 = \V199(0)  & (\V199(1)  & \V64(12) ),
  V341 = \V199(0)  & (\V199(1)  & \V64(11) ),
  V342 = \V199(0)  & (\V199(1)  & \V64(10) ),
  V343 = \V199(0)  & (\V199(1)  & \V64(9) ),
  V344 = \V199(0)  & (\V199(1)  & \V64(8) ),
  V345 = \V199(0)  & (\V199(1)  & \V64(7) ),
  V346 = \V199(0)  & (\V199(1)  & \V64(6) ),
  V347 = \V199(0)  & (\V199(1)  & \V64(5) ),
  V348 = \V199(0)  & (\V199(1)  & \V64(4) ),
  \V538(21)  = ~\V192(21) ,
  V349 = \V199(0)  & (\V199(1)  & \V64(3) ),
  V350 = \V199(0)  & (\V199(1)  & \V64(2) ),
  V351 = \V199(0)  & (\V199(1)  & \V64(1) ),
  V352 = \V199(0)  & (\V199(1)  & \V64(0) ),
  \V538(20)  = ~\V192(20) ,
  \V538(23)  = ~\V192(23) ,
  \V538(22)  = ~\V192(22) ,
  V381 = V296 & (\V199(1)  & \V380(27) ),
  V382 = V296 & (\V199(1)  & \V380(26) ),
  V383 = V296 & (\V199(1)  & \V380(25) ),
  V384 = V296 & (\V199(1)  & \V380(24) ),
  V385 = V296 & (\V199(1)  & \V380(23) ),
  V386 = V296 & (\V199(1)  & \V380(22) ),
  V387 = V296 & (\V199(1)  & \V380(21) ),
  V388 = V296 & (\V199(1)  & \V380(20) ),
  \V538(25)  = ~\V192(25) ,
  V389 = V296 & (\V199(1)  & \V380(19) ),
  V390 = V296 & (\V199(1)  & \V380(18) ),
  V391 = V296 & (\V199(1)  & \V380(17) ),
  V392 = V296 & (\V199(1)  & \V380(16) ),
  V393 = V296 & (\V199(1)  & \V380(15) ),
  V394 = V296 & (\V199(1)  & \V380(14) ),
  V395 = V296 & (\V199(1)  & \V380(13) ),
  V396 = V296 & (\V199(1)  & \V380(12) ),
  V397 = V296 & (\V199(1)  & \V380(11) ),
  V398 = V296 & (\V199(1)  & \V380(10) ),
  \V538(24)  = ~\V192(24) ,
  V399 = V296 & (\V199(1)  & \V380(9) ),
  \V538(17)  = ~\V192(17) ,
  \V538(16)  = ~\V192(16) ,
  \V227(21)  = \[6] ,
  \V538(19)  = ~\V192(19) ,
  \V227(20)  = \[7] ,
  \V538(18)  = ~\V192(18) ,
  \V227(23)  = \[4] ,
  \V227(22)  = \[5] ,
  \V227(25)  = \[2] ,
  V400 = V296 & (\V199(1)  & \V380(8) ),
  V401 = V296 & (\V199(1)  & \V380(7) ),
  V402 = V296 & (\V199(1)  & \V380(6) ),
  V403 = V296 & (\V199(1)  & \V380(5) ),
  V404 = V296 & (\V199(1)  & \V380(4) ),
  V405 = V296 & (\V199(1)  & \V380(3) ),
  V406 = V296 & (\V199(1)  & \V380(2) ),
  V407 = V296 & (\V199(1)  & \V380(1) ),
  V408 = V296 & (\V199(1)  & \V380(0) ),
  V409 = ~\V199(1) ,
  \V227(24)  = \[3] ,
  V410 = \V199(4)  & (V409 & (\V199(0)  & \V128(27) )),
  V411 = \V199(4)  & (V409 & (\V199(0)  & \V128(26) )),
  V412 = \V199(4)  & (V409 & (\V199(0)  & \V128(25) )),
  V413 = \V199(4)  & (V409 & (\V199(0)  & \V128(24) )),
  V414 = \V199(4)  & (V409 & (\V199(0)  & \V128(23) )),
  V415 = \V199(4)  & (V409 & (\V199(0)  & \V128(22) )),
  V416 = \V199(4)  & (V409 & (\V199(0)  & \V128(21) )),
  V417 = \V199(4)  & (V409 & (\V199(0)  & \V128(20) )),
  V418 = \V199(4)  & (V409 & (\V199(0)  & \V128(19) )),
  V419 = \V199(4)  & (V409 & (\V199(0)  & \V128(18) )),
  \V227(17)  = \[10] ,
  V420 = \V199(4)  & (V409 & (\V199(0)  & \V128(17) )),
  V421 = \V199(4)  & (V409 & (\V199(0)  & \V128(16) )),
  V422 = \V199(4)  & (V409 & (\V199(0)  & \V128(15) )),
  V423 = \V199(4)  & (V409 & (\V199(0)  & \V128(14) )),
  V424 = \V199(4)  & (V409 & (\V199(0)  & \V128(13) )),
  V425 = \V199(4)  & (V409 & (\V199(0)  & \V128(12) )),
  V426 = \V199(4)  & (V409 & (\V199(0)  & \V128(11) )),
  V427 = \V199(4)  & (V409 & (\V199(0)  & \V128(10) )),
  V428 = \V199(4)  & (V409 & (\V199(0)  & \V128(9) )),
  V429 = \V199(4)  & (V409 & (\V199(0)  & \V128(8) )),
  \V227(16)  = \[11] ,
  V430 = \V199(4)  & (V409 & (\V199(0)  & \V128(7) )),
  V431 = \V199(4)  & (V409 & (\V199(0)  & \V128(6) )),
  V432 = \V199(4)  & (V409 & (\V199(0)  & \V128(5) )),
  V433 = \V199(4)  & (V409 & (\V199(0)  & \V128(4) )),
  V434 = \V199(4)  & (V409 & (\V199(0)  & \V128(3) )),
  V435 = \V199(4)  & (V409 & (\V199(0)  & \V128(2) )),
  V436 = \V199(4)  & (V409 & (\V199(0)  & \V128(1) )),
  V437 = \V199(4)  & (V409 & (\V199(0)  & \V128(0) )),
  V438 = \V199(4)  & (V409 & (\V199(0)  & \V32(31) )),
  V439 = \V199(4)  & (V409 & (\V199(0)  & \V32(30) )),
  \V227(19)  = \[8] ,
  V440 = \V199(4)  & (V409 & (\V199(0)  & \V32(29) )),
  V441 = \V199(4)  & (V409 & (\V199(0)  & \V32(28) )),
  V442 = ~\V199(0) ,
  V443 = \V199(4)  & (V409 & (V442 & \V192(27) )),
  V444 = \V199(4)  & (V409 & (V442 & \V192(26) )),
  V445 = \V199(4)  & (V409 & (V442 & \V192(25) )),
  V446 = \V199(4)  & (V409 & (V442 & \V192(24) )),
  V447 = \V199(4)  & (V409 & (V442 & \V192(23) )),
  V448 = \V199(4)  & (V409 & (V442 & \V192(22) )),
  \V538(11)  = ~\V192(11) ,
  V449 = \V199(4)  & (V409 & (V442 & \V192(21) )),
  \V227(18)  = \[9] ,
  V450 = \V199(4)  & (V409 & (V442 & \V192(20) )),
  V451 = \V199(4)  & (V409 & (V442 & \V192(19) )),
  V452 = \V199(4)  & (V409 & (V442 & \V192(18) )),
  V453 = \V199(4)  & (V409 & (V442 & \V192(17) )),
  V454 = \V199(4)  & (V409 & (V442 & \V192(16) )),
  V455 = \V199(4)  & (V409 & (V442 & \V192(15) )),
  V456 = \V199(4)  & (V409 & (V442 & \V192(14) )),
  V457 = \V199(4)  & (V409 & (V442 & \V192(13) )),
  V458 = \V199(4)  & (V409 & (V442 & \V192(12) )),
  \V538(10)  = ~\V192(10) ,
  V459 = \V199(4)  & (V409 & (V442 & \V192(11) )),
  V460 = \V199(4)  & (V409 & (V442 & \V192(10) )),
  V461 = \V199(4)  & (V409 & (V442 & \V192(9) )),
  V462 = \V199(4)  & (V409 & (V442 & \V192(8) )),
  V463 = \V199(4)  & (V409 & (V442 & \V192(7) )),
  V464 = \V199(4)  & (V409 & (V442 & \V192(6) )),
  V465 = \V199(4)  & (V409 & (V442 & \V192(5) )),
  V466 = \V199(4)  & (V409 & (V442 & \V192(4) )),
  V467 = \V199(4)  & (V409 & (V442 & \V192(3) )),
  V468 = \V199(4)  & (V409 & (V442 & \V192(2) )),
  \V538(13)  = ~\V192(13) ,
  V469 = \V199(4)  & (V409 & (V442 & \V192(1) )),
  V470 = \V199(4)  & (V409 & (V442 & \V192(0) )),
  V471 = \V199(4)  & (V409 & (V442 & \V96(31) )),
  V472 = \V199(4)  & (V409 & (V442 & \V96(30) )),
  V473 = \V199(4)  & (V409 & (V442 & \V96(29) )),
  V474 = \V199(4)  & (V409 & (V442 & \V96(28) )),
  V475 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(27) )),
  V476 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(26) )),
  V477 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(25) )),
  V478 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(24) )),
  \V538(12)  = ~\V192(12) ,
  V479 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(23) )),
  V480 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(22) )),
  V481 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(21) )),
  V482 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(20) )),
  V483 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(19) )),
  V484 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(18) )),
  V485 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(17) )),
  V486 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(16) )),
  V487 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(15) )),
  V488 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(14) )),
  \V538(15)  = ~\V192(15) ,
  V489 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(13) )),
  V490 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(12) )),
  V491 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(11) )),
  V492 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(10) )),
  V493 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(9) )),
  V494 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(8) )),
  V495 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(7) )),
  V496 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(6) )),
  V497 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(5) )),
  V498 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(4) )),
  \V538(14)  = ~\V192(14) ,
  V499 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(3) )),
  \[10]  = V391 | (V335 | (V307 | V278)),
  \[11]  = V392 | (V336 | (V308 | V279)),
  \V227(11)  = \[16] ,
  \[12]  = V393 | (V337 | (V309 | V280)),
  \V227(10)  = \[17] ,
  \[13]  = V394 | (V338 | (V310 | V281)),
  \V227(13)  = \[14] ,
  \[14]  = V395 | (V339 | (V311 | V282)),
  \V227(12)  = \[15] ,
  \[15]  = V396 | (V340 | (V312 | V283)),
  \V227(15)  = \[12] ,
  V500 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(2) )),
  V501 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(1) )),
  V502 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V160(0) )),
  V503 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V64(31) )),
  V504 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V64(30) )),
  V505 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V64(29) )),
  V506 = \V199(4)  & (\V199(1)  & (\V199(0)  & \V64(28) )),
  \[16]  = V397 | (V341 | (V313 | V284)),
  \V227(14)  = \[13] ,
  \[17]  = V398 | (V342 | (V314 | V285)),
  \[18]  = V399 | (V343 | (V315 | V286)),
  V539 = \V199(4)  & (\V199(1)  & (V442 & \V538(27) )),
  \[19]  = V400 | (V344 | (V316 | V287)),
  V540 = \V199(4)  & (\V199(1)  & (V442 & \V538(26) )),
  V541 = \V199(4)  & (\V199(1)  & (V442 & \V538(25) )),
  V542 = \V199(4)  & (\V199(1)  & (V442 & \V538(24) )),
  V543 = \V199(4)  & (\V199(1)  & (V442 & \V538(23) )),
  V544 = \V199(4)  & (\V199(1)  & (V442 & \V538(22) )),
  V545 = \V199(4)  & (\V199(1)  & (V442 & \V538(21) )),
  V546 = \V199(4)  & (\V199(1)  & (V442 & \V538(20) )),
  V547 = \V199(4)  & (\V199(1)  & (V442 & \V538(19) )),
  V548 = \V199(4)  & (\V199(1)  & (V442 & \V538(18) )),
  V549 = \V199(4)  & (\V199(1)  & (V442 & \V538(17) )),
  V550 = \V199(4)  & (\V199(1)  & (V442 & \V538(16) )),
  V551 = \V199(4)  & (\V199(1)  & (V442 & \V538(15) )),
  V552 = \V199(4)  & (\V199(1)  & (V442 & \V538(14) )),
  V553 = \V199(4)  & (\V199(1)  & (V442 & \V538(13) )),
  V554 = \V199(4)  & (\V199(1)  & (V442 & \V538(12) )),
  V555 = \V199(4)  & (\V199(1)  & (V442 & \V538(11) )),
  V556 = \V199(4)  & (\V199(1)  & (V442 & \V538(10) )),
  V557 = \V199(4)  & (\V199(1)  & (V442 & \V538(9) )),
  V558 = \V199(4)  & (\V199(1)  & (V442 & \V538(8) )),
  V559 = \V199(4)  & (\V199(1)  & (V442 & \V538(7) )),
  V560 = \V199(4)  & (\V199(1)  & (V442 & \V538(6) )),
  V561 = \V199(4)  & (\V199(1)  & (V442 & \V538(5) )),
  V562 = \V199(4)  & (\V199(1)  & (V442 & \V538(4) )),
  V563 = \V199(4)  & (\V199(1)  & (V442 & \V538(3) )),
  V564 = \V199(4)  & (\V199(1)  & (V442 & \V538(2) )),
  V565 = \V199(4)  & (\V199(1)  & (V442 & \V538(1) )),
  V566 = \V199(4)  & (\V199(1)  & (V442 & \V538(0) )),
  V567 = \V199(4)  & (\V199(1)  & (V442 & \V510(3) )),
  V568 = \V199(4)  & (\V199(1)  & (V442 & \V510(2) )),
  V569 = \V199(4)  & (\V199(1)  & (V442 & \V510(1) )),
  V570 = \V199(4)  & (\V199(1)  & (V442 & \V510(0) )),
  V571 = ~\V199(4) ,
  V572 = V571 & \V199(1) ,
  V573 = ~\V199(1) ,
  V574 = \V199(3)  & (V573 & (\V199(0)  & \V128(31) )),
  V575 = \V199(3)  & (V573 & (\V199(0)  & \V128(30) )),
  V576 = \V199(3)  & (V573 & (\V199(0)  & \V128(29) )),
  V577 = \V199(3)  & (V573 & (\V199(0)  & \V128(28) )),
  V578 = ~\V199(0) ,
  V579 = \V199(3)  & (V573 & (V578 & \V195(0) )),
  V580 = \V199(3)  & (V573 & (V578 & \V194(1) )),
  V581 = \V199(3)  & (V573 & (V578 & \V194(0) )),
  V582 = \V199(3)  & (V573 & (V578 & \V192(31) )),
  V583 = \V199(3)  & (V573 & (V578 & \V192(30) )),
  V584 = \V199(3)  & (V573 & (V578 & \V192(29) )),
  V585 = \V199(3)  & (V573 & (V578 & \V192(28) )),
  V586 = \V199(0)  & (\V199(1)  & \V199(3) ),
  V587 = \V160(31)  & V586,
  V588 = \V160(30)  & V586,
  V589 = \V160(29)  & V586,
  V590 = \V160(28)  & V586,
  V597 = \V199(3)  & (\V199(1)  & (V578 & \V195(0) )),
  V598 = \V199(3)  & (\V199(1)  & (V578 & \V596(1) )),
  V599 = \V199(3)  & (\V199(1)  & (V578 & \V596(0) )),
  \[20]  = V401 | (V345 | (V317 | V288)),
  \[21]  = V402 | (V346 | (V318 | V289)),
  \[22]  = V403 | (V347 | (V319 | V290)),
  \[23]  = V404 | (V348 | (V320 | V291)),
  \[24]  = V405 | (V349 | (V321 | V292)),
  \[25]  = V406 | (V350 | (V322 | V293)),
  V600 = \V199(3)  & (\V199(1)  & (V578 & \V594(3) )),
  V601 = \V199(3)  & (\V199(1)  & (V578 & \V594(2) )),
  \V380(3)  = ~\V96(3) ,
  V602 = \V199(3)  & (\V199(1)  & (V578 & \V594(1) )),
  V603 = \V199(3)  & (\V199(1)  & (V578 & \V594(0) )),
  V604 = ~\V199(3) ,
  V605 = V604 & \V199(1) ,
  \[26]  = V407 | (V351 | (V323 | V294)),
  \V380(2)  = ~\V96(2) ,
  \[27]  = V408 | (V352 | (V324 | V295)),
  \V380(5)  = ~\V96(5) ,
  \[28]  = V572 | (V539 | (V475 | (V443 | V410))),
  \V380(4)  = ~\V96(4) ,
  \[29]  = V572 | (V540 | (V476 | (V444 | V411))),
  \V380(1)  = ~\V96(1) ,
  \V380(0)  = ~\V96(0) ,
  \[30]  = V572 | (V541 | (V477 | (V445 | V412))),
  \[31]  = V572 | (V542 | (V478 | (V446 | V413))),
  \V380(7)  = ~\V96(7) ,
  \[32]  = V572 | (V543 | (V479 | (V447 | V414))),
  \V380(6)  = ~\V96(6) ,
  \[33]  = V572 | (V544 | (V480 | (V448 | V415))),
  \V380(9)  = ~\V96(9) ,
  \[34]  = V572 | (V545 | (V481 | (V449 | V416))),
  \V380(8)  = ~\V96(8) ,
  \[35]  = V572 | (V546 | (V482 | (V450 | V417))),
  \V380(27)  = ~\V96(27) ,
  \[36]  = V572 | (V547 | (V483 | (V451 | V418))),
  \V380(26)  = ~\V96(26) ,
  \[37]  = V572 | (V548 | (V484 | (V452 | V419))),
  \[38]  = V572 | (V549 | (V485 | (V453 | V420))),
  \[39]  = V572 | (V550 | (V486 | (V454 | V421))),
  \V380(21)  = ~\V96(21) ,
  \V538(3)  = ~\V192(3) ,
  \[40]  = V572 | (V551 | (V487 | (V455 | V422))),
  \V380(20)  = ~\V96(20) ,
  \V538(2)  = ~\V192(2) ,
  \[41]  = V572 | (V552 | (V488 | (V456 | V423))),
  \V266(3)  = \[63] ,
  \V380(23)  = ~\V96(23) ,
  \V538(5)  = ~\V192(5) ,
  \[42]  = V572 | (V553 | (V489 | (V457 | V424))),
  \V266(2)  = \[64] ,
  \V380(22)  = ~\V96(22) ,
  \V538(4)  = ~\V192(4) ,
  \[43]  = V572 | (V554 | (V490 | (V458 | V425))),
  \V266(5)  = \[61] ,
  \V380(25)  = ~\V96(25) ,
  \[44]  = V572 | (V555 | (V491 | (V459 | V426))),
  \V266(4)  = \[62] ,
  \V380(24)  = ~\V96(24) ,
  \[45]  = V572 | (V556 | (V492 | (V460 | V427))),
  \V380(17)  = ~\V96(17) ,
  \V538(1)  = ~\V192(1) ,
  \[46]  = V572 | (V557 | (V493 | (V461 | V428))),
  \V380(16)  = ~\V96(16) ,
  \V538(0)  = ~\V192(0) ,
  \[47]  = V572 | (V558 | (V494 | (V462 | V429))),
  \V266(1)  = \[65] ,
  \V380(19)  = ~\V96(19) ,
  \[48]  = V572 | (V559 | (V495 | (V463 | V430))),
  \V266(0)  = \[66] ,
  \V380(18)  = ~\V96(18) ,
  \[49]  = V572 | (V560 | (V496 | (V464 | V431))),
  \V538(7)  = ~\V192(7) ,
  \V538(6)  = ~\V192(6) ,
  \V538(9)  = ~\V192(9) ,
  \V266(6)  = \[60] ,
  \V538(8)  = ~\V192(8) ,
  \V380(11)  = ~\V96(11) ,
  \[50]  = V572 | (V561 | (V497 | (V465 | V432))),
  \V380(10)  = ~\V96(10) ,
  \[51]  = V572 | (V562 | (V498 | (V466 | V433))),
  \V380(13)  = ~\V96(13) ,
  \[52]  = V572 | (V563 | (V499 | (V467 | V434))),
  \V380(12)  = ~\V96(12) ,
  \[53]  = V572 | (V564 | (V500 | (V468 | V435))),
  \V380(15)  = ~\V96(15) ,
  \[54]  = V572 | (V565 | (V501 | (V469 | V436))),
  \V380(14)  = ~\V96(14) ,
  \[55]  = V572 | (V566 | (V502 | (V470 | V437))),
  \[56]  = V572 | (V567 | (V503 | (V471 | V438))),
  \[57]  = V572 | (V568 | (V504 | (V472 | V439))),
  \[58]  = V572 | (V569 | (V505 | (V473 | V440))),
  \[59]  = V572 | (V570 | (V506 | (V474 | V441))),
  \V227(3)  = \[24] ,
  \V227(2)  = \[25] ,
  \[60]  = V579 | V597,
  \V227(5)  = \[22] ,
  \[61]  = V598 | (V586 | (V580 | V605)),
  \V227(4)  = \[23] ,
  \[62]  = V599 | (V586 | (V581 | V605)),
  \[63]  = V605 | (V600 | (V587 | (V582 | V574))),
  \[64]  = V605 | (V601 | (V588 | (V583 | V575))),
  \V227(1)  = \[26] ,
  \[65]  = V605 | (V602 | (V589 | (V584 | V576))),
  \V227(0)  = \[27] ,
  \[66]  = V605 | (V603 | (V590 | (V585 | V577))),
  \V510(3)  = ~\V96(31) ,
  \V227(7)  = \[20] ,
  \V510(2)  = ~\V96(30) ,
  \V227(6)  = \[21] ,
  \V227(9)  = \[18] ,
  \V227(8)  = \[19] ,
  \V510(1)  = ~\V96(29) ,
  \V510(0)  = ~\V96(28) ,
  \V594(3)  = ~\V192(31) ,
  \V594(2)  = ~\V192(30) ;
endmodule

