// IWLS benchmark module "MultiplierB_32" printed on Wed May 29 22:12:35 2002
module MultiplierB_32(\1 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \13 , \14 , \15 , \16 , \17 , \18 , \19 , \20 , \21 , \22 , \23 , \24 , \25 , \26 , \27 , \28 , \29 , \30 , \31 , \32 , \33 , \98 );
input
  \1 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ,
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ,
  \19 ,
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ;
output
  \98 ;
reg
  \2 ,
  \36 ,
  \37 ,
  \38 ,
  \39 ,
  \40 ,
  \41 ,
  \42 ,
  \43 ,
  \44 ,
  \45 ,
  \46 ,
  \47 ,
  \48 ,
  \49 ,
  \50 ,
  \51 ,
  \52 ,
  \53 ,
  \54 ,
  \55 ,
  \56 ,
  \57 ,
  \58 ,
  \59 ,
  \60 ,
  \61 ,
  \62 ,
  \63 ,
  \64 ,
  \65 ,
  \66 ,
  \67 ,
  \68 ,
  \69 ,
  \70 ,
  \71 ,
  \72 ,
  \73 ,
  \74 ,
  \75 ,
  \76 ,
  \77 ,
  \78 ,
  \79 ,
  \80 ,
  \81 ,
  \82 ,
  \83 ,
  \84 ,
  \85 ,
  \86 ,
  \87 ,
  \88 ,
  \89 ,
  \90 ,
  \91 ,
  \92 ,
  \93 ,
  \94 ,
  \95 ;
wire
  \370 ,
  \371 ,
  \372 ,
  \373 ,
  \374 ,
  \375 ,
  \376 ,
  \377 ,
  \383 ,
  \384 ,
  \386 ,
  \387 ,
  \389 ,
  \390 ,
  \392 ,
  \393 ,
  \395 ,
  \396 ,
  \398 ,
  \399 ,
  \[64] ,
  \[65] ,
  \[66] ,
  \[67] ,
  \[68] ,
  \[69] ,
  \401 ,
  \402 ,
  \404 ,
  \405 ,
  \407 ,
  \408 ,
  \410 ,
  \411 ,
  \413 ,
  \414 ,
  \416 ,
  \417 ,
  \419 ,
  \420 ,
  \422 ,
  \423 ,
  \425 ,
  \426 ,
  \428 ,
  \429 ,
  \431 ,
  \432 ,
  \434 ,
  \435 ,
  \437 ,
  \438 ,
  \440 ,
  \441 ,
  \443 ,
  \444 ,
  \446 ,
  \447 ,
  \449 ,
  \450 ,
  \452 ,
  \453 ,
  \455 ,
  \456 ,
  \458 ,
  \459 ,
  \461 ,
  \462 ,
  \464 ,
  \465 ,
  \467 ,
  \468 ,
  \[70] ,
  \470 ,
  \471 ,
  \477 ,
  \479 ,
  \[71] ,
  \481 ,
  \483 ,
  \485 ,
  \487 ,
  \489 ,
  \[72] ,
  \491 ,
  \493 ,
  \495 ,
  \497 ,
  \499 ,
  \[73] ,
  \[74] ,
  \[75] ,
  \[76] ,
  \[77] ,
  \[78] ,
  \[79] ,
  \501 ,
  \503 ,
  \505 ,
  \507 ,
  \509 ,
  \511 ,
  \513 ,
  \515 ,
  \517 ,
  \519 ,
  \521 ,
  \523 ,
  \525 ,
  \527 ,
  \529 ,
  \531 ,
  \533 ,
  \535 ,
  \537 ,
  \[80] ,
  \[81] ,
  \[82] ,
  \[83] ,
  \[84] ,
  \[85] ,
  \[86] ,
  \[87] ,
  \[88] ,
  \[89] ,
  \[90] ,
  \[91] ,
  \[92] ,
  \[93] ,
  \[94] ,
  \[95] ,
  \[96] ,
  \[97] ,
  \[98] ,
  \[100] ,
  \[99] ,
  \[101] ,
  \[102] ,
  \[103] ,
  \[104] ,
  \[105] ,
  \[106] ,
  \[107] ,
  \[108] ,
  \[109] ,
  \[110] ,
  \[111] ,
  \[112] ,
  \[113] ,
  \[114] ,
  \[115] ,
  \[116] ,
  \[117] ,
  \[118] ,
  \[119] ,
  \[120] ,
  \[121] ,
  \[122] ,
  \[123] ,
  \[124] ,
  \226 ,
  \227 ,
  \228 ,
  \229 ,
  \230 ,
  \231 ,
  \232 ,
  \233 ,
  \234 ,
  \235 ,
  \236 ,
  \237 ,
  \238 ,
  \239 ,
  \240 ,
  \241 ,
  \242 ,
  \243 ,
  \244 ,
  \245 ,
  \246 ,
  \247 ,
  \248 ,
  \249 ,
  \250 ,
  \251 ,
  \252 ,
  \253 ,
  \254 ,
  \255 ,
  \256 ,
  \257 ,
  \258 ,
  \259 ,
  \260 ,
  \261 ,
  \262 ,
  \263 ,
  \264 ,
  \265 ,
  \266 ,
  \267 ,
  \268 ,
  \269 ,
  \270 ,
  \271 ,
  \272 ,
  \273 ,
  \274 ,
  \275 ,
  \276 ,
  \277 ,
  \278 ,
  \279 ,
  \280 ,
  \281 ,
  \282 ,
  \283 ,
  \284 ,
  \285 ,
  \286 ,
  \287 ,
  \288 ,
  \289 ,
  \290 ,
  \291 ,
  \292 ,
  \293 ,
  \294 ,
  \295 ,
  \296 ,
  \297 ,
  \298 ,
  \299 ,
  \300 ,
  \301 ,
  \302 ,
  \303 ,
  \304 ,
  \305 ,
  \306 ,
  \307 ,
  \308 ,
  \309 ,
  \310 ,
  \311 ,
  \312 ,
  \313 ,
  \314 ,
  \315 ,
  \316 ,
  \317 ,
  \318 ,
  \319 ,
  \320 ,
  \321 ,
  \322 ,
  \323 ,
  \324 ,
  \325 ,
  \326 ,
  \327 ,
  \328 ,
  \329 ,
  \330 ,
  \331 ,
  \332 ,
  \333 ,
  \334 ,
  \335 ,
  \336 ,
  \337 ,
  \338 ,
  \339 ,
  \340 ,
  \341 ,
  \342 ,
  \343 ,
  \344 ,
  \345 ,
  \346 ,
  \347 ,
  \348 ,
  \349 ,
  \350 ,
  \351 ,
  \352 ,
  \353 ,
  \354 ,
  \355 ,
  \356 ,
  \357 ,
  \358 ,
  \359 ,
  \360 ,
  \361 ,
  \362 ,
  \363 ,
  \364 ,
  \365 ,
  \366 ,
  \367 ,
  \368 ,
  \369 ;
assign
  \370  = \468  | \369 ,
  \371  = (~\479  & \470 ) | (\479  & ~\470 ),
  \372  = \479  & \65 ,
  \373  = \479  & \95 ,
  \374  = \65  & \95 ,
  \375  = \471  | \374 ,
  \376  = (~\477  & \2 ) | (\477  & ~\2 ),
  \377  = \477  & \2 ,
  \383  = (~\36  & \66 ) | (\36  & ~\66 ),
  \384  = \228  | \227 ,
  \386  = (~\37  & \67 ) | (\37  & ~\67 ),
  \387  = \233  | \232 ,
  \389  = (~\38  & \68 ) | (\38  & ~\68 ),
  \390  = \238  | \237 ,
  \392  = (~\39  & \69 ) | (\39  & ~\69 ),
  \393  = \243  | \242 ,
  \395  = (~\40  & \70 ) | (\40  & ~\70 ),
  \396  = \248  | \247 ,
  \398  = (~\41  & \71 ) | (\41  & ~\71 ),
  \399  = \253  | \252 ,
  \[64]  = \231 ,
  \[65]  = \236 ,
  \[66]  = \241 ,
  \[67]  = \246 ,
  \[68]  = \251 ,
  \[69]  = \256 ,
  \401  = (~\42  & \72 ) | (\42  & ~\72 ),
  \402  = \258  | \257 ,
  \404  = (~\43  & \73 ) | (\43  & ~\73 ),
  \405  = \263  | \262 ,
  \407  = (~\44  & \74 ) | (\44  & ~\74 ),
  \408  = \268  | \267 ,
  \410  = (~\45  & \75 ) | (\45  & ~\75 ),
  \411  = \273  | \272 ,
  \413  = (~\46  & \76 ) | (\46  & ~\76 ),
  \414  = \278  | \277 ,
  \416  = (~\47  & \77 ) | (\47  & ~\77 ),
  \417  = \283  | \282 ,
  \419  = (~\48  & \78 ) | (\48  & ~\78 ),
  \420  = \288  | \287 ,
  \422  = (~\49  & \79 ) | (\49  & ~\79 ),
  \423  = \293  | \292 ,
  \425  = (~\50  & \80 ) | (\50  & ~\80 ),
  \426  = \298  | \297 ,
  \428  = (~\51  & \81 ) | (\51  & ~\81 ),
  \429  = \303  | \302 ,
  \431  = (~\52  & \82 ) | (\52  & ~\82 ),
  \432  = \308  | \307 ,
  \434  = (~\53  & \83 ) | (\53  & ~\83 ),
  \435  = \313  | \312 ,
  \437  = (~\54  & \84 ) | (\54  & ~\84 ),
  \438  = \318  | \317 ,
  \440  = (~\55  & \85 ) | (\55  & ~\85 ),
  \441  = \323  | \322 ,
  \443  = (~\56  & \86 ) | (\56  & ~\86 ),
  \444  = \328  | \327 ,
  \446  = (~\57  & \87 ) | (\57  & ~\87 ),
  \447  = \333  | \332 ,
  \449  = (~\58  & \88 ) | (\58  & ~\88 ),
  \450  = \338  | \337 ,
  \452  = (~\59  & \89 ) | (\59  & ~\89 ),
  \453  = \343  | \342 ,
  \455  = (~\60  & \90 ) | (\60  & ~\90 ),
  \456  = \348  | \347 ,
  \458  = (~\61  & \91 ) | (\61  & ~\91 ),
  \459  = \353  | \352 ,
  \461  = (~\62  & \92 ) | (\62  & ~\92 ),
  \462  = \358  | \357 ,
  \464  = (~\63  & \93 ) | (\63  & ~\93 ),
  \465  = \363  | \362 ,
  \467  = (~\64  & \94 ) | (\64  & ~\94 ),
  \468  = \368  | \367 ,
  \[70]  = \261 ,
  \470  = (~\65  & \95 ) | (\65  & ~\95 ),
  \471  = \373  | \372 ,
  \477  = \33  & \1 ,
  \479  = \32  & \1 ,
  \[71]  = \266 ,
  \481  = \31  & \1 ,
  \483  = \30  & \1 ,
  \485  = \29  & \1 ,
  \487  = \28  & \1 ,
  \489  = \27  & \1 ,
  \[72]  = \271 ,
  \491  = \26  & \1 ,
  \493  = \25  & \1 ,
  \495  = \24  & \1 ,
  \497  = \23  & \1 ,
  \499  = \22  & \1 ,
  \[73]  = \276 ,
  \[74]  = \281 ,
  \[75]  = \286 ,
  \[76]  = \291 ,
  \[77]  = \296 ,
  \[78]  = \301 ,
  \[79]  = \306 ,
  \501  = \21  & \1 ,
  \503  = \20  & \1 ,
  \505  = \19  & \1 ,
  \507  = \18  & \1 ,
  \509  = \17  & \1 ,
  \511  = \16  & \1 ,
  \513  = \15  & \1 ,
  \515  = \14  & \1 ,
  \517  = \13  & \1 ,
  \519  = \12  & \1 ,
  \521  = \11  & \1 ,
  \523  = \10  & \1 ,
  \525  = \9  & \1 ,
  \527  = \8  & \1 ,
  \529  = \7  & \1 ,
  \531  = \6  & \1 ,
  \533  = \5  & \1 ,
  \535  = \4  & \1 ,
  \537  = \3  & \1 ,
  \[80]  = \311 ,
  \[81]  = \316 ,
  \[82]  = \321 ,
  \[83]  = \326 ,
  \[84]  = \331 ,
  \[85]  = \336 ,
  \[86]  = \341 ,
  \[87]  = \346 ,
  \[88]  = \351 ,
  \[89]  = \356 ,
  \[90]  = \361 ,
  \[91]  = \366 ,
  \[92]  = \371 ,
  \[93]  = \376 ,
  \[94]  = \230 ,
  \[95]  = \235 ,
  \[96]  = \240 ,
  \[97]  = \245 ,
  \[98]  = \250 ,
  \[100]  = \260 ,
  \[99]  = \255 ,
  \[101]  = \265 ,
  \[102]  = \270 ,
  \[103]  = \275 ,
  \98  = \226 ,
  \[104]  = \280 ,
  \[105]  = \285 ,
  \[106]  = \290 ,
  \[107]  = \295 ,
  \[108]  = \300 ,
  \[109]  = \305 ,
  \[110]  = \310 ,
  \[111]  = \315 ,
  \[112]  = \320 ,
  \[113]  = \325 ,
  \[114]  = \330 ,
  \[115]  = \335 ,
  \[116]  = \340 ,
  \[117]  = \345 ,
  \[118]  = \350 ,
  \[119]  = \355 ,
  \[120]  = \360 ,
  \[121]  = \365 ,
  \[122]  = \370 ,
  \[123]  = \375 ,
  \[124]  = \377 ,
  \226  = (~\537  & \383 ) | (\537  & ~\383 ),
  \227  = \537  & \36 ,
  \228  = \537  & \66 ,
  \229  = \36  & \66 ,
  \230  = \384  | \229 ,
  \231  = (~\535  & \386 ) | (\535  & ~\386 ),
  \232  = \535  & \37 ,
  \233  = \535  & \67 ,
  \234  = \37  & \67 ,
  \235  = \387  | \234 ,
  \236  = (~\533  & \389 ) | (\533  & ~\389 ),
  \237  = \533  & \38 ,
  \238  = \533  & \68 ,
  \239  = \38  & \68 ,
  \240  = \390  | \239 ,
  \241  = (~\531  & \392 ) | (\531  & ~\392 ),
  \242  = \531  & \39 ,
  \243  = \531  & \69 ,
  \244  = \39  & \69 ,
  \245  = \393  | \244 ,
  \246  = (~\529  & \395 ) | (\529  & ~\395 ),
  \247  = \529  & \40 ,
  \248  = \529  & \70 ,
  \249  = \40  & \70 ,
  \250  = \396  | \249 ,
  \251  = (~\527  & \398 ) | (\527  & ~\398 ),
  \252  = \527  & \41 ,
  \253  = \527  & \71 ,
  \254  = \41  & \71 ,
  \255  = \399  | \254 ,
  \256  = (~\525  & \401 ) | (\525  & ~\401 ),
  \257  = \525  & \42 ,
  \258  = \525  & \72 ,
  \259  = \42  & \72 ,
  \260  = \402  | \259 ,
  \261  = (~\523  & \404 ) | (\523  & ~\404 ),
  \262  = \523  & \43 ,
  \263  = \523  & \73 ,
  \264  = \43  & \73 ,
  \265  = \405  | \264 ,
  \266  = (~\521  & \407 ) | (\521  & ~\407 ),
  \267  = \521  & \44 ,
  \268  = \521  & \74 ,
  \269  = \44  & \74 ,
  \270  = \408  | \269 ,
  \271  = (~\519  & \410 ) | (\519  & ~\410 ),
  \272  = \519  & \45 ,
  \273  = \519  & \75 ,
  \274  = \45  & \75 ,
  \275  = \411  | \274 ,
  \276  = (~\517  & \413 ) | (\517  & ~\413 ),
  \277  = \517  & \46 ,
  \278  = \517  & \76 ,
  \279  = \46  & \76 ,
  \280  = \414  | \279 ,
  \281  = (~\515  & \416 ) | (\515  & ~\416 ),
  \282  = \515  & \47 ,
  \283  = \515  & \77 ,
  \284  = \47  & \77 ,
  \285  = \417  | \284 ,
  \286  = (~\513  & \419 ) | (\513  & ~\419 ),
  \287  = \513  & \48 ,
  \288  = \513  & \78 ,
  \289  = \48  & \78 ,
  \290  = \420  | \289 ,
  \291  = (~\511  & \422 ) | (\511  & ~\422 ),
  \292  = \511  & \49 ,
  \293  = \511  & \79 ,
  \294  = \49  & \79 ,
  \295  = \423  | \294 ,
  \296  = (~\509  & \425 ) | (\509  & ~\425 ),
  \297  = \509  & \50 ,
  \298  = \509  & \80 ,
  \299  = \50  & \80 ,
  \300  = \426  | \299 ,
  \301  = (~\507  & \428 ) | (\507  & ~\428 ),
  \302  = \507  & \51 ,
  \303  = \507  & \81 ,
  \304  = \51  & \81 ,
  \305  = \429  | \304 ,
  \306  = (~\505  & \431 ) | (\505  & ~\431 ),
  \307  = \505  & \52 ,
  \308  = \505  & \82 ,
  \309  = \52  & \82 ,
  \310  = \432  | \309 ,
  \311  = (~\503  & \434 ) | (\503  & ~\434 ),
  \312  = \503  & \53 ,
  \313  = \503  & \83 ,
  \314  = \53  & \83 ,
  \315  = \435  | \314 ,
  \316  = (~\501  & \437 ) | (\501  & ~\437 ),
  \317  = \501  & \54 ,
  \318  = \501  & \84 ,
  \319  = \54  & \84 ,
  \320  = \438  | \319 ,
  \321  = (~\499  & \440 ) | (\499  & ~\440 ),
  \322  = \499  & \55 ,
  \323  = \499  & \85 ,
  \324  = \55  & \85 ,
  \325  = \441  | \324 ,
  \326  = (~\497  & \443 ) | (\497  & ~\443 ),
  \327  = \497  & \56 ,
  \328  = \497  & \86 ,
  \329  = \56  & \86 ,
  \330  = \444  | \329 ,
  \331  = (~\495  & \446 ) | (\495  & ~\446 ),
  \332  = \495  & \57 ,
  \333  = \495  & \87 ,
  \334  = \57  & \87 ,
  \335  = \447  | \334 ,
  \336  = (~\493  & \449 ) | (\493  & ~\449 ),
  \337  = \493  & \58 ,
  \338  = \493  & \88 ,
  \339  = \58  & \88 ,
  \340  = \450  | \339 ,
  \341  = (~\491  & \452 ) | (\491  & ~\452 ),
  \342  = \491  & \59 ,
  \343  = \491  & \89 ,
  \344  = \59  & \89 ,
  \345  = \453  | \344 ,
  \346  = (~\489  & \455 ) | (\489  & ~\455 ),
  \347  = \489  & \60 ,
  \348  = \489  & \90 ,
  \349  = \60  & \90 ,
  \350  = \456  | \349 ,
  \351  = (~\487  & \458 ) | (\487  & ~\458 ),
  \352  = \487  & \61 ,
  \353  = \487  & \91 ,
  \354  = \61  & \91 ,
  \355  = \459  | \354 ,
  \356  = (~\485  & \461 ) | (\485  & ~\461 ),
  \357  = \485  & \62 ,
  \358  = \485  & \92 ,
  \359  = \62  & \92 ,
  \360  = \462  | \359 ,
  \361  = (~\483  & \464 ) | (\483  & ~\464 ),
  \362  = \483  & \63 ,
  \363  = \483  & \93 ,
  \364  = \63  & \93 ,
  \365  = \465  | \364 ,
  \366  = (~\481  & \467 ) | (\481  & ~\467 ),
  \367  = \481  & \64 ,
  \368  = \481  & \94 ,
  \369  = \64  & \94 ;
always begin
  \2  = \[64] ;
  \36  = \[65] ;
  \37  = \[66] ;
  \38  = \[67] ;
  \39  = \[68] ;
  \40  = \[69] ;
  \41  = \[70] ;
  \42  = \[71] ;
  \43  = \[72] ;
  \44  = \[73] ;
  \45  = \[74] ;
  \46  = \[75] ;
  \47  = \[76] ;
  \48  = \[77] ;
  \49  = \[78] ;
  \50  = \[79] ;
  \51  = \[80] ;
  \52  = \[81] ;
  \53  = \[82] ;
  \54  = \[83] ;
  \55  = \[84] ;
  \56  = \[85] ;
  \57  = \[86] ;
  \58  = \[87] ;
  \59  = \[88] ;
  \60  = \[89] ;
  \61  = \[90] ;
  \62  = \[91] ;
  \63  = \[92] ;
  \64  = \[93] ;
  \65  = \[94] ;
  \66  = \[95] ;
  \67  = \[96] ;
  \68  = \[97] ;
  \69  = \[98] ;
  \70  = \[99] ;
  \71  = \[100] ;
  \72  = \[101] ;
  \73  = \[102] ;
  \74  = \[103] ;
  \75  = \[104] ;
  \76  = \[105] ;
  \77  = \[106] ;
  \78  = \[107] ;
  \79  = \[108] ;
  \80  = \[109] ;
  \81  = \[110] ;
  \82  = \[111] ;
  \83  = \[112] ;
  \84  = \[113] ;
  \85  = \[114] ;
  \86  = \[115] ;
  \87  = \[116] ;
  \88  = \[117] ;
  \89  = \[118] ;
  \90  = \[119] ;
  \91  = \[120] ;
  \92  = \[121] ;
  \93  = \[122] ;
  \94  = \[123] ;
  \95  = \[124] ;
end
initial begin
  \2  = 0;
  \36  = 0;
  \37  = 0;
  \38  = 0;
  \39  = 0;
  \40  = 0;
  \41  = 0;
  \42  = 0;
  \43  = 0;
  \44  = 0;
  \45  = 0;
  \46  = 0;
  \47  = 0;
  \48  = 0;
  \49  = 0;
  \50  = 0;
  \51  = 0;
  \52  = 0;
  \53  = 0;
  \54  = 0;
  \55  = 0;
  \56  = 0;
  \57  = 0;
  \58  = 0;
  \59  = 0;
  \60  = 0;
  \61  = 0;
  \62  = 0;
  \63  = 0;
  \64  = 0;
  \65  = 0;
  \66  = 0;
  \67  = 0;
  \68  = 0;
  \69  = 0;
  \70  = 0;
  \71  = 0;
  \72  = 0;
  \73  = 0;
  \74  = 0;
  \75  = 0;
  \76  = 0;
  \77  = 0;
  \78  = 0;
  \79  = 0;
  \80  = 0;
  \81  = 0;
  \82  = 0;
  \83  = 0;
  \84  = 0;
  \85  = 0;
  \86  = 0;
  \87  = 0;
  \88  = 0;
  \89  = 0;
  \90  = 0;
  \91  = 0;
  \92  = 0;
  \93  = 0;
  \94  = 0;
  \95  = 0;
end
endmodule

