//NOTE: no-implementation module stub

module REG12LC (
    input wire DSPCLK,
    input wire MMR_web,
    input wire AUTO_we,
    input wire [11:0] DMD,
    output reg [11:0] AUTO_b,
    input wire RST
);

endmodule
