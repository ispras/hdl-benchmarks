module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
 n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
 n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
 n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
 n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
 n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , 
 n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , 
 n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , 
 n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , 
 n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , 
 n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , 
 n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , 
 n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , 
 n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , 
 n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , 
 n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , 
 n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , 
 n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , 
 n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , 
 n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , 
 n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , 
 n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , 
 n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , 
 n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , 
 n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , 
 n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , 
 n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , 
 n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , 
 n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , 
 n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , 
 n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , 
 n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , 
 n541 , n542 , n543 , n544 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 ;
output n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
 n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
 n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
 n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
 n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
 n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , 
 n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , 
 n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , 
 n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , 
 n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , 
 n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , 
 n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , 
 n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , 
 n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , 
 n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , 
 n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , 
 n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , 
 n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , 
 n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , 
 n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , 
 n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , 
 n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , 
 n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , 
 n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , 
 n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , 
 n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , 
 n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , 
 n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , 
 n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , 
 n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , 
 n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , 
 n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , 
 n541 , n542 , n543 , n544 ;
wire n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , 
 n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , 
 n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , 
 n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , 
 n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , 
 n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , 
 n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , 
 n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , 
 n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , 
 n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , 
 n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , 
 n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , 
 n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , 
 n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , 
 n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , 
 n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , 
 n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , 
 n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , 
 n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , 
 n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , 
 n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , 
 n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , 
 n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , 
 n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , 
 n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , 
 n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , 
 n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , 
 n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , 
 n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , 
 n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , 
 n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , 
 n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , 
 n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , 
 n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , 
 n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , 
 n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , 
 n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , 
 n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , 
 n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , 
 n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , 
 n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , 
 n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , 
 n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , 
 n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , 
 n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , 
 n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , 
 n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , 
 n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , 
 n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , 
 n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , 
 n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , 
 n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , 
 n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , 
 n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , 
 n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , 
 n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , 
 n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , 
 n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , 
 n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , 
 n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , 
 n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , 
 n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , 
 n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , 
 n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , 
 n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , 
 n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , 
 n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , 
 n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , 
 n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , 
 n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , 
 n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , 
 n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , 
 n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , 
 n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , 
 n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , 
 n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , 
 n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , 
 n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , 
 n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , 
 n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , 
 n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , 
 n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , 
 n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , 
 n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , 
 n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , 
 n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , 
 n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , 
 n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , 
 n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , 
 n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , 
 n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , 
 n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , 
 n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , 
 n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , 
 n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , 
 n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , 
 n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , 
 n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , 
 n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , 
 n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , 
 n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , 
 n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , 
 n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , 
 n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , 
 n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , 
 n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , 
 n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , 
 n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , 
 n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , 
 n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , 
 n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , 
 n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , 
 n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , 
 n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , 
 n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , 
 n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , 
 n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , 
 n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , 
 n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , 
 n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , 
 n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , 
 n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , 
 n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , 
 n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , 
 n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , 
 n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , 
 n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , 
 n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , 
 n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , 
 n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , 
 n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , 
 n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , 
 n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , 
 n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , 
 n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , 
 n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , 
 n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , 
 n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , 
 n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , 
 n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , 
 n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , 
 n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , 
 n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , 
 n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , 
 n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , 
 n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , 
 n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , 
 n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , 
 n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , 
 n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , 
 n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , 
 n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , 
 n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , 
 n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , 
 n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , 
 n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , 
 n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , 
 n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , 
 n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , 
 n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , 
 n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , 
 n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , 
 n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , 
 n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , 
 n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , 
 n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , 
 n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , 
 n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , 
 n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , 
 n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , 
 n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , 
 n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , 
 n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , 
 n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , 
 n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , 
 n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , 
 n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , 
 n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , 
 n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , 
 n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , 
 n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , 
 n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , 
 n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , 
 n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , 
 n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , 
 n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , 
 n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , 
 n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , 
 n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , 
 n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , 
 n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , 
 n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , 
 n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , 
 n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , 
 n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , 
 n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , 
 n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , 
 n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , 
 n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , 
 n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , 
 n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , 
 n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , 
 n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , 
 n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , 
 n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , 
 n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , 
 n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , 
 n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , 
 n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , 
 n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , 
 n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , 
 n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , 
 n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , 
 n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , 
 n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , 
 n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , 
 n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , 
 n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , 
 n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , 
 n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , 
 n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , 
 n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , 
 n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , 
 n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , 
 n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , 
 n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , 
 n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , 
 n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , 
 n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , 
 n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , 
 n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , 
 n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , 
 n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , 
 n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , 
 n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , 
 n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , 
 n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , 
 n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , 
 n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , 
 n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , 
 n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , 
 n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , 
 n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , 
 n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , 
 n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , 
 n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , 
 n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , 
 n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , 
 n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , 
 n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , 
 n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , 
 n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , 
 n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , 
 n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , 
 n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , 
 n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , 
 n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , 
 n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , 
 n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , 
 n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , 
 n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , 
 n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , 
 n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , 
 n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , 
 n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , 
 n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , 
 n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , 
 n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , 
 n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , 
 n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , 
 n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , 
 n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , 
 n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , 
 n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , 
 n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , 
 n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , 
 n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , 
 n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , 
 n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , 
 n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , 
 n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , 
 n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , 
 n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , 
 n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , 
 n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , 
 n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , 
 n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , 
 n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , 
 n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , 
 n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , 
 n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , 
 n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , 
 n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , 
 n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , 
 n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , 
 n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , 
 n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , 
 n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , 
 n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , 
 n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , 
 n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , 
 n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , 
 n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , 
 n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , 
 n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , 
 n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , 
 n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , 
 n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , 
 n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , 
 n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , 
 n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , 
 n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , 
 n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , 
 n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , 
 n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , 
 n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , 
 n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , 
 n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , 
 n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , 
 n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , 
 n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , 
 n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , 
 n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , 
 n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , 
 n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , 
 n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , 
 n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , 
 n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , 
 n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , 
 n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , 
 n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , 
 n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , 
 n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , 
 n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , 
 n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , 
 n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , 
 n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , 
 n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , 
 n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , 
 n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , 
 n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , 
 n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , 
 n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , 
 n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , 
 n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , 
 n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , 
 n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , 
 n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , 
 n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , 
 n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , 
 n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , 
 n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , 
 n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , 
 n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , 
 n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , 
 n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , 
 n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , 
 n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , 
 n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , 
 n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , 
 n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , 
 n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , 
 n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , 
 n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , 
 n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , 
 n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , 
 n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , 
 n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , 
 n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , 
 n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , 
 n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , 
 n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , 
 n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , 
 n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , 
 n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , 
 n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , 
 n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , 
 n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , 
 n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , 
 n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , 
 n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , 
 n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , 
 n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , 
 n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , 
 n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , 
 n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , 
 n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , 
 n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , 
 n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , 
 n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , 
 n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , 
 n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , 
 n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , 
 n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , 
 n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , 
 n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , 
 n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , 
 n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , 
 n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , 
 n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , 
 n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , 
 n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , 
 n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , 
 n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , 
 n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , 
 n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , 
 n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , 
 n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , 
 n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , 
 n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , 
 n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , 
 n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , 
 n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , 
 n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , 
 n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , 
 n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , 
 n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , 
 n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , 
 n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , 
 n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , 
 n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , 
 n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , 
 n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , 
 n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , 
 n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , 
 n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , 
 n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , 
 n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , 
 n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , 
 n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , 
 n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , 
 n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , 
 n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , 
 n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , 
 n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , 
 n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , 
 n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , 
 n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , 
 n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , 
 n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , 
 n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , 
 n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , 
 n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , 
 n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , 
 n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , 
 n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , 
 n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , 
 n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , 
 n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , 
 n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , 
 n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , 
 n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , 
 n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , 
 n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , 
 n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , 
 n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , 
 n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , 
 n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , 
 n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , 
 n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , 
 n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , 
 n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , 
 n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , 
 n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , 
 n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , 
 n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , 
 n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , 
 n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , 
 n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , 
 n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , 
 n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , 
 n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , 
 n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , 
 n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , 
 n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , 
 n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , 
 n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , 
 n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , 
 n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , 
 n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , 
 n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , 
 n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , 
 n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , 
 n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , 
 n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , 
 n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , 
 n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , 
 n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , 
 n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , 
 n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , 
 n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , 
 n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , 
 n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , 
 n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , 
 n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , 
 n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , 
 n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , 
 n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , 
 n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , 
 n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , 
 n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , 
 n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , 
 n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , 
 n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , 
 n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , 
 n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , 
 n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , 
 n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , 
 n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , 
 n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , 
 n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , 
 n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , 
 n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , 
 n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , 
 n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , 
 n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , 
 n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , 
 n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , 
 n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , 
 n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , 
 n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , 
 n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , 
 n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , 
 n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , 
 n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , 
 n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , 
 n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , 
 n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , 
 n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , 
 n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , 
 n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , 
 n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , 
 n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , 
 n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , 
 n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , 
 n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , 
 n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , 
 n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , 
 n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , 
 n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , 
 n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , 
 n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , 
 n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , 
 n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , 
 n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , 
 n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , 
 n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , 
 n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , 
 n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , 
 n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , 
 n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , 
 n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , 
 n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , 
 n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , 
 n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , 
 n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , 
 n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , 
 n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , 
 n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , 
 n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , 
 n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , 
 n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , 
 n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , 
 n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , 
 n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , 
 n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , 
 n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , 
 n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , 
 n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , 
 n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , 
 n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , 
 n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , 
 n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , 
 n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , 
 n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , 
 n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , 
 n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , 
 n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , 
 n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , 
 n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , 
 n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , 
 n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , 
 n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , 
 n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , 
 n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , 
 n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , 
 n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , 
 n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , 
 n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , 
 n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , 
 n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , 
 n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , 
 n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , 
 n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , 
 n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , 
 n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , 
 n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , 
 n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , 
 n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , 
 n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , 
 n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , 
 n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , 
 n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , 
 n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , 
 n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , 
 n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , 
 n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , 
 n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , 
 n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , 
 n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , 
 n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , 
 n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , 
 n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , 
 n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , 
 n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , 
 n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , 
 n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , 
 n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , 
 n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , 
 n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , 
 n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , 
 n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , 
 n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , 
 n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , 
 n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , 
 n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , 
 n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , 
 n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , 
 n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , 
 n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , 
 n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , 
 n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , 
 n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , 
 n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , 
 n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , 
 n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , 
 n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , 
 n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , 
 n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , 
 n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , 
 n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , 
 n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , 
 n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , 
 n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , 
 n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , 
 n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , 
 n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , 
 n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , 
 n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , 
 n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , 
 n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , 
 n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , 
 n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , 
 n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , 
 n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , 
 n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , 
 n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , 
 n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , 
 n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , 
 n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , 
 n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , 
 n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , 
 n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , 
 n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , 
 n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , 
 n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , 
 n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , 
 n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , 
 n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , 
 n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , 
 n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , 
 n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , 
 n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , 
 n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , 
 n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , 
 n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , 
 n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , 
 n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , 
 n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , 
 n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , 
 n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , 
 n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , 
 n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , 
 n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , 
 n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , 
 n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , 
 n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , 
 n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , 
 n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , 
 n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , 
 n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , 
 n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , 
 n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , 
 n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , 
 n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , 
 n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , 
 n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , 
 n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , 
 n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , 
 n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , 
 n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , 
 n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , 
 n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , 
 n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , 
 n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , 
 n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , 
 n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , 
 n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , 
 n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , 
 n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , 
 n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , 
 n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , 
 n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , 
 n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , 
 n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , 
 n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , 
 n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , 
 n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , 
 n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , 
 n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , 
 n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , 
 n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , 
 n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , 
 n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , 
 n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , 
 n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , 
 n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , 
 n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , 
 n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , 
 n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , 
 n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , 
 n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , 
 n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , 
 n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , 
 n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , 
 n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , 
 n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , 
 n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , 
 n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , 
 n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , 
 n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , 
 n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , 
 n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , 
 n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , 
 n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , 
 n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , 
 n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , 
 n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , 
 n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , 
 n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , 
 n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , 
 n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , 
 n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , 
 n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , 
 n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , 
 n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , 
 n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , 
 n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , 
 n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , 
 n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , 
 n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , 
 n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , 
 n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , 
 n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , 
 n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , 
 n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , 
 n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , 
 n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , 
 n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , 
 n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , 
 n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , 
 n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , 
 n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , 
 n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , 
 n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , 
 n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , 
 n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , 
 n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , 
 n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , 
 n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , 
 n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , 
 n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , 
 n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , 
 n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , 
 n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , 
 n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , 
 n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , 
 n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , 
 n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , 
 n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , 
 n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , 
 n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , 
 n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , 
 n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , 
 n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , 
 n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , 
 n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , 
 n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , 
 n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , 
 n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , 
 n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , 
 n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , 
 n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , 
 n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , 
 n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , 
 n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , 
 n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , 
 n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , 
 n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , 
 n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , 
 n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , 
 n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , 
 n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , 
 n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , 
 n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , 
 n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , 
 n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , 
 n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , 
 n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , 
 n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , 
 n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , 
 n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , 
 n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , 
 n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , 
 n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , 
 n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , 
 n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , 
 n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , 
 n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , 
 n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , 
 n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , 
 n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , 
 n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , 
 n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , 
 n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , 
 n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , 
 n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , 
 n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , 
 n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , 
 n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , 
 n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , 
 n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , 
 n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , 
 n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , 
 n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , 
 n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , 
 n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , 
 n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , 
 n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , 
 n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , 
 n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , 
 n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , 
 n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , 
 n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , 
 n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , 
 n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , 
 n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , 
 n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , 
 n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , 
 n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , 
 n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , 
 n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , 
 n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , 
 n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , 
 n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , 
 n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , 
 n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , 
 n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , 
 n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , 
 n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , 
 n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , 
 n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , 
 n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , 
 n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , 
 n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , 
 n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , 
 n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , 
 n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , 
 n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , 
 n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , 
 n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , 
 n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , 
 n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , 
 n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , 
 n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , 
 n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , 
 n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , 
 n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , 
 n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , 
 n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , 
 n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , 
 n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , 
 n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , 
 n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , 
 n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , 
 n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , 
 n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , 
 n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , 
 n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , 
 n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , 
 n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , 
 n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , 
 n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , 
 n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , 
 n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , 
 n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , 
 n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , 
 n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , 
 n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , 
 n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , 
 n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , 
 n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , 
 n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , 
 n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , 
 n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , 
 n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , 
 n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , 
 n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , 
 n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , 
 n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , 
 n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , 
 n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , 
 n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , 
 n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , 
 n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , 
 n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , 
 n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , 
 n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , 
 n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , 
 n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , 
 n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , 
 n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , 
 n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , 
 n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , 
 n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , 
 n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , 
 n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , 
 n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , 
 n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , 
 n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , 
 n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , 
 n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , 
 n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , 
 n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , 
 n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , 
 n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , 
 n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , 
 n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , 
 n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , 
 n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , 
 n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , 
 n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , 
 n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , 
 n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , 
 n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , 
 n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , 
 n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , 
 n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , 
 n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , 
 n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , 
 n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , 
 n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , 
 n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , 
 n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , 
 n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , 
 n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , 
 n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , 
 n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , 
 n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , 
 n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , 
 n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , 
 n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , 
 n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , 
 n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , 
 n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , 
 n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , 
 n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , 
 n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , 
 n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , 
 n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , 
 n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , 
 n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , 
 n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , 
 n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , 
 n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , 
 n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , 
 n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , 
 n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , 
 n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , 
 n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , 
 n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , 
 n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , 
 n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , 
 n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , 
 n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , 
 n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , 
 n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , 
 n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , 
 n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , 
 n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , 
 n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , 
 n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , 
 n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , 
 n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , 
 n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , 
 n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , 
 n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , 
 n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , 
 n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , 
 n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , 
 n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , 
 n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , 
 n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , 
 n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , 
 n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , 
 n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , 
 n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , 
 n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , 
 n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , 
 n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , 
 n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , 
 n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , 
 n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , 
 n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , 
 n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , 
 n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , 
 n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , 
 n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , 
 n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , 
 n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , 
 n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , 
 n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , 
 n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , 
 n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , 
 n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , 
 n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , 
 n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , 
 n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , 
 n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , 
 n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , 
 n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , 
 n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , 
 n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , 
 n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , 
 n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , 
 n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , 
 n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , 
 n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , 
 n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , 
 n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , 
 n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , 
 n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , 
 n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , 
 n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , 
 n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , 
 n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , 
 n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , 
 n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , 
 n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , 
 n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , 
 n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , 
 n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , 
 n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , 
 n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , 
 n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , 
 n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , 
 n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , 
 n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , 
 n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , 
 n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , 
 n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , 
 n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , 
 n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , 
 n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , 
 n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , 
 n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , 
 n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , 
 n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , 
 n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , 
 n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , 
 n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , 
 n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , 
 n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , 
 n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , 
 n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , 
 n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , 
 n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , 
 n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , 
 n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , 
 n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , 
 n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , 
 n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , 
 n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , 
 n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , 
 n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , 
 n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , 
 n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , 
 n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , 
 n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , 
 n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , 
 n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , 
 n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , 
 n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , 
 n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , 
 n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , 
 n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , 
 n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , 
 n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , 
 n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , 
 n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , 
 n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , 
 n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , 
 n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , 
 n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , 
 n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , 
 n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , 
 n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , 
 n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , 
 n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , 
 n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , 
 n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , 
 n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , 
 n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , 
 n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , 
 n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , 
 n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , 
 n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , 
 n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , 
 n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , 
 n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , 
 n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , 
 n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , 
 n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , 
 n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , 
 n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , 
 n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , 
 n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , 
 n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , 
 n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , 
 n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , 
 n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , 
 n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , 
 n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , 
 n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , 
 n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , 
 n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , 
 n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , 
 n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , 
 n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , 
 n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , 
 n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , 
 n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , 
 n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , 
 n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , 
 n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , 
 n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , 
 n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , 
 n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , 
 n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , 
 n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , 
 n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , 
 n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , 
 n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , 
 n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , 
 n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , 
 n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , 
 n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , 
 n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , 
 n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , 
 n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , 
 n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , 
 n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , 
 n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , 
 n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , 
 n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , 
 n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , 
 n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , 
 n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , 
 n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , 
 n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , 
 n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , 
 n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , 
 n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , 
 n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , 
 n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , 
 n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , 
 n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , 
 n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , 
 n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , 
 n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , 
 n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , 
 n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , 
 n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , 
 n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , 
 n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , 
 n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , 
 n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , 
 n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , 
 n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , 
 n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , 
 n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , 
 n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , 
 n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , 
 n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , 
 n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , 
 n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , 
 n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , 
 n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , 
 n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , 
 n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , 
 n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , 
 n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , 
 n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , 
 n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , 
 n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , 
 n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , 
 n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , 
 n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , 
 n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , 
 n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , 
 n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , 
 n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , 
 n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , 
 n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , 
 n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , 
 n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , 
 n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , 
 n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , 
 n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , 
 n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , 
 n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , 
 n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , 
 n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , 
 n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , 
 n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , 
 n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , 
 n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , 
 n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , 
 n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , 
 n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , 
 n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , 
 n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , 
 n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , 
 n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , 
 n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , 
 n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , 
 n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , 
 n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , 
 n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , 
 n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , 
 n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , 
 n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , 
 n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , 
 n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , 
 n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , 
 n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , 
 n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , 
 n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , 
 n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , 
 n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , 
 n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , 
 n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , 
 n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , 
 n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , 
 n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , 
 n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , 
 n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , 
 n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , 
 n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , 
 n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , 
 n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , 
 n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , 
 n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , 
 n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , 
 n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , 
 n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , 
 n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , 
 n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , 
 n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , 
 n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , 
 n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , 
 n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , 
 n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , 
 n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , 
 n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , 
 n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , 
 n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , 
 n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , 
 n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , 
 n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , 
 n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , 
 n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , 
 n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , 
 n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , 
 n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , 
 n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , 
 n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , 
 n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , 
 n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , 
 n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , 
 n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , 
 n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , 
 n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , 
 n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , 
 n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , 
 n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , 
 n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , 
 n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , 
 n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , 
 n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , 
 n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , 
 n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , 
 n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , 
 n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , 
 n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , 
 n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , 
 n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , 
 n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , 
 n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , 
 n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , 
 n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , 
 n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , 
 n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , 
 n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , 
 n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , 
 n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , 
 n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , 
 n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , 
 n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , 
 n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , 
 n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , 
 n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , 
 n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , 
 n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , 
 n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , 
 n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , 
 n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , 
 n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , 
 n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , 
 n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , 
 n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , 
 n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , 
 n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , 
 n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , 
 n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , 
 n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , 
 n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , 
 n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , 
 n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , 
 n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , 
 n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , 
 n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , 
 n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , 
 n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , 
 n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , 
 n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , 
 n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , 
 n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , 
 n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , 
 n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , 
 n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , 
 n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , 
 n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , 
 n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , 
 n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , 
 n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , 
 n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , 
 n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , 
 n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , 
 n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , 
 n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , 
 n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , 
 n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , 
 n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , 
 n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , 
 n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , 
 n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , 
 n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , 
 n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , 
 n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , 
 n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , 
 n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , 
 n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , 
 n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , 
 n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , 
 n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , 
 n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , 
 n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , 
 n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , 
 n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , 
 n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , 
 n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , 
 n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , 
 n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , 
 n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , 
 n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , 
 n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , 
 n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , 
 n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , 
 n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , 
 n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , 
 n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , 
 n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , 
 n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , 
 n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , 
 n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , 
 n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , 
 n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , 
 n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , 
 n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , 
 n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , 
 n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , 
 n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , 
 n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , 
 n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , 
 n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , 
 n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , 
 n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , 
 n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , 
 n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , 
 n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , 
 n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , 
 n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , 
 n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , 
 n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , 
 n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , 
 n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , 
 n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , 
 n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , 
 n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , 
 n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , 
 n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , 
 n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , 
 n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , 
 n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , 
 n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , 
 n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , 
 n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , 
 n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , 
 n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , 
 n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , 
 n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , 
 n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , 
 n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , 
 n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , 
 n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , 
 n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , 
 n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , 
 n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , 
 n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , 
 n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , 
 n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , 
 n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , 
 n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , 
 n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , 
 n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , 
 n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , 
 n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , 
 n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , 
 n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , 
 n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , 
 n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , 
 n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , 
 n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , 
 n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , 
 n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , 
 n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , 
 n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , 
 n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , 
 n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , 
 n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , 
 n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , 
 n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , 
 n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , 
 n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , 
 n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , 
 n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , 
 n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , 
 n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , 
 n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , 
 n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , 
 n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , 
 n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , 
 n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , 
 n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , 
 n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , 
 n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , 
 n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , 
 n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , 
 n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , 
 n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , 
 n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , 
 n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , 
 n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , 
 n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , 
 n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , 
 n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , 
 n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , 
 n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , 
 n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , 
 n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , 
 n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , 
 n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , 
 n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , 
 n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , 
 n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , 
 n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , 
 n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , 
 n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , 
 n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , 
 n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , 
 n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , 
 n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , 
 n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , 
 n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , 
 n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , 
 n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , 
 n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , 
 n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , 
 n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , 
 n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , 
 n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , 
 n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , 
 n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , 
 n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , 
 n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , 
 n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , 
 n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , 
 n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , 
 n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , 
 n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , 
 n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , 
 n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , 
 n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , 
 n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , 
 n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , 
 n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , 
 n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , 
 n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , 
 n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , 
 n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , 
 n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , 
 n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , 
 n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , 
 n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , 
 n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , 
 n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , 
 n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , 
 n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , 
 n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , 
 n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , 
 n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , 
 n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , 
 n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , 
 n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , 
 n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , 
 n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , 
 n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , 
 n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , 
 n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , 
 n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , 
 n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , 
 n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , 
 n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , 
 n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , 
 n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , 
 n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , 
 n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , 
 n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , 
 n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , 
 n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , 
 n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , 
 n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , 
 n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , 
 n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , 
 n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , 
 n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , 
 n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , 
 n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , 
 n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , 
 n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , 
 n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , 
 n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , 
 n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , 
 n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , 
 n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , 
 n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , 
 n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , 
 n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , 
 n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , 
 n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , 
 n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , 
 n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , 
 n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , 
 n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , 
 n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , 
 n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , 
 n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , 
 n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , 
 n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , 
 n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , 
 n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , 
 n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , 
 n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , 
 n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , 
 n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , 
 n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , 
 n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , 
 n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , 
 n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , 
 n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , 
 n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , 
 n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , 
 n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , 
 n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , 
 n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , 
 n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , 
 n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , 
 n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , 
 n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , 
 n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , 
 n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , 
 n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , 
 n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , 
 n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , 
 n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , 
 n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , 
 n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , 
 n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , 
 n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , 
 n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , 
 n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , 
 n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , 
 n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , 
 n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , 
 n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , 
 n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , 
 n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , 
 n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , 
 n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , 
 n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , 
 n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , 
 n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , 
 n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , 
 n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , 
 n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , 
 n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , 
 n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , 
 n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , 
 n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , 
 n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , 
 n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , 
 n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , 
 n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , 
 n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , 
 n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , 
 n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , 
 n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , 
 n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , 
 n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , 
 n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , 
 n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , 
 n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , 
 n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , 
 n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , 
 n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , 
 n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , 
 n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , 
 n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , 
 n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , 
 n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , 
 n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , 
 n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , 
 n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , 
 n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , 
 n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , 
 n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , 
 n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , 
 n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , 
 n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , 
 n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , 
 n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , 
 n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , 
 n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , 
 n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , 
 n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , 
 n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , 
 n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , 
 n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , 
 n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , 
 n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , 
 n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , 
 n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , 
 n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , 
 n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , 
 n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , 
 n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , 
 n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , 
 n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , 
 n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , 
 n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , 
 n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , 
 n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , 
 n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , 
 n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , 
 n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , 
 n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , 
 n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , 
 n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , 
 n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , 
 n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , 
 n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , 
 n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , 
 n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , 
 n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , 
 n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , 
 n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , 
 n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , 
 n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , 
 n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , 
 n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , 
 n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , 
 n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , 
 n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , 
 n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , 
 n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , 
 n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , 
 n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , 
 n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , 
 n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , 
 n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , 
 n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , 
 n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , 
 n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , 
 n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , 
 n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , 
 n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , 
 n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , 
 n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , 
 n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , 
 n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , 
 n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , 
 n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , 
 n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , 
 n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , 
 n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , 
 n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , 
 n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , 
 n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , 
 n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , 
 n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , 
 n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , 
 n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , 
 n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , 
 n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , 
 n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , 
 n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , 
 n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , 
 n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , 
 n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , 
 n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , 
 n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , 
 n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , 
 n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , 
 n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , 
 n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , 
 n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , 
 n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , 
 n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , 
 n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , 
 n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , 
 n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , 
 n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , 
 n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , 
 n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , 
 n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , 
 n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , 
 n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , 
 n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , 
 n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , 
 n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , 
 n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , 
 n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , 
 n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , 
 n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , 
 n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , 
 n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , 
 n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , 
 n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , 
 n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , 
 n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , 
 n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , 
 n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , 
 n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , 
 n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , 
 n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , 
 n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , 
 n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , 
 n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , 
 n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , 
 n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , 
 n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , 
 n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , 
 n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , 
 n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , 
 n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , 
 n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , 
 n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , 
 n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , 
 n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , 
 n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , 
 n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , 
 n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , 
 n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , 
 n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , 
 n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , 
 n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , 
 n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , 
 n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , 
 n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , 
 n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , 
 n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , 
 n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , 
 n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , 
 n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , 
 n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , 
 n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , 
 n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , 
 n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , 
 n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , 
 n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , 
 n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , 
 n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , 
 n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , 
 n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , 
 n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , 
 n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , 
 n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , 
 n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , 
 n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , 
 n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , 
 n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , 
 n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , 
 n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , 
 n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , 
 n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , 
 n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , 
 n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , 
 n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , 
 n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , 
 n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , 
 n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , 
 n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , 
 n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , 
 n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , 
 n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , 
 n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , 
 n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , 
 n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , 
 n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , 
 n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , 
 n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , 
 n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , 
 n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , 
 n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , 
 n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , 
 n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , 
 n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , 
 n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , 
 n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , 
 n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , 
 n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , 
 n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , 
 n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , 
 n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , 
 n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , 
 n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , 
 n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , 
 n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , 
 n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , 
 n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , 
 n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , 
 n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , 
 n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , 
 n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , 
 n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , 
 n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , 
 n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , 
 n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , 
 n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , 
 n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , 
 n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , 
 n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , 
 n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , 
 n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , 
 n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , 
 n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , 
 n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , 
 n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , 
 n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , 
 n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , 
 n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , 
 n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , 
 n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , 
 n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , 
 n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , 
 n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , 
 n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , 
 n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , 
 n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , 
 n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , 
 n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , 
 n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , 
 n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , 
 n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , 
 n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , 
 n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , 
 n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , 
 n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , 
 n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , 
 n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , 
 n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , 
 n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , 
 n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , 
 n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , 
 n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , 
 n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , 
 n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , 
 n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , 
 n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , 
 n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , 
 n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , 
 n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , 
 n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , 
 n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , 
 n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , 
 n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , 
 n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , 
 n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , 
 n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , 
 n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , 
 n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , 
 n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , 
 n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , 
 n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , 
 n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , 
 n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , 
 n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , 
 n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , 
 n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , 
 n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , 
 n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , 
 n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , 
 n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , 
 n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , 
 n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , 
 n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , 
 n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , 
 n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , 
 n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , 
 n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , 
 n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , 
 n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , 
 n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , 
 n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , 
 n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , 
 n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , 
 n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , 
 n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , 
 n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , 
 n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , 
 n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , 
 n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , 
 n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , 
 n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , 
 n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , 
 n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , 
 n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , 
 n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , 
 n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , 
 n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , 
 n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , 
 n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , 
 n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , 
 n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , 
 n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , 
 n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , 
 n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , 
 n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , 
 n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , 
 n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , 
 n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , 
 n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , 
 n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , 
 n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , 
 n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , 
 n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , 
 n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , 
 n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , 
 n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , 
 n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , 
 n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , 
 n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , 
 n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , 
 n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , 
 n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , 
 n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , 
 n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , 
 n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , 
 n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , 
 n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , 
 n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , 
 n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , 
 n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , 
 n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , 
 n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , 
 n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , 
 n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , 
 n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , 
 n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , 
 n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , 
 n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , 
 n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , 
 n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , 
 n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , 
 n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , 
 n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , 
 n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , 
 n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , 
 n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , 
 n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , 
 n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , 
 n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , 
 n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , 
 n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , 
 n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , 
 n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , 
 n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , 
 n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , 
 n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , 
 n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , 
 n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , 
 n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , 
 n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , 
 n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , 
 n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , 
 n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , 
 n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , 
 n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , 
 n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , 
 n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , 
 n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , 
 n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , 
 n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , 
 n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , 
 n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , 
 n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , 
 n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , 
 n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , 
 n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , 
 n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , 
 n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , 
 n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , 
 n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , 
 n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , 
 n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , 
 n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , 
 n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , 
 n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , 
 n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , 
 n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , 
 n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , 
 n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , 
 n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , 
 n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , 
 n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , 
 n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , 
 n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , 
 n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , 
 n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , 
 n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , 
 n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , 
 n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , 
 n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , 
 n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , 
 n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , 
 n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , 
 n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , 
 n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , 
 n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , 
 n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , 
 n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , 
 n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , 
 n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , 
 n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , 
 n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , 
 n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , 
 n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , 
 n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , 
 n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , 
 n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , 
 n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , 
 n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , 
 n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , 
 n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , 
 n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , 
 n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , 
 n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , 
 n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , 
 n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , 
 n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , 
 n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , 
 n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , 
 n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , 
 n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , 
 n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , 
 n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , 
 n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , 
 n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , 
 n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , 
 n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , 
 n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , 
 n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , 
 n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , 
 n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , 
 n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , 
 n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , 
 n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , 
 n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , 
 n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , 
 n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , 
 n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , 
 n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , 
 n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , 
 n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , 
 n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , 
 n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , 
 n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , 
 n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , 
 n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , 
 n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , 
 n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , 
 n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , 
 n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , 
 n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , 
 n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , 
 n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , 
 n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , 
 n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , 
 n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , 
 n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , 
 n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , 
 n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , 
 n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , 
 n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , 
 n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , 
 n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , 
 n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , 
 n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , 
 n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , 
 n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , 
 n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , 
 n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , 
 n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , 
 n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , 
 n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , 
 n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , 
 n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , 
 n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , 
 n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , 
 n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , 
 n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , 
 n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , 
 n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , 
 n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , 
 n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , 
 n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , 
 n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , 
 n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , 
 n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , 
 n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , 
 n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , 
 n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , 
 n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , 
 n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , 
 n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , 
 n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , 
 n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , 
 n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , 
 n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , 
 n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , 
 n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , 
 n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , 
 n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , 
 n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , 
 n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , 
 n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , 
 n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , 
 n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , 
 n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , 
 n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , 
 n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , 
 n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , 
 n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , 
 n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , 
 n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , 
 n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , 
 n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , 
 n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , 
 n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , 
 n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , 
 n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , 
 n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , 
 n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , 
 n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , 
 n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , 
 n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , 
 n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , 
 n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , 
 n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , 
 n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , 
 n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , 
 n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , 
 n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , 
 n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , 
 n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , 
 n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , 
 n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , 
 n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , 
 n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , 
 n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , 
 n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , 
 n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , 
 n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , 
 n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , 
 n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , 
 n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , 
 n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , 
 n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , 
 n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , 
 n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , 
 n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , 
 n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , 
 n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , 
 n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , 
 n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , 
 n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , 
 n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , 
 n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , 
 n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , 
 n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , 
 n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , 
 n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , 
 n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , 
 n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , 
 n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , 
 n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , 
 n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , 
 n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , 
 n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , 
 n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , 
 n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , 
 n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , 
 n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , 
 n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , 
 n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , 
 n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , 
 n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , 
 n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , 
 n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , 
 n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , 
 n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , 
 n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , 
 n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , 
 n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , 
 n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , 
 n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , 
 n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , 
 n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , 
 n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , 
 n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , 
 n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , 
 n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , 
 n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , 
 n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , 
 n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , 
 n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , 
 n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , 
 n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , 
 n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , 
 n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , 
 n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , 
 n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , 
 n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , 
 n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , 
 n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , 
 n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , 
 n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , 
 n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , 
 n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , 
 n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , 
 n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , 
 n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , 
 n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , 
 n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , 
 n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , 
 n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , 
 n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , 
 n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , 
 n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , 
 n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , 
 n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , 
 n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , 
 n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , 
 n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , 
 n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , 
 n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , 
 n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , 
 n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , 
 n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , 
 n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , 
 n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , 
 n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , 
 n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , 
 n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , 
 n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , 
 n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , 
 n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , 
 n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , 
 n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , 
 n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , 
 n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , 
 n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , 
 n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , 
 n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , 
 n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , 
 n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , 
 n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , 
 n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , 
 n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , 
 n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , 
 n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , 
 n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , 
 n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , 
 n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , 
 n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , 
 n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , 
 n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , 
 n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , 
 n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , 
 n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , 
 n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , 
 n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , 
 n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , 
 n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , 
 n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , 
 n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , 
 n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , 
 n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , 
 n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , 
 n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , 
 n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , 
 n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , 
 n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , 
 n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , 
 n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , 
 n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , 
 n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , 
 n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , 
 n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , 
 n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , 
 n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , 
 n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , 
 n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , 
 n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , 
 n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , 
 n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , 
 n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , 
 n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , 
 n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , 
 n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , 
 n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , 
 n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , 
 n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , 
 n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , 
 n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , 
 n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , 
 n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , 
 n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , 
 n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , 
 n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , 
 n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , 
 n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , 
 n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , 
 n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , 
 n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , 
 n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , 
 n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , 
 n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , 
 n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , 
 n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , 
 n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , 
 n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , 
 n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , 
 n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , 
 n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , 
 n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , 
 n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , 
 n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , 
 n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , 
 n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , 
 n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , 
 n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , 
 n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , 
 n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , 
 n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , 
 n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , 
 n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , 
 n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , 
 n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , 
 n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , 
 n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , 
 n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , 
 n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , 
 n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , 
 n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , 
 n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , 
 n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , 
 n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , 
 n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , 
 n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , 
 n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , 
 n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , 
 n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , 
 n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , 
 n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , 
 n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , 
 n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , 
 n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , 
 n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , 
 n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , 
 n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , 
 n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , 
 n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , 
 n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , 
 n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , 
 n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , 
 n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , 
 n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , 
 n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , 
 n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , 
 n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , 
 n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , 
 n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , 
 n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , 
 n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , 
 n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , 
 n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , 
 n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , 
 n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , 
 n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , 
 n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , 
 n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , 
 n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , 
 n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , 
 n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , 
 n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , 
 n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , 
 n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , 
 n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , 
 n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , 
 n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , 
 n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , 
 n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , 
 n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , 
 n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , 
 n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , 
 n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , 
 n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , 
 n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , 
 n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , 
 n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , 
 n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , 
 n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , 
 n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , 
 n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , 
 n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , 
 n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , 
 n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , 
 n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , 
 n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , 
 n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , 
 n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , 
 n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , 
 n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , 
 n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , 
 n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , 
 n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , 
 n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , 
 n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , 
 n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , 
 n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , 
 n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , 
 n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , 
 n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , 
 n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , 
 n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , 
 n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , 
 n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , 
 n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , 
 n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , 
 n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , 
 n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , 
 n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , 
 n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , 
 n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , 
 n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , 
 n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , 
 n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , 
 n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , 
 n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , 
 n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , 
 n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , 
 n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , 
 n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , 
 n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , 
 n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , 
 n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , 
 n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , 
 n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , 
 n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , 
 n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , 
 n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , 
 n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , 
 n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , 
 n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , 
 n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , 
 n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , 
 n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , 
 n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , 
 n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , 
 n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , 
 n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , 
 n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , 
 n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , 
 n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , 
 n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , 
 n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , 
 n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , 
 n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , 
 n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , 
 n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , 
 n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , 
 n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , 
 n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , 
 n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , 
 n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , 
 n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , 
 n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , 
 n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , 
 n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , 
 n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , 
 n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , 
 n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , 
 n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , 
 n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , 
 n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , 
 n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , 
 n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , 
 n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , 
 n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , 
 n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , 
 n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , 
 n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , 
 n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , 
 n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , 
 n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , 
 n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , 
 n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , 
 n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , 
 n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , 
 n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , 
 n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , 
 n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , 
 n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , 
 n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , 
 n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , 
 n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , 
 n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , 
 n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , 
 n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , 
 n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , 
 n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , 
 n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , 
 n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , 
 n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , 
 n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , 
 n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , 
 n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , 
 n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , 
 n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , 
 n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , 
 n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , 
 n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , 
 n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , 
 n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , 
 n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , 
 n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , 
 n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , 
 n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , 
 n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , 
 n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , 
 n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , 
 n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , 
 n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , 
 n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , 
 n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , 
 n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , 
 n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , 
 n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , 
 n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , 
 n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , 
 n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , 
 n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , 
 n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , 
 n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , 
 n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , 
 n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , 
 n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , 
 n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , 
 n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , 
 n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , 
 n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , 
 n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , 
 n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , 
 n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , 
 n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , 
 n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , 
 n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , 
 n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , 
 n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , 
 n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , 
 n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , 
 n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , 
 n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , 
 n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , 
 n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , 
 n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , 
 n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , 
 n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , 
 n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , 
 n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , 
 n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , 
 n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , 
 n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , 
 n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , 
 n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , 
 n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , 
 n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , 
 n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , 
 n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , 
 n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , 
 n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , 
 n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , 
 n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , 
 n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , 
 n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , 
 n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , 
 n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , 
 n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , 
 n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , 
 n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , 
 n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , 
 n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , 
 n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , 
 n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , 
 n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , 
 n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , 
 n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , 
 n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , 
 n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , 
 n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , 
 n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , 
 n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , 
 n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , 
 n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , 
 n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , 
 n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , 
 n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , 
 n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , 
 n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , 
 n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , 
 n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , 
 n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , 
 n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , 
 n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , 
 n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , 
 n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , 
 n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , 
 n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , 
 n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , 
 n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , 
 n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , 
 n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , 
 n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , 
 n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , 
 n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , 
 n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , 
 n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , 
 n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , 
 n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , 
 n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , 
 n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , 
 n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , 
 n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , 
 n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , 
 n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , 
 n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , 
 n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , 
 n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , 
 n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , 
 n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , 
 n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , 
 n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , 
 n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , 
 n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , 
 n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , 
 n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , 
 n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , 
 n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , 
 n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , 
 n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , 
 n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , 
 n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , 
 n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , 
 n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , 
 n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , 
 n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , 
 n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , 
 n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , 
 n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , 
 n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , 
 n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , 
 n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , 
 n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , 
 n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , 
 n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , 
 n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , 
 n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , 
 n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , 
 n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , 
 n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , 
 n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , 
 n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , 
 n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , 
 n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , 
 n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , 
 n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , 
 n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , 
 n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , 
 n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , 
 n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , 
 n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , 
 n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , 
 n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , 
 n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , 
 n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , 
 n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , 
 n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , 
 n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , 
 n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , 
 n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , 
 n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , 
 n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , 
 n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , 
 n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , 
 n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , 
 n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , 
 n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , 
 n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , 
 n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , 
 n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , 
 n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , 
 n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , 
 n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , 
 n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , 
 n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , 
 n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , 
 n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , 
 n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , 
 n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , 
 n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , 
 n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , 
 n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , 
 n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , 
 n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , 
 n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , 
 n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , 
 n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , 
 n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , 
 n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , 
 n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , 
 n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , 
 n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , 
 n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , 
 n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , 
 n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , 
 n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , 
 n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , 
 n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , 
 n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , 
 n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , 
 n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , 
 n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , 
 n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , 
 n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , 
 n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , 
 n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , 
 n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , 
 n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , 
 n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , 
 n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , 
 n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , 
 n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , 
 n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , 
 n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , 
 n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , 
 n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , 
 n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , 
 n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , 
 n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , 
 n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , 
 n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , 
 n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , 
 n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , 
 n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , 
 n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , 
 n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , 
 n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , 
 n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , 
 n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , 
 n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , 
 n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , 
 n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , 
 n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , 
 n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , 
 n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , 
 n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , 
 n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , 
 n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , 
 n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , 
 n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , 
 n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , 
 n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , 
 n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , 
 n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , 
 n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , 
 n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , 
 n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , 
 n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , 
 n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , 
 n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , 
 n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , 
 n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , 
 n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , 
 n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , 
 n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , 
 n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , 
 n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , 
 n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , 
 n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , 
 n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , 
 n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , 
 n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , 
 n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , 
 n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , 
 n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , 
 n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , 
 n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , 
 n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , 
 n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , 
 n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , 
 n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , 
 n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , 
 n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , 
 n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , 
 n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , 
 n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , 
 n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , 
 n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , 
 n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , 
 n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , 
 n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , 
 n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , 
 n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , 
 n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , 
 n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , 
 n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , 
 n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , 
 n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , 
 n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , 
 n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , 
 n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , 
 n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , 
 n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , 
 n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , 
 n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , 
 n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , 
 n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , 
 n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , 
 n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , 
 n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , 
 n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , 
 n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , 
 n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , 
 n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , 
 n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , 
 n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , 
 n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , 
 n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , 
 n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , 
 n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , 
 n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , 
 n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , 
 n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , 
 n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , 
 n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , 
 n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , 
 n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , 
 n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , 
 n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , 
 n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , 
 n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , 
 n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , 
 n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , 
 n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , 
 n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , 
 n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , 
 n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , 
 n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , 
 n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , 
 n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , 
 n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , 
 n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , 
 n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , 
 n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , 
 n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , 
 n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , 
 n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , 
 n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , 
 n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , 
 n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , 
 n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , 
 n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , 
 n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , 
 n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , 
 n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , 
 n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , 
 n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , 
 n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , 
 n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , 
 n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , 
 n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , 
 n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , 
 n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , 
 n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , 
 n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , 
 n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , 
 n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , 
 n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , 
 n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , 
 n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , 
 n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , 
 n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , 
 n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , 
 n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , 
 n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , 
 n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , 
 n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , 
 n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , 
 n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , 
 n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , 
 n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , 
 n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , 
 n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , 
 n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , 
 n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , 
 n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , 
 n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , 
 n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , 
 n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , 
 n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , 
 n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , 
 n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , 
 n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , 
 n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , 
 n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , 
 n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , 
 n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , 
 n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , 
 n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , 
 n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , 
 n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , 
 n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , 
 n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , 
 n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , 
 n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , 
 n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , 
 n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , 
 n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , 
 n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , 
 n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , 
 n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , 
 n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , 
 n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , 
 n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , 
 n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , 
 n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , 
 n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , 
 n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , 
 n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , 
 n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , 
 n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , 
 n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , 
 n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , 
 n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , 
 n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , 
 n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , 
 n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , 
 n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , 
 n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , 
 n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , 
 n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , 
 n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , 
 n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , 
 n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , 
 n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , 
 n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , 
 n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , 
 n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , 
 n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , 
 n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , 
 n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , 
 n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , 
 n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , 
 n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , 
 n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , 
 n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , 
 n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , 
 n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , 
 n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , 
 n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , 
 n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , 
 n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , 
 n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , 
 n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , 
 n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , 
 n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , 
 n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , 
 n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , 
 n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , 
 n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , 
 n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , 
 n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , 
 n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , 
 n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , 
 n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , 
 n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , 
 n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , 
 n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , 
 n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , 
 n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , 
 n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , 
 n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , 
 n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , 
 n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , 
 n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , 
 n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , 
 n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , 
 n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , 
 n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , 
 n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , 
 n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , 
 n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , 
 n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , 
 n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , 
 n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , 
 n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , 
 n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , 
 n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , 
 n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , 
 n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , 
 n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , 
 n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , 
 n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , 
 n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , 
 n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , 
 n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , 
 n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , 
 n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , 
 n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , 
 n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , 
 n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , 
 n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , 
 n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , 
 n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , 
 n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , 
 n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , 
 n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , 
 n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , 
 n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , 
 n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , 
 n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , 
 n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , 
 n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , 
 n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , 
 n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , 
 n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , 
 n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , 
 n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , 
 n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , 
 n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , 
 n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , 
 n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , 
 n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , 
 n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , 
 n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , 
 n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , 
 n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , 
 n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , 
 n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , 
 n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , 
 n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , 
 n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , 
 n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , 
 n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , 
 n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , 
 n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , 
 n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , 
 n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , 
 n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , 
 n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , 
 n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , 
 n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , 
 n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , 
 n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , 
 n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , 
 n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , 
 n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , 
 n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , 
 n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , 
 n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , 
 n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , 
 n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , 
 n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , 
 n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , 
 n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , 
 n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , 
 n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , 
 n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , 
 n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , 
 n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , 
 n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , 
 n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , 
 n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , 
 n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , 
 n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , 
 n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , 
 n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , 
 n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , 
 n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , 
 n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , 
 n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , 
 n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , 
 n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , 
 n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , 
 n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , 
 n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , 
 n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , 
 n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , 
 n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , 
 n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , 
 n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , 
 n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , 
 n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , 
 n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , 
 n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , 
 n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , 
 n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , 
 n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , 
 n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , 
 n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , 
 n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , 
 n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , 
 n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , 
 n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , 
 n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , 
 n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , 
 n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , 
 n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , 
 n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , 
 n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , 
 n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , 
 n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , 
 n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , 
 n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , 
 n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , 
 n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , 
 n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , 
 n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , 
 n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , 
 n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , 
 n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , 
 n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , 
 n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , 
 n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , 
 n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , 
 n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , 
 n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , 
 n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , 
 n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , 
 n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , 
 n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , 
 n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , 
 n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , 
 n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , 
 n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , 
 n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , 
 n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , 
 n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , 
 n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , 
 n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , 
 n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , 
 n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , 
 n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , 
 n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , 
 n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , 
 n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , 
 n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , 
 n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , 
 n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , 
 n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , 
 n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , 
 n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , 
 n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , 
 n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , 
 n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , 
 n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , 
 n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , 
 n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , 
 n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , 
 n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , 
 n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , 
 n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , 
 n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , 
 n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , 
 n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , 
 n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , 
 n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , 
 n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , 
 n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , 
 n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , 
 n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , 
 n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , 
 n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , 
 n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , 
 n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , 
 n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , 
 n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , 
 n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , 
 n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , 
 n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , 
 n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , 
 n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , 
 n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , 
 n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , 
 n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , 
 n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , 
 n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , 
 n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , 
 n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , 
 n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , 
 n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , 
 n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , 
 n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , 
 n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , 
 n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , 
 n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , 
 n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , 
 n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , 
 n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , 
 n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , 
 n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , 
 n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , 
 n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , 
 n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , 
 n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , 
 n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , 
 n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , 
 n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , 
 n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , 
 n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , 
 n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , 
 n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , 
 n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , 
 n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , 
 n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , 
 n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , 
 n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , 
 n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , 
 n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , 
 n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , 
 n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , 
 n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , 
 n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , 
 n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , 
 n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , 
 n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , 
 n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , 
 n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , 
 n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , 
 n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , 
 n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , 
 n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , 
 n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , 
 n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , 
 n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , 
 n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , 
 n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , 
 n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , 
 n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , 
 n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , 
 n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , 
 n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , 
 n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , 
 n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , 
 n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , 
 n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , 
 n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , 
 n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , 
 n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , 
 n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , 
 n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , 
 n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , 
 n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , 
 n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , 
 n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , 
 n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , 
 n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , 
 n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , 
 n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , 
 n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , 
 n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , 
 n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , 
 n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , 
 n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , 
 n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , 
 n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , 
 n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , 
 n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , 
 n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , 
 n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , 
 n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , 
 n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , 
 n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , 
 n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , 
 n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , 
 n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , 
 n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , 
 n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , 
 n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , 
 n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , 
 n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , 
 n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , 
 n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , 
 n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , 
 n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , 
 n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , 
 n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , 
 n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , 
 n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , 
 n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , 
 n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , 
 n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , 
 n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , 
 n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , 
 n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , 
 n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , 
 n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , 
 n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , 
 n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , 
 n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , 
 n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , 
 n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , 
 n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , 
 n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , 
 n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , 
 n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , 
 n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , 
 n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , 
 n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , 
 n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , 
 n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , 
 n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , 
 n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , 
 n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , 
 n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , 
 n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , 
 n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , 
 n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , 
 n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , 
 n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , 
 n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , 
 n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , 
 n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , 
 n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , 
 n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , 
 n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , 
 n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , 
 n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , 
 n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , 
 n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , 
 n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , 
 n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , 
 n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , 
 n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , 
 n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , 
 n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , 
 n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , 
 n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , 
 n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , 
 n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , 
 n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , 
 n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , 
 n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , 
 n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , 
 n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , 
 n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , 
 n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , 
 n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , 
 n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , 
 n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , 
 n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , 
 n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , 
 n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , 
 n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , 
 n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , 
 n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , 
 n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , 
 n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , 
 n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , 
 n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , 
 n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , 
 n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , 
 n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , 
 n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , 
 n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , 
 n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , 
 n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , 
 n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , 
 n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , 
 n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , 
 n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , 
 n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , 
 n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , 
 n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , 
 n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , 
 n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , 
 n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , 
 n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , 
 n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , 
 n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , 
 n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , 
 n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , 
 n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , 
 n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , 
 n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , 
 n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , 
 n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , 
 n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , 
 n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , 
 n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , 
 n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , 
 n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , 
 n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , 
 n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , 
 n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , 
 n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , 
 n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , 
 n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , 
 n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , 
 n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , 
 n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , 
 n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , 
 n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , 
 n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , 
 n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , 
 n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , 
 n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , 
 n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , 
 n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , 
 n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , 
 n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , 
 n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , 
 n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , 
 n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , 
 n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , 
 n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , 
 n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , 
 n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , 
 n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , 
 n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , 
 n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , 
 n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , 
 n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , 
 n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , 
 n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , 
 n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , 
 n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , 
 n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , 
 n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , 
 n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , 
 n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , 
 n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , 
 n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , 
 n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , 
 n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , 
 n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , 
 n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , 
 n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , 
 n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , 
 n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , 
 n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , 
 n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , 
 n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , 
 n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , 
 n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , 
 n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , 
 n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , 
 n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , 
 n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , 
 n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , 
 n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , 
 n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , 
 n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , 
 n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , 
 n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , 
 n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , 
 n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , 
 n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , 
 n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , 
 n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , 
 n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , 
 n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , 
 n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , 
 n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , 
 n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , 
 n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , 
 n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , 
 n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , 
 n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , 
 n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , 
 n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , 
 n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , 
 n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , 
 n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , 
 n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , 
 n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , 
 n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , 
 n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , 
 n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , 
 n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , 
 n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , 
 n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , 
 n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , 
 n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , 
 n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , 
 n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , 
 n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , 
 n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , 
 n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , 
 n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , 
 n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , 
 n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , 
 n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , 
 n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , 
 n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , 
 n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , 
 n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , 
 n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , 
 n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , 
 n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , 
 n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , 
 n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , 
 n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , 
 n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , 
 n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , 
 n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , 
 n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , 
 n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , 
 n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , 
 n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , 
 n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , 
 n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , 
 n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , 
 n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , 
 n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , 
 n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , 
 n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , 
 n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , 
 n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , 
 n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , 
 n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , 
 n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , 
 n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , 
 n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , 
 n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , 
 n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , 
 n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , 
 n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , 
 n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , 
 n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , 
 n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , 
 n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , 
 n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , 
 n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , 
 n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , 
 n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , 
 n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , 
 n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , 
 n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , 
 n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , 
 n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , 
 n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , 
 n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , 
 n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , 
 n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , 
 n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , 
 n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , 
 n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , 
 n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , 
 n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , 
 n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , 
 n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , 
 n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , 
 n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , 
 n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , 
 n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , 
 n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , 
 n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , 
 n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , 
 n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , 
 n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , 
 n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , 
 n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , 
 n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , 
 n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , 
 n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , 
 n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , 
 n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , 
 n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , 
 n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , 
 n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , 
 n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , 
 n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , 
 n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , 
 n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , 
 n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , 
 n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , 
 n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , 
 n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , 
 n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , 
 n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , 
 n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , 
 n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , 
 n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , 
 n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , 
 n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , 
 n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , 
 n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , 
 n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , 
 n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , 
 n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , 
 n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , 
 n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , 
 n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , 
 n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , 
 n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , 
 n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , 
 n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , 
 n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , 
 n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , 
 n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , 
 n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , 
 n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , 
 n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , 
 n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , 
 n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , 
 n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , 
 n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , 
 n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , 
 n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , 
 n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , 
 n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , 
 n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , 
 n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , 
 n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , 
 n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , 
 n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , 
 n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , 
 n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , 
 n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , 
 n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , 
 n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , 
 n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , 
 n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , 
 n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , 
 n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , 
 n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , 
 n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , 
 n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , 
 n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , 
 n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , 
 n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , 
 n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , 
 n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , 
 n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , 
 n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , 
 n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , 
 n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , 
 n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , 
 n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , 
 n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , 
 n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , 
 n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , 
 n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , 
 n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , 
 n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , 
 n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , 
 n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , 
 n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , 
 n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , 
 n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , 
 n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , 
 n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , 
 n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , 
 n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , 
 n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , 
 n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , 
 n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , 
 n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , 
 n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , 
 n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , 
 n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , 
 n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , 
 n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , 
 n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , 
 n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , 
 n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , 
 n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , 
 n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , 
 n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , 
 n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , 
 n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , 
 n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , 
 n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , 
 n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , 
 n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , 
 n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , 
 n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , 
 n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , 
 n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , 
 n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , 
 n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , 
 n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , 
 n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , 
 n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , 
 n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , 
 n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , 
 n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , 
 n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , 
 n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , 
 n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , 
 n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , 
 n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , 
 n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , 
 n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , 
 n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , 
 n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , 
 n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , 
 n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , 
 n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , 
 n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , 
 n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , 
 n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , 
 n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , 
 n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , 
 n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , 
 n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , 
 n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , 
 n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , 
 n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , 
 n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , 
 n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , 
 n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , 
 n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , 
 n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , 
 n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , 
 n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , 
 n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , 
 n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , 
 n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , 
 n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , 
 n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , 
 n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , 
 n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , 
 n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , 
 n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , 
 n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , 
 n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , 
 n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , 
 n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , 
 n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , 
 n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , 
 n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , 
 n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , 
 n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , 
 n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , 
 n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , 
 n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , 
 n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , 
 n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , 
 n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , 
 n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , 
 n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , 
 n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , 
 n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , 
 n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , 
 n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , 
 n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , 
 n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , 
 n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , 
 n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , 
 n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , 
 n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , 
 n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , 
 n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , 
 n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , 
 n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , 
 n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , 
 n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , 
 n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , 
 n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , 
 n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , 
 n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , 
 n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , 
 n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , 
 n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , 
 n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , 
 n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , 
 n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , 
 n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , 
 n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , 
 n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , 
 n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , 
 n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , 
 n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , 
 n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , 
 n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , 
 n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , 
 n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , 
 n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , 
 n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , 
 n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , 
 n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , 
 n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , 
 n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , 
 n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , 
 n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , 
 n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , 
 n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , 
 n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , 
 n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , 
 n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , 
 n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , 
 n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , 
 n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , 
 n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , 
 n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , 
 n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , 
 n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , 
 n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , 
 n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , 
 n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , 
 n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , 
 n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , 
 n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , 
 n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , 
 n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , 
 n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , 
 n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , 
 n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , 
 n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , 
 n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , 
 n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , 
 n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , 
 n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , 
 n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , 
 n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , 
 n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , 
 n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , 
 n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , 
 n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , 
 n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , 
 n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , 
 n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , 
 n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , 
 n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , 
 n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , 
 n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , 
 n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , 
 n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , 
 n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , 
 n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , 
 n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , 
 n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , 
 n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , 
 n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , 
 n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , 
 n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , 
 n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , 
 n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , 
 n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , 
 n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , 
 n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , 
 n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , 
 n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , 
 n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , 
 n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , 
 n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , 
 n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , 
 n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , 
 n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , 
 n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , 
 n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , 
 n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , 
 n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , 
 n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , 
 n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , 
 n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , 
 n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , 
 n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , 
 n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , 
 n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , 
 n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , 
 n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , 
 n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , 
 n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , 
 n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , 
 n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , 
 n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , 
 n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , 
 n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , 
 n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , 
 n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , 
 n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , 
 n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , 
 n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , 
 n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , 
 n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , 
 n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , 
 n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , 
 n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , 
 n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , 
 n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , 
 n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , 
 n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , 
 n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , 
 n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , 
 n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , 
 n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , 
 n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , 
 n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , 
 n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , 
 n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , 
 n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , 
 n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , 
 n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , 
 n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , 
 n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , 
 n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , 
 n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , 
 n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , 
 n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , 
 n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , 
 n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , 
 n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , 
 n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , 
 n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , 
 n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , 
 n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , 
 n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , 
 n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , 
 n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , 
 n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , 
 n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , 
 n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , 
 n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , 
 n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , 
 n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , 
 n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , 
 n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , 
 n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , 
 n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , 
 n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , 
 n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , 
 n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , 
 n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , 
 n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , 
 n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , 
 n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , 
 n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , 
 n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , 
 n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , 
 n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , 
 n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , 
 n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , 
 n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , 
 n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , 
 n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , 
 n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , 
 n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , 
 n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , 
 n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , 
 n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , 
 n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , 
 n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , 
 n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , 
 n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , 
 n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , 
 n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , 
 n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , 
 n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , 
 n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , 
 n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , 
 n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , 
 n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , 
 n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , 
 n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , 
 n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , 
 n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , 
 n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , 
 n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , 
 n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , 
 n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , 
 n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , 
 n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , 
 n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , 
 n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , 
 n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , 
 n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , 
 n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , 
 n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , 
 n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , 
 n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , 
 n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , 
 n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , 
 n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , 
 n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , 
 n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , 
 n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , 
 n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , 
 n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , 
 n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , 
 n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , 
 n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , 
 n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , 
 n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , 
 n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , 
 n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , 
 n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , 
 n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , 
 n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , 
 n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , 
 n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , 
 n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , 
 n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , 
 n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , 
 n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , 
 n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , 
 n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , 
 n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , 
 n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , 
 n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , 
 n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , 
 n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , 
 n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , 
 n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , 
 n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , 
 n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , 
 n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , 
 n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , 
 n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , 
 n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , 
 n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , 
 n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , 
 n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , 
 n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , 
 n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , 
 n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , 
 n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , 
 n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , 
 n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , 
 n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , 
 n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , 
 n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , 
 n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , 
 n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , 
 n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , 
 n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , 
 n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , 
 n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , 
 n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , 
 n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , 
 n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , 
 n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , 
 n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , 
 n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , 
 n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , 
 n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , 
 n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , 
 n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , 
 n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , 
 n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , 
 n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , 
 n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , 
 n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , 
 n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , 
 n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , 
 n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , 
 n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , 
 n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , 
 n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , 
 n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , 
 n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , 
 n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , 
 n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , 
 n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , 
 n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , 
 n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , 
 n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , 
 n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , 
 n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , 
 n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , 
 n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , 
 n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , 
 n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , 
 n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , 
 n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , 
 n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , 
 n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , 
 n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , 
 n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , 
 n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , 
 n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , 
 n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , 
 n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , 
 n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , 
 n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , 
 n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , 
 n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , 
 n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , 
 n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , 
 n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , 
 n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , 
 n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , 
 n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , 
 n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , 
 n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , 
 n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , 
 n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , 
 n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , 
 n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , 
 n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , 
 n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , 
 n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , 
 n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , 
 n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , 
 n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , 
 n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , 
 n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , 
 n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , 
 n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , 
 n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , 
 n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , 
 n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , 
 n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , 
 n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , 
 n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , 
 n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , 
 n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , 
 n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , 
 n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , 
 n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , 
 n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , 
 n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , 
 n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , 
 n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , 
 n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , 
 n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , 
 n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , 
 n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , 
 n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , 
 n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , 
 n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , 
 n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , 
 n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , 
 n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , 
 n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , 
 n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , 
 n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , 
 n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , 
 n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , 
 n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , 
 n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , 
 n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , 
 n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , 
 n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , 
 n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , 
 n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , 
 n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , 
 n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , 
 n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , 
 n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , 
 n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , 
 n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , 
 n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , 
 n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , 
 n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , 
 n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , 
 n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , 
 n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , 
 n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , 
 n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , 
 n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , 
 n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , 
 n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , 
 n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , 
 n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , 
 n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , 
 n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , 
 n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , 
 n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , 
 n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , 
 n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , 
 n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , 
 n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , 
 n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , 
 n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , 
 n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , 
 n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , 
 n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , 
 n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , 
 n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , 
 n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , 
 n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , 
 n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , 
 n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , 
 n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , 
 n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , 
 n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , 
 n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , 
 n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , 
 n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , 
 n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , 
 n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , 
 n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , 
 n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , 
 n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , 
 n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , 
 n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , 
 n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , 
 n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , 
 n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , 
 n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , 
 n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , 
 n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , 
 n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , 
 n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , 
 n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , 
 n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , 
 n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , 
 n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , 
 n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , 
 n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , 
 n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , 
 n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , 
 n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , 
 n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , 
 n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , 
 n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , 
 n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , 
 n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , 
 n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , 
 n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , 
 n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , 
 n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , 
 n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , 
 n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , 
 n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , 
 n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , 
 n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , 
 n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , 
 n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , 
 n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , 
 n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , 
 n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , 
 n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , 
 n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , 
 n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , 
 n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , 
 n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , 
 n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , 
 n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , 
 n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , 
 n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , 
 n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , 
 n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , 
 n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , 
 n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , 
 n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , 
 n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , 
 n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , 
 n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , 
 n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , 
 n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , 
 n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , 
 n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , 
 n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , 
 n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , 
 n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , 
 n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , 
 n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , 
 n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , 
 n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , 
 n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , 
 n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , 
 n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , 
 n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , 
 n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , 
 n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , 
 n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , 
 n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , 
 n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , 
 n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , 
 n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , 
 n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , 
 n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , 
 n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , 
 n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , 
 n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , 
 n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , 
 n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , 
 n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , 
 n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , 
 n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , 
 n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , 
 n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , 
 n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , 
 n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , 
 n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , 
 n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , 
 n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , 
 n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , 
 n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , 
 n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , 
 n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , 
 n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , 
 n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , 
 n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , 
 n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , 
 n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , 
 n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , 
 n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , 
 n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , 
 n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , 
 n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , 
 n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , 
 n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , 
 n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , 
 n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , 
 n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , 
 n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , 
 n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , 
 n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , 
 n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , 
 n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , 
 n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , 
 n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , 
 n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , 
 n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , 
 n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , 
 n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , 
 n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , 
 n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , 
 n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , 
 n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , 
 n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , 
 n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , 
 n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , 
 n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , 
 n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , 
 n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , 
 n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , 
 n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , 
 n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , 
 n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , 
 n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , 
 n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , 
 n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , 
 n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , 
 n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , 
 n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , 
 n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , 
 n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , 
 n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , 
 n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , 
 n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , 
 n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , 
 n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , 
 n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , 
 n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , 
 n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , 
 n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , 
 n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , 
 n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , 
 n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , 
 n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , 
 n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , 
 n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , 
 n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , 
 n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , 
 n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , 
 n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , 
 n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , 
 n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , 
 n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , 
 n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , 
 n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , 
 n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , 
 n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , 
 n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , 
 n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , 
 n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , 
 n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , 
 n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , 
 n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , 
 n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , 
 n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , 
 n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , 
 n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , 
 n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , 
 n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , 
 n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , 
 n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , 
 n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , 
 n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , 
 n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , 
 n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , 
 n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , 
 n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , 
 n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , 
 n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , 
 n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , 
 n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , 
 n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , 
 n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , 
 n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , 
 n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , 
 n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , 
 n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , 
 n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , 
 n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , 
 n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , 
 n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , 
 n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , 
 n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , 
 n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , 
 n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , 
 n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , 
 n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , 
 n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , 
 n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , 
 n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , 
 n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , 
 n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , 
 n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , 
 n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , 
 n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , 
 n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , 
 n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , 
 n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , 
 n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , 
 n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , 
 n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , 
 n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , 
 n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , 
 n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , 
 n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , 
 n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , 
 n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , 
 n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , 
 n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , 
 n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , 
 n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , 
 n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , 
 n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , 
 n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , 
 n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , 
 n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , 
 n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , 
 n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , 
 n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , 
 n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , 
 n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , 
 n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , 
 n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , 
 n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , 
 n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , 
 n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , 
 n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , 
 n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , 
 n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , 
 n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , 
 n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , 
 n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , 
 n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , 
 n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , 
 n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , 
 n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , 
 n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , 
 n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , 
 n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , 
 n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , 
 n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , 
 n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , 
 n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , 
 n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , 
 n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , 
 n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , 
 n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , 
 n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , 
 n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , 
 n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , 
 n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , 
 n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , 
 n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , 
 n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , 
 n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , 
 n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , 
 n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , 
 n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , 
 n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , 
 n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , 
 n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , 
 n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , 
 n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , 
 n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , 
 n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , 
 n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , 
 n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , 
 n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , 
 n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , 
 n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , 
 n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , 
 n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , 
 n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , 
 n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , 
 n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , 
 n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , 
 n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , 
 n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , 
 n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , 
 n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , 
 n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , 
 n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , 
 n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , 
 n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , 
 n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , 
 n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , 
 n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , 
 n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , 
 n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , 
 n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , 
 n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , 
 n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , 
 n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , 
 n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , 
 n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , 
 n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , 
 n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , 
 n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , 
 n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , 
 n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , 
 n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , 
 n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , 
 n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , 
 n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , 
 n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , 
 n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , 
 n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , 
 n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , 
 n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , 
 n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , 
 n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , 
 n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , 
 n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , 
 n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , 
 n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , 
 n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , 
 n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , 
 n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , 
 n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , 
 n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , 
 n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , 
 n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , 
 n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , 
 n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , 
 n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , 
 n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , 
 n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , 
 n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , 
 n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , 
 n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , 
 n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , 
 n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , 
 n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , 
 n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , 
 n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , 
 n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , 
 n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , 
 n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , 
 n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , 
 n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , 
 n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , 
 n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , 
 n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , 
 n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , 
 n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , 
 n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , 
 n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , 
 n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , 
 n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , 
 n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , 
 n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , 
 n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , 
 n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , 
 n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , 
 n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , 
 n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , 
 n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , 
 n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , 
 n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , 
 n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , 
 n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , 
 n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , 
 n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , 
 n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , 
 n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , 
 n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , 
 n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , 
 n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , 
 n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , 
 n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , 
 n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , 
 n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , 
 n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , 
 n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , 
 n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , 
 n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , 
 n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , 
 n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , 
 n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , 
 n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , 
 n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , 
 n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , 
 n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , 
 n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , 
 n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , 
 n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , 
 n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , 
 n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , 
 n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , 
 n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , 
 n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , 
 n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , 
 n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , 
 n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , 
 n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , 
 n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , 
 n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , 
 n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , 
 n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , 
 n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , 
 n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , 
 n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , 
 n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , 
 n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , 
 n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , 
 n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , 
 n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , 
 n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , 
 n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , 
 n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , 
 n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , 
 n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , 
 n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , 
 n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , 
 n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , 
 n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , 
 n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , 
 n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , 
 n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , 
 n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , 
 n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , 
 n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , 
 n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , 
 n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , 
 n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , 
 n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , 
 n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , 
 n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , 
 n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , 
 n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , 
 n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , 
 n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , 
 n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , 
 n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , 
 n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , 
 n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , 
 n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , 
 n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , 
 n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , 
 n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , 
 n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , 
 n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , 
 n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , 
 n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , 
 n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , 
 n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , 
 n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , 
 n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , 
 n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , 
 n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , 
 n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , 
 n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , 
 n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , 
 n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , 
 n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , 
 n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , 
 n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , 
 n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , 
 n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , 
 n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , 
 n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , 
 n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , 
 n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , 
 n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , 
 n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , 
 n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , 
 n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , 
 n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , 
 n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , 
 n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , 
 n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , 
 n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , 
 n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , 
 n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , 
 n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , 
 n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , 
 n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , 
 n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , 
 n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , 
 n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , 
 n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , 
 n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , 
 n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , 
 n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , 
 n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , 
 n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , 
 n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , 
 n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , 
 n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , 
 n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , 
 n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , 
 n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , 
 n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , 
 n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , 
 n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , 
 n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , 
 n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , 
 n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , 
 n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , 
 n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , 
 n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , 
 n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , 
 n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , 
 n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , 
 n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , 
 n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , 
 n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , 
 n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , 
 n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , 
 n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , 
 n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , 
 n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , 
 n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , 
 n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , 
 n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , 
 n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , 
 n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , 
 n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , 
 n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , 
 n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , 
 n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , 
 n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , 
 n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , 
 n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , 
 n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , 
 n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , 
 n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , 
 n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , 
 n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , 
 n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , 
 n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , 
 n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , 
 n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , 
 n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , 
 n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , 
 n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , 
 n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , 
 n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , 
 n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , 
 n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , 
 n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , 
 n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , 
 n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , 
 n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , 
 n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , 
 n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , 
 n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , 
 n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , 
 n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , 
 n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , 
 n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , 
 n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , 
 n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , 
 n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , 
 n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , 
 n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , 
 n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , 
 n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , 
 n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , 
 n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , 
 n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , 
 n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , 
 n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , 
 n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , 
 n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , 
 n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , 
 n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , 
 n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , 
 n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , 
 n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , 
 n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , 
 n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , 
 n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , 
 n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , 
 n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , 
 n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , 
 n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , 
 n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , 
 n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , 
 n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , 
 n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , 
 n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , 
 n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , 
 n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , 
 n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , 
 n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , 
 n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , 
 n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , 
 n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , 
 n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , 
 n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , 
 n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , 
 n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , 
 n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , 
 n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , 
 n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , 
 n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , 
 n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , 
 n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , 
 n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , 
 n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , 
 n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , 
 n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , 
 n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , 
 n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , 
 n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , 
 n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , 
 n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , 
 n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , 
 n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , 
 n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , 
 n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , 
 n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , 
 n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , 
 n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , 
 n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , 
 n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , 
 n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , 
 n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , 
 n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , 
 n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , 
 n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , 
 n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , 
 n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , 
 n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , 
 n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , 
 n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , 
 n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , 
 n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , 
 n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , 
 n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , 
 n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , 
 n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , 
 n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , 
 n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , 
 n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , 
 n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , 
 n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , 
 n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , 
 n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , 
 n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , 
 n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , 
 n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , 
 n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , 
 n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , 
 n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , 
 n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , 
 n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , 
 n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , 
 n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , 
 n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , 
 n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , 
 n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , 
 n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , 
 n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , 
 n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , 
 n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , 
 n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , 
 n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , 
 n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , 
 n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , 
 n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , 
 n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , 
 n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , 
 n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , 
 n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , 
 n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , 
 n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , 
 n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , 
 n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , 
 n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , 
 n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , 
 n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , 
 n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , 
 n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , 
 n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , 
 n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , 
 n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , 
 n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , 
 n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , 
 n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , 
 n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , 
 n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , 
 n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , 
 n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , 
 n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , 
 n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , 
 n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , 
 n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , 
 n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , 
 n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , 
 n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , 
 n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , 
 n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , 
 n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , 
 n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , 
 n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , 
 n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , 
 n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , 
 n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , 
 n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , 
 n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , 
 n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , 
 n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , 
 n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , 
 n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , 
 n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , 
 n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , 
 n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , 
 n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , 
 n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , 
 n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , 
 n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , 
 n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , 
 n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , 
 n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , 
 n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , 
 n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , 
 n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , 
 n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , 
 n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , 
 n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , 
 n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , 
 n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , 
 n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , 
 n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , 
 n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , 
 n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , 
 n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , 
 n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , 
 n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , 
 n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , 
 n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , 
 n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , 
 n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , 
 n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , 
 n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , 
 n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , 
 n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , 
 n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , 
 n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , 
 n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , 
 n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , 
 n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , 
 n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , 
 n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , 
 n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , 
 n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , 
 n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , 
 n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , 
 n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , 
 n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , 
 n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , 
 n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , 
 n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , 
 n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , 
 n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , 
 n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , 
 n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , 
 n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , 
 n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , 
 n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , 
 n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , 
 n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , 
 n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , 
 n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , 
 n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , 
 n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , 
 n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , 
 n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , 
 n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , 
 n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , 
 n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , 
 n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , 
 n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , 
 n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , 
 n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , 
 n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , 
 n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , 
 n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , 
 n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , 
 n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , 
 n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , 
 n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , 
 n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , 
 n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , 
 n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , 
 n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , 
 n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , 
 n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , 
 n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , 
 n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , 
 n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , 
 n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , 
 n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , 
 n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , 
 n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , 
 n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , 
 n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , 
 n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , 
 n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , 
 n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , 
 n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , 
 n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , 
 n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , 
 n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , 
 n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , 
 n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , 
 n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , 
 n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , 
 n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , 
 n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , 
 n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , 
 n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , 
 n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , 
 n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , 
 n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , 
 n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , 
 n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , 
 n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , 
 n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , 
 n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , 
 n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , 
 n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , 
 n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , 
 n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , 
 n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , 
 n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , 
 n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , 
 n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , 
 n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , 
 n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , 
 n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , 
 n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , 
 n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , 
 n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , 
 n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , 
 n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , 
 n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , 
 n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , 
 n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , 
 n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , 
 n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , 
 n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , 
 n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , 
 n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , 
 n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , 
 n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , 
 n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , 
 n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , 
 n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , 
 n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , 
 n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , 
 n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , 
 n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , 
 n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , 
 n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , 
 n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , 
 n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , 
 n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , 
 n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , 
 n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , 
 n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , 
 n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , 
 n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , 
 n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , 
 n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , 
 n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , 
 n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , 
 n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , 
 n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , 
 n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , 
 n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , 
 n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , 
 n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , 
 n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , 
 n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , 
 n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , 
 n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , 
 n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , 
 n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , 
 n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , 
 n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , 
 n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , 
 n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , 
 n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , 
 n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , 
 n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , 
 n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , 
 n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , 
 n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , 
 n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , 
 n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , 
 n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , 
 n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , 
 n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , 
 n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , 
 n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , 
 n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , 
 n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , 
 n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , 
 n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , 
 n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , 
 n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , 
 n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , 
 n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , 
 n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , 
 n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , 
 n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , 
 n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , 
 n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , 
 n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , 
 n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , 
 n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , 
 n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , 
 n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , 
 n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , 
 n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , 
 n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , 
 n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , 
 n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , 
 n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , 
 n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , 
 n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , 
 n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , 
 n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , 
 n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , 
 n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , 
 n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , 
 n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , 
 n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , 
 n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , 
 n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , 
 n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , 
 n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , 
 n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , 
 n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , 
 n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , 
 n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , 
 n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , 
 n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , 
 n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , 
 n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , 
 n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , 
 n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , 
 n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , 
 n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , 
 n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , 
 n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , 
 n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , 
 n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , 
 n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , 
 n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , 
 n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , 
 n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , 
 n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , 
 n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , 
 n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , 
 n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , 
 n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , 
 n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , 
 n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , 
 n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , 
 n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , 
 n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , 
 n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , 
 n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , 
 n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , 
 n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , 
 n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , 
 n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , 
 n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , 
 n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , 
 n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , 
 n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , 
 n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , 
 n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , 
 n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , 
 n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , 
 n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , 
 n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , 
 n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , 
 n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , 
 n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , 
 n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , 
 n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , 
 n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , 
 n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , 
 n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , 
 n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , 
 n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , 
 n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , 
 n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , 
 n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , 
 n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , 
 n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , 
 n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , 
 n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , 
 n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , 
 n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , 
 n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , 
 n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , n54147 , n54148 , n54149 , n54150 , 
 n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , 
 n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , 
 n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , 
 n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , 
 n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , 
 n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , 
 n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , 
 n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , 
 n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , n54239 , n54240 , 
 n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , 
 n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , 
 n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , n54267 , n54268 , n54269 , n54270 , 
 n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , n54277 , n54278 , n54279 , n54280 , 
 n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , n54287 , n54288 , n54289 , n54290 , 
 n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , n54297 , n54298 , n54299 , n54300 , 
 n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , n54307 , n54308 , n54309 , n54310 , 
 n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , n54317 , n54318 , n54319 , n54320 , 
 n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , n54327 , n54328 , n54329 , n54330 , 
 n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , n54337 , n54338 , n54339 , n54340 , 
 n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , n54347 , n54348 , n54349 , n54350 , 
 n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , n54357 , n54358 , n54359 , n54360 , 
 n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , n54367 , n54368 , n54369 , n54370 , 
 n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , n54377 , n54378 , n54379 , n54380 , 
 n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , n54387 , n54388 , n54389 , n54390 , 
 n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , n54397 , n54398 , n54399 , n54400 , 
 n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , n54407 , n54408 , n54409 , n54410 , 
 n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , n54417 , n54418 , n54419 , n54420 , 
 n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , n54427 , n54428 , n54429 , n54430 , 
 n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , n54437 , n54438 , n54439 , n54440 , 
 n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , n54447 , n54448 , n54449 , n54450 , 
 n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , n54457 , n54458 , n54459 , n54460 , 
 n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , n54467 , n54468 , n54469 , n54470 , 
 n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , n54477 , n54478 , n54479 , n54480 , 
 n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , n54487 , n54488 , n54489 , n54490 , 
 n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , n54497 , n54498 , n54499 , n54500 , 
 n54501 , n54502 , n54503 , n54504 , n54505 , n54506 , n54507 , n54508 , n54509 , n54510 , 
 n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , n54517 , n54518 , n54519 , n54520 , 
 n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , n54527 , n54528 , n54529 , n54530 , 
 n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , n54537 , n54538 , n54539 , n54540 , 
 n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , n54547 , n54548 , n54549 , n54550 , 
 n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , n54557 , n54558 , n54559 , n54560 , 
 n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , n54567 , n54568 , n54569 , n54570 , 
 n54571 , n54572 , n54573 , n54574 , n54575 , n54576 , n54577 , n54578 , n54579 , n54580 , 
 n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , n54587 , n54588 , n54589 , n54590 , 
 n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , 
 n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , n54607 , n54608 , n54609 , n54610 , 
 n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , n54617 , n54618 , n54619 , n54620 , 
 n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , n54627 , n54628 , n54629 , n54630 , 
 n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , n54637 , n54638 , n54639 , n54640 , 
 n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , n54647 , n54648 , n54649 , n54650 , 
 n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , n54657 , n54658 , n54659 , n54660 , 
 n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , n54667 , n54668 , n54669 , n54670 , 
 n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , n54677 , n54678 , n54679 , n54680 , 
 n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , n54687 , n54688 , n54689 , n54690 , 
 n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , n54697 , n54698 , n54699 , n54700 , 
 n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , n54707 , n54708 , n54709 , n54710 , 
 n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , n54717 , n54718 , n54719 , n54720 , 
 n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , n54727 , n54728 , n54729 , n54730 , 
 n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , n54737 , n54738 , n54739 , n54740 , 
 n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , 
 n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , n54757 , n54758 , n54759 , n54760 , 
 n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , n54767 , n54768 , n54769 , n54770 , 
 n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , n54777 , n54778 , n54779 , n54780 , 
 n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , 
 n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , n54797 , n54798 , n54799 , n54800 , 
 n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , n54807 , n54808 , n54809 , n54810 , 
 n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , n54817 , n54818 , n54819 , n54820 , 
 n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , n54827 , n54828 , n54829 , n54830 , 
 n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , n54837 , n54838 , n54839 , n54840 , 
 n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , n54847 , n54848 , n54849 , n54850 , 
 n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , n54857 , n54858 , n54859 , n54860 , 
 n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , n54867 , n54868 , n54869 , n54870 , 
 n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , n54877 , n54878 , n54879 , n54880 , 
 n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , n54887 , n54888 , n54889 , n54890 , 
 n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , n54897 , n54898 , n54899 , n54900 , 
 n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , n54907 , n54908 , n54909 , n54910 , 
 n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , n54917 , n54918 , n54919 , n54920 , 
 n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , n54927 , n54928 , n54929 , n54930 , 
 n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , n54937 , n54938 , n54939 , n54940 , 
 n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , n54947 , n54948 , n54949 , n54950 , 
 n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , n54957 , n54958 , n54959 , n54960 , 
 n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , n54967 , n54968 , n54969 , n54970 , 
 n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , n54977 , n54978 , n54979 , n54980 , 
 n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , n54987 , n54988 , n54989 , n54990 , 
 n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , 
 n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , 
 n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , n55017 , n55018 , n55019 , n55020 , 
 n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , n55027 , n55028 , n55029 , n55030 , 
 n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , n55037 , n55038 , n55039 , n55040 , 
 n55041 , n55042 , n55043 , n55044 , n55045 , n55046 , n55047 , n55048 , n55049 , n55050 , 
 n55051 , n55052 , n55053 , n55054 , n55055 , n55056 , n55057 , n55058 , n55059 , n55060 , 
 n55061 , n55062 , n55063 , n55064 , n55065 , n55066 , n55067 , n55068 , n55069 , n55070 , 
 n55071 , n55072 , n55073 , n55074 , n55075 , n55076 , n55077 , n55078 , n55079 , n55080 , 
 n55081 , n55082 , n55083 , n55084 , n55085 , n55086 , n55087 , n55088 , n55089 , n55090 , 
 n55091 , n55092 , n55093 , n55094 , n55095 , n55096 , n55097 , n55098 , n55099 , n55100 , 
 n55101 , n55102 , n55103 , n55104 , n55105 , n55106 , n55107 , n55108 , n55109 , n55110 , 
 n55111 , n55112 , n55113 , n55114 , n55115 , n55116 , n55117 , n55118 , n55119 , n55120 , 
 n55121 , n55122 , n55123 , n55124 , n55125 , n55126 , n55127 , n55128 , n55129 , n55130 , 
 n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , n55137 , n55138 , n55139 , n55140 , 
 n55141 , n55142 , n55143 , n55144 , n55145 , n55146 , n55147 , n55148 , n55149 , n55150 , 
 n55151 , n55152 , n55153 , n55154 , n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , 
 n55161 , n55162 , n55163 , n55164 , n55165 , n55166 , n55167 , n55168 , n55169 , n55170 , 
 n55171 , n55172 , n55173 , n55174 , n55175 , n55176 , n55177 , n55178 , n55179 , n55180 , 
 n55181 , n55182 , n55183 , n55184 , n55185 , n55186 , n55187 , n55188 , n55189 , n55190 , 
 n55191 , n55192 , n55193 , n55194 , n55195 , n55196 , n55197 , n55198 , n55199 , n55200 , 
 n55201 , n55202 , n55203 , n55204 , n55205 , n55206 , n55207 , n55208 , n55209 , n55210 , 
 n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , n55217 , n55218 , n55219 , n55220 , 
 n55221 , n55222 , n55223 , n55224 , n55225 , n55226 , n55227 , n55228 , n55229 , n55230 , 
 n55231 , n55232 , n55233 , n55234 , n55235 , n55236 , n55237 , n55238 , n55239 , n55240 , 
 n55241 , n55242 , n55243 , n55244 , n55245 , n55246 , n55247 , n55248 , n55249 , n55250 , 
 n55251 , n55252 , n55253 , n55254 , n55255 , n55256 , n55257 , n55258 , n55259 , n55260 , 
 n55261 , n55262 , n55263 , n55264 , n55265 , n55266 , n55267 , n55268 , n55269 , n55270 , 
 n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , n55277 , n55278 , n55279 , n55280 , 
 n55281 , n55282 , n55283 , n55284 , n55285 , n55286 , n55287 , n55288 , n55289 , n55290 , 
 n55291 , n55292 , n55293 , n55294 , n55295 , n55296 , n55297 , n55298 , n55299 , n55300 , 
 n55301 , n55302 , n55303 , n55304 , n55305 , n55306 , n55307 , n55308 , n55309 , n55310 , 
 n55311 , n55312 , n55313 , n55314 , n55315 , n55316 , n55317 , n55318 , n55319 , n55320 , 
 n55321 , n55322 , n55323 , n55324 , n55325 , n55326 , n55327 , n55328 , n55329 , n55330 , 
 n55331 , n55332 , n55333 , n55334 , n55335 , n55336 , n55337 , n55338 , n55339 , n55340 , 
 n55341 , n55342 , n55343 , n55344 , n55345 , n55346 , n55347 , n55348 , n55349 , n55350 , 
 n55351 , n55352 , n55353 , n55354 , n55355 , n55356 , n55357 , n55358 , n55359 , n55360 , 
 n55361 , n55362 , n55363 , n55364 , n55365 , n55366 , n55367 , n55368 , n55369 , n55370 , 
 n55371 , n55372 , n55373 , n55374 , n55375 , n55376 , n55377 , n55378 , n55379 , n55380 , 
 n55381 , n55382 , n55383 , n55384 , n55385 , n55386 , n55387 , n55388 , n55389 , n55390 , 
 n55391 , n55392 , n55393 , n55394 , n55395 , n55396 , n55397 , n55398 , n55399 , n55400 , 
 n55401 , n55402 , n55403 , n55404 , n55405 , n55406 , n55407 , n55408 , n55409 , n55410 , 
 n55411 , n55412 , n55413 , n55414 , n55415 , n55416 , n55417 , n55418 , n55419 , n55420 , 
 n55421 , n55422 , n55423 , n55424 , n55425 , n55426 , n55427 , n55428 , n55429 , n55430 , 
 n55431 , n55432 , n55433 , n55434 , n55435 , n55436 , n55437 , n55438 , n55439 , n55440 , 
 n55441 , n55442 , n55443 , n55444 , n55445 , n55446 , n55447 , n55448 , n55449 , n55450 , 
 n55451 , n55452 , n55453 , n55454 , n55455 , n55456 , n55457 , n55458 , n55459 , n55460 , 
 n55461 , n55462 , n55463 , n55464 , n55465 , n55466 , n55467 , n55468 , n55469 , n55470 , 
 n55471 , n55472 , n55473 , n55474 , n55475 , n55476 , n55477 , n55478 , n55479 , n55480 , 
 n55481 , n55482 , n55483 , n55484 , n55485 , n55486 , n55487 , n55488 , n55489 , n55490 , 
 n55491 , n55492 , n55493 , n55494 , n55495 , n55496 , n55497 , n55498 , n55499 , n55500 , 
 n55501 , n55502 , n55503 , n55504 , n55505 , n55506 , n55507 , n55508 , n55509 , n55510 , 
 n55511 , n55512 , n55513 , n55514 , n55515 , n55516 , n55517 , n55518 , n55519 , n55520 , 
 n55521 , n55522 , n55523 , n55524 , n55525 , n55526 , n55527 , n55528 , n55529 , n55530 , 
 n55531 , n55532 , n55533 , n55534 , n55535 , n55536 , n55537 , n55538 , n55539 , n55540 , 
 n55541 , n55542 , n55543 , n55544 , n55545 , n55546 , n55547 , n55548 , n55549 , n55550 , 
 n55551 , n55552 , n55553 , n55554 , n55555 , n55556 , n55557 , n55558 , n55559 , n55560 , 
 n55561 , n55562 , n55563 , n55564 , n55565 , n55566 , n55567 , n55568 , n55569 , n55570 , 
 n55571 , n55572 , n55573 , n55574 , n55575 , n55576 , n55577 , n55578 , n55579 , n55580 , 
 n55581 , n55582 , n55583 , n55584 , n55585 , n55586 , n55587 , n55588 , n55589 , n55590 , 
 n55591 , n55592 , n55593 , n55594 , n55595 , n55596 , n55597 , n55598 , n55599 , n55600 , 
 n55601 , n55602 , n55603 , n55604 , n55605 , n55606 , n55607 , n55608 , n55609 , n55610 , 
 n55611 , n55612 , n55613 , n55614 , n55615 , n55616 , n55617 , n55618 , n55619 , n55620 , 
 n55621 , n55622 , n55623 , n55624 , n55625 , n55626 , n55627 , n55628 , n55629 , n55630 , 
 n55631 , n55632 , n55633 , n55634 , n55635 , n55636 , n55637 , n55638 , n55639 , n55640 , 
 n55641 , n55642 , n55643 , n55644 , n55645 , n55646 , n55647 , n55648 , n55649 , n55650 , 
 n55651 , n55652 , n55653 , n55654 , n55655 , n55656 , n55657 , n55658 , n55659 , n55660 , 
 n55661 , n55662 , n55663 , n55664 , n55665 , n55666 , n55667 , n55668 , n55669 , n55670 , 
 n55671 , n55672 , n55673 , n55674 , n55675 , n55676 , n55677 , n55678 , n55679 , n55680 , 
 n55681 , n55682 , n55683 , n55684 , n55685 , n55686 , n55687 , n55688 , n55689 , n55690 , 
 n55691 , n55692 , n55693 , n55694 , n55695 , n55696 , n55697 , n55698 , n55699 , n55700 , 
 n55701 , n55702 , n55703 , n55704 , n55705 , n55706 , n55707 , n55708 , n55709 , n55710 , 
 n55711 , n55712 , n55713 , n55714 , n55715 , n55716 , n55717 , n55718 , n55719 , n55720 , 
 n55721 , n55722 , n55723 , n55724 , n55725 , n55726 , n55727 , n55728 , n55729 , n55730 , 
 n55731 , n55732 , n55733 , n55734 , n55735 , n55736 , n55737 , n55738 , n55739 , n55740 , 
 n55741 , n55742 , n55743 , n55744 , n55745 , n55746 , n55747 , n55748 , n55749 , n55750 , 
 n55751 , n55752 , n55753 , n55754 , n55755 , n55756 , n55757 , n55758 , n55759 , n55760 , 
 n55761 , n55762 , n55763 , n55764 , n55765 , n55766 , n55767 , n55768 , n55769 , n55770 , 
 n55771 , n55772 , n55773 , n55774 , n55775 , n55776 , n55777 , n55778 , n55779 , n55780 , 
 n55781 , n55782 , n55783 , n55784 , n55785 , n55786 , n55787 , n55788 , n55789 , n55790 , 
 n55791 , n55792 , n55793 , n55794 , n55795 , n55796 , n55797 , n55798 , n55799 , n55800 , 
 n55801 , n55802 , n55803 , n55804 , n55805 , n55806 , n55807 , n55808 , n55809 , n55810 , 
 n55811 , n55812 , n55813 , n55814 , n55815 , n55816 , n55817 , n55818 , n55819 , n55820 , 
 n55821 , n55822 , n55823 , n55824 , n55825 , n55826 , n55827 , n55828 , n55829 , n55830 , 
 n55831 , n55832 , n55833 , n55834 , n55835 , n55836 , n55837 , n55838 , n55839 , n55840 , 
 n55841 , n55842 , n55843 , n55844 , n55845 , n55846 , n55847 , n55848 , n55849 , n55850 , 
 n55851 , n55852 , n55853 , n55854 , n55855 , n55856 , n55857 , n55858 , n55859 , n55860 , 
 n55861 , n55862 , n55863 , n55864 , n55865 , n55866 , n55867 , n55868 , n55869 , n55870 , 
 n55871 , n55872 , n55873 , n55874 , n55875 , n55876 , n55877 , n55878 , n55879 , n55880 , 
 n55881 , n55882 , n55883 , n55884 , n55885 , n55886 , n55887 , n55888 , n55889 , n55890 , 
 n55891 , n55892 , n55893 , n55894 , n55895 , n55896 , n55897 , n55898 , n55899 , n55900 , 
 n55901 , n55902 , n55903 , n55904 , n55905 , n55906 , n55907 , n55908 , n55909 , n55910 , 
 n55911 , n55912 , n55913 , n55914 , n55915 , n55916 , n55917 , n55918 , n55919 , n55920 , 
 n55921 , n55922 , n55923 , n55924 , n55925 , n55926 , n55927 , n55928 , n55929 , n55930 , 
 n55931 , n55932 , n55933 , n55934 , n55935 , n55936 , n55937 , n55938 , n55939 , n55940 , 
 n55941 , n55942 , n55943 , n55944 , n55945 , n55946 , n55947 , n55948 , n55949 , n55950 , 
 n55951 , n55952 , n55953 , n55954 , n55955 , n55956 , n55957 , n55958 , n55959 , n55960 , 
 n55961 , n55962 , n55963 , n55964 , n55965 , n55966 , n55967 , n55968 , n55969 , n55970 , 
 n55971 , n55972 , n55973 , n55974 , n55975 , n55976 , n55977 , n55978 , n55979 , n55980 , 
 n55981 , n55982 , n55983 , n55984 , n55985 , n55986 , n55987 , n55988 , n55989 , n55990 , 
 n55991 , n55992 , n55993 , n55994 , n55995 , n55996 , n55997 , n55998 , n55999 , n56000 , 
 n56001 , n56002 , n56003 , n56004 , n56005 , n56006 , n56007 , n56008 , n56009 , n56010 , 
 n56011 , n56012 , n56013 , n56014 , n56015 , n56016 , n56017 , n56018 , n56019 , n56020 , 
 n56021 , n56022 , n56023 , n56024 , n56025 , n56026 , n56027 , n56028 , n56029 , n56030 , 
 n56031 , n56032 , n56033 , n56034 , n56035 , n56036 , n56037 , n56038 , n56039 , n56040 , 
 n56041 , n56042 , n56043 , n56044 , n56045 , n56046 , n56047 , n56048 , n56049 , n56050 , 
 n56051 , n56052 , n56053 , n56054 , n56055 , n56056 , n56057 , n56058 , n56059 , n56060 , 
 n56061 , n56062 , n56063 , n56064 , n56065 , n56066 , n56067 , n56068 , n56069 , n56070 , 
 n56071 , n56072 , n56073 , n56074 , n56075 , n56076 , n56077 , n56078 , n56079 , n56080 , 
 n56081 , n56082 , n56083 , n56084 , n56085 , n56086 , n56087 , n56088 , n56089 , n56090 , 
 n56091 , n56092 , n56093 , n56094 , n56095 , n56096 , n56097 , n56098 , n56099 , n56100 , 
 n56101 , n56102 , n56103 , n56104 , n56105 , n56106 , n56107 , n56108 , n56109 , n56110 , 
 n56111 , n56112 , n56113 , n56114 , n56115 , n56116 , n56117 , n56118 , n56119 , n56120 , 
 n56121 , n56122 , n56123 , n56124 , n56125 , n56126 , n56127 , n56128 , n56129 , n56130 , 
 n56131 , n56132 , n56133 , n56134 , n56135 , n56136 , n56137 , n56138 , n56139 , n56140 , 
 n56141 , n56142 , n56143 , n56144 , n56145 , n56146 , n56147 , n56148 , n56149 , n56150 , 
 n56151 , n56152 , n56153 , n56154 , n56155 , n56156 , n56157 , n56158 , n56159 , n56160 , 
 n56161 , n56162 , n56163 , n56164 , n56165 , n56166 , n56167 , n56168 , n56169 , n56170 , 
 n56171 , n56172 , n56173 , n56174 , n56175 , n56176 , n56177 , n56178 , n56179 , n56180 , 
 n56181 , n56182 , n56183 , n56184 , n56185 , n56186 , n56187 , n56188 , n56189 , n56190 , 
 n56191 , n56192 , n56193 , n56194 , n56195 , n56196 , n56197 , n56198 , n56199 , n56200 , 
 n56201 , n56202 , n56203 , n56204 , n56205 , n56206 , n56207 , n56208 , n56209 , n56210 , 
 n56211 , n56212 , n56213 , n56214 , n56215 , n56216 , n56217 , n56218 , n56219 , n56220 , 
 n56221 , n56222 , n56223 , n56224 , n56225 , n56226 , n56227 , n56228 , n56229 , n56230 , 
 n56231 , n56232 , n56233 , n56234 , n56235 , n56236 , n56237 , n56238 , n56239 , n56240 , 
 n56241 , n56242 , n56243 , n56244 , n56245 , n56246 , n56247 , n56248 , n56249 , n56250 , 
 n56251 , n56252 , n56253 , n56254 , n56255 , n56256 , n56257 , n56258 , n56259 , n56260 , 
 n56261 , n56262 , n56263 , n56264 , n56265 , n56266 , n56267 , n56268 , n56269 , n56270 , 
 n56271 , n56272 , n56273 , n56274 , n56275 , n56276 , n56277 , n56278 , n56279 , n56280 , 
 n56281 , n56282 , n56283 , n56284 , n56285 , n56286 , n56287 , n56288 , n56289 , n56290 , 
 n56291 , n56292 , n56293 , n56294 , n56295 , n56296 , n56297 , n56298 , n56299 , n56300 , 
 n56301 , n56302 , n56303 , n56304 , n56305 , n56306 , n56307 , n56308 , n56309 , n56310 , 
 n56311 , n56312 , n56313 , n56314 , n56315 , n56316 , n56317 , n56318 , n56319 , n56320 , 
 n56321 , n56322 , n56323 , n56324 , n56325 , n56326 , n56327 , n56328 , n56329 , n56330 , 
 n56331 , n56332 , n56333 , n56334 , n56335 , n56336 , n56337 , n56338 , n56339 , n56340 , 
 n56341 , n56342 , n56343 , n56344 , n56345 , n56346 , n56347 , n56348 , n56349 , n56350 , 
 n56351 , n56352 , n56353 , n56354 , n56355 , n56356 , n56357 , n56358 , n56359 , n56360 , 
 n56361 , n56362 , n56363 , n56364 , n56365 , n56366 , n56367 , n56368 , n56369 , n56370 , 
 n56371 , n56372 , n56373 , n56374 , n56375 , n56376 , n56377 , n56378 , n56379 , n56380 , 
 n56381 , n56382 , n56383 , n56384 , n56385 , n56386 , n56387 , n56388 , n56389 , n56390 , 
 n56391 , n56392 , n56393 , n56394 , n56395 , n56396 , n56397 , n56398 , n56399 , n56400 , 
 n56401 , n56402 , n56403 , n56404 , n56405 , n56406 , n56407 , n56408 , n56409 , n56410 , 
 n56411 , n56412 , n56413 , n56414 , n56415 , n56416 , n56417 , n56418 , n56419 , n56420 , 
 n56421 , n56422 , n56423 , n56424 , n56425 , n56426 , n56427 , n56428 , n56429 , n56430 , 
 n56431 , n56432 , n56433 , n56434 , n56435 , n56436 , n56437 , n56438 , n56439 , n56440 , 
 n56441 , n56442 , n56443 , n56444 , n56445 , n56446 , n56447 , n56448 , n56449 , n56450 , 
 n56451 , n56452 , n56453 , n56454 , n56455 , n56456 , n56457 , n56458 , n56459 , n56460 , 
 n56461 , n56462 , n56463 , n56464 , n56465 , n56466 , n56467 , n56468 , n56469 , n56470 , 
 n56471 , n56472 , n56473 , n56474 , n56475 , n56476 , n56477 , n56478 , n56479 , n56480 , 
 n56481 , n56482 , n56483 , n56484 , n56485 , n56486 , n56487 , n56488 , n56489 , n56490 , 
 n56491 , n56492 , n56493 , n56494 , n56495 , n56496 , n56497 , n56498 , n56499 , n56500 , 
 n56501 , n56502 , n56503 , n56504 , n56505 , n56506 , n56507 , n56508 , n56509 , n56510 , 
 n56511 , n56512 , n56513 , n56514 , n56515 , n56516 , n56517 , n56518 , n56519 , n56520 , 
 n56521 , n56522 , n56523 , n56524 , n56525 , n56526 , n56527 , n56528 , n56529 , n56530 , 
 n56531 , n56532 , n56533 , n56534 , n56535 , n56536 , n56537 , n56538 , n56539 , n56540 , 
 n56541 , n56542 , n56543 , n56544 , n56545 , n56546 , n56547 , n56548 , n56549 , n56550 , 
 n56551 , n56552 , n56553 , n56554 , n56555 , n56556 , n56557 , n56558 , n56559 , n56560 , 
 n56561 , n56562 , n56563 , n56564 , n56565 , n56566 , n56567 , n56568 , n56569 , n56570 , 
 n56571 , n56572 , n56573 , n56574 , n56575 , n56576 , n56577 , n56578 , n56579 , n56580 , 
 n56581 , n56582 , n56583 , n56584 , n56585 , n56586 , n56587 , n56588 , n56589 , n56590 , 
 n56591 , n56592 , n56593 , n56594 , n56595 , n56596 , n56597 , n56598 , n56599 , n56600 , 
 n56601 , n56602 , n56603 , n56604 , n56605 , n56606 , n56607 , n56608 , n56609 , n56610 , 
 n56611 , n56612 , n56613 , n56614 , n56615 , n56616 , n56617 , n56618 , n56619 , n56620 , 
 n56621 , n56622 , n56623 , n56624 , n56625 , n56626 , n56627 , n56628 , n56629 , n56630 , 
 n56631 , n56632 , n56633 , n56634 , n56635 , n56636 , n56637 , n56638 , n56639 , n56640 , 
 n56641 , n56642 , n56643 , n56644 , n56645 , n56646 , n56647 , n56648 , n56649 , n56650 , 
 n56651 , n56652 , n56653 , n56654 , n56655 , n56656 , n56657 , n56658 , n56659 , n56660 , 
 n56661 , n56662 , n56663 , n56664 , n56665 , n56666 , n56667 , n56668 , n56669 , n56670 , 
 n56671 , n56672 , n56673 , n56674 , n56675 , n56676 , n56677 , n56678 , n56679 , n56680 , 
 n56681 , n56682 , n56683 , n56684 , n56685 , n56686 , n56687 , n56688 , n56689 , n56690 , 
 n56691 , n56692 , n56693 , n56694 , n56695 , n56696 , n56697 , n56698 , n56699 , n56700 , 
 n56701 , n56702 , n56703 , n56704 , n56705 , n56706 , n56707 , n56708 , n56709 , n56710 , 
 n56711 , n56712 , n56713 , n56714 , n56715 , n56716 , n56717 , n56718 , n56719 , n56720 , 
 n56721 , n56722 , n56723 , n56724 , n56725 , n56726 , n56727 , n56728 , n56729 , n56730 , 
 n56731 , n56732 , n56733 , n56734 , n56735 , n56736 , n56737 , n56738 , n56739 , n56740 , 
 n56741 , n56742 , n56743 , n56744 , n56745 , n56746 , n56747 , n56748 , n56749 , n56750 , 
 n56751 , n56752 , n56753 , n56754 , n56755 , n56756 , n56757 , n56758 , n56759 , n56760 , 
 n56761 , n56762 , n56763 , n56764 , n56765 , n56766 , n56767 , n56768 , n56769 , n56770 , 
 n56771 , n56772 , n56773 , n56774 , n56775 , n56776 , n56777 , n56778 , n56779 , n56780 , 
 n56781 , n56782 , n56783 , n56784 , n56785 , n56786 , n56787 , n56788 , n56789 , n56790 , 
 n56791 , n56792 , n56793 , n56794 , n56795 , n56796 , n56797 , n56798 , n56799 , n56800 , 
 n56801 , n56802 , n56803 , n56804 , n56805 , n56806 , n56807 , n56808 , n56809 , n56810 , 
 n56811 , n56812 , n56813 , n56814 , n56815 , n56816 , n56817 , n56818 , n56819 , n56820 , 
 n56821 , n56822 , n56823 , n56824 , n56825 , n56826 , n56827 , n56828 , n56829 , n56830 , 
 n56831 , n56832 , n56833 , n56834 , n56835 , n56836 , n56837 , n56838 , n56839 , n56840 , 
 n56841 , n56842 , n56843 , n56844 , n56845 , n56846 , n56847 , n56848 , n56849 , n56850 , 
 n56851 , n56852 , n56853 , n56854 , n56855 , n56856 , n56857 , n56858 , n56859 , n56860 , 
 n56861 , n56862 , n56863 , n56864 , n56865 , n56866 , n56867 , n56868 , n56869 , n56870 , 
 n56871 , n56872 , n56873 , n56874 , n56875 , n56876 , n56877 , n56878 , n56879 , n56880 , 
 n56881 , n56882 , n56883 , n56884 , n56885 , n56886 , n56887 , n56888 , n56889 , n56890 , 
 n56891 , n56892 , n56893 , n56894 , n56895 , n56896 , n56897 , n56898 , n56899 , n56900 , 
 n56901 , n56902 , n56903 , n56904 , n56905 , n56906 , n56907 , n56908 , n56909 , n56910 , 
 n56911 , n56912 , n56913 , n56914 , n56915 , n56916 , n56917 , n56918 , n56919 , n56920 , 
 n56921 , n56922 , n56923 , n56924 , n56925 , n56926 , n56927 , n56928 , n56929 , n56930 , 
 n56931 , n56932 , n56933 , n56934 , n56935 , n56936 , n56937 , n56938 , n56939 , n56940 , 
 n56941 , n56942 , n56943 , n56944 , n56945 , n56946 , n56947 , n56948 , n56949 , n56950 , 
 n56951 , n56952 , n56953 , n56954 , n56955 , n56956 , n56957 , n56958 , n56959 , n56960 , 
 n56961 , n56962 , n56963 , n56964 , n56965 , n56966 , n56967 , n56968 , n56969 , n56970 , 
 n56971 , n56972 , n56973 , n56974 , n56975 , n56976 , n56977 , n56978 , n56979 , n56980 , 
 n56981 , n56982 , n56983 , n56984 , n56985 , n56986 , n56987 , n56988 , n56989 , n56990 , 
 n56991 , n56992 , n56993 , n56994 , n56995 , n56996 , n56997 , n56998 , n56999 , n57000 , 
 n57001 , n57002 , n57003 , n57004 , n57005 , n57006 , n57007 , n57008 , n57009 , n57010 , 
 n57011 , n57012 , n57013 , n57014 , n57015 , n57016 , n57017 , n57018 , n57019 , n57020 , 
 n57021 , n57022 , n57023 , n57024 , n57025 , n57026 , n57027 , n57028 , n57029 , n57030 , 
 n57031 , n57032 , n57033 , n57034 , n57035 , n57036 , n57037 , n57038 , n57039 , n57040 , 
 n57041 , n57042 , n57043 , n57044 , n57045 , n57046 , n57047 , n57048 , n57049 , n57050 , 
 n57051 , n57052 , n57053 , n57054 , n57055 , n57056 , n57057 , n57058 , n57059 , n57060 , 
 n57061 , n57062 , n57063 , n57064 , n57065 , n57066 , n57067 , n57068 , n57069 , n57070 , 
 n57071 , n57072 , n57073 , n57074 , n57075 , n57076 , n57077 , n57078 , n57079 , n57080 , 
 n57081 , n57082 , n57083 , n57084 , n57085 , n57086 , n57087 , n57088 , n57089 , n57090 , 
 n57091 , n57092 , n57093 , n57094 , n57095 , n57096 , n57097 , n57098 , n57099 , n57100 , 
 n57101 , n57102 , n57103 , n57104 , n57105 , n57106 , n57107 , n57108 , n57109 , n57110 , 
 n57111 , n57112 , n57113 , n57114 , n57115 , n57116 , n57117 , n57118 , n57119 , n57120 , 
 n57121 , n57122 , n57123 , n57124 , n57125 , n57126 , n57127 , n57128 , n57129 , n57130 , 
 n57131 , n57132 , n57133 , n57134 , n57135 , n57136 , n57137 , n57138 , n57139 , n57140 , 
 n57141 , n57142 , n57143 , n57144 , n57145 , n57146 , n57147 , n57148 , n57149 , n57150 , 
 n57151 , n57152 , n57153 , n57154 , n57155 , n57156 , n57157 , n57158 , n57159 , n57160 , 
 n57161 , n57162 , n57163 , n57164 , n57165 , n57166 , n57167 , n57168 , n57169 , n57170 , 
 n57171 , n57172 , n57173 , n57174 , n57175 , n57176 , n57177 , n57178 , n57179 , n57180 , 
 n57181 , n57182 , n57183 , n57184 , n57185 , n57186 , n57187 , n57188 , n57189 , n57190 , 
 n57191 , n57192 , n57193 , n57194 , n57195 , n57196 , n57197 , n57198 , n57199 , n57200 , 
 n57201 , n57202 , n57203 , n57204 , n57205 , n57206 , n57207 , n57208 , n57209 , n57210 , 
 n57211 , n57212 , n57213 , n57214 , n57215 , n57216 , n57217 , n57218 , n57219 , n57220 , 
 n57221 , n57222 , n57223 , n57224 , n57225 , n57226 , n57227 , n57228 , n57229 , n57230 , 
 n57231 , n57232 , n57233 , n57234 , n57235 , n57236 , n57237 , n57238 , n57239 , n57240 , 
 n57241 , n57242 , n57243 , n57244 , n57245 , n57246 , n57247 , n57248 , n57249 , n57250 , 
 n57251 , n57252 , n57253 , n57254 , n57255 , n57256 , n57257 , n57258 , n57259 , n57260 , 
 n57261 , n57262 , n57263 , n57264 , n57265 , n57266 , n57267 , n57268 , n57269 , n57270 , 
 n57271 , n57272 , n57273 , n57274 , n57275 , n57276 , n57277 , n57278 , n57279 , n57280 , 
 n57281 , n57282 , n57283 , n57284 , n57285 , n57286 , n57287 , n57288 , n57289 , n57290 , 
 n57291 , n57292 , n57293 , n57294 , n57295 , n57296 , n57297 , n57298 , n57299 , n57300 , 
 n57301 , n57302 , n57303 , n57304 , n57305 , n57306 , n57307 , n57308 , n57309 , n57310 , 
 n57311 , n57312 , n57313 , n57314 , n57315 , n57316 , n57317 , n57318 , n57319 , n57320 , 
 n57321 , n57322 , n57323 , n57324 , n57325 , n57326 , n57327 , n57328 , n57329 , n57330 , 
 n57331 , n57332 , n57333 , n57334 , n57335 , n57336 , n57337 , n57338 , n57339 , n57340 , 
 n57341 , n57342 , n57343 , n57344 , n57345 , n57346 , n57347 , n57348 , n57349 , n57350 , 
 n57351 , n57352 , n57353 , n57354 , n57355 , n57356 , n57357 , n57358 , n57359 , n57360 , 
 n57361 , n57362 , n57363 , n57364 , n57365 , n57366 , n57367 , n57368 , n57369 , n57370 , 
 n57371 , n57372 , n57373 , n57374 , n57375 , n57376 , n57377 , n57378 , n57379 , n57380 , 
 n57381 , n57382 , n57383 , n57384 , n57385 , n57386 , n57387 , n57388 , n57389 , n57390 , 
 n57391 , n57392 , n57393 , n57394 , n57395 , n57396 , n57397 , n57398 , n57399 , n57400 , 
 n57401 , n57402 , n57403 , n57404 , n57405 , n57406 , n57407 , n57408 , n57409 , n57410 , 
 n57411 , n57412 , n57413 , n57414 , n57415 , n57416 , n57417 , n57418 , n57419 , n57420 , 
 n57421 , n57422 , n57423 , n57424 , n57425 , n57426 , n57427 , n57428 , n57429 , n57430 , 
 n57431 , n57432 , n57433 , n57434 , n57435 , n57436 , n57437 , n57438 , n57439 , n57440 , 
 n57441 , n57442 , n57443 , n57444 , n57445 , n57446 , n57447 , n57448 , n57449 , n57450 , 
 n57451 , n57452 , n57453 , n57454 , n57455 , n57456 , n57457 , n57458 , n57459 , n57460 , 
 n57461 , n57462 , n57463 , n57464 , n57465 , n57466 , n57467 , n57468 , n57469 , n57470 , 
 n57471 , n57472 , n57473 , n57474 , n57475 , n57476 , n57477 , n57478 , n57479 , n57480 , 
 n57481 , n57482 , n57483 , n57484 , n57485 , n57486 , n57487 , n57488 , n57489 , n57490 , 
 n57491 , n57492 , n57493 , n57494 , n57495 , n57496 , n57497 , n57498 , n57499 , n57500 , 
 n57501 , n57502 , n57503 , n57504 , n57505 , n57506 , n57507 , n57508 , n57509 , n57510 , 
 n57511 , n57512 , n57513 , n57514 , n57515 , n57516 , n57517 , n57518 , n57519 , n57520 , 
 n57521 , n57522 , n57523 , n57524 , n57525 , n57526 , n57527 , n57528 , n57529 , n57530 , 
 n57531 , n57532 , n57533 , n57534 , n57535 , n57536 , n57537 , n57538 , n57539 , n57540 , 
 n57541 , n57542 , n57543 , n57544 , n57545 , n57546 , n57547 , n57548 , n57549 , n57550 , 
 n57551 , n57552 , n57553 , n57554 , n57555 , n57556 , n57557 , n57558 , n57559 , n57560 , 
 n57561 , n57562 , n57563 , n57564 , n57565 , n57566 , n57567 , n57568 , n57569 , n57570 , 
 n57571 , n57572 , n57573 , n57574 , n57575 , n57576 , n57577 , n57578 , n57579 , n57580 , 
 n57581 , n57582 , n57583 , n57584 , n57585 , n57586 , n57587 , n57588 , n57589 , n57590 , 
 n57591 , n57592 , n57593 , n57594 , n57595 , n57596 , n57597 , n57598 , n57599 , n57600 , 
 n57601 , n57602 , n57603 , n57604 , n57605 , n57606 , n57607 , n57608 , n57609 , n57610 , 
 n57611 , n57612 , n57613 , n57614 , n57615 , n57616 , n57617 , n57618 , n57619 , n57620 , 
 n57621 , n57622 , n57623 , n57624 , n57625 , n57626 , n57627 , n57628 , n57629 , n57630 , 
 n57631 , n57632 , n57633 , n57634 , n57635 , n57636 , n57637 , n57638 , n57639 , n57640 , 
 n57641 , n57642 , n57643 , n57644 , n57645 , n57646 , n57647 , n57648 , n57649 , n57650 , 
 n57651 , n57652 , n57653 , n57654 , n57655 , n57656 , n57657 , n57658 , n57659 , n57660 , 
 n57661 , n57662 , n57663 , n57664 , n57665 , n57666 , n57667 , n57668 , n57669 , n57670 , 
 n57671 , n57672 , n57673 , n57674 , n57675 , n57676 , n57677 , n57678 , n57679 , n57680 , 
 n57681 , n57682 , n57683 , n57684 , n57685 , n57686 , n57687 , n57688 , n57689 , n57690 , 
 n57691 , n57692 , n57693 , n57694 , n57695 , n57696 , n57697 , n57698 , n57699 , n57700 , 
 n57701 , n57702 , n57703 , n57704 , n57705 , n57706 , n57707 , n57708 , n57709 , n57710 , 
 n57711 , n57712 , n57713 , n57714 , n57715 , n57716 , n57717 , n57718 , n57719 , n57720 , 
 n57721 , n57722 , n57723 , n57724 , n57725 , n57726 , n57727 , n57728 , n57729 , n57730 , 
 n57731 , n57732 , n57733 , n57734 , n57735 , n57736 , n57737 , n57738 , n57739 , n57740 , 
 n57741 , n57742 , n57743 , n57744 , n57745 , n57746 , n57747 , n57748 , n57749 , n57750 , 
 n57751 , n57752 , n57753 , n57754 , n57755 , n57756 , n57757 , n57758 , n57759 , n57760 , 
 n57761 , n57762 , n57763 , n57764 , n57765 , n57766 , n57767 , n57768 , n57769 , n57770 , 
 n57771 , n57772 , n57773 , n57774 , n57775 , n57776 , n57777 , n57778 , n57779 , n57780 , 
 n57781 , n57782 , n57783 , n57784 , n57785 , n57786 , n57787 , n57788 , n57789 , n57790 , 
 n57791 , n57792 , n57793 , n57794 , n57795 , n57796 , n57797 , n57798 , n57799 , n57800 , 
 n57801 , n57802 , n57803 , n57804 , n57805 , n57806 , n57807 , n57808 , n57809 , n57810 , 
 n57811 , n57812 , n57813 , n57814 , n57815 , n57816 , n57817 , n57818 , n57819 , n57820 , 
 n57821 , n57822 , n57823 , n57824 , n57825 , n57826 , n57827 , n57828 , n57829 , n57830 , 
 n57831 , n57832 , n57833 , n57834 , n57835 , n57836 , n57837 , n57838 , n57839 , n57840 , 
 n57841 , n57842 , n57843 , n57844 , n57845 , n57846 , n57847 , n57848 , n57849 , n57850 , 
 n57851 , n57852 , n57853 , n57854 , n57855 , n57856 , n57857 , n57858 , n57859 , n57860 , 
 n57861 , n57862 , n57863 , n57864 , n57865 , n57866 , n57867 , n57868 , n57869 , n57870 , 
 n57871 , n57872 , n57873 , n57874 , n57875 , n57876 , n57877 , n57878 , n57879 , n57880 , 
 n57881 , n57882 , n57883 , n57884 , n57885 , n57886 , n57887 , n57888 , n57889 , n57890 , 
 n57891 , n57892 , n57893 , n57894 , n57895 , n57896 , n57897 , n57898 , n57899 , n57900 , 
 n57901 , n57902 , n57903 , n57904 , n57905 , n57906 , n57907 , n57908 , n57909 , n57910 , 
 n57911 , n57912 , n57913 , n57914 , n57915 , n57916 , n57917 , n57918 , n57919 , n57920 , 
 n57921 , n57922 , n57923 , n57924 , n57925 , n57926 , n57927 , n57928 , n57929 , n57930 , 
 n57931 , n57932 , n57933 , n57934 , n57935 , n57936 , n57937 , n57938 , n57939 , n57940 , 
 n57941 , n57942 , n57943 , n57944 , n57945 , n57946 , n57947 , n57948 , n57949 , n57950 , 
 n57951 , n57952 , n57953 , n57954 , n57955 , n57956 , n57957 , n57958 , n57959 , n57960 , 
 n57961 , n57962 , n57963 , n57964 , n57965 , n57966 , n57967 , n57968 , n57969 , n57970 , 
 n57971 , n57972 , n57973 , n57974 , n57975 , n57976 , n57977 , n57978 , n57979 , n57980 , 
 n57981 , n57982 , n57983 , n57984 , n57985 , n57986 , n57987 , n57988 , n57989 , n57990 , 
 n57991 , n57992 , n57993 , n57994 , n57995 , n57996 , n57997 , n57998 , n57999 , n58000 , 
 n58001 , n58002 , n58003 , n58004 , n58005 , n58006 , n58007 , n58008 , n58009 , n58010 , 
 n58011 , n58012 , n58013 , n58014 , n58015 , n58016 , n58017 , n58018 , n58019 , n58020 , 
 n58021 , n58022 , n58023 , n58024 , n58025 , n58026 , n58027 , n58028 , n58029 , n58030 , 
 n58031 , n58032 , n58033 , n58034 , n58035 , n58036 , n58037 , n58038 , n58039 , n58040 , 
 n58041 , n58042 , n58043 , n58044 , n58045 , n58046 , n58047 , n58048 , n58049 , n58050 , 
 n58051 , n58052 , n58053 , n58054 , n58055 , n58056 , n58057 , n58058 , n58059 , n58060 , 
 n58061 , n58062 , n58063 , n58064 , n58065 , n58066 , n58067 , n58068 , n58069 , n58070 , 
 n58071 , n58072 , n58073 , n58074 , n58075 , n58076 , n58077 , n58078 , n58079 , n58080 , 
 n58081 , n58082 , n58083 , n58084 , n58085 , n58086 , n58087 , n58088 , n58089 , n58090 , 
 n58091 , n58092 , n58093 , n58094 , n58095 , n58096 , n58097 , n58098 , n58099 , n58100 , 
 n58101 , n58102 , n58103 , n58104 , n58105 , n58106 , n58107 , n58108 , n58109 , n58110 , 
 n58111 , n58112 , n58113 , n58114 , n58115 , n58116 , n58117 , n58118 , n58119 , n58120 , 
 n58121 , n58122 , n58123 , n58124 , n58125 , n58126 , n58127 , n58128 , n58129 , n58130 , 
 n58131 , n58132 , n58133 , n58134 , n58135 , n58136 , n58137 , n58138 , n58139 , n58140 , 
 n58141 , n58142 , n58143 , n58144 , n58145 , n58146 , n58147 , n58148 , n58149 , n58150 , 
 n58151 , n58152 , n58153 , n58154 , n58155 , n58156 , n58157 , n58158 , n58159 , n58160 , 
 n58161 , n58162 , n58163 , n58164 , n58165 , n58166 , n58167 , n58168 , n58169 , n58170 , 
 n58171 , n58172 , n58173 , n58174 , n58175 , n58176 , n58177 , n58178 , n58179 , n58180 , 
 n58181 , n58182 , n58183 , n58184 , n58185 , n58186 , n58187 , n58188 , n58189 , n58190 , 
 n58191 , n58192 , n58193 , n58194 , n58195 , n58196 , n58197 , n58198 , n58199 , n58200 , 
 n58201 , n58202 , n58203 , n58204 , n58205 , n58206 , n58207 , n58208 , n58209 , n58210 , 
 n58211 , n58212 , n58213 , n58214 , n58215 , n58216 , n58217 , n58218 , n58219 , n58220 , 
 n58221 , n58222 , n58223 , n58224 , n58225 , n58226 , n58227 , n58228 , n58229 , n58230 , 
 n58231 , n58232 , n58233 , n58234 , n58235 , n58236 , n58237 , n58238 , n58239 , n58240 , 
 n58241 , n58242 , n58243 , n58244 , n58245 , n58246 , n58247 , n58248 , n58249 , n58250 , 
 n58251 , n58252 , n58253 , n58254 , n58255 , n58256 , n58257 , n58258 , n58259 , n58260 , 
 n58261 , n58262 , n58263 , n58264 , n58265 , n58266 , n58267 , n58268 , n58269 , n58270 , 
 n58271 , n58272 , n58273 , n58274 , n58275 , n58276 , n58277 , n58278 , n58279 , n58280 , 
 n58281 , n58282 , n58283 , n58284 , n58285 , n58286 , n58287 , n58288 , n58289 , n58290 , 
 n58291 , n58292 , n58293 , n58294 , n58295 , n58296 , n58297 , n58298 , n58299 , n58300 , 
 n58301 , n58302 , n58303 , n58304 , n58305 , n58306 , n58307 , n58308 , n58309 , n58310 , 
 n58311 , n58312 , n58313 , n58314 , n58315 , n58316 , n58317 , n58318 , n58319 , n58320 , 
 n58321 , n58322 , n58323 , n58324 , n58325 , n58326 , n58327 , n58328 , n58329 , n58330 , 
 n58331 , n58332 , n58333 , n58334 , n58335 , n58336 , n58337 , n58338 , n58339 , n58340 , 
 n58341 , n58342 , n58343 , n58344 , n58345 , n58346 , n58347 , n58348 , n58349 , n58350 , 
 n58351 , n58352 , n58353 , n58354 , n58355 , n58356 , n58357 , n58358 , n58359 , n58360 , 
 n58361 , n58362 , n58363 , n58364 , n58365 , n58366 , n58367 , n58368 , n58369 , n58370 , 
 n58371 , n58372 , n58373 , n58374 , n58375 , n58376 , n58377 , n58378 , n58379 , n58380 , 
 n58381 , n58382 , n58383 , n58384 , n58385 , n58386 , n58387 , n58388 , n58389 , n58390 , 
 n58391 , n58392 , n58393 , n58394 , n58395 , n58396 , n58397 , n58398 , n58399 , n58400 , 
 n58401 , n58402 , n58403 , n58404 , n58405 , n58406 , n58407 , n58408 , n58409 , n58410 , 
 n58411 , n58412 , n58413 , n58414 , n58415 , n58416 , n58417 , n58418 , n58419 , n58420 , 
 n58421 , n58422 , n58423 , n58424 , n58425 , n58426 , n58427 , n58428 , n58429 , n58430 , 
 n58431 , n58432 , n58433 , n58434 , n58435 , n58436 , n58437 , n58438 , n58439 , n58440 , 
 n58441 , n58442 , n58443 , n58444 , n58445 , n58446 , n58447 , n58448 , n58449 , n58450 , 
 n58451 , n58452 , n58453 , n58454 , n58455 , n58456 , n58457 , n58458 , n58459 , n58460 , 
 n58461 , n58462 , n58463 , n58464 , n58465 , n58466 , n58467 , n58468 , n58469 , n58470 , 
 n58471 , n58472 , n58473 , n58474 , n58475 , n58476 , n58477 , n58478 , n58479 , n58480 , 
 n58481 , n58482 , n58483 , n58484 , n58485 , n58486 , n58487 , n58488 , n58489 , n58490 , 
 n58491 , n58492 , n58493 , n58494 , n58495 , n58496 , n58497 , n58498 , n58499 , n58500 , 
 n58501 , n58502 , n58503 , n58504 , n58505 , n58506 , n58507 , n58508 , n58509 , n58510 , 
 n58511 , n58512 , n58513 , n58514 , n58515 , n58516 , n58517 , n58518 , n58519 , n58520 , 
 n58521 , n58522 , n58523 , n58524 , n58525 , n58526 , n58527 , n58528 , n58529 , n58530 , 
 n58531 , n58532 , n58533 , n58534 , n58535 , n58536 , n58537 , n58538 , n58539 , n58540 , 
 n58541 , n58542 , n58543 , n58544 , n58545 , n58546 , n58547 , n58548 , n58549 , n58550 , 
 n58551 , n58552 , n58553 , n58554 , n58555 , n58556 , n58557 , n58558 , n58559 , n58560 , 
 n58561 , n58562 , n58563 , n58564 , n58565 , n58566 , n58567 , n58568 , n58569 , n58570 , 
 n58571 , n58572 , n58573 , n58574 , n58575 , n58576 , n58577 , n58578 , n58579 , n58580 , 
 n58581 , n58582 , n58583 , n58584 , n58585 , n58586 , n58587 , n58588 , n58589 , n58590 , 
 n58591 , n58592 , n58593 , n58594 , n58595 , n58596 , n58597 , n58598 , n58599 , n58600 , 
 n58601 , n58602 , n58603 , n58604 , n58605 , n58606 , n58607 , n58608 , n58609 , n58610 , 
 n58611 , n58612 , n58613 , n58614 , n58615 , n58616 , n58617 , n58618 , n58619 , n58620 , 
 n58621 , n58622 , n58623 , n58624 , n58625 , n58626 , n58627 , n58628 , n58629 , n58630 , 
 n58631 , n58632 , n58633 , n58634 , n58635 , n58636 , n58637 , n58638 , n58639 , n58640 , 
 n58641 , n58642 , n58643 , n58644 , n58645 , n58646 , n58647 , n58648 , n58649 , n58650 , 
 n58651 , n58652 , n58653 , n58654 , n58655 , n58656 , n58657 , n58658 , n58659 , n58660 , 
 n58661 , n58662 , n58663 , n58664 , n58665 , n58666 , n58667 , n58668 , n58669 , n58670 , 
 n58671 , n58672 , n58673 , n58674 , n58675 , n58676 , n58677 , n58678 , n58679 , n58680 , 
 n58681 , n58682 , n58683 , n58684 , n58685 , n58686 , n58687 , n58688 , n58689 , n58690 , 
 n58691 , n58692 , n58693 , n58694 , n58695 , n58696 , n58697 , n58698 , n58699 , n58700 , 
 n58701 , n58702 , n58703 , n58704 , n58705 , n58706 , n58707 , n58708 , n58709 , n58710 , 
 n58711 , n58712 , n58713 , n58714 , n58715 , n58716 , n58717 , n58718 , n58719 , n58720 , 
 n58721 , n58722 , n58723 , n58724 , n58725 , n58726 , n58727 , n58728 , n58729 , n58730 , 
 n58731 , n58732 , n58733 , n58734 , n58735 , n58736 , n58737 , n58738 , n58739 , n58740 , 
 n58741 , n58742 , n58743 , n58744 , n58745 , n58746 , n58747 , n58748 , n58749 , n58750 , 
 n58751 , n58752 , n58753 , n58754 , n58755 , n58756 , n58757 , n58758 , n58759 , n58760 , 
 n58761 , n58762 , n58763 , n58764 , n58765 , n58766 , n58767 , n58768 , n58769 , n58770 , 
 n58771 , n58772 , n58773 , n58774 , n58775 , n58776 , n58777 , n58778 , n58779 , n58780 , 
 n58781 , n58782 , n58783 , n58784 , n58785 , n58786 , n58787 , n58788 , n58789 , n58790 , 
 n58791 , n58792 , n58793 , n58794 , n58795 , n58796 , n58797 , n58798 , n58799 , n58800 , 
 n58801 , n58802 , n58803 , n58804 , n58805 , n58806 , n58807 , n58808 , n58809 , n58810 , 
 n58811 , n58812 , n58813 , n58814 , n58815 , n58816 , n58817 , n58818 , n58819 , n58820 , 
 n58821 , n58822 , n58823 , n58824 , n58825 , n58826 , n58827 , n58828 , n58829 , n58830 , 
 n58831 , n58832 , n58833 , n58834 , n58835 , n58836 , n58837 , n58838 , n58839 , n58840 , 
 n58841 , n58842 , n58843 , n58844 , n58845 , n58846 , n58847 , n58848 , n58849 , n58850 , 
 n58851 , n58852 , n58853 , n58854 , n58855 , n58856 , n58857 , n58858 , n58859 , n58860 , 
 n58861 , n58862 , n58863 , n58864 , n58865 , n58866 , n58867 , n58868 , n58869 , n58870 , 
 n58871 , n58872 , n58873 , n58874 , n58875 , n58876 , n58877 , n58878 , n58879 , n58880 , 
 n58881 , n58882 , n58883 , n58884 , n58885 , n58886 , n58887 , n58888 , n58889 , n58890 , 
 n58891 , n58892 , n58893 , n58894 , n58895 , n58896 , n58897 , n58898 , n58899 , n58900 , 
 n58901 , n58902 , n58903 , n58904 , n58905 , n58906 , n58907 , n58908 , n58909 , n58910 , 
 n58911 , n58912 , n58913 , n58914 , n58915 , n58916 , n58917 , n58918 , n58919 , n58920 , 
 n58921 , n58922 , n58923 , n58924 , n58925 , n58926 , n58927 , n58928 , n58929 , n58930 , 
 n58931 , n58932 , n58933 , n58934 , n58935 , n58936 , n58937 , n58938 , n58939 , n58940 , 
 n58941 , n58942 , n58943 , n58944 , n58945 , n58946 , n58947 , n58948 , n58949 , n58950 , 
 n58951 , n58952 , n58953 , n58954 , n58955 , n58956 , n58957 , n58958 , n58959 , n58960 , 
 n58961 , n58962 , n58963 , n58964 , n58965 , n58966 , n58967 , n58968 , n58969 , n58970 , 
 n58971 , n58972 , n58973 , n58974 , n58975 , n58976 , n58977 , n58978 , n58979 , n58980 , 
 n58981 , n58982 , n58983 , n58984 , n58985 , n58986 , n58987 , n58988 , n58989 , n58990 , 
 n58991 , n58992 , n58993 , n58994 , n58995 , n58996 , n58997 , n58998 , n58999 , n59000 , 
 n59001 , n59002 , n59003 , n59004 , n59005 , n59006 , n59007 , n59008 , n59009 , n59010 , 
 n59011 , n59012 , n59013 , n59014 , n59015 , n59016 , n59017 , n59018 , n59019 , n59020 , 
 n59021 , n59022 , n59023 , n59024 , n59025 , n59026 , n59027 , n59028 , n59029 , n59030 , 
 n59031 , n59032 , n59033 , n59034 , n59035 , n59036 , n59037 , n59038 , n59039 , n59040 , 
 n59041 , n59042 , n59043 , n59044 , n59045 , n59046 , n59047 , n59048 , n59049 , n59050 , 
 n59051 , n59052 , n59053 , n59054 , n59055 , n59056 , n59057 , n59058 , n59059 , n59060 , 
 n59061 , n59062 , n59063 , n59064 , n59065 , n59066 , n59067 , n59068 , n59069 , n59070 , 
 n59071 , n59072 , n59073 , n59074 , n59075 , n59076 , n59077 , n59078 , n59079 , n59080 , 
 n59081 , n59082 , n59083 , n59084 , n59085 , n59086 , n59087 , n59088 , n59089 , n59090 , 
 n59091 , n59092 , n59093 , n59094 , n59095 , n59096 , n59097 , n59098 , n59099 , n59100 , 
 n59101 , n59102 , n59103 , n59104 , n59105 , n59106 , n59107 , n59108 , n59109 , n59110 , 
 n59111 , n59112 , n59113 , n59114 , n59115 , n59116 , n59117 , n59118 , n59119 , n59120 , 
 n59121 , n59122 , n59123 , n59124 , n59125 , n59126 , n59127 , n59128 , n59129 , n59130 , 
 n59131 , n59132 , n59133 , n59134 , n59135 , n59136 , n59137 , n59138 , n59139 , n59140 , 
 n59141 , n59142 , n59143 , n59144 , n59145 , n59146 , n59147 , n59148 , n59149 , n59150 , 
 n59151 , n59152 , n59153 , n59154 , n59155 , n59156 , n59157 , n59158 , n59159 , n59160 , 
 n59161 , n59162 , n59163 , n59164 , n59165 , n59166 , n59167 , n59168 , n59169 , n59170 , 
 n59171 , n59172 , n59173 , n59174 , n59175 , n59176 , n59177 , n59178 , n59179 , n59180 , 
 n59181 , n59182 , n59183 , n59184 , n59185 , n59186 , n59187 , n59188 , n59189 , n59190 , 
 n59191 , n59192 , n59193 , n59194 , n59195 , n59196 , n59197 , n59198 , n59199 , n59200 , 
 n59201 , n59202 , n59203 , n59204 , n59205 , n59206 , n59207 , n59208 , n59209 , n59210 , 
 n59211 , n59212 , n59213 , n59214 , n59215 , n59216 , n59217 , n59218 , n59219 , n59220 , 
 n59221 , n59222 , n59223 , n59224 , n59225 , n59226 , n59227 , n59228 , n59229 , n59230 , 
 n59231 , n59232 , n59233 , n59234 , n59235 , n59236 , n59237 , n59238 , n59239 , n59240 , 
 n59241 , n59242 , n59243 , n59244 , n59245 , n59246 , n59247 , n59248 , n59249 , n59250 , 
 n59251 , n59252 , n59253 , n59254 , n59255 , n59256 , n59257 , n59258 , n59259 , n59260 , 
 n59261 , n59262 , n59263 , n59264 , n59265 , n59266 , n59267 , n59268 , n59269 , n59270 , 
 n59271 , n59272 , n59273 , n59274 , n59275 , n59276 , n59277 , n59278 , n59279 , n59280 , 
 n59281 , n59282 , n59283 , n59284 , n59285 , n59286 , n59287 , n59288 , n59289 , n59290 , 
 n59291 , n59292 , n59293 , n59294 , n59295 , n59296 , n59297 , n59298 , n59299 , n59300 , 
 n59301 , n59302 , n59303 , n59304 , n59305 , n59306 , n59307 , n59308 , n59309 , n59310 , 
 n59311 , n59312 , n59313 , n59314 , n59315 , n59316 , n59317 , n59318 , n59319 , n59320 , 
 n59321 , n59322 , n59323 , n59324 , n59325 , n59326 , n59327 , n59328 , n59329 , n59330 , 
 n59331 , n59332 , n59333 , n59334 , n59335 , n59336 , n59337 , n59338 , n59339 , n59340 , 
 n59341 , n59342 , n59343 , n59344 , n59345 , n59346 , n59347 , n59348 , n59349 , n59350 , 
 n59351 , n59352 , n59353 , n59354 , n59355 , n59356 , n59357 , n59358 , n59359 , n59360 , 
 n59361 , n59362 , n59363 , n59364 , n59365 , n59366 , n59367 , n59368 , n59369 , n59370 , 
 n59371 , n59372 , n59373 , n59374 , n59375 , n59376 , n59377 , n59378 , n59379 , n59380 , 
 n59381 , n59382 , n59383 , n59384 , n59385 , n59386 , n59387 , n59388 , n59389 , n59390 , 
 n59391 , n59392 , n59393 , n59394 , n59395 , n59396 , n59397 , n59398 , n59399 , n59400 , 
 n59401 , n59402 , n59403 , n59404 , n59405 , n59406 , n59407 , n59408 , n59409 , n59410 , 
 n59411 , n59412 , n59413 , n59414 , n59415 , n59416 , n59417 , n59418 , n59419 , n59420 , 
 n59421 , n59422 , n59423 , n59424 , n59425 , n59426 , n59427 , n59428 , n59429 , n59430 , 
 n59431 , n59432 , n59433 , n59434 , n59435 , n59436 , n59437 , n59438 , n59439 , n59440 , 
 n59441 , n59442 , n59443 , n59444 , n59445 , n59446 , n59447 , n59448 , n59449 , n59450 , 
 n59451 , n59452 , n59453 , n59454 , n59455 , n59456 , n59457 , n59458 , n59459 , n59460 , 
 n59461 , n59462 , n59463 , n59464 , n59465 , n59466 , n59467 , n59468 , n59469 , n59470 , 
 n59471 , n59472 , n59473 , n59474 , n59475 , n59476 , n59477 , n59478 , n59479 , n59480 , 
 n59481 , n59482 , n59483 , n59484 , n59485 , n59486 , n59487 , n59488 , n59489 , n59490 , 
 n59491 , n59492 , n59493 , n59494 , n59495 , n59496 , n59497 , n59498 , n59499 , n59500 , 
 n59501 , n59502 , n59503 , n59504 , n59505 , n59506 , n59507 , n59508 , n59509 , n59510 , 
 n59511 , n59512 , n59513 , n59514 , n59515 , n59516 , n59517 , n59518 , n59519 , n59520 , 
 n59521 , n59522 , n59523 , n59524 , n59525 , n59526 , n59527 , n59528 , n59529 , n59530 , 
 n59531 , n59532 , n59533 , n59534 , n59535 , n59536 , n59537 , n59538 , n59539 , n59540 , 
 n59541 , n59542 , n59543 , n59544 , n59545 , n59546 , n59547 , n59548 , n59549 , n59550 , 
 n59551 , n59552 , n59553 , n59554 , n59555 , n59556 , n59557 , n59558 , n59559 , n59560 , 
 n59561 , n59562 , n59563 , n59564 , n59565 , n59566 , n59567 , n59568 , n59569 , n59570 , 
 n59571 , n59572 , n59573 , n59574 , n59575 , n59576 , n59577 , n59578 , n59579 , n59580 , 
 n59581 , n59582 , n59583 , n59584 , n59585 , n59586 , n59587 , n59588 , n59589 , n59590 , 
 n59591 , n59592 , n59593 , n59594 , n59595 , n59596 , n59597 , n59598 , n59599 , n59600 , 
 n59601 , n59602 , n59603 , n59604 , n59605 , n59606 , n59607 , n59608 , n59609 , n59610 , 
 n59611 , n59612 , n59613 , n59614 , n59615 , n59616 , n59617 , n59618 , n59619 , n59620 , 
 n59621 , n59622 , n59623 , n59624 , n59625 , n59626 , n59627 , n59628 , n59629 , n59630 , 
 n59631 , n59632 , n59633 , n59634 , n59635 , n59636 , n59637 , n59638 , n59639 , n59640 , 
 n59641 , n59642 , n59643 , n59644 , n59645 , n59646 , n59647 , n59648 , n59649 , n59650 , 
 n59651 , n59652 , n59653 , n59654 , n59655 , n59656 , n59657 , n59658 , n59659 , n59660 , 
 n59661 , n59662 , n59663 , n59664 , n59665 , n59666 , n59667 , n59668 , n59669 , n59670 , 
 n59671 , n59672 , n59673 , n59674 , n59675 , n59676 , n59677 , n59678 , n59679 , n59680 , 
 n59681 , n59682 , n59683 , n59684 , n59685 , n59686 , n59687 , n59688 , n59689 , n59690 , 
 n59691 , n59692 , n59693 , n59694 , n59695 , n59696 , n59697 , n59698 , n59699 , n59700 , 
 n59701 , n59702 , n59703 , n59704 , n59705 , n59706 , n59707 , n59708 , n59709 , n59710 , 
 n59711 , n59712 , n59713 , n59714 , n59715 , n59716 , n59717 , n59718 , n59719 , n59720 , 
 n59721 , n59722 , n59723 , n59724 , n59725 , n59726 , n59727 , n59728 , n59729 , n59730 , 
 n59731 , n59732 , n59733 , n59734 , n59735 , n59736 , n59737 , n59738 , n59739 , n59740 , 
 n59741 , n59742 , n59743 , n59744 , n59745 , n59746 , n59747 , n59748 , n59749 , n59750 , 
 n59751 , n59752 , n59753 , n59754 , n59755 , n59756 , n59757 , n59758 , n59759 , n59760 , 
 n59761 , n59762 , n59763 , n59764 , n59765 , n59766 , n59767 , n59768 , n59769 , n59770 , 
 n59771 , n59772 , n59773 , n59774 , n59775 , n59776 , n59777 , n59778 , n59779 , n59780 , 
 n59781 , n59782 , n59783 , n59784 , n59785 , n59786 , n59787 , n59788 , n59789 , n59790 , 
 n59791 , n59792 , n59793 , n59794 , n59795 , n59796 , n59797 , n59798 , n59799 , n59800 , 
 n59801 , n59802 , n59803 , n59804 , n59805 , n59806 , n59807 , n59808 , n59809 , n59810 , 
 n59811 , n59812 , n59813 , n59814 , n59815 , n59816 , n59817 , n59818 , n59819 , n59820 , 
 n59821 , n59822 , n59823 , n59824 , n59825 , n59826 , n59827 , n59828 , n59829 , n59830 , 
 n59831 , n59832 , n59833 , n59834 , n59835 , n59836 , n59837 , n59838 , n59839 , n59840 , 
 n59841 , n59842 , n59843 , n59844 , n59845 , n59846 , n59847 , n59848 , n59849 , n59850 , 
 n59851 , n59852 , n59853 , n59854 , n59855 , n59856 , n59857 , n59858 , n59859 , n59860 , 
 n59861 , n59862 , n59863 , n59864 , n59865 , n59866 , n59867 , n59868 , n59869 , n59870 , 
 n59871 , n59872 , n59873 , n59874 , n59875 , n59876 , n59877 , n59878 , n59879 , n59880 , 
 n59881 , n59882 , n59883 , n59884 , n59885 , n59886 , n59887 , n59888 , n59889 , n59890 , 
 n59891 , n59892 , n59893 , n59894 , n59895 , n59896 , n59897 , n59898 , n59899 , n59900 , 
 n59901 , n59902 , n59903 , n59904 , n59905 , n59906 , n59907 , n59908 , n59909 , n59910 , 
 n59911 , n59912 , n59913 , n59914 , n59915 , n59916 , n59917 , n59918 , n59919 , n59920 , 
 n59921 , n59922 , n59923 , n59924 , n59925 , n59926 , n59927 , n59928 , n59929 , n59930 , 
 n59931 , n59932 , n59933 , n59934 , n59935 , n59936 , n59937 , n59938 , n59939 , n59940 , 
 n59941 , n59942 , n59943 , n59944 , n59945 , n59946 , n59947 , n59948 , n59949 , n59950 , 
 n59951 , n59952 , n59953 , n59954 , n59955 , n59956 , n59957 , n59958 , n59959 , n59960 , 
 n59961 , n59962 , n59963 , n59964 , n59965 , n59966 , n59967 , n59968 , n59969 , n59970 , 
 n59971 , n59972 , n59973 , n59974 , n59975 , n59976 , n59977 , n59978 , n59979 , n59980 , 
 n59981 , n59982 , n59983 , n59984 , n59985 , n59986 , n59987 , n59988 , n59989 , n59990 , 
 n59991 , n59992 , n59993 , n59994 , n59995 , n59996 , n59997 , n59998 , n59999 , n60000 , 
 n60001 , n60002 , n60003 , n60004 , n60005 , n60006 , n60007 , n60008 , n60009 , n60010 , 
 n60011 , n60012 , n60013 , n60014 , n60015 , n60016 , n60017 , n60018 , n60019 , n60020 , 
 n60021 , n60022 , n60023 , n60024 , n60025 , n60026 , n60027 , n60028 , n60029 , n60030 , 
 n60031 , n60032 , n60033 , n60034 , n60035 , n60036 , n60037 , n60038 , n60039 , n60040 , 
 n60041 , n60042 , n60043 , n60044 , n60045 , n60046 , n60047 , n60048 , n60049 , n60050 , 
 n60051 , n60052 , n60053 , n60054 , n60055 , n60056 , n60057 , n60058 , n60059 , n60060 , 
 n60061 , n60062 , n60063 , n60064 , n60065 , n60066 , n60067 , n60068 , n60069 , n60070 , 
 n60071 , n60072 , n60073 , n60074 , n60075 , n60076 , n60077 , n60078 , n60079 , n60080 , 
 n60081 , n60082 , n60083 , n60084 , n60085 , n60086 , n60087 , n60088 , n60089 , n60090 , 
 n60091 , n60092 , n60093 , n60094 , n60095 , n60096 , n60097 , n60098 , n60099 , n60100 , 
 n60101 , n60102 , n60103 , n60104 , n60105 , n60106 , n60107 , n60108 , n60109 , n60110 , 
 n60111 , n60112 , n60113 , n60114 , n60115 , n60116 , n60117 , n60118 , n60119 , n60120 , 
 n60121 , n60122 , n60123 , n60124 , n60125 , n60126 , n60127 , n60128 , n60129 , n60130 , 
 n60131 , n60132 , n60133 , n60134 , n60135 , n60136 , n60137 , n60138 , n60139 , n60140 , 
 n60141 , n60142 , n60143 , n60144 , n60145 , n60146 , n60147 , n60148 , n60149 , n60150 , 
 n60151 , n60152 , n60153 , n60154 , n60155 , n60156 , n60157 , n60158 , n60159 , n60160 , 
 n60161 , n60162 , n60163 , n60164 , n60165 , n60166 , n60167 , n60168 , n60169 , n60170 , 
 n60171 , n60172 , n60173 , n60174 , n60175 , n60176 , n60177 , n60178 , n60179 , n60180 , 
 n60181 , n60182 , n60183 , n60184 , n60185 , n60186 , n60187 , n60188 , n60189 , n60190 , 
 n60191 , n60192 , n60193 , n60194 , n60195 , n60196 , n60197 , n60198 , n60199 , n60200 , 
 n60201 , n60202 , n60203 , n60204 , n60205 , n60206 , n60207 , n60208 , n60209 , n60210 , 
 n60211 , n60212 , n60213 , n60214 , n60215 , n60216 , n60217 , n60218 , n60219 , n60220 , 
 n60221 , n60222 , n60223 , n60224 , n60225 , n60226 , n60227 , n60228 , n60229 , n60230 , 
 n60231 , n60232 , n60233 , n60234 , n60235 , n60236 , n60237 , n60238 , n60239 , n60240 , 
 n60241 , n60242 , n60243 , n60244 , n60245 , n60246 , n60247 , n60248 , n60249 , n60250 , 
 n60251 , n60252 , n60253 , n60254 , n60255 , n60256 , n60257 , n60258 , n60259 , n60260 , 
 n60261 , n60262 , n60263 , n60264 , n60265 , n60266 , n60267 , n60268 , n60269 , n60270 , 
 n60271 , n60272 , n60273 , n60274 , n60275 , n60276 , n60277 , n60278 , n60279 , n60280 , 
 n60281 , n60282 , n60283 , n60284 , n60285 , n60286 , n60287 , n60288 , n60289 , n60290 , 
 n60291 , n60292 , n60293 , n60294 , n60295 , n60296 , n60297 , n60298 , n60299 , n60300 , 
 n60301 , n60302 , n60303 , n60304 , n60305 , n60306 , n60307 , n60308 , n60309 , n60310 , 
 n60311 , n60312 , n60313 , n60314 , n60315 , n60316 , n60317 , n60318 , n60319 , n60320 , 
 n60321 , n60322 , n60323 , n60324 , n60325 , n60326 , n60327 , n60328 , n60329 , n60330 , 
 n60331 , n60332 , n60333 , n60334 , n60335 , n60336 , n60337 , n60338 , n60339 , n60340 , 
 n60341 , n60342 , n60343 , n60344 , n60345 , n60346 , n60347 , n60348 , n60349 , n60350 , 
 n60351 , n60352 , n60353 , n60354 , n60355 , n60356 , n60357 , n60358 , n60359 , n60360 , 
 n60361 , n60362 , n60363 , n60364 , n60365 , n60366 , n60367 , n60368 , n60369 , n60370 , 
 n60371 , n60372 , n60373 , n60374 , n60375 , n60376 , n60377 , n60378 , n60379 , n60380 , 
 n60381 , n60382 , n60383 , n60384 , n60385 , n60386 , n60387 , n60388 , n60389 , n60390 , 
 n60391 , n60392 , n60393 , n60394 , n60395 , n60396 , n60397 , n60398 , n60399 , n60400 , 
 n60401 , n60402 , n60403 , n60404 , n60405 , n60406 , n60407 , n60408 , n60409 , n60410 , 
 n60411 , n60412 , n60413 , n60414 , n60415 , n60416 , n60417 , n60418 , n60419 , n60420 , 
 n60421 , n60422 , n60423 , n60424 , n60425 , n60426 , n60427 , n60428 , n60429 , n60430 , 
 n60431 , n60432 , n60433 , n60434 , n60435 , n60436 , n60437 , n60438 , n60439 , n60440 , 
 n60441 , n60442 , n60443 , n60444 , n60445 , n60446 , n60447 , n60448 , n60449 , n60450 , 
 n60451 , n60452 , n60453 , n60454 , n60455 , n60456 , n60457 , n60458 , n60459 , n60460 , 
 n60461 , n60462 , n60463 , n60464 , n60465 , n60466 , n60467 , n60468 , n60469 , n60470 , 
 n60471 , n60472 , n60473 , n60474 , n60475 , n60476 , n60477 , n60478 , n60479 , n60480 , 
 n60481 , n60482 , n60483 , n60484 , n60485 , n60486 , n60487 , n60488 , n60489 , n60490 , 
 n60491 , n60492 , n60493 , n60494 , n60495 , n60496 , n60497 , n60498 , n60499 , n60500 , 
 n60501 , n60502 , n60503 , n60504 , n60505 , n60506 , n60507 , n60508 , n60509 , n60510 , 
 n60511 , n60512 , n60513 , n60514 , n60515 , n60516 , n60517 , n60518 , n60519 , n60520 , 
 n60521 , n60522 , n60523 , n60524 , n60525 , n60526 , n60527 , n60528 , n60529 , n60530 , 
 n60531 , n60532 , n60533 , n60534 , n60535 , n60536 , n60537 , n60538 , n60539 , n60540 , 
 n60541 , n60542 , n60543 , n60544 , n60545 , n60546 , n60547 , n60548 , n60549 , n60550 , 
 n60551 , n60552 , n60553 , n60554 , n60555 , n60556 , n60557 , n60558 , n60559 , n60560 , 
 n60561 , n60562 , n60563 , n60564 , n60565 , n60566 , n60567 , n60568 , n60569 , n60570 , 
 n60571 , n60572 , n60573 , n60574 , n60575 , n60576 , n60577 , n60578 , n60579 , n60580 , 
 n60581 , n60582 , n60583 , n60584 , n60585 , n60586 , n60587 , n60588 , n60589 , n60590 , 
 n60591 , n60592 , n60593 , n60594 , n60595 , n60596 , n60597 , n60598 , n60599 , n60600 , 
 n60601 , n60602 , n60603 , n60604 , n60605 , n60606 , n60607 , n60608 , n60609 , n60610 , 
 n60611 , n60612 , n60613 , n60614 , n60615 , n60616 , n60617 , n60618 , n60619 , n60620 , 
 n60621 , n60622 , n60623 , n60624 , n60625 , n60626 , n60627 , n60628 , n60629 , n60630 , 
 n60631 , n60632 , n60633 , n60634 , n60635 , n60636 , n60637 , n60638 , n60639 , n60640 , 
 n60641 , n60642 , n60643 , n60644 , n60645 , n60646 , n60647 , n60648 , n60649 , n60650 , 
 n60651 , n60652 , n60653 , n60654 , n60655 , n60656 , n60657 , n60658 , n60659 , n60660 , 
 n60661 , n60662 , n60663 , n60664 , n60665 , n60666 , n60667 , n60668 , n60669 , n60670 , 
 n60671 , n60672 , n60673 , n60674 , n60675 , n60676 , n60677 , n60678 , n60679 , n60680 , 
 n60681 , n60682 , n60683 , n60684 , n60685 , n60686 , n60687 , n60688 , n60689 , n60690 , 
 n60691 , n60692 , n60693 , n60694 , n60695 , n60696 , n60697 , n60698 , n60699 , n60700 , 
 n60701 , n60702 , n60703 , n60704 , n60705 , n60706 , n60707 , n60708 , n60709 , n60710 , 
 n60711 , n60712 , n60713 , n60714 , n60715 , n60716 , n60717 , n60718 , n60719 , n60720 , 
 n60721 , n60722 , n60723 , n60724 , n60725 , n60726 , n60727 , n60728 , n60729 , n60730 , 
 n60731 , n60732 , n60733 , n60734 , n60735 , n60736 , n60737 , n60738 , n60739 , n60740 , 
 n60741 , n60742 , n60743 , n60744 , n60745 , n60746 , n60747 , n60748 , n60749 , n60750 , 
 n60751 , n60752 , n60753 , n60754 , n60755 , n60756 , n60757 , n60758 , n60759 , n60760 , 
 n60761 , n60762 , n60763 , n60764 , n60765 , n60766 , n60767 , n60768 , n60769 , n60770 , 
 n60771 , n60772 , n60773 , n60774 , n60775 , n60776 , n60777 , n60778 , n60779 , n60780 , 
 n60781 , n60782 , n60783 , n60784 , n60785 , n60786 , n60787 , n60788 , n60789 , n60790 , 
 n60791 , n60792 , n60793 , n60794 , n60795 , n60796 , n60797 , n60798 , n60799 , n60800 , 
 n60801 , n60802 , n60803 , n60804 , n60805 , n60806 , n60807 , n60808 , n60809 , n60810 , 
 n60811 , n60812 , n60813 , n60814 , n60815 , n60816 , n60817 , n60818 , n60819 , n60820 , 
 n60821 , n60822 , n60823 , n60824 , n60825 , n60826 , n60827 , n60828 , n60829 , n60830 , 
 n60831 , n60832 , n60833 , n60834 , n60835 , n60836 , n60837 , n60838 , n60839 , n60840 , 
 n60841 , n60842 , n60843 , n60844 , n60845 , n60846 , n60847 , n60848 , n60849 , n60850 , 
 n60851 , n60852 , n60853 , n60854 , n60855 , n60856 , n60857 , n60858 , n60859 , n60860 , 
 n60861 , n60862 , n60863 , n60864 , n60865 , n60866 , n60867 , n60868 , n60869 , n60870 , 
 n60871 , n60872 , n60873 , n60874 , n60875 , n60876 , n60877 , n60878 , n60879 , n60880 , 
 n60881 , n60882 , n60883 , n60884 , n60885 , n60886 , n60887 , n60888 , n60889 , n60890 , 
 n60891 , n60892 , n60893 , n60894 , n60895 , n60896 , n60897 , n60898 , n60899 , n60900 , 
 n60901 , n60902 , n60903 , n60904 , n60905 , n60906 , n60907 , n60908 , n60909 , n60910 , 
 n60911 , n60912 , n60913 , n60914 , n60915 , n60916 , n60917 , n60918 , n60919 , n60920 , 
 n60921 , n60922 , n60923 , n60924 , n60925 , n60926 , n60927 , n60928 , n60929 , n60930 , 
 n60931 , n60932 , n60933 , n60934 , n60935 , n60936 , n60937 , n60938 , n60939 , n60940 , 
 n60941 , n60942 , n60943 , n60944 , n60945 , n60946 , n60947 , n60948 , n60949 , n60950 , 
 n60951 , n60952 , n60953 , n60954 , n60955 , n60956 , n60957 , n60958 , n60959 , n60960 , 
 n60961 , n60962 , n60963 , n60964 , n60965 , n60966 , n60967 , n60968 , n60969 , n60970 , 
 n60971 , n60972 , n60973 , n60974 , n60975 , n60976 , n60977 , n60978 , n60979 , n60980 , 
 n60981 , n60982 , n60983 , n60984 , n60985 , n60986 , n60987 , n60988 , n60989 , n60990 , 
 n60991 , n60992 , n60993 , n60994 , n60995 , n60996 , n60997 , n60998 , n60999 , n61000 , 
 n61001 , n61002 , n61003 , n61004 , n61005 , n61006 , n61007 , n61008 , n61009 , n61010 , 
 n61011 , n61012 , n61013 , n61014 , n61015 , n61016 , n61017 , n61018 , n61019 , n61020 , 
 n61021 , n61022 , n61023 , n61024 , n61025 , n61026 , n61027 , n61028 , n61029 , n61030 , 
 n61031 , n61032 , n61033 , n61034 , n61035 , n61036 , n61037 , n61038 , n61039 , n61040 , 
 n61041 , n61042 , n61043 , n61044 , n61045 , n61046 , n61047 , n61048 , n61049 , n61050 , 
 n61051 , n61052 , n61053 , n61054 , n61055 , n61056 , n61057 , n61058 , n61059 , n61060 , 
 n61061 , n61062 , n61063 , n61064 , n61065 , n61066 , n61067 , n61068 , n61069 , n61070 , 
 n61071 , n61072 , n61073 , n61074 , n61075 , n61076 , n61077 , n61078 , n61079 , n61080 , 
 n61081 , n61082 , n61083 , n61084 , n61085 , n61086 , n61087 , n61088 , n61089 , n61090 , 
 n61091 , n61092 , n61093 , n61094 , n61095 , n61096 , n61097 , n61098 , n61099 , n61100 , 
 n61101 , n61102 , n61103 , n61104 , n61105 , n61106 , n61107 , n61108 , n61109 , n61110 , 
 n61111 , n61112 , n61113 , n61114 , n61115 , n61116 , n61117 , n61118 , n61119 , n61120 , 
 n61121 , n61122 , n61123 , n61124 , n61125 , n61126 , n61127 , n61128 , n61129 , n61130 , 
 n61131 , n61132 , n61133 , n61134 , n61135 , n61136 , n61137 , n61138 , n61139 , n61140 , 
 n61141 , n61142 , n61143 , n61144 , n61145 , n61146 , n61147 , n61148 , n61149 , n61150 , 
 n61151 , n61152 , n61153 , n61154 , n61155 , n61156 , n61157 , n61158 , n61159 , n61160 , 
 n61161 , n61162 , n61163 , n61164 , n61165 , n61166 , n61167 , n61168 , n61169 , n61170 , 
 n61171 , n61172 , n61173 , n61174 , n61175 , n61176 , n61177 , n61178 , n61179 , n61180 , 
 n61181 , n61182 , n61183 , n61184 , n61185 , n61186 , n61187 , n61188 , n61189 , n61190 , 
 n61191 , n61192 , n61193 , n61194 , n61195 , n61196 , n61197 , n61198 , n61199 , n61200 , 
 n61201 , n61202 , n61203 , n61204 , n61205 , n61206 , n61207 , n61208 , n61209 , n61210 , 
 n61211 , n61212 , n61213 , n61214 , n61215 , n61216 , n61217 , n61218 , n61219 , n61220 , 
 n61221 , n61222 , n61223 , n61224 , n61225 , n61226 , n61227 , n61228 , n61229 , n61230 , 
 n61231 , n61232 , n61233 , n61234 , n61235 , n61236 , n61237 , n61238 , n61239 , n61240 , 
 n61241 , n61242 , n61243 , n61244 , n61245 , n61246 , n61247 , n61248 , n61249 , n61250 , 
 n61251 , n61252 , n61253 , n61254 , n61255 , n61256 , n61257 , n61258 , n61259 , n61260 , 
 n61261 , n61262 , n61263 , n61264 , n61265 , n61266 , n61267 , n61268 , n61269 , n61270 , 
 n61271 , n61272 , n61273 , n61274 , n61275 , n61276 , n61277 , n61278 , n61279 , n61280 , 
 n61281 , n61282 , n61283 , n61284 , n61285 , n61286 , n61287 , n61288 , n61289 , n61290 , 
 n61291 , n61292 , n61293 , n61294 , n61295 , n61296 , n61297 , n61298 , n61299 , n61300 , 
 n61301 , n61302 , n61303 , n61304 , n61305 , n61306 , n61307 , n61308 , n61309 , n61310 , 
 n61311 , n61312 , n61313 , n61314 , n61315 , n61316 , n61317 , n61318 , n61319 , n61320 , 
 n61321 , n61322 , n61323 , n61324 , n61325 , n61326 , n61327 , n61328 , n61329 , n61330 , 
 n61331 , n61332 , n61333 , n61334 , n61335 , n61336 , n61337 , n61338 , n61339 , n61340 , 
 n61341 , n61342 , n61343 , n61344 , n61345 , n61346 , n61347 , n61348 , n61349 , n61350 , 
 n61351 , n61352 , n61353 , n61354 , n61355 , n61356 , n61357 , n61358 , n61359 , n61360 , 
 n61361 , n61362 , n61363 , n61364 , n61365 , n61366 , n61367 , n61368 , n61369 , n61370 , 
 n61371 , n61372 , n61373 , n61374 , n61375 , n61376 , n61377 , n61378 , n61379 , n61380 , 
 n61381 , n61382 , n61383 , n61384 , n61385 , n61386 , n61387 , n61388 , n61389 , n61390 , 
 n61391 , n61392 , n61393 , n61394 , n61395 , n61396 , n61397 , n61398 , n61399 , n61400 , 
 n61401 , n61402 , n61403 , n61404 , n61405 , n61406 , n61407 , n61408 , n61409 , n61410 , 
 n61411 , n61412 , n61413 , n61414 , n61415 , n61416 , n61417 , n61418 , n61419 , n61420 , 
 n61421 , n61422 , n61423 , n61424 , n61425 , n61426 , n61427 , n61428 , n61429 , n61430 , 
 n61431 , n61432 , n61433 , n61434 , n61435 , n61436 , n61437 , n61438 , n61439 , n61440 , 
 n61441 , n61442 , n61443 , n61444 , n61445 , n61446 , n61447 , n61448 , n61449 , n61450 , 
 n61451 , n61452 , n61453 , n61454 , n61455 , n61456 , n61457 , n61458 , n61459 , n61460 , 
 n61461 , n61462 , n61463 , n61464 , n61465 , n61466 , n61467 , n61468 , n61469 , n61470 , 
 n61471 , n61472 , n61473 , n61474 , n61475 , n61476 , n61477 , n61478 , n61479 , n61480 , 
 n61481 , n61482 , n61483 , n61484 , n61485 , n61486 , n61487 , n61488 , n61489 , n61490 , 
 n61491 , n61492 , n61493 , n61494 , n61495 , n61496 , n61497 , n61498 , n61499 , n61500 , 
 n61501 , n61502 , n61503 , n61504 , n61505 , n61506 , n61507 , n61508 , n61509 , n61510 , 
 n61511 , n61512 , n61513 , n61514 , n61515 , n61516 , n61517 , n61518 , n61519 , n61520 , 
 n61521 , n61522 , n61523 , n61524 , n61525 , n61526 , n61527 , n61528 , n61529 , n61530 , 
 n61531 , n61532 , n61533 , n61534 , n61535 , n61536 , n61537 , n61538 , n61539 , n61540 , 
 n61541 , n61542 , n61543 , n61544 , n61545 , n61546 , n61547 , n61548 , n61549 , n61550 , 
 n61551 , n61552 , n61553 , n61554 , n61555 , n61556 , n61557 , n61558 , n61559 , n61560 , 
 n61561 , n61562 , n61563 , n61564 , n61565 , n61566 , n61567 , n61568 , n61569 , n61570 , 
 n61571 , n61572 , n61573 , n61574 , n61575 , n61576 , n61577 , n61578 , n61579 , n61580 , 
 n61581 , n61582 , n61583 , n61584 , n61585 , n61586 , n61587 , n61588 , n61589 , n61590 , 
 n61591 , n61592 , n61593 , n61594 , n61595 , n61596 , n61597 , n61598 , n61599 , n61600 , 
 n61601 , n61602 , n61603 , n61604 , n61605 , n61606 , n61607 , n61608 , n61609 , n61610 , 
 n61611 , n61612 , n61613 , n61614 , n61615 , n61616 , n61617 , n61618 , n61619 , n61620 , 
 n61621 , n61622 , n61623 , n61624 , n61625 , n61626 , n61627 , n61628 , n61629 , n61630 , 
 n61631 , n61632 , n61633 , n61634 , n61635 , n61636 , n61637 , n61638 , n61639 , n61640 , 
 n61641 , n61642 , n61643 , n61644 , n61645 , n61646 , n61647 , n61648 , n61649 , n61650 , 
 n61651 , n61652 , n61653 , n61654 , n61655 , n61656 , n61657 , n61658 , n61659 , n61660 , 
 n61661 , n61662 , n61663 , n61664 , n61665 , n61666 , n61667 , n61668 , n61669 , n61670 , 
 n61671 , n61672 , n61673 , n61674 , n61675 , n61676 , n61677 , n61678 , n61679 , n61680 , 
 n61681 , n61682 , n61683 , n61684 , n61685 , n61686 , n61687 , n61688 , n61689 , n61690 , 
 n61691 , n61692 , n61693 , n61694 , n61695 , n61696 , n61697 , n61698 , n61699 , n61700 , 
 n61701 , n61702 , n61703 , n61704 , n61705 , n61706 , n61707 , n61708 , n61709 , n61710 , 
 n61711 , n61712 , n61713 , n61714 , n61715 , n61716 , n61717 , n61718 , n61719 , n61720 , 
 n61721 , n61722 , n61723 , n61724 , n61725 , n61726 , n61727 , n61728 , n61729 , n61730 , 
 n61731 , n61732 , n61733 , n61734 , n61735 , n61736 , n61737 , n61738 , n61739 , n61740 , 
 n61741 , n61742 , n61743 , n61744 , n61745 , n61746 , n61747 , n61748 , n61749 , n61750 , 
 n61751 , n61752 , n61753 , n61754 , n61755 , n61756 , n61757 , n61758 , n61759 , n61760 , 
 n61761 , n61762 , n61763 , n61764 , n61765 , n61766 , n61767 , n61768 , n61769 , n61770 , 
 n61771 , n61772 , n61773 , n61774 , n61775 , n61776 , n61777 , n61778 , n61779 , n61780 , 
 n61781 , n61782 , n61783 , n61784 , n61785 , n61786 , n61787 , n61788 , n61789 , n61790 , 
 n61791 , n61792 , n61793 , n61794 , n61795 , n61796 , n61797 , n61798 , n61799 , n61800 , 
 n61801 , n61802 , n61803 , n61804 , n61805 , n61806 , n61807 , n61808 , n61809 , n61810 , 
 n61811 , n61812 , n61813 , n61814 , n61815 , n61816 , n61817 , n61818 , n61819 , n61820 , 
 n61821 , n61822 , n61823 , n61824 , n61825 , n61826 , n61827 , n61828 , n61829 , n61830 , 
 n61831 , n61832 , n61833 , n61834 , n61835 , n61836 , n61837 , n61838 , n61839 , n61840 , 
 n61841 , n61842 , n61843 , n61844 , n61845 , n61846 , n61847 , n61848 , n61849 , n61850 , 
 n61851 , n61852 , n61853 , n61854 , n61855 , n61856 , n61857 , n61858 , n61859 , n61860 , 
 n61861 , n61862 , n61863 , n61864 , n61865 , n61866 , n61867 , n61868 , n61869 , n61870 , 
 n61871 , n61872 , n61873 , n61874 , n61875 , n61876 , n61877 , n61878 , n61879 , n61880 , 
 n61881 , n61882 , n61883 , n61884 , n61885 , n61886 , n61887 , n61888 , n61889 , n61890 , 
 n61891 , n61892 , n61893 , n61894 , n61895 , n61896 , n61897 , n61898 , n61899 , n61900 , 
 n61901 , n61902 , n61903 , n61904 , n61905 , n61906 , n61907 , n61908 , n61909 , n61910 , 
 n61911 , n61912 , n61913 , n61914 , n61915 , n61916 , n61917 , n61918 , n61919 , n61920 , 
 n61921 , n61922 , n61923 , n61924 , n61925 , n61926 , n61927 , n61928 , n61929 , n61930 , 
 n61931 , n61932 , n61933 , n61934 , n61935 , n61936 , n61937 , n61938 , n61939 , n61940 , 
 n61941 , n61942 , n61943 , n61944 , n61945 , n61946 , n61947 , n61948 , n61949 , n61950 , 
 n61951 , n61952 , n61953 , n61954 , n61955 , n61956 , n61957 , n61958 , n61959 , n61960 , 
 n61961 , n61962 , n61963 , n61964 , n61965 , n61966 , n61967 , n61968 , n61969 , n61970 , 
 n61971 , n61972 , n61973 , n61974 , n61975 , n61976 , n61977 , n61978 , n61979 , n61980 , 
 n61981 , n61982 , n61983 , n61984 , n61985 , n61986 , n61987 , n61988 , n61989 , n61990 , 
 n61991 , n61992 , n61993 , n61994 , n61995 , n61996 , n61997 , n61998 , n61999 , n62000 , 
 n62001 , n62002 , n62003 , n62004 , n62005 , n62006 , n62007 , n62008 , n62009 , n62010 , 
 n62011 , n62012 , n62013 , n62014 , n62015 , n62016 , n62017 , n62018 , n62019 , n62020 , 
 n62021 , n62022 , n62023 , n62024 , n62025 , n62026 , n62027 , n62028 , n62029 , n62030 , 
 n62031 , n62032 , n62033 , n62034 , n62035 , n62036 , n62037 , n62038 , n62039 , n62040 , 
 n62041 , n62042 , n62043 , n62044 , n62045 , n62046 , n62047 , n62048 , n62049 , n62050 , 
 n62051 , n62052 , n62053 , n62054 , n62055 , n62056 , n62057 , n62058 , n62059 , n62060 , 
 n62061 , n62062 , n62063 , n62064 , n62065 , n62066 , n62067 , n62068 , n62069 , n62070 , 
 n62071 , n62072 , n62073 , n62074 , n62075 , n62076 , n62077 , n62078 , n62079 , n62080 , 
 n62081 , n62082 , n62083 , n62084 , n62085 , n62086 , n62087 , n62088 , n62089 , n62090 , 
 n62091 , n62092 , n62093 , n62094 , n62095 , n62096 , n62097 , n62098 , n62099 , n62100 , 
 n62101 , n62102 , n62103 , n62104 , n62105 , n62106 , n62107 , n62108 , n62109 , n62110 , 
 n62111 , n62112 , n62113 , n62114 , n62115 , n62116 , n62117 , n62118 , n62119 , n62120 , 
 n62121 , n62122 , n62123 , n62124 , n62125 , n62126 , n62127 , n62128 , n62129 , n62130 , 
 n62131 , n62132 , n62133 , n62134 , n62135 , n62136 , n62137 , n62138 , n62139 , n62140 , 
 n62141 , n62142 , n62143 , n62144 , n62145 , n62146 , n62147 , n62148 , n62149 , n62150 , 
 n62151 , n62152 , n62153 , n62154 , n62155 , n62156 , n62157 , n62158 , n62159 , n62160 , 
 n62161 , n62162 , n62163 , n62164 , n62165 , n62166 , n62167 , n62168 , n62169 , n62170 , 
 n62171 , n62172 , n62173 , n62174 , n62175 , n62176 , n62177 , n62178 , n62179 , n62180 , 
 n62181 , n62182 , n62183 , n62184 , n62185 , n62186 , n62187 , n62188 , n62189 , n62190 , 
 n62191 , n62192 , n62193 , n62194 , n62195 , n62196 , n62197 , n62198 , n62199 , n62200 , 
 n62201 , n62202 , n62203 , n62204 , n62205 , n62206 , n62207 , n62208 , n62209 , n62210 , 
 n62211 , n62212 , n62213 , n62214 , n62215 , n62216 , n62217 , n62218 , n62219 , n62220 , 
 n62221 , n62222 , n62223 , n62224 , n62225 , n62226 , n62227 , n62228 , n62229 , n62230 , 
 n62231 , n62232 , n62233 , n62234 , n62235 , n62236 , n62237 , n62238 , n62239 , n62240 , 
 n62241 , n62242 , n62243 , n62244 , n62245 , n62246 , n62247 , n62248 , n62249 , n62250 , 
 n62251 , n62252 , n62253 , n62254 , n62255 , n62256 , n62257 , n62258 , n62259 , n62260 , 
 n62261 , n62262 , n62263 , n62264 , n62265 , n62266 , n62267 , n62268 , n62269 , n62270 , 
 n62271 , n62272 , n62273 , n62274 , n62275 , n62276 , n62277 , n62278 , n62279 , n62280 , 
 n62281 , n62282 , n62283 , n62284 , n62285 , n62286 , n62287 , n62288 , n62289 , n62290 , 
 n62291 , n62292 , n62293 , n62294 , n62295 , n62296 , n62297 , n62298 , n62299 , n62300 , 
 n62301 , n62302 , n62303 , n62304 , n62305 , n62306 , n62307 , n62308 , n62309 , n62310 , 
 n62311 , n62312 , n62313 , n62314 , n62315 , n62316 , n62317 , n62318 , n62319 , n62320 , 
 n62321 , n62322 , n62323 , n62324 , n62325 , n62326 , n62327 , n62328 , n62329 , n62330 , 
 n62331 , n62332 , n62333 , n62334 , n62335 , n62336 , n62337 , n62338 , n62339 , n62340 , 
 n62341 , n62342 , n62343 , n62344 , n62345 , n62346 , n62347 , n62348 , n62349 , n62350 , 
 n62351 , n62352 , n62353 , n62354 , n62355 , n62356 , n62357 , n62358 , n62359 , n62360 , 
 n62361 , n62362 , n62363 , n62364 , n62365 , n62366 , n62367 , n62368 , n62369 , n62370 , 
 n62371 , n62372 , n62373 , n62374 , n62375 , n62376 , n62377 , n62378 , n62379 , n62380 , 
 n62381 , n62382 , n62383 , n62384 , n62385 , n62386 , n62387 , n62388 , n62389 , n62390 , 
 n62391 , n62392 , n62393 , n62394 , n62395 , n62396 , n62397 , n62398 , n62399 , n62400 , 
 n62401 , n62402 , n62403 , n62404 , n62405 , n62406 , n62407 , n62408 , n62409 , n62410 , 
 n62411 , n62412 , n62413 , n62414 , n62415 , n62416 , n62417 , n62418 , n62419 , n62420 , 
 n62421 , n62422 , n62423 , n62424 , n62425 , n62426 , n62427 , n62428 , n62429 , n62430 , 
 n62431 , n62432 , n62433 , n62434 , n62435 , n62436 , n62437 , n62438 , n62439 , n62440 , 
 n62441 , n62442 , n62443 , n62444 , n62445 , n62446 , n62447 , n62448 , n62449 , n62450 , 
 n62451 , n62452 , n62453 , n62454 , n62455 , n62456 , n62457 , n62458 , n62459 , n62460 , 
 n62461 , n62462 , n62463 , n62464 , n62465 , n62466 , n62467 , n62468 , n62469 , n62470 , 
 n62471 , n62472 , n62473 , n62474 , n62475 , n62476 , n62477 , n62478 , n62479 , n62480 , 
 n62481 , n62482 , n62483 , n62484 , n62485 , n62486 , n62487 , n62488 , n62489 , n62490 , 
 n62491 , n62492 , n62493 , n62494 , n62495 , n62496 , n62497 , n62498 , n62499 , n62500 , 
 n62501 , n62502 , n62503 , n62504 , n62505 , n62506 , n62507 , n62508 , n62509 , n62510 , 
 n62511 , n62512 , n62513 , n62514 , n62515 , n62516 , n62517 , n62518 , n62519 , n62520 , 
 n62521 , n62522 , n62523 , n62524 , n62525 , n62526 , n62527 , n62528 , n62529 , n62530 , 
 n62531 , n62532 , n62533 , n62534 , n62535 , n62536 , n62537 , n62538 , n62539 , n62540 , 
 n62541 , n62542 , n62543 , n62544 , n62545 , n62546 , n62547 , n62548 , n62549 , n62550 , 
 n62551 , n62552 , n62553 , n62554 , n62555 , n62556 , n62557 , n62558 , n62559 , n62560 , 
 n62561 , n62562 , n62563 , n62564 , n62565 , n62566 , n62567 , n62568 , n62569 , n62570 , 
 n62571 , n62572 , n62573 , n62574 , n62575 , n62576 , n62577 , n62578 , n62579 , n62580 , 
 n62581 , n62582 , n62583 , n62584 , n62585 , n62586 , n62587 , n62588 , n62589 , n62590 , 
 n62591 , n62592 , n62593 , n62594 , n62595 , n62596 , n62597 , n62598 , n62599 , n62600 , 
 n62601 , n62602 , n62603 , n62604 , n62605 , n62606 , n62607 , n62608 , n62609 , n62610 , 
 n62611 , n62612 , n62613 , n62614 , n62615 , n62616 , n62617 , n62618 , n62619 , n62620 , 
 n62621 , n62622 , n62623 , n62624 , n62625 , n62626 , n62627 , n62628 , n62629 , n62630 , 
 n62631 , n62632 , n62633 , n62634 , n62635 , n62636 , n62637 , n62638 , n62639 , n62640 , 
 n62641 , n62642 , n62643 , n62644 , n62645 , n62646 , n62647 , n62648 , n62649 , n62650 , 
 n62651 , n62652 , n62653 , n62654 , n62655 , n62656 , n62657 , n62658 , n62659 , n62660 , 
 n62661 , n62662 , n62663 , n62664 , n62665 , n62666 , n62667 , n62668 , n62669 , n62670 , 
 n62671 , n62672 , n62673 , n62674 , n62675 , n62676 , n62677 , n62678 , n62679 , n62680 , 
 n62681 , n62682 , n62683 , n62684 , n62685 , n62686 , n62687 , n62688 , n62689 , n62690 , 
 n62691 , n62692 , n62693 , n62694 , n62695 , n62696 , n62697 , n62698 , n62699 , n62700 , 
 n62701 , n62702 , n62703 , n62704 , n62705 , n62706 , n62707 , n62708 , n62709 , n62710 , 
 n62711 , n62712 , n62713 , n62714 , n62715 , n62716 , n62717 , n62718 , n62719 , n62720 , 
 n62721 , n62722 , n62723 , n62724 , n62725 , n62726 , n62727 , n62728 , n62729 , n62730 , 
 n62731 , n62732 , n62733 , n62734 , n62735 , n62736 , n62737 , n62738 , n62739 , n62740 , 
 n62741 , n62742 , n62743 , n62744 , n62745 , n62746 , n62747 , n62748 , n62749 , n62750 , 
 n62751 , n62752 , n62753 , n62754 , n62755 , n62756 , n62757 , n62758 , n62759 , n62760 , 
 n62761 , n62762 , n62763 , n62764 , n62765 , n62766 , n62767 , n62768 , n62769 , n62770 , 
 n62771 , n62772 , n62773 , n62774 , n62775 , n62776 , n62777 , n62778 , n62779 , n62780 , 
 n62781 , n62782 , n62783 , n62784 , n62785 , n62786 , n62787 , n62788 , n62789 , n62790 , 
 n62791 , n62792 , n62793 , n62794 , n62795 , n62796 , n62797 , n62798 , n62799 , n62800 , 
 n62801 , n62802 , n62803 , n62804 , n62805 , n62806 , n62807 , n62808 , n62809 , n62810 , 
 n62811 , n62812 , n62813 , n62814 , n62815 , n62816 , n62817 , n62818 , n62819 , n62820 , 
 n62821 , n62822 , n62823 , n62824 , n62825 , n62826 , n62827 , n62828 , n62829 , n62830 , 
 n62831 , n62832 , n62833 , n62834 , n62835 , n62836 , n62837 , n62838 , n62839 , n62840 , 
 n62841 , n62842 , n62843 , n62844 , n62845 , n62846 , n62847 , n62848 , n62849 , n62850 , 
 n62851 , n62852 , n62853 , n62854 , n62855 , n62856 , n62857 , n62858 , n62859 , n62860 , 
 n62861 , n62862 , n62863 , n62864 , n62865 , n62866 , n62867 , n62868 , n62869 , n62870 , 
 n62871 , n62872 , n62873 , n62874 , n62875 , n62876 , n62877 , n62878 , n62879 , n62880 , 
 n62881 , n62882 , n62883 , n62884 , n62885 , n62886 , n62887 , n62888 , n62889 , n62890 , 
 n62891 , n62892 , n62893 , n62894 , n62895 , n62896 , n62897 , n62898 , n62899 , n62900 , 
 n62901 , n62902 , n62903 , n62904 , n62905 , n62906 , n62907 , n62908 , n62909 , n62910 , 
 n62911 , n62912 , n62913 , n62914 , n62915 , n62916 , n62917 , n62918 , n62919 , n62920 , 
 n62921 , n62922 , n62923 , n62924 , n62925 , n62926 , n62927 , n62928 , n62929 , n62930 , 
 n62931 , n62932 , n62933 , n62934 , n62935 , n62936 , n62937 , n62938 , n62939 , n62940 , 
 n62941 , n62942 , n62943 , n62944 , n62945 , n62946 , n62947 , n62948 , n62949 , n62950 , 
 n62951 , n62952 , n62953 , n62954 , n62955 , n62956 , n62957 , n62958 , n62959 , n62960 , 
 n62961 , n62962 , n62963 , n62964 , n62965 , n62966 , n62967 , n62968 , n62969 , n62970 , 
 n62971 , n62972 , n62973 , n62974 , n62975 , n62976 , n62977 , n62978 , n62979 , n62980 , 
 n62981 , n62982 , n62983 , n62984 , n62985 , n62986 , n62987 , n62988 , n62989 , n62990 , 
 n62991 , n62992 , n62993 , n62994 , n62995 , n62996 , n62997 , n62998 , n62999 , n63000 , 
 n63001 , n63002 , n63003 , n63004 , n63005 , n63006 , n63007 , n63008 , n63009 , n63010 , 
 n63011 , n63012 , n63013 , n63014 , n63015 , n63016 , n63017 , n63018 , n63019 , n63020 , 
 n63021 , n63022 , n63023 , n63024 , n63025 , n63026 , n63027 , n63028 , n63029 , n63030 , 
 n63031 , n63032 , n63033 , n63034 , n63035 , n63036 , n63037 , n63038 , n63039 , n63040 , 
 n63041 , n63042 , n63043 , n63044 , n63045 , n63046 , n63047 , n63048 , n63049 , n63050 , 
 n63051 , n63052 , n63053 , n63054 , n63055 , n63056 , n63057 , n63058 , n63059 , n63060 , 
 n63061 , n63062 , n63063 , n63064 , n63065 , n63066 , n63067 , n63068 , n63069 , n63070 , 
 n63071 , n63072 , n63073 , n63074 , n63075 , n63076 , n63077 , n63078 , n63079 , n63080 , 
 n63081 , n63082 , n63083 , n63084 , n63085 , n63086 , n63087 , n63088 , n63089 , n63090 , 
 n63091 , n63092 , n63093 , n63094 , n63095 , n63096 , n63097 , n63098 , n63099 , n63100 , 
 n63101 , n63102 , n63103 , n63104 , n63105 , n63106 , n63107 , n63108 , n63109 , n63110 , 
 n63111 , n63112 , n63113 , n63114 , n63115 , n63116 , n63117 , n63118 , n63119 , n63120 , 
 n63121 , n63122 , n63123 , n63124 , n63125 , n63126 , n63127 , n63128 , n63129 , n63130 , 
 n63131 , n63132 , n63133 , n63134 , n63135 , n63136 , n63137 , n63138 , n63139 , n63140 , 
 n63141 , n63142 , n63143 , n63144 , n63145 , n63146 , n63147 , n63148 , n63149 , n63150 , 
 n63151 , n63152 , n63153 , n63154 , n63155 , n63156 , n63157 , n63158 , n63159 , n63160 , 
 n63161 , n63162 , n63163 , n63164 , n63165 , n63166 , n63167 , n63168 , n63169 , n63170 , 
 n63171 , n63172 , n63173 , n63174 , n63175 , n63176 , n63177 , n63178 , n63179 , n63180 , 
 n63181 , n63182 , n63183 , n63184 , n63185 , n63186 , n63187 , n63188 , n63189 , n63190 , 
 n63191 , n63192 , n63193 , n63194 , n63195 , n63196 , n63197 , n63198 , n63199 , n63200 , 
 n63201 , n63202 , n63203 , n63204 , n63205 , n63206 , n63207 , n63208 , n63209 , n63210 , 
 n63211 , n63212 , n63213 , n63214 , n63215 , n63216 , n63217 , n63218 , n63219 , n63220 , 
 n63221 , n63222 , n63223 , n63224 , n63225 , n63226 , n63227 , n63228 , n63229 , n63230 , 
 n63231 , n63232 , n63233 , n63234 , n63235 , n63236 , n63237 , n63238 , n63239 , n63240 , 
 n63241 , n63242 , n63243 , n63244 , n63245 , n63246 , n63247 , n63248 , n63249 , n63250 , 
 n63251 , n63252 , n63253 , n63254 , n63255 , n63256 , n63257 , n63258 , n63259 , n63260 , 
 n63261 , n63262 , n63263 , n63264 , n63265 , n63266 , n63267 , n63268 , n63269 , n63270 , 
 n63271 , n63272 , n63273 , n63274 , n63275 , n63276 , n63277 , n63278 , n63279 , n63280 , 
 n63281 , n63282 , n63283 , n63284 , n63285 , n63286 , n63287 , n63288 , n63289 , n63290 , 
 n63291 , n63292 , n63293 , n63294 , n63295 , n63296 , n63297 , n63298 , n63299 , n63300 , 
 n63301 , n63302 , n63303 , n63304 , n63305 , n63306 , n63307 , n63308 , n63309 , n63310 , 
 n63311 , n63312 , n63313 , n63314 , n63315 , n63316 , n63317 , n63318 , n63319 , n63320 , 
 n63321 , n63322 , n63323 , n63324 , n63325 , n63326 , n63327 , n63328 , n63329 , n63330 , 
 n63331 , n63332 , n63333 , n63334 , n63335 , n63336 , n63337 , n63338 , n63339 , n63340 , 
 n63341 , n63342 , n63343 , n63344 , n63345 , n63346 , n63347 , n63348 , n63349 , n63350 , 
 n63351 , n63352 , n63353 , n63354 , n63355 , n63356 , n63357 , n63358 , n63359 , n63360 , 
 n63361 , n63362 , n63363 , n63364 , n63365 , n63366 , n63367 , n63368 , n63369 , n63370 , 
 n63371 , n63372 , n63373 , n63374 , n63375 , n63376 , n63377 , n63378 , n63379 , n63380 , 
 n63381 , n63382 , n63383 , n63384 , n63385 , n63386 , n63387 , n63388 , n63389 , n63390 , 
 n63391 , n63392 , n63393 , n63394 , n63395 , n63396 , n63397 , n63398 , n63399 , n63400 , 
 n63401 , n63402 , n63403 , n63404 , n63405 , n63406 , n63407 , n63408 , n63409 , n63410 , 
 n63411 , n63412 , n63413 , n63414 , n63415 , n63416 , n63417 , n63418 , n63419 , n63420 , 
 n63421 , n63422 , n63423 , n63424 , n63425 , n63426 , n63427 , n63428 , n63429 , n63430 , 
 n63431 , n63432 , n63433 , n63434 , n63435 , n63436 , n63437 , n63438 , n63439 , n63440 , 
 n63441 , n63442 , n63443 , n63444 , n63445 , n63446 , n63447 , n63448 , n63449 , n63450 , 
 n63451 , n63452 , n63453 , n63454 , n63455 , n63456 , n63457 , n63458 , n63459 , n63460 , 
 n63461 , n63462 , n63463 , n63464 , n63465 , n63466 , n63467 , n63468 , n63469 , n63470 , 
 n63471 , n63472 , n63473 , n63474 , n63475 , n63476 , n63477 , n63478 , n63479 , n63480 , 
 n63481 , n63482 , n63483 , n63484 , n63485 , n63486 , n63487 , n63488 , n63489 , n63490 , 
 n63491 , n63492 , n63493 , n63494 , n63495 , n63496 , n63497 , n63498 , n63499 , n63500 , 
 n63501 , n63502 , n63503 , n63504 , n63505 , n63506 , n63507 , n63508 , n63509 , n63510 , 
 n63511 , n63512 , n63513 , n63514 , n63515 , n63516 , n63517 , n63518 , n63519 , n63520 , 
 n63521 , n63522 , n63523 , n63524 , n63525 , n63526 , n63527 , n63528 , n63529 , n63530 , 
 n63531 , n63532 , n63533 , n63534 , n63535 , n63536 , n63537 , n63538 , n63539 , n63540 , 
 n63541 , n63542 , n63543 , n63544 , n63545 , n63546 , n63547 , n63548 , n63549 , n63550 , 
 n63551 , n63552 , n63553 , n63554 , n63555 , n63556 , n63557 , n63558 , n63559 , n63560 , 
 n63561 , n63562 , n63563 , n63564 , n63565 , n63566 , n63567 , n63568 , n63569 , n63570 , 
 n63571 , n63572 , n63573 , n63574 , n63575 , n63576 , n63577 , n63578 , n63579 , n63580 , 
 n63581 , n63582 , n63583 , n63584 , n63585 , n63586 , n63587 , n63588 , n63589 , n63590 , 
 n63591 , n63592 , n63593 , n63594 , n63595 , n63596 , n63597 , n63598 , n63599 , n63600 , 
 n63601 , n63602 , n63603 , n63604 , n63605 , n63606 , n63607 , n63608 , n63609 , n63610 , 
 n63611 , n63612 , n63613 , n63614 , n63615 , n63616 , n63617 , n63618 , n63619 , n63620 , 
 n63621 , n63622 , n63623 , n63624 , n63625 , n63626 , n63627 , n63628 , n63629 , n63630 , 
 n63631 , n63632 , n63633 , n63634 , n63635 , n63636 , n63637 , n63638 , n63639 , n63640 , 
 n63641 , n63642 , n63643 , n63644 , n63645 , n63646 , n63647 , n63648 , n63649 , n63650 , 
 n63651 , n63652 , n63653 , n63654 , n63655 , n63656 , n63657 , n63658 , n63659 , n63660 , 
 n63661 , n63662 , n63663 , n63664 , n63665 , n63666 , n63667 , n63668 , n63669 , n63670 , 
 n63671 , n63672 , n63673 , n63674 , n63675 , n63676 , n63677 , n63678 , n63679 , n63680 , 
 n63681 , n63682 , n63683 , n63684 , n63685 , n63686 , n63687 , n63688 , n63689 , n63690 , 
 n63691 , n63692 , n63693 , n63694 , n63695 , n63696 , n63697 , n63698 , n63699 , n63700 , 
 n63701 , n63702 , n63703 , n63704 , n63705 , n63706 , n63707 , n63708 , n63709 , n63710 , 
 n63711 , n63712 , n63713 , n63714 , n63715 , n63716 , n63717 , n63718 , n63719 , n63720 , 
 n63721 , n63722 , n63723 , n63724 , n63725 , n63726 , n63727 , n63728 , n63729 , n63730 , 
 n63731 , n63732 , n63733 , n63734 , n63735 , n63736 , n63737 , n63738 , n63739 , n63740 , 
 n63741 , n63742 , n63743 , n63744 , n63745 , n63746 , n63747 , n63748 , n63749 , n63750 , 
 n63751 , n63752 , n63753 , n63754 , n63755 , n63756 , n63757 , n63758 , n63759 , n63760 , 
 n63761 , n63762 , n63763 , n63764 , n63765 , n63766 , n63767 , n63768 , n63769 , n63770 , 
 n63771 , n63772 , n63773 , n63774 , n63775 , n63776 , n63777 , n63778 , n63779 , n63780 , 
 n63781 , n63782 , n63783 , n63784 , n63785 , n63786 , n63787 , n63788 , n63789 , n63790 , 
 n63791 , n63792 , n63793 , n63794 , n63795 , n63796 , n63797 , n63798 , n63799 , n63800 , 
 n63801 , n63802 , n63803 , n63804 , n63805 , n63806 , n63807 , n63808 , n63809 , n63810 , 
 n63811 , n63812 , n63813 , n63814 , n63815 , n63816 , n63817 , n63818 , n63819 , n63820 , 
 n63821 , n63822 , n63823 , n63824 , n63825 , n63826 , n63827 , n63828 , n63829 , n63830 , 
 n63831 , n63832 , n63833 , n63834 , n63835 , n63836 , n63837 , n63838 , n63839 , n63840 , 
 n63841 , n63842 , n63843 , n63844 , n63845 , n63846 , n63847 , n63848 , n63849 , n63850 , 
 n63851 , n63852 , n63853 , n63854 , n63855 , n63856 , n63857 , n63858 , n63859 , n63860 , 
 n63861 , n63862 , n63863 , n63864 , n63865 , n63866 , n63867 , n63868 , n63869 , n63870 , 
 n63871 , n63872 , n63873 , n63874 , n63875 , n63876 , n63877 , n63878 , n63879 , n63880 , 
 n63881 , n63882 , n63883 , n63884 , n63885 , n63886 , n63887 , n63888 , n63889 , n63890 , 
 n63891 , n63892 , n63893 , n63894 , n63895 , n63896 , n63897 , n63898 , n63899 , n63900 , 
 n63901 , n63902 , n63903 , n63904 , n63905 , n63906 , n63907 , n63908 , n63909 , n63910 , 
 n63911 , n63912 , n63913 , n63914 , n63915 , n63916 , n63917 , n63918 , n63919 , n63920 , 
 n63921 , n63922 , n63923 , n63924 , n63925 , n63926 , n63927 , n63928 , n63929 , n63930 , 
 n63931 , n63932 , n63933 , n63934 , n63935 , n63936 , n63937 , n63938 , n63939 , n63940 , 
 n63941 , n63942 , n63943 , n63944 , n63945 , n63946 , n63947 , n63948 , n63949 , n63950 , 
 n63951 , n63952 , n63953 , n63954 , n63955 , n63956 , n63957 , n63958 , n63959 , n63960 , 
 n63961 , n63962 , n63963 , n63964 , n63965 , n63966 , n63967 , n63968 , n63969 , n63970 , 
 n63971 , n63972 , n63973 , n63974 , n63975 , n63976 , n63977 , n63978 , n63979 , n63980 , 
 n63981 , n63982 , n63983 , n63984 , n63985 , n63986 , n63987 , n63988 , n63989 , n63990 , 
 n63991 , n63992 , n63993 , n63994 , n63995 , n63996 , n63997 , n63998 , n63999 , n64000 , 
 n64001 , n64002 , n64003 , n64004 , n64005 , n64006 , n64007 , n64008 , n64009 , n64010 , 
 n64011 , n64012 , n64013 , n64014 , n64015 , n64016 , n64017 , n64018 , n64019 , n64020 , 
 n64021 , n64022 , n64023 , n64024 , n64025 , n64026 , n64027 , n64028 , n64029 , n64030 , 
 n64031 , n64032 , n64033 , n64034 , n64035 , n64036 , n64037 , n64038 , n64039 , n64040 , 
 n64041 , n64042 , n64043 , n64044 , n64045 , n64046 , n64047 , n64048 , n64049 , n64050 , 
 n64051 , n64052 , n64053 , n64054 , n64055 , n64056 , n64057 , n64058 , n64059 , n64060 , 
 n64061 , n64062 , n64063 , n64064 , n64065 , n64066 , n64067 , n64068 , n64069 , n64070 , 
 n64071 , n64072 , n64073 , n64074 , n64075 , n64076 , n64077 , n64078 , n64079 , n64080 , 
 n64081 , n64082 , n64083 , n64084 , n64085 , n64086 , n64087 , n64088 , n64089 , n64090 , 
 n64091 , n64092 , n64093 , n64094 , n64095 , n64096 , n64097 , n64098 , n64099 , n64100 , 
 n64101 , n64102 , n64103 , n64104 , n64105 , n64106 , n64107 , n64108 , n64109 , n64110 , 
 n64111 , n64112 , n64113 , n64114 , n64115 , n64116 , n64117 , n64118 , n64119 , n64120 , 
 n64121 , n64122 , n64123 , n64124 , n64125 , n64126 , n64127 , n64128 , n64129 , n64130 , 
 n64131 , n64132 , n64133 , n64134 , n64135 , n64136 , n64137 , n64138 , n64139 , n64140 , 
 n64141 , n64142 , n64143 , n64144 , n64145 , n64146 , n64147 , n64148 , n64149 , n64150 , 
 n64151 , n64152 , n64153 , n64154 , n64155 , n64156 , n64157 , n64158 , n64159 , n64160 , 
 n64161 , n64162 , n64163 , n64164 , n64165 , n64166 , n64167 , n64168 , n64169 , n64170 , 
 n64171 , n64172 , n64173 , n64174 , n64175 , n64176 , n64177 , n64178 , n64179 , n64180 , 
 n64181 , n64182 , n64183 , n64184 , n64185 , n64186 , n64187 , n64188 , n64189 , n64190 , 
 n64191 , n64192 , n64193 , n64194 , n64195 , n64196 , n64197 , n64198 , n64199 , n64200 , 
 n64201 , n64202 , n64203 , n64204 , n64205 , n64206 , n64207 , n64208 , n64209 , n64210 , 
 n64211 , n64212 , n64213 , n64214 , n64215 , n64216 , n64217 , n64218 , n64219 , n64220 , 
 n64221 , n64222 , n64223 , n64224 , n64225 , n64226 , n64227 , n64228 , n64229 , n64230 , 
 n64231 , n64232 , n64233 , n64234 , n64235 , n64236 , n64237 , n64238 , n64239 , n64240 , 
 n64241 , n64242 , n64243 , n64244 , n64245 , n64246 , n64247 , n64248 , n64249 , n64250 , 
 n64251 , n64252 , n64253 , n64254 , n64255 , n64256 , n64257 , n64258 , n64259 , n64260 , 
 n64261 , n64262 , n64263 , n64264 , n64265 , n64266 , n64267 , n64268 , n64269 , n64270 , 
 n64271 , n64272 , n64273 , n64274 , n64275 , n64276 , n64277 , n64278 , n64279 , n64280 , 
 n64281 , n64282 , n64283 , n64284 , n64285 , n64286 , n64287 , n64288 , n64289 , n64290 , 
 n64291 , n64292 , n64293 , n64294 , n64295 , n64296 , n64297 , n64298 , n64299 , n64300 , 
 n64301 , n64302 , n64303 , n64304 , n64305 , n64306 , n64307 , n64308 , n64309 , n64310 , 
 n64311 , n64312 , n64313 , n64314 , n64315 , n64316 , n64317 , n64318 , n64319 , n64320 , 
 n64321 , n64322 , n64323 , n64324 , n64325 , n64326 , n64327 , n64328 , n64329 , n64330 , 
 n64331 , n64332 , n64333 , n64334 , n64335 , n64336 , n64337 , n64338 , n64339 , n64340 , 
 n64341 , n64342 , n64343 , n64344 , n64345 , n64346 , n64347 , n64348 , n64349 , n64350 , 
 n64351 , n64352 , n64353 , n64354 , n64355 , n64356 , n64357 , n64358 , n64359 , n64360 , 
 n64361 , n64362 , n64363 , n64364 , n64365 , n64366 , n64367 , n64368 , n64369 , n64370 , 
 n64371 , n64372 , n64373 , n64374 , n64375 , n64376 , n64377 , n64378 , n64379 , n64380 , 
 n64381 , n64382 , n64383 , n64384 , n64385 , n64386 , n64387 , n64388 , n64389 , n64390 , 
 n64391 , n64392 , n64393 , n64394 , n64395 , n64396 , n64397 , n64398 , n64399 , n64400 , 
 n64401 , n64402 , n64403 , n64404 , n64405 , n64406 , n64407 , n64408 , n64409 , n64410 , 
 n64411 , n64412 , n64413 , n64414 , n64415 , n64416 , n64417 , n64418 , n64419 , n64420 , 
 n64421 , n64422 , n64423 , n64424 , n64425 , n64426 , n64427 , n64428 , n64429 , n64430 , 
 n64431 , n64432 , n64433 , n64434 , n64435 , n64436 , n64437 , n64438 , n64439 , n64440 , 
 n64441 , n64442 , n64443 , n64444 , n64445 , n64446 , n64447 , n64448 , n64449 , n64450 , 
 n64451 , n64452 , n64453 , n64454 , n64455 , n64456 , n64457 , n64458 , n64459 , n64460 , 
 n64461 , n64462 , n64463 , n64464 , n64465 , n64466 , n64467 , n64468 , n64469 , n64470 , 
 n64471 , n64472 , n64473 , n64474 , n64475 , n64476 , n64477 , n64478 , n64479 , n64480 , 
 n64481 , n64482 , n64483 , n64484 , n64485 , n64486 , n64487 , n64488 , n64489 , n64490 , 
 n64491 , n64492 , n64493 , n64494 , n64495 , n64496 , n64497 , n64498 , n64499 , n64500 , 
 n64501 , n64502 , n64503 , n64504 , n64505 , n64506 , n64507 , n64508 , n64509 , n64510 , 
 n64511 , n64512 , n64513 , n64514 , n64515 , n64516 , n64517 , n64518 , n64519 , n64520 , 
 n64521 , n64522 , n64523 , n64524 , n64525 , n64526 , n64527 , n64528 , n64529 , n64530 , 
 n64531 , n64532 , n64533 , n64534 , n64535 , n64536 , n64537 , n64538 , n64539 , n64540 , 
 n64541 , n64542 , n64543 , n64544 , n64545 , n64546 , n64547 , n64548 , n64549 , n64550 , 
 n64551 , n64552 , n64553 , n64554 , n64555 , n64556 , n64557 , n64558 , n64559 , n64560 , 
 n64561 , n64562 , n64563 , n64564 , n64565 , n64566 , n64567 , n64568 , n64569 , n64570 , 
 n64571 , n64572 , n64573 , n64574 , n64575 , n64576 , n64577 , n64578 , n64579 , n64580 , 
 n64581 , n64582 , n64583 , n64584 , n64585 , n64586 , n64587 , n64588 , n64589 , n64590 , 
 n64591 , n64592 , n64593 , n64594 , n64595 , n64596 , n64597 , n64598 , n64599 , n64600 , 
 n64601 , n64602 , n64603 , n64604 , n64605 , n64606 , n64607 , n64608 , n64609 , n64610 , 
 n64611 , n64612 , n64613 , n64614 , n64615 , n64616 , n64617 , n64618 , n64619 , n64620 , 
 n64621 , n64622 , n64623 , n64624 , n64625 , n64626 , n64627 , n64628 , n64629 , n64630 , 
 n64631 , n64632 , n64633 , n64634 , n64635 , n64636 , n64637 , n64638 , n64639 , n64640 , 
 n64641 , n64642 , n64643 , n64644 , n64645 , n64646 , n64647 , n64648 , n64649 , n64650 , 
 n64651 , n64652 , n64653 , n64654 , n64655 , n64656 , n64657 , n64658 , n64659 , n64660 , 
 n64661 , n64662 , n64663 , n64664 , n64665 , n64666 , n64667 , n64668 , n64669 , n64670 , 
 n64671 , n64672 , n64673 , n64674 , n64675 , n64676 , n64677 , n64678 , n64679 , n64680 , 
 n64681 , n64682 , n64683 , n64684 , n64685 , n64686 , n64687 , n64688 , n64689 , n64690 , 
 n64691 , n64692 , n64693 , n64694 , n64695 , n64696 , n64697 , n64698 , n64699 , n64700 , 
 n64701 , n64702 , n64703 , n64704 , n64705 , n64706 , n64707 , n64708 , n64709 , n64710 , 
 n64711 , n64712 , n64713 , n64714 , n64715 , n64716 , n64717 , n64718 , n64719 , n64720 , 
 n64721 , n64722 , n64723 , n64724 , n64725 , n64726 , n64727 , n64728 , n64729 , n64730 , 
 n64731 , n64732 , n64733 , n64734 , n64735 , n64736 , n64737 , n64738 , n64739 , n64740 , 
 n64741 , n64742 , n64743 , n64744 , n64745 , n64746 , n64747 , n64748 , n64749 , n64750 , 
 n64751 , n64752 , n64753 , n64754 , n64755 , n64756 , n64757 , n64758 , n64759 , n64760 , 
 n64761 , n64762 , n64763 , n64764 , n64765 , n64766 , n64767 , n64768 , n64769 , n64770 , 
 n64771 , n64772 , n64773 , n64774 , n64775 , n64776 , n64777 , n64778 , n64779 , n64780 , 
 n64781 , n64782 , n64783 , n64784 , n64785 , n64786 , n64787 , n64788 , n64789 , n64790 , 
 n64791 , n64792 , n64793 , n64794 , n64795 , n64796 , n64797 , n64798 , n64799 , n64800 , 
 n64801 , n64802 , n64803 , n64804 , n64805 , n64806 , n64807 , n64808 , n64809 , n64810 , 
 n64811 , n64812 , n64813 , n64814 , n64815 , n64816 , n64817 , n64818 , n64819 , n64820 , 
 n64821 , n64822 , n64823 , n64824 , n64825 , n64826 , n64827 , n64828 , n64829 , n64830 , 
 n64831 , n64832 , n64833 , n64834 , n64835 , n64836 , n64837 , n64838 , n64839 , n64840 , 
 n64841 , n64842 , n64843 , n64844 , n64845 , n64846 , n64847 , n64848 , n64849 , n64850 , 
 n64851 , n64852 , n64853 , n64854 , n64855 , n64856 , n64857 , n64858 , n64859 , n64860 , 
 n64861 , n64862 , n64863 , n64864 , n64865 , n64866 , n64867 , n64868 , n64869 , n64870 , 
 n64871 , n64872 , n64873 , n64874 , n64875 , n64876 , n64877 , n64878 , n64879 , n64880 , 
 n64881 , n64882 , n64883 , n64884 , n64885 , n64886 , n64887 , n64888 , n64889 , n64890 , 
 n64891 , n64892 , n64893 , n64894 , n64895 , n64896 , n64897 , n64898 , n64899 , n64900 , 
 n64901 , n64902 , n64903 , n64904 , n64905 , n64906 , n64907 , n64908 , n64909 , n64910 , 
 n64911 , n64912 , n64913 , n64914 , n64915 , n64916 , n64917 , n64918 , n64919 , n64920 , 
 n64921 , n64922 , n64923 , n64924 , n64925 , n64926 , n64927 , n64928 , n64929 , n64930 , 
 n64931 , n64932 , n64933 , n64934 , n64935 , n64936 , n64937 , n64938 , n64939 , n64940 , 
 n64941 , n64942 , n64943 , n64944 , n64945 , n64946 , n64947 , n64948 , n64949 , n64950 , 
 n64951 , n64952 , n64953 , n64954 , n64955 , n64956 , n64957 , n64958 , n64959 , n64960 , 
 n64961 , n64962 , n64963 , n64964 , n64965 , n64966 , n64967 , n64968 , n64969 , n64970 , 
 n64971 , n64972 , n64973 , n64974 , n64975 , n64976 , n64977 , n64978 , n64979 , n64980 , 
 n64981 , n64982 , n64983 , n64984 , n64985 , n64986 , n64987 , n64988 , n64989 , n64990 , 
 n64991 , n64992 , n64993 , n64994 , n64995 , n64996 , n64997 , n64998 , n64999 , n65000 , 
 n65001 , n65002 , n65003 , n65004 , n65005 , n65006 , n65007 , n65008 , n65009 , n65010 , 
 n65011 , n65012 , n65013 , n65014 , n65015 , n65016 , n65017 , n65018 , n65019 , n65020 , 
 n65021 , n65022 , n65023 , n65024 , n65025 , n65026 , n65027 , n65028 , n65029 , n65030 , 
 n65031 , n65032 , n65033 , n65034 , n65035 , n65036 , n65037 , n65038 , n65039 , n65040 , 
 n65041 , n65042 , n65043 , n65044 , n65045 , n65046 , n65047 , n65048 , n65049 , n65050 , 
 n65051 , n65052 , n65053 , n65054 , n65055 , n65056 , n65057 , n65058 , n65059 , n65060 , 
 n65061 , n65062 , n65063 , n65064 , n65065 , n65066 , n65067 , n65068 , n65069 , n65070 , 
 n65071 , n65072 , n65073 , n65074 , n65075 , n65076 , n65077 , n65078 , n65079 , n65080 , 
 n65081 , n65082 , n65083 , n65084 , n65085 , n65086 , n65087 , n65088 , n65089 , n65090 , 
 n65091 , n65092 , n65093 , n65094 , n65095 , n65096 , n65097 , n65098 , n65099 , n65100 , 
 n65101 , n65102 , n65103 , n65104 , n65105 , n65106 , n65107 , n65108 , n65109 , n65110 , 
 n65111 , n65112 , n65113 , n65114 , n65115 , n65116 , n65117 , n65118 , n65119 , n65120 , 
 n65121 , n65122 , n65123 , n65124 , n65125 , n65126 , n65127 , n65128 , n65129 , n65130 , 
 n65131 , n65132 , n65133 , n65134 , n65135 , n65136 , n65137 , n65138 , n65139 , n65140 , 
 n65141 , n65142 , n65143 , n65144 , n65145 , n65146 , n65147 , n65148 , n65149 , n65150 , 
 n65151 , n65152 , n65153 , n65154 , n65155 , n65156 , n65157 , n65158 , n65159 , n65160 , 
 n65161 , n65162 , n65163 , n65164 , n65165 , n65166 , n65167 , n65168 , n65169 , n65170 , 
 n65171 , n65172 , n65173 , n65174 , n65175 , n65176 , n65177 , n65178 , n65179 , n65180 , 
 n65181 , n65182 , n65183 , n65184 , n65185 , n65186 , n65187 , n65188 , n65189 , n65190 , 
 n65191 , n65192 , n65193 , n65194 , n65195 , n65196 , n65197 , n65198 , n65199 , n65200 , 
 n65201 , n65202 , n65203 , n65204 , n65205 , n65206 , n65207 , n65208 , n65209 , n65210 , 
 n65211 , n65212 , n65213 , n65214 , n65215 , n65216 , n65217 , n65218 , n65219 , n65220 , 
 n65221 , n65222 , n65223 , n65224 , n65225 , n65226 , n65227 , n65228 , n65229 , n65230 , 
 n65231 , n65232 , n65233 , n65234 , n65235 , n65236 , n65237 , n65238 , n65239 , n65240 , 
 n65241 , n65242 , n65243 , n65244 , n65245 , n65246 , n65247 , n65248 , n65249 , n65250 , 
 n65251 , n65252 , n65253 , n65254 , n65255 , n65256 , n65257 , n65258 , n65259 , n65260 , 
 n65261 , n65262 , n65263 , n65264 , n65265 , n65266 , n65267 , n65268 , n65269 , n65270 , 
 n65271 , n65272 , n65273 , n65274 , n65275 , n65276 , n65277 , n65278 , n65279 , n65280 , 
 n65281 , n65282 , n65283 , n65284 , n65285 , n65286 , n65287 , n65288 , n65289 , n65290 , 
 n65291 , n65292 , n65293 , n65294 , n65295 , n65296 , n65297 , n65298 , n65299 , n65300 , 
 n65301 , n65302 , n65303 , n65304 , n65305 , n65306 , n65307 , n65308 , n65309 , n65310 , 
 n65311 , n65312 , n65313 , n65314 , n65315 , n65316 , n65317 , n65318 , n65319 , n65320 , 
 n65321 , n65322 , n65323 , n65324 , n65325 , n65326 , n65327 , n65328 , n65329 , n65330 , 
 n65331 , n65332 , n65333 , n65334 , n65335 , n65336 , n65337 , n65338 , n65339 , n65340 , 
 n65341 , n65342 , n65343 , n65344 , n65345 , n65346 , n65347 , n65348 , n65349 , n65350 , 
 n65351 , n65352 , n65353 , n65354 , n65355 , n65356 , n65357 , n65358 , n65359 , n65360 , 
 n65361 , n65362 , n65363 , n65364 , n65365 , n65366 , n65367 , n65368 , n65369 , n65370 , 
 n65371 , n65372 , n65373 , n65374 , n65375 , n65376 , n65377 , n65378 , n65379 , n65380 , 
 n65381 , n65382 , n65383 , n65384 , n65385 , n65386 , n65387 , n65388 , n65389 , n65390 , 
 n65391 , n65392 , n65393 , n65394 , n65395 , n65396 , n65397 , n65398 , n65399 , n65400 , 
 n65401 , n65402 , n65403 , n65404 , n65405 , n65406 , n65407 , n65408 , n65409 , n65410 , 
 n65411 , n65412 , n65413 , n65414 , n65415 , n65416 , n65417 , n65418 , n65419 , n65420 , 
 n65421 , n65422 , n65423 , n65424 , n65425 , n65426 , n65427 , n65428 , n65429 , n65430 , 
 n65431 , n65432 , n65433 , n65434 , n65435 , n65436 , n65437 , n65438 , n65439 , n65440 , 
 n65441 , n65442 , n65443 , n65444 , n65445 , n65446 , n65447 , n65448 , n65449 , n65450 , 
 n65451 , n65452 , n65453 , n65454 , n65455 , n65456 , n65457 , n65458 , n65459 , n65460 , 
 n65461 , n65462 , n65463 , n65464 , n65465 , n65466 , n65467 , n65468 , n65469 , n65470 , 
 n65471 , n65472 , n65473 , n65474 , n65475 , n65476 , n65477 , n65478 , n65479 , n65480 , 
 n65481 , n65482 , n65483 , n65484 , n65485 , n65486 , n65487 , n65488 , n65489 , n65490 , 
 n65491 , n65492 , n65493 , n65494 , n65495 , n65496 , n65497 , n65498 , n65499 , n65500 , 
 n65501 , n65502 , n65503 , n65504 , n65505 , n65506 , n65507 , n65508 , n65509 , n65510 , 
 n65511 , n65512 , n65513 , n65514 , n65515 , n65516 , n65517 , n65518 , n65519 , n65520 , 
 n65521 , n65522 , n65523 , n65524 , n65525 , n65526 , n65527 , n65528 , n65529 , n65530 , 
 n65531 , n65532 , n65533 , n65534 , n65535 , n65536 , n65537 , n65538 , n65539 , n65540 , 
 n65541 , n65542 , n65543 , n65544 , n65545 , n65546 , n65547 , n65548 , n65549 , n65550 , 
 n65551 , n65552 , n65553 , n65554 , n65555 , n65556 , n65557 , n65558 , n65559 , n65560 , 
 n65561 , n65562 , n65563 , n65564 , n65565 , n65566 , n65567 , n65568 , n65569 , n65570 , 
 n65571 , n65572 , n65573 , n65574 , n65575 , n65576 , n65577 , n65578 , n65579 , n65580 , 
 n65581 , n65582 , n65583 , n65584 , n65585 , n65586 , n65587 , n65588 , n65589 , n65590 , 
 n65591 , n65592 , n65593 , n65594 , n65595 , n65596 , n65597 , n65598 , n65599 , n65600 , 
 n65601 , n65602 , n65603 , n65604 , n65605 , n65606 , n65607 , n65608 , n65609 , n65610 , 
 n65611 , n65612 , n65613 , n65614 , n65615 , n65616 , n65617 , n65618 , n65619 , n65620 , 
 n65621 , n65622 , n65623 , n65624 , n65625 , n65626 , n65627 , n65628 , n65629 , n65630 , 
 n65631 , n65632 , n65633 , n65634 , n65635 , n65636 , n65637 , n65638 , n65639 , n65640 , 
 n65641 , n65642 , n65643 , n65644 , n65645 , n65646 , n65647 , n65648 , n65649 , n65650 , 
 n65651 , n65652 , n65653 , n65654 , n65655 , n65656 , n65657 , n65658 , n65659 , n65660 , 
 n65661 , n65662 , n65663 , n65664 , n65665 , n65666 , n65667 , n65668 , n65669 , n65670 , 
 n65671 , n65672 , n65673 , n65674 , n65675 , n65676 , n65677 , n65678 , n65679 , n65680 , 
 n65681 , n65682 , n65683 , n65684 , n65685 , n65686 , n65687 , n65688 , n65689 , n65690 , 
 n65691 , n65692 , n65693 , n65694 , n65695 , n65696 , n65697 , n65698 , n65699 , n65700 , 
 n65701 , n65702 , n65703 , n65704 , n65705 , n65706 , n65707 , n65708 , n65709 , n65710 , 
 n65711 , n65712 , n65713 , n65714 , n65715 , n65716 , n65717 , n65718 , n65719 , n65720 , 
 n65721 , n65722 , n65723 , n65724 , n65725 , n65726 , n65727 , n65728 , n65729 , n65730 , 
 n65731 , n65732 , n65733 , n65734 , n65735 , n65736 , n65737 , n65738 , n65739 , n65740 , 
 n65741 , n65742 , n65743 , n65744 , n65745 , n65746 , n65747 , n65748 , n65749 , n65750 , 
 n65751 , n65752 , n65753 , n65754 , n65755 , n65756 , n65757 , n65758 , n65759 , n65760 , 
 n65761 , n65762 , n65763 , n65764 , n65765 , n65766 , n65767 , n65768 , n65769 , n65770 , 
 n65771 , n65772 , n65773 , n65774 , n65775 , n65776 , n65777 , n65778 , n65779 , n65780 , 
 n65781 , n65782 , n65783 , n65784 , n65785 , n65786 , n65787 , n65788 , n65789 , n65790 , 
 n65791 , n65792 , n65793 , n65794 , n65795 , n65796 , n65797 , n65798 , n65799 , n65800 , 
 n65801 , n65802 , n65803 , n65804 , n65805 , n65806 , n65807 , n65808 , n65809 , n65810 , 
 n65811 , n65812 , n65813 , n65814 , n65815 , n65816 , n65817 , n65818 , n65819 , n65820 , 
 n65821 , n65822 , n65823 , n65824 , n65825 , n65826 , n65827 , n65828 , n65829 , n65830 , 
 n65831 , n65832 , n65833 , n65834 , n65835 , n65836 , n65837 , n65838 , n65839 , n65840 , 
 n65841 , n65842 , n65843 , n65844 , n65845 , n65846 , n65847 , n65848 , n65849 , n65850 , 
 n65851 , n65852 , n65853 , n65854 , n65855 , n65856 , n65857 , n65858 , n65859 , n65860 , 
 n65861 , n65862 , n65863 , n65864 , n65865 , n65866 , n65867 , n65868 , n65869 , n65870 , 
 n65871 , n65872 , n65873 , n65874 , n65875 , n65876 , n65877 , n65878 , n65879 , n65880 , 
 n65881 , n65882 , n65883 , n65884 , n65885 , n65886 , n65887 , n65888 , n65889 , n65890 , 
 n65891 , n65892 , n65893 , n65894 , n65895 , n65896 , n65897 , n65898 , n65899 , n65900 , 
 n65901 , n65902 , n65903 , n65904 , n65905 , n65906 , n65907 , n65908 , n65909 , n65910 , 
 n65911 , n65912 , n65913 , n65914 , n65915 , n65916 , n65917 , n65918 , n65919 , n65920 , 
 n65921 , n65922 , n65923 , n65924 , n65925 , n65926 , n65927 , n65928 , n65929 , n65930 , 
 n65931 , n65932 , n65933 , n65934 , n65935 , n65936 , n65937 , n65938 , n65939 , n65940 , 
 n65941 , n65942 , n65943 , n65944 , n65945 , n65946 , n65947 , n65948 , n65949 , n65950 , 
 n65951 , n65952 , n65953 , n65954 , n65955 , n65956 , n65957 , n65958 , n65959 , n65960 , 
 n65961 , n65962 , n65963 , n65964 , n65965 , n65966 , n65967 , n65968 , n65969 , n65970 , 
 n65971 , n65972 , n65973 , n65974 , n65975 , n65976 , n65977 , n65978 , n65979 , n65980 , 
 n65981 , n65982 , n65983 , n65984 , n65985 , n65986 , n65987 , n65988 , n65989 , n65990 , 
 n65991 , n65992 , n65993 , n65994 , n65995 , n65996 , n65997 , n65998 , n65999 , n66000 , 
 n66001 , n66002 , n66003 , n66004 , n66005 , n66006 , n66007 , n66008 , n66009 , n66010 , 
 n66011 , n66012 , n66013 , n66014 , n66015 , n66016 , n66017 , n66018 , n66019 , n66020 , 
 n66021 , n66022 , n66023 , n66024 , n66025 , n66026 , n66027 , n66028 , n66029 , n66030 , 
 n66031 , n66032 , n66033 , n66034 , n66035 , n66036 , n66037 , n66038 , n66039 , n66040 , 
 n66041 , n66042 , n66043 , n66044 , n66045 , n66046 , n66047 , n66048 , n66049 , n66050 , 
 n66051 , n66052 , n66053 , n66054 , n66055 , n66056 , n66057 , n66058 , n66059 , n66060 , 
 n66061 , n66062 , n66063 , n66064 , n66065 , n66066 , n66067 , n66068 , n66069 , n66070 , 
 n66071 , n66072 , n66073 , n66074 , n66075 , n66076 , n66077 , n66078 , n66079 , n66080 , 
 n66081 , n66082 , n66083 , n66084 , n66085 , n66086 , n66087 , n66088 , n66089 , n66090 , 
 n66091 , n66092 , n66093 , n66094 , n66095 , n66096 , n66097 , n66098 , n66099 , n66100 , 
 n66101 , n66102 , n66103 , n66104 , n66105 , n66106 , n66107 , n66108 , n66109 , n66110 , 
 n66111 , n66112 , n66113 , n66114 , n66115 , n66116 , n66117 , n66118 , n66119 , n66120 , 
 n66121 , n66122 , n66123 , n66124 , n66125 , n66126 , n66127 , n66128 , n66129 , n66130 , 
 n66131 , n66132 , n66133 , n66134 , n66135 , n66136 , n66137 , n66138 , n66139 , n66140 , 
 n66141 , n66142 , n66143 , n66144 , n66145 , n66146 , n66147 , n66148 , n66149 , n66150 , 
 n66151 , n66152 , n66153 , n66154 , n66155 , n66156 , n66157 , n66158 , n66159 , n66160 , 
 n66161 , n66162 , n66163 , n66164 , n66165 , n66166 , n66167 , n66168 , n66169 , n66170 , 
 n66171 , n66172 , n66173 , n66174 , n66175 , n66176 , n66177 , n66178 , n66179 , n66180 , 
 n66181 , n66182 , n66183 , n66184 , n66185 , n66186 , n66187 , n66188 , n66189 , n66190 , 
 n66191 , n66192 , n66193 , n66194 , n66195 , n66196 , n66197 , n66198 , n66199 , n66200 , 
 n66201 , n66202 , n66203 , n66204 , n66205 , n66206 , n66207 , n66208 , n66209 , n66210 , 
 n66211 , n66212 , n66213 , n66214 , n66215 , n66216 , n66217 , n66218 , n66219 , n66220 , 
 n66221 , n66222 , n66223 , n66224 , n66225 , n66226 , n66227 , n66228 , n66229 , n66230 , 
 n66231 , n66232 , n66233 , n66234 , n66235 , n66236 , n66237 , n66238 , n66239 , n66240 , 
 n66241 , n66242 , n66243 , n66244 , n66245 , n66246 , n66247 , n66248 , n66249 , n66250 , 
 n66251 , n66252 , n66253 , n66254 , n66255 , n66256 , n66257 , n66258 , n66259 , n66260 , 
 n66261 , n66262 , n66263 , n66264 , n66265 , n66266 , n66267 , n66268 , n66269 , n66270 , 
 n66271 , n66272 , n66273 , n66274 , n66275 , n66276 , n66277 , n66278 , n66279 , n66280 , 
 n66281 , n66282 , n66283 , n66284 , n66285 , n66286 , n66287 , n66288 , n66289 , n66290 , 
 n66291 , n66292 , n66293 , n66294 , n66295 , n66296 , n66297 , n66298 , n66299 , n66300 , 
 n66301 , n66302 , n66303 , n66304 , n66305 , n66306 , n66307 , n66308 , n66309 , n66310 , 
 n66311 , n66312 , n66313 , n66314 , n66315 , n66316 , n66317 , n66318 , n66319 , n66320 , 
 n66321 , n66322 , n66323 , n66324 , n66325 , n66326 , n66327 , n66328 , n66329 , n66330 , 
 n66331 , n66332 , n66333 , n66334 , n66335 , n66336 , n66337 , n66338 , n66339 , n66340 , 
 n66341 , n66342 , n66343 , n66344 , n66345 , n66346 , n66347 , n66348 , n66349 , n66350 , 
 n66351 , n66352 , n66353 , n66354 , n66355 , n66356 , n66357 , n66358 , n66359 , n66360 , 
 n66361 , n66362 , n66363 , n66364 , n66365 , n66366 , n66367 , n66368 , n66369 , n66370 , 
 n66371 , n66372 , n66373 , n66374 , n66375 , n66376 , n66377 , n66378 , n66379 , n66380 , 
 n66381 , n66382 , n66383 , n66384 , n66385 , n66386 , n66387 , n66388 , n66389 , n66390 , 
 n66391 , n66392 , n66393 , n66394 , n66395 , n66396 , n66397 , n66398 , n66399 , n66400 , 
 n66401 , n66402 , n66403 , n66404 , n66405 , n66406 , n66407 , n66408 , n66409 , n66410 , 
 n66411 , n66412 , n66413 , n66414 , n66415 , n66416 , n66417 , n66418 , n66419 , n66420 , 
 n66421 , n66422 , n66423 , n66424 , n66425 , n66426 , n66427 , n66428 , n66429 , n66430 , 
 n66431 , n66432 , n66433 , n66434 , n66435 , n66436 , n66437 , n66438 , n66439 , n66440 , 
 n66441 , n66442 , n66443 , n66444 , n66445 , n66446 , n66447 , n66448 , n66449 , n66450 , 
 n66451 , n66452 , n66453 , n66454 , n66455 , n66456 , n66457 , n66458 , n66459 , n66460 , 
 n66461 , n66462 , n66463 , n66464 , n66465 , n66466 , n66467 , n66468 , n66469 , n66470 , 
 n66471 , n66472 , n66473 , n66474 , n66475 , n66476 , n66477 , n66478 , n66479 , n66480 , 
 n66481 , n66482 , n66483 , n66484 , n66485 , n66486 , n66487 , n66488 , n66489 , n66490 , 
 n66491 , n66492 , n66493 , n66494 , n66495 , n66496 , n66497 , n66498 , n66499 , n66500 , 
 n66501 , n66502 , n66503 , n66504 , n66505 , n66506 , n66507 , n66508 , n66509 , n66510 , 
 n66511 , n66512 , n66513 , n66514 , n66515 , n66516 , n66517 , n66518 , n66519 , n66520 , 
 n66521 , n66522 , n66523 , n66524 , n66525 , n66526 , n66527 , n66528 , n66529 , n66530 , 
 n66531 , n66532 , n66533 , n66534 , n66535 , n66536 , n66537 , n66538 , n66539 , n66540 , 
 n66541 , n66542 , n66543 , n66544 , n66545 , n66546 , n66547 , n66548 , n66549 , n66550 , 
 n66551 , n66552 , n66553 , n66554 , n66555 , n66556 , n66557 , n66558 , n66559 , n66560 , 
 n66561 , n66562 , n66563 , n66564 , n66565 , n66566 , n66567 , n66568 , n66569 , n66570 , 
 n66571 , n66572 , n66573 , n66574 , n66575 , n66576 , n66577 , n66578 , n66579 , n66580 , 
 n66581 , n66582 , n66583 , n66584 , n66585 , n66586 , n66587 , n66588 , n66589 , n66590 , 
 n66591 , n66592 , n66593 , n66594 , n66595 , n66596 , n66597 , n66598 , n66599 , n66600 , 
 n66601 , n66602 , n66603 , n66604 , n66605 , n66606 , n66607 , n66608 , n66609 , n66610 , 
 n66611 , n66612 , n66613 , n66614 , n66615 , n66616 , n66617 , n66618 , n66619 , n66620 , 
 n66621 , n66622 , n66623 , n66624 , n66625 , n66626 , n66627 , n66628 , n66629 , n66630 , 
 n66631 , n66632 , n66633 , n66634 , n66635 , n66636 , n66637 , n66638 , n66639 , n66640 , 
 n66641 , n66642 , n66643 , n66644 , n66645 , n66646 , n66647 , n66648 , n66649 , n66650 , 
 n66651 , n66652 , n66653 , n66654 , n66655 , n66656 , n66657 , n66658 , n66659 , n66660 , 
 n66661 , n66662 , n66663 , n66664 , n66665 , n66666 , n66667 , n66668 , n66669 , n66670 , 
 n66671 , n66672 , n66673 , n66674 , n66675 , n66676 , n66677 , n66678 , n66679 , n66680 , 
 n66681 , n66682 , n66683 , n66684 , n66685 , n66686 , n66687 , n66688 , n66689 , n66690 , 
 n66691 , n66692 , n66693 , n66694 , n66695 , n66696 , n66697 , n66698 , n66699 , n66700 , 
 n66701 , n66702 , n66703 , n66704 , n66705 , n66706 , n66707 , n66708 , n66709 , n66710 , 
 n66711 , n66712 , n66713 , n66714 , n66715 , n66716 , n66717 , n66718 , n66719 , n66720 , 
 n66721 , n66722 , n66723 , n66724 , n66725 , n66726 , n66727 , n66728 , n66729 , n66730 , 
 n66731 , n66732 , n66733 , n66734 , n66735 , n66736 , n66737 , n66738 , n66739 , n66740 , 
 n66741 , n66742 , n66743 , n66744 , n66745 , n66746 , n66747 , n66748 , n66749 , n66750 , 
 n66751 , n66752 , n66753 , n66754 , n66755 , n66756 , n66757 , n66758 , n66759 , n66760 , 
 n66761 , n66762 , n66763 , n66764 , n66765 , n66766 , n66767 , n66768 , n66769 , n66770 , 
 n66771 , n66772 , n66773 , n66774 , n66775 , n66776 , n66777 , n66778 , n66779 , n66780 , 
 n66781 , n66782 , n66783 , n66784 , n66785 , n66786 , n66787 , n66788 , n66789 , n66790 , 
 n66791 , n66792 , n66793 , n66794 , n66795 , n66796 , n66797 , n66798 , n66799 , n66800 , 
 n66801 , n66802 , n66803 , n66804 , n66805 , n66806 , n66807 , n66808 , n66809 , n66810 , 
 n66811 , n66812 , n66813 , n66814 , n66815 , n66816 , n66817 , n66818 , n66819 , n66820 , 
 n66821 , n66822 , n66823 , n66824 , n66825 , n66826 , n66827 , n66828 , n66829 , n66830 , 
 n66831 , n66832 , n66833 , n66834 , n66835 , n66836 , n66837 , n66838 , n66839 , n66840 , 
 n66841 , n66842 , n66843 , n66844 , n66845 , n66846 , n66847 , n66848 , n66849 , n66850 , 
 n66851 , n66852 , n66853 , n66854 , n66855 , n66856 , n66857 , n66858 , n66859 , n66860 , 
 n66861 , n66862 , n66863 , n66864 , n66865 , n66866 , n66867 , n66868 , n66869 , n66870 , 
 n66871 , n66872 , n66873 , n66874 , n66875 , n66876 , n66877 , n66878 , n66879 , n66880 , 
 n66881 , n66882 , n66883 , n66884 , n66885 , n66886 , n66887 , n66888 , n66889 , n66890 , 
 n66891 , n66892 , n66893 , n66894 , n66895 , n66896 , n66897 , n66898 , n66899 , n66900 , 
 n66901 , n66902 , n66903 , n66904 , n66905 , n66906 , n66907 , n66908 , n66909 , n66910 , 
 n66911 , n66912 , n66913 , n66914 , n66915 , n66916 , n66917 , n66918 , n66919 , n66920 , 
 n66921 , n66922 , n66923 , n66924 , n66925 , n66926 , n66927 , n66928 , n66929 , n66930 , 
 n66931 , n66932 , n66933 , n66934 , n66935 , n66936 , n66937 , n66938 , n66939 , n66940 , 
 n66941 , n66942 , n66943 , n66944 , n66945 , n66946 , n66947 , n66948 , n66949 , n66950 , 
 n66951 , n66952 , n66953 , n66954 , n66955 , n66956 , n66957 , n66958 , n66959 , n66960 , 
 n66961 , n66962 , n66963 , n66964 , n66965 , n66966 , n66967 , n66968 , n66969 , n66970 , 
 n66971 , n66972 , n66973 , n66974 , n66975 , n66976 , n66977 , n66978 , n66979 , n66980 , 
 n66981 , n66982 , n66983 , n66984 , n66985 , n66986 , n66987 , n66988 , n66989 , n66990 , 
 n66991 , n66992 , n66993 , n66994 , n66995 , n66996 , n66997 , n66998 , n66999 , n67000 , 
 n67001 , n67002 , n67003 , n67004 , n67005 , n67006 , n67007 , n67008 , n67009 , n67010 , 
 n67011 , n67012 , n67013 , n67014 , n67015 , n67016 , n67017 , n67018 , n67019 , n67020 , 
 n67021 , n67022 , n67023 , n67024 , n67025 , n67026 , n67027 , n67028 , n67029 , n67030 , 
 n67031 , n67032 , n67033 , n67034 , n67035 , n67036 , n67037 , n67038 , n67039 , n67040 , 
 n67041 , n67042 , n67043 , n67044 , n67045 , n67046 , n67047 , n67048 , n67049 , n67050 , 
 n67051 , n67052 , n67053 , n67054 , n67055 , n67056 , n67057 , n67058 , n67059 , n67060 , 
 n67061 , n67062 , n67063 , n67064 , n67065 , n67066 , n67067 , n67068 , n67069 , n67070 , 
 n67071 , n67072 , n67073 , n67074 , n67075 , n67076 , n67077 , n67078 , n67079 , n67080 , 
 n67081 , n67082 , n67083 , n67084 , n67085 , n67086 , n67087 , n67088 , n67089 , n67090 , 
 n67091 , n67092 , n67093 , n67094 , n67095 , n67096 , n67097 , n67098 , n67099 , n67100 , 
 n67101 , n67102 , n67103 , n67104 , n67105 , n67106 , n67107 , n67108 , n67109 , n67110 , 
 n67111 , n67112 , n67113 , n67114 , n67115 , n67116 , n67117 , n67118 , n67119 , n67120 , 
 n67121 , n67122 , n67123 , n67124 , n67125 , n67126 , n67127 , n67128 , n67129 , n67130 , 
 n67131 , n67132 , n67133 , n67134 , n67135 , n67136 , n67137 , n67138 , n67139 , n67140 , 
 n67141 , n67142 , n67143 , n67144 , n67145 , n67146 , n67147 , n67148 , n67149 , n67150 , 
 n67151 , n67152 , n67153 , n67154 , n67155 , n67156 , n67157 , n67158 , n67159 , n67160 , 
 n67161 , n67162 , n67163 , n67164 , n67165 , n67166 , n67167 , n67168 , n67169 , n67170 , 
 n67171 , n67172 , n67173 , n67174 , n67175 , n67176 , n67177 , n67178 , n67179 , n67180 , 
 n67181 , n67182 , n67183 , n67184 , n67185 , n67186 , n67187 , n67188 , n67189 , n67190 , 
 n67191 , n67192 , n67193 , n67194 , n67195 , n67196 , n67197 , n67198 , n67199 , n67200 , 
 n67201 , n67202 , n67203 , n67204 , n67205 , n67206 , n67207 , n67208 , n67209 , n67210 , 
 n67211 , n67212 , n67213 , n67214 , n67215 , n67216 , n67217 , n67218 , n67219 , n67220 , 
 n67221 , n67222 , n67223 , n67224 , n67225 , n67226 , n67227 , n67228 , n67229 , n67230 , 
 n67231 , n67232 , n67233 , n67234 , n67235 , n67236 , n67237 , n67238 , n67239 , n67240 , 
 n67241 , n67242 , n67243 , n67244 , n67245 , n67246 , n67247 , n67248 , n67249 , n67250 , 
 n67251 , n67252 , n67253 , n67254 , n67255 , n67256 , n67257 , n67258 , n67259 , n67260 , 
 n67261 , n67262 , n67263 , n67264 , n67265 , n67266 , n67267 , n67268 , n67269 , n67270 , 
 n67271 , n67272 , n67273 , n67274 , n67275 , n67276 , n67277 , n67278 , n67279 , n67280 , 
 n67281 , n67282 , n67283 , n67284 , n67285 , n67286 , n67287 , n67288 , n67289 , n67290 , 
 n67291 , n67292 , n67293 , n67294 , n67295 , n67296 , n67297 , n67298 , n67299 , n67300 , 
 n67301 , n67302 , n67303 , n67304 , n67305 , n67306 , n67307 , n67308 , n67309 , n67310 , 
 n67311 , n67312 , n67313 , n67314 , n67315 , n67316 , n67317 , n67318 , n67319 , n67320 , 
 n67321 , n67322 , n67323 , n67324 , n67325 , n67326 , n67327 , n67328 , n67329 , n67330 , 
 n67331 , n67332 , n67333 , n67334 , n67335 , n67336 , n67337 , n67338 , n67339 , n67340 , 
 n67341 , n67342 , n67343 , n67344 , n67345 , n67346 , n67347 , n67348 , n67349 , n67350 , 
 n67351 , n67352 , n67353 , n67354 , n67355 , n67356 , n67357 , n67358 , n67359 , n67360 , 
 n67361 , n67362 , n67363 , n67364 , n67365 , n67366 , n67367 , n67368 , n67369 , n67370 , 
 n67371 , n67372 , n67373 , n67374 , n67375 , n67376 , n67377 , n67378 , n67379 , n67380 , 
 n67381 , n67382 , n67383 , n67384 , n67385 , n67386 , n67387 , n67388 , n67389 , n67390 , 
 n67391 , n67392 , n67393 , n67394 , n67395 , n67396 , n67397 , n67398 , n67399 , n67400 , 
 n67401 , n67402 , n67403 , n67404 , n67405 , n67406 , n67407 , n67408 , n67409 , n67410 , 
 n67411 , n67412 , n67413 , n67414 , n67415 , n67416 , n67417 , n67418 , n67419 , n67420 , 
 n67421 , n67422 , n67423 , n67424 , n67425 , n67426 , n67427 , n67428 , n67429 , n67430 , 
 n67431 , n67432 , n67433 , n67434 , n67435 , n67436 , n67437 , n67438 , n67439 , n67440 , 
 n67441 , n67442 , n67443 , n67444 , n67445 , n67446 , n67447 , n67448 , n67449 , n67450 , 
 n67451 , n67452 , n67453 , n67454 , n67455 , n67456 , n67457 , n67458 , n67459 , n67460 , 
 n67461 , n67462 , n67463 , n67464 , n67465 , n67466 , n67467 , n67468 , n67469 , n67470 , 
 n67471 , n67472 , n67473 , n67474 , n67475 , n67476 , n67477 , n67478 , n67479 , n67480 , 
 n67481 , n67482 , n67483 , n67484 , n67485 , n67486 , n67487 , n67488 , n67489 , n67490 , 
 n67491 , n67492 , n67493 , n67494 , n67495 , n67496 , n67497 , n67498 , n67499 , n67500 , 
 n67501 , n67502 , n67503 , n67504 , n67505 , n67506 , n67507 , n67508 , n67509 , n67510 , 
 n67511 , n67512 , n67513 , n67514 , n67515 , n67516 , n67517 , n67518 , n67519 , n67520 , 
 n67521 , n67522 , n67523 , n67524 , n67525 , n67526 , n67527 , n67528 , n67529 , n67530 , 
 n67531 , n67532 , n67533 , n67534 , n67535 , n67536 , n67537 , n67538 , n67539 , n67540 , 
 n67541 , n67542 , n67543 , n67544 , n67545 , n67546 , n67547 , n67548 , n67549 , n67550 , 
 n67551 , n67552 , n67553 , n67554 , n67555 , n67556 , n67557 , n67558 , n67559 , n67560 , 
 n67561 , n67562 , n67563 , n67564 , n67565 , n67566 , n67567 , n67568 , n67569 , n67570 , 
 n67571 , n67572 , n67573 , n67574 , n67575 , n67576 , n67577 , n67578 , n67579 , n67580 , 
 n67581 , n67582 , n67583 , n67584 , n67585 , n67586 , n67587 , n67588 , n67589 , n67590 , 
 n67591 , n67592 , n67593 , n67594 , n67595 , n67596 , n67597 , n67598 , n67599 , n67600 , 
 n67601 , n67602 , n67603 , n67604 , n67605 , n67606 , n67607 , n67608 , n67609 , n67610 , 
 n67611 , n67612 , n67613 , n67614 , n67615 , n67616 , n67617 , n67618 , n67619 , n67620 , 
 n67621 , n67622 , n67623 , n67624 , n67625 , n67626 , n67627 , n67628 , n67629 , n67630 , 
 n67631 , n67632 , n67633 , n67634 , n67635 , n67636 , n67637 , n67638 , n67639 , n67640 , 
 n67641 , n67642 , n67643 , n67644 , n67645 , n67646 , n67647 , n67648 , n67649 , n67650 , 
 n67651 , n67652 , n67653 , n67654 , n67655 , n67656 , n67657 , n67658 , n67659 , n67660 , 
 n67661 , n67662 , n67663 , n67664 , n67665 , n67666 , n67667 , n67668 , n67669 , n67670 , 
 n67671 , n67672 , n67673 , n67674 , n67675 , n67676 , n67677 , n67678 , n67679 , n67680 , 
 n67681 , n67682 , n67683 , n67684 , n67685 , n67686 , n67687 , n67688 , n67689 , n67690 , 
 n67691 , n67692 , n67693 , n67694 , n67695 , n67696 , n67697 , n67698 , n67699 , n67700 , 
 n67701 , n67702 , n67703 , n67704 , n67705 , n67706 , n67707 , n67708 , n67709 , n67710 , 
 n67711 , n67712 , n67713 , n67714 , n67715 , n67716 , n67717 , n67718 , n67719 , n67720 , 
 n67721 , n67722 , n67723 , n67724 , n67725 , n67726 , n67727 , n67728 , n67729 , n67730 , 
 n67731 , n67732 , n67733 , n67734 , n67735 , n67736 , n67737 , n67738 , n67739 , n67740 , 
 n67741 , n67742 , n67743 , n67744 , n67745 , n67746 , n67747 , n67748 , n67749 , n67750 , 
 n67751 , n67752 , n67753 , n67754 , n67755 , n67756 , n67757 , n67758 , n67759 , n67760 , 
 n67761 , n67762 , n67763 , n67764 , n67765 , n67766 , n67767 , n67768 , n67769 , n67770 , 
 n67771 , n67772 , n67773 , n67774 , n67775 , n67776 , n67777 , n67778 , n67779 , n67780 , 
 n67781 , n67782 , n67783 , n67784 , n67785 , n67786 , n67787 , n67788 , n67789 , n67790 , 
 n67791 , n67792 , n67793 , n67794 , n67795 , n67796 , n67797 , n67798 , n67799 , n67800 , 
 n67801 , n67802 , n67803 , n67804 , n67805 , n67806 , n67807 , n67808 , n67809 , n67810 , 
 n67811 , n67812 , n67813 , n67814 , n67815 , n67816 , n67817 , n67818 , n67819 , n67820 , 
 n67821 , n67822 , n67823 , n67824 , n67825 , n67826 , n67827 , n67828 , n67829 , n67830 , 
 n67831 , n67832 , n67833 , n67834 , n67835 , n67836 , n67837 , n67838 , n67839 , n67840 , 
 n67841 , n67842 , n67843 , n67844 , n67845 , n67846 , n67847 , n67848 , n67849 , n67850 , 
 n67851 , n67852 , n67853 , n67854 , n67855 , n67856 , n67857 , n67858 , n67859 , n67860 , 
 n67861 , n67862 , n67863 , n67864 , n67865 , n67866 , n67867 , n67868 , n67869 , n67870 , 
 n67871 , n67872 , n67873 , n67874 , n67875 , n67876 , n67877 , n67878 , n67879 , n67880 , 
 n67881 , n67882 , n67883 , n67884 , n67885 , n67886 , n67887 , n67888 , n67889 , n67890 , 
 n67891 , n67892 , n67893 , n67894 , n67895 , n67896 , n67897 , n67898 , n67899 , n67900 , 
 n67901 , n67902 , n67903 , n67904 , n67905 , n67906 , n67907 , n67908 , n67909 , n67910 , 
 n67911 , n67912 , n67913 , n67914 , n67915 , n67916 , n67917 , n67918 , n67919 , n67920 , 
 n67921 , n67922 , n67923 , n67924 , n67925 , n67926 , n67927 , n67928 , n67929 , n67930 , 
 n67931 , n67932 , n67933 , n67934 , n67935 , n67936 , n67937 , n67938 , n67939 , n67940 , 
 n67941 , n67942 , n67943 , n67944 , n67945 , n67946 , n67947 , n67948 , n67949 , n67950 , 
 n67951 , n67952 , n67953 , n67954 , n67955 , n67956 , n67957 , n67958 , n67959 , n67960 , 
 n67961 , n67962 , n67963 , n67964 , n67965 , n67966 , n67967 , n67968 , n67969 , n67970 , 
 n67971 , n67972 , n67973 , n67974 , n67975 , n67976 , n67977 , n67978 , n67979 , n67980 , 
 n67981 , n67982 , n67983 , n67984 , n67985 , n67986 , n67987 , n67988 , n67989 , n67990 , 
 n67991 , n67992 , n67993 , n67994 , n67995 , n67996 , n67997 , n67998 , n67999 , n68000 , 
 n68001 , n68002 , n68003 , n68004 , n68005 , n68006 , n68007 , n68008 , n68009 , n68010 , 
 n68011 , n68012 , n68013 , n68014 , n68015 , n68016 , n68017 , n68018 , n68019 , n68020 , 
 n68021 , n68022 , n68023 , n68024 , n68025 , n68026 , n68027 , n68028 , n68029 , n68030 , 
 n68031 , n68032 , n68033 , n68034 , n68035 , n68036 , n68037 , n68038 , n68039 , n68040 , 
 n68041 , n68042 , n68043 , n68044 , n68045 , n68046 , n68047 , n68048 , n68049 , n68050 , 
 n68051 , n68052 , n68053 , n68054 , n68055 , n68056 , n68057 , n68058 , n68059 , n68060 , 
 n68061 , n68062 , n68063 , n68064 , n68065 , n68066 , n68067 , n68068 , n68069 , n68070 , 
 n68071 , n68072 , n68073 , n68074 , n68075 , n68076 , n68077 , n68078 , n68079 , n68080 , 
 n68081 , n68082 , n68083 , n68084 , n68085 , n68086 , n68087 , n68088 , n68089 , n68090 , 
 n68091 , n68092 , n68093 , n68094 , n68095 , n68096 , n68097 , n68098 , n68099 , n68100 , 
 n68101 , n68102 , n68103 , n68104 , n68105 , n68106 , n68107 , n68108 , n68109 , n68110 , 
 n68111 , n68112 , n68113 , n68114 , n68115 , n68116 , n68117 , n68118 , n68119 , n68120 , 
 n68121 , n68122 , n68123 , n68124 , n68125 , n68126 , n68127 , n68128 , n68129 , n68130 , 
 n68131 , n68132 , n68133 , n68134 , n68135 , n68136 , n68137 , n68138 , n68139 , n68140 , 
 n68141 , n68142 , n68143 , n68144 , n68145 , n68146 , n68147 , n68148 , n68149 , n68150 , 
 n68151 , n68152 , n68153 , n68154 , n68155 , n68156 , n68157 , n68158 , n68159 , n68160 , 
 n68161 , n68162 , n68163 , n68164 , n68165 , n68166 , n68167 , n68168 , n68169 , n68170 , 
 n68171 , n68172 , n68173 , n68174 , n68175 , n68176 , n68177 , n68178 , n68179 , n68180 , 
 n68181 , n68182 , n68183 , n68184 , n68185 , n68186 , n68187 , n68188 , n68189 , n68190 , 
 n68191 , n68192 , n68193 , n68194 , n68195 , n68196 , n68197 , n68198 , n68199 , n68200 , 
 n68201 , n68202 , n68203 , n68204 , n68205 , n68206 , n68207 , n68208 , n68209 , n68210 , 
 n68211 , n68212 , n68213 , n68214 , n68215 , n68216 , n68217 , n68218 , n68219 , n68220 , 
 n68221 , n68222 , n68223 , n68224 , n68225 , n68226 , n68227 , n68228 , n68229 , n68230 , 
 n68231 , n68232 , n68233 , n68234 , n68235 , n68236 , n68237 , n68238 , n68239 , n68240 , 
 n68241 , n68242 , n68243 , n68244 , n68245 , n68246 , n68247 , n68248 , n68249 , n68250 , 
 n68251 , n68252 , n68253 , n68254 , n68255 , n68256 , n68257 , n68258 , n68259 , n68260 , 
 n68261 , n68262 , n68263 , n68264 , n68265 , n68266 , n68267 , n68268 , n68269 , n68270 , 
 n68271 , n68272 , n68273 , n68274 , n68275 , n68276 , n68277 , n68278 , n68279 , n68280 , 
 n68281 , n68282 , n68283 , n68284 , n68285 , n68286 , n68287 , n68288 , n68289 , n68290 , 
 n68291 , n68292 , n68293 , n68294 , n68295 , n68296 , n68297 , n68298 , n68299 , n68300 , 
 n68301 , n68302 , n68303 , n68304 , n68305 , n68306 , n68307 , n68308 , n68309 , n68310 , 
 n68311 , n68312 , n68313 , n68314 , n68315 , n68316 , n68317 , n68318 , n68319 , n68320 , 
 n68321 , n68322 , n68323 , n68324 , n68325 , n68326 , n68327 , n68328 , n68329 , n68330 , 
 n68331 , n68332 , n68333 , n68334 , n68335 , n68336 , n68337 , n68338 , n68339 , n68340 , 
 n68341 , n68342 , n68343 , n68344 , n68345 , n68346 , n68347 , n68348 , n68349 , n68350 , 
 n68351 , n68352 , n68353 , n68354 , n68355 , n68356 , n68357 , n68358 , n68359 , n68360 , 
 n68361 , n68362 , n68363 , n68364 , n68365 , n68366 , n68367 , n68368 , n68369 , n68370 , 
 n68371 , n68372 , n68373 , n68374 , n68375 , n68376 , n68377 , n68378 , n68379 , n68380 , 
 n68381 , n68382 , n68383 , n68384 , n68385 , n68386 , n68387 , n68388 , n68389 , n68390 , 
 n68391 , n68392 , n68393 , n68394 , n68395 , n68396 , n68397 , n68398 , n68399 , n68400 , 
 n68401 , n68402 , n68403 , n68404 , n68405 , n68406 , n68407 , n68408 , n68409 , n68410 , 
 n68411 , n68412 , n68413 , n68414 , n68415 , n68416 , n68417 , n68418 , n68419 , n68420 , 
 n68421 , n68422 , n68423 , n68424 , n68425 , n68426 , n68427 , n68428 , n68429 , n68430 , 
 n68431 , n68432 , n68433 , n68434 , n68435 , n68436 , n68437 , n68438 , n68439 , n68440 , 
 n68441 , n68442 , n68443 , n68444 , n68445 , n68446 , n68447 , n68448 , n68449 , n68450 , 
 n68451 , n68452 , n68453 , n68454 , n68455 , n68456 , n68457 , n68458 , n68459 , n68460 , 
 n68461 , n68462 , n68463 , n68464 , n68465 , n68466 , n68467 , n68468 , n68469 , n68470 , 
 n68471 , n68472 , n68473 , n68474 , n68475 , n68476 , n68477 , n68478 , n68479 , n68480 , 
 n68481 , n68482 , n68483 , n68484 , n68485 , n68486 , n68487 , n68488 , n68489 , n68490 , 
 n68491 , n68492 , n68493 , n68494 , n68495 , n68496 , n68497 , n68498 , n68499 , n68500 , 
 n68501 , n68502 , n68503 , n68504 , n68505 , n68506 , n68507 , n68508 , n68509 , n68510 , 
 n68511 , n68512 , n68513 , n68514 , n68515 , n68516 , n68517 , n68518 , n68519 , n68520 , 
 n68521 , n68522 , n68523 , n68524 , n68525 , n68526 , n68527 , n68528 , n68529 , n68530 , 
 n68531 , n68532 , n68533 , n68534 , n68535 , n68536 , n68537 , n68538 , n68539 , n68540 , 
 n68541 , n68542 , n68543 , n68544 , n68545 , n68546 , n68547 , n68548 , n68549 , n68550 , 
 n68551 , n68552 , n68553 , n68554 , n68555 , n68556 , n68557 , n68558 , n68559 , n68560 , 
 n68561 , n68562 , n68563 , n68564 , n68565 , n68566 , n68567 , n68568 , n68569 , n68570 , 
 n68571 , n68572 , n68573 , n68574 , n68575 , n68576 , n68577 , n68578 , n68579 , n68580 , 
 n68581 , n68582 , n68583 , n68584 , n68585 , n68586 , n68587 , n68588 , n68589 , n68590 , 
 n68591 , n68592 , n68593 , n68594 , n68595 , n68596 , n68597 , n68598 , n68599 , n68600 , 
 n68601 , n68602 , n68603 , n68604 , n68605 , n68606 , n68607 , n68608 , n68609 , n68610 , 
 n68611 , n68612 , n68613 , n68614 , n68615 , n68616 , n68617 , n68618 , n68619 , n68620 , 
 n68621 , n68622 , n68623 , n68624 , n68625 , n68626 , n68627 , n68628 , n68629 , n68630 , 
 n68631 , n68632 , n68633 , n68634 , n68635 , n68636 , n68637 , n68638 , n68639 , n68640 , 
 n68641 , n68642 , n68643 , n68644 , n68645 , n68646 , n68647 , n68648 , n68649 , n68650 , 
 n68651 , n68652 , n68653 , n68654 , n68655 , n68656 , n68657 , n68658 , n68659 , n68660 , 
 n68661 , n68662 , n68663 , n68664 , n68665 , n68666 , n68667 , n68668 , n68669 , n68670 , 
 n68671 , n68672 , n68673 , n68674 , n68675 , n68676 , n68677 , n68678 , n68679 , n68680 , 
 n68681 , n68682 , n68683 , n68684 , n68685 , n68686 , n68687 , n68688 , n68689 , n68690 , 
 n68691 , n68692 , n68693 , n68694 , n68695 , n68696 , n68697 , n68698 , n68699 , n68700 , 
 n68701 , n68702 , n68703 , n68704 , n68705 , n68706 , n68707 , n68708 , n68709 , n68710 , 
 n68711 , n68712 , n68713 , n68714 , n68715 , n68716 , n68717 , n68718 , n68719 , n68720 , 
 n68721 , n68722 , n68723 , n68724 , n68725 , n68726 , n68727 , n68728 , n68729 , n68730 , 
 n68731 , n68732 , n68733 , n68734 , n68735 , n68736 , n68737 , n68738 , n68739 , n68740 , 
 n68741 , n68742 , n68743 , n68744 , n68745 , n68746 , n68747 , n68748 , n68749 , n68750 , 
 n68751 , n68752 , n68753 , n68754 , n68755 , n68756 , n68757 , n68758 , n68759 , n68760 , 
 n68761 , n68762 , n68763 , n68764 , n68765 , n68766 , n68767 , n68768 , n68769 , n68770 , 
 n68771 , n68772 , n68773 , n68774 , n68775 , n68776 , n68777 , n68778 , n68779 , n68780 , 
 n68781 , n68782 , n68783 , n68784 , n68785 , n68786 , n68787 , n68788 , n68789 , n68790 , 
 n68791 , n68792 , n68793 , n68794 , n68795 , n68796 , n68797 , n68798 , n68799 , n68800 , 
 n68801 , n68802 , n68803 , n68804 , n68805 , n68806 , n68807 , n68808 , n68809 , n68810 , 
 n68811 , n68812 , n68813 , n68814 , n68815 , n68816 , n68817 , n68818 , n68819 , n68820 , 
 n68821 , n68822 , n68823 , n68824 , n68825 , n68826 , n68827 , n68828 , n68829 , n68830 , 
 n68831 , n68832 , n68833 , n68834 , n68835 , n68836 , n68837 , n68838 , n68839 , n68840 , 
 n68841 , n68842 , n68843 , n68844 , n68845 , n68846 , n68847 , n68848 , n68849 , n68850 , 
 n68851 , n68852 , n68853 , n68854 , n68855 , n68856 , n68857 , n68858 , n68859 , n68860 , 
 n68861 , n68862 , n68863 , n68864 , n68865 , n68866 , n68867 , n68868 , n68869 , n68870 , 
 n68871 , n68872 , n68873 , n68874 , n68875 , n68876 , n68877 , n68878 , n68879 , n68880 , 
 n68881 , n68882 , n68883 , n68884 , n68885 , n68886 , n68887 , n68888 , n68889 , n68890 , 
 n68891 , n68892 , n68893 , n68894 , n68895 , n68896 , n68897 , n68898 , n68899 , n68900 , 
 n68901 , n68902 , n68903 , n68904 , n68905 , n68906 , n68907 , n68908 , n68909 , n68910 , 
 n68911 , n68912 , n68913 , n68914 , n68915 , n68916 , n68917 , n68918 , n68919 , n68920 , 
 n68921 , n68922 , n68923 , n68924 , n68925 , n68926 , n68927 , n68928 , n68929 , n68930 , 
 n68931 , n68932 , n68933 , n68934 , n68935 , n68936 , n68937 , n68938 , n68939 , n68940 , 
 n68941 , n68942 , n68943 , n68944 , n68945 , n68946 , n68947 , n68948 , n68949 , n68950 , 
 n68951 , n68952 , n68953 , n68954 , n68955 , n68956 , n68957 , n68958 , n68959 , n68960 , 
 n68961 , n68962 , n68963 , n68964 , n68965 , n68966 , n68967 , n68968 , n68969 , n68970 , 
 n68971 , n68972 , n68973 , n68974 , n68975 , n68976 , n68977 , n68978 , n68979 , n68980 , 
 n68981 , n68982 , n68983 , n68984 , n68985 , n68986 , n68987 , n68988 , n68989 , n68990 , 
 n68991 , n68992 , n68993 , n68994 , n68995 , n68996 , n68997 , n68998 , n68999 , n69000 , 
 n69001 , n69002 , n69003 , n69004 , n69005 , n69006 , n69007 , n69008 , n69009 , n69010 , 
 n69011 , n69012 , n69013 , n69014 , n69015 , n69016 , n69017 , n69018 , n69019 , n69020 , 
 n69021 , n69022 , n69023 , n69024 , n69025 , n69026 , n69027 , n69028 , n69029 , n69030 , 
 n69031 , n69032 , n69033 , n69034 , n69035 , n69036 , n69037 , n69038 , n69039 , n69040 , 
 n69041 , n69042 , n69043 , n69044 , n69045 , n69046 , n69047 , n69048 , n69049 , n69050 , 
 n69051 , n69052 , n69053 , n69054 , n69055 , n69056 , n69057 , n69058 , n69059 , n69060 , 
 n69061 , n69062 , n69063 , n69064 , n69065 , n69066 , n69067 , n69068 , n69069 , n69070 , 
 n69071 , n69072 , n69073 , n69074 , n69075 , n69076 , n69077 , n69078 , n69079 , n69080 , 
 n69081 , n69082 , n69083 , n69084 , n69085 , n69086 , n69087 , n69088 , n69089 , n69090 , 
 n69091 , n69092 , n69093 , n69094 , n69095 , n69096 , n69097 , n69098 , n69099 , n69100 , 
 n69101 , n69102 , n69103 , n69104 , n69105 , n69106 , n69107 , n69108 , n69109 , n69110 , 
 n69111 , n69112 , n69113 , n69114 , n69115 , n69116 , n69117 , n69118 , n69119 , n69120 , 
 n69121 , n69122 , n69123 , n69124 , n69125 , n69126 , n69127 , n69128 , n69129 , n69130 , 
 n69131 , n69132 , n69133 , n69134 , n69135 , n69136 , n69137 , n69138 , n69139 , n69140 , 
 n69141 , n69142 , n69143 , n69144 , n69145 , n69146 , n69147 , n69148 , n69149 , n69150 , 
 n69151 , n69152 , n69153 , n69154 , n69155 , n69156 , n69157 , n69158 , n69159 , n69160 , 
 n69161 , n69162 , n69163 , n69164 , n69165 , n69166 , n69167 , n69168 , n69169 , n69170 , 
 n69171 , n69172 , n69173 , n69174 , n69175 , n69176 , n69177 , n69178 , n69179 , n69180 , 
 n69181 , n69182 , n69183 , n69184 , n69185 , n69186 , n69187 , n69188 , n69189 , n69190 , 
 n69191 , n69192 , n69193 , n69194 , n69195 , n69196 , n69197 , n69198 , n69199 , n69200 , 
 n69201 , n69202 , n69203 , n69204 , n69205 , n69206 , n69207 , n69208 , n69209 , n69210 , 
 n69211 , n69212 , n69213 , n69214 , n69215 , n69216 , n69217 , n69218 , n69219 , n69220 , 
 n69221 , n69222 , n69223 , n69224 , n69225 , n69226 , n69227 , n69228 , n69229 , n69230 , 
 n69231 , n69232 , n69233 , n69234 , n69235 , n69236 , n69237 , n69238 , n69239 , n69240 , 
 n69241 , n69242 , n69243 , n69244 , n69245 , n69246 , n69247 , n69248 , n69249 , n69250 , 
 n69251 , n69252 , n69253 , n69254 , n69255 , n69256 , n69257 , n69258 , n69259 , n69260 , 
 n69261 , n69262 , n69263 , n69264 , n69265 , n69266 , n69267 , n69268 , n69269 , n69270 , 
 n69271 , n69272 , n69273 , n69274 , n69275 , n69276 , n69277 , n69278 , n69279 , n69280 , 
 n69281 , n69282 , n69283 , n69284 , n69285 , n69286 , n69287 , n69288 , n69289 , n69290 , 
 n69291 , n69292 , n69293 , n69294 , n69295 , n69296 , n69297 , n69298 , n69299 , n69300 , 
 n69301 , n69302 , n69303 , n69304 , n69305 , n69306 , n69307 , n69308 , n69309 , n69310 , 
 n69311 , n69312 , n69313 , n69314 , n69315 , n69316 , n69317 , n69318 , n69319 , n69320 , 
 n69321 , n69322 , n69323 , n69324 , n69325 , n69326 , n69327 , n69328 , n69329 , n69330 , 
 n69331 , n69332 , n69333 , n69334 , n69335 , n69336 , n69337 , n69338 , n69339 , n69340 , 
 n69341 , n69342 , n69343 , n69344 , n69345 , n69346 , n69347 , n69348 , n69349 , n69350 , 
 n69351 , n69352 , n69353 , n69354 , n69355 , n69356 , n69357 , n69358 , n69359 , n69360 , 
 n69361 , n69362 , n69363 , n69364 , n69365 , n69366 , n69367 , n69368 , n69369 , n69370 , 
 n69371 , n69372 , n69373 , n69374 , n69375 , n69376 , n69377 , n69378 , n69379 , n69380 , 
 n69381 , n69382 , n69383 , n69384 , n69385 , n69386 , n69387 , n69388 , n69389 , n69390 , 
 n69391 , n69392 , n69393 , n69394 , n69395 , n69396 , n69397 , n69398 , n69399 , n69400 , 
 n69401 , n69402 , n69403 , n69404 , n69405 , n69406 , n69407 , n69408 , n69409 , n69410 , 
 n69411 , n69412 , n69413 , n69414 , n69415 , n69416 , n69417 , n69418 , n69419 , n69420 , 
 n69421 , n69422 , n69423 , n69424 , n69425 , n69426 , n69427 , n69428 , n69429 , n69430 , 
 n69431 , n69432 , n69433 , n69434 , n69435 , n69436 , n69437 , n69438 , n69439 , n69440 , 
 n69441 , n69442 , n69443 , n69444 , n69445 , n69446 , n69447 , n69448 , n69449 , n69450 , 
 n69451 , n69452 , n69453 , n69454 , n69455 , n69456 , n69457 , n69458 , n69459 , n69460 , 
 n69461 , n69462 , n69463 , n69464 , n69465 , n69466 , n69467 , n69468 , n69469 , n69470 , 
 n69471 , n69472 , n69473 , n69474 , n69475 , n69476 , n69477 , n69478 , n69479 , n69480 , 
 n69481 , n69482 , n69483 , n69484 , n69485 , n69486 , n69487 , n69488 , n69489 , n69490 , 
 n69491 , n69492 , n69493 , n69494 , n69495 , n69496 , n69497 , n69498 , n69499 , n69500 , 
 n69501 , n69502 , n69503 , n69504 , n69505 , n69506 , n69507 , n69508 , n69509 , n69510 , 
 n69511 , n69512 , n69513 , n69514 , n69515 , n69516 , n69517 , n69518 , n69519 , n69520 , 
 n69521 , n69522 , n69523 , n69524 , n69525 , n69526 , n69527 , n69528 , n69529 , n69530 , 
 n69531 , n69532 , n69533 , n69534 , n69535 , n69536 , n69537 , n69538 , n69539 , n69540 , 
 n69541 , n69542 , n69543 , n69544 , n69545 , n69546 , n69547 , n69548 , n69549 , n69550 , 
 n69551 , n69552 , n69553 , n69554 , n69555 , n69556 , n69557 , n69558 , n69559 , n69560 , 
 n69561 , n69562 , n69563 , n69564 , n69565 , n69566 , n69567 , n69568 , n69569 , n69570 , 
 n69571 , n69572 , n69573 , n69574 , n69575 , n69576 , n69577 , n69578 , n69579 , n69580 , 
 n69581 , n69582 , n69583 , n69584 , n69585 , n69586 , n69587 , n69588 , n69589 , n69590 , 
 n69591 , n69592 , n69593 , n69594 , n69595 , n69596 , n69597 , n69598 , n69599 , n69600 , 
 n69601 , n69602 , n69603 , n69604 , n69605 , n69606 , n69607 , n69608 , n69609 , n69610 , 
 n69611 , n69612 , n69613 , n69614 , n69615 , n69616 , n69617 , n69618 , n69619 , n69620 , 
 n69621 , n69622 , n69623 , n69624 , n69625 , n69626 , n69627 , n69628 , n69629 , n69630 , 
 n69631 , n69632 , n69633 , n69634 , n69635 , n69636 , n69637 , n69638 , n69639 , n69640 , 
 n69641 , n69642 , n69643 , n69644 , n69645 , n69646 , n69647 , n69648 , n69649 , n69650 , 
 n69651 , n69652 , n69653 , n69654 , n69655 , n69656 , n69657 , n69658 , n69659 , n69660 , 
 n69661 , n69662 , n69663 , n69664 , n69665 , n69666 , n69667 , n69668 , n69669 , n69670 , 
 n69671 , n69672 , n69673 , n69674 , n69675 , n69676 , n69677 , n69678 , n69679 , n69680 , 
 n69681 , n69682 , n69683 , n69684 , n69685 , n69686 , n69687 , n69688 , n69689 , n69690 , 
 n69691 , n69692 , n69693 , n69694 , n69695 , n69696 , n69697 , n69698 , n69699 , n69700 , 
 n69701 , n69702 , n69703 , n69704 , n69705 , n69706 , n69707 , n69708 , n69709 , n69710 , 
 n69711 , n69712 , n69713 , n69714 , n69715 , n69716 , n69717 , n69718 , n69719 , n69720 , 
 n69721 , n69722 , n69723 , n69724 , n69725 , n69726 , n69727 , n69728 , n69729 , n69730 , 
 n69731 , n69732 , n69733 , n69734 , n69735 , n69736 , n69737 , n69738 , n69739 , n69740 , 
 n69741 , n69742 , n69743 , n69744 , n69745 , n69746 , n69747 , n69748 , n69749 , n69750 , 
 n69751 , n69752 , n69753 , n69754 , n69755 , n69756 , n69757 , n69758 , n69759 , n69760 , 
 n69761 , n69762 , n69763 , n69764 , n69765 , n69766 , n69767 , n69768 , n69769 , n69770 , 
 n69771 , n69772 , n69773 , n69774 , n69775 , n69776 , n69777 , n69778 , n69779 , n69780 , 
 n69781 , n69782 , n69783 , n69784 , n69785 , n69786 , n69787 , n69788 , n69789 , n69790 , 
 n69791 , n69792 , n69793 , n69794 , n69795 , n69796 , n69797 , n69798 , n69799 , n69800 , 
 n69801 , n69802 , n69803 , n69804 , n69805 , n69806 , n69807 , n69808 , n69809 , n69810 , 
 n69811 , n69812 , n69813 , n69814 , n69815 , n69816 , n69817 , n69818 , n69819 , n69820 , 
 n69821 , n69822 , n69823 , n69824 , n69825 , n69826 , n69827 , n69828 , n69829 , n69830 , 
 n69831 , n69832 , n69833 , n69834 , n69835 , n69836 , n69837 , n69838 , n69839 , n69840 , 
 n69841 , n69842 , n69843 , n69844 , n69845 , n69846 , n69847 , n69848 , n69849 , n69850 , 
 n69851 , n69852 , n69853 , n69854 , n69855 , n69856 , n69857 , n69858 , n69859 , n69860 , 
 n69861 , n69862 , n69863 , n69864 , n69865 , n69866 , n69867 , n69868 , n69869 , n69870 , 
 n69871 , n69872 , n69873 , n69874 , n69875 , n69876 , n69877 , n69878 , n69879 , n69880 , 
 n69881 , n69882 , n69883 , n69884 , n69885 , n69886 , n69887 , n69888 , n69889 , n69890 , 
 n69891 , n69892 , n69893 , n69894 , n69895 , n69896 , n69897 , n69898 , n69899 , n69900 , 
 n69901 , n69902 , n69903 , n69904 , n69905 , n69906 , n69907 , n69908 , n69909 , n69910 , 
 n69911 , n69912 , n69913 , n69914 , n69915 , n69916 , n69917 , n69918 , n69919 , n69920 , 
 n69921 , n69922 , n69923 , n69924 , n69925 , n69926 , n69927 , n69928 , n69929 , n69930 , 
 n69931 , n69932 , n69933 , n69934 , n69935 , n69936 , n69937 , n69938 , n69939 , n69940 , 
 n69941 , n69942 , n69943 , n69944 , n69945 , n69946 , n69947 , n69948 , n69949 , n69950 , 
 n69951 , n69952 , n69953 , n69954 , n69955 , n69956 , n69957 , n69958 , n69959 , n69960 , 
 n69961 , n69962 , n69963 , n69964 , n69965 , n69966 , n69967 , n69968 , n69969 , n69970 , 
 n69971 , n69972 , n69973 , n69974 , n69975 , n69976 , n69977 , n69978 , n69979 , n69980 , 
 n69981 , n69982 , n69983 , n69984 , n69985 , n69986 , n69987 , n69988 , n69989 , n69990 , 
 n69991 , n69992 , n69993 , n69994 , n69995 , n69996 , n69997 , n69998 , n69999 , n70000 , 
 n70001 , n70002 , n70003 , n70004 , n70005 , n70006 , n70007 , n70008 , n70009 , n70010 , 
 n70011 , n70012 , n70013 , n70014 , n70015 , n70016 , n70017 , n70018 , n70019 , n70020 , 
 n70021 , n70022 , n70023 , n70024 , n70025 , n70026 , n70027 , n70028 , n70029 , n70030 , 
 n70031 , n70032 , n70033 , n70034 , n70035 , n70036 , n70037 , n70038 , n70039 , n70040 , 
 n70041 , n70042 , n70043 , n70044 , n70045 , n70046 , n70047 , n70048 , n70049 , n70050 , 
 n70051 , n70052 , n70053 , n70054 , n70055 , n70056 , n70057 , n70058 , n70059 , n70060 , 
 n70061 , n70062 , n70063 , n70064 , n70065 , n70066 , n70067 , n70068 , n70069 , n70070 , 
 n70071 , n70072 , n70073 , n70074 , n70075 , n70076 , n70077 , n70078 , n70079 , n70080 , 
 n70081 , n70082 , n70083 , n70084 , n70085 , n70086 , n70087 , n70088 , n70089 , n70090 , 
 n70091 , n70092 , n70093 , n70094 , n70095 , n70096 , n70097 , n70098 , n70099 , n70100 , 
 n70101 , n70102 , n70103 , n70104 , n70105 , n70106 , n70107 , n70108 , n70109 , n70110 , 
 n70111 , n70112 , n70113 , n70114 , n70115 , n70116 , n70117 , n70118 , n70119 , n70120 , 
 n70121 , n70122 , n70123 , n70124 , n70125 , n70126 , n70127 , n70128 , n70129 , n70130 , 
 n70131 , n70132 , n70133 , n70134 , n70135 , n70136 , n70137 , n70138 , n70139 , n70140 , 
 n70141 , n70142 , n70143 , n70144 , n70145 , n70146 , n70147 , n70148 , n70149 , n70150 , 
 n70151 , n70152 , n70153 , n70154 , n70155 , n70156 , n70157 , n70158 , n70159 , n70160 , 
 n70161 , n70162 , n70163 , n70164 , n70165 , n70166 , n70167 , n70168 , n70169 , n70170 , 
 n70171 , n70172 , n70173 , n70174 , n70175 , n70176 , n70177 , n70178 , n70179 , n70180 , 
 n70181 , n70182 , n70183 , n70184 , n70185 , n70186 , n70187 , n70188 , n70189 , n70190 , 
 n70191 , n70192 , n70193 , n70194 , n70195 , n70196 , n70197 , n70198 , n70199 , n70200 , 
 n70201 , n70202 , n70203 , n70204 , n70205 , n70206 , n70207 , n70208 , n70209 , n70210 , 
 n70211 , n70212 , n70213 , n70214 , n70215 , n70216 , n70217 , n70218 , n70219 , n70220 , 
 n70221 , n70222 , n70223 , n70224 , n70225 , n70226 , n70227 , n70228 , n70229 , n70230 , 
 n70231 , n70232 , n70233 , n70234 , n70235 , n70236 , n70237 , n70238 , n70239 , n70240 , 
 n70241 , n70242 , n70243 , n70244 , n70245 , n70246 , n70247 , n70248 , n70249 , n70250 , 
 n70251 , n70252 , n70253 , n70254 , n70255 , n70256 , n70257 , n70258 , n70259 , n70260 , 
 n70261 , n70262 , n70263 , n70264 , n70265 , n70266 , n70267 , n70268 , n70269 , n70270 , 
 n70271 , n70272 , n70273 , n70274 , n70275 , n70276 , n70277 , n70278 , n70279 , n70280 , 
 n70281 , n70282 , n70283 , n70284 , n70285 , n70286 , n70287 , n70288 , n70289 , n70290 , 
 n70291 , n70292 , n70293 , n70294 , n70295 , n70296 , n70297 , n70298 , n70299 , n70300 , 
 n70301 , n70302 , n70303 , n70304 , n70305 , n70306 , n70307 , n70308 , n70309 , n70310 , 
 n70311 , n70312 , n70313 , n70314 , n70315 , n70316 , n70317 , n70318 , n70319 , n70320 , 
 n70321 , n70322 , n70323 , n70324 , n70325 , n70326 , n70327 , n70328 , n70329 , n70330 , 
 n70331 , n70332 , n70333 , n70334 , n70335 , n70336 , n70337 , n70338 , n70339 , n70340 , 
 n70341 , n70342 , n70343 , n70344 , n70345 , n70346 , n70347 , n70348 , n70349 , n70350 , 
 n70351 , n70352 , n70353 , n70354 , n70355 , n70356 , n70357 , n70358 , n70359 , n70360 , 
 n70361 , n70362 , n70363 , n70364 , n70365 , n70366 , n70367 , n70368 , n70369 , n70370 , 
 n70371 , n70372 , n70373 , n70374 , n70375 , n70376 , n70377 , n70378 , n70379 , n70380 , 
 n70381 , n70382 , n70383 , n70384 , n70385 , n70386 , n70387 , n70388 , n70389 , n70390 , 
 n70391 , n70392 , n70393 , n70394 , n70395 , n70396 , n70397 , n70398 , n70399 , n70400 , 
 n70401 , n70402 , n70403 , n70404 , n70405 , n70406 , n70407 , n70408 , n70409 , n70410 , 
 n70411 , n70412 , n70413 , n70414 , n70415 , n70416 , n70417 , n70418 , n70419 , n70420 , 
 n70421 , n70422 , n70423 , n70424 , n70425 , n70426 , n70427 , n70428 , n70429 , n70430 , 
 n70431 , n70432 , n70433 , n70434 , n70435 , n70436 , n70437 , n70438 , n70439 , n70440 , 
 n70441 , n70442 , n70443 , n70444 , n70445 , n70446 , n70447 , n70448 , n70449 , n70450 , 
 n70451 , n70452 , n70453 , n70454 , n70455 , n70456 , n70457 , n70458 , n70459 , n70460 , 
 n70461 , n70462 , n70463 , n70464 , n70465 , n70466 , n70467 , n70468 , n70469 , n70470 , 
 n70471 , n70472 , n70473 , n70474 , n70475 , n70476 , n70477 , n70478 , n70479 , n70480 , 
 n70481 , n70482 , n70483 , n70484 , n70485 , n70486 , n70487 , n70488 , n70489 , n70490 , 
 n70491 , n70492 , n70493 , n70494 , n70495 , n70496 , n70497 , n70498 , n70499 , n70500 , 
 n70501 , n70502 , n70503 , n70504 , n70505 , n70506 , n70507 , n70508 , n70509 , n70510 , 
 n70511 , n70512 , n70513 , n70514 , n70515 , n70516 , n70517 , n70518 , n70519 , n70520 , 
 n70521 , n70522 , n70523 , n70524 , n70525 , n70526 , n70527 , n70528 , n70529 , n70530 , 
 n70531 , n70532 , n70533 , n70534 , n70535 , n70536 , n70537 , n70538 , n70539 , n70540 , 
 n70541 , n70542 , n70543 , n70544 , n70545 , n70546 , n70547 , n70548 , n70549 , n70550 , 
 n70551 , n70552 , n70553 , n70554 , n70555 , n70556 , n70557 , n70558 , n70559 , n70560 , 
 n70561 , n70562 , n70563 , n70564 , n70565 , n70566 , n70567 , n70568 , n70569 , n70570 , 
 n70571 , n70572 , n70573 , n70574 , n70575 , n70576 , n70577 , n70578 , n70579 , n70580 , 
 n70581 , n70582 , n70583 , n70584 , n70585 , n70586 , n70587 , n70588 , n70589 , n70590 , 
 n70591 , n70592 , n70593 , n70594 , n70595 , n70596 , n70597 , n70598 , n70599 , n70600 , 
 n70601 , n70602 , n70603 , n70604 , n70605 , n70606 , n70607 , n70608 , n70609 , n70610 , 
 n70611 , n70612 , n70613 , n70614 , n70615 , n70616 , n70617 , n70618 , n70619 , n70620 , 
 n70621 , n70622 , n70623 , n70624 , n70625 , n70626 , n70627 , n70628 , n70629 , n70630 , 
 n70631 , n70632 , n70633 , n70634 , n70635 , n70636 , n70637 , n70638 , n70639 , n70640 , 
 n70641 , n70642 , n70643 , n70644 , n70645 , n70646 , n70647 , n70648 , n70649 , n70650 , 
 n70651 , n70652 , n70653 , n70654 , n70655 , n70656 , n70657 , n70658 , n70659 , n70660 , 
 n70661 , n70662 , n70663 , n70664 , n70665 , n70666 , n70667 , n70668 , n70669 , n70670 , 
 n70671 , n70672 , n70673 , n70674 , n70675 , n70676 , n70677 , n70678 , n70679 , n70680 , 
 n70681 , n70682 , n70683 , n70684 , n70685 , n70686 , n70687 , n70688 , n70689 , n70690 , 
 n70691 , n70692 , n70693 , n70694 , n70695 , n70696 , n70697 , n70698 , n70699 , n70700 , 
 n70701 , n70702 , n70703 , n70704 , n70705 , n70706 , n70707 , n70708 , n70709 , n70710 , 
 n70711 , n70712 , n70713 , n70714 , n70715 , n70716 , n70717 , n70718 , n70719 , n70720 , 
 n70721 , n70722 , n70723 , n70724 , n70725 , n70726 , n70727 , n70728 , n70729 , n70730 , 
 n70731 , n70732 , n70733 , n70734 , n70735 , n70736 , n70737 , n70738 , n70739 , n70740 , 
 n70741 , n70742 , n70743 , n70744 , n70745 , n70746 , n70747 , n70748 , n70749 , n70750 , 
 n70751 , n70752 , n70753 , n70754 , n70755 , n70756 , n70757 , n70758 , n70759 , n70760 , 
 n70761 , n70762 , n70763 , n70764 , n70765 , n70766 , n70767 , n70768 , n70769 , n70770 , 
 n70771 , n70772 , n70773 , n70774 , n70775 , n70776 , n70777 , n70778 , n70779 , n70780 , 
 n70781 , n70782 , n70783 , n70784 , n70785 , n70786 , n70787 , n70788 , n70789 , n70790 , 
 n70791 , n70792 , n70793 , n70794 , n70795 , n70796 , n70797 , n70798 , n70799 , n70800 , 
 n70801 , n70802 , n70803 , n70804 , n70805 , n70806 , n70807 , n70808 , n70809 , n70810 , 
 n70811 , n70812 , n70813 , n70814 , n70815 , n70816 , n70817 , n70818 , n70819 , n70820 , 
 n70821 , n70822 , n70823 , n70824 , n70825 , n70826 , n70827 , n70828 , n70829 , n70830 , 
 n70831 , n70832 , n70833 , n70834 , n70835 , n70836 , n70837 , n70838 , n70839 , n70840 , 
 n70841 , n70842 , n70843 , n70844 , n70845 , n70846 , n70847 , n70848 , n70849 , n70850 , 
 n70851 , n70852 , n70853 , n70854 , n70855 , n70856 , n70857 , n70858 , n70859 , n70860 , 
 n70861 , n70862 , n70863 , n70864 , n70865 , n70866 , n70867 , n70868 , n70869 , n70870 , 
 n70871 , n70872 , n70873 , n70874 , n70875 , n70876 , n70877 , n70878 , n70879 , n70880 , 
 n70881 , n70882 , n70883 , n70884 , n70885 , n70886 , n70887 , n70888 , n70889 , n70890 , 
 n70891 , n70892 , n70893 , n70894 , n70895 , n70896 , n70897 , n70898 , n70899 , n70900 , 
 n70901 , n70902 , n70903 , n70904 , n70905 , n70906 , n70907 , n70908 , n70909 , n70910 , 
 n70911 , n70912 , n70913 , n70914 , n70915 , n70916 , n70917 , n70918 , n70919 , n70920 , 
 n70921 , n70922 , n70923 , n70924 , n70925 , n70926 , n70927 , n70928 , n70929 , n70930 , 
 n70931 , n70932 , n70933 , n70934 , n70935 , n70936 , n70937 , n70938 , n70939 , n70940 , 
 n70941 , n70942 , n70943 , n70944 , n70945 , n70946 , n70947 , n70948 , n70949 , n70950 , 
 n70951 , n70952 , n70953 , n70954 , n70955 , n70956 , n70957 , n70958 , n70959 , n70960 , 
 n70961 , n70962 , n70963 , n70964 , n70965 , n70966 , n70967 , n70968 , n70969 , n70970 , 
 n70971 , n70972 , n70973 , n70974 , n70975 , n70976 , n70977 , n70978 , n70979 , n70980 , 
 n70981 , n70982 , n70983 , n70984 , n70985 , n70986 , n70987 , n70988 , n70989 , n70990 , 
 n70991 , n70992 , n70993 , n70994 , n70995 , n70996 , n70997 , n70998 , n70999 , n71000 , 
 n71001 , n71002 , n71003 , n71004 , n71005 , n71006 , n71007 , n71008 , n71009 , n71010 , 
 n71011 , n71012 , n71013 , n71014 , n71015 , n71016 , n71017 , n71018 , n71019 , n71020 , 
 n71021 , n71022 , n71023 , n71024 , n71025 , n71026 , n71027 , n71028 , n71029 , n71030 , 
 n71031 , n71032 , n71033 , n71034 , n71035 , n71036 , n71037 , n71038 , n71039 , n71040 , 
 n71041 , n71042 , n71043 , n71044 , n71045 , n71046 , n71047 , n71048 , n71049 , n71050 , 
 n71051 , n71052 , n71053 , n71054 , n71055 , n71056 , n71057 , n71058 , n71059 , n71060 , 
 n71061 , n71062 , n71063 , n71064 , n71065 , n71066 , n71067 , n71068 , n71069 , n71070 , 
 n71071 , n71072 , n71073 , n71074 , n71075 , n71076 , n71077 , n71078 , n71079 , n71080 , 
 n71081 , n71082 , n71083 , n71084 , n71085 , n71086 , n71087 , n71088 , n71089 , n71090 , 
 n71091 , n71092 , n71093 , n71094 , n71095 , n71096 , n71097 , n71098 , n71099 , n71100 , 
 n71101 , n71102 , n71103 , n71104 , n71105 , n71106 , n71107 , n71108 , n71109 , n71110 , 
 n71111 , n71112 , n71113 , n71114 , n71115 , n71116 , n71117 , n71118 , n71119 , n71120 , 
 n71121 , n71122 , n71123 , n71124 , n71125 , n71126 , n71127 , n71128 , n71129 , n71130 , 
 n71131 , n71132 , n71133 , n71134 , n71135 , n71136 , n71137 , n71138 , n71139 , n71140 , 
 n71141 , n71142 , n71143 , n71144 , n71145 , n71146 , n71147 , n71148 , n71149 , n71150 , 
 n71151 , n71152 , n71153 , n71154 , n71155 , n71156 , n71157 , n71158 , n71159 , n71160 , 
 n71161 , n71162 , n71163 , n71164 , n71165 , n71166 , n71167 , n71168 , n71169 , n71170 , 
 n71171 , n71172 , n71173 , n71174 , n71175 , n71176 , n71177 , n71178 , n71179 , n71180 , 
 n71181 , n71182 , n71183 , n71184 , n71185 , n71186 , n71187 , n71188 , n71189 , n71190 , 
 n71191 , n71192 , n71193 , n71194 , n71195 , n71196 , n71197 , n71198 , n71199 , n71200 , 
 n71201 , n71202 , n71203 , n71204 , n71205 , n71206 , n71207 , n71208 , n71209 , n71210 , 
 n71211 , n71212 , n71213 , n71214 , n71215 , n71216 , n71217 , n71218 , n71219 , n71220 , 
 n71221 , n71222 , n71223 , n71224 , n71225 , n71226 , n71227 , n71228 , n71229 , n71230 , 
 n71231 , n71232 , n71233 , n71234 , n71235 , n71236 , n71237 , n71238 , n71239 , n71240 , 
 n71241 , n71242 , n71243 , n71244 , n71245 , n71246 , n71247 , n71248 , n71249 , n71250 , 
 n71251 , n71252 , n71253 , n71254 , n71255 , n71256 , n71257 , n71258 , n71259 , n71260 , 
 n71261 , n71262 , n71263 , n71264 , n71265 , n71266 , n71267 , n71268 , n71269 , n71270 , 
 n71271 , n71272 , n71273 , n71274 , n71275 , n71276 , n71277 , n71278 , n71279 , n71280 , 
 n71281 , n71282 , n71283 , n71284 , n71285 , n71286 , n71287 , n71288 , n71289 , n71290 , 
 n71291 , n71292 , n71293 , n71294 , n71295 , n71296 , n71297 , n71298 , n71299 , n71300 , 
 n71301 , n71302 , n71303 , n71304 , n71305 , n71306 , n71307 , n71308 , n71309 , n71310 , 
 n71311 , n71312 , n71313 , n71314 , n71315 , n71316 , n71317 , n71318 , n71319 , n71320 , 
 n71321 , n71322 , n71323 , n71324 , n71325 , n71326 , n71327 , n71328 , n71329 , n71330 , 
 n71331 , n71332 , n71333 , n71334 , n71335 , n71336 , n71337 , n71338 , n71339 , n71340 , 
 n71341 , n71342 , n71343 , n71344 , n71345 , n71346 , n71347 , n71348 , n71349 , n71350 , 
 n71351 , n71352 , n71353 , n71354 , n71355 , n71356 , n71357 , n71358 , n71359 , n71360 , 
 n71361 , n71362 , n71363 , n71364 , n71365 , n71366 , n71367 , n71368 , n71369 , n71370 , 
 n71371 , n71372 , n71373 , n71374 , n71375 , n71376 , n71377 , n71378 , n71379 , n71380 , 
 n71381 , n71382 , n71383 , n71384 , n71385 , n71386 , n71387 , n71388 , n71389 , n71390 , 
 n71391 , n71392 , n71393 , n71394 , n71395 , n71396 , n71397 , n71398 , n71399 , n71400 , 
 n71401 , n71402 , n71403 , n71404 , n71405 , n71406 , n71407 , n71408 , n71409 , n71410 , 
 n71411 , n71412 , n71413 , n71414 , n71415 , n71416 , n71417 , n71418 , n71419 , n71420 , 
 n71421 , n71422 , n71423 , n71424 , n71425 , n71426 , n71427 , n71428 , n71429 , n71430 , 
 n71431 , n71432 , n71433 , n71434 , n71435 , n71436 , n71437 , n71438 , n71439 , n71440 , 
 n71441 , n71442 , n71443 , n71444 , n71445 , n71446 , n71447 , n71448 , n71449 , n71450 , 
 n71451 , n71452 , n71453 , n71454 , n71455 , n71456 , n71457 , n71458 , n71459 , n71460 , 
 n71461 , n71462 , n71463 , n71464 , n71465 , n71466 , n71467 , n71468 , n71469 , n71470 , 
 n71471 , n71472 , n71473 , n71474 , n71475 , n71476 , n71477 , n71478 , n71479 , n71480 , 
 n71481 , n71482 , n71483 , n71484 , n71485 , n71486 , n71487 , n71488 , n71489 , n71490 , 
 n71491 , n71492 , n71493 , n71494 , n71495 , n71496 , n71497 , n71498 , n71499 , n71500 , 
 n71501 , n71502 , n71503 , n71504 , n71505 , n71506 , n71507 , n71508 , n71509 , n71510 , 
 n71511 , n71512 , n71513 , n71514 , n71515 , n71516 , n71517 , n71518 , n71519 , n71520 , 
 n71521 , n71522 , n71523 , n71524 , n71525 , n71526 , n71527 , n71528 , n71529 , n71530 , 
 n71531 , n71532 , n71533 , n71534 , n71535 , n71536 , n71537 , n71538 , n71539 , n71540 , 
 n71541 , n71542 , n71543 , n71544 , n71545 , n71546 , n71547 , n71548 , n71549 , n71550 , 
 n71551 , n71552 , n71553 , n71554 , n71555 , n71556 , n71557 , n71558 , n71559 , n71560 , 
 n71561 , n71562 , n71563 , n71564 , n71565 , n71566 , n71567 , n71568 , n71569 , n71570 , 
 n71571 , n71572 , n71573 , n71574 , n71575 , n71576 , n71577 , n71578 , n71579 , n71580 , 
 n71581 , n71582 , n71583 , n71584 , n71585 , n71586 , n71587 , n71588 , n71589 , n71590 , 
 n71591 , n71592 , n71593 , n71594 , n71595 , n71596 , n71597 , n71598 , n71599 , n71600 , 
 n71601 , n71602 , n71603 , n71604 , n71605 , n71606 , n71607 , n71608 , n71609 , n71610 , 
 n71611 , n71612 , n71613 , n71614 , n71615 , n71616 , n71617 , n71618 , n71619 , n71620 , 
 n71621 , n71622 , n71623 , n71624 , n71625 , n71626 , n71627 , n71628 , n71629 , n71630 , 
 n71631 , n71632 , n71633 , n71634 , n71635 , n71636 , n71637 , n71638 , n71639 , n71640 , 
 n71641 , n71642 , n71643 , n71644 , n71645 , n71646 , n71647 , n71648 , n71649 , n71650 , 
 n71651 , n71652 , n71653 , n71654 , n71655 , n71656 , n71657 , n71658 , n71659 , n71660 , 
 n71661 , n71662 , n71663 , n71664 , n71665 , n71666 , n71667 , n71668 , n71669 , n71670 , 
 n71671 , n71672 , n71673 , n71674 , n71675 , n71676 , n71677 , n71678 , n71679 , n71680 , 
 n71681 , n71682 , n71683 , n71684 , n71685 , n71686 , n71687 , n71688 , n71689 , n71690 , 
 n71691 , n71692 , n71693 , n71694 , n71695 , n71696 , n71697 , n71698 , n71699 , n71700 , 
 n71701 , n71702 , n71703 , n71704 , n71705 , n71706 , n71707 , n71708 , n71709 , n71710 , 
 n71711 , n71712 , n71713 , n71714 , n71715 , n71716 , n71717 , n71718 , n71719 , n71720 , 
 n71721 , n71722 , n71723 , n71724 , n71725 , n71726 , n71727 , n71728 , n71729 , n71730 , 
 n71731 , n71732 , n71733 , n71734 , n71735 , n71736 , n71737 , n71738 , n71739 , n71740 , 
 n71741 , n71742 , n71743 , n71744 , n71745 , n71746 , n71747 , n71748 , n71749 , n71750 , 
 n71751 , n71752 , n71753 , n71754 , n71755 , n71756 , n71757 , n71758 , n71759 , n71760 , 
 n71761 , n71762 , n71763 , n71764 , n71765 , n71766 , n71767 , n71768 , n71769 , n71770 , 
 n71771 , n71772 , n71773 , n71774 , n71775 , n71776 , n71777 , n71778 , n71779 , n71780 , 
 n71781 , n71782 , n71783 , n71784 , n71785 , n71786 , n71787 , n71788 , n71789 , n71790 , 
 n71791 , n71792 , n71793 , n71794 , n71795 , n71796 , n71797 , n71798 , n71799 , n71800 , 
 n71801 , n71802 , n71803 , n71804 , n71805 , n71806 , n71807 , n71808 , n71809 , n71810 , 
 n71811 , n71812 , n71813 , n71814 , n71815 , n71816 , n71817 , n71818 , n71819 , n71820 , 
 n71821 , n71822 , n71823 , n71824 , n71825 , n71826 , n71827 , n71828 , n71829 , n71830 , 
 n71831 , n71832 , n71833 , n71834 , n71835 , n71836 , n71837 , n71838 , n71839 , n71840 , 
 n71841 , n71842 , n71843 , n71844 , n71845 , n71846 , n71847 , n71848 , n71849 , n71850 , 
 n71851 , n71852 , n71853 , n71854 , n71855 , n71856 , n71857 , n71858 , n71859 , n71860 , 
 n71861 , n71862 , n71863 , n71864 , n71865 , n71866 , n71867 , n71868 , n71869 , n71870 , 
 n71871 , n71872 , n71873 , n71874 , n71875 , n71876 , n71877 , n71878 , n71879 , n71880 , 
 n71881 , n71882 , n71883 , n71884 , n71885 , n71886 , n71887 , n71888 , n71889 , n71890 , 
 n71891 , n71892 , n71893 , n71894 , n71895 , n71896 , n71897 , n71898 , n71899 , n71900 , 
 n71901 , n71902 , n71903 , n71904 , n71905 , n71906 , n71907 , n71908 , n71909 , n71910 , 
 n71911 , n71912 , n71913 , n71914 , n71915 , n71916 , n71917 , n71918 , n71919 , n71920 , 
 n71921 , n71922 , n71923 , n71924 , n71925 , n71926 , n71927 , n71928 , n71929 , n71930 , 
 n71931 , n71932 , n71933 , n71934 , n71935 , n71936 , n71937 , n71938 , n71939 , n71940 , 
 n71941 , n71942 , n71943 , n71944 , n71945 , n71946 , n71947 , n71948 , n71949 , n71950 , 
 n71951 , n71952 , n71953 , n71954 , n71955 , n71956 , n71957 , n71958 , n71959 , n71960 , 
 n71961 , n71962 , n71963 , n71964 , n71965 , n71966 , n71967 , n71968 , n71969 , n71970 , 
 n71971 , n71972 , n71973 , n71974 , n71975 , n71976 , n71977 , n71978 , n71979 , n71980 , 
 n71981 , n71982 , n71983 , n71984 , n71985 , n71986 , n71987 , n71988 , n71989 , n71990 , 
 n71991 , n71992 , n71993 , n71994 , n71995 , n71996 , n71997 , n71998 , n71999 , n72000 , 
 n72001 , n72002 , n72003 , n72004 , n72005 , n72006 , n72007 , n72008 , n72009 , n72010 , 
 n72011 , n72012 , n72013 , n72014 , n72015 , n72016 , n72017 , n72018 , n72019 , n72020 , 
 n72021 , n72022 , n72023 , n72024 , n72025 , n72026 , n72027 , n72028 , n72029 , n72030 , 
 n72031 , n72032 , n72033 , n72034 , n72035 , n72036 , n72037 , n72038 , n72039 , n72040 , 
 n72041 , n72042 , n72043 , n72044 , n72045 , n72046 , n72047 , n72048 , n72049 , n72050 , 
 n72051 , n72052 , n72053 , n72054 , n72055 , n72056 , n72057 , n72058 , n72059 , n72060 , 
 n72061 , n72062 , n72063 , n72064 , n72065 , n72066 , n72067 , n72068 , n72069 , n72070 , 
 n72071 , n72072 , n72073 , n72074 , n72075 , n72076 , n72077 , n72078 , n72079 , n72080 , 
 n72081 , n72082 , n72083 , n72084 , n72085 , n72086 , n72087 , n72088 , n72089 , n72090 , 
 n72091 , n72092 , n72093 , n72094 , n72095 , n72096 , n72097 , n72098 , n72099 , n72100 , 
 n72101 , n72102 , n72103 , n72104 , n72105 , n72106 , n72107 , n72108 , n72109 , n72110 , 
 n72111 , n72112 , n72113 , n72114 , n72115 , n72116 , n72117 , n72118 , n72119 , n72120 , 
 n72121 , n72122 , n72123 , n72124 , n72125 , n72126 , n72127 , n72128 , n72129 , n72130 , 
 n72131 , n72132 , n72133 , n72134 , n72135 , n72136 , n72137 , n72138 , n72139 , n72140 , 
 n72141 , n72142 , n72143 , n72144 , n72145 , n72146 , n72147 , n72148 , n72149 , n72150 , 
 n72151 , n72152 , n72153 , n72154 , n72155 , n72156 , n72157 , n72158 , n72159 , n72160 , 
 n72161 , n72162 , n72163 , n72164 , n72165 , n72166 , n72167 , n72168 , n72169 , n72170 , 
 n72171 , n72172 , n72173 , n72174 , n72175 , n72176 , n72177 , n72178 , n72179 , n72180 , 
 n72181 , n72182 , n72183 , n72184 , n72185 , n72186 , n72187 , n72188 , n72189 , n72190 , 
 n72191 , n72192 , n72193 , n72194 , n72195 , n72196 , n72197 , n72198 , n72199 , n72200 , 
 n72201 , n72202 , n72203 , n72204 , n72205 , n72206 , n72207 , n72208 , n72209 , n72210 , 
 n72211 , n72212 , n72213 , n72214 , n72215 , n72216 , n72217 , n72218 , n72219 , n72220 , 
 n72221 , n72222 , n72223 , n72224 , n72225 , n72226 , n72227 , n72228 , n72229 , n72230 , 
 n72231 , n72232 , n72233 , n72234 , n72235 , n72236 , n72237 , n72238 , n72239 , n72240 , 
 n72241 , n72242 , n72243 , n72244 , n72245 , n72246 , n72247 , n72248 , n72249 , n72250 , 
 n72251 , n72252 , n72253 , n72254 , n72255 , n72256 , n72257 , n72258 , n72259 , n72260 , 
 n72261 , n72262 , n72263 , n72264 , n72265 , n72266 , n72267 , n72268 , n72269 , n72270 , 
 n72271 , n72272 , n72273 , n72274 , n72275 , n72276 , n72277 , n72278 , n72279 , n72280 , 
 n72281 , n72282 , n72283 , n72284 , n72285 , n72286 , n72287 , n72288 , n72289 , n72290 , 
 n72291 , n72292 , n72293 , n72294 , n72295 , n72296 , n72297 , n72298 , n72299 , n72300 , 
 n72301 , n72302 , n72303 , n72304 , n72305 , n72306 , n72307 , n72308 , n72309 , n72310 , 
 n72311 , n72312 , n72313 , n72314 , n72315 , n72316 , n72317 , n72318 , n72319 , n72320 , 
 n72321 , n72322 , n72323 , n72324 , n72325 , n72326 , n72327 , n72328 , n72329 , n72330 , 
 n72331 , n72332 , n72333 , n72334 , n72335 , n72336 , n72337 , n72338 , n72339 , n72340 , 
 n72341 , n72342 , n72343 , n72344 , n72345 , n72346 , n72347 , n72348 , n72349 , n72350 , 
 n72351 , n72352 , n72353 , n72354 , n72355 , n72356 , n72357 , n72358 , n72359 , n72360 , 
 n72361 , n72362 , n72363 , n72364 , n72365 , n72366 , n72367 , n72368 , n72369 , n72370 , 
 n72371 , n72372 , n72373 , n72374 , n72375 , n72376 , n72377 , n72378 , n72379 , n72380 , 
 n72381 , n72382 , n72383 , n72384 , n72385 , n72386 , n72387 , n72388 , n72389 , n72390 , 
 n72391 , n72392 , n72393 , n72394 , n72395 , n72396 , n72397 , n72398 , n72399 , n72400 , 
 n72401 , n72402 , n72403 , n72404 , n72405 , n72406 , n72407 , n72408 , n72409 , n72410 , 
 n72411 , n72412 , n72413 , n72414 , n72415 , n72416 , n72417 , n72418 , n72419 , n72420 , 
 n72421 , n72422 , n72423 , n72424 , n72425 , n72426 , n72427 , n72428 , n72429 , n72430 , 
 n72431 , n72432 , n72433 , n72434 , n72435 , n72436 , n72437 , n72438 , n72439 , n72440 , 
 n72441 , n72442 , n72443 , n72444 , n72445 , n72446 , n72447 , n72448 , n72449 , n72450 , 
 n72451 , n72452 , n72453 , n72454 , n72455 , n72456 , n72457 , n72458 , n72459 , n72460 , 
 n72461 , n72462 , n72463 , n72464 , n72465 , n72466 , n72467 , n72468 , n72469 , n72470 , 
 n72471 , n72472 , n72473 , n72474 , n72475 , n72476 , n72477 , n72478 , n72479 , n72480 , 
 n72481 , n72482 , n72483 , n72484 , n72485 , n72486 , n72487 , n72488 , n72489 , n72490 , 
 n72491 , n72492 , n72493 , n72494 , n72495 , n72496 , n72497 , n72498 , n72499 , n72500 , 
 n72501 , n72502 , n72503 , n72504 , n72505 , n72506 , n72507 , n72508 , n72509 , n72510 , 
 n72511 , n72512 , n72513 , n72514 , n72515 , n72516 , n72517 , n72518 , n72519 , n72520 , 
 n72521 , n72522 , n72523 , n72524 , n72525 , n72526 , n72527 , n72528 , n72529 , n72530 , 
 n72531 , n72532 , n72533 , n72534 , n72535 , n72536 , n72537 , n72538 , n72539 , n72540 , 
 n72541 , n72542 , n72543 , n72544 , n72545 , n72546 , n72547 , n72548 , n72549 , n72550 , 
 n72551 , n72552 , n72553 , n72554 , n72555 , n72556 , n72557 , n72558 , n72559 , n72560 , 
 n72561 , n72562 , n72563 , n72564 , n72565 , n72566 , n72567 , n72568 , n72569 , n72570 , 
 n72571 , n72572 , n72573 , n72574 , n72575 , n72576 , n72577 , n72578 , n72579 , n72580 , 
 n72581 , n72582 , n72583 , n72584 , n72585 , n72586 , n72587 , n72588 , n72589 , n72590 , 
 n72591 , n72592 , n72593 , n72594 , n72595 , n72596 , n72597 , n72598 , n72599 , n72600 , 
 n72601 , n72602 , n72603 , n72604 , n72605 , n72606 , n72607 , n72608 , n72609 , n72610 , 
 n72611 , n72612 , n72613 , n72614 , n72615 , n72616 , n72617 , n72618 , n72619 , n72620 , 
 n72621 , n72622 , n72623 , n72624 , n72625 , n72626 , n72627 , n72628 , n72629 , n72630 , 
 n72631 , n72632 , n72633 , n72634 , n72635 , n72636 , n72637 , n72638 , n72639 , n72640 , 
 n72641 , n72642 , n72643 , n72644 , n72645 , n72646 , n72647 , n72648 , n72649 , n72650 , 
 n72651 , n72652 , n72653 , n72654 , n72655 , n72656 , n72657 , n72658 , n72659 , n72660 , 
 n72661 , n72662 , n72663 , n72664 , n72665 , n72666 , n72667 , n72668 , n72669 , n72670 , 
 n72671 , n72672 , n72673 , n72674 , n72675 , n72676 , n72677 , n72678 , n72679 , n72680 , 
 n72681 , n72682 , n72683 , n72684 , n72685 , n72686 , n72687 , n72688 , n72689 , n72690 , 
 n72691 , n72692 , n72693 , n72694 , n72695 , n72696 , n72697 , n72698 , n72699 , n72700 , 
 n72701 , n72702 , n72703 , n72704 , n72705 , n72706 , n72707 , n72708 , n72709 , n72710 , 
 n72711 , n72712 , n72713 , n72714 , n72715 , n72716 , n72717 , n72718 , n72719 , n72720 , 
 n72721 , n72722 , n72723 , n72724 , n72725 , n72726 , n72727 , n72728 , n72729 , n72730 , 
 n72731 , n72732 , n72733 , n72734 , n72735 , n72736 , n72737 , n72738 , n72739 , n72740 , 
 n72741 , n72742 , n72743 , n72744 , n72745 , n72746 , n72747 , n72748 , n72749 , n72750 , 
 n72751 , n72752 , n72753 , n72754 , n72755 , n72756 , n72757 , n72758 , n72759 , n72760 , 
 n72761 , n72762 , n72763 , n72764 , n72765 , n72766 , n72767 , n72768 , n72769 , n72770 , 
 n72771 , n72772 , n72773 , n72774 , n72775 , n72776 , n72777 , n72778 , n72779 , n72780 , 
 n72781 , n72782 , n72783 , n72784 , n72785 , n72786 , n72787 , n72788 , n72789 , n72790 , 
 n72791 , n72792 , n72793 , n72794 , n72795 , n72796 , n72797 , n72798 , n72799 , n72800 , 
 n72801 , n72802 , n72803 , n72804 , n72805 , n72806 , n72807 , n72808 , n72809 , n72810 , 
 n72811 , n72812 , n72813 , n72814 , n72815 , n72816 , n72817 , n72818 , n72819 , n72820 , 
 n72821 , n72822 , n72823 , n72824 , n72825 , n72826 , n72827 , n72828 , n72829 , n72830 , 
 n72831 , n72832 , n72833 , n72834 , n72835 , n72836 , n72837 , n72838 , n72839 , n72840 , 
 n72841 , n72842 , n72843 , n72844 , n72845 , n72846 , n72847 , n72848 , n72849 , n72850 , 
 n72851 , n72852 , n72853 , n72854 , n72855 , n72856 , n72857 , n72858 , n72859 , n72860 , 
 n72861 , n72862 , n72863 , n72864 , n72865 , n72866 , n72867 , n72868 , n72869 , n72870 , 
 n72871 , n72872 , n72873 , n72874 , n72875 , n72876 , n72877 , n72878 , n72879 , n72880 , 
 n72881 , n72882 , n72883 , n72884 , n72885 , n72886 , n72887 , n72888 , n72889 , n72890 , 
 n72891 , n72892 , n72893 , n72894 , n72895 , n72896 , n72897 , n72898 , n72899 , n72900 , 
 n72901 , n72902 , n72903 , n72904 , n72905 , n72906 , n72907 , n72908 , n72909 , n72910 , 
 n72911 , n72912 , n72913 , n72914 , n72915 , n72916 , n72917 , n72918 , n72919 , n72920 , 
 n72921 , n72922 , n72923 , n72924 , n72925 , n72926 , n72927 , n72928 , n72929 , n72930 , 
 n72931 , n72932 , n72933 , n72934 , n72935 , n72936 , n72937 , n72938 , n72939 , n72940 , 
 n72941 , n72942 , n72943 , n72944 , n72945 , n72946 , n72947 , n72948 , n72949 , n72950 , 
 n72951 , n72952 , n72953 , n72954 , n72955 , n72956 , n72957 , n72958 , n72959 , n72960 , 
 n72961 , n72962 , n72963 , n72964 , n72965 , n72966 , n72967 , n72968 , n72969 , n72970 , 
 n72971 , n72972 , n72973 , n72974 , n72975 , n72976 , n72977 , n72978 , n72979 , n72980 , 
 n72981 , n72982 , n72983 , n72984 , n72985 , n72986 , n72987 , n72988 , n72989 , n72990 , 
 n72991 , n72992 , n72993 , n72994 , n72995 , n72996 , n72997 , n72998 , n72999 , n73000 , 
 n73001 , n73002 , n73003 , n73004 , n73005 , n73006 , n73007 , n73008 , n73009 , n73010 , 
 n73011 , n73012 , n73013 , n73014 , n73015 , n73016 , n73017 , n73018 , n73019 , n73020 , 
 n73021 , n73022 , n73023 , n73024 , n73025 , n73026 , n73027 , n73028 , n73029 , n73030 , 
 n73031 , n73032 , n73033 , n73034 , n73035 , n73036 , n73037 , n73038 , n73039 , n73040 , 
 n73041 , n73042 , n73043 , n73044 , n73045 , n73046 , n73047 , n73048 , n73049 , n73050 , 
 n73051 , n73052 , n73053 , n73054 , n73055 , n73056 , n73057 , n73058 , n73059 , n73060 , 
 n73061 , n73062 , n73063 , n73064 , n73065 , n73066 , n73067 , n73068 , n73069 , n73070 , 
 n73071 , n73072 , n73073 , n73074 , n73075 , n73076 , n73077 , n73078 , n73079 , n73080 , 
 n73081 , n73082 , n73083 , n73084 , n73085 , n73086 , n73087 , n73088 , n73089 , n73090 , 
 n73091 , n73092 , n73093 , n73094 , n73095 , n73096 , n73097 , n73098 , n73099 , n73100 , 
 n73101 , n73102 , n73103 , n73104 , n73105 , n73106 , n73107 , n73108 , n73109 , n73110 , 
 n73111 , n73112 , n73113 , n73114 , n73115 , n73116 , n73117 , n73118 , n73119 , n73120 , 
 n73121 , n73122 , n73123 , n73124 , n73125 , n73126 , n73127 , n73128 , n73129 , n73130 , 
 n73131 , n73132 , n73133 , n73134 , n73135 , n73136 , n73137 , n73138 , n73139 , n73140 , 
 n73141 , n73142 , n73143 , n73144 , n73145 , n73146 , n73147 , n73148 , n73149 , n73150 , 
 n73151 , n73152 , n73153 , n73154 , n73155 , n73156 , n73157 , n73158 , n73159 , n73160 , 
 n73161 , n73162 , n73163 , n73164 , n73165 , n73166 , n73167 , n73168 , n73169 , n73170 , 
 n73171 , n73172 , n73173 , n73174 , n73175 , n73176 , n73177 , n73178 , n73179 , n73180 , 
 n73181 , n73182 , n73183 , n73184 , n73185 , n73186 , n73187 , n73188 , n73189 , n73190 , 
 n73191 , n73192 , n73193 , n73194 , n73195 , n73196 , n73197 , n73198 , n73199 , n73200 , 
 n73201 , n73202 , n73203 , n73204 , n73205 , n73206 , n73207 , n73208 , n73209 , n73210 , 
 n73211 , n73212 , n73213 , n73214 , n73215 , n73216 , n73217 , n73218 , n73219 , n73220 , 
 n73221 , n73222 , n73223 , n73224 , n73225 , n73226 , n73227 , n73228 , n73229 , n73230 , 
 n73231 , n73232 , n73233 , n73234 , n73235 , n73236 , n73237 , n73238 , n73239 , n73240 , 
 n73241 , n73242 , n73243 , n73244 , n73245 , n73246 , n73247 , n73248 , n73249 , n73250 , 
 n73251 , n73252 , n73253 , n73254 , n73255 , n73256 , n73257 , n73258 , n73259 , n73260 , 
 n73261 , n73262 , n73263 , n73264 , n73265 , n73266 , n73267 , n73268 , n73269 , n73270 , 
 n73271 , n73272 , n73273 , n73274 , n73275 , n73276 , n73277 , n73278 , n73279 , n73280 , 
 n73281 , n73282 , n73283 , n73284 , n73285 , n73286 , n73287 , n73288 , n73289 , n73290 , 
 n73291 , n73292 , n73293 , n73294 , n73295 , n73296 , n73297 , n73298 , n73299 , n73300 , 
 n73301 , n73302 , n73303 , n73304 , n73305 , n73306 , n73307 , n73308 , n73309 , n73310 , 
 n73311 , n73312 , n73313 , n73314 , n73315 , n73316 , n73317 , n73318 , n73319 , n73320 , 
 n73321 , n73322 , n73323 , n73324 , n73325 , n73326 , n73327 , n73328 , n73329 , n73330 , 
 n73331 , n73332 , n73333 , n73334 , n73335 , n73336 , n73337 , n73338 , n73339 , n73340 , 
 n73341 , n73342 , n73343 , n73344 , n73345 , n73346 , n73347 , n73348 , n73349 , n73350 , 
 n73351 , n73352 , n73353 , n73354 , n73355 , n73356 , n73357 , n73358 , n73359 , n73360 , 
 n73361 , n73362 , n73363 , n73364 , n73365 , n73366 , n73367 , n73368 , n73369 , n73370 , 
 n73371 , n73372 , n73373 , n73374 , n73375 , n73376 , n73377 , n73378 , n73379 , n73380 , 
 n73381 , n73382 , n73383 , n73384 , n73385 , n73386 , n73387 , n73388 , n73389 , n73390 , 
 n73391 , n73392 , n73393 , n73394 , n73395 , n73396 , n73397 , n73398 , n73399 , n73400 , 
 n73401 , n73402 , n73403 , n73404 , n73405 , n73406 , n73407 , n73408 , n73409 , n73410 , 
 n73411 , n73412 , n73413 , n73414 , n73415 , n73416 , n73417 , n73418 , n73419 , n73420 , 
 n73421 , n73422 , n73423 , n73424 , n73425 , n73426 , n73427 , n73428 , n73429 , n73430 , 
 n73431 , n73432 , n73433 , n73434 , n73435 , n73436 , n73437 , n73438 , n73439 , n73440 , 
 n73441 , n73442 , n73443 , n73444 , n73445 , n73446 , n73447 , n73448 , n73449 , n73450 , 
 n73451 , n73452 , n73453 , n73454 , n73455 , n73456 , n73457 , n73458 , n73459 , n73460 , 
 n73461 , n73462 , n73463 , n73464 , n73465 , n73466 , n73467 , n73468 , n73469 , n73470 , 
 n73471 , n73472 , n73473 , n73474 , n73475 , n73476 , n73477 , n73478 , n73479 , n73480 , 
 n73481 , n73482 , n73483 , n73484 , n73485 , n73486 , n73487 , n73488 , n73489 , n73490 , 
 n73491 , n73492 , n73493 , n73494 , n73495 , n73496 , n73497 , n73498 , n73499 , n73500 , 
 n73501 , n73502 , n73503 , n73504 , n73505 , n73506 , n73507 , n73508 , n73509 , n73510 , 
 n73511 , n73512 , n73513 , n73514 , n73515 , n73516 , n73517 , n73518 , n73519 , n73520 , 
 n73521 , n73522 , n73523 , n73524 , n73525 , n73526 , n73527 , n73528 , n73529 , n73530 , 
 n73531 , n73532 , n73533 , n73534 , n73535 , n73536 , n73537 , n73538 , n73539 , n73540 , 
 n73541 , n73542 , n73543 , n73544 , n73545 , n73546 , n73547 , n73548 , n73549 , n73550 , 
 n73551 , n73552 , n73553 , n73554 , n73555 , n73556 , n73557 , n73558 , n73559 , n73560 , 
 n73561 , n73562 , n73563 , n73564 , n73565 , n73566 , n73567 , n73568 , n73569 , n73570 , 
 n73571 , n73572 , n73573 , n73574 , n73575 , n73576 , n73577 , n73578 , n73579 , n73580 , 
 n73581 , n73582 , n73583 , n73584 , n73585 , n73586 , n73587 , n73588 , n73589 , n73590 , 
 n73591 , n73592 , n73593 , n73594 , n73595 , n73596 , n73597 , n73598 , n73599 , n73600 , 
 n73601 , n73602 , n73603 , n73604 , n73605 , n73606 , n73607 , n73608 , n73609 , n73610 , 
 n73611 , n73612 , n73613 , n73614 , n73615 , n73616 , n73617 , n73618 , n73619 , n73620 , 
 n73621 , n73622 , n73623 , n73624 , n73625 , n73626 , n73627 , n73628 , n73629 , n73630 , 
 n73631 , n73632 , n73633 , n73634 , n73635 , n73636 , n73637 , n73638 , n73639 , n73640 , 
 n73641 , n73642 , n73643 , n73644 , n73645 , n73646 , n73647 , n73648 , n73649 , n73650 , 
 n73651 , n73652 , n73653 , n73654 , n73655 , n73656 , n73657 , n73658 , n73659 , n73660 , 
 n73661 , n73662 , n73663 , n73664 , n73665 , n73666 , n73667 , n73668 , n73669 , n73670 , 
 n73671 , n73672 , n73673 , n73674 , n73675 , n73676 , n73677 , n73678 , n73679 , n73680 , 
 n73681 , n73682 , n73683 , n73684 , n73685 , n73686 , n73687 , n73688 , n73689 , n73690 , 
 n73691 , n73692 , n73693 , n73694 , n73695 , n73696 , n73697 , n73698 , n73699 , n73700 , 
 n73701 , n73702 , n73703 , n73704 , n73705 , n73706 , n73707 , n73708 , n73709 , n73710 , 
 n73711 , n73712 , n73713 , n73714 , n73715 , n73716 , n73717 , n73718 , n73719 , n73720 , 
 n73721 , n73722 , n73723 , n73724 , n73725 , n73726 , n73727 , n73728 , n73729 , n73730 , 
 n73731 , n73732 , n73733 , n73734 , n73735 , n73736 , n73737 , n73738 , n73739 , n73740 , 
 n73741 , n73742 , n73743 , n73744 , n73745 , n73746 , n73747 , n73748 , n73749 , n73750 , 
 n73751 , n73752 , n73753 , n73754 , n73755 , n73756 , n73757 , n73758 , n73759 , n73760 , 
 n73761 , n73762 , n73763 , n73764 , n73765 , n73766 , n73767 , n73768 , n73769 , n73770 , 
 n73771 , n73772 , n73773 , n73774 , n73775 , n73776 , n73777 , n73778 , n73779 , n73780 , 
 n73781 , n73782 , n73783 , n73784 , n73785 , n73786 , n73787 , n73788 , n73789 , n73790 , 
 n73791 , n73792 , n73793 , n73794 , n73795 , n73796 , n73797 , n73798 , n73799 , n73800 , 
 n73801 , n73802 , n73803 , n73804 , n73805 , n73806 , n73807 , n73808 , n73809 , n73810 , 
 n73811 , n73812 , n73813 , n73814 , n73815 , n73816 , n73817 , n73818 , n73819 , n73820 , 
 n73821 , n73822 , n73823 , n73824 , n73825 , n73826 , n73827 , n73828 , n73829 , n73830 , 
 n73831 , n73832 , n73833 , n73834 , n73835 , n73836 , n73837 , n73838 , n73839 , n73840 , 
 n73841 , n73842 , n73843 , n73844 , n73845 , n73846 , n73847 , n73848 , n73849 , n73850 , 
 n73851 , n73852 , n73853 , n73854 , n73855 , n73856 , n73857 , n73858 , n73859 , n73860 , 
 n73861 , n73862 , n73863 , n73864 , n73865 , n73866 , n73867 , n73868 , n73869 , n73870 , 
 n73871 , n73872 , n73873 , n73874 , n73875 , n73876 , n73877 , n73878 , n73879 , n73880 , 
 n73881 , n73882 , n73883 , n73884 , n73885 , n73886 , n73887 , n73888 , n73889 , n73890 , 
 n73891 , n73892 , n73893 , n73894 , n73895 , n73896 , n73897 , n73898 , n73899 , n73900 , 
 n73901 , n73902 , n73903 , n73904 , n73905 , n73906 , n73907 , n73908 , n73909 , n73910 , 
 n73911 , n73912 , n73913 , n73914 , n73915 , n73916 , n73917 , n73918 , n73919 , n73920 , 
 n73921 , n73922 , n73923 , n73924 , n73925 , n73926 , n73927 , n73928 , n73929 , n73930 , 
 n73931 , n73932 , n73933 , n73934 , n73935 , n73936 , n73937 , n73938 , n73939 , n73940 , 
 n73941 , n73942 , n73943 , n73944 , n73945 , n73946 , n73947 , n73948 , n73949 , n73950 , 
 n73951 , n73952 , n73953 , n73954 , n73955 , n73956 , n73957 , n73958 , n73959 , n73960 , 
 n73961 , n73962 , n73963 , n73964 , n73965 , n73966 , n73967 , n73968 , n73969 , n73970 , 
 n73971 , n73972 , n73973 , n73974 , n73975 , n73976 , n73977 , n73978 , n73979 , n73980 , 
 n73981 , n73982 , n73983 , n73984 , n73985 , n73986 , n73987 , n73988 , n73989 , n73990 , 
 n73991 , n73992 , n73993 , n73994 , n73995 , n73996 , n73997 , n73998 , n73999 , n74000 , 
 n74001 , n74002 , n74003 , n74004 , n74005 , n74006 , n74007 , n74008 , n74009 , n74010 , 
 n74011 , n74012 , n74013 , n74014 , n74015 , n74016 , n74017 , n74018 , n74019 , n74020 , 
 n74021 , n74022 , n74023 , n74024 , n74025 , n74026 , n74027 , n74028 , n74029 , n74030 , 
 n74031 , n74032 , n74033 , n74034 , n74035 , n74036 , n74037 , n74038 , n74039 , n74040 , 
 n74041 , n74042 , n74043 , n74044 , n74045 , n74046 , n74047 , n74048 , n74049 , n74050 , 
 n74051 , n74052 , n74053 , n74054 , n74055 , n74056 , n74057 , n74058 , n74059 , n74060 , 
 n74061 , n74062 , n74063 , n74064 , n74065 , n74066 , n74067 , n74068 , n74069 , n74070 , 
 n74071 , n74072 , n74073 , n74074 , n74075 , n74076 , n74077 , n74078 , n74079 , n74080 , 
 n74081 , n74082 , n74083 , n74084 , n74085 , n74086 , n74087 , n74088 , n74089 , n74090 , 
 n74091 , n74092 , n74093 , n74094 , n74095 , n74096 , n74097 , n74098 , n74099 , n74100 , 
 n74101 , n74102 , n74103 , n74104 , n74105 , n74106 , n74107 , n74108 , n74109 , n74110 , 
 n74111 , n74112 , n74113 , n74114 , n74115 , n74116 , n74117 , n74118 , n74119 , n74120 , 
 n74121 , n74122 , n74123 , n74124 , n74125 , n74126 , n74127 , n74128 , n74129 , n74130 , 
 n74131 , n74132 , n74133 , n74134 , n74135 , n74136 , n74137 , n74138 , n74139 , n74140 , 
 n74141 , n74142 , n74143 , n74144 , n74145 , n74146 , n74147 , n74148 , n74149 , n74150 , 
 n74151 , n74152 , n74153 , n74154 , n74155 , n74156 , n74157 , n74158 , n74159 , n74160 , 
 n74161 , n74162 , n74163 , n74164 , n74165 , n74166 , n74167 , n74168 , n74169 , n74170 , 
 n74171 , n74172 , n74173 , n74174 , n74175 , n74176 , n74177 , n74178 , n74179 , n74180 , 
 n74181 , n74182 , n74183 , n74184 , n74185 , n74186 , n74187 , n74188 , n74189 , n74190 , 
 n74191 , n74192 , n74193 , n74194 , n74195 , n74196 , n74197 , n74198 , n74199 , n74200 , 
 n74201 , n74202 , n74203 , n74204 , n74205 , n74206 , n74207 , n74208 , n74209 , n74210 , 
 n74211 , n74212 , n74213 , n74214 , n74215 , n74216 , n74217 , n74218 , n74219 , n74220 , 
 n74221 , n74222 , n74223 , n74224 , n74225 , n74226 , n74227 , n74228 , n74229 , n74230 , 
 n74231 , n74232 , n74233 , n74234 , n74235 , n74236 , n74237 , n74238 , n74239 , n74240 , 
 n74241 , n74242 , n74243 , n74244 , n74245 , n74246 , n74247 , n74248 , n74249 , n74250 , 
 n74251 , n74252 , n74253 , n74254 , n74255 , n74256 , n74257 , n74258 , n74259 , n74260 , 
 n74261 , n74262 , n74263 , n74264 , n74265 , n74266 , n74267 , n74268 , n74269 , n74270 , 
 n74271 , n74272 , n74273 , n74274 , n74275 , n74276 , n74277 , n74278 , n74279 , n74280 , 
 n74281 , n74282 , n74283 , n74284 , n74285 , n74286 , n74287 , n74288 , n74289 , n74290 , 
 n74291 , n74292 , n74293 , n74294 , n74295 , n74296 , n74297 , n74298 , n74299 , n74300 , 
 n74301 , n74302 , n74303 , n74304 , n74305 , n74306 , n74307 , n74308 , n74309 , n74310 , 
 n74311 , n74312 , n74313 , n74314 , n74315 , n74316 , n74317 , n74318 , n74319 , n74320 , 
 n74321 , n74322 , n74323 , n74324 , n74325 , n74326 , n74327 , n74328 , n74329 , n74330 , 
 n74331 , n74332 , n74333 , n74334 , n74335 , n74336 , n74337 , n74338 , n74339 , n74340 , 
 n74341 , n74342 , n74343 , n74344 , n74345 , n74346 , n74347 , n74348 , n74349 , n74350 , 
 n74351 , n74352 , n74353 , n74354 , n74355 , n74356 , n74357 , n74358 , n74359 , n74360 , 
 n74361 , n74362 , n74363 , n74364 , n74365 , n74366 , n74367 , n74368 , n74369 , n74370 , 
 n74371 , n74372 , n74373 , n74374 , n74375 , n74376 , n74377 , n74378 , n74379 , n74380 , 
 n74381 , n74382 , n74383 , n74384 , n74385 , n74386 , n74387 , n74388 , n74389 , n74390 , 
 n74391 , n74392 , n74393 , n74394 , n74395 , n74396 , n74397 , n74398 , n74399 , n74400 , 
 n74401 , n74402 , n74403 , n74404 , n74405 , n74406 , n74407 , n74408 , n74409 , n74410 , 
 n74411 , n74412 , n74413 , n74414 , n74415 , n74416 , n74417 , n74418 , n74419 , n74420 , 
 n74421 , n74422 , n74423 , n74424 , n74425 , n74426 , n74427 , n74428 , n74429 , n74430 , 
 n74431 , n74432 , n74433 , n74434 , n74435 , n74436 , n74437 , n74438 , n74439 , n74440 , 
 n74441 , n74442 , n74443 , n74444 , n74445 , n74446 , n74447 , n74448 , n74449 , n74450 , 
 n74451 , n74452 , n74453 , n74454 , n74455 , n74456 , n74457 , n74458 , n74459 , n74460 , 
 n74461 , n74462 , n74463 , n74464 , n74465 , n74466 , n74467 , n74468 , n74469 , n74470 , 
 n74471 , n74472 , n74473 , n74474 , n74475 , n74476 , n74477 , n74478 , n74479 , n74480 , 
 n74481 , n74482 , n74483 , n74484 , n74485 , n74486 , n74487 , n74488 , n74489 , n74490 , 
 n74491 , n74492 , n74493 , n74494 , n74495 , n74496 , n74497 , n74498 , n74499 , n74500 , 
 n74501 , n74502 , n74503 , n74504 , n74505 , n74506 , n74507 , n74508 , n74509 , n74510 , 
 n74511 , n74512 , n74513 , n74514 , n74515 , n74516 , n74517 , n74518 , n74519 , n74520 , 
 n74521 , n74522 , n74523 , n74524 , n74525 , n74526 , n74527 , n74528 , n74529 , n74530 , 
 n74531 , n74532 , n74533 , n74534 , n74535 , n74536 , n74537 , n74538 , n74539 , n74540 , 
 n74541 , n74542 , n74543 , n74544 , n74545 , n74546 , n74547 , n74548 , n74549 , n74550 , 
 n74551 , n74552 , n74553 , n74554 , n74555 , n74556 , n74557 , n74558 , n74559 , n74560 , 
 n74561 , n74562 , n74563 , n74564 , n74565 , n74566 , n74567 , n74568 , n74569 , n74570 , 
 n74571 , n74572 , n74573 , n74574 , n74575 , n74576 , n74577 , n74578 , n74579 , n74580 , 
 n74581 , n74582 , n74583 , n74584 , n74585 , n74586 , n74587 , n74588 , n74589 , n74590 , 
 n74591 , n74592 , n74593 , n74594 , n74595 , n74596 , n74597 , n74598 , n74599 , n74600 , 
 n74601 , n74602 , n74603 , n74604 , n74605 , n74606 , n74607 , n74608 , n74609 , n74610 , 
 n74611 , n74612 , n74613 , n74614 , n74615 , n74616 , n74617 , n74618 , n74619 , n74620 , 
 n74621 , n74622 , n74623 , n74624 , n74625 , n74626 , n74627 , n74628 , n74629 , n74630 , 
 n74631 , n74632 , n74633 , n74634 , n74635 , n74636 , n74637 , n74638 , n74639 , n74640 , 
 n74641 , n74642 , n74643 , n74644 , n74645 , n74646 , n74647 , n74648 , n74649 , n74650 , 
 n74651 , n74652 , n74653 , n74654 , n74655 , n74656 , n74657 , n74658 , n74659 , n74660 , 
 n74661 , n74662 , n74663 , n74664 , n74665 , n74666 , n74667 , n74668 , n74669 , n74670 , 
 n74671 , n74672 , n74673 , n74674 , n74675 , n74676 , n74677 , n74678 , n74679 , n74680 , 
 n74681 , n74682 , n74683 , n74684 , n74685 , n74686 , n74687 , n74688 , n74689 , n74690 , 
 n74691 , n74692 , n74693 , n74694 , n74695 , n74696 , n74697 , n74698 , n74699 , n74700 , 
 n74701 , n74702 , n74703 , n74704 , n74705 , n74706 , n74707 , n74708 , n74709 , n74710 , 
 n74711 , n74712 , n74713 , n74714 , n74715 , n74716 , n74717 , n74718 , n74719 , n74720 , 
 n74721 , n74722 , n74723 , n74724 , n74725 , n74726 , n74727 , n74728 , n74729 , n74730 , 
 n74731 , n74732 , n74733 , n74734 , n74735 , n74736 , n74737 , n74738 , n74739 , n74740 , 
 n74741 , n74742 , n74743 , n74744 , n74745 , n74746 , n74747 , n74748 , n74749 , n74750 , 
 n74751 , n74752 , n74753 , n74754 , n74755 , n74756 , n74757 , n74758 , n74759 , n74760 , 
 n74761 , n74762 , n74763 , n74764 , n74765 , n74766 , n74767 , n74768 , n74769 , n74770 , 
 n74771 , n74772 , n74773 , n74774 , n74775 , n74776 , n74777 , n74778 , n74779 , n74780 , 
 n74781 , n74782 , n74783 , n74784 , n74785 , n74786 , n74787 , n74788 , n74789 , n74790 , 
 n74791 , n74792 , n74793 , n74794 , n74795 , n74796 , n74797 , n74798 , n74799 , n74800 , 
 n74801 , n74802 , n74803 , n74804 , n74805 , n74806 , n74807 , n74808 , n74809 , n74810 , 
 n74811 , n74812 , n74813 , n74814 , n74815 , n74816 , n74817 , n74818 , n74819 , n74820 , 
 n74821 , n74822 , n74823 , n74824 , n74825 , n74826 , n74827 , n74828 , n74829 , n74830 , 
 n74831 , n74832 , n74833 , n74834 , n74835 , n74836 , n74837 , n74838 , n74839 , n74840 , 
 n74841 , n74842 , n74843 , n74844 , n74845 , n74846 , n74847 , n74848 , n74849 , n74850 , 
 n74851 , n74852 , n74853 , n74854 , n74855 , n74856 , n74857 , n74858 , n74859 , n74860 , 
 n74861 , n74862 , n74863 , n74864 , n74865 , n74866 , n74867 , n74868 , n74869 , n74870 , 
 n74871 , n74872 , n74873 , n74874 , n74875 , n74876 , n74877 , n74878 , n74879 , n74880 , 
 n74881 , n74882 , n74883 , n74884 , n74885 , n74886 , n74887 , n74888 , n74889 , n74890 , 
 n74891 , n74892 , n74893 , n74894 , n74895 , n74896 , n74897 , n74898 , n74899 , n74900 , 
 n74901 , n74902 , n74903 , n74904 , n74905 , n74906 , n74907 , n74908 , n74909 , n74910 , 
 n74911 , n74912 , n74913 , n74914 , n74915 , n74916 , n74917 , n74918 , n74919 , n74920 , 
 n74921 , n74922 , n74923 , n74924 , n74925 , n74926 , n74927 , n74928 , n74929 , n74930 , 
 n74931 , n74932 , n74933 , n74934 , n74935 , n74936 , n74937 , n74938 , n74939 , n74940 , 
 n74941 , n74942 , n74943 , n74944 , n74945 , n74946 , n74947 , n74948 , n74949 , n74950 , 
 n74951 , n74952 , n74953 , n74954 , n74955 , n74956 , n74957 , n74958 , n74959 , n74960 , 
 n74961 , n74962 , n74963 , n74964 , n74965 , n74966 , n74967 , n74968 , n74969 , n74970 , 
 n74971 , n74972 , n74973 , n74974 , n74975 , n74976 , n74977 , n74978 , n74979 , n74980 , 
 n74981 , n74982 , n74983 , n74984 , n74985 , n74986 , n74987 , n74988 , n74989 , n74990 , 
 n74991 , n74992 , n74993 , n74994 , n74995 , n74996 , n74997 , n74998 , n74999 , n75000 , 
 n75001 , n75002 , n75003 , n75004 , n75005 , n75006 , n75007 , n75008 , n75009 , n75010 , 
 n75011 , n75012 , n75013 , n75014 , n75015 , n75016 , n75017 , n75018 , n75019 , n75020 , 
 n75021 , n75022 , n75023 , n75024 , n75025 , n75026 , n75027 , n75028 , n75029 , n75030 , 
 n75031 , n75032 , n75033 , n75034 , n75035 , n75036 , n75037 , n75038 , n75039 , n75040 , 
 n75041 , n75042 , n75043 , n75044 , n75045 , n75046 , n75047 , n75048 , n75049 , n75050 , 
 n75051 , n75052 , n75053 , n75054 , n75055 , n75056 , n75057 , n75058 , n75059 , n75060 , 
 n75061 , n75062 , n75063 , n75064 , n75065 , n75066 , n75067 , n75068 , n75069 , n75070 , 
 n75071 , n75072 , n75073 , n75074 , n75075 , n75076 , n75077 , n75078 , n75079 , n75080 , 
 n75081 , n75082 , n75083 , n75084 , n75085 , n75086 , n75087 , n75088 , n75089 , n75090 , 
 n75091 , n75092 , n75093 , n75094 , n75095 , n75096 , n75097 , n75098 , n75099 , n75100 , 
 n75101 , n75102 , n75103 , n75104 , n75105 , n75106 , n75107 , n75108 , n75109 , n75110 , 
 n75111 , n75112 , n75113 , n75114 , n75115 , n75116 , n75117 , n75118 , n75119 , n75120 , 
 n75121 , n75122 , n75123 , n75124 , n75125 , n75126 , n75127 , n75128 , n75129 , n75130 , 
 n75131 , n75132 , n75133 , n75134 , n75135 , n75136 , n75137 , n75138 , n75139 , n75140 , 
 n75141 , n75142 , n75143 , n75144 , n75145 , n75146 , n75147 , n75148 , n75149 , n75150 , 
 n75151 , n75152 , n75153 , n75154 , n75155 , n75156 , n75157 , n75158 , n75159 , n75160 , 
 n75161 , n75162 , n75163 , n75164 , n75165 , n75166 , n75167 , n75168 , n75169 , n75170 , 
 n75171 , n75172 , n75173 , n75174 , n75175 , n75176 , n75177 , n75178 , n75179 , n75180 , 
 n75181 , n75182 , n75183 , n75184 , n75185 , n75186 , n75187 , n75188 , n75189 , n75190 , 
 n75191 , n75192 , n75193 , n75194 , n75195 , n75196 , n75197 , n75198 , n75199 , n75200 , 
 n75201 , n75202 , n75203 , n75204 , n75205 , n75206 , n75207 , n75208 , n75209 , n75210 , 
 n75211 , n75212 , n75213 , n75214 , n75215 , n75216 , n75217 , n75218 , n75219 , n75220 , 
 n75221 , n75222 , n75223 , n75224 , n75225 , n75226 , n75227 , n75228 , n75229 , n75230 , 
 n75231 , n75232 , n75233 , n75234 , n75235 , n75236 , n75237 , n75238 , n75239 , n75240 , 
 n75241 , n75242 , n75243 , n75244 , n75245 , n75246 , n75247 , n75248 , n75249 , n75250 , 
 n75251 , n75252 , n75253 , n75254 , n75255 , n75256 , n75257 , n75258 , n75259 , n75260 , 
 n75261 , n75262 , n75263 , n75264 , n75265 , n75266 , n75267 , n75268 , n75269 , n75270 , 
 n75271 , n75272 , n75273 , n75274 , n75275 , n75276 , n75277 , n75278 , n75279 , n75280 , 
 n75281 , n75282 , n75283 , n75284 , n75285 , n75286 , n75287 , n75288 , n75289 , n75290 , 
 n75291 , n75292 , n75293 , n75294 , n75295 , n75296 , n75297 , n75298 , n75299 , n75300 , 
 n75301 , n75302 , n75303 , n75304 , n75305 , n75306 , n75307 , n75308 , n75309 , n75310 , 
 n75311 , n75312 , n75313 , n75314 , n75315 , n75316 , n75317 , n75318 , n75319 , n75320 , 
 n75321 , n75322 , n75323 , n75324 , n75325 , n75326 , n75327 , n75328 , n75329 , n75330 , 
 n75331 , n75332 , n75333 , n75334 , n75335 , n75336 , n75337 , n75338 , n75339 , n75340 , 
 n75341 , n75342 , n75343 , n75344 , n75345 , n75346 , n75347 , n75348 , n75349 , n75350 , 
 n75351 , n75352 , n75353 , n75354 , n75355 , n75356 , n75357 , n75358 , n75359 , n75360 , 
 n75361 , n75362 , n75363 , n75364 , n75365 , n75366 , n75367 , n75368 , n75369 , n75370 , 
 n75371 , n75372 , n75373 , n75374 , n75375 , n75376 , n75377 , n75378 , n75379 , n75380 , 
 n75381 , n75382 , n75383 , n75384 , n75385 , n75386 , n75387 , n75388 , n75389 , n75390 , 
 n75391 , n75392 , n75393 , n75394 , n75395 , n75396 , n75397 , n75398 , n75399 , n75400 , 
 n75401 , n75402 , n75403 , n75404 , n75405 , n75406 , n75407 , n75408 , n75409 , n75410 , 
 n75411 , n75412 , n75413 , n75414 , n75415 , n75416 , n75417 , n75418 , n75419 , n75420 , 
 n75421 , n75422 , n75423 , n75424 , n75425 , n75426 , n75427 , n75428 , n75429 , n75430 , 
 n75431 , n75432 , n75433 , n75434 , n75435 , n75436 , n75437 , n75438 , n75439 , n75440 , 
 n75441 , n75442 , n75443 , n75444 , n75445 , n75446 , n75447 , n75448 , n75449 , n75450 , 
 n75451 , n75452 , n75453 , n75454 , n75455 , n75456 , n75457 , n75458 , n75459 , n75460 , 
 n75461 , n75462 , n75463 , n75464 , n75465 , n75466 , n75467 , n75468 , n75469 , n75470 , 
 n75471 , n75472 , n75473 , n75474 , n75475 , n75476 , n75477 , n75478 , n75479 , n75480 , 
 n75481 , n75482 , n75483 , n75484 , n75485 , n75486 , n75487 , n75488 , n75489 , n75490 , 
 n75491 , n75492 , n75493 , n75494 , n75495 , n75496 , n75497 , n75498 , n75499 , n75500 , 
 n75501 , n75502 , n75503 , n75504 , n75505 , n75506 , n75507 , n75508 , n75509 , n75510 , 
 n75511 , n75512 , n75513 , n75514 , n75515 , n75516 , n75517 , n75518 , n75519 , n75520 , 
 n75521 , n75522 , n75523 , n75524 , n75525 , n75526 , n75527 , n75528 , n75529 , n75530 , 
 n75531 , n75532 , n75533 , n75534 , n75535 , n75536 , n75537 , n75538 , n75539 , n75540 , 
 n75541 , n75542 , n75543 , n75544 , n75545 , n75546 , n75547 , n75548 , n75549 , n75550 , 
 n75551 , n75552 , n75553 , n75554 , n75555 , n75556 , n75557 , n75558 , n75559 , n75560 , 
 n75561 , n75562 , n75563 , n75564 , n75565 , n75566 , n75567 , n75568 , n75569 , n75570 , 
 n75571 , n75572 , n75573 , n75574 , n75575 , n75576 , n75577 , n75578 , n75579 , n75580 , 
 n75581 , n75582 , n75583 , n75584 , n75585 , n75586 , n75587 , n75588 , n75589 , n75590 , 
 n75591 , C0n , C0 ;
buf ( n1090 , n0 );
buf ( n1091 , n1 );
buf ( n1092 , n2 );
buf ( n1093 , n3 );
buf ( n1094 , n4 );
buf ( n1095 , n5 );
buf ( n1096 , n6 );
buf ( n1097 , n7 );
buf ( n1098 , n8 );
buf ( n1099 , n9 );
buf ( n1100 , n10 );
buf ( n1101 , n11 );
buf ( n1102 , n12 );
buf ( n1103 , n13 );
buf ( n1104 , n14 );
buf ( n1105 , n15 );
buf ( n1106 , n16 );
buf ( n1107 , n17 );
buf ( n1108 , n18 );
buf ( n1109 , n19 );
buf ( n1110 , n20 );
buf ( n1111 , n21 );
buf ( n1112 , n22 );
buf ( n1113 , n23 );
buf ( n1114 , n24 );
buf ( n1115 , n25 );
buf ( n1116 , n26 );
buf ( n1117 , n27 );
buf ( n1118 , n28 );
buf ( n1119 , n29 );
buf ( n1120 , n30 );
buf ( n1121 , n31 );
buf ( n1122 , n32 );
buf ( n1123 , n33 );
buf ( n1124 , n34 );
buf ( n1125 , n35 );
buf ( n1126 , n36 );
buf ( n1127 , n37 );
buf ( n1128 , n38 );
buf ( n1129 , n39 );
buf ( n1130 , n40 );
buf ( n1131 , n41 );
buf ( n1132 , n42 );
buf ( n1133 , n43 );
buf ( n1134 , n44 );
buf ( n1135 , n45 );
buf ( n1136 , n46 );
buf ( n1137 , n47 );
buf ( n1138 , n48 );
buf ( n1139 , n49 );
buf ( n1140 , n50 );
buf ( n1141 , n51 );
buf ( n1142 , n52 );
buf ( n1143 , n53 );
buf ( n1144 , n54 );
buf ( n1145 , n55 );
buf ( n1146 , n56 );
buf ( n1147 , n57 );
buf ( n1148 , n58 );
buf ( n1149 , n59 );
buf ( n1150 , n60 );
buf ( n1151 , n61 );
buf ( n1152 , n62 );
buf ( n1153 , n63 );
buf ( n1154 , n64 );
buf ( n1155 , n65 );
buf ( n1156 , n66 );
buf ( n1157 , n67 );
buf ( n1158 , n68 );
buf ( n1159 , n69 );
buf ( n1160 , n70 );
buf ( n1161 , n71 );
buf ( n1162 , n72 );
buf ( n1163 , n73 );
buf ( n1164 , n74 );
buf ( n1165 , n75 );
buf ( n1166 , n76 );
buf ( n1167 , n77 );
buf ( n1168 , n78 );
buf ( n1169 , n79 );
buf ( n1170 , n80 );
buf ( n1171 , n81 );
buf ( n1172 , n82 );
buf ( n1173 , n83 );
buf ( n1174 , n84 );
buf ( n1175 , n85 );
buf ( n1176 , n86 );
buf ( n1177 , n87 );
buf ( n1178 , n88 );
buf ( n1179 , n89 );
buf ( n1180 , n90 );
buf ( n1181 , n91 );
buf ( n1182 , n92 );
buf ( n1183 , n93 );
buf ( n1184 , n94 );
buf ( n1185 , n95 );
buf ( n1186 , n96 );
buf ( n1187 , n97 );
buf ( n1188 , n98 );
buf ( n1189 , n99 );
buf ( n1190 , n100 );
buf ( n1191 , n101 );
buf ( n1192 , n102 );
buf ( n1193 , n103 );
buf ( n1194 , n104 );
buf ( n1195 , n105 );
buf ( n1196 , n106 );
buf ( n1197 , n107 );
buf ( n1198 , n108 );
buf ( n1199 , n109 );
buf ( n1200 , n110 );
buf ( n1201 , n111 );
buf ( n1202 , n112 );
buf ( n1203 , n113 );
buf ( n1204 , n114 );
buf ( n1205 , n115 );
buf ( n1206 , n116 );
buf ( n1207 , n117 );
buf ( n1208 , n118 );
buf ( n1209 , n119 );
buf ( n1210 , n120 );
buf ( n1211 , n121 );
buf ( n1212 , n122 );
buf ( n1213 , n123 );
buf ( n1214 , n124 );
buf ( n1215 , n125 );
buf ( n1216 , n126 );
buf ( n1217 , n127 );
buf ( n1218 , n128 );
buf ( n1219 , n129 );
buf ( n1220 , n130 );
buf ( n1221 , n131 );
buf ( n1222 , n132 );
buf ( n1223 , n133 );
buf ( n1224 , n134 );
buf ( n1225 , n135 );
buf ( n1226 , n136 );
buf ( n1227 , n137 );
buf ( n1228 , n138 );
buf ( n1229 , n139 );
buf ( n1230 , n140 );
buf ( n1231 , n141 );
buf ( n1232 , n142 );
buf ( n1233 , n143 );
buf ( n1234 , n144 );
buf ( n1235 , n145 );
buf ( n1236 , n146 );
buf ( n1237 , n147 );
buf ( n1238 , n148 );
buf ( n1239 , n149 );
buf ( n1240 , n150 );
buf ( n1241 , n151 );
buf ( n1242 , n152 );
buf ( n1243 , n153 );
buf ( n1244 , n154 );
buf ( n1245 , n155 );
buf ( n1246 , n156 );
buf ( n1247 , n157 );
buf ( n1248 , n158 );
buf ( n1249 , n159 );
buf ( n160 , n1250 );
buf ( n161 , n1251 );
buf ( n162 , n1252 );
buf ( n163 , n1253 );
buf ( n164 , n1254 );
buf ( n165 , n1255 );
buf ( n166 , n1256 );
buf ( n167 , n1257 );
buf ( n168 , n1258 );
buf ( n169 , n1259 );
buf ( n170 , n1260 );
buf ( n171 , n1261 );
buf ( n172 , n1262 );
buf ( n173 , n1263 );
buf ( n174 , n1264 );
buf ( n175 , n1265 );
buf ( n176 , n1266 );
buf ( n177 , n1267 );
buf ( n178 , n1268 );
buf ( n179 , n1269 );
buf ( n180 , n1270 );
buf ( n181 , n1271 );
buf ( n182 , n1272 );
buf ( n183 , n1273 );
buf ( n184 , n1274 );
buf ( n185 , n1275 );
buf ( n186 , n1276 );
buf ( n187 , n1277 );
buf ( n188 , n1278 );
buf ( n189 , n1279 );
buf ( n190 , n1280 );
buf ( n191 , n1281 );
buf ( n192 , n1282 );
buf ( n193 , n1283 );
buf ( n194 , n1284 );
buf ( n195 , n1285 );
buf ( n196 , n1286 );
buf ( n197 , n1287 );
buf ( n198 , n1288 );
buf ( n199 , n1289 );
buf ( n200 , n1290 );
buf ( n201 , n1291 );
buf ( n202 , n1292 );
buf ( n203 , n1293 );
buf ( n204 , n1294 );
buf ( n205 , n1295 );
buf ( n206 , n1296 );
buf ( n207 , n1297 );
buf ( n208 , n1298 );
buf ( n209 , n1299 );
buf ( n210 , n1300 );
buf ( n211 , n1301 );
buf ( n212 , n1302 );
buf ( n213 , n1303 );
buf ( n214 , n1304 );
buf ( n215 , n1305 );
buf ( n216 , n1306 );
buf ( n217 , n1307 );
buf ( n218 , n1308 );
buf ( n219 , n1309 );
buf ( n220 , n1310 );
buf ( n221 , n1311 );
buf ( n222 , n1312 );
buf ( n223 , n1313 );
buf ( n224 , n1314 );
buf ( n225 , n1315 );
buf ( n226 , n1316 );
buf ( n227 , n1317 );
buf ( n228 , n1318 );
buf ( n229 , n1319 );
buf ( n230 , n1320 );
buf ( n231 , n1321 );
buf ( n232 , n1322 );
buf ( n233 , n1323 );
buf ( n234 , n1324 );
buf ( n235 , n1325 );
buf ( n236 , n1326 );
buf ( n237 , n1327 );
buf ( n238 , n1328 );
buf ( n239 , n1329 );
buf ( n240 , n1330 );
buf ( n241 , n1331 );
buf ( n242 , n1332 );
buf ( n243 , n1333 );
buf ( n244 , n1334 );
buf ( n245 , n1335 );
buf ( n246 , n1336 );
buf ( n247 , n1337 );
buf ( n248 , n1338 );
buf ( n249 , n1339 );
buf ( n250 , n1340 );
buf ( n251 , n1341 );
buf ( n252 , n1342 );
buf ( n253 , n1343 );
buf ( n254 , n1344 );
buf ( n255 , n1345 );
buf ( n256 , n1346 );
buf ( n257 , n1347 );
buf ( n258 , n1348 );
buf ( n259 , n1349 );
buf ( n260 , n1350 );
buf ( n261 , n1351 );
buf ( n262 , n1352 );
buf ( n263 , n1353 );
buf ( n264 , n1354 );
buf ( n265 , n1355 );
buf ( n266 , n1356 );
buf ( n267 , n1357 );
buf ( n268 , n1358 );
buf ( n269 , n1359 );
buf ( n270 , n1360 );
buf ( n271 , n1361 );
buf ( n272 , n1362 );
buf ( n273 , n1363 );
buf ( n274 , n1364 );
buf ( n275 , n1365 );
buf ( n276 , n1366 );
buf ( n277 , n1367 );
buf ( n278 , n1368 );
buf ( n279 , n1369 );
buf ( n280 , n1370 );
buf ( n281 , n1371 );
buf ( n282 , n1372 );
buf ( n283 , n1373 );
buf ( n284 , n1374 );
buf ( n285 , n1375 );
buf ( n286 , n1376 );
buf ( n287 , n1377 );
buf ( n288 , n1378 );
buf ( n289 , n1379 );
buf ( n290 , n1380 );
buf ( n291 , n1381 );
buf ( n292 , n1382 );
buf ( n293 , n1383 );
buf ( n294 , n1384 );
buf ( n295 , n1385 );
buf ( n296 , n1386 );
buf ( n297 , n1387 );
buf ( n298 , n1388 );
buf ( n299 , n1389 );
buf ( n300 , n1390 );
buf ( n301 , n1391 );
buf ( n302 , n1392 );
buf ( n303 , n1393 );
buf ( n304 , n1394 );
buf ( n305 , n1395 );
buf ( n306 , n1396 );
buf ( n307 , n1397 );
buf ( n308 , n1398 );
buf ( n309 , n1399 );
buf ( n310 , n1400 );
buf ( n311 , n1401 );
buf ( n312 , n1402 );
buf ( n313 , n1403 );
buf ( n314 , n1404 );
buf ( n315 , n1405 );
buf ( n316 , n1406 );
buf ( n317 , n1407 );
buf ( n318 , n1408 );
buf ( n319 , n1409 );
buf ( n320 , n1410 );
buf ( n321 , n1411 );
buf ( n322 , n1412 );
buf ( n323 , n1413 );
buf ( n324 , n1414 );
buf ( n325 , n1415 );
buf ( n326 , n1416 );
buf ( n327 , n1417 );
buf ( n328 , n1418 );
buf ( n329 , n1419 );
buf ( n330 , n1420 );
buf ( n331 , n1421 );
buf ( n332 , n1422 );
buf ( n333 , n1423 );
buf ( n334 , n1424 );
buf ( n335 , n1425 );
buf ( n336 , n1426 );
buf ( n337 , n1427 );
buf ( n338 , n1428 );
buf ( n339 , n1429 );
buf ( n340 , n1430 );
buf ( n341 , n1431 );
buf ( n342 , n1432 );
buf ( n343 , n1433 );
buf ( n344 , n1434 );
buf ( n345 , n1435 );
buf ( n346 , n1436 );
buf ( n347 , n1437 );
buf ( n348 , n1438 );
buf ( n349 , n1439 );
buf ( n350 , n1440 );
buf ( n351 , n1441 );
buf ( n352 , n1442 );
buf ( n353 , n1443 );
buf ( n354 , n1444 );
buf ( n355 , n1445 );
buf ( n356 , n1446 );
buf ( n357 , n1447 );
buf ( n358 , n1448 );
buf ( n359 , n1449 );
buf ( n360 , n1450 );
buf ( n361 , n1451 );
buf ( n362 , n1452 );
buf ( n363 , n1453 );
buf ( n364 , n1454 );
buf ( n365 , n1455 );
buf ( n366 , n1456 );
buf ( n367 , n1457 );
buf ( n368 , n1458 );
buf ( n369 , n1459 );
buf ( n370 , n1460 );
buf ( n371 , n1461 );
buf ( n372 , n1462 );
buf ( n373 , n1463 );
buf ( n374 , n1464 );
buf ( n375 , n1465 );
buf ( n376 , n1466 );
buf ( n377 , n1467 );
buf ( n378 , n1468 );
buf ( n379 , n1469 );
buf ( n380 , n1470 );
buf ( n381 , n1471 );
buf ( n382 , n1472 );
buf ( n383 , n1473 );
buf ( n384 , n1474 );
buf ( n385 , n1475 );
buf ( n386 , n1476 );
buf ( n387 , n1477 );
buf ( n388 , n1478 );
buf ( n389 , n1479 );
buf ( n390 , n1480 );
buf ( n391 , n1481 );
buf ( n392 , n1482 );
buf ( n393 , n1483 );
buf ( n394 , n1484 );
buf ( n395 , n1485 );
buf ( n396 , n1486 );
buf ( n397 , n1487 );
buf ( n398 , n1488 );
buf ( n399 , n1489 );
buf ( n400 , n1490 );
buf ( n401 , n1491 );
buf ( n402 , n1492 );
buf ( n403 , n1493 );
buf ( n404 , n1494 );
buf ( n405 , n1495 );
buf ( n406 , n1496 );
buf ( n407 , n1497 );
buf ( n408 , n1498 );
buf ( n409 , n1499 );
buf ( n410 , n1500 );
buf ( n411 , n1501 );
buf ( n412 , n1502 );
buf ( n413 , n1503 );
buf ( n414 , n1504 );
buf ( n415 , n1505 );
buf ( n416 , n1506 );
buf ( n417 , n1507 );
buf ( n418 , n1508 );
buf ( n419 , n1509 );
buf ( n420 , n1510 );
buf ( n421 , n1511 );
buf ( n422 , n1512 );
buf ( n423 , n1513 );
buf ( n424 , n1514 );
buf ( n425 , n1515 );
buf ( n426 , n1516 );
buf ( n427 , n1517 );
buf ( n428 , n1518 );
buf ( n429 , n1519 );
buf ( n430 , n1520 );
buf ( n431 , n1521 );
buf ( n432 , n1522 );
buf ( n433 , n1523 );
buf ( n434 , n1524 );
buf ( n435 , n1525 );
buf ( n436 , n1526 );
buf ( n437 , n1527 );
buf ( n438 , n1528 );
buf ( n439 , n1529 );
buf ( n440 , n1530 );
buf ( n441 , n1531 );
buf ( n442 , n1532 );
buf ( n443 , n1533 );
buf ( n444 , n1534 );
buf ( n445 , n1535 );
buf ( n446 , n1536 );
buf ( n447 , n1537 );
buf ( n448 , n1538 );
buf ( n449 , n1539 );
buf ( n450 , n1540 );
buf ( n451 , n1541 );
buf ( n452 , n1542 );
buf ( n453 , n1543 );
buf ( n454 , n1544 );
buf ( n455 , n1545 );
buf ( n456 , n1546 );
buf ( n457 , n1547 );
buf ( n458 , n1548 );
buf ( n459 , n1549 );
buf ( n460 , n1550 );
buf ( n461 , n1551 );
buf ( n462 , n1552 );
buf ( n463 , n1553 );
buf ( n464 , n1554 );
buf ( n465 , n1555 );
buf ( n466 , n1556 );
buf ( n467 , n1557 );
buf ( n468 , n1558 );
buf ( n469 , n1559 );
buf ( n470 , n1560 );
buf ( n471 , n1561 );
buf ( n472 , n1562 );
buf ( n473 , n1563 );
buf ( n474 , n1564 );
buf ( n475 , n1565 );
buf ( n476 , n1566 );
buf ( n477 , n1567 );
buf ( n478 , n1568 );
buf ( n479 , n1569 );
buf ( n480 , n1570 );
buf ( n481 , n1571 );
buf ( n482 , n1572 );
buf ( n483 , n1573 );
buf ( n484 , n1574 );
buf ( n485 , n1575 );
buf ( n486 , n1576 );
buf ( n487 , n1577 );
buf ( n488 , n1578 );
buf ( n489 , n1579 );
buf ( n490 , n1580 );
buf ( n491 , n1581 );
buf ( n492 , n1582 );
buf ( n493 , n1583 );
buf ( n494 , n1584 );
buf ( n495 , n1585 );
buf ( n496 , n1586 );
buf ( n497 , n1587 );
buf ( n498 , n1588 );
buf ( n499 , n1589 );
buf ( n500 , n1590 );
buf ( n501 , n1591 );
buf ( n502 , n1592 );
buf ( n503 , n1593 );
buf ( n504 , n1594 );
buf ( n505 , n1595 );
buf ( n506 , n1596 );
buf ( n507 , n1597 );
buf ( n508 , n1598 );
buf ( n509 , n1599 );
buf ( n510 , n1600 );
buf ( n511 , n1601 );
buf ( n512 , n1602 );
buf ( n513 , n1603 );
buf ( n514 , n1604 );
buf ( n515 , n1605 );
buf ( n516 , n1606 );
buf ( n517 , n1607 );
buf ( n518 , n1608 );
buf ( n519 , n1609 );
buf ( n520 , n1610 );
buf ( n521 , n1611 );
buf ( n522 , n1612 );
buf ( n523 , n1613 );
buf ( n524 , n1614 );
buf ( n525 , n1615 );
buf ( n526 , n1616 );
buf ( n527 , n1617 );
buf ( n528 , n1618 );
buf ( n529 , n1619 );
buf ( n530 , n1620 );
buf ( n531 , n1621 );
buf ( n532 , n1622 );
buf ( n533 , n1623 );
buf ( n534 , n1624 );
buf ( n535 , n1625 );
buf ( n536 , n1626 );
buf ( n537 , n1627 );
buf ( n538 , n1628 );
buf ( n539 , n1629 );
buf ( n540 , n1630 );
buf ( n541 , n1631 );
buf ( n542 , n1632 );
buf ( n543 , n1633 );
buf ( n544 , n1634 );
buf ( n1250 , C0 );
buf ( n1251 , C0 );
buf ( n1252 , C0 );
buf ( n1253 , C0 );
buf ( n1254 , C0 );
buf ( n1255 , C0 );
buf ( n1256 , C0 );
buf ( n1257 , C0 );
buf ( n1258 , C0 );
buf ( n1259 , C0 );
buf ( n1260 , C0 );
buf ( n1261 , C0 );
buf ( n1262 , C0 );
buf ( n1263 , C0 );
buf ( n1264 , C0 );
buf ( n1265 , C0 );
buf ( n1266 , C0 );
buf ( n1267 , C0 );
buf ( n1268 , C0 );
buf ( n1269 , C0 );
buf ( n1270 , C0 );
buf ( n1271 , C0 );
buf ( n1272 , C0 );
buf ( n1273 , C0 );
buf ( n1274 , C0 );
buf ( n1275 , C0 );
buf ( n1276 , C0 );
buf ( n1277 , C0 );
buf ( n1278 , C0 );
buf ( n1279 , C0 );
buf ( n1280 , C0 );
buf ( n1281 , n75399 );
buf ( n1282 , n75401 );
buf ( n1283 , n75403 );
buf ( n1284 , n75405 );
buf ( n1285 , n75407 );
buf ( n1286 , n75409 );
buf ( n1287 , n75411 );
buf ( n1288 , n75413 );
buf ( n1289 , n75415 );
buf ( n1290 , n75417 );
buf ( n1291 , n75419 );
buf ( n1292 , n75421 );
buf ( n1293 , n75423 );
buf ( n1294 , n75425 );
buf ( n1295 , n75427 );
buf ( n1296 , n75429 );
buf ( n1297 , n75431 );
buf ( n1298 , n75433 );
buf ( n1299 , n75435 );
buf ( n1300 , n75437 );
buf ( n1301 , n75439 );
buf ( n1302 , n75441 );
buf ( n1303 , n75443 );
buf ( n1304 , n75445 );
buf ( n1305 , n75447 );
buf ( n1306 , n75449 );
buf ( n1307 , n75451 );
buf ( n1308 , n75453 );
buf ( n1309 , n75455 );
buf ( n1310 , n75457 );
buf ( n1311 , n75459 );
buf ( n1312 , n75461 );
buf ( n1313 , n75463 );
buf ( n1314 , n75465 );
buf ( n1315 , n75467 );
buf ( n1316 , n75469 );
buf ( n1317 , n75471 );
buf ( n1318 , n75473 );
buf ( n1319 , n75475 );
buf ( n1320 , n75477 );
buf ( n1321 , n75479 );
buf ( n1322 , n75481 );
buf ( n1323 , n75483 );
buf ( n1324 , n75485 );
buf ( n1325 , n75487 );
buf ( n1326 , n75489 );
buf ( n1327 , n75491 );
buf ( n1328 , n75493 );
buf ( n1329 , n75495 );
buf ( n1330 , n75497 );
buf ( n1331 , n75499 );
buf ( n1332 , n75501 );
buf ( n1333 , n75503 );
buf ( n1334 , n75505 );
buf ( n1335 , n75507 );
buf ( n1336 , n75509 );
buf ( n1337 , n75511 );
buf ( n1338 , n75513 );
buf ( n1339 , n75515 );
buf ( n1340 , n75517 );
buf ( n1341 , n75519 );
buf ( n1342 , n75521 );
buf ( n1343 , n75523 );
buf ( n1344 , n75525 );
buf ( n1345 , n75527 );
buf ( n1346 , n75529 );
buf ( n1347 , n75531 );
buf ( n1348 , n75533 );
buf ( n1349 , n75535 );
buf ( n1350 , n75537 );
buf ( n1351 , n75539 );
buf ( n1352 , n75541 );
buf ( n1353 , n75543 );
buf ( n1354 , n75545 );
buf ( n1355 , n75547 );
buf ( n1356 , n75549 );
buf ( n1357 , n75551 );
buf ( n1358 , n75553 );
buf ( n1359 , n75555 );
buf ( n1360 , n75557 );
buf ( n1361 , n75559 );
buf ( n1362 , n75561 );
buf ( n1363 , n75563 );
buf ( n1364 , n75565 );
buf ( n1365 , n75567 );
buf ( n1366 , n75569 );
buf ( n1367 , n75571 );
buf ( n1368 , n75573 );
buf ( n1369 , n75575 );
buf ( n1370 , n75577 );
buf ( n1371 , n75579 );
buf ( n1372 , n75581 );
buf ( n1373 , n75583 );
buf ( n1374 , n75585 );
buf ( n1375 , n75587 );
buf ( n1376 , n75589 );
buf ( n1377 , n75591 );
buf ( n1378 , C0 );
buf ( n1379 , C0 );
buf ( n1380 , C0 );
buf ( n1381 , C0 );
buf ( n1382 , C0 );
buf ( n1383 , C0 );
buf ( n1384 , C0 );
buf ( n1385 , C0 );
buf ( n1386 , C0 );
buf ( n1387 , C0 );
buf ( n1388 , C0 );
buf ( n1389 , C0 );
buf ( n1390 , C0 );
buf ( n1391 , C0 );
buf ( n1392 , C0 );
buf ( n1393 , C0 );
buf ( n1394 , C0 );
buf ( n1395 , C0 );
buf ( n1396 , C0 );
buf ( n1397 , C0 );
buf ( n1398 , C0 );
buf ( n1399 , C0 );
buf ( n1400 , n64296 );
buf ( n1401 , n64298 );
buf ( n1402 , n64300 );
buf ( n1403 , n64302 );
buf ( n1404 , n64304 );
buf ( n1405 , n64306 );
buf ( n1406 , n64308 );
buf ( n1407 , n64310 );
buf ( n1408 , n64312 );
buf ( n1409 , n64314 );
buf ( n1410 , n64316 );
buf ( n1411 , n64318 );
buf ( n1412 , n64320 );
buf ( n1413 , n64322 );
buf ( n1414 , n64324 );
buf ( n1415 , n64326 );
buf ( n1416 , n64328 );
buf ( n1417 , n64330 );
buf ( n1418 , n64332 );
buf ( n1419 , n64334 );
buf ( n1420 , n64336 );
buf ( n1421 , n64338 );
buf ( n1422 , n64340 );
buf ( n1423 , n64342 );
buf ( n1424 , n64344 );
buf ( n1425 , n64346 );
buf ( n1426 , n64348 );
buf ( n1427 , n64350 );
buf ( n1428 , n64352 );
buf ( n1429 , n64354 );
buf ( n1430 , n64356 );
buf ( n1431 , n64358 );
buf ( n1432 , n64360 );
buf ( n1433 , n64362 );
buf ( n1434 , n64364 );
buf ( n1435 , n64366 );
buf ( n1436 , n64368 );
buf ( n1437 , n64370 );
buf ( n1438 , n64372 );
buf ( n1439 , n64374 );
buf ( n1440 , n64376 );
buf ( n1441 , n64378 );
buf ( n1442 , n64380 );
buf ( n1443 , n64382 );
buf ( n1444 , n64384 );
buf ( n1445 , n64386 );
buf ( n1446 , n64388 );
buf ( n1447 , n64390 );
buf ( n1448 , n64392 );
buf ( n1449 , n64394 );
buf ( n1450 , n64396 );
buf ( n1451 , n64398 );
buf ( n1452 , n64400 );
buf ( n1453 , n64402 );
buf ( n1454 , n64404 );
buf ( n1455 , n64406 );
buf ( n1456 , n64408 );
buf ( n1457 , n64410 );
buf ( n1458 , n64412 );
buf ( n1459 , n64414 );
buf ( n1460 , n64416 );
buf ( n1461 , n64418 );
buf ( n1462 , n64420 );
buf ( n1463 , n64422 );
buf ( n1464 , n64424 );
buf ( n1465 , n64426 );
buf ( n1466 , n64428 );
buf ( n1467 , n64430 );
buf ( n1468 , n64432 );
buf ( n1469 , n64434 );
buf ( n1470 , n64436 );
buf ( n1471 , n64438 );
buf ( n1472 , n64440 );
buf ( n1473 , n64442 );
buf ( n1474 , n64444 );
buf ( n1475 , n64446 );
buf ( n1476 , n64448 );
buf ( n1477 , n64450 );
buf ( n1478 , n64452 );
buf ( n1479 , n64454 );
buf ( n1480 , n64456 );
buf ( n1481 , n64458 );
buf ( n1482 , n64460 );
buf ( n1483 , n64462 );
buf ( n1484 , n64464 );
buf ( n1485 , n64466 );
buf ( n1486 , n64468 );
buf ( n1487 , n64470 );
buf ( n1488 , n64472 );
buf ( n1489 , n64474 );
buf ( n1490 , n64476 );
buf ( n1491 , n64478 );
buf ( n1492 , n64480 );
buf ( n1493 , n64482 );
buf ( n1494 , n64484 );
buf ( n1495 , n64486 );
buf ( n1496 , n64488 );
buf ( n1497 , n64490 );
buf ( n1498 , n64492 );
buf ( n1499 , n64494 );
buf ( n1500 , n64496 );
buf ( n1501 , n64498 );
buf ( n1502 , n64500 );
buf ( n1503 , n64502 );
buf ( n1504 , n64504 );
buf ( n1505 , n64506 );
buf ( n1506 , n51393 );
buf ( n1507 , n51395 );
buf ( n1508 , n51397 );
buf ( n1509 , n51399 );
buf ( n1510 , n51401 );
buf ( n1511 , n51403 );
buf ( n1512 , n51405 );
buf ( n1513 , n51407 );
buf ( n1514 , n51409 );
buf ( n1515 , n51411 );
buf ( n1516 , n51413 );
buf ( n1517 , n51415 );
buf ( n1518 , n51417 );
buf ( n1519 , n51419 );
buf ( n1520 , n51421 );
buf ( n1521 , n51423 );
buf ( n1522 , n51425 );
buf ( n1523 , n51427 );
buf ( n1524 , n51429 );
buf ( n1525 , n51431 );
buf ( n1526 , n51433 );
buf ( n1527 , n51435 );
buf ( n1528 , n51437 );
buf ( n1529 , n51439 );
buf ( n1530 , n51441 );
buf ( n1531 , n51443 );
buf ( n1532 , n51445 );
buf ( n1533 , n51447 );
buf ( n1534 , n51449 );
buf ( n1535 , n51451 );
buf ( n1536 , n51453 );
buf ( n1537 , n51455 );
buf ( n1538 , n51457 );
buf ( n1539 , n51459 );
buf ( n1540 , n51461 );
buf ( n1541 , n51463 );
buf ( n1542 , n51465 );
buf ( n1543 , n51467 );
buf ( n1544 , n51469 );
buf ( n1545 , n51471 );
buf ( n1546 , n51473 );
buf ( n1547 , n51475 );
buf ( n1548 , n51477 );
buf ( n1549 , n51479 );
buf ( n1550 , n51481 );
buf ( n1551 , n51483 );
buf ( n1552 , n51485 );
buf ( n1553 , n51487 );
buf ( n1554 , n51489 );
buf ( n1555 , n51491 );
buf ( n1556 , n51493 );
buf ( n1557 , n51495 );
buf ( n1558 , n51497 );
buf ( n1559 , n51499 );
buf ( n1560 , n51501 );
buf ( n1561 , n51503 );
buf ( n1562 , n51505 );
buf ( n1563 , n51507 );
buf ( n1564 , n51509 );
buf ( n1565 , n51511 );
buf ( n1566 , n51513 );
buf ( n1567 , n51515 );
buf ( n1568 , n51517 );
buf ( n1569 , n51519 );
buf ( n1570 , n51521 );
buf ( n1571 , n51523 );
buf ( n1572 , n51525 );
buf ( n1573 , n51527 );
buf ( n1574 , n51529 );
buf ( n1575 , n51531 );
buf ( n1576 , n51533 );
buf ( n1577 , n51535 );
buf ( n1578 , n51537 );
buf ( n1579 , n51539 );
buf ( n1580 , n51541 );
buf ( n1581 , n51543 );
buf ( n1582 , n51545 );
buf ( n1583 , n51547 );
buf ( n1584 , n51549 );
buf ( n1585 , n51551 );
buf ( n1586 , n51553 );
buf ( n1587 , n51555 );
buf ( n1588 , n51557 );
buf ( n1589 , n51559 );
buf ( n1590 , n51561 );
buf ( n1591 , n51563 );
buf ( n1592 , n51565 );
buf ( n1593 , n51567 );
buf ( n1594 , n51569 );
buf ( n1595 , n51571 );
buf ( n1596 , n51573 );
buf ( n1597 , n51575 );
buf ( n1598 , n51577 );
buf ( n1599 , n51579 );
buf ( n1600 , n51581 );
buf ( n1601 , n51583 );
buf ( n1602 , n51585 );
buf ( n1603 , n51587 );
buf ( n1604 , n51589 );
buf ( n1605 , n51591 );
buf ( n1606 , n51593 );
buf ( n1607 , n51595 );
buf ( n1608 , n51597 );
buf ( n1609 , n51599 );
buf ( n1610 , n51601 );
buf ( n1611 , n51603 );
buf ( n1612 , n51605 );
buf ( n1613 , n51608 );
buf ( n1614 , n51611 );
buf ( n1615 , n51614 );
buf ( n1616 , n51617 );
buf ( n1617 , n51620 );
buf ( n1618 , n51623 );
buf ( n1619 , n51626 );
buf ( n1620 , n51629 );
buf ( n1621 , n51632 );
buf ( n1622 , n51635 );
buf ( n1623 , n51638 );
buf ( n1624 , n51641 );
buf ( n1625 , n51644 );
buf ( n1626 , n51647 );
buf ( n1627 , n51650 );
buf ( n1628 , n51653 );
buf ( n1629 , n51656 );
buf ( n1630 , n51659 );
buf ( n1631 , n51662 );
buf ( n1632 , n51665 );
buf ( n1633 , n51668 );
buf ( n1634 , n51670 );
buf ( n1635 , n1122 );
buf ( n1636 , n1635 );
buf ( n1637 , n1156 );
buf ( n1638 , n1637 );
buf ( n1639 , n1157 );
buf ( n1640 , n1639 );
xor ( n1641 , n1638 , n1640 );
buf ( n1642 , n1158 );
buf ( n1643 , n1642 );
xor ( n1644 , n1640 , n1643 );
not ( n1645 , n1644 );
and ( n1646 , n1641 , n1645 );
and ( n1647 , n1636 , n1646 );
not ( n1648 , n1647 );
and ( n1649 , n1640 , n1643 );
not ( n1650 , n1649 );
and ( n1651 , n1638 , n1650 );
xnor ( n1652 , n1648 , n1651 );
not ( n1653 , n1652 );
buf ( n1654 , n1124 );
buf ( n1655 , n1654 );
buf ( n1656 , n1154 );
buf ( n1657 , n1656 );
buf ( n1658 , n1155 );
buf ( n1659 , n1658 );
xor ( n1660 , n1657 , n1659 );
xor ( n1661 , n1659 , n1638 );
not ( n1662 , n1661 );
and ( n1663 , n1660 , n1662 );
and ( n1664 , n1655 , n1663 );
buf ( n1665 , n1123 );
buf ( n1666 , n1665 );
and ( n1667 , n1666 , n1661 );
nor ( n1668 , n1664 , n1667 );
and ( n1669 , n1659 , n1638 );
not ( n1670 , n1669 );
and ( n1671 , n1657 , n1670 );
xnor ( n1672 , n1668 , n1671 );
and ( n1673 , n1653 , n1672 );
buf ( n1674 , n1125 );
buf ( n1675 , n1674 );
and ( n1676 , n1675 , n1657 );
and ( n1677 , n1672 , n1676 );
and ( n1678 , n1653 , n1676 );
or ( n1679 , n1673 , n1677 , n1678 );
buf ( n1680 , n1652 );
xor ( n1681 , n1679 , n1680 );
not ( n1682 , n1651 );
and ( n1683 , n1666 , n1663 );
and ( n1684 , n1636 , n1661 );
nor ( n1685 , n1683 , n1684 );
xnor ( n1686 , n1685 , n1671 );
xor ( n1687 , n1682 , n1686 );
and ( n1688 , n1655 , n1657 );
xor ( n1689 , n1687 , n1688 );
xor ( n1690 , n1681 , n1689 );
buf ( n1691 , n1159 );
buf ( n1692 , n1691 );
buf ( n1693 , n1160 );
buf ( n1694 , n1693 );
and ( n1695 , n1692 , n1694 );
not ( n1696 , n1695 );
and ( n1697 , n1643 , n1696 );
not ( n1698 , n1697 );
and ( n1699 , n1666 , n1646 );
and ( n1700 , n1636 , n1644 );
nor ( n1701 , n1699 , n1700 );
xnor ( n1702 , n1701 , n1651 );
and ( n1703 , n1698 , n1702 );
buf ( n1704 , n1126 );
buf ( n1705 , n1704 );
and ( n1706 , n1705 , n1657 );
and ( n1707 , n1702 , n1706 );
and ( n1708 , n1698 , n1706 );
or ( n1709 , n1703 , n1707 , n1708 );
and ( n1710 , n1655 , n1646 );
and ( n1711 , n1666 , n1644 );
nor ( n1712 , n1710 , n1711 );
xnor ( n1713 , n1712 , n1651 );
and ( n1714 , n1705 , n1663 );
and ( n1715 , n1675 , n1661 );
nor ( n1716 , n1714 , n1715 );
xnor ( n1717 , n1716 , n1671 );
and ( n1718 , n1713 , n1717 );
buf ( n1719 , n1127 );
buf ( n1720 , n1719 );
and ( n1721 , n1720 , n1657 );
and ( n1722 , n1717 , n1721 );
and ( n1723 , n1713 , n1721 );
or ( n1724 , n1718 , n1722 , n1723 );
xor ( n1725 , n1643 , n1692 );
xor ( n1726 , n1692 , n1694 );
not ( n1727 , n1726 );
and ( n1728 , n1725 , n1727 );
and ( n1729 , n1636 , n1728 );
not ( n1730 , n1729 );
xnor ( n1731 , n1730 , n1697 );
buf ( n1732 , n1731 );
and ( n1733 , n1724 , n1732 );
and ( n1734 , n1675 , n1663 );
and ( n1735 , n1655 , n1661 );
nor ( n1736 , n1734 , n1735 );
xnor ( n1737 , n1736 , n1671 );
and ( n1738 , n1732 , n1737 );
and ( n1739 , n1724 , n1737 );
or ( n1740 , n1733 , n1738 , n1739 );
and ( n1741 , n1709 , n1740 );
xor ( n1742 , n1653 , n1672 );
xor ( n1743 , n1742 , n1676 );
and ( n1744 , n1740 , n1743 );
and ( n1745 , n1709 , n1743 );
or ( n1746 , n1741 , n1744 , n1745 );
xor ( n1747 , n1690 , n1746 );
xor ( n1748 , n1709 , n1740 );
xor ( n1749 , n1748 , n1743 );
buf ( n1750 , n1161 );
buf ( n1751 , n1750 );
buf ( n1752 , n1162 );
buf ( n1753 , n1752 );
and ( n1754 , n1751 , n1753 );
not ( n1755 , n1754 );
and ( n1756 , n1694 , n1755 );
not ( n1757 , n1756 );
and ( n1758 , n1666 , n1728 );
and ( n1759 , n1636 , n1726 );
nor ( n1760 , n1758 , n1759 );
xnor ( n1761 , n1760 , n1697 );
and ( n1762 , n1757 , n1761 );
and ( n1763 , n1720 , n1663 );
and ( n1764 , n1705 , n1661 );
nor ( n1765 , n1763 , n1764 );
xnor ( n1766 , n1765 , n1671 );
and ( n1767 , n1761 , n1766 );
and ( n1768 , n1757 , n1766 );
or ( n1769 , n1762 , n1767 , n1768 );
not ( n1770 , n1731 );
and ( n1771 , n1769 , n1770 );
xor ( n1772 , n1713 , n1717 );
xor ( n1773 , n1772 , n1721 );
and ( n1774 , n1770 , n1773 );
and ( n1775 , n1769 , n1773 );
or ( n1776 , n1771 , n1774 , n1775 );
xor ( n1777 , n1698 , n1702 );
xor ( n1778 , n1777 , n1706 );
and ( n1779 , n1776 , n1778 );
xor ( n1780 , n1724 , n1732 );
xor ( n1781 , n1780 , n1737 );
and ( n1782 , n1778 , n1781 );
and ( n1783 , n1776 , n1781 );
or ( n1784 , n1779 , n1782 , n1783 );
and ( n1785 , n1749 , n1784 );
xor ( n1786 , n1776 , n1778 );
xor ( n1787 , n1786 , n1781 );
and ( n1788 , n1655 , n1728 );
and ( n1789 , n1666 , n1726 );
nor ( n1790 , n1788 , n1789 );
xnor ( n1791 , n1790 , n1697 );
buf ( n1792 , n1791 );
and ( n1793 , n1675 , n1646 );
and ( n1794 , n1655 , n1644 );
nor ( n1795 , n1793 , n1794 );
xnor ( n1796 , n1795 , n1651 );
and ( n1797 , n1792 , n1796 );
buf ( n1798 , n1128 );
buf ( n1799 , n1798 );
and ( n1800 , n1799 , n1657 );
and ( n1801 , n1796 , n1800 );
and ( n1802 , n1792 , n1800 );
or ( n1803 , n1797 , n1801 , n1802 );
xor ( n1804 , n1694 , n1751 );
xor ( n1805 , n1751 , n1753 );
not ( n1806 , n1805 );
and ( n1807 , n1804 , n1806 );
and ( n1808 , n1636 , n1807 );
not ( n1809 , n1808 );
xnor ( n1810 , n1809 , n1756 );
and ( n1811 , n1799 , n1663 );
and ( n1812 , n1720 , n1661 );
nor ( n1813 , n1811 , n1812 );
xnor ( n1814 , n1813 , n1671 );
and ( n1815 , n1810 , n1814 );
buf ( n1816 , n1129 );
buf ( n1817 , n1816 );
and ( n1818 , n1817 , n1657 );
and ( n1819 , n1814 , n1818 );
and ( n1820 , n1810 , n1818 );
or ( n1821 , n1815 , n1819 , n1820 );
xor ( n1822 , n1757 , n1761 );
xor ( n1823 , n1822 , n1766 );
and ( n1824 , n1821 , n1823 );
xor ( n1825 , n1792 , n1796 );
xor ( n1826 , n1825 , n1800 );
and ( n1827 , n1823 , n1826 );
and ( n1828 , n1821 , n1826 );
or ( n1829 , n1824 , n1827 , n1828 );
and ( n1830 , n1803 , n1829 );
xor ( n1831 , n1769 , n1770 );
xor ( n1832 , n1831 , n1773 );
and ( n1833 , n1829 , n1832 );
and ( n1834 , n1803 , n1832 );
or ( n1835 , n1830 , n1833 , n1834 );
and ( n1836 , n1787 , n1835 );
xor ( n1837 , n1803 , n1829 );
xor ( n1838 , n1837 , n1832 );
and ( n1839 , n1675 , n1728 );
and ( n1840 , n1655 , n1726 );
nor ( n1841 , n1839 , n1840 );
xnor ( n1842 , n1841 , n1697 );
and ( n1843 , n1817 , n1663 );
and ( n1844 , n1799 , n1661 );
nor ( n1845 , n1843 , n1844 );
xnor ( n1846 , n1845 , n1671 );
and ( n1847 , n1842 , n1846 );
buf ( n1848 , n1130 );
buf ( n1849 , n1848 );
and ( n1850 , n1849 , n1657 );
and ( n1851 , n1846 , n1850 );
and ( n1852 , n1842 , n1850 );
or ( n1853 , n1847 , n1851 , n1852 );
not ( n1854 , n1791 );
and ( n1855 , n1853 , n1854 );
and ( n1856 , n1705 , n1646 );
and ( n1857 , n1675 , n1644 );
nor ( n1858 , n1856 , n1857 );
xnor ( n1859 , n1858 , n1651 );
and ( n1860 , n1854 , n1859 );
and ( n1861 , n1853 , n1859 );
or ( n1862 , n1855 , n1860 , n1861 );
buf ( n1863 , n1163 );
buf ( n1864 , n1863 );
buf ( n1865 , n1164 );
buf ( n1866 , n1865 );
and ( n1867 , n1864 , n1866 );
not ( n1868 , n1867 );
and ( n1869 , n1753 , n1868 );
not ( n1870 , n1869 );
and ( n1871 , n1666 , n1807 );
and ( n1872 , n1636 , n1805 );
nor ( n1873 , n1871 , n1872 );
xnor ( n1874 , n1873 , n1756 );
and ( n1875 , n1870 , n1874 );
and ( n1876 , n1720 , n1646 );
and ( n1877 , n1705 , n1644 );
nor ( n1878 , n1876 , n1877 );
xnor ( n1879 , n1878 , n1651 );
and ( n1880 , n1874 , n1879 );
and ( n1881 , n1870 , n1879 );
or ( n1882 , n1875 , n1880 , n1881 );
xor ( n1883 , n1810 , n1814 );
xor ( n1884 , n1883 , n1818 );
and ( n1885 , n1882 , n1884 );
xor ( n1886 , n1853 , n1854 );
xor ( n1887 , n1886 , n1859 );
and ( n1888 , n1884 , n1887 );
and ( n1889 , n1882 , n1887 );
or ( n1890 , n1885 , n1888 , n1889 );
and ( n1891 , n1862 , n1890 );
xor ( n1892 , n1821 , n1823 );
xor ( n1893 , n1892 , n1826 );
and ( n1894 , n1890 , n1893 );
and ( n1895 , n1862 , n1893 );
or ( n1896 , n1891 , n1894 , n1895 );
and ( n1897 , n1838 , n1896 );
xor ( n1898 , n1753 , n1864 );
xor ( n1899 , n1864 , n1866 );
not ( n1900 , n1899 );
and ( n1901 , n1898 , n1900 );
and ( n1902 , n1636 , n1901 );
not ( n1903 , n1902 );
xnor ( n1904 , n1903 , n1869 );
and ( n1905 , n1799 , n1646 );
and ( n1906 , n1720 , n1644 );
nor ( n1907 , n1905 , n1906 );
xnor ( n1908 , n1907 , n1651 );
and ( n1909 , n1904 , n1908 );
and ( n1910 , n1849 , n1663 );
and ( n1911 , n1817 , n1661 );
nor ( n1912 , n1910 , n1911 );
xnor ( n1913 , n1912 , n1671 );
and ( n1914 , n1908 , n1913 );
and ( n1915 , n1904 , n1913 );
or ( n1916 , n1909 , n1914 , n1915 );
and ( n1917 , n1655 , n1807 );
and ( n1918 , n1666 , n1805 );
nor ( n1919 , n1917 , n1918 );
xnor ( n1920 , n1919 , n1756 );
buf ( n1921 , n1920 );
and ( n1922 , n1916 , n1921 );
xor ( n1923 , n1842 , n1846 );
xor ( n1924 , n1923 , n1850 );
and ( n1925 , n1921 , n1924 );
and ( n1926 , n1916 , n1924 );
or ( n1927 , n1922 , n1925 , n1926 );
not ( n1928 , n1920 );
and ( n1929 , n1705 , n1728 );
and ( n1930 , n1675 , n1726 );
nor ( n1931 , n1929 , n1930 );
xnor ( n1932 , n1931 , n1697 );
and ( n1933 , n1928 , n1932 );
buf ( n1934 , n1131 );
buf ( n1935 , n1934 );
and ( n1936 , n1935 , n1657 );
and ( n1937 , n1932 , n1936 );
and ( n1938 , n1928 , n1936 );
or ( n1939 , n1933 , n1937 , n1938 );
xor ( n1940 , n1870 , n1874 );
xor ( n1941 , n1940 , n1879 );
and ( n1942 , n1939 , n1941 );
xor ( n1943 , n1916 , n1921 );
xor ( n1944 , n1943 , n1924 );
and ( n1945 , n1941 , n1944 );
and ( n1946 , n1939 , n1944 );
or ( n1947 , n1942 , n1945 , n1946 );
and ( n1948 , n1927 , n1947 );
xor ( n1949 , n1882 , n1884 );
xor ( n1950 , n1949 , n1887 );
and ( n1951 , n1947 , n1950 );
and ( n1952 , n1927 , n1950 );
or ( n1953 , n1948 , n1951 , n1952 );
xor ( n1954 , n1862 , n1890 );
xor ( n1955 , n1954 , n1893 );
and ( n1956 , n1953 , n1955 );
xor ( n1957 , n1927 , n1947 );
xor ( n1958 , n1957 , n1950 );
and ( n1959 , n1675 , n1807 );
and ( n1960 , n1655 , n1805 );
nor ( n1961 , n1959 , n1960 );
xnor ( n1962 , n1961 , n1756 );
and ( n1963 , n1817 , n1646 );
and ( n1964 , n1799 , n1644 );
nor ( n1965 , n1963 , n1964 );
xnor ( n1966 , n1965 , n1651 );
and ( n1967 , n1962 , n1966 );
and ( n1968 , n1935 , n1663 );
and ( n1969 , n1849 , n1661 );
nor ( n1970 , n1968 , n1969 );
xnor ( n1971 , n1970 , n1671 );
and ( n1972 , n1966 , n1971 );
and ( n1973 , n1962 , n1971 );
or ( n1974 , n1967 , n1972 , n1973 );
buf ( n1975 , n1165 );
buf ( n1976 , n1975 );
buf ( n1977 , n1166 );
buf ( n1978 , n1977 );
and ( n1979 , n1976 , n1978 );
not ( n1980 , n1979 );
and ( n1981 , n1866 , n1980 );
not ( n1982 , n1981 );
and ( n1983 , n1666 , n1901 );
and ( n1984 , n1636 , n1899 );
nor ( n1985 , n1983 , n1984 );
xnor ( n1986 , n1985 , n1869 );
and ( n1987 , n1982 , n1986 );
and ( n1988 , n1720 , n1728 );
and ( n1989 , n1705 , n1726 );
nor ( n1990 , n1988 , n1989 );
xnor ( n1991 , n1990 , n1697 );
and ( n1992 , n1986 , n1991 );
and ( n1993 , n1982 , n1991 );
or ( n1994 , n1987 , n1992 , n1993 );
and ( n1995 , n1974 , n1994 );
xor ( n1996 , n1904 , n1908 );
xor ( n1997 , n1996 , n1913 );
and ( n1998 , n1994 , n1997 );
and ( n1999 , n1974 , n1997 );
or ( n2000 , n1995 , n1998 , n1999 );
and ( n2001 , n1655 , n1901 );
and ( n2002 , n1666 , n1899 );
nor ( n2003 , n2001 , n2002 );
xnor ( n2004 , n2003 , n1869 );
and ( n2005 , n1799 , n1728 );
and ( n2006 , n1720 , n1726 );
nor ( n2007 , n2005 , n2006 );
xnor ( n2008 , n2007 , n1697 );
and ( n2009 , n2004 , n2008 );
and ( n2010 , n1849 , n1646 );
and ( n2011 , n1817 , n1644 );
nor ( n2012 , n2010 , n2011 );
xnor ( n2013 , n2012 , n1651 );
and ( n2014 , n2008 , n2013 );
and ( n2015 , n2004 , n2013 );
or ( n2016 , n2009 , n2014 , n2015 );
xor ( n2017 , n1866 , n1976 );
xor ( n2018 , n1976 , n1978 );
not ( n2019 , n2018 );
and ( n2020 , n2017 , n2019 );
and ( n2021 , n1636 , n2020 );
not ( n2022 , n2021 );
xnor ( n2023 , n2022 , n1981 );
buf ( n2024 , n2023 );
and ( n2025 , n2016 , n2024 );
buf ( n2026 , n1132 );
buf ( n2027 , n2026 );
and ( n2028 , n2027 , n1657 );
and ( n2029 , n2024 , n2028 );
and ( n2030 , n2016 , n2028 );
or ( n2031 , n2025 , n2029 , n2030 );
and ( n2032 , n1705 , n1807 );
and ( n2033 , n1675 , n1805 );
nor ( n2034 , n2032 , n2033 );
xnor ( n2035 , n2034 , n1756 );
and ( n2036 , n2027 , n1663 );
and ( n2037 , n1935 , n1661 );
nor ( n2038 , n2036 , n2037 );
xnor ( n2039 , n2038 , n1671 );
and ( n2040 , n2035 , n2039 );
buf ( n2041 , n1133 );
buf ( n2042 , n2041 );
and ( n2043 , n2042 , n1657 );
and ( n2044 , n2039 , n2043 );
and ( n2045 , n2035 , n2043 );
or ( n2046 , n2040 , n2044 , n2045 );
xor ( n2047 , n1962 , n1966 );
xor ( n2048 , n2047 , n1971 );
and ( n2049 , n2046 , n2048 );
xor ( n2050 , n1982 , n1986 );
xor ( n2051 , n2050 , n1991 );
and ( n2052 , n2048 , n2051 );
and ( n2053 , n2046 , n2051 );
or ( n2054 , n2049 , n2052 , n2053 );
and ( n2055 , n2031 , n2054 );
xor ( n2056 , n1928 , n1932 );
xor ( n2057 , n2056 , n1936 );
and ( n2058 , n2054 , n2057 );
and ( n2059 , n2031 , n2057 );
or ( n2060 , n2055 , n2058 , n2059 );
and ( n2061 , n2000 , n2060 );
xor ( n2062 , n1939 , n1941 );
xor ( n2063 , n2062 , n1944 );
and ( n2064 , n2060 , n2063 );
and ( n2065 , n2000 , n2063 );
or ( n2066 , n2061 , n2064 , n2065 );
and ( n2067 , n1958 , n2066 );
xor ( n2068 , n2000 , n2060 );
xor ( n2069 , n2068 , n2063 );
and ( n2070 , n1675 , n1901 );
and ( n2071 , n1655 , n1899 );
nor ( n2072 , n2070 , n2071 );
xnor ( n2073 , n2072 , n1869 );
and ( n2074 , n1817 , n1728 );
and ( n2075 , n1799 , n1726 );
nor ( n2076 , n2074 , n2075 );
xnor ( n2077 , n2076 , n1697 );
and ( n2078 , n2073 , n2077 );
buf ( n2079 , n1134 );
buf ( n2080 , n2079 );
and ( n2081 , n2080 , n1657 );
and ( n2082 , n2077 , n2081 );
and ( n2083 , n2073 , n2081 );
or ( n2084 , n2078 , n2082 , n2083 );
buf ( n2085 , n1167 );
buf ( n2086 , n2085 );
buf ( n2087 , n1168 );
buf ( n2088 , n2087 );
and ( n2089 , n2086 , n2088 );
not ( n2090 , n2089 );
and ( n2091 , n1978 , n2090 );
not ( n2092 , n2091 );
and ( n2093 , n1666 , n2020 );
and ( n2094 , n1636 , n2018 );
nor ( n2095 , n2093 , n2094 );
xnor ( n2096 , n2095 , n1981 );
and ( n2097 , n2092 , n2096 );
and ( n2098 , n1720 , n1807 );
and ( n2099 , n1705 , n1805 );
nor ( n2100 , n2098 , n2099 );
xnor ( n2101 , n2100 , n1756 );
and ( n2102 , n2096 , n2101 );
and ( n2103 , n2092 , n2101 );
or ( n2104 , n2097 , n2102 , n2103 );
and ( n2105 , n2084 , n2104 );
not ( n2106 , n2023 );
and ( n2107 , n2104 , n2106 );
and ( n2108 , n2084 , n2106 );
or ( n2109 , n2105 , n2107 , n2108 );
xor ( n2110 , n1978 , n2086 );
xor ( n2111 , n2086 , n2088 );
not ( n2112 , n2111 );
and ( n2113 , n2110 , n2112 );
and ( n2114 , n1636 , n2113 );
not ( n2115 , n2114 );
xnor ( n2116 , n2115 , n2091 );
buf ( n2117 , n2116 );
and ( n2118 , n1935 , n1646 );
and ( n2119 , n1849 , n1644 );
nor ( n2120 , n2118 , n2119 );
xnor ( n2121 , n2120 , n1651 );
and ( n2122 , n2117 , n2121 );
and ( n2123 , n2042 , n1663 );
and ( n2124 , n2027 , n1661 );
nor ( n2125 , n2123 , n2124 );
xnor ( n2126 , n2125 , n1671 );
and ( n2127 , n2121 , n2126 );
and ( n2128 , n2117 , n2126 );
or ( n2129 , n2122 , n2127 , n2128 );
xor ( n2130 , n2035 , n2039 );
xor ( n2131 , n2130 , n2043 );
and ( n2132 , n2129 , n2131 );
xor ( n2133 , n2004 , n2008 );
xor ( n2134 , n2133 , n2013 );
and ( n2135 , n2131 , n2134 );
and ( n2136 , n2129 , n2134 );
or ( n2137 , n2132 , n2135 , n2136 );
and ( n2138 , n2109 , n2137 );
xor ( n2139 , n2016 , n2024 );
xor ( n2140 , n2139 , n2028 );
and ( n2141 , n2137 , n2140 );
and ( n2142 , n2109 , n2140 );
or ( n2143 , n2138 , n2141 , n2142 );
xor ( n2144 , n1974 , n1994 );
xor ( n2145 , n2144 , n1997 );
and ( n2146 , n2143 , n2145 );
xor ( n2147 , n2031 , n2054 );
xor ( n2148 , n2147 , n2057 );
and ( n2149 , n2145 , n2148 );
and ( n2150 , n2143 , n2148 );
or ( n2151 , n2146 , n2149 , n2150 );
and ( n2152 , n2069 , n2151 );
xor ( n2153 , n2143 , n2145 );
xor ( n2154 , n2153 , n2148 );
and ( n2155 , n1705 , n1901 );
and ( n2156 , n1675 , n1899 );
nor ( n2157 , n2155 , n2156 );
xnor ( n2158 , n2157 , n1869 );
and ( n2159 , n1849 , n1728 );
and ( n2160 , n1817 , n1726 );
nor ( n2161 , n2159 , n2160 );
xnor ( n2162 , n2161 , n1697 );
and ( n2163 , n2158 , n2162 );
and ( n2164 , n2027 , n1646 );
and ( n2165 , n1935 , n1644 );
nor ( n2166 , n2164 , n2165 );
xnor ( n2167 , n2166 , n1651 );
and ( n2168 , n2162 , n2167 );
and ( n2169 , n2158 , n2167 );
or ( n2170 , n2163 , n2168 , n2169 );
and ( n2171 , n1655 , n2020 );
and ( n2172 , n1666 , n2018 );
nor ( n2173 , n2171 , n2172 );
xnor ( n2174 , n2173 , n1981 );
and ( n2175 , n1799 , n1807 );
and ( n2176 , n1720 , n1805 );
nor ( n2177 , n2175 , n2176 );
xnor ( n2178 , n2177 , n1756 );
and ( n2179 , n2174 , n2178 );
buf ( n2180 , n1135 );
buf ( n2181 , n2180 );
and ( n2182 , n2181 , n1657 );
and ( n2183 , n2178 , n2182 );
and ( n2184 , n2174 , n2182 );
or ( n2185 , n2179 , n2183 , n2184 );
and ( n2186 , n2170 , n2185 );
xor ( n2187 , n2092 , n2096 );
xor ( n2188 , n2187 , n2101 );
and ( n2189 , n2185 , n2188 );
and ( n2190 , n2170 , n2188 );
or ( n2191 , n2186 , n2189 , n2190 );
xor ( n2192 , n2084 , n2104 );
xor ( n2193 , n2192 , n2106 );
and ( n2194 , n2191 , n2193 );
xor ( n2195 , n2129 , n2131 );
xor ( n2196 , n2195 , n2134 );
and ( n2197 , n2193 , n2196 );
and ( n2198 , n2191 , n2196 );
or ( n2199 , n2194 , n2197 , n2198 );
xor ( n2200 , n2046 , n2048 );
xor ( n2201 , n2200 , n2051 );
and ( n2202 , n2199 , n2201 );
xor ( n2203 , n2109 , n2137 );
xor ( n2204 , n2203 , n2140 );
and ( n2205 , n2201 , n2204 );
and ( n2206 , n2199 , n2204 );
or ( n2207 , n2202 , n2205 , n2206 );
and ( n2208 , n2154 , n2207 );
xor ( n2209 , n2199 , n2201 );
xor ( n2210 , n2209 , n2204 );
buf ( n2211 , n1169 );
buf ( n2212 , n2211 );
buf ( n2213 , n1170 );
buf ( n2214 , n2213 );
and ( n2215 , n2212 , n2214 );
not ( n2216 , n2215 );
and ( n2217 , n2088 , n2216 );
not ( n2218 , n2217 );
and ( n2219 , n1666 , n2113 );
and ( n2220 , n1636 , n2111 );
nor ( n2221 , n2219 , n2220 );
xnor ( n2222 , n2221 , n2091 );
and ( n2223 , n2218 , n2222 );
and ( n2224 , n1720 , n1901 );
and ( n2225 , n1705 , n1899 );
nor ( n2226 , n2224 , n2225 );
xnor ( n2227 , n2226 , n1869 );
and ( n2228 , n2222 , n2227 );
and ( n2229 , n2218 , n2227 );
or ( n2230 , n2223 , n2228 , n2229 );
not ( n2231 , n2116 );
and ( n2232 , n2230 , n2231 );
and ( n2233 , n2080 , n1663 );
and ( n2234 , n2042 , n1661 );
nor ( n2235 , n2233 , n2234 );
xnor ( n2236 , n2235 , n1671 );
and ( n2237 , n2231 , n2236 );
and ( n2238 , n2230 , n2236 );
or ( n2239 , n2232 , n2237 , n2238 );
xor ( n2240 , n2073 , n2077 );
xor ( n2241 , n2240 , n2081 );
and ( n2242 , n2239 , n2241 );
xor ( n2243 , n2117 , n2121 );
xor ( n2244 , n2243 , n2126 );
and ( n2245 , n2241 , n2244 );
and ( n2246 , n2239 , n2244 );
or ( n2247 , n2242 , n2245 , n2246 );
and ( n2248 , n1817 , n1807 );
and ( n2249 , n1799 , n1805 );
nor ( n2250 , n2248 , n2249 );
xnor ( n2251 , n2250 , n1756 );
and ( n2252 , n2181 , n1663 );
and ( n2253 , n2080 , n1661 );
nor ( n2254 , n2252 , n2253 );
xnor ( n2255 , n2254 , n1671 );
and ( n2256 , n2251 , n2255 );
buf ( n2257 , n1136 );
buf ( n2258 , n2257 );
and ( n2259 , n2258 , n1657 );
and ( n2260 , n2255 , n2259 );
and ( n2261 , n2251 , n2259 );
or ( n2262 , n2256 , n2260 , n2261 );
and ( n2263 , n1675 , n2020 );
and ( n2264 , n1655 , n2018 );
nor ( n2265 , n2263 , n2264 );
xnor ( n2266 , n2265 , n1981 );
and ( n2267 , n1935 , n1728 );
and ( n2268 , n1849 , n1726 );
nor ( n2269 , n2267 , n2268 );
xnor ( n2270 , n2269 , n1697 );
and ( n2271 , n2266 , n2270 );
and ( n2272 , n2042 , n1646 );
and ( n2273 , n2027 , n1644 );
nor ( n2274 , n2272 , n2273 );
xnor ( n2275 , n2274 , n1651 );
and ( n2276 , n2270 , n2275 );
and ( n2277 , n2266 , n2275 );
or ( n2278 , n2271 , n2276 , n2277 );
and ( n2279 , n2262 , n2278 );
xor ( n2280 , n2158 , n2162 );
xor ( n2281 , n2280 , n2167 );
and ( n2282 , n2278 , n2281 );
and ( n2283 , n2262 , n2281 );
or ( n2284 , n2279 , n2282 , n2283 );
and ( n2285 , n1799 , n1901 );
and ( n2286 , n1720 , n1899 );
nor ( n2287 , n2285 , n2286 );
xnor ( n2288 , n2287 , n1869 );
and ( n2289 , n2258 , n1663 );
and ( n2290 , n2181 , n1661 );
nor ( n2291 , n2289 , n2290 );
xnor ( n2292 , n2291 , n1671 );
and ( n2293 , n2288 , n2292 );
buf ( n2294 , n1137 );
buf ( n2295 , n2294 );
and ( n2296 , n2295 , n1657 );
and ( n2297 , n2292 , n2296 );
and ( n2298 , n2288 , n2296 );
or ( n2299 , n2293 , n2297 , n2298 );
and ( n2300 , n1655 , n2113 );
and ( n2301 , n1666 , n2111 );
nor ( n2302 , n2300 , n2301 );
xnor ( n2303 , n2302 , n2091 );
and ( n2304 , n1705 , n2020 );
and ( n2305 , n1675 , n2018 );
nor ( n2306 , n2304 , n2305 );
xnor ( n2307 , n2306 , n1981 );
and ( n2308 , n2303 , n2307 );
and ( n2309 , n1849 , n1807 );
and ( n2310 , n1817 , n1805 );
nor ( n2311 , n2309 , n2310 );
xnor ( n2312 , n2311 , n1756 );
and ( n2313 , n2307 , n2312 );
and ( n2314 , n2303 , n2312 );
or ( n2315 , n2308 , n2313 , n2314 );
and ( n2316 , n2299 , n2315 );
xor ( n2317 , n2088 , n2212 );
xor ( n2318 , n2212 , n2214 );
not ( n2319 , n2318 );
and ( n2320 , n2317 , n2319 );
and ( n2321 , n1636 , n2320 );
not ( n2322 , n2321 );
xnor ( n2323 , n2322 , n2217 );
buf ( n2324 , n2323 );
and ( n2325 , n2315 , n2324 );
and ( n2326 , n2299 , n2324 );
or ( n2327 , n2316 , n2325 , n2326 );
xor ( n2328 , n2174 , n2178 );
xor ( n2329 , n2328 , n2182 );
and ( n2330 , n2327 , n2329 );
xor ( n2331 , n2230 , n2231 );
xor ( n2332 , n2331 , n2236 );
and ( n2333 , n2329 , n2332 );
and ( n2334 , n2327 , n2332 );
or ( n2335 , n2330 , n2333 , n2334 );
and ( n2336 , n2284 , n2335 );
xor ( n2337 , n2170 , n2185 );
xor ( n2338 , n2337 , n2188 );
and ( n2339 , n2335 , n2338 );
and ( n2340 , n2284 , n2338 );
or ( n2341 , n2336 , n2339 , n2340 );
and ( n2342 , n2247 , n2341 );
xor ( n2343 , n2191 , n2193 );
xor ( n2344 , n2343 , n2196 );
and ( n2345 , n2341 , n2344 );
and ( n2346 , n2247 , n2344 );
or ( n2347 , n2342 , n2345 , n2346 );
and ( n2348 , n2210 , n2347 );
xor ( n2349 , n2251 , n2255 );
xor ( n2350 , n2349 , n2259 );
xor ( n2351 , n2266 , n2270 );
xor ( n2352 , n2351 , n2275 );
and ( n2353 , n2350 , n2352 );
xor ( n2354 , n2218 , n2222 );
xor ( n2355 , n2354 , n2227 );
and ( n2356 , n2352 , n2355 );
and ( n2357 , n2350 , n2355 );
or ( n2358 , n2353 , n2356 , n2357 );
xor ( n2359 , n2262 , n2278 );
xor ( n2360 , n2359 , n2281 );
and ( n2361 , n2358 , n2360 );
xor ( n2362 , n2327 , n2329 );
xor ( n2363 , n2362 , n2332 );
and ( n2364 , n2360 , n2363 );
and ( n2365 , n2358 , n2363 );
or ( n2366 , n2361 , n2364 , n2365 );
xor ( n2367 , n2239 , n2241 );
xor ( n2368 , n2367 , n2244 );
and ( n2369 , n2366 , n2368 );
xor ( n2370 , n2284 , n2335 );
xor ( n2371 , n2370 , n2338 );
and ( n2372 , n2368 , n2371 );
and ( n2373 , n2366 , n2371 );
or ( n2374 , n2369 , n2372 , n2373 );
xor ( n2375 , n2247 , n2341 );
xor ( n2376 , n2375 , n2344 );
and ( n2377 , n2374 , n2376 );
xor ( n2378 , n2366 , n2368 );
xor ( n2379 , n2378 , n2371 );
and ( n2380 , n1675 , n2113 );
and ( n2381 , n1655 , n2111 );
nor ( n2382 , n2380 , n2381 );
xnor ( n2383 , n2382 , n2091 );
and ( n2384 , n1935 , n1807 );
and ( n2385 , n1849 , n1805 );
nor ( n2386 , n2384 , n2385 );
xnor ( n2387 , n2386 , n1756 );
and ( n2388 , n2383 , n2387 );
buf ( n2389 , n1138 );
buf ( n2390 , n2389 );
and ( n2391 , n2390 , n1657 );
and ( n2392 , n2387 , n2391 );
and ( n2393 , n2383 , n2391 );
or ( n2394 , n2388 , n2392 , n2393 );
and ( n2395 , n1817 , n1901 );
and ( n2396 , n1799 , n1899 );
nor ( n2397 , n2395 , n2396 );
xnor ( n2398 , n2397 , n1869 );
and ( n2399 , n2181 , n1646 );
and ( n2400 , n2080 , n1644 );
nor ( n2401 , n2399 , n2400 );
xnor ( n2402 , n2401 , n1651 );
and ( n2403 , n2398 , n2402 );
and ( n2404 , n2295 , n1663 );
and ( n2405 , n2258 , n1661 );
nor ( n2406 , n2404 , n2405 );
xnor ( n2407 , n2406 , n1671 );
and ( n2408 , n2402 , n2407 );
and ( n2409 , n2398 , n2407 );
or ( n2410 , n2403 , n2408 , n2409 );
and ( n2411 , n2394 , n2410 );
buf ( n2412 , n1171 );
buf ( n2413 , n2412 );
buf ( n2414 , n1172 );
buf ( n2415 , n2414 );
and ( n2416 , n2413 , n2415 );
not ( n2417 , n2416 );
and ( n2418 , n2214 , n2417 );
not ( n2419 , n2418 );
and ( n2420 , n1666 , n2320 );
and ( n2421 , n1636 , n2318 );
nor ( n2422 , n2420 , n2421 );
xnor ( n2423 , n2422 , n2217 );
and ( n2424 , n2419 , n2423 );
and ( n2425 , n1720 , n2020 );
and ( n2426 , n1705 , n2018 );
nor ( n2427 , n2425 , n2426 );
xnor ( n2428 , n2427 , n1981 );
and ( n2429 , n2423 , n2428 );
and ( n2430 , n2419 , n2428 );
or ( n2431 , n2424 , n2429 , n2430 );
and ( n2432 , n2410 , n2431 );
and ( n2433 , n2394 , n2431 );
or ( n2434 , n2411 , n2432 , n2433 );
not ( n2435 , n2323 );
and ( n2436 , n2027 , n1728 );
and ( n2437 , n1935 , n1726 );
nor ( n2438 , n2436 , n2437 );
xnor ( n2439 , n2438 , n1697 );
and ( n2440 , n2435 , n2439 );
and ( n2441 , n2080 , n1646 );
and ( n2442 , n2042 , n1644 );
nor ( n2443 , n2441 , n2442 );
xnor ( n2444 , n2443 , n1651 );
and ( n2445 , n2439 , n2444 );
and ( n2446 , n2435 , n2444 );
or ( n2447 , n2440 , n2445 , n2446 );
and ( n2448 , n2434 , n2447 );
xor ( n2449 , n2299 , n2315 );
xor ( n2450 , n2449 , n2324 );
and ( n2451 , n2447 , n2450 );
and ( n2452 , n2434 , n2450 );
or ( n2453 , n2448 , n2451 , n2452 );
xor ( n2454 , n2288 , n2292 );
xor ( n2455 , n2454 , n2296 );
xor ( n2456 , n2303 , n2307 );
xor ( n2457 , n2456 , n2312 );
and ( n2458 , n2455 , n2457 );
xor ( n2459 , n2435 , n2439 );
xor ( n2460 , n2459 , n2444 );
and ( n2461 , n2457 , n2460 );
and ( n2462 , n2455 , n2460 );
or ( n2463 , n2458 , n2461 , n2462 );
and ( n2464 , n1799 , n2020 );
and ( n2465 , n1720 , n2018 );
nor ( n2466 , n2464 , n2465 );
xnor ( n2467 , n2466 , n1981 );
and ( n2468 , n2258 , n1646 );
and ( n2469 , n2181 , n1644 );
nor ( n2470 , n2468 , n2469 );
xnor ( n2471 , n2470 , n1651 );
and ( n2472 , n2467 , n2471 );
and ( n2473 , n2390 , n1663 );
and ( n2474 , n2295 , n1661 );
nor ( n2475 , n2473 , n2474 );
xnor ( n2476 , n2475 , n1671 );
and ( n2477 , n2471 , n2476 );
and ( n2478 , n2467 , n2476 );
or ( n2479 , n2472 , n2477 , n2478 );
xor ( n2480 , n2214 , n2413 );
xor ( n2481 , n2413 , n2415 );
not ( n2482 , n2481 );
and ( n2483 , n2480 , n2482 );
and ( n2484 , n1636 , n2483 );
not ( n2485 , n2484 );
xnor ( n2486 , n2485 , n2418 );
buf ( n2487 , n2486 );
and ( n2488 , n2479 , n2487 );
and ( n2489 , n2042 , n1728 );
and ( n2490 , n2027 , n1726 );
nor ( n2491 , n2489 , n2490 );
xnor ( n2492 , n2491 , n1697 );
and ( n2493 , n2487 , n2492 );
and ( n2494 , n2479 , n2492 );
or ( n2495 , n2488 , n2493 , n2494 );
and ( n2496 , n1655 , n2320 );
and ( n2497 , n1666 , n2318 );
nor ( n2498 , n2496 , n2497 );
xnor ( n2499 , n2498 , n2217 );
and ( n2500 , n1849 , n1901 );
and ( n2501 , n1817 , n1899 );
nor ( n2502 , n2500 , n2501 );
xnor ( n2503 , n2502 , n1869 );
and ( n2504 , n2499 , n2503 );
buf ( n2505 , n1139 );
buf ( n2506 , n2505 );
and ( n2507 , n2506 , n1657 );
and ( n2508 , n2503 , n2507 );
and ( n2509 , n2499 , n2507 );
or ( n2510 , n2504 , n2508 , n2509 );
and ( n2511 , n1705 , n2113 );
and ( n2512 , n1675 , n2111 );
nor ( n2513 , n2511 , n2512 );
xnor ( n2514 , n2513 , n2091 );
and ( n2515 , n2027 , n1807 );
and ( n2516 , n1935 , n1805 );
nor ( n2517 , n2515 , n2516 );
xnor ( n2518 , n2517 , n1756 );
and ( n2519 , n2514 , n2518 );
and ( n2520 , n2080 , n1728 );
and ( n2521 , n2042 , n1726 );
nor ( n2522 , n2520 , n2521 );
xnor ( n2523 , n2522 , n1697 );
and ( n2524 , n2518 , n2523 );
and ( n2525 , n2514 , n2523 );
or ( n2526 , n2519 , n2524 , n2525 );
and ( n2527 , n2510 , n2526 );
xor ( n2528 , n2383 , n2387 );
xor ( n2529 , n2528 , n2391 );
and ( n2530 , n2526 , n2529 );
and ( n2531 , n2510 , n2529 );
or ( n2532 , n2527 , n2530 , n2531 );
and ( n2533 , n2495 , n2532 );
xor ( n2534 , n2394 , n2410 );
xor ( n2535 , n2534 , n2431 );
and ( n2536 , n2532 , n2535 );
and ( n2537 , n2495 , n2535 );
or ( n2538 , n2533 , n2536 , n2537 );
and ( n2539 , n2463 , n2538 );
xor ( n2540 , n2350 , n2352 );
xor ( n2541 , n2540 , n2355 );
and ( n2542 , n2538 , n2541 );
and ( n2543 , n2463 , n2541 );
or ( n2544 , n2539 , n2542 , n2543 );
and ( n2545 , n2453 , n2544 );
xor ( n2546 , n2358 , n2360 );
xor ( n2547 , n2546 , n2363 );
and ( n2548 , n2544 , n2547 );
and ( n2549 , n2453 , n2547 );
or ( n2550 , n2545 , n2548 , n2549 );
and ( n2551 , n2379 , n2550 );
xor ( n2552 , n2453 , n2544 );
xor ( n2553 , n2552 , n2547 );
xor ( n2554 , n2398 , n2402 );
xor ( n2555 , n2554 , n2407 );
xor ( n2556 , n2419 , n2423 );
xor ( n2557 , n2556 , n2428 );
and ( n2558 , n2555 , n2557 );
xor ( n2559 , n2479 , n2487 );
xor ( n2560 , n2559 , n2492 );
and ( n2561 , n2557 , n2560 );
and ( n2562 , n2555 , n2560 );
or ( n2563 , n2558 , n2561 , n2562 );
buf ( n2564 , n1173 );
buf ( n2565 , n2564 );
buf ( n2566 , n1174 );
buf ( n2567 , n2566 );
and ( n2568 , n2565 , n2567 );
not ( n2569 , n2568 );
and ( n2570 , n2415 , n2569 );
not ( n2571 , n2570 );
and ( n2572 , n1666 , n2483 );
and ( n2573 , n1636 , n2481 );
nor ( n2574 , n2572 , n2573 );
xnor ( n2575 , n2574 , n2418 );
and ( n2576 , n2571 , n2575 );
and ( n2577 , n1720 , n2113 );
and ( n2578 , n1705 , n2111 );
nor ( n2579 , n2577 , n2578 );
xnor ( n2580 , n2579 , n2091 );
and ( n2581 , n2575 , n2580 );
and ( n2582 , n2571 , n2580 );
or ( n2583 , n2576 , n2581 , n2582 );
and ( n2584 , n1817 , n2020 );
and ( n2585 , n1799 , n2018 );
nor ( n2586 , n2584 , n2585 );
xnor ( n2587 , n2586 , n1981 );
and ( n2588 , n2181 , n1728 );
and ( n2589 , n2080 , n1726 );
nor ( n2590 , n2588 , n2589 );
xnor ( n2591 , n2590 , n1697 );
and ( n2592 , n2587 , n2591 );
and ( n2593 , n2295 , n1646 );
and ( n2594 , n2258 , n1644 );
nor ( n2595 , n2593 , n2594 );
xnor ( n2596 , n2595 , n1651 );
and ( n2597 , n2591 , n2596 );
and ( n2598 , n2587 , n2596 );
or ( n2599 , n2592 , n2597 , n2598 );
and ( n2600 , n2583 , n2599 );
not ( n2601 , n2486 );
and ( n2602 , n2599 , n2601 );
and ( n2603 , n2583 , n2601 );
or ( n2604 , n2600 , n2602 , n2603 );
and ( n2605 , n1675 , n2320 );
and ( n2606 , n1655 , n2318 );
nor ( n2607 , n2605 , n2606 );
xnor ( n2608 , n2607 , n2217 );
and ( n2609 , n2506 , n1663 );
and ( n2610 , n2390 , n1661 );
nor ( n2611 , n2609 , n2610 );
xnor ( n2612 , n2611 , n1671 );
and ( n2613 , n2608 , n2612 );
buf ( n2614 , n1140 );
buf ( n2615 , n2614 );
and ( n2616 , n2615 , n1657 );
and ( n2617 , n2612 , n2616 );
and ( n2618 , n2608 , n2616 );
or ( n2619 , n2613 , n2617 , n2618 );
xor ( n2620 , n2499 , n2503 );
xor ( n2621 , n2620 , n2507 );
and ( n2622 , n2619 , n2621 );
xor ( n2623 , n2467 , n2471 );
xor ( n2624 , n2623 , n2476 );
and ( n2625 , n2621 , n2624 );
and ( n2626 , n2619 , n2624 );
or ( n2627 , n2622 , n2625 , n2626 );
and ( n2628 , n2604 , n2627 );
xor ( n2629 , n2510 , n2526 );
xor ( n2630 , n2629 , n2529 );
and ( n2631 , n2627 , n2630 );
and ( n2632 , n2604 , n2630 );
or ( n2633 , n2628 , n2631 , n2632 );
and ( n2634 , n2563 , n2633 );
xor ( n2635 , n2455 , n2457 );
xor ( n2636 , n2635 , n2460 );
and ( n2637 , n2633 , n2636 );
and ( n2638 , n2563 , n2636 );
or ( n2639 , n2634 , n2637 , n2638 );
xor ( n2640 , n2434 , n2447 );
xor ( n2641 , n2640 , n2450 );
and ( n2642 , n2639 , n2641 );
xor ( n2643 , n2463 , n2538 );
xor ( n2644 , n2643 , n2541 );
and ( n2645 , n2641 , n2644 );
and ( n2646 , n2639 , n2644 );
or ( n2647 , n2642 , n2645 , n2646 );
and ( n2648 , n2553 , n2647 );
xor ( n2649 , n2639 , n2641 );
xor ( n2650 , n2649 , n2644 );
xor ( n2651 , n2415 , n2565 );
xor ( n2652 , n2565 , n2567 );
not ( n2653 , n2652 );
and ( n2654 , n2651 , n2653 );
and ( n2655 , n1636 , n2654 );
not ( n2656 , n2655 );
xnor ( n2657 , n2656 , n2570 );
and ( n2658 , n1705 , n2320 );
and ( n2659 , n1675 , n2318 );
nor ( n2660 , n2658 , n2659 );
xnor ( n2661 , n2660 , n2217 );
and ( n2662 , n2657 , n2661 );
and ( n2663 , n2027 , n1901 );
and ( n2664 , n1935 , n1899 );
nor ( n2665 , n2663 , n2664 );
xnor ( n2666 , n2665 , n1869 );
and ( n2667 , n2661 , n2666 );
and ( n2668 , n2657 , n2666 );
or ( n2669 , n2662 , n2667 , n2668 );
and ( n2670 , n1799 , n2113 );
and ( n2671 , n1720 , n2111 );
nor ( n2672 , n2670 , n2671 );
xnor ( n2673 , n2672 , n2091 );
and ( n2674 , n2258 , n1728 );
and ( n2675 , n2181 , n1726 );
nor ( n2676 , n2674 , n2675 );
xnor ( n2677 , n2676 , n1697 );
and ( n2678 , n2673 , n2677 );
and ( n2679 , n2390 , n1646 );
and ( n2680 , n2295 , n1644 );
nor ( n2681 , n2679 , n2680 );
xnor ( n2682 , n2681 , n1651 );
and ( n2683 , n2677 , n2682 );
and ( n2684 , n2673 , n2682 );
or ( n2685 , n2678 , n2683 , n2684 );
and ( n2686 , n2669 , n2685 );
and ( n2687 , n1849 , n2020 );
and ( n2688 , n1817 , n2018 );
nor ( n2689 , n2687 , n2688 );
xnor ( n2690 , n2689 , n1981 );
and ( n2691 , n2615 , n1663 );
and ( n2692 , n2506 , n1661 );
nor ( n2693 , n2691 , n2692 );
xnor ( n2694 , n2693 , n1671 );
and ( n2695 , n2690 , n2694 );
buf ( n2696 , n1141 );
buf ( n2697 , n2696 );
and ( n2698 , n2697 , n1657 );
and ( n2699 , n2694 , n2698 );
and ( n2700 , n2690 , n2698 );
or ( n2701 , n2695 , n2699 , n2700 );
and ( n2702 , n2685 , n2701 );
and ( n2703 , n2669 , n2701 );
or ( n2704 , n2686 , n2702 , n2703 );
and ( n2705 , n1655 , n2483 );
and ( n2706 , n1666 , n2481 );
nor ( n2707 , n2705 , n2706 );
xnor ( n2708 , n2707 , n2418 );
buf ( n2709 , n2708 );
and ( n2710 , n1935 , n1901 );
and ( n2711 , n1849 , n1899 );
nor ( n2712 , n2710 , n2711 );
xnor ( n2713 , n2712 , n1869 );
and ( n2714 , n2709 , n2713 );
and ( n2715 , n2042 , n1807 );
and ( n2716 , n2027 , n1805 );
nor ( n2717 , n2715 , n2716 );
xnor ( n2718 , n2717 , n1756 );
and ( n2719 , n2713 , n2718 );
and ( n2720 , n2709 , n2718 );
or ( n2721 , n2714 , n2719 , n2720 );
and ( n2722 , n2704 , n2721 );
xor ( n2723 , n2514 , n2518 );
xor ( n2724 , n2723 , n2523 );
and ( n2725 , n2721 , n2724 );
and ( n2726 , n2704 , n2724 );
or ( n2727 , n2722 , n2725 , n2726 );
xor ( n2728 , n2571 , n2575 );
xor ( n2729 , n2728 , n2580 );
xor ( n2730 , n2587 , n2591 );
xor ( n2731 , n2730 , n2596 );
and ( n2732 , n2729 , n2731 );
xor ( n2733 , n2608 , n2612 );
xor ( n2734 , n2733 , n2616 );
and ( n2735 , n2731 , n2734 );
and ( n2736 , n2729 , n2734 );
or ( n2737 , n2732 , n2735 , n2736 );
xor ( n2738 , n2583 , n2599 );
xor ( n2739 , n2738 , n2601 );
and ( n2740 , n2737 , n2739 );
xor ( n2741 , n2619 , n2621 );
xor ( n2742 , n2741 , n2624 );
and ( n2743 , n2739 , n2742 );
and ( n2744 , n2737 , n2742 );
or ( n2745 , n2740 , n2743 , n2744 );
and ( n2746 , n2727 , n2745 );
xor ( n2747 , n2555 , n2557 );
xor ( n2748 , n2747 , n2560 );
and ( n2749 , n2745 , n2748 );
and ( n2750 , n2727 , n2748 );
or ( n2751 , n2746 , n2749 , n2750 );
xor ( n2752 , n2495 , n2532 );
xor ( n2753 , n2752 , n2535 );
and ( n2754 , n2751 , n2753 );
xor ( n2755 , n2563 , n2633 );
xor ( n2756 , n2755 , n2636 );
and ( n2757 , n2753 , n2756 );
and ( n2758 , n2751 , n2756 );
or ( n2759 , n2754 , n2757 , n2758 );
and ( n2760 , n2650 , n2759 );
xor ( n2761 , n2751 , n2753 );
xor ( n2762 , n2761 , n2756 );
and ( n2763 , n1935 , n2020 );
and ( n2764 , n1849 , n2018 );
nor ( n2765 , n2763 , n2764 );
xnor ( n2766 , n2765 , n1981 );
and ( n2767 , n2042 , n1901 );
and ( n2768 , n2027 , n1899 );
nor ( n2769 , n2767 , n2768 );
xnor ( n2770 , n2769 , n1869 );
and ( n2771 , n2766 , n2770 );
buf ( n2772 , n1142 );
buf ( n2773 , n2772 );
and ( n2774 , n2773 , n1657 );
and ( n2775 , n2770 , n2774 );
and ( n2776 , n2766 , n2774 );
or ( n2777 , n2771 , n2775 , n2776 );
and ( n2778 , n1817 , n2113 );
and ( n2779 , n1799 , n2111 );
nor ( n2780 , n2778 , n2779 );
xnor ( n2781 , n2780 , n2091 );
and ( n2782 , n2181 , n1807 );
and ( n2783 , n2080 , n1805 );
nor ( n2784 , n2782 , n2783 );
xnor ( n2785 , n2784 , n1756 );
and ( n2786 , n2781 , n2785 );
and ( n2787 , n2295 , n1728 );
and ( n2788 , n2258 , n1726 );
nor ( n2789 , n2787 , n2788 );
xnor ( n2790 , n2789 , n1697 );
and ( n2791 , n2785 , n2790 );
and ( n2792 , n2781 , n2790 );
or ( n2793 , n2786 , n2791 , n2792 );
and ( n2794 , n2777 , n2793 );
buf ( n2795 , n1175 );
buf ( n2796 , n2795 );
buf ( n2797 , n1176 );
buf ( n2798 , n2797 );
and ( n2799 , n2796 , n2798 );
not ( n2800 , n2799 );
and ( n2801 , n2567 , n2800 );
not ( n2802 , n2801 );
and ( n2803 , n1666 , n2654 );
and ( n2804 , n1636 , n2652 );
nor ( n2805 , n2803 , n2804 );
xnor ( n2806 , n2805 , n2570 );
and ( n2807 , n2802 , n2806 );
and ( n2808 , n1720 , n2320 );
and ( n2809 , n1705 , n2318 );
nor ( n2810 , n2808 , n2809 );
xnor ( n2811 , n2810 , n2217 );
and ( n2812 , n2806 , n2811 );
and ( n2813 , n2802 , n2811 );
or ( n2814 , n2807 , n2812 , n2813 );
and ( n2815 , n2793 , n2814 );
and ( n2816 , n2777 , n2814 );
or ( n2817 , n2794 , n2815 , n2816 );
and ( n2818 , n1675 , n2483 );
and ( n2819 , n1655 , n2481 );
nor ( n2820 , n2818 , n2819 );
xnor ( n2821 , n2820 , n2418 );
and ( n2822 , n2506 , n1646 );
and ( n2823 , n2390 , n1644 );
nor ( n2824 , n2822 , n2823 );
xnor ( n2825 , n2824 , n1651 );
and ( n2826 , n2821 , n2825 );
and ( n2827 , n2697 , n1663 );
and ( n2828 , n2615 , n1661 );
nor ( n2829 , n2827 , n2828 );
xnor ( n2830 , n2829 , n1671 );
and ( n2831 , n2825 , n2830 );
and ( n2832 , n2821 , n2830 );
or ( n2833 , n2826 , n2831 , n2832 );
not ( n2834 , n2708 );
and ( n2835 , n2833 , n2834 );
and ( n2836 , n2080 , n1807 );
and ( n2837 , n2042 , n1805 );
nor ( n2838 , n2836 , n2837 );
xnor ( n2839 , n2838 , n1756 );
and ( n2840 , n2834 , n2839 );
and ( n2841 , n2833 , n2839 );
or ( n2842 , n2835 , n2840 , n2841 );
and ( n2843 , n2817 , n2842 );
xor ( n2844 , n2709 , n2713 );
xor ( n2845 , n2844 , n2718 );
and ( n2846 , n2842 , n2845 );
and ( n2847 , n2817 , n2845 );
or ( n2848 , n2843 , n2846 , n2847 );
xor ( n2849 , n2657 , n2661 );
xor ( n2850 , n2849 , n2666 );
xor ( n2851 , n2673 , n2677 );
xor ( n2852 , n2851 , n2682 );
and ( n2853 , n2850 , n2852 );
xor ( n2854 , n2690 , n2694 );
xor ( n2855 , n2854 , n2698 );
and ( n2856 , n2852 , n2855 );
and ( n2857 , n2850 , n2855 );
or ( n2858 , n2853 , n2856 , n2857 );
xor ( n2859 , n2669 , n2685 );
xor ( n2860 , n2859 , n2701 );
and ( n2861 , n2858 , n2860 );
xor ( n2862 , n2729 , n2731 );
xor ( n2863 , n2862 , n2734 );
and ( n2864 , n2860 , n2863 );
and ( n2865 , n2858 , n2863 );
or ( n2866 , n2861 , n2864 , n2865 );
and ( n2867 , n2848 , n2866 );
xor ( n2868 , n2704 , n2721 );
xor ( n2869 , n2868 , n2724 );
and ( n2870 , n2866 , n2869 );
and ( n2871 , n2848 , n2869 );
or ( n2872 , n2867 , n2870 , n2871 );
xor ( n2873 , n2604 , n2627 );
xor ( n2874 , n2873 , n2630 );
and ( n2875 , n2872 , n2874 );
xor ( n2876 , n2727 , n2745 );
xor ( n2877 , n2876 , n2748 );
and ( n2878 , n2874 , n2877 );
and ( n2879 , n2872 , n2877 );
or ( n2880 , n2875 , n2878 , n2879 );
and ( n2881 , n2762 , n2880 );
xor ( n2882 , n2872 , n2874 );
xor ( n2883 , n2882 , n2877 );
xor ( n2884 , n2567 , n2796 );
xor ( n2885 , n2796 , n2798 );
not ( n2886 , n2885 );
and ( n2887 , n2884 , n2886 );
and ( n2888 , n1636 , n2887 );
not ( n2889 , n2888 );
xnor ( n2890 , n2889 , n2801 );
and ( n2891 , n1705 , n2483 );
and ( n2892 , n1675 , n2481 );
nor ( n2893 , n2891 , n2892 );
xnor ( n2894 , n2893 , n2418 );
and ( n2895 , n2890 , n2894 );
buf ( n2896 , n1143 );
buf ( n2897 , n2896 );
and ( n2898 , n2897 , n1657 );
and ( n2899 , n2894 , n2898 );
and ( n2900 , n2890 , n2898 );
or ( n2901 , n2895 , n2899 , n2900 );
and ( n2902 , n1799 , n2320 );
and ( n2903 , n1720 , n2318 );
nor ( n2904 , n2902 , n2903 );
xnor ( n2905 , n2904 , n2217 );
and ( n2906 , n2258 , n1807 );
and ( n2907 , n2181 , n1805 );
nor ( n2908 , n2906 , n2907 );
xnor ( n2909 , n2908 , n1756 );
and ( n2910 , n2905 , n2909 );
and ( n2911 , n2390 , n1728 );
and ( n2912 , n2295 , n1726 );
nor ( n2913 , n2911 , n2912 );
xnor ( n2914 , n2913 , n1697 );
and ( n2915 , n2909 , n2914 );
and ( n2916 , n2905 , n2914 );
or ( n2917 , n2910 , n2915 , n2916 );
and ( n2918 , n2901 , n2917 );
and ( n2919 , n1655 , n2654 );
and ( n2920 , n1666 , n2652 );
nor ( n2921 , n2919 , n2920 );
xnor ( n2922 , n2921 , n2570 );
buf ( n2923 , n2922 );
and ( n2924 , n2917 , n2923 );
and ( n2925 , n2901 , n2923 );
or ( n2926 , n2918 , n2924 , n2925 );
xor ( n2927 , n2777 , n2793 );
xor ( n2928 , n2927 , n2814 );
and ( n2929 , n2926 , n2928 );
xor ( n2930 , n2833 , n2834 );
xor ( n2931 , n2930 , n2839 );
and ( n2932 , n2928 , n2931 );
and ( n2933 , n2926 , n2931 );
or ( n2934 , n2929 , n2932 , n2933 );
xor ( n2935 , n2817 , n2842 );
xor ( n2936 , n2935 , n2845 );
and ( n2937 , n2934 , n2936 );
xor ( n2938 , n2858 , n2860 );
xor ( n2939 , n2938 , n2863 );
and ( n2940 , n2936 , n2939 );
and ( n2941 , n2934 , n2939 );
or ( n2942 , n2937 , n2940 , n2941 );
xor ( n2943 , n2737 , n2739 );
xor ( n2944 , n2943 , n2742 );
and ( n2945 , n2942 , n2944 );
xor ( n2946 , n2848 , n2866 );
xor ( n2947 , n2946 , n2869 );
and ( n2948 , n2944 , n2947 );
and ( n2949 , n2942 , n2947 );
or ( n2950 , n2945 , n2948 , n2949 );
and ( n2951 , n2883 , n2950 );
xor ( n2952 , n2942 , n2944 );
xor ( n2953 , n2952 , n2947 );
and ( n2954 , n1849 , n2113 );
and ( n2955 , n1817 , n2111 );
nor ( n2956 , n2954 , n2955 );
xnor ( n2957 , n2956 , n2091 );
and ( n2958 , n2615 , n1646 );
and ( n2959 , n2506 , n1644 );
nor ( n2960 , n2958 , n2959 );
xnor ( n2961 , n2960 , n1651 );
and ( n2962 , n2957 , n2961 );
and ( n2963 , n2773 , n1663 );
and ( n2964 , n2697 , n1661 );
nor ( n2965 , n2963 , n2964 );
xnor ( n2966 , n2965 , n1671 );
and ( n2967 , n2961 , n2966 );
and ( n2968 , n2957 , n2966 );
or ( n2969 , n2962 , n2967 , n2968 );
xor ( n2970 , n2766 , n2770 );
xor ( n2971 , n2970 , n2774 );
and ( n2972 , n2969 , n2971 );
xor ( n2973 , n2821 , n2825 );
xor ( n2974 , n2973 , n2830 );
and ( n2975 , n2971 , n2974 );
and ( n2976 , n2969 , n2974 );
or ( n2977 , n2972 , n2975 , n2976 );
not ( n2978 , n2922 );
and ( n2979 , n2027 , n2020 );
and ( n2980 , n1935 , n2018 );
nor ( n2981 , n2979 , n2980 );
xnor ( n2982 , n2981 , n1981 );
and ( n2983 , n2978 , n2982 );
and ( n2984 , n2080 , n1901 );
and ( n2985 , n2042 , n1899 );
nor ( n2986 , n2984 , n2985 );
xnor ( n2987 , n2986 , n1869 );
and ( n2988 , n2982 , n2987 );
and ( n2989 , n2978 , n2987 );
or ( n2990 , n2983 , n2988 , n2989 );
xor ( n2991 , n2781 , n2785 );
xor ( n2992 , n2991 , n2790 );
and ( n2993 , n2990 , n2992 );
xor ( n2994 , n2802 , n2806 );
xor ( n2995 , n2994 , n2811 );
and ( n2996 , n2992 , n2995 );
and ( n2997 , n2990 , n2995 );
or ( n2998 , n2993 , n2996 , n2997 );
and ( n2999 , n2977 , n2998 );
xor ( n3000 , n2850 , n2852 );
xor ( n3001 , n3000 , n2855 );
and ( n3002 , n2998 , n3001 );
and ( n3003 , n2977 , n3001 );
or ( n3004 , n2999 , n3002 , n3003 );
and ( n3005 , n1675 , n2654 );
and ( n3006 , n1655 , n2652 );
nor ( n3007 , n3005 , n3006 );
xnor ( n3008 , n3007 , n2570 );
and ( n3009 , n2506 , n1728 );
and ( n3010 , n2390 , n1726 );
nor ( n3011 , n3009 , n3010 );
xnor ( n3012 , n3011 , n1697 );
and ( n3013 , n3008 , n3012 );
and ( n3014 , n2697 , n1646 );
and ( n3015 , n2615 , n1644 );
nor ( n3016 , n3014 , n3015 );
xnor ( n3017 , n3016 , n1651 );
and ( n3018 , n3012 , n3017 );
and ( n3019 , n3008 , n3017 );
or ( n3020 , n3013 , n3018 , n3019 );
buf ( n3021 , n1177 );
buf ( n3022 , n3021 );
buf ( n3023 , n1178 );
buf ( n3024 , n3023 );
and ( n3025 , n3022 , n3024 );
not ( n3026 , n3025 );
and ( n3027 , n2798 , n3026 );
not ( n3028 , n3027 );
and ( n3029 , n1666 , n2887 );
and ( n3030 , n1636 , n2885 );
nor ( n3031 , n3029 , n3030 );
xnor ( n3032 , n3031 , n2801 );
and ( n3033 , n3028 , n3032 );
and ( n3034 , n1720 , n2483 );
and ( n3035 , n1705 , n2481 );
nor ( n3036 , n3034 , n3035 );
xnor ( n3037 , n3036 , n2418 );
and ( n3038 , n3032 , n3037 );
and ( n3039 , n3028 , n3037 );
or ( n3040 , n3033 , n3038 , n3039 );
and ( n3041 , n3020 , n3040 );
and ( n3042 , n1935 , n2113 );
and ( n3043 , n1849 , n2111 );
nor ( n3044 , n3042 , n3043 );
xnor ( n3045 , n3044 , n2091 );
and ( n3046 , n2897 , n1663 );
and ( n3047 , n2773 , n1661 );
nor ( n3048 , n3046 , n3047 );
xnor ( n3049 , n3048 , n1671 );
and ( n3050 , n3045 , n3049 );
buf ( n3051 , n1144 );
buf ( n3052 , n3051 );
and ( n3053 , n3052 , n1657 );
and ( n3054 , n3049 , n3053 );
and ( n3055 , n3045 , n3053 );
or ( n3056 , n3050 , n3054 , n3055 );
and ( n3057 , n3040 , n3056 );
and ( n3058 , n3020 , n3056 );
or ( n3059 , n3041 , n3057 , n3058 );
and ( n3060 , n1817 , n2320 );
and ( n3061 , n1799 , n2318 );
nor ( n3062 , n3060 , n3061 );
xnor ( n3063 , n3062 , n2217 );
and ( n3064 , n2181 , n1901 );
and ( n3065 , n2080 , n1899 );
nor ( n3066 , n3064 , n3065 );
xnor ( n3067 , n3066 , n1869 );
and ( n3068 , n3063 , n3067 );
and ( n3069 , n2295 , n1807 );
and ( n3070 , n2258 , n1805 );
nor ( n3071 , n3069 , n3070 );
xnor ( n3072 , n3071 , n1756 );
and ( n3073 , n3067 , n3072 );
and ( n3074 , n3063 , n3072 );
or ( n3075 , n3068 , n3073 , n3074 );
xor ( n3076 , n2890 , n2894 );
xor ( n3077 , n3076 , n2898 );
and ( n3078 , n3075 , n3077 );
xor ( n3079 , n2905 , n2909 );
xor ( n3080 , n3079 , n2914 );
and ( n3081 , n3077 , n3080 );
and ( n3082 , n3075 , n3080 );
or ( n3083 , n3078 , n3081 , n3082 );
and ( n3084 , n3059 , n3083 );
xor ( n3085 , n2901 , n2917 );
xor ( n3086 , n3085 , n2923 );
and ( n3087 , n3083 , n3086 );
and ( n3088 , n3059 , n3086 );
or ( n3089 , n3084 , n3087 , n3088 );
xor ( n3090 , n2798 , n3022 );
xor ( n3091 , n3022 , n3024 );
not ( n3092 , n3091 );
and ( n3093 , n3090 , n3092 );
and ( n3094 , n1636 , n3093 );
not ( n3095 , n3094 );
xnor ( n3096 , n3095 , n3027 );
and ( n3097 , n2027 , n2113 );
and ( n3098 , n1935 , n2111 );
nor ( n3099 , n3097 , n3098 );
xnor ( n3100 , n3099 , n2091 );
and ( n3101 , n3096 , n3100 );
and ( n3102 , n3052 , n1663 );
and ( n3103 , n2897 , n1661 );
nor ( n3104 , n3102 , n3103 );
xnor ( n3105 , n3104 , n1671 );
and ( n3106 , n3100 , n3105 );
and ( n3107 , n3096 , n3105 );
or ( n3108 , n3101 , n3106 , n3107 );
and ( n3109 , n1799 , n2483 );
and ( n3110 , n1720 , n2481 );
nor ( n3111 , n3109 , n3110 );
xnor ( n3112 , n3111 , n2418 );
and ( n3113 , n2258 , n1901 );
and ( n3114 , n2181 , n1899 );
nor ( n3115 , n3113 , n3114 );
xnor ( n3116 , n3115 , n1869 );
and ( n3117 , n3112 , n3116 );
and ( n3118 , n2390 , n1807 );
and ( n3119 , n2295 , n1805 );
nor ( n3120 , n3118 , n3119 );
xnor ( n3121 , n3120 , n1756 );
and ( n3122 , n3116 , n3121 );
and ( n3123 , n3112 , n3121 );
or ( n3124 , n3117 , n3122 , n3123 );
and ( n3125 , n3108 , n3124 );
and ( n3126 , n1705 , n2654 );
and ( n3127 , n1675 , n2652 );
nor ( n3128 , n3126 , n3127 );
xnor ( n3129 , n3128 , n2570 );
and ( n3130 , n2080 , n2020 );
and ( n3131 , n2042 , n2018 );
nor ( n3132 , n3130 , n3131 );
xnor ( n3133 , n3132 , n1981 );
and ( n3134 , n3129 , n3133 );
buf ( n3135 , n1145 );
buf ( n3136 , n3135 );
and ( n3137 , n3136 , n1657 );
and ( n3138 , n3133 , n3137 );
and ( n3139 , n3129 , n3137 );
or ( n3140 , n3134 , n3138 , n3139 );
and ( n3141 , n3124 , n3140 );
and ( n3142 , n3108 , n3140 );
or ( n3143 , n3125 , n3141 , n3142 );
xor ( n3144 , n2957 , n2961 );
xor ( n3145 , n3144 , n2966 );
and ( n3146 , n3143 , n3145 );
xor ( n3147 , n2978 , n2982 );
xor ( n3148 , n3147 , n2987 );
and ( n3149 , n3145 , n3148 );
and ( n3150 , n3143 , n3148 );
or ( n3151 , n3146 , n3149 , n3150 );
xor ( n3152 , n2969 , n2971 );
xor ( n3153 , n3152 , n2974 );
and ( n3154 , n3151 , n3153 );
xor ( n3155 , n2990 , n2992 );
xor ( n3156 , n3155 , n2995 );
and ( n3157 , n3153 , n3156 );
and ( n3158 , n3151 , n3156 );
or ( n3159 , n3154 , n3157 , n3158 );
and ( n3160 , n3089 , n3159 );
xor ( n3161 , n2926 , n2928 );
xor ( n3162 , n3161 , n2931 );
and ( n3163 , n3159 , n3162 );
and ( n3164 , n3089 , n3162 );
or ( n3165 , n3160 , n3163 , n3164 );
and ( n3166 , n3004 , n3165 );
xor ( n3167 , n2934 , n2936 );
xor ( n3168 , n3167 , n2939 );
and ( n3169 , n3165 , n3168 );
and ( n3170 , n3004 , n3168 );
or ( n3171 , n3166 , n3169 , n3170 );
and ( n3172 , n2953 , n3171 );
xor ( n3173 , n3004 , n3165 );
xor ( n3174 , n3173 , n3168 );
and ( n3175 , n1849 , n2320 );
and ( n3176 , n1817 , n2318 );
nor ( n3177 , n3175 , n3176 );
xnor ( n3178 , n3177 , n2217 );
and ( n3179 , n2615 , n1728 );
and ( n3180 , n2506 , n1726 );
nor ( n3181 , n3179 , n3180 );
xnor ( n3182 , n3181 , n1697 );
and ( n3183 , n3178 , n3182 );
and ( n3184 , n2773 , n1646 );
and ( n3185 , n2697 , n1644 );
nor ( n3186 , n3184 , n3185 );
xnor ( n3187 , n3186 , n1651 );
and ( n3188 , n3182 , n3187 );
and ( n3189 , n3178 , n3187 );
or ( n3190 , n3183 , n3188 , n3189 );
and ( n3191 , n1655 , n2887 );
and ( n3192 , n1666 , n2885 );
nor ( n3193 , n3191 , n3192 );
xnor ( n3194 , n3193 , n2801 );
buf ( n3195 , n3194 );
and ( n3196 , n3190 , n3195 );
and ( n3197 , n2042 , n2020 );
and ( n3198 , n2027 , n2018 );
nor ( n3199 , n3197 , n3198 );
xnor ( n3200 , n3199 , n1981 );
and ( n3201 , n3195 , n3200 );
and ( n3202 , n3190 , n3200 );
or ( n3203 , n3196 , n3201 , n3202 );
xor ( n3204 , n3063 , n3067 );
xor ( n3205 , n3204 , n3072 );
xor ( n3206 , n3008 , n3012 );
xor ( n3207 , n3206 , n3017 );
and ( n3208 , n3205 , n3207 );
xor ( n3209 , n3028 , n3032 );
xor ( n3210 , n3209 , n3037 );
and ( n3211 , n3207 , n3210 );
and ( n3212 , n3205 , n3210 );
or ( n3213 , n3208 , n3211 , n3212 );
and ( n3214 , n3203 , n3213 );
xor ( n3215 , n3020 , n3040 );
xor ( n3216 , n3215 , n3056 );
and ( n3217 , n3213 , n3216 );
and ( n3218 , n3203 , n3216 );
or ( n3219 , n3214 , n3217 , n3218 );
and ( n3220 , n1817 , n2483 );
and ( n3221 , n1799 , n2481 );
nor ( n3222 , n3220 , n3221 );
xnor ( n3223 , n3222 , n2418 );
and ( n3224 , n2181 , n2020 );
and ( n3225 , n2080 , n2018 );
nor ( n3226 , n3224 , n3225 );
xnor ( n3227 , n3226 , n1981 );
and ( n3228 , n3223 , n3227 );
and ( n3229 , n2295 , n1901 );
and ( n3230 , n2258 , n1899 );
nor ( n3231 , n3229 , n3230 );
xnor ( n3232 , n3231 , n1869 );
and ( n3233 , n3227 , n3232 );
and ( n3234 , n3223 , n3232 );
or ( n3235 , n3228 , n3233 , n3234 );
and ( n3236 , n1675 , n2887 );
and ( n3237 , n1655 , n2885 );
nor ( n3238 , n3236 , n3237 );
xnor ( n3239 , n3238 , n2801 );
and ( n3240 , n2506 , n1807 );
and ( n3241 , n2390 , n1805 );
nor ( n3242 , n3240 , n3241 );
xnor ( n3243 , n3242 , n1756 );
and ( n3244 , n3239 , n3243 );
and ( n3245 , n2697 , n1728 );
and ( n3246 , n2615 , n1726 );
nor ( n3247 , n3245 , n3246 );
xnor ( n3248 , n3247 , n1697 );
and ( n3249 , n3243 , n3248 );
and ( n3250 , n3239 , n3248 );
or ( n3251 , n3244 , n3249 , n3250 );
and ( n3252 , n3235 , n3251 );
not ( n3253 , n3194 );
and ( n3254 , n3251 , n3253 );
and ( n3255 , n3235 , n3253 );
or ( n3256 , n3252 , n3254 , n3255 );
xor ( n3257 , n3045 , n3049 );
xor ( n3258 , n3257 , n3053 );
and ( n3259 , n3256 , n3258 );
xor ( n3260 , n3190 , n3195 );
xor ( n3261 , n3260 , n3200 );
and ( n3262 , n3258 , n3261 );
and ( n3263 , n3256 , n3261 );
or ( n3264 , n3259 , n3262 , n3263 );
xor ( n3265 , n3075 , n3077 );
xor ( n3266 , n3265 , n3080 );
and ( n3267 , n3264 , n3266 );
xor ( n3268 , n3143 , n3145 );
xor ( n3269 , n3268 , n3148 );
and ( n3270 , n3266 , n3269 );
and ( n3271 , n3264 , n3269 );
or ( n3272 , n3267 , n3270 , n3271 );
and ( n3273 , n3219 , n3272 );
xor ( n3274 , n3059 , n3083 );
xor ( n3275 , n3274 , n3086 );
and ( n3276 , n3272 , n3275 );
and ( n3277 , n3219 , n3275 );
or ( n3278 , n3273 , n3276 , n3277 );
xor ( n3279 , n2977 , n2998 );
xor ( n3280 , n3279 , n3001 );
and ( n3281 , n3278 , n3280 );
xor ( n3282 , n3089 , n3159 );
xor ( n3283 , n3282 , n3162 );
and ( n3284 , n3280 , n3283 );
and ( n3285 , n3278 , n3283 );
or ( n3286 , n3281 , n3284 , n3285 );
and ( n3287 , n3174 , n3286 );
xor ( n3288 , n3278 , n3280 );
xor ( n3289 , n3288 , n3283 );
xor ( n3290 , n3096 , n3100 );
xor ( n3291 , n3290 , n3105 );
xor ( n3292 , n3112 , n3116 );
xor ( n3293 , n3292 , n3121 );
and ( n3294 , n3291 , n3293 );
xor ( n3295 , n3178 , n3182 );
xor ( n3296 , n3295 , n3187 );
and ( n3297 , n3293 , n3296 );
and ( n3298 , n3291 , n3296 );
or ( n3299 , n3294 , n3297 , n3298 );
buf ( n3300 , n1179 );
buf ( n3301 , n3300 );
buf ( n3302 , n1180 );
buf ( n3303 , n3302 );
and ( n3304 , n3301 , n3303 );
not ( n3305 , n3304 );
and ( n3306 , n3024 , n3305 );
not ( n3307 , n3306 );
and ( n3308 , n1666 , n3093 );
and ( n3309 , n1636 , n3091 );
nor ( n3310 , n3308 , n3309 );
xnor ( n3311 , n3310 , n3027 );
and ( n3312 , n3307 , n3311 );
and ( n3313 , n1720 , n2654 );
and ( n3314 , n1705 , n2652 );
nor ( n3315 , n3313 , n3314 );
xnor ( n3316 , n3315 , n2570 );
and ( n3317 , n3311 , n3316 );
and ( n3318 , n3307 , n3316 );
or ( n3319 , n3312 , n3317 , n3318 );
and ( n3320 , n1935 , n2320 );
and ( n3321 , n1849 , n2318 );
nor ( n3322 , n3320 , n3321 );
xnor ( n3323 , n3322 , n2217 );
and ( n3324 , n2897 , n1646 );
and ( n3325 , n2773 , n1644 );
nor ( n3326 , n3324 , n3325 );
xnor ( n3327 , n3326 , n1651 );
and ( n3328 , n3323 , n3327 );
and ( n3329 , n3136 , n1663 );
and ( n3330 , n3052 , n1661 );
nor ( n3331 , n3329 , n3330 );
xnor ( n3332 , n3331 , n1671 );
and ( n3333 , n3327 , n3332 );
and ( n3334 , n3323 , n3332 );
or ( n3335 , n3328 , n3333 , n3334 );
and ( n3336 , n3319 , n3335 );
xor ( n3337 , n3129 , n3133 );
xor ( n3338 , n3337 , n3137 );
and ( n3339 , n3335 , n3338 );
and ( n3340 , n3319 , n3338 );
or ( n3341 , n3336 , n3339 , n3340 );
and ( n3342 , n3299 , n3341 );
xor ( n3343 , n3108 , n3124 );
xor ( n3344 , n3343 , n3140 );
and ( n3345 , n3341 , n3344 );
and ( n3346 , n3299 , n3344 );
or ( n3347 , n3342 , n3345 , n3346 );
and ( n3348 , n1799 , n2654 );
and ( n3349 , n1720 , n2652 );
nor ( n3350 , n3348 , n3349 );
xnor ( n3351 , n3350 , n2570 );
and ( n3352 , n2258 , n2020 );
and ( n3353 , n2181 , n2018 );
nor ( n3354 , n3352 , n3353 );
xnor ( n3355 , n3354 , n1981 );
and ( n3356 , n3351 , n3355 );
and ( n3357 , n2390 , n1901 );
and ( n3358 , n2295 , n1899 );
nor ( n3359 , n3357 , n3358 );
xnor ( n3360 , n3359 , n1869 );
and ( n3361 , n3355 , n3360 );
and ( n3362 , n3351 , n3360 );
or ( n3363 , n3356 , n3361 , n3362 );
xor ( n3364 , n3024 , n3301 );
xor ( n3365 , n3301 , n3303 );
not ( n3366 , n3365 );
and ( n3367 , n3364 , n3366 );
and ( n3368 , n1636 , n3367 );
not ( n3369 , n3368 );
xnor ( n3370 , n3369 , n3306 );
and ( n3371 , n2027 , n2320 );
and ( n3372 , n1935 , n2318 );
nor ( n3373 , n3371 , n3372 );
xnor ( n3374 , n3373 , n2217 );
and ( n3375 , n3370 , n3374 );
and ( n3376 , n3052 , n1646 );
and ( n3377 , n2897 , n1644 );
nor ( n3378 , n3376 , n3377 );
xnor ( n3379 , n3378 , n1651 );
and ( n3380 , n3374 , n3379 );
and ( n3381 , n3370 , n3379 );
or ( n3382 , n3375 , n3380 , n3381 );
and ( n3383 , n3363 , n3382 );
and ( n3384 , n1849 , n2483 );
and ( n3385 , n1817 , n2481 );
nor ( n3386 , n3384 , n3385 );
xnor ( n3387 , n3386 , n2418 );
and ( n3388 , n2615 , n1807 );
and ( n3389 , n2506 , n1805 );
nor ( n3390 , n3388 , n3389 );
xnor ( n3391 , n3390 , n1756 );
and ( n3392 , n3387 , n3391 );
and ( n3393 , n2773 , n1728 );
and ( n3394 , n2697 , n1726 );
nor ( n3395 , n3393 , n3394 );
xnor ( n3396 , n3395 , n1697 );
and ( n3397 , n3391 , n3396 );
and ( n3398 , n3387 , n3396 );
or ( n3399 , n3392 , n3397 , n3398 );
and ( n3400 , n3382 , n3399 );
and ( n3401 , n3363 , n3399 );
or ( n3402 , n3383 , n3400 , n3401 );
and ( n3403 , n1655 , n3093 );
and ( n3404 , n1666 , n3091 );
nor ( n3405 , n3403 , n3404 );
xnor ( n3406 , n3405 , n3027 );
buf ( n3407 , n3406 );
and ( n3408 , n2042 , n2113 );
and ( n3409 , n2027 , n2111 );
nor ( n3410 , n3408 , n3409 );
xnor ( n3411 , n3410 , n2091 );
and ( n3412 , n3407 , n3411 );
buf ( n3413 , n1146 );
buf ( n3414 , n3413 );
and ( n3415 , n3414 , n1657 );
and ( n3416 , n3411 , n3415 );
and ( n3417 , n3407 , n3415 );
or ( n3418 , n3412 , n3416 , n3417 );
and ( n3419 , n3402 , n3418 );
xor ( n3420 , n3235 , n3251 );
xor ( n3421 , n3420 , n3253 );
and ( n3422 , n3418 , n3421 );
and ( n3423 , n3402 , n3421 );
or ( n3424 , n3419 , n3422 , n3423 );
xor ( n3425 , n3205 , n3207 );
xor ( n3426 , n3425 , n3210 );
and ( n3427 , n3424 , n3426 );
xor ( n3428 , n3256 , n3258 );
xor ( n3429 , n3428 , n3261 );
and ( n3430 , n3426 , n3429 );
and ( n3431 , n3424 , n3429 );
or ( n3432 , n3427 , n3430 , n3431 );
and ( n3433 , n3347 , n3432 );
xor ( n3434 , n3203 , n3213 );
xor ( n3435 , n3434 , n3216 );
and ( n3436 , n3432 , n3435 );
and ( n3437 , n3347 , n3435 );
or ( n3438 , n3433 , n3436 , n3437 );
xor ( n3439 , n3151 , n3153 );
xor ( n3440 , n3439 , n3156 );
and ( n3441 , n3438 , n3440 );
xor ( n3442 , n3219 , n3272 );
xor ( n3443 , n3442 , n3275 );
and ( n3444 , n3440 , n3443 );
and ( n3445 , n3438 , n3443 );
or ( n3446 , n3441 , n3444 , n3445 );
and ( n3447 , n3289 , n3446 );
xor ( n3448 , n3438 , n3440 );
xor ( n3449 , n3448 , n3443 );
xor ( n3450 , n3264 , n3266 );
xor ( n3451 , n3450 , n3269 );
xor ( n3452 , n3347 , n3432 );
xor ( n3453 , n3452 , n3435 );
and ( n3454 , n3451 , n3453 );
and ( n3455 , n3449 , n3454 );
and ( n3456 , n1705 , n2887 );
and ( n3457 , n1675 , n2885 );
nor ( n3458 , n3456 , n3457 );
xnor ( n3459 , n3458 , n2801 );
and ( n3460 , n3414 , n1663 );
and ( n3461 , n3136 , n1661 );
nor ( n3462 , n3460 , n3461 );
xnor ( n3463 , n3462 , n1671 );
and ( n3464 , n3459 , n3463 );
buf ( n3465 , n1147 );
buf ( n3466 , n3465 );
and ( n3467 , n3466 , n1657 );
and ( n3468 , n3463 , n3467 );
and ( n3469 , n3459 , n3467 );
or ( n3470 , n3464 , n3468 , n3469 );
xor ( n3471 , n3223 , n3227 );
xor ( n3472 , n3471 , n3232 );
and ( n3473 , n3470 , n3472 );
xor ( n3474 , n3307 , n3311 );
xor ( n3475 , n3474 , n3316 );
and ( n3476 , n3472 , n3475 );
and ( n3477 , n3470 , n3475 );
or ( n3478 , n3473 , n3476 , n3477 );
xor ( n3479 , n3239 , n3243 );
xor ( n3480 , n3479 , n3248 );
xor ( n3481 , n3323 , n3327 );
xor ( n3482 , n3481 , n3332 );
and ( n3483 , n3480 , n3482 );
xor ( n3484 , n3407 , n3411 );
xor ( n3485 , n3484 , n3415 );
and ( n3486 , n3482 , n3485 );
and ( n3487 , n3480 , n3485 );
or ( n3488 , n3483 , n3486 , n3487 );
and ( n3489 , n3478 , n3488 );
xor ( n3490 , n3319 , n3335 );
xor ( n3491 , n3490 , n3338 );
and ( n3492 , n3488 , n3491 );
and ( n3493 , n3478 , n3491 );
or ( n3494 , n3489 , n3492 , n3493 );
xor ( n3495 , n3299 , n3341 );
xor ( n3496 , n3495 , n3344 );
and ( n3497 , n3494 , n3496 );
xor ( n3498 , n3451 , n3453 );
and ( n3499 , n3497 , n3498 );
xor ( n3500 , n3424 , n3426 );
xor ( n3501 , n3500 , n3429 );
xor ( n3502 , n3291 , n3293 );
xor ( n3503 , n3502 , n3296 );
xor ( n3504 , n3363 , n3382 );
xor ( n3505 , n3504 , n3399 );
and ( n3506 , n1935 , n2483 );
and ( n3507 , n1849 , n2481 );
nor ( n3508 , n3506 , n3507 );
xnor ( n3509 , n3508 , n2418 );
and ( n3510 , n2897 , n1728 );
and ( n3511 , n2773 , n1726 );
nor ( n3512 , n3510 , n3511 );
xnor ( n3513 , n3512 , n1697 );
and ( n3514 , n3509 , n3513 );
and ( n3515 , n3136 , n1646 );
and ( n3516 , n3052 , n1644 );
nor ( n3517 , n3515 , n3516 );
xnor ( n3518 , n3517 , n1651 );
and ( n3519 , n3513 , n3518 );
and ( n3520 , n3509 , n3518 );
or ( n3521 , n3514 , n3519 , n3520 );
not ( n3522 , n3406 );
and ( n3523 , n3521 , n3522 );
and ( n3524 , n2080 , n2113 );
and ( n3525 , n2042 , n2111 );
nor ( n3526 , n3524 , n3525 );
xnor ( n3527 , n3526 , n2091 );
and ( n3528 , n3522 , n3527 );
and ( n3529 , n3521 , n3527 );
or ( n3530 , n3523 , n3528 , n3529 );
and ( n3531 , n3505 , n3530 );
buf ( n3532 , n1181 );
buf ( n3533 , n3532 );
buf ( n3534 , n1182 );
buf ( n3535 , n3534 );
and ( n3536 , n3533 , n3535 );
not ( n3537 , n3536 );
and ( n3538 , n3303 , n3537 );
not ( n3539 , n3538 );
and ( n3540 , n1666 , n3367 );
and ( n3541 , n1636 , n3365 );
nor ( n3542 , n3540 , n3541 );
xnor ( n3543 , n3542 , n3306 );
and ( n3544 , n3539 , n3543 );
and ( n3545 , n1720 , n2887 );
and ( n3546 , n1705 , n2885 );
nor ( n3547 , n3545 , n3546 );
xnor ( n3548 , n3547 , n2801 );
and ( n3549 , n3543 , n3548 );
and ( n3550 , n3539 , n3548 );
or ( n3551 , n3544 , n3549 , n3550 );
and ( n3552 , n1675 , n3093 );
and ( n3553 , n1655 , n3091 );
nor ( n3554 , n3552 , n3553 );
xnor ( n3555 , n3554 , n3027 );
and ( n3556 , n2506 , n1901 );
and ( n3557 , n2390 , n1899 );
nor ( n3558 , n3556 , n3557 );
xnor ( n3559 , n3558 , n1869 );
and ( n3560 , n3555 , n3559 );
and ( n3561 , n2697 , n1807 );
and ( n3562 , n2615 , n1805 );
nor ( n3563 , n3561 , n3562 );
xnor ( n3564 , n3563 , n1756 );
and ( n3565 , n3559 , n3564 );
and ( n3566 , n3555 , n3564 );
or ( n3567 , n3560 , n3565 , n3566 );
and ( n3568 , n3551 , n3567 );
and ( n3569 , n1817 , n2654 );
and ( n3570 , n1799 , n2652 );
nor ( n3571 , n3569 , n3570 );
xnor ( n3572 , n3571 , n2570 );
and ( n3573 , n2181 , n2113 );
and ( n3574 , n2080 , n2111 );
nor ( n3575 , n3573 , n3574 );
xnor ( n3576 , n3575 , n2091 );
and ( n3577 , n3572 , n3576 );
and ( n3578 , n2295 , n2020 );
and ( n3579 , n2258 , n2018 );
nor ( n3580 , n3578 , n3579 );
xnor ( n3581 , n3580 , n1981 );
and ( n3582 , n3576 , n3581 );
and ( n3583 , n3572 , n3581 );
or ( n3584 , n3577 , n3582 , n3583 );
and ( n3585 , n3567 , n3584 );
and ( n3586 , n3551 , n3584 );
or ( n3587 , n3568 , n3585 , n3586 );
and ( n3588 , n3530 , n3587 );
and ( n3589 , n3505 , n3587 );
or ( n3590 , n3531 , n3588 , n3589 );
and ( n3591 , n3503 , n3590 );
xor ( n3592 , n3402 , n3418 );
xor ( n3593 , n3592 , n3421 );
and ( n3594 , n3590 , n3593 );
and ( n3595 , n3503 , n3593 );
or ( n3596 , n3591 , n3594 , n3595 );
and ( n3597 , n3501 , n3596 );
xor ( n3598 , n3494 , n3496 );
and ( n3599 , n3596 , n3598 );
and ( n3600 , n3501 , n3598 );
or ( n3601 , n3597 , n3599 , n3600 );
and ( n3602 , n3498 , n3601 );
and ( n3603 , n3497 , n3601 );
or ( n3604 , n3499 , n3602 , n3603 );
and ( n3605 , n3454 , n3604 );
and ( n3606 , n3449 , n3604 );
or ( n3607 , n3455 , n3605 , n3606 );
and ( n3608 , n3446 , n3607 );
and ( n3609 , n3289 , n3607 );
or ( n3610 , n3447 , n3608 , n3609 );
and ( n3611 , n3286 , n3610 );
and ( n3612 , n3174 , n3610 );
or ( n3613 , n3287 , n3611 , n3612 );
and ( n3614 , n3171 , n3613 );
and ( n3615 , n2953 , n3613 );
or ( n3616 , n3172 , n3614 , n3615 );
and ( n3617 , n2950 , n3616 );
and ( n3618 , n2883 , n3616 );
or ( n3619 , n2951 , n3617 , n3618 );
and ( n3620 , n2880 , n3619 );
and ( n3621 , n2762 , n3619 );
or ( n3622 , n2881 , n3620 , n3621 );
and ( n3623 , n2759 , n3622 );
and ( n3624 , n2650 , n3622 );
or ( n3625 , n2760 , n3623 , n3624 );
and ( n3626 , n2647 , n3625 );
and ( n3627 , n2553 , n3625 );
or ( n3628 , n2648 , n3626 , n3627 );
and ( n3629 , n2550 , n3628 );
and ( n3630 , n2379 , n3628 );
or ( n3631 , n2551 , n3629 , n3630 );
and ( n3632 , n2376 , n3631 );
and ( n3633 , n2374 , n3631 );
or ( n3634 , n2377 , n3632 , n3633 );
and ( n3635 , n2347 , n3634 );
and ( n3636 , n2210 , n3634 );
or ( n3637 , n2348 , n3635 , n3636 );
and ( n3638 , n2207 , n3637 );
and ( n3639 , n2154 , n3637 );
or ( n3640 , n2208 , n3638 , n3639 );
and ( n3641 , n2151 , n3640 );
and ( n3642 , n2069 , n3640 );
or ( n3643 , n2152 , n3641 , n3642 );
and ( n3644 , n2066 , n3643 );
and ( n3645 , n1958 , n3643 );
or ( n3646 , n2067 , n3644 , n3645 );
and ( n3647 , n1955 , n3646 );
and ( n3648 , n1953 , n3646 );
or ( n3649 , n1956 , n3647 , n3648 );
and ( n3650 , n1896 , n3649 );
and ( n3651 , n1838 , n3649 );
or ( n3652 , n1897 , n3650 , n3651 );
and ( n3653 , n1835 , n3652 );
and ( n3654 , n1787 , n3652 );
or ( n3655 , n1836 , n3653 , n3654 );
and ( n3656 , n1784 , n3655 );
and ( n3657 , n1749 , n3655 );
or ( n3658 , n1785 , n3656 , n3657 );
xor ( n3659 , n1747 , n3658 );
xor ( n3660 , n1749 , n1784 );
xor ( n3661 , n3660 , n3655 );
xor ( n3662 , n1787 , n1835 );
xor ( n3663 , n3662 , n3652 );
xor ( n3664 , n1838 , n1896 );
xor ( n3665 , n3664 , n3649 );
xor ( n3666 , n1953 , n1955 );
xor ( n3667 , n3666 , n3646 );
xor ( n3668 , n1958 , n2066 );
xor ( n3669 , n3668 , n3643 );
xor ( n3670 , n2069 , n2151 );
xor ( n3671 , n3670 , n3640 );
xor ( n3672 , n2154 , n2207 );
xor ( n3673 , n3672 , n3637 );
xor ( n3674 , n2210 , n2347 );
xor ( n3675 , n3674 , n3634 );
xor ( n3676 , n2374 , n2376 );
xor ( n3677 , n3676 , n3631 );
xor ( n3678 , n2379 , n2550 );
xor ( n3679 , n3678 , n3628 );
xor ( n3680 , n2553 , n2647 );
xor ( n3681 , n3680 , n3625 );
xor ( n3682 , n2650 , n2759 );
xor ( n3683 , n3682 , n3622 );
xor ( n3684 , n2762 , n2880 );
xor ( n3685 , n3684 , n3619 );
xor ( n3686 , n2883 , n2950 );
xor ( n3687 , n3686 , n3616 );
xor ( n3688 , n2953 , n3171 );
xor ( n3689 , n3688 , n3613 );
xor ( n3690 , n3174 , n3286 );
xor ( n3691 , n3690 , n3610 );
xor ( n3692 , n3289 , n3446 );
xor ( n3693 , n3692 , n3607 );
xor ( n3694 , n3449 , n3454 );
xor ( n3695 , n3694 , n3604 );
xor ( n3696 , n3370 , n3374 );
xor ( n3697 , n3696 , n3379 );
xor ( n3698 , n3387 , n3391 );
xor ( n3699 , n3698 , n3396 );
and ( n3700 , n3697 , n3699 );
xor ( n3701 , n3521 , n3522 );
xor ( n3702 , n3701 , n3527 );
and ( n3703 , n3699 , n3702 );
and ( n3704 , n3697 , n3702 );
or ( n3705 , n3700 , n3703 , n3704 );
and ( n3706 , n1655 , n3367 );
and ( n3707 , n1666 , n3365 );
nor ( n3708 , n3706 , n3707 );
xnor ( n3709 , n3708 , n3306 );
and ( n3710 , n1799 , n2887 );
and ( n3711 , n1720 , n2885 );
nor ( n3712 , n3710 , n3711 );
xnor ( n3713 , n3712 , n2801 );
and ( n3714 , n3709 , n3713 );
and ( n3715 , n2258 , n2113 );
and ( n3716 , n2181 , n2111 );
nor ( n3717 , n3715 , n3716 );
xnor ( n3718 , n3717 , n2091 );
and ( n3719 , n3713 , n3718 );
and ( n3720 , n3709 , n3718 );
or ( n3721 , n3714 , n3719 , n3720 );
and ( n3722 , n1849 , n2654 );
and ( n3723 , n1817 , n2652 );
nor ( n3724 , n3722 , n3723 );
xnor ( n3725 , n3724 , n2570 );
and ( n3726 , n2390 , n2020 );
and ( n3727 , n2295 , n2018 );
nor ( n3728 , n3726 , n3727 );
xnor ( n3729 , n3728 , n1981 );
and ( n3730 , n3725 , n3729 );
and ( n3731 , n2615 , n1901 );
and ( n3732 , n2506 , n1899 );
nor ( n3733 , n3731 , n3732 );
xnor ( n3734 , n3733 , n1869 );
and ( n3735 , n3729 , n3734 );
and ( n3736 , n3725 , n3734 );
or ( n3737 , n3730 , n3735 , n3736 );
and ( n3738 , n3721 , n3737 );
xor ( n3739 , n3303 , n3533 );
xor ( n3740 , n3533 , n3535 );
not ( n3741 , n3740 );
and ( n3742 , n3739 , n3741 );
and ( n3743 , n1636 , n3742 );
not ( n3744 , n3743 );
xnor ( n3745 , n3744 , n3538 );
buf ( n3746 , n3745 );
and ( n3747 , n3737 , n3746 );
and ( n3748 , n3721 , n3746 );
or ( n3749 , n3738 , n3747 , n3748 );
and ( n3750 , n2080 , n2320 );
and ( n3751 , n2042 , n2318 );
nor ( n3752 , n3750 , n3751 );
xnor ( n3753 , n3752 , n2217 );
and ( n3754 , n3052 , n1728 );
and ( n3755 , n2897 , n1726 );
nor ( n3756 , n3754 , n3755 );
xnor ( n3757 , n3756 , n1697 );
and ( n3758 , n3753 , n3757 );
and ( n3759 , n3414 , n1646 );
and ( n3760 , n3136 , n1644 );
nor ( n3761 , n3759 , n3760 );
xnor ( n3762 , n3761 , n1651 );
and ( n3763 , n3757 , n3762 );
and ( n3764 , n3753 , n3762 );
or ( n3765 , n3758 , n3763 , n3764 );
and ( n3766 , n1705 , n3093 );
and ( n3767 , n1675 , n3091 );
nor ( n3768 , n3766 , n3767 );
xnor ( n3769 , n3768 , n3027 );
and ( n3770 , n2027 , n2483 );
and ( n3771 , n1935 , n2481 );
nor ( n3772 , n3770 , n3771 );
xnor ( n3773 , n3772 , n2418 );
and ( n3774 , n3769 , n3773 );
and ( n3775 , n2773 , n1807 );
and ( n3776 , n2697 , n1805 );
nor ( n3777 , n3775 , n3776 );
xnor ( n3778 , n3777 , n1756 );
and ( n3779 , n3773 , n3778 );
and ( n3780 , n3769 , n3778 );
or ( n3781 , n3774 , n3779 , n3780 );
and ( n3782 , n3765 , n3781 );
xor ( n3783 , n3572 , n3576 );
xor ( n3784 , n3783 , n3581 );
and ( n3785 , n3781 , n3784 );
and ( n3786 , n3765 , n3784 );
or ( n3787 , n3782 , n3785 , n3786 );
and ( n3788 , n3749 , n3787 );
xor ( n3789 , n3551 , n3567 );
xor ( n3790 , n3789 , n3584 );
and ( n3791 , n3787 , n3790 );
and ( n3792 , n3749 , n3790 );
or ( n3793 , n3788 , n3791 , n3792 );
and ( n3794 , n3705 , n3793 );
xor ( n3795 , n3505 , n3530 );
xor ( n3796 , n3795 , n3587 );
and ( n3797 , n3793 , n3796 );
and ( n3798 , n3705 , n3796 );
or ( n3799 , n3794 , n3797 , n3798 );
xor ( n3800 , n3478 , n3488 );
xor ( n3801 , n3800 , n3491 );
and ( n3802 , n3799 , n3801 );
and ( n3803 , n2042 , n2320 );
and ( n3804 , n2027 , n2318 );
nor ( n3805 , n3803 , n3804 );
xnor ( n3806 , n3805 , n2217 );
and ( n3807 , n3466 , n1663 );
and ( n3808 , n3414 , n1661 );
nor ( n3809 , n3807 , n3808 );
xnor ( n3810 , n3809 , n1671 );
and ( n3811 , n3806 , n3810 );
buf ( n3812 , n1148 );
buf ( n3813 , n3812 );
and ( n3814 , n3813 , n1657 );
and ( n3815 , n3810 , n3814 );
and ( n3816 , n3806 , n3814 );
or ( n3817 , n3811 , n3815 , n3816 );
xor ( n3818 , n3459 , n3463 );
xor ( n3819 , n3818 , n3467 );
and ( n3820 , n3817 , n3819 );
xor ( n3821 , n3351 , n3355 );
xor ( n3822 , n3821 , n3360 );
and ( n3823 , n3819 , n3822 );
and ( n3824 , n3817 , n3822 );
or ( n3825 , n3820 , n3823 , n3824 );
xor ( n3826 , n3470 , n3472 );
xor ( n3827 , n3826 , n3475 );
and ( n3828 , n3825 , n3827 );
xor ( n3829 , n3480 , n3482 );
xor ( n3830 , n3829 , n3485 );
and ( n3831 , n3827 , n3830 );
and ( n3832 , n3825 , n3830 );
or ( n3833 , n3828 , n3831 , n3832 );
and ( n3834 , n3801 , n3833 );
and ( n3835 , n3799 , n3833 );
or ( n3836 , n3802 , n3834 , n3835 );
xor ( n3837 , n3503 , n3590 );
xor ( n3838 , n3837 , n3593 );
xor ( n3839 , n3806 , n3810 );
xor ( n3840 , n3839 , n3814 );
xor ( n3841 , n3539 , n3543 );
xor ( n3842 , n3841 , n3548 );
and ( n3843 , n3840 , n3842 );
xor ( n3844 , n3509 , n3513 );
xor ( n3845 , n3844 , n3518 );
and ( n3846 , n3842 , n3845 );
and ( n3847 , n3840 , n3845 );
or ( n3848 , n3843 , n3846 , n3847 );
and ( n3849 , n2181 , n2320 );
and ( n3850 , n2080 , n2318 );
nor ( n3851 , n3849 , n3850 );
xnor ( n3852 , n3851 , n2217 );
and ( n3853 , n2295 , n2113 );
and ( n3854 , n2258 , n2111 );
nor ( n3855 , n3853 , n3854 );
xnor ( n3856 , n3855 , n2091 );
and ( n3857 , n3852 , n3856 );
buf ( n3858 , n1150 );
buf ( n3859 , n3858 );
and ( n3860 , n3859 , n1657 );
and ( n3861 , n3856 , n3860 );
and ( n3862 , n3852 , n3860 );
or ( n3863 , n3857 , n3861 , n3862 );
buf ( n3864 , n1183 );
buf ( n3865 , n3864 );
buf ( n3866 , n1184 );
buf ( n3867 , n3866 );
and ( n3868 , n3865 , n3867 );
not ( n3869 , n3868 );
and ( n3870 , n3535 , n3869 );
not ( n3871 , n3870 );
and ( n3872 , n1666 , n3742 );
and ( n3873 , n1636 , n3740 );
nor ( n3874 , n3872 , n3873 );
xnor ( n3875 , n3874 , n3538 );
and ( n3876 , n3871 , n3875 );
and ( n3877 , n1720 , n3093 );
and ( n3878 , n1705 , n3091 );
nor ( n3879 , n3877 , n3878 );
xnor ( n3880 , n3879 , n3027 );
and ( n3881 , n3875 , n3880 );
and ( n3882 , n3871 , n3880 );
or ( n3883 , n3876 , n3881 , n3882 );
and ( n3884 , n3863 , n3883 );
and ( n3885 , n1817 , n2887 );
and ( n3886 , n1799 , n2885 );
nor ( n3887 , n3885 , n3886 );
xnor ( n3888 , n3887 , n2801 );
and ( n3889 , n2506 , n2020 );
and ( n3890 , n2390 , n2018 );
nor ( n3891 , n3889 , n3890 );
xnor ( n3892 , n3891 , n1981 );
and ( n3893 , n3888 , n3892 );
and ( n3894 , n2697 , n1901 );
and ( n3895 , n2615 , n1899 );
nor ( n3896 , n3894 , n3895 );
xnor ( n3897 , n3896 , n1869 );
and ( n3898 , n3892 , n3897 );
and ( n3899 , n3888 , n3897 );
or ( n3900 , n3893 , n3898 , n3899 );
and ( n3901 , n3883 , n3900 );
and ( n3902 , n3863 , n3900 );
or ( n3903 , n3884 , n3901 , n3902 );
not ( n3904 , n3745 );
and ( n3905 , n3813 , n1663 );
and ( n3906 , n3466 , n1661 );
nor ( n3907 , n3905 , n3906 );
xnor ( n3908 , n3907 , n1671 );
and ( n3909 , n3904 , n3908 );
buf ( n3910 , n1149 );
buf ( n3911 , n3910 );
and ( n3912 , n3911 , n1657 );
and ( n3913 , n3908 , n3912 );
and ( n3914 , n3904 , n3912 );
or ( n3915 , n3909 , n3913 , n3914 );
and ( n3916 , n3903 , n3915 );
xor ( n3917 , n3555 , n3559 );
xor ( n3918 , n3917 , n3564 );
and ( n3919 , n3915 , n3918 );
and ( n3920 , n3903 , n3918 );
or ( n3921 , n3916 , n3919 , n3920 );
and ( n3922 , n3848 , n3921 );
xor ( n3923 , n3817 , n3819 );
xor ( n3924 , n3923 , n3822 );
and ( n3925 , n3921 , n3924 );
and ( n3926 , n3848 , n3924 );
or ( n3927 , n3922 , n3925 , n3926 );
xor ( n3928 , n3825 , n3827 );
xor ( n3929 , n3928 , n3830 );
and ( n3930 , n3927 , n3929 );
and ( n3931 , n3838 , n3930 );
xor ( n3932 , n3697 , n3699 );
xor ( n3933 , n3932 , n3702 );
and ( n3934 , n2042 , n2483 );
and ( n3935 , n2027 , n2481 );
nor ( n3936 , n3934 , n3935 );
xnor ( n3937 , n3936 , n2418 );
and ( n3938 , n3136 , n1728 );
and ( n3939 , n3052 , n1726 );
nor ( n3940 , n3938 , n3939 );
xnor ( n3941 , n3940 , n1697 );
and ( n3942 , n3937 , n3941 );
and ( n3943 , n3466 , n1646 );
and ( n3944 , n3414 , n1644 );
nor ( n3945 , n3943 , n3944 );
xnor ( n3946 , n3945 , n1651 );
and ( n3947 , n3941 , n3946 );
and ( n3948 , n3937 , n3946 );
or ( n3949 , n3942 , n3947 , n3948 );
and ( n3950 , n1675 , n3367 );
and ( n3951 , n1655 , n3365 );
nor ( n3952 , n3950 , n3951 );
xnor ( n3953 , n3952 , n3306 );
and ( n3954 , n1935 , n2654 );
and ( n3955 , n1849 , n2652 );
nor ( n3956 , n3954 , n3955 );
xnor ( n3957 , n3956 , n2570 );
and ( n3958 , n3953 , n3957 );
and ( n3959 , n2897 , n1807 );
and ( n3960 , n2773 , n1805 );
nor ( n3961 , n3959 , n3960 );
xnor ( n3962 , n3961 , n1756 );
and ( n3963 , n3957 , n3962 );
and ( n3964 , n3953 , n3962 );
or ( n3965 , n3958 , n3963 , n3964 );
and ( n3966 , n3949 , n3965 );
xor ( n3967 , n3709 , n3713 );
xor ( n3968 , n3967 , n3718 );
and ( n3969 , n3965 , n3968 );
and ( n3970 , n3949 , n3968 );
or ( n3971 , n3966 , n3969 , n3970 );
xor ( n3972 , n3721 , n3737 );
xor ( n3973 , n3972 , n3746 );
and ( n3974 , n3971 , n3973 );
xor ( n3975 , n3765 , n3781 );
xor ( n3976 , n3975 , n3784 );
and ( n3977 , n3973 , n3976 );
and ( n3978 , n3971 , n3976 );
or ( n3979 , n3974 , n3977 , n3978 );
and ( n3980 , n3933 , n3979 );
xor ( n3981 , n3749 , n3787 );
xor ( n3982 , n3981 , n3790 );
and ( n3983 , n3979 , n3982 );
and ( n3984 , n3933 , n3982 );
or ( n3985 , n3980 , n3983 , n3984 );
xor ( n3986 , n3705 , n3793 );
xor ( n3987 , n3986 , n3796 );
and ( n3988 , n3985 , n3987 );
xor ( n3989 , n3753 , n3757 );
xor ( n3990 , n3989 , n3762 );
xor ( n3991 , n3725 , n3729 );
xor ( n3992 , n3991 , n3734 );
and ( n3993 , n3990 , n3992 );
xor ( n3994 , n3769 , n3773 );
xor ( n3995 , n3994 , n3778 );
and ( n3996 , n3992 , n3995 );
and ( n3997 , n3990 , n3995 );
or ( n3998 , n3993 , n3996 , n3997 );
xor ( n3999 , n3840 , n3842 );
xor ( n4000 , n3999 , n3845 );
and ( n4001 , n3998 , n4000 );
xor ( n4002 , n3903 , n3915 );
xor ( n4003 , n4002 , n3918 );
and ( n4004 , n4000 , n4003 );
and ( n4005 , n3998 , n4003 );
or ( n4006 , n4001 , n4004 , n4005 );
xor ( n4007 , n3848 , n3921 );
xor ( n4008 , n4007 , n3924 );
and ( n4009 , n4006 , n4008 );
and ( n4010 , n3987 , n4009 );
and ( n4011 , n3985 , n4009 );
or ( n4012 , n3988 , n4010 , n4011 );
and ( n4013 , n3930 , n4012 );
and ( n4014 , n3838 , n4012 );
or ( n4015 , n3931 , n4013 , n4014 );
and ( n4016 , n3836 , n4015 );
xor ( n4017 , n3501 , n3596 );
xor ( n4018 , n4017 , n3598 );
and ( n4019 , n4015 , n4018 );
and ( n4020 , n3836 , n4018 );
or ( n4021 , n4016 , n4019 , n4020 );
xor ( n4022 , n3497 , n3498 );
xor ( n4023 , n4022 , n3601 );
and ( n4024 , n4021 , n4023 );
xor ( n4025 , n4021 , n4023 );
xor ( n4026 , n3836 , n4015 );
xor ( n4027 , n4026 , n4018 );
xor ( n4028 , n3799 , n3801 );
xor ( n4029 , n4028 , n3833 );
xor ( n4030 , n3838 , n3930 );
xor ( n4031 , n4030 , n4012 );
and ( n4032 , n4029 , n4031 );
xor ( n4033 , n3927 , n3929 );
xor ( n4034 , n3985 , n3987 );
xor ( n4035 , n4034 , n4009 );
and ( n4036 , n4033 , n4035 );
and ( n4037 , n1849 , n2887 );
and ( n4038 , n1817 , n2885 );
nor ( n4039 , n4037 , n4038 );
xnor ( n4040 , n4039 , n2801 );
and ( n4041 , n2258 , n2320 );
and ( n4042 , n2181 , n2318 );
nor ( n4043 , n4041 , n4042 );
xnor ( n4044 , n4043 , n2217 );
and ( n4045 , n4040 , n4044 );
and ( n4046 , n2390 , n2113 );
and ( n4047 , n2295 , n2111 );
nor ( n4048 , n4046 , n4047 );
xnor ( n4049 , n4048 , n2091 );
and ( n4050 , n4044 , n4049 );
and ( n4051 , n4040 , n4049 );
or ( n4052 , n4045 , n4050 , n4051 );
and ( n4053 , n1705 , n3367 );
and ( n4054 , n1675 , n3365 );
nor ( n4055 , n4053 , n4054 );
xnor ( n4056 , n4055 , n3306 );
and ( n4057 , n2615 , n2020 );
and ( n4058 , n2506 , n2018 );
nor ( n4059 , n4057 , n4058 );
xnor ( n4060 , n4059 , n1981 );
and ( n4061 , n4056 , n4060 );
and ( n4062 , n2773 , n1901 );
and ( n4063 , n2697 , n1899 );
nor ( n4064 , n4062 , n4063 );
xnor ( n4065 , n4064 , n1869 );
and ( n4066 , n4060 , n4065 );
and ( n4067 , n4056 , n4065 );
or ( n4068 , n4061 , n4066 , n4067 );
and ( n4069 , n4052 , n4068 );
and ( n4070 , n2027 , n2654 );
and ( n4071 , n1935 , n2652 );
nor ( n4072 , n4070 , n4071 );
xnor ( n4073 , n4072 , n2570 );
and ( n4074 , n3052 , n1807 );
and ( n4075 , n2897 , n1805 );
nor ( n4076 , n4074 , n4075 );
xnor ( n4077 , n4076 , n1756 );
and ( n4078 , n4073 , n4077 );
and ( n4079 , n3414 , n1728 );
and ( n4080 , n3136 , n1726 );
nor ( n4081 , n4079 , n4080 );
xnor ( n4082 , n4081 , n1697 );
and ( n4083 , n4077 , n4082 );
and ( n4084 , n4073 , n4082 );
or ( n4085 , n4078 , n4083 , n4084 );
and ( n4086 , n4068 , n4085 );
and ( n4087 , n4052 , n4085 );
or ( n4088 , n4069 , n4086 , n4087 );
and ( n4089 , n1655 , n3742 );
and ( n4090 , n1666 , n3740 );
nor ( n4091 , n4089 , n4090 );
xnor ( n4092 , n4091 , n3538 );
and ( n4093 , n1799 , n3093 );
and ( n4094 , n1720 , n3091 );
nor ( n4095 , n4093 , n4094 );
xnor ( n4096 , n4095 , n3027 );
and ( n4097 , n4092 , n4096 );
buf ( n4098 , n1151 );
buf ( n4099 , n4098 );
and ( n4100 , n4099 , n1657 );
and ( n4101 , n4096 , n4100 );
and ( n4102 , n4092 , n4100 );
or ( n4103 , n4097 , n4101 , n4102 );
xor ( n4104 , n3535 , n3865 );
xor ( n4105 , n3865 , n3867 );
not ( n4106 , n4105 );
and ( n4107 , n4104 , n4106 );
and ( n4108 , n1636 , n4107 );
not ( n4109 , n4108 );
xnor ( n4110 , n4109 , n3870 );
buf ( n4111 , n4110 );
and ( n4112 , n4103 , n4111 );
and ( n4113 , n3911 , n1663 );
and ( n4114 , n3813 , n1661 );
nor ( n4115 , n4113 , n4114 );
xnor ( n4116 , n4115 , n1671 );
and ( n4117 , n4111 , n4116 );
and ( n4118 , n4103 , n4116 );
or ( n4119 , n4112 , n4117 , n4118 );
and ( n4120 , n4088 , n4119 );
xor ( n4121 , n3904 , n3908 );
xor ( n4122 , n4121 , n3912 );
and ( n4123 , n4119 , n4122 );
and ( n4124 , n4088 , n4122 );
or ( n4125 , n4120 , n4123 , n4124 );
and ( n4126 , n2080 , n2483 );
and ( n4127 , n2042 , n2481 );
nor ( n4128 , n4126 , n4127 );
xnor ( n4129 , n4128 , n2418 );
and ( n4130 , n3813 , n1646 );
and ( n4131 , n3466 , n1644 );
nor ( n4132 , n4130 , n4131 );
xnor ( n4133 , n4132 , n1651 );
and ( n4134 , n4129 , n4133 );
and ( n4135 , n3859 , n1663 );
and ( n4136 , n3911 , n1661 );
nor ( n4137 , n4135 , n4136 );
xnor ( n4138 , n4137 , n1671 );
and ( n4139 , n4133 , n4138 );
and ( n4140 , n4129 , n4138 );
or ( n4141 , n4134 , n4139 , n4140 );
xor ( n4142 , n3852 , n3856 );
xor ( n4143 , n4142 , n3860 );
and ( n4144 , n4141 , n4143 );
xor ( n4145 , n3871 , n3875 );
xor ( n4146 , n4145 , n3880 );
and ( n4147 , n4143 , n4146 );
and ( n4148 , n4141 , n4146 );
or ( n4149 , n4144 , n4147 , n4148 );
xor ( n4150 , n3863 , n3883 );
xor ( n4151 , n4150 , n3900 );
and ( n4152 , n4149 , n4151 );
xor ( n4153 , n3949 , n3965 );
xor ( n4154 , n4153 , n3968 );
and ( n4155 , n4151 , n4154 );
and ( n4156 , n4149 , n4154 );
or ( n4157 , n4152 , n4155 , n4156 );
and ( n4158 , n4125 , n4157 );
xor ( n4159 , n3971 , n3973 );
xor ( n4160 , n4159 , n3976 );
and ( n4161 , n4157 , n4160 );
and ( n4162 , n4125 , n4160 );
or ( n4163 , n4158 , n4161 , n4162 );
xor ( n4164 , n3888 , n3892 );
xor ( n4165 , n4164 , n3897 );
xor ( n4166 , n3937 , n3941 );
xor ( n4167 , n4166 , n3946 );
and ( n4168 , n4165 , n4167 );
xor ( n4169 , n3953 , n3957 );
xor ( n4170 , n4169 , n3962 );
and ( n4171 , n4167 , n4170 );
and ( n4172 , n4165 , n4170 );
or ( n4173 , n4168 , n4171 , n4172 );
and ( n4174 , n1666 , n4107 );
and ( n4175 , n1636 , n4105 );
nor ( n4176 , n4174 , n4175 );
xnor ( n4177 , n4176 , n3870 );
and ( n4178 , n1720 , n3367 );
and ( n4179 , n1705 , n3365 );
nor ( n4180 , n4178 , n4179 );
xnor ( n4181 , n4180 , n3306 );
and ( n4182 , n4177 , n4181 );
and ( n4183 , n2295 , n2320 );
and ( n4184 , n2258 , n2318 );
nor ( n4185 , n4183 , n4184 );
xnor ( n4186 , n4185 , n2217 );
and ( n4187 , n4181 , n4186 );
and ( n4188 , n4177 , n4186 );
or ( n4189 , n4182 , n4187 , n4188 );
and ( n4190 , n1675 , n3742 );
and ( n4191 , n1655 , n3740 );
nor ( n4192 , n4190 , n4191 );
xnor ( n4193 , n4192 , n3538 );
and ( n4194 , n1935 , n2887 );
and ( n4195 , n1849 , n2885 );
nor ( n4196 , n4194 , n4195 );
xnor ( n4197 , n4196 , n2801 );
and ( n4198 , n4193 , n4197 );
and ( n4199 , n2897 , n1901 );
and ( n4200 , n2773 , n1899 );
nor ( n4201 , n4199 , n4200 );
xnor ( n4202 , n4201 , n1869 );
and ( n4203 , n4197 , n4202 );
and ( n4204 , n4193 , n4202 );
or ( n4205 , n4198 , n4203 , n4204 );
and ( n4206 , n4189 , n4205 );
and ( n4207 , n1817 , n3093 );
and ( n4208 , n1799 , n3091 );
nor ( n4209 , n4207 , n4208 );
xnor ( n4210 , n4209 , n3027 );
and ( n4211 , n2506 , n2113 );
and ( n4212 , n2390 , n2111 );
nor ( n4213 , n4211 , n4212 );
xnor ( n4214 , n4213 , n2091 );
and ( n4215 , n4210 , n4214 );
and ( n4216 , n2697 , n2020 );
and ( n4217 , n2615 , n2018 );
nor ( n4218 , n4216 , n4217 );
xnor ( n4219 , n4218 , n1981 );
and ( n4220 , n4214 , n4219 );
and ( n4221 , n4210 , n4219 );
or ( n4222 , n4215 , n4220 , n4221 );
and ( n4223 , n4205 , n4222 );
and ( n4224 , n4189 , n4222 );
or ( n4225 , n4206 , n4223 , n4224 );
and ( n4226 , n2181 , n2483 );
and ( n4227 , n2080 , n2481 );
nor ( n4228 , n4226 , n4227 );
xnor ( n4229 , n4228 , n2418 );
and ( n4230 , n4099 , n1663 );
and ( n4231 , n3859 , n1661 );
nor ( n4232 , n4230 , n4231 );
xnor ( n4233 , n4232 , n1671 );
and ( n4234 , n4229 , n4233 );
buf ( n4235 , n1152 );
buf ( n4236 , n4235 );
and ( n4237 , n4236 , n1657 );
and ( n4238 , n4233 , n4237 );
and ( n4239 , n4229 , n4237 );
or ( n4240 , n4234 , n4238 , n4239 );
not ( n4241 , n3867 );
buf ( n4242 , n4241 );
and ( n4243 , n4240 , n4242 );
not ( n4244 , n4110 );
and ( n4245 , n4242 , n4244 );
and ( n4246 , n4240 , n4244 );
or ( n4247 , n4243 , n4245 , n4246 );
and ( n4248 , n4225 , n4247 );
xor ( n4249 , n4103 , n4111 );
xor ( n4250 , n4249 , n4116 );
and ( n4251 , n4247 , n4250 );
and ( n4252 , n4225 , n4250 );
or ( n4253 , n4248 , n4251 , n4252 );
and ( n4254 , n4173 , n4253 );
xor ( n4255 , n3990 , n3992 );
xor ( n4256 , n4255 , n3995 );
and ( n4257 , n4253 , n4256 );
and ( n4258 , n4173 , n4256 );
or ( n4259 , n4254 , n4257 , n4258 );
and ( n4260 , n2042 , n2654 );
and ( n4261 , n2027 , n2652 );
nor ( n4262 , n4260 , n4261 );
xnor ( n4263 , n4262 , n2570 );
and ( n4264 , n3136 , n1807 );
and ( n4265 , n3052 , n1805 );
nor ( n4266 , n4264 , n4265 );
xnor ( n4267 , n4266 , n1756 );
and ( n4268 , n4263 , n4267 );
and ( n4269 , n3466 , n1728 );
and ( n4270 , n3414 , n1726 );
nor ( n4271 , n4269 , n4270 );
xnor ( n4272 , n4271 , n1697 );
and ( n4273 , n4267 , n4272 );
and ( n4274 , n4263 , n4272 );
or ( n4275 , n4268 , n4273 , n4274 );
xor ( n4276 , n4040 , n4044 );
xor ( n4277 , n4276 , n4049 );
and ( n4278 , n4275 , n4277 );
xor ( n4279 , n4129 , n4133 );
xor ( n4280 , n4279 , n4138 );
and ( n4281 , n4277 , n4280 );
and ( n4282 , n4275 , n4280 );
or ( n4283 , n4278 , n4281 , n4282 );
xor ( n4284 , n4092 , n4096 );
xor ( n4285 , n4284 , n4100 );
xor ( n4286 , n4056 , n4060 );
xor ( n4287 , n4286 , n4065 );
and ( n4288 , n4285 , n4287 );
xor ( n4289 , n4073 , n4077 );
xor ( n4290 , n4289 , n4082 );
and ( n4291 , n4287 , n4290 );
and ( n4292 , n4285 , n4290 );
or ( n4293 , n4288 , n4291 , n4292 );
and ( n4294 , n4283 , n4293 );
xor ( n4295 , n4052 , n4068 );
xor ( n4296 , n4295 , n4085 );
and ( n4297 , n4293 , n4296 );
and ( n4298 , n4283 , n4296 );
or ( n4299 , n4294 , n4297 , n4298 );
xor ( n4300 , n4088 , n4119 );
xor ( n4301 , n4300 , n4122 );
and ( n4302 , n4299 , n4301 );
xor ( n4303 , n4149 , n4151 );
xor ( n4304 , n4303 , n4154 );
and ( n4305 , n4301 , n4304 );
and ( n4306 , n4299 , n4304 );
or ( n4307 , n4302 , n4305 , n4306 );
and ( n4308 , n4259 , n4307 );
xor ( n4309 , n3998 , n4000 );
xor ( n4310 , n4309 , n4003 );
and ( n4311 , n4307 , n4310 );
and ( n4312 , n4259 , n4310 );
or ( n4313 , n4308 , n4311 , n4312 );
and ( n4314 , n4163 , n4313 );
and ( n4315 , n4035 , n4314 );
and ( n4316 , n4033 , n4314 );
or ( n4317 , n4036 , n4315 , n4316 );
and ( n4318 , n4031 , n4317 );
and ( n4319 , n4029 , n4317 );
or ( n4320 , n4032 , n4318 , n4319 );
and ( n4321 , n4027 , n4320 );
xor ( n4322 , n4027 , n4320 );
xor ( n4323 , n4029 , n4031 );
xor ( n4324 , n4323 , n4317 );
xor ( n4325 , n3933 , n3979 );
xor ( n4326 , n4325 , n3982 );
xor ( n4327 , n4006 , n4008 );
and ( n4328 , n4326 , n4327 );
xor ( n4329 , n4163 , n4313 );
and ( n4330 , n4327 , n4329 );
and ( n4331 , n4326 , n4329 );
or ( n4332 , n4328 , n4330 , n4331 );
xor ( n4333 , n4033 , n4035 );
xor ( n4334 , n4333 , n4314 );
and ( n4335 , n4332 , n4334 );
and ( n4336 , n2080 , n2654 );
and ( n4337 , n2042 , n2652 );
nor ( n4338 , n4336 , n4337 );
xnor ( n4339 , n4338 , n2570 );
and ( n4340 , n3052 , n1901 );
and ( n4341 , n2897 , n1899 );
nor ( n4342 , n4340 , n4341 );
xnor ( n4343 , n4342 , n1869 );
and ( n4344 , n4339 , n4343 );
and ( n4345 , n3414 , n1807 );
and ( n4346 , n3136 , n1805 );
nor ( n4347 , n4345 , n4346 );
xnor ( n4348 , n4347 , n1756 );
and ( n4349 , n4343 , n4348 );
and ( n4350 , n4339 , n4348 );
or ( n4351 , n4344 , n4349 , n4350 );
and ( n4352 , n1849 , n3093 );
and ( n4353 , n1817 , n3091 );
nor ( n4354 , n4352 , n4353 );
xnor ( n4355 , n4354 , n3027 );
and ( n4356 , n2390 , n2320 );
and ( n4357 , n2295 , n2318 );
nor ( n4358 , n4356 , n4357 );
xnor ( n4359 , n4358 , n2217 );
and ( n4360 , n4355 , n4359 );
and ( n4361 , n2615 , n2113 );
and ( n4362 , n2506 , n2111 );
nor ( n4363 , n4361 , n4362 );
xnor ( n4364 , n4363 , n2091 );
and ( n4365 , n4359 , n4364 );
and ( n4366 , n4355 , n4364 );
or ( n4367 , n4360 , n4365 , n4366 );
and ( n4368 , n4351 , n4367 );
and ( n4369 , n1799 , n3367 );
and ( n4370 , n1720 , n3365 );
nor ( n4371 , n4369 , n4370 );
xnor ( n4372 , n4371 , n3306 );
and ( n4373 , n2258 , n2483 );
and ( n4374 , n2181 , n2481 );
nor ( n4375 , n4373 , n4374 );
xnor ( n4376 , n4375 , n2418 );
and ( n4377 , n4372 , n4376 );
and ( n4378 , n4236 , n1663 );
and ( n4379 , n4099 , n1661 );
nor ( n4380 , n4378 , n4379 );
xnor ( n4381 , n4380 , n1671 );
and ( n4382 , n4376 , n4381 );
and ( n4383 , n4372 , n4381 );
or ( n4384 , n4377 , n4382 , n4383 );
and ( n4385 , n4367 , n4384 );
and ( n4386 , n4351 , n4384 );
or ( n4387 , n4368 , n4385 , n4386 );
buf ( n4388 , n1185 );
buf ( n4389 , n4388 );
xor ( n4390 , n3867 , n4389 );
not ( n4391 , n4389 );
and ( n4392 , n4390 , n4391 );
and ( n4393 , n1636 , n4392 );
not ( n4394 , n4393 );
xnor ( n4395 , n4394 , n3867 );
and ( n4396 , n1655 , n4107 );
and ( n4397 , n1666 , n4105 );
nor ( n4398 , n4396 , n4397 );
xnor ( n4399 , n4398 , n3870 );
and ( n4400 , n4395 , n4399 );
buf ( n4401 , n1153 );
buf ( n4402 , n4401 );
and ( n4403 , n4402 , n1657 );
and ( n4404 , n4399 , n4403 );
and ( n4405 , n4395 , n4403 );
or ( n4406 , n4400 , n4404 , n4405 );
and ( n4407 , n4406 , n3867 );
and ( n4408 , n3911 , n1646 );
and ( n4409 , n3813 , n1644 );
nor ( n4410 , n4408 , n4409 );
xnor ( n4411 , n4410 , n1651 );
and ( n4412 , n3867 , n4411 );
and ( n4413 , n4406 , n4411 );
or ( n4414 , n4407 , n4412 , n4413 );
and ( n4415 , n4387 , n4414 );
xor ( n4416 , n4189 , n4205 );
xor ( n4417 , n4416 , n4222 );
and ( n4418 , n4414 , n4417 );
and ( n4419 , n4387 , n4417 );
or ( n4420 , n4415 , n4418 , n4419 );
and ( n4421 , n1705 , n3742 );
and ( n4422 , n1675 , n3740 );
nor ( n4423 , n4421 , n4422 );
xnor ( n4424 , n4423 , n3538 );
and ( n4425 , n2027 , n2887 );
and ( n4426 , n1935 , n2885 );
nor ( n4427 , n4425 , n4426 );
xnor ( n4428 , n4427 , n2801 );
and ( n4429 , n4424 , n4428 );
and ( n4430 , n2773 , n2020 );
and ( n4431 , n2697 , n2018 );
nor ( n4432 , n4430 , n4431 );
xnor ( n4433 , n4432 , n1981 );
and ( n4434 , n4428 , n4433 );
and ( n4435 , n4424 , n4433 );
or ( n4436 , n4429 , n4434 , n4435 );
xor ( n4437 , n4229 , n4233 );
xor ( n4438 , n4437 , n4237 );
and ( n4439 , n4436 , n4438 );
xor ( n4440 , n4263 , n4267 );
xor ( n4441 , n4440 , n4272 );
and ( n4442 , n4438 , n4441 );
and ( n4443 , n4436 , n4441 );
or ( n4444 , n4439 , n4442 , n4443 );
xor ( n4445 , n4177 , n4181 );
xor ( n4446 , n4445 , n4186 );
xor ( n4447 , n4193 , n4197 );
xor ( n4448 , n4447 , n4202 );
and ( n4449 , n4446 , n4448 );
xor ( n4450 , n4210 , n4214 );
xor ( n4451 , n4450 , n4219 );
and ( n4452 , n4448 , n4451 );
and ( n4453 , n4446 , n4451 );
or ( n4454 , n4449 , n4452 , n4453 );
and ( n4455 , n4444 , n4454 );
xor ( n4456 , n4240 , n4242 );
xor ( n4457 , n4456 , n4244 );
and ( n4458 , n4454 , n4457 );
and ( n4459 , n4444 , n4457 );
or ( n4460 , n4455 , n4458 , n4459 );
and ( n4461 , n4420 , n4460 );
xor ( n4462 , n4283 , n4293 );
xor ( n4463 , n4462 , n4296 );
and ( n4464 , n4460 , n4463 );
and ( n4465 , n4420 , n4463 );
or ( n4466 , n4461 , n4464 , n4465 );
xor ( n4467 , n4141 , n4143 );
xor ( n4468 , n4467 , n4146 );
xor ( n4469 , n4165 , n4167 );
xor ( n4470 , n4469 , n4170 );
and ( n4471 , n4468 , n4470 );
xor ( n4472 , n4225 , n4247 );
xor ( n4473 , n4472 , n4250 );
and ( n4474 , n4470 , n4473 );
and ( n4475 , n4468 , n4473 );
or ( n4476 , n4471 , n4474 , n4475 );
and ( n4477 , n4466 , n4476 );
xor ( n4478 , n4173 , n4253 );
xor ( n4479 , n4478 , n4256 );
and ( n4480 , n4476 , n4479 );
and ( n4481 , n4466 , n4479 );
or ( n4482 , n4477 , n4480 , n4481 );
xor ( n4483 , n4125 , n4157 );
xor ( n4484 , n4483 , n4160 );
and ( n4485 , n4482 , n4484 );
xor ( n4486 , n4259 , n4307 );
xor ( n4487 , n4486 , n4310 );
and ( n4488 , n4484 , n4487 );
and ( n4489 , n4482 , n4487 );
or ( n4490 , n4485 , n4488 , n4489 );
xor ( n4491 , n4326 , n4327 );
xor ( n4492 , n4491 , n4329 );
and ( n4493 , n4490 , n4492 );
xor ( n4494 , n4482 , n4484 );
xor ( n4495 , n4494 , n4487 );
xor ( n4496 , n4339 , n4343 );
xor ( n4497 , n4496 , n4348 );
xor ( n4498 , n4424 , n4428 );
xor ( n4499 , n4498 , n4433 );
and ( n4500 , n4497 , n4499 );
xor ( n4501 , n4355 , n4359 );
xor ( n4502 , n4501 , n4364 );
and ( n4503 , n4499 , n4502 );
and ( n4504 , n4497 , n4502 );
or ( n4505 , n4500 , n4503 , n4504 );
xor ( n4506 , n4351 , n4367 );
xor ( n4507 , n4506 , n4384 );
and ( n4508 , n4505 , n4507 );
xor ( n4509 , n4406 , n3867 );
xor ( n4510 , n4509 , n4411 );
and ( n4511 , n4507 , n4510 );
and ( n4512 , n4505 , n4510 );
or ( n4513 , n4508 , n4511 , n4512 );
xor ( n4514 , n4275 , n4277 );
xor ( n4515 , n4514 , n4280 );
and ( n4516 , n4513 , n4515 );
xor ( n4517 , n4285 , n4287 );
xor ( n4518 , n4517 , n4290 );
and ( n4519 , n4515 , n4518 );
and ( n4520 , n4513 , n4518 );
or ( n4521 , n4516 , n4519 , n4520 );
and ( n4522 , n1720 , n3742 );
and ( n4523 , n1705 , n3740 );
nor ( n4524 , n4522 , n4523 );
xnor ( n4525 , n4524 , n3538 );
and ( n4526 , n2697 , n2113 );
and ( n4527 , n2615 , n2111 );
nor ( n4528 , n4526 , n4527 );
xnor ( n4529 , n4528 , n2091 );
and ( n4530 , n4525 , n4529 );
and ( n4531 , n2897 , n2020 );
and ( n4532 , n2773 , n2018 );
nor ( n4533 , n4531 , n4532 );
xnor ( n4534 , n4533 , n1981 );
and ( n4535 , n4529 , n4534 );
and ( n4536 , n4525 , n4534 );
or ( n4537 , n4530 , n4535 , n4536 );
and ( n4538 , n1675 , n4107 );
and ( n4539 , n1655 , n4105 );
nor ( n4540 , n4538 , n4539 );
xnor ( n4541 , n4540 , n3870 );
and ( n4542 , n1817 , n3367 );
and ( n4543 , n1799 , n3365 );
nor ( n4544 , n4542 , n4543 );
xnor ( n4545 , n4544 , n3306 );
and ( n4546 , n4541 , n4545 );
and ( n4547 , n4402 , n1663 );
and ( n4548 , n4236 , n1661 );
nor ( n4549 , n4547 , n4548 );
xnor ( n4550 , n4549 , n1671 );
and ( n4551 , n4545 , n4550 );
and ( n4552 , n4541 , n4550 );
or ( n4553 , n4546 , n4551 , n4552 );
and ( n4554 , n4537 , n4553 );
and ( n4555 , n1935 , n3093 );
and ( n4556 , n1849 , n3091 );
nor ( n4557 , n4555 , n4556 );
xnor ( n4558 , n4557 , n3027 );
and ( n4559 , n2295 , n2483 );
and ( n4560 , n2258 , n2481 );
nor ( n4561 , n4559 , n4560 );
xnor ( n4562 , n4561 , n2418 );
and ( n4563 , n4558 , n4562 );
and ( n4564 , n2506 , n2320 );
and ( n4565 , n2390 , n2318 );
nor ( n4566 , n4564 , n4565 );
xnor ( n4567 , n4566 , n2217 );
and ( n4568 , n4562 , n4567 );
and ( n4569 , n4558 , n4567 );
or ( n4570 , n4563 , n4568 , n4569 );
and ( n4571 , n4553 , n4570 );
and ( n4572 , n4537 , n4570 );
or ( n4573 , n4554 , n4571 , n4572 );
and ( n4574 , n1666 , n4392 );
and ( n4575 , n1636 , n4389 );
nor ( n4576 , n4574 , n4575 );
xnor ( n4577 , n4576 , n3867 );
and ( n4578 , n4402 , n1661 );
not ( n4579 , n4578 );
and ( n4580 , n4579 , n1671 );
and ( n4581 , n4577 , n4580 );
and ( n4582 , n3813 , n1728 );
and ( n4583 , n3466 , n1726 );
nor ( n4584 , n4582 , n4583 );
xnor ( n4585 , n4584 , n1697 );
and ( n4586 , n4581 , n4585 );
and ( n4587 , n3859 , n1646 );
and ( n4588 , n3911 , n1644 );
nor ( n4589 , n4587 , n4588 );
xnor ( n4590 , n4589 , n1651 );
and ( n4591 , n4585 , n4590 );
and ( n4592 , n4581 , n4590 );
or ( n4593 , n4586 , n4591 , n4592 );
and ( n4594 , n4573 , n4593 );
and ( n4595 , n2042 , n2887 );
and ( n4596 , n2027 , n2885 );
nor ( n4597 , n4595 , n4596 );
xnor ( n4598 , n4597 , n2801 );
and ( n4599 , n3136 , n1901 );
and ( n4600 , n3052 , n1899 );
nor ( n4601 , n4599 , n4600 );
xnor ( n4602 , n4601 , n1869 );
and ( n4603 , n4598 , n4602 );
and ( n4604 , n3466 , n1807 );
and ( n4605 , n3414 , n1805 );
nor ( n4606 , n4604 , n4605 );
xnor ( n4607 , n4606 , n1756 );
and ( n4608 , n4602 , n4607 );
and ( n4609 , n4598 , n4607 );
or ( n4610 , n4603 , n4608 , n4609 );
and ( n4611 , n2181 , n2654 );
and ( n4612 , n2080 , n2652 );
nor ( n4613 , n4611 , n4612 );
xnor ( n4614 , n4613 , n2570 );
and ( n4615 , n3911 , n1728 );
and ( n4616 , n3813 , n1726 );
nor ( n4617 , n4615 , n4616 );
xnor ( n4618 , n4617 , n1697 );
and ( n4619 , n4614 , n4618 );
and ( n4620 , n4099 , n1646 );
and ( n4621 , n3859 , n1644 );
nor ( n4622 , n4620 , n4621 );
xnor ( n4623 , n4622 , n1651 );
and ( n4624 , n4618 , n4623 );
and ( n4625 , n4614 , n4623 );
or ( n4626 , n4619 , n4624 , n4625 );
and ( n4627 , n4610 , n4626 );
xor ( n4628 , n4395 , n4399 );
xor ( n4629 , n4628 , n4403 );
and ( n4630 , n4626 , n4629 );
and ( n4631 , n4610 , n4629 );
or ( n4632 , n4627 , n4630 , n4631 );
and ( n4633 , n4593 , n4632 );
and ( n4634 , n4573 , n4632 );
or ( n4635 , n4594 , n4633 , n4634 );
xor ( n4636 , n4387 , n4414 );
xor ( n4637 , n4636 , n4417 );
and ( n4638 , n4635 , n4637 );
xor ( n4639 , n4444 , n4454 );
xor ( n4640 , n4639 , n4457 );
and ( n4641 , n4637 , n4640 );
and ( n4642 , n4635 , n4640 );
or ( n4643 , n4638 , n4641 , n4642 );
and ( n4644 , n4521 , n4643 );
xor ( n4645 , n4468 , n4470 );
xor ( n4646 , n4645 , n4473 );
and ( n4647 , n4643 , n4646 );
and ( n4648 , n4521 , n4646 );
or ( n4649 , n4644 , n4647 , n4648 );
xor ( n4650 , n4299 , n4301 );
xor ( n4651 , n4650 , n4304 );
and ( n4652 , n4649 , n4651 );
xor ( n4653 , n4466 , n4476 );
xor ( n4654 , n4653 , n4479 );
and ( n4655 , n4651 , n4654 );
and ( n4656 , n4649 , n4654 );
or ( n4657 , n4652 , n4655 , n4656 );
and ( n4658 , n4495 , n4657 );
xor ( n4659 , n4649 , n4651 );
xor ( n4660 , n4659 , n4654 );
xor ( n4661 , n4420 , n4460 );
xor ( n4662 , n4661 , n4463 );
and ( n4663 , n1799 , n3742 );
and ( n4664 , n1720 , n3740 );
nor ( n4665 , n4663 , n4664 );
xnor ( n4666 , n4665 , n3538 );
and ( n4667 , n2080 , n2887 );
and ( n4668 , n2042 , n2885 );
nor ( n4669 , n4667 , n4668 );
xnor ( n4670 , n4669 , n2801 );
and ( n4671 , n4666 , n4670 );
and ( n4672 , n3414 , n1901 );
and ( n4673 , n3136 , n1899 );
nor ( n4674 , n4672 , n4673 );
xnor ( n4675 , n4674 , n1869 );
and ( n4676 , n4670 , n4675 );
and ( n4677 , n4666 , n4675 );
or ( n4678 , n4671 , n4676 , n4677 );
and ( n4679 , n2258 , n2654 );
and ( n4680 , n2181 , n2652 );
nor ( n4681 , n4679 , n4680 );
xnor ( n4682 , n4681 , n2570 );
and ( n4683 , n3813 , n1807 );
and ( n4684 , n3466 , n1805 );
nor ( n4685 , n4683 , n4684 );
xnor ( n4686 , n4685 , n1756 );
and ( n4687 , n4682 , n4686 );
and ( n4688 , n3859 , n1728 );
and ( n4689 , n3911 , n1726 );
nor ( n4690 , n4688 , n4689 );
xnor ( n4691 , n4690 , n1697 );
and ( n4692 , n4686 , n4691 );
and ( n4693 , n4682 , n4691 );
or ( n4694 , n4687 , n4692 , n4693 );
and ( n4695 , n4678 , n4694 );
and ( n4696 , n2027 , n3093 );
and ( n4697 , n1935 , n3091 );
nor ( n4698 , n4696 , n4697 );
xnor ( n4699 , n4698 , n3027 );
and ( n4700 , n2773 , n2113 );
and ( n4701 , n2697 , n2111 );
nor ( n4702 , n4700 , n4701 );
xnor ( n4703 , n4702 , n2091 );
and ( n4704 , n4699 , n4703 );
and ( n4705 , n3052 , n2020 );
and ( n4706 , n2897 , n2018 );
nor ( n4707 , n4705 , n4706 );
xnor ( n4708 , n4707 , n1981 );
and ( n4709 , n4703 , n4708 );
and ( n4710 , n4699 , n4708 );
or ( n4711 , n4704 , n4709 , n4710 );
and ( n4712 , n4694 , n4711 );
and ( n4713 , n4678 , n4711 );
or ( n4714 , n4695 , n4712 , n4713 );
xor ( n4715 , n4372 , n4376 );
xor ( n4716 , n4715 , n4381 );
and ( n4717 , n4714 , n4716 );
xor ( n4718 , n4581 , n4585 );
xor ( n4719 , n4718 , n4590 );
and ( n4720 , n4716 , n4719 );
and ( n4721 , n4714 , n4719 );
or ( n4722 , n4717 , n4720 , n4721 );
xor ( n4723 , n4436 , n4438 );
xor ( n4724 , n4723 , n4441 );
and ( n4725 , n4722 , n4724 );
xor ( n4726 , n4446 , n4448 );
xor ( n4727 , n4726 , n4451 );
and ( n4728 , n4724 , n4727 );
and ( n4729 , n4722 , n4727 );
or ( n4730 , n4725 , n4728 , n4729 );
xor ( n4731 , n4577 , n4580 );
and ( n4732 , n1655 , n4392 );
and ( n4733 , n1666 , n4389 );
nor ( n4734 , n4732 , n4733 );
xnor ( n4735 , n4734 , n3867 );
and ( n4736 , n1705 , n4107 );
and ( n4737 , n1675 , n4105 );
nor ( n4738 , n4736 , n4737 );
xnor ( n4739 , n4738 , n3870 );
and ( n4740 , n4735 , n4739 );
and ( n4741 , n4739 , n4578 );
and ( n4742 , n4735 , n4578 );
or ( n4743 , n4740 , n4741 , n4742 );
and ( n4744 , n4731 , n4743 );
and ( n4745 , n1849 , n3367 );
and ( n4746 , n1817 , n3365 );
nor ( n4747 , n4745 , n4746 );
xnor ( n4748 , n4747 , n3306 );
and ( n4749 , n2390 , n2483 );
and ( n4750 , n2295 , n2481 );
nor ( n4751 , n4749 , n4750 );
xnor ( n4752 , n4751 , n2418 );
and ( n4753 , n4748 , n4752 );
and ( n4754 , n2615 , n2320 );
and ( n4755 , n2506 , n2318 );
nor ( n4756 , n4754 , n4755 );
xnor ( n4757 , n4756 , n2217 );
and ( n4758 , n4752 , n4757 );
and ( n4759 , n4748 , n4757 );
or ( n4760 , n4753 , n4758 , n4759 );
and ( n4761 , n4743 , n4760 );
and ( n4762 , n4731 , n4760 );
or ( n4763 , n4744 , n4761 , n4762 );
xor ( n4764 , n4614 , n4618 );
xor ( n4765 , n4764 , n4623 );
xor ( n4766 , n4541 , n4545 );
xor ( n4767 , n4766 , n4550 );
and ( n4768 , n4765 , n4767 );
xor ( n4769 , n4558 , n4562 );
xor ( n4770 , n4769 , n4567 );
and ( n4771 , n4767 , n4770 );
and ( n4772 , n4765 , n4770 );
or ( n4773 , n4768 , n4771 , n4772 );
and ( n4774 , n4763 , n4773 );
xor ( n4775 , n4610 , n4626 );
xor ( n4776 , n4775 , n4629 );
and ( n4777 , n4773 , n4776 );
and ( n4778 , n4763 , n4776 );
or ( n4779 , n4774 , n4777 , n4778 );
xor ( n4780 , n4573 , n4593 );
xor ( n4781 , n4780 , n4632 );
and ( n4782 , n4779 , n4781 );
xor ( n4783 , n4505 , n4507 );
xor ( n4784 , n4783 , n4510 );
and ( n4785 , n4781 , n4784 );
and ( n4786 , n4779 , n4784 );
or ( n4787 , n4782 , n4785 , n4786 );
and ( n4788 , n4730 , n4787 );
xor ( n4789 , n4513 , n4515 );
xor ( n4790 , n4789 , n4518 );
and ( n4791 , n4787 , n4790 );
and ( n4792 , n4730 , n4790 );
or ( n4793 , n4788 , n4791 , n4792 );
and ( n4794 , n4662 , n4793 );
xor ( n4795 , n4521 , n4643 );
xor ( n4796 , n4795 , n4646 );
and ( n4797 , n4793 , n4796 );
and ( n4798 , n4662 , n4796 );
or ( n4799 , n4794 , n4797 , n4798 );
and ( n4800 , n4660 , n4799 );
and ( n4801 , n1817 , n3742 );
and ( n4802 , n1799 , n3740 );
nor ( n4803 , n4801 , n4802 );
xnor ( n4804 , n4803 , n3538 );
and ( n4805 , n2181 , n2887 );
and ( n4806 , n2080 , n2885 );
nor ( n4807 , n4805 , n4806 );
xnor ( n4808 , n4807 , n2801 );
and ( n4809 , n4804 , n4808 );
and ( n4810 , n3136 , n2020 );
and ( n4811 , n3052 , n2018 );
nor ( n4812 , n4810 , n4811 );
xnor ( n4813 , n4812 , n1981 );
and ( n4814 , n4808 , n4813 );
and ( n4815 , n4804 , n4813 );
or ( n4816 , n4809 , n4814 , n4815 );
and ( n4817 , n2295 , n2654 );
and ( n4818 , n2258 , n2652 );
nor ( n4819 , n4817 , n4818 );
xnor ( n4820 , n4819 , n2570 );
and ( n4821 , n3466 , n1901 );
and ( n4822 , n3414 , n1899 );
nor ( n4823 , n4821 , n4822 );
xnor ( n4824 , n4823 , n1869 );
and ( n4825 , n4820 , n4824 );
and ( n4826 , n3911 , n1807 );
and ( n4827 , n3813 , n1805 );
nor ( n4828 , n4826 , n4827 );
xnor ( n4829 , n4828 , n1756 );
and ( n4830 , n4824 , n4829 );
and ( n4831 , n4820 , n4829 );
or ( n4832 , n4825 , n4830 , n4831 );
and ( n4833 , n4816 , n4832 );
and ( n4834 , n2042 , n3093 );
and ( n4835 , n2027 , n3091 );
nor ( n4836 , n4834 , n4835 );
xnor ( n4837 , n4836 , n3027 );
and ( n4838 , n2697 , n2320 );
and ( n4839 , n2615 , n2318 );
nor ( n4840 , n4838 , n4839 );
xnor ( n4841 , n4840 , n2217 );
and ( n4842 , n4837 , n4841 );
and ( n4843 , n2897 , n2113 );
and ( n4844 , n2773 , n2111 );
nor ( n4845 , n4843 , n4844 );
xnor ( n4846 , n4845 , n2091 );
and ( n4847 , n4841 , n4846 );
and ( n4848 , n4837 , n4846 );
or ( n4849 , n4842 , n4847 , n4848 );
and ( n4850 , n4832 , n4849 );
and ( n4851 , n4816 , n4849 );
or ( n4852 , n4833 , n4850 , n4851 );
xor ( n4853 , n4525 , n4529 );
xor ( n4854 , n4853 , n4534 );
and ( n4855 , n4852 , n4854 );
xor ( n4856 , n4598 , n4602 );
xor ( n4857 , n4856 , n4607 );
and ( n4858 , n4854 , n4857 );
and ( n4859 , n4852 , n4857 );
or ( n4860 , n4855 , n4858 , n4859 );
xor ( n4861 , n4537 , n4553 );
xor ( n4862 , n4861 , n4570 );
and ( n4863 , n4860 , n4862 );
xor ( n4864 , n4497 , n4499 );
xor ( n4865 , n4864 , n4502 );
and ( n4866 , n4862 , n4865 );
and ( n4867 , n4860 , n4865 );
or ( n4868 , n4863 , n4866 , n4867 );
and ( n4869 , n1720 , n4107 );
and ( n4870 , n1705 , n4105 );
nor ( n4871 , n4869 , n4870 );
xnor ( n4872 , n4871 , n3870 );
and ( n4873 , n1935 , n3367 );
and ( n4874 , n1849 , n3365 );
nor ( n4875 , n4873 , n4874 );
xnor ( n4876 , n4875 , n3306 );
and ( n4877 , n4872 , n4876 );
and ( n4878 , n2506 , n2483 );
and ( n4879 , n2390 , n2481 );
nor ( n4880 , n4878 , n4879 );
xnor ( n4881 , n4880 , n2418 );
and ( n4882 , n4876 , n4881 );
and ( n4883 , n4872 , n4881 );
or ( n4884 , n4877 , n4882 , n4883 );
and ( n4885 , n1675 , n4392 );
and ( n4886 , n1655 , n4389 );
nor ( n4887 , n4885 , n4886 );
xnor ( n4888 , n4887 , n3867 );
and ( n4889 , n4402 , n1644 );
not ( n4890 , n4889 );
and ( n4891 , n4890 , n1651 );
and ( n4892 , n4888 , n4891 );
and ( n4893 , n4884 , n4892 );
and ( n4894 , n4236 , n1646 );
and ( n4895 , n4099 , n1644 );
nor ( n4896 , n4894 , n4895 );
xnor ( n4897 , n4896 , n1651 );
and ( n4898 , n4892 , n4897 );
and ( n4899 , n4884 , n4897 );
or ( n4900 , n4893 , n4898 , n4899 );
xor ( n4901 , n4678 , n4694 );
xor ( n4902 , n4901 , n4711 );
and ( n4903 , n4900 , n4902 );
xor ( n4904 , n4731 , n4743 );
xor ( n4905 , n4904 , n4760 );
and ( n4906 , n4902 , n4905 );
and ( n4907 , n4900 , n4905 );
or ( n4908 , n4903 , n4906 , n4907 );
xor ( n4909 , n4666 , n4670 );
xor ( n4910 , n4909 , n4675 );
xor ( n4911 , n4735 , n4739 );
xor ( n4912 , n4911 , n4578 );
and ( n4913 , n4910 , n4912 );
xor ( n4914 , n4682 , n4686 );
xor ( n4915 , n4914 , n4691 );
and ( n4916 , n4912 , n4915 );
and ( n4917 , n4910 , n4915 );
or ( n4918 , n4913 , n4916 , n4917 );
xor ( n4919 , n4888 , n4891 );
and ( n4920 , n4099 , n1728 );
and ( n4921 , n3859 , n1726 );
nor ( n4922 , n4920 , n4921 );
xnor ( n4923 , n4922 , n1697 );
and ( n4924 , n4919 , n4923 );
and ( n4925 , n4402 , n1646 );
and ( n4926 , n4236 , n1644 );
nor ( n4927 , n4925 , n4926 );
xnor ( n4928 , n4927 , n1651 );
and ( n4929 , n4923 , n4928 );
and ( n4930 , n4919 , n4928 );
or ( n4931 , n4924 , n4929 , n4930 );
xor ( n4932 , n4748 , n4752 );
xor ( n4933 , n4932 , n4757 );
and ( n4934 , n4931 , n4933 );
xor ( n4935 , n4699 , n4703 );
xor ( n4936 , n4935 , n4708 );
and ( n4937 , n4933 , n4936 );
and ( n4938 , n4931 , n4936 );
or ( n4939 , n4934 , n4937 , n4938 );
and ( n4940 , n4918 , n4939 );
xor ( n4941 , n4765 , n4767 );
xor ( n4942 , n4941 , n4770 );
and ( n4943 , n4939 , n4942 );
and ( n4944 , n4918 , n4942 );
or ( n4945 , n4940 , n4943 , n4944 );
and ( n4946 , n4908 , n4945 );
xor ( n4947 , n4714 , n4716 );
xor ( n4948 , n4947 , n4719 );
and ( n4949 , n4945 , n4948 );
and ( n4950 , n4908 , n4948 );
or ( n4951 , n4946 , n4949 , n4950 );
and ( n4952 , n4868 , n4951 );
xor ( n4953 , n4722 , n4724 );
xor ( n4954 , n4953 , n4727 );
and ( n4955 , n4951 , n4954 );
and ( n4956 , n4868 , n4954 );
or ( n4957 , n4952 , n4955 , n4956 );
xor ( n4958 , n4635 , n4637 );
xor ( n4959 , n4958 , n4640 );
and ( n4960 , n4957 , n4959 );
xor ( n4961 , n4730 , n4787 );
xor ( n4962 , n4961 , n4790 );
and ( n4963 , n4959 , n4962 );
and ( n4964 , n4957 , n4962 );
or ( n4965 , n4960 , n4963 , n4964 );
xor ( n4966 , n4662 , n4793 );
xor ( n4967 , n4966 , n4796 );
and ( n4968 , n4965 , n4967 );
xor ( n4969 , n4957 , n4959 );
xor ( n4970 , n4969 , n4962 );
xor ( n4971 , n4763 , n4773 );
xor ( n4972 , n4971 , n4776 );
xor ( n4973 , n4860 , n4862 );
xor ( n4974 , n4973 , n4865 );
and ( n4975 , n4972 , n4974 );
xor ( n4976 , n4908 , n4945 );
xor ( n4977 , n4976 , n4948 );
and ( n4978 , n4974 , n4977 );
and ( n4979 , n4972 , n4977 );
or ( n4980 , n4975 , n4978 , n4979 );
xor ( n4981 , n4779 , n4781 );
xor ( n4982 , n4981 , n4784 );
and ( n4983 , n4980 , n4982 );
xor ( n4984 , n4868 , n4951 );
xor ( n4985 , n4984 , n4954 );
and ( n4986 , n4982 , n4985 );
and ( n4987 , n4980 , n4985 );
or ( n4988 , n4983 , n4986 , n4987 );
and ( n4989 , n4970 , n4988 );
xor ( n4990 , n4980 , n4982 );
xor ( n4991 , n4990 , n4985 );
and ( n4992 , n1799 , n4107 );
and ( n4993 , n1720 , n4105 );
nor ( n4994 , n4992 , n4993 );
xnor ( n4995 , n4994 , n3870 );
and ( n4996 , n2027 , n3367 );
and ( n4997 , n1935 , n3365 );
nor ( n4998 , n4996 , n4997 );
xnor ( n4999 , n4998 , n3306 );
and ( n5000 , n4995 , n4999 );
and ( n5001 , n4999 , n4889 );
and ( n5002 , n4995 , n4889 );
or ( n5003 , n5000 , n5001 , n5002 );
and ( n5004 , n1705 , n4392 );
and ( n5005 , n1675 , n4389 );
nor ( n5006 , n5004 , n5005 );
xnor ( n5007 , n5006 , n3867 );
and ( n5008 , n3052 , n2113 );
and ( n5009 , n2897 , n2111 );
nor ( n5010 , n5008 , n5009 );
xnor ( n5011 , n5010 , n2091 );
and ( n5012 , n5007 , n5011 );
and ( n5013 , n3414 , n2020 );
and ( n5014 , n3136 , n2018 );
nor ( n5015 , n5013 , n5014 );
xnor ( n5016 , n5015 , n1981 );
and ( n5017 , n5011 , n5016 );
and ( n5018 , n5007 , n5016 );
or ( n5019 , n5012 , n5017 , n5018 );
and ( n5020 , n5003 , n5019 );
and ( n5021 , n2080 , n3093 );
and ( n5022 , n2042 , n3091 );
nor ( n5023 , n5021 , n5022 );
xnor ( n5024 , n5023 , n3027 );
and ( n5025 , n2615 , n2483 );
and ( n5026 , n2506 , n2481 );
nor ( n5027 , n5025 , n5026 );
xnor ( n5028 , n5027 , n2418 );
and ( n5029 , n5024 , n5028 );
and ( n5030 , n2773 , n2320 );
and ( n5031 , n2697 , n2318 );
nor ( n5032 , n5030 , n5031 );
xnor ( n5033 , n5032 , n2217 );
and ( n5034 , n5028 , n5033 );
and ( n5035 , n5024 , n5033 );
or ( n5036 , n5029 , n5034 , n5035 );
and ( n5037 , n5019 , n5036 );
and ( n5038 , n5003 , n5036 );
or ( n5039 , n5020 , n5037 , n5038 );
xor ( n5040 , n4804 , n4808 );
xor ( n5041 , n5040 , n4813 );
xor ( n5042 , n4820 , n4824 );
xor ( n5043 , n5042 , n4829 );
and ( n5044 , n5041 , n5043 );
xor ( n5045 , n4837 , n4841 );
xor ( n5046 , n5045 , n4846 );
and ( n5047 , n5043 , n5046 );
and ( n5048 , n5041 , n5046 );
or ( n5049 , n5044 , n5047 , n5048 );
and ( n5050 , n5039 , n5049 );
xor ( n5051 , n4884 , n4892 );
xor ( n5052 , n5051 , n4897 );
and ( n5053 , n5049 , n5052 );
and ( n5054 , n5039 , n5052 );
or ( n5055 , n5050 , n5053 , n5054 );
and ( n5056 , n1849 , n3742 );
and ( n5057 , n1817 , n3740 );
nor ( n5058 , n5056 , n5057 );
xnor ( n5059 , n5058 , n3538 );
and ( n5060 , n2390 , n2654 );
and ( n5061 , n2295 , n2652 );
nor ( n5062 , n5060 , n5061 );
xnor ( n5063 , n5062 , n2570 );
and ( n5064 , n5059 , n5063 );
and ( n5065 , n4236 , n1728 );
and ( n5066 , n4099 , n1726 );
nor ( n5067 , n5065 , n5066 );
xnor ( n5068 , n5067 , n1697 );
and ( n5069 , n5063 , n5068 );
and ( n5070 , n5059 , n5068 );
or ( n5071 , n5064 , n5069 , n5070 );
and ( n5072 , n2258 , n2887 );
and ( n5073 , n2181 , n2885 );
nor ( n5074 , n5072 , n5073 );
xnor ( n5075 , n5074 , n2801 );
and ( n5076 , n3813 , n1901 );
and ( n5077 , n3466 , n1899 );
nor ( n5078 , n5076 , n5077 );
xnor ( n5079 , n5078 , n1869 );
and ( n5080 , n5075 , n5079 );
and ( n5081 , n3859 , n1807 );
and ( n5082 , n3911 , n1805 );
nor ( n5083 , n5081 , n5082 );
xnor ( n5084 , n5083 , n1756 );
and ( n5085 , n5079 , n5084 );
and ( n5086 , n5075 , n5084 );
or ( n5087 , n5080 , n5085 , n5086 );
and ( n5088 , n5071 , n5087 );
xor ( n5089 , n4872 , n4876 );
xor ( n5090 , n5089 , n4881 );
and ( n5091 , n5087 , n5090 );
and ( n5092 , n5071 , n5090 );
or ( n5093 , n5088 , n5091 , n5092 );
xor ( n5094 , n4816 , n4832 );
xor ( n5095 , n5094 , n4849 );
and ( n5096 , n5093 , n5095 );
xor ( n5097 , n4931 , n4933 );
xor ( n5098 , n5097 , n4936 );
and ( n5099 , n5095 , n5098 );
and ( n5100 , n5093 , n5098 );
or ( n5101 , n5096 , n5099 , n5100 );
and ( n5102 , n5055 , n5101 );
xor ( n5103 , n4852 , n4854 );
xor ( n5104 , n5103 , n4857 );
and ( n5105 , n5101 , n5104 );
and ( n5106 , n5055 , n5104 );
or ( n5107 , n5102 , n5105 , n5106 );
and ( n5108 , n2042 , n3367 );
and ( n5109 , n2027 , n3365 );
nor ( n5110 , n5108 , n5109 );
xnor ( n5111 , n5110 , n3306 );
and ( n5112 , n2697 , n2483 );
and ( n5113 , n2615 , n2481 );
nor ( n5114 , n5112 , n5113 );
xnor ( n5115 , n5114 , n2418 );
and ( n5116 , n5111 , n5115 );
and ( n5117 , n2897 , n2320 );
and ( n5118 , n2773 , n2318 );
nor ( n5119 , n5117 , n5118 );
xnor ( n5120 , n5119 , n2217 );
and ( n5121 , n5115 , n5120 );
and ( n5122 , n5111 , n5120 );
or ( n5123 , n5116 , n5121 , n5122 );
and ( n5124 , n2181 , n3093 );
and ( n5125 , n2080 , n3091 );
nor ( n5126 , n5124 , n5125 );
xnor ( n5127 , n5126 , n3027 );
and ( n5128 , n3136 , n2113 );
and ( n5129 , n3052 , n2111 );
nor ( n5130 , n5128 , n5129 );
xnor ( n5131 , n5130 , n2091 );
and ( n5132 , n5127 , n5131 );
and ( n5133 , n3466 , n2020 );
and ( n5134 , n3414 , n2018 );
nor ( n5135 , n5133 , n5134 );
xnor ( n5136 , n5135 , n1981 );
and ( n5137 , n5131 , n5136 );
and ( n5138 , n5127 , n5136 );
or ( n5139 , n5132 , n5137 , n5138 );
and ( n5140 , n5123 , n5139 );
and ( n5141 , n1817 , n4107 );
and ( n5142 , n1799 , n4105 );
nor ( n5143 , n5141 , n5142 );
xnor ( n5144 , n5143 , n3870 );
and ( n5145 , n4402 , n1726 );
not ( n5146 , n5145 );
and ( n5147 , n5146 , n1697 );
and ( n5148 , n5144 , n5147 );
and ( n5149 , n5139 , n5148 );
and ( n5150 , n5123 , n5148 );
or ( n5151 , n5140 , n5149 , n5150 );
xor ( n5152 , n4995 , n4999 );
xor ( n5153 , n5152 , n4889 );
xor ( n5154 , n5059 , n5063 );
xor ( n5155 , n5154 , n5068 );
and ( n5156 , n5153 , n5155 );
xor ( n5157 , n5007 , n5011 );
xor ( n5158 , n5157 , n5016 );
and ( n5159 , n5155 , n5158 );
and ( n5160 , n5153 , n5158 );
or ( n5161 , n5156 , n5159 , n5160 );
and ( n5162 , n5151 , n5161 );
xor ( n5163 , n4919 , n4923 );
xor ( n5164 , n5163 , n4928 );
and ( n5165 , n5161 , n5164 );
and ( n5166 , n5151 , n5164 );
or ( n5167 , n5162 , n5165 , n5166 );
and ( n5168 , n1720 , n4392 );
and ( n5169 , n1705 , n4389 );
nor ( n5170 , n5168 , n5169 );
xnor ( n5171 , n5170 , n3867 );
and ( n5172 , n2295 , n2887 );
and ( n5173 , n2258 , n2885 );
nor ( n5174 , n5172 , n5173 );
xnor ( n5175 , n5174 , n2801 );
and ( n5176 , n5171 , n5175 );
and ( n5177 , n3911 , n1901 );
and ( n5178 , n3813 , n1899 );
nor ( n5179 , n5177 , n5178 );
xnor ( n5180 , n5179 , n1869 );
and ( n5181 , n5175 , n5180 );
and ( n5182 , n5171 , n5180 );
or ( n5183 , n5176 , n5181 , n5182 );
and ( n5184 , n1935 , n3742 );
and ( n5185 , n1849 , n3740 );
nor ( n5186 , n5184 , n5185 );
xnor ( n5187 , n5186 , n3538 );
and ( n5188 , n4099 , n1807 );
and ( n5189 , n3859 , n1805 );
nor ( n5190 , n5188 , n5189 );
xnor ( n5191 , n5190 , n1756 );
and ( n5192 , n5187 , n5191 );
and ( n5193 , n4402 , n1728 );
and ( n5194 , n4236 , n1726 );
nor ( n5195 , n5193 , n5194 );
xnor ( n5196 , n5195 , n1697 );
and ( n5197 , n5191 , n5196 );
and ( n5198 , n5187 , n5196 );
or ( n5199 , n5192 , n5197 , n5198 );
and ( n5200 , n5183 , n5199 );
xor ( n5201 , n5024 , n5028 );
xor ( n5202 , n5201 , n5033 );
and ( n5203 , n5199 , n5202 );
and ( n5204 , n5183 , n5202 );
or ( n5205 , n5200 , n5203 , n5204 );
xor ( n5206 , n5003 , n5019 );
xor ( n5207 , n5206 , n5036 );
and ( n5208 , n5205 , n5207 );
xor ( n5209 , n5071 , n5087 );
xor ( n5210 , n5209 , n5090 );
and ( n5211 , n5207 , n5210 );
and ( n5212 , n5205 , n5210 );
or ( n5213 , n5208 , n5211 , n5212 );
and ( n5214 , n5167 , n5213 );
xor ( n5215 , n4910 , n4912 );
xor ( n5216 , n5215 , n4915 );
and ( n5217 , n5213 , n5216 );
and ( n5218 , n5167 , n5216 );
or ( n5219 , n5214 , n5217 , n5218 );
xor ( n5220 , n4900 , n4902 );
xor ( n5221 , n5220 , n4905 );
and ( n5222 , n5219 , n5221 );
xor ( n5223 , n4918 , n4939 );
xor ( n5224 , n5223 , n4942 );
and ( n5225 , n5221 , n5224 );
and ( n5226 , n5219 , n5224 );
or ( n5227 , n5222 , n5225 , n5226 );
and ( n5228 , n5107 , n5227 );
xor ( n5229 , n4972 , n4974 );
xor ( n5230 , n5229 , n4977 );
and ( n5231 , n5227 , n5230 );
and ( n5232 , n5107 , n5230 );
or ( n5233 , n5228 , n5231 , n5232 );
and ( n5234 , n4991 , n5233 );
and ( n5235 , n1799 , n4392 );
and ( n5236 , n1720 , n4389 );
nor ( n5237 , n5235 , n5236 );
xnor ( n5238 , n5237 , n3867 );
and ( n5239 , n3414 , n2113 );
and ( n5240 , n3136 , n2111 );
nor ( n5241 , n5239 , n5240 );
xnor ( n5242 , n5241 , n2091 );
and ( n5243 , n5238 , n5242 );
and ( n5244 , n3813 , n2020 );
and ( n5245 , n3466 , n2018 );
nor ( n5246 , n5244 , n5245 );
xnor ( n5247 , n5246 , n1981 );
and ( n5248 , n5242 , n5247 );
and ( n5249 , n5238 , n5247 );
or ( n5250 , n5243 , n5248 , n5249 );
and ( n5251 , n2390 , n2887 );
and ( n5252 , n2295 , n2885 );
nor ( n5253 , n5251 , n5252 );
xnor ( n5254 , n5253 , n2801 );
and ( n5255 , n3859 , n1901 );
and ( n5256 , n3911 , n1899 );
nor ( n5257 , n5255 , n5256 );
xnor ( n5258 , n5257 , n1869 );
and ( n5259 , n5254 , n5258 );
and ( n5260 , n4236 , n1807 );
and ( n5261 , n4099 , n1805 );
nor ( n5262 , n5260 , n5261 );
xnor ( n5263 , n5262 , n1756 );
and ( n5264 , n5258 , n5263 );
and ( n5265 , n5254 , n5263 );
or ( n5266 , n5259 , n5264 , n5265 );
and ( n5267 , n5250 , n5266 );
and ( n5268 , n2258 , n3093 );
and ( n5269 , n2181 , n3091 );
nor ( n5270 , n5268 , n5269 );
xnor ( n5271 , n5270 , n3027 );
and ( n5272 , n2773 , n2483 );
and ( n5273 , n2697 , n2481 );
nor ( n5274 , n5272 , n5273 );
xnor ( n5275 , n5274 , n2418 );
and ( n5276 , n5271 , n5275 );
and ( n5277 , n3052 , n2320 );
and ( n5278 , n2897 , n2318 );
nor ( n5279 , n5277 , n5278 );
xnor ( n5280 , n5279 , n2217 );
and ( n5281 , n5275 , n5280 );
and ( n5282 , n5271 , n5280 );
or ( n5283 , n5276 , n5281 , n5282 );
and ( n5284 , n5266 , n5283 );
and ( n5285 , n5250 , n5283 );
or ( n5286 , n5267 , n5284 , n5285 );
xor ( n5287 , n5144 , n5147 );
and ( n5288 , n1849 , n4107 );
and ( n5289 , n1817 , n4105 );
nor ( n5290 , n5288 , n5289 );
xnor ( n5291 , n5290 , n3870 );
and ( n5292 , n2080 , n3367 );
and ( n5293 , n2042 , n3365 );
nor ( n5294 , n5292 , n5293 );
xnor ( n5295 , n5294 , n3306 );
and ( n5296 , n5291 , n5295 );
and ( n5297 , n5295 , n5145 );
and ( n5298 , n5291 , n5145 );
or ( n5299 , n5296 , n5297 , n5298 );
and ( n5300 , n5287 , n5299 );
and ( n5301 , n2506 , n2654 );
and ( n5302 , n2390 , n2652 );
nor ( n5303 , n5301 , n5302 );
xnor ( n5304 , n5303 , n2570 );
and ( n5305 , n5299 , n5304 );
and ( n5306 , n5287 , n5304 );
or ( n5307 , n5300 , n5305 , n5306 );
and ( n5308 , n5286 , n5307 );
xor ( n5309 , n5075 , n5079 );
xor ( n5310 , n5309 , n5084 );
and ( n5311 , n5307 , n5310 );
and ( n5312 , n5286 , n5310 );
or ( n5313 , n5308 , n5311 , n5312 );
xor ( n5314 , n5171 , n5175 );
xor ( n5315 , n5314 , n5180 );
xor ( n5316 , n5187 , n5191 );
xor ( n5317 , n5316 , n5196 );
and ( n5318 , n5315 , n5317 );
xor ( n5319 , n5111 , n5115 );
xor ( n5320 , n5319 , n5120 );
and ( n5321 , n5317 , n5320 );
and ( n5322 , n5315 , n5320 );
or ( n5323 , n5318 , n5321 , n5322 );
xor ( n5324 , n5123 , n5139 );
xor ( n5325 , n5324 , n5148 );
and ( n5326 , n5323 , n5325 );
xor ( n5327 , n5183 , n5199 );
xor ( n5328 , n5327 , n5202 );
and ( n5329 , n5325 , n5328 );
and ( n5330 , n5323 , n5328 );
or ( n5331 , n5326 , n5329 , n5330 );
and ( n5332 , n5313 , n5331 );
xor ( n5333 , n5041 , n5043 );
xor ( n5334 , n5333 , n5046 );
and ( n5335 , n5331 , n5334 );
and ( n5336 , n5313 , n5334 );
or ( n5337 , n5332 , n5335 , n5336 );
xor ( n5338 , n5039 , n5049 );
xor ( n5339 , n5338 , n5052 );
and ( n5340 , n5337 , n5339 );
xor ( n5341 , n5093 , n5095 );
xor ( n5342 , n5341 , n5098 );
and ( n5343 , n5339 , n5342 );
and ( n5344 , n5337 , n5342 );
or ( n5345 , n5340 , n5343 , n5344 );
xor ( n5346 , n5055 , n5101 );
xor ( n5347 , n5346 , n5104 );
and ( n5348 , n5345 , n5347 );
xor ( n5349 , n5219 , n5221 );
xor ( n5350 , n5349 , n5224 );
and ( n5351 , n5347 , n5350 );
and ( n5352 , n5345 , n5350 );
or ( n5353 , n5348 , n5351 , n5352 );
xor ( n5354 , n5107 , n5227 );
xor ( n5355 , n5354 , n5230 );
and ( n5356 , n5353 , n5355 );
xor ( n5357 , n5345 , n5347 );
xor ( n5358 , n5357 , n5350 );
xor ( n5359 , n5151 , n5161 );
xor ( n5360 , n5359 , n5164 );
xor ( n5361 , n5205 , n5207 );
xor ( n5362 , n5361 , n5210 );
and ( n5363 , n5360 , n5362 );
xor ( n5364 , n5313 , n5331 );
xor ( n5365 , n5364 , n5334 );
and ( n5366 , n5362 , n5365 );
and ( n5367 , n5360 , n5365 );
or ( n5368 , n5363 , n5366 , n5367 );
xor ( n5369 , n5167 , n5213 );
xor ( n5370 , n5369 , n5216 );
and ( n5371 , n5368 , n5370 );
xor ( n5372 , n5337 , n5339 );
xor ( n5373 , n5372 , n5342 );
and ( n5374 , n5370 , n5373 );
and ( n5375 , n5368 , n5373 );
or ( n5376 , n5371 , n5374 , n5375 );
and ( n5377 , n5358 , n5376 );
xor ( n5378 , n5368 , n5370 );
xor ( n5379 , n5378 , n5373 );
and ( n5380 , n1935 , n4107 );
and ( n5381 , n1849 , n4105 );
nor ( n5382 , n5380 , n5381 );
xnor ( n5383 , n5382 , n3870 );
and ( n5384 , n4402 , n1805 );
not ( n5385 , n5384 );
and ( n5386 , n5385 , n1756 );
and ( n5387 , n5383 , n5386 );
and ( n5388 , n2027 , n3742 );
and ( n5389 , n1935 , n3740 );
nor ( n5390 , n5388 , n5389 );
xnor ( n5391 , n5390 , n3538 );
and ( n5392 , n5387 , n5391 );
and ( n5393 , n2615 , n2654 );
and ( n5394 , n2506 , n2652 );
nor ( n5395 , n5393 , n5394 );
xnor ( n5396 , n5395 , n2570 );
and ( n5397 , n5391 , n5396 );
and ( n5398 , n5387 , n5396 );
or ( n5399 , n5392 , n5397 , n5398 );
xor ( n5400 , n5127 , n5131 );
xor ( n5401 , n5400 , n5136 );
and ( n5402 , n5399 , n5401 );
xor ( n5403 , n5287 , n5299 );
xor ( n5404 , n5403 , n5304 );
and ( n5405 , n5401 , n5404 );
and ( n5406 , n5399 , n5404 );
or ( n5407 , n5402 , n5405 , n5406 );
and ( n5408 , n2181 , n3367 );
and ( n5409 , n2080 , n3365 );
nor ( n5410 , n5408 , n5409 );
xnor ( n5411 , n5410 , n3306 );
and ( n5412 , n2897 , n2483 );
and ( n5413 , n2773 , n2481 );
nor ( n5414 , n5412 , n5413 );
xnor ( n5415 , n5414 , n2418 );
and ( n5416 , n5411 , n5415 );
and ( n5417 , n3136 , n2320 );
and ( n5418 , n3052 , n2318 );
nor ( n5419 , n5417 , n5418 );
xnor ( n5420 , n5419 , n2217 );
and ( n5421 , n5415 , n5420 );
and ( n5422 , n5411 , n5420 );
or ( n5423 , n5416 , n5421 , n5422 );
and ( n5424 , n1817 , n4392 );
and ( n5425 , n1799 , n4389 );
nor ( n5426 , n5424 , n5425 );
xnor ( n5427 , n5426 , n3867 );
and ( n5428 , n2506 , n2887 );
and ( n5429 , n2390 , n2885 );
nor ( n5430 , n5428 , n5429 );
xnor ( n5431 , n5430 , n2801 );
and ( n5432 , n5427 , n5431 );
and ( n5433 , n4099 , n1901 );
and ( n5434 , n3859 , n1899 );
nor ( n5435 , n5433 , n5434 );
xnor ( n5436 , n5435 , n1869 );
and ( n5437 , n5431 , n5436 );
and ( n5438 , n5427 , n5436 );
or ( n5439 , n5432 , n5437 , n5438 );
and ( n5440 , n5423 , n5439 );
and ( n5441 , n2295 , n3093 );
and ( n5442 , n2258 , n3091 );
nor ( n5443 , n5441 , n5442 );
xnor ( n5444 , n5443 , n3027 );
and ( n5445 , n3466 , n2113 );
and ( n5446 , n3414 , n2111 );
nor ( n5447 , n5445 , n5446 );
xnor ( n5448 , n5447 , n2091 );
and ( n5449 , n5444 , n5448 );
and ( n5450 , n3911 , n2020 );
and ( n5451 , n3813 , n2018 );
nor ( n5452 , n5450 , n5451 );
xnor ( n5453 , n5452 , n1981 );
and ( n5454 , n5448 , n5453 );
and ( n5455 , n5444 , n5453 );
or ( n5456 , n5449 , n5454 , n5455 );
and ( n5457 , n5439 , n5456 );
and ( n5458 , n5423 , n5456 );
or ( n5459 , n5440 , n5457 , n5458 );
and ( n5460 , n2042 , n3742 );
and ( n5461 , n2027 , n3740 );
nor ( n5462 , n5460 , n5461 );
xnor ( n5463 , n5462 , n3538 );
and ( n5464 , n2697 , n2654 );
and ( n5465 , n2615 , n2652 );
nor ( n5466 , n5464 , n5465 );
xnor ( n5467 , n5466 , n2570 );
and ( n5468 , n5463 , n5467 );
and ( n5469 , n4402 , n1807 );
and ( n5470 , n4236 , n1805 );
nor ( n5471 , n5469 , n5470 );
xnor ( n5472 , n5471 , n1756 );
and ( n5473 , n5467 , n5472 );
and ( n5474 , n5463 , n5472 );
or ( n5475 , n5468 , n5473 , n5474 );
xor ( n5476 , n5291 , n5295 );
xor ( n5477 , n5476 , n5145 );
and ( n5478 , n5475 , n5477 );
xor ( n5479 , n5238 , n5242 );
xor ( n5480 , n5479 , n5247 );
and ( n5481 , n5477 , n5480 );
and ( n5482 , n5475 , n5480 );
or ( n5483 , n5478 , n5481 , n5482 );
and ( n5484 , n5459 , n5483 );
xor ( n5485 , n5250 , n5266 );
xor ( n5486 , n5485 , n5283 );
and ( n5487 , n5483 , n5486 );
and ( n5488 , n5459 , n5486 );
or ( n5489 , n5484 , n5487 , n5488 );
and ( n5490 , n5407 , n5489 );
xor ( n5491 , n5153 , n5155 );
xor ( n5492 , n5491 , n5158 );
and ( n5493 , n5489 , n5492 );
and ( n5494 , n5407 , n5492 );
or ( n5495 , n5490 , n5493 , n5494 );
xor ( n5496 , n5254 , n5258 );
xor ( n5497 , n5496 , n5263 );
xor ( n5498 , n5271 , n5275 );
xor ( n5499 , n5498 , n5280 );
and ( n5500 , n5497 , n5499 );
xor ( n5501 , n5387 , n5391 );
xor ( n5502 , n5501 , n5396 );
and ( n5503 , n5499 , n5502 );
and ( n5504 , n5497 , n5502 );
or ( n5505 , n5500 , n5503 , n5504 );
xor ( n5506 , n5315 , n5317 );
xor ( n5507 , n5506 , n5320 );
and ( n5508 , n5505 , n5507 );
xor ( n5509 , n5399 , n5401 );
xor ( n5510 , n5509 , n5404 );
and ( n5511 , n5507 , n5510 );
and ( n5512 , n5505 , n5510 );
or ( n5513 , n5508 , n5511 , n5512 );
xor ( n5514 , n5286 , n5307 );
xor ( n5515 , n5514 , n5310 );
and ( n5516 , n5513 , n5515 );
xor ( n5517 , n5323 , n5325 );
xor ( n5518 , n5517 , n5328 );
and ( n5519 , n5515 , n5518 );
and ( n5520 , n5513 , n5518 );
or ( n5521 , n5516 , n5519 , n5520 );
and ( n5522 , n5495 , n5521 );
xor ( n5523 , n5360 , n5362 );
xor ( n5524 , n5523 , n5365 );
and ( n5525 , n5521 , n5524 );
and ( n5526 , n5495 , n5524 );
or ( n5527 , n5522 , n5525 , n5526 );
and ( n5528 , n5379 , n5527 );
xor ( n5529 , n5495 , n5521 );
xor ( n5530 , n5529 , n5524 );
xor ( n5531 , n5383 , n5386 );
and ( n5532 , n1849 , n4392 );
and ( n5533 , n1817 , n4389 );
nor ( n5534 , n5532 , n5533 );
xnor ( n5535 , n5534 , n3867 );
and ( n5536 , n3813 , n2113 );
and ( n5537 , n3466 , n2111 );
nor ( n5538 , n5536 , n5537 );
xnor ( n5539 , n5538 , n2091 );
and ( n5540 , n5535 , n5539 );
and ( n5541 , n3859 , n2020 );
and ( n5542 , n3911 , n2018 );
nor ( n5543 , n5541 , n5542 );
xnor ( n5544 , n5543 , n1981 );
and ( n5545 , n5539 , n5544 );
and ( n5546 , n5535 , n5544 );
or ( n5547 , n5540 , n5545 , n5546 );
and ( n5548 , n5531 , n5547 );
and ( n5549 , n2390 , n3093 );
and ( n5550 , n2295 , n3091 );
nor ( n5551 , n5549 , n5550 );
xnor ( n5552 , n5551 , n3027 );
and ( n5553 , n3052 , n2483 );
and ( n5554 , n2897 , n2481 );
nor ( n5555 , n5553 , n5554 );
xnor ( n5556 , n5555 , n2418 );
and ( n5557 , n5552 , n5556 );
and ( n5558 , n3414 , n2320 );
and ( n5559 , n3136 , n2318 );
nor ( n5560 , n5558 , n5559 );
xnor ( n5561 , n5560 , n2217 );
and ( n5562 , n5556 , n5561 );
and ( n5563 , n5552 , n5561 );
or ( n5564 , n5557 , n5562 , n5563 );
and ( n5565 , n5547 , n5564 );
and ( n5566 , n5531 , n5564 );
or ( n5567 , n5548 , n5565 , n5566 );
and ( n5568 , n2027 , n4107 );
and ( n5569 , n1935 , n4105 );
nor ( n5570 , n5568 , n5569 );
xnor ( n5571 , n5570 , n3870 );
and ( n5572 , n2258 , n3367 );
and ( n5573 , n2181 , n3365 );
nor ( n5574 , n5572 , n5573 );
xnor ( n5575 , n5574 , n3306 );
and ( n5576 , n5571 , n5575 );
and ( n5577 , n5575 , n5384 );
and ( n5578 , n5571 , n5384 );
or ( n5579 , n5576 , n5577 , n5578 );
and ( n5580 , n2080 , n3742 );
and ( n5581 , n2042 , n3740 );
nor ( n5582 , n5580 , n5581 );
xnor ( n5583 , n5582 , n3538 );
and ( n5584 , n2615 , n2887 );
and ( n5585 , n2506 , n2885 );
nor ( n5586 , n5584 , n5585 );
xnor ( n5587 , n5586 , n2801 );
and ( n5588 , n5583 , n5587 );
and ( n5589 , n4236 , n1901 );
and ( n5590 , n4099 , n1899 );
nor ( n5591 , n5589 , n5590 );
xnor ( n5592 , n5591 , n1869 );
and ( n5593 , n5587 , n5592 );
and ( n5594 , n5583 , n5592 );
or ( n5595 , n5588 , n5593 , n5594 );
and ( n5596 , n5579 , n5595 );
xor ( n5597 , n5463 , n5467 );
xor ( n5598 , n5597 , n5472 );
and ( n5599 , n5595 , n5598 );
and ( n5600 , n5579 , n5598 );
or ( n5601 , n5596 , n5599 , n5600 );
and ( n5602 , n5567 , n5601 );
xor ( n5603 , n5411 , n5415 );
xor ( n5604 , n5603 , n5420 );
xor ( n5605 , n5427 , n5431 );
xor ( n5606 , n5605 , n5436 );
and ( n5607 , n5604 , n5606 );
xor ( n5608 , n5444 , n5448 );
xor ( n5609 , n5608 , n5453 );
and ( n5610 , n5606 , n5609 );
and ( n5611 , n5604 , n5609 );
or ( n5612 , n5607 , n5610 , n5611 );
and ( n5613 , n5601 , n5612 );
and ( n5614 , n5567 , n5612 );
or ( n5615 , n5602 , n5613 , n5614 );
xor ( n5616 , n5423 , n5439 );
xor ( n5617 , n5616 , n5456 );
xor ( n5618 , n5475 , n5477 );
xor ( n5619 , n5618 , n5480 );
and ( n5620 , n5617 , n5619 );
xor ( n5621 , n5497 , n5499 );
xor ( n5622 , n5621 , n5502 );
and ( n5623 , n5619 , n5622 );
and ( n5624 , n5617 , n5622 );
or ( n5625 , n5620 , n5623 , n5624 );
and ( n5626 , n5615 , n5625 );
xor ( n5627 , n5459 , n5483 );
xor ( n5628 , n5627 , n5486 );
and ( n5629 , n5625 , n5628 );
and ( n5630 , n5615 , n5628 );
or ( n5631 , n5626 , n5629 , n5630 );
xor ( n5632 , n5407 , n5489 );
xor ( n5633 , n5632 , n5492 );
and ( n5634 , n5631 , n5633 );
xor ( n5635 , n5513 , n5515 );
xor ( n5636 , n5635 , n5518 );
and ( n5637 , n5633 , n5636 );
and ( n5638 , n5631 , n5636 );
or ( n5639 , n5634 , n5637 , n5638 );
and ( n5640 , n5530 , n5639 );
xor ( n5641 , n5631 , n5633 );
xor ( n5642 , n5641 , n5636 );
and ( n5643 , n2506 , n3093 );
and ( n5644 , n2390 , n3091 );
nor ( n5645 , n5643 , n5644 );
xnor ( n5646 , n5645 , n3027 );
and ( n5647 , n3911 , n2113 );
and ( n5648 , n3813 , n2111 );
nor ( n5649 , n5647 , n5648 );
xnor ( n5650 , n5649 , n2091 );
and ( n5651 , n5646 , n5650 );
and ( n5652 , n4099 , n2020 );
and ( n5653 , n3859 , n2018 );
nor ( n5654 , n5652 , n5653 );
xnor ( n5655 , n5654 , n1981 );
and ( n5656 , n5650 , n5655 );
and ( n5657 , n5646 , n5655 );
or ( n5658 , n5651 , n5656 , n5657 );
and ( n5659 , n2042 , n4107 );
and ( n5660 , n2027 , n4105 );
nor ( n5661 , n5659 , n5660 );
xnor ( n5662 , n5661 , n3870 );
and ( n5663 , n4402 , n1899 );
not ( n5664 , n5663 );
and ( n5665 , n5664 , n1869 );
and ( n5666 , n5662 , n5665 );
and ( n5667 , n5658 , n5666 );
and ( n5668 , n2773 , n2654 );
and ( n5669 , n2697 , n2652 );
nor ( n5670 , n5668 , n5669 );
xnor ( n5671 , n5670 , n2570 );
and ( n5672 , n5666 , n5671 );
and ( n5673 , n5658 , n5671 );
or ( n5674 , n5667 , n5672 , n5673 );
xor ( n5675 , n5571 , n5575 );
xor ( n5676 , n5675 , n5384 );
xor ( n5677 , n5535 , n5539 );
xor ( n5678 , n5677 , n5544 );
and ( n5679 , n5676 , n5678 );
xor ( n5680 , n5552 , n5556 );
xor ( n5681 , n5680 , n5561 );
and ( n5682 , n5678 , n5681 );
and ( n5683 , n5676 , n5681 );
or ( n5684 , n5679 , n5682 , n5683 );
and ( n5685 , n5674 , n5684 );
xor ( n5686 , n5579 , n5595 );
xor ( n5687 , n5686 , n5598 );
and ( n5688 , n5684 , n5687 );
and ( n5689 , n5674 , n5687 );
or ( n5690 , n5685 , n5688 , n5689 );
and ( n5691 , n2295 , n3367 );
and ( n5692 , n2258 , n3365 );
nor ( n5693 , n5691 , n5692 );
xnor ( n5694 , n5693 , n3306 );
and ( n5695 , n3136 , n2483 );
and ( n5696 , n3052 , n2481 );
nor ( n5697 , n5695 , n5696 );
xnor ( n5698 , n5697 , n2418 );
and ( n5699 , n5694 , n5698 );
and ( n5700 , n3466 , n2320 );
and ( n5701 , n3414 , n2318 );
nor ( n5702 , n5700 , n5701 );
xnor ( n5703 , n5702 , n2217 );
and ( n5704 , n5698 , n5703 );
and ( n5705 , n5694 , n5703 );
or ( n5706 , n5699 , n5704 , n5705 );
and ( n5707 , n1935 , n4392 );
and ( n5708 , n1849 , n4389 );
nor ( n5709 , n5707 , n5708 );
xnor ( n5710 , n5709 , n3867 );
and ( n5711 , n2181 , n3742 );
and ( n5712 , n2080 , n3740 );
nor ( n5713 , n5711 , n5712 );
xnor ( n5714 , n5713 , n3538 );
and ( n5715 , n5710 , n5714 );
and ( n5716 , n4402 , n1901 );
and ( n5717 , n4236 , n1899 );
nor ( n5718 , n5716 , n5717 );
xnor ( n5719 , n5718 , n1869 );
and ( n5720 , n5714 , n5719 );
and ( n5721 , n5710 , n5719 );
or ( n5722 , n5715 , n5720 , n5721 );
and ( n5723 , n5706 , n5722 );
xor ( n5724 , n5583 , n5587 );
xor ( n5725 , n5724 , n5592 );
and ( n5726 , n5722 , n5725 );
and ( n5727 , n5706 , n5725 );
or ( n5728 , n5723 , n5726 , n5727 );
xor ( n5729 , n5531 , n5547 );
xor ( n5730 , n5729 , n5564 );
and ( n5731 , n5728 , n5730 );
xor ( n5732 , n5604 , n5606 );
xor ( n5733 , n5732 , n5609 );
and ( n5734 , n5730 , n5733 );
and ( n5735 , n5728 , n5733 );
or ( n5736 , n5731 , n5734 , n5735 );
and ( n5737 , n5690 , n5736 );
xor ( n5738 , n5567 , n5601 );
xor ( n5739 , n5738 , n5612 );
and ( n5740 , n5736 , n5739 );
and ( n5741 , n5690 , n5739 );
or ( n5742 , n5737 , n5740 , n5741 );
xor ( n5743 , n5505 , n5507 );
xor ( n5744 , n5743 , n5510 );
and ( n5745 , n5742 , n5744 );
xor ( n5746 , n5615 , n5625 );
xor ( n5747 , n5746 , n5628 );
and ( n5748 , n5744 , n5747 );
and ( n5749 , n5742 , n5747 );
or ( n5750 , n5745 , n5748 , n5749 );
and ( n5751 , n5642 , n5750 );
and ( n5752 , n2027 , n4392 );
and ( n5753 , n1935 , n4389 );
nor ( n5754 , n5752 , n5753 );
xnor ( n5755 , n5754 , n3867 );
and ( n5756 , n3859 , n2113 );
and ( n5757 , n3911 , n2111 );
nor ( n5758 , n5756 , n5757 );
xnor ( n5759 , n5758 , n2091 );
and ( n5760 , n5755 , n5759 );
and ( n5761 , n4236 , n2020 );
and ( n5762 , n4099 , n2018 );
nor ( n5763 , n5761 , n5762 );
xnor ( n5764 , n5763 , n1981 );
and ( n5765 , n5759 , n5764 );
and ( n5766 , n5755 , n5764 );
or ( n5767 , n5760 , n5765 , n5766 );
and ( n5768 , n2080 , n4107 );
and ( n5769 , n2042 , n4105 );
nor ( n5770 , n5768 , n5769 );
xnor ( n5771 , n5770 , n3870 );
and ( n5772 , n2390 , n3367 );
and ( n5773 , n2295 , n3365 );
nor ( n5774 , n5772 , n5773 );
xnor ( n5775 , n5774 , n3306 );
and ( n5776 , n5771 , n5775 );
and ( n5777 , n5775 , n5663 );
and ( n5778 , n5771 , n5663 );
or ( n5779 , n5776 , n5777 , n5778 );
and ( n5780 , n5767 , n5779 );
and ( n5781 , n2258 , n3742 );
and ( n5782 , n2181 , n3740 );
nor ( n5783 , n5781 , n5782 );
xnor ( n5784 , n5783 , n3538 );
and ( n5785 , n2773 , n2887 );
and ( n5786 , n2697 , n2885 );
nor ( n5787 , n5785 , n5786 );
xnor ( n5788 , n5787 , n2801 );
and ( n5789 , n5784 , n5788 );
and ( n5790 , n3052 , n2654 );
and ( n5791 , n2897 , n2652 );
nor ( n5792 , n5790 , n5791 );
xnor ( n5793 , n5792 , n2570 );
and ( n5794 , n5788 , n5793 );
and ( n5795 , n5784 , n5793 );
or ( n5796 , n5789 , n5794 , n5795 );
and ( n5797 , n5779 , n5796 );
and ( n5798 , n5767 , n5796 );
or ( n5799 , n5780 , n5797 , n5798 );
xor ( n5800 , n5662 , n5665 );
and ( n5801 , n2697 , n2887 );
and ( n5802 , n2615 , n2885 );
nor ( n5803 , n5801 , n5802 );
xnor ( n5804 , n5803 , n2801 );
and ( n5805 , n5800 , n5804 );
and ( n5806 , n2897 , n2654 );
and ( n5807 , n2773 , n2652 );
nor ( n5808 , n5806 , n5807 );
xnor ( n5809 , n5808 , n2570 );
and ( n5810 , n5804 , n5809 );
and ( n5811 , n5800 , n5809 );
or ( n5812 , n5805 , n5810 , n5811 );
and ( n5813 , n5799 , n5812 );
xor ( n5814 , n5658 , n5666 );
xor ( n5815 , n5814 , n5671 );
and ( n5816 , n5812 , n5815 );
and ( n5817 , n5799 , n5815 );
or ( n5818 , n5813 , n5816 , n5817 );
and ( n5819 , n2615 , n3093 );
and ( n5820 , n2506 , n3091 );
nor ( n5821 , n5819 , n5820 );
xnor ( n5822 , n5821 , n3027 );
and ( n5823 , n3414 , n2483 );
and ( n5824 , n3136 , n2481 );
nor ( n5825 , n5823 , n5824 );
xnor ( n5826 , n5825 , n2418 );
and ( n5827 , n5822 , n5826 );
and ( n5828 , n3813 , n2320 );
and ( n5829 , n3466 , n2318 );
nor ( n5830 , n5828 , n5829 );
xnor ( n5831 , n5830 , n2217 );
and ( n5832 , n5826 , n5831 );
and ( n5833 , n5822 , n5831 );
or ( n5834 , n5827 , n5832 , n5833 );
xor ( n5835 , n5646 , n5650 );
xor ( n5836 , n5835 , n5655 );
and ( n5837 , n5834 , n5836 );
xor ( n5838 , n5710 , n5714 );
xor ( n5839 , n5838 , n5719 );
and ( n5840 , n5836 , n5839 );
and ( n5841 , n5834 , n5839 );
or ( n5842 , n5837 , n5840 , n5841 );
xor ( n5843 , n5706 , n5722 );
xor ( n5844 , n5843 , n5725 );
and ( n5845 , n5842 , n5844 );
xor ( n5846 , n5676 , n5678 );
xor ( n5847 , n5846 , n5681 );
and ( n5848 , n5844 , n5847 );
and ( n5849 , n5842 , n5847 );
or ( n5850 , n5845 , n5848 , n5849 );
and ( n5851 , n5818 , n5850 );
xor ( n5852 , n5674 , n5684 );
xor ( n5853 , n5852 , n5687 );
and ( n5854 , n5850 , n5853 );
and ( n5855 , n5818 , n5853 );
or ( n5856 , n5851 , n5854 , n5855 );
xor ( n5857 , n5690 , n5736 );
xor ( n5858 , n5857 , n5739 );
and ( n5859 , n5856 , n5858 );
xor ( n5860 , n5617 , n5619 );
xor ( n5861 , n5860 , n5622 );
and ( n5862 , n5858 , n5861 );
and ( n5863 , n5856 , n5861 );
or ( n5864 , n5859 , n5862 , n5863 );
xor ( n5865 , n5742 , n5744 );
xor ( n5866 , n5865 , n5747 );
and ( n5867 , n5864 , n5866 );
xor ( n5868 , n5856 , n5858 );
xor ( n5869 , n5868 , n5861 );
and ( n5870 , n2697 , n3093 );
and ( n5871 , n2615 , n3091 );
nor ( n5872 , n5870 , n5871 );
xnor ( n5873 , n5872 , n3027 );
and ( n5874 , n4099 , n2113 );
and ( n5875 , n3859 , n2111 );
nor ( n5876 , n5874 , n5875 );
xnor ( n5877 , n5876 , n2091 );
and ( n5878 , n5873 , n5877 );
and ( n5879 , n4402 , n2020 );
and ( n5880 , n4236 , n2018 );
nor ( n5881 , n5879 , n5880 );
xnor ( n5882 , n5881 , n1981 );
and ( n5883 , n5877 , n5882 );
and ( n5884 , n5873 , n5882 );
or ( n5885 , n5878 , n5883 , n5884 );
and ( n5886 , n2042 , n4392 );
and ( n5887 , n2027 , n4389 );
nor ( n5888 , n5886 , n5887 );
xnor ( n5889 , n5888 , n3867 );
and ( n5890 , n2295 , n3742 );
and ( n5891 , n2258 , n3740 );
nor ( n5892 , n5890 , n5891 );
xnor ( n5893 , n5892 , n3538 );
and ( n5894 , n5889 , n5893 );
and ( n5895 , n2897 , n2887 );
and ( n5896 , n2773 , n2885 );
nor ( n5897 , n5895 , n5896 );
xnor ( n5898 , n5897 , n2801 );
and ( n5899 , n5893 , n5898 );
and ( n5900 , n5889 , n5898 );
or ( n5901 , n5894 , n5899 , n5900 );
and ( n5902 , n5885 , n5901 );
and ( n5903 , n2181 , n4107 );
and ( n5904 , n2080 , n4105 );
nor ( n5905 , n5903 , n5904 );
xnor ( n5906 , n5905 , n3870 );
and ( n5907 , n4402 , n2018 );
not ( n5908 , n5907 );
and ( n5909 , n5908 , n1981 );
and ( n5910 , n5906 , n5909 );
and ( n5911 , n5901 , n5910 );
and ( n5912 , n5885 , n5910 );
or ( n5913 , n5902 , n5911 , n5912 );
xor ( n5914 , n5694 , n5698 );
xor ( n5915 , n5914 , n5703 );
and ( n5916 , n5913 , n5915 );
xor ( n5917 , n5800 , n5804 );
xor ( n5918 , n5917 , n5809 );
and ( n5919 , n5915 , n5918 );
and ( n5920 , n5913 , n5918 );
or ( n5921 , n5916 , n5919 , n5920 );
and ( n5922 , n2506 , n3367 );
and ( n5923 , n2390 , n3365 );
nor ( n5924 , n5922 , n5923 );
xnor ( n5925 , n5924 , n3306 );
and ( n5926 , n3466 , n2483 );
and ( n5927 , n3414 , n2481 );
nor ( n5928 , n5926 , n5927 );
xnor ( n5929 , n5928 , n2418 );
and ( n5930 , n5925 , n5929 );
and ( n5931 , n3911 , n2320 );
and ( n5932 , n3813 , n2318 );
nor ( n5933 , n5931 , n5932 );
xnor ( n5934 , n5933 , n2217 );
and ( n5935 , n5929 , n5934 );
and ( n5936 , n5925 , n5934 );
or ( n5937 , n5930 , n5935 , n5936 );
xor ( n5938 , n5784 , n5788 );
xor ( n5939 , n5938 , n5793 );
and ( n5940 , n5937 , n5939 );
xor ( n5941 , n5822 , n5826 );
xor ( n5942 , n5941 , n5831 );
and ( n5943 , n5939 , n5942 );
and ( n5944 , n5937 , n5942 );
or ( n5945 , n5940 , n5943 , n5944 );
xor ( n5946 , n5767 , n5779 );
xor ( n5947 , n5946 , n5796 );
and ( n5948 , n5945 , n5947 );
xor ( n5949 , n5834 , n5836 );
xor ( n5950 , n5949 , n5839 );
and ( n5951 , n5947 , n5950 );
and ( n5952 , n5945 , n5950 );
or ( n5953 , n5948 , n5951 , n5952 );
and ( n5954 , n5921 , n5953 );
xor ( n5955 , n5799 , n5812 );
xor ( n5956 , n5955 , n5815 );
and ( n5957 , n5953 , n5956 );
and ( n5958 , n5921 , n5956 );
or ( n5959 , n5954 , n5957 , n5958 );
xor ( n5960 , n5728 , n5730 );
xor ( n5961 , n5960 , n5733 );
and ( n5962 , n5959 , n5961 );
xor ( n5963 , n5818 , n5850 );
xor ( n5964 , n5963 , n5853 );
and ( n5965 , n5961 , n5964 );
and ( n5966 , n5959 , n5964 );
or ( n5967 , n5962 , n5965 , n5966 );
and ( n5968 , n5869 , n5967 );
xor ( n5969 , n5959 , n5961 );
xor ( n5970 , n5969 , n5964 );
xor ( n5971 , n5906 , n5909 );
and ( n5972 , n2258 , n4107 );
and ( n5973 , n2181 , n4105 );
nor ( n5974 , n5972 , n5973 );
xnor ( n5975 , n5974 , n3870 );
and ( n5976 , n3813 , n2483 );
and ( n5977 , n3466 , n2481 );
nor ( n5978 , n5976 , n5977 );
xnor ( n5979 , n5978 , n2418 );
and ( n5980 , n5975 , n5979 );
and ( n5981 , n3859 , n2320 );
and ( n5982 , n3911 , n2318 );
nor ( n5983 , n5981 , n5982 );
xnor ( n5984 , n5983 , n2217 );
and ( n5985 , n5979 , n5984 );
and ( n5986 , n5975 , n5984 );
or ( n5987 , n5980 , n5985 , n5986 );
and ( n5988 , n5971 , n5987 );
and ( n5989 , n3136 , n2654 );
and ( n5990 , n3052 , n2652 );
nor ( n5991 , n5989 , n5990 );
xnor ( n5992 , n5991 , n2570 );
and ( n5993 , n5987 , n5992 );
and ( n5994 , n5971 , n5992 );
or ( n5995 , n5988 , n5993 , n5994 );
xor ( n5996 , n5755 , n5759 );
xor ( n5997 , n5996 , n5764 );
and ( n5998 , n5995 , n5997 );
xor ( n5999 , n5771 , n5775 );
xor ( n6000 , n5999 , n5663 );
and ( n6001 , n5997 , n6000 );
and ( n6002 , n5995 , n6000 );
or ( n6003 , n5998 , n6001 , n6002 );
xor ( n6004 , n5913 , n5915 );
xor ( n6005 , n6004 , n5918 );
and ( n6006 , n6003 , n6005 );
xor ( n6007 , n5945 , n5947 );
xor ( n6008 , n6007 , n5950 );
and ( n6009 , n6005 , n6008 );
and ( n6010 , n6003 , n6008 );
or ( n6011 , n6006 , n6009 , n6010 );
xor ( n6012 , n5842 , n5844 );
xor ( n6013 , n6012 , n5847 );
and ( n6014 , n6011 , n6013 );
xor ( n6015 , n5921 , n5953 );
xor ( n6016 , n6015 , n5956 );
and ( n6017 , n6013 , n6016 );
and ( n6018 , n6011 , n6016 );
or ( n6019 , n6014 , n6017 , n6018 );
and ( n6020 , n5970 , n6019 );
xor ( n6021 , n6011 , n6013 );
xor ( n6022 , n6021 , n6016 );
and ( n6023 , n2080 , n4392 );
and ( n6024 , n2042 , n4389 );
nor ( n6025 , n6023 , n6024 );
xnor ( n6026 , n6025 , n3867 );
and ( n6027 , n2615 , n3367 );
and ( n6028 , n2506 , n3365 );
nor ( n6029 , n6027 , n6028 );
xnor ( n6030 , n6029 , n3306 );
and ( n6031 , n6026 , n6030 );
and ( n6032 , n6030 , n5907 );
and ( n6033 , n6026 , n5907 );
or ( n6034 , n6031 , n6032 , n6033 );
and ( n6035 , n2390 , n3742 );
and ( n6036 , n2295 , n3740 );
nor ( n6037 , n6035 , n6036 );
xnor ( n6038 , n6037 , n3538 );
and ( n6039 , n2773 , n3093 );
and ( n6040 , n2697 , n3091 );
nor ( n6041 , n6039 , n6040 );
xnor ( n6042 , n6041 , n3027 );
and ( n6043 , n6038 , n6042 );
and ( n6044 , n4236 , n2113 );
and ( n6045 , n4099 , n2111 );
nor ( n6046 , n6044 , n6045 );
xnor ( n6047 , n6046 , n2091 );
and ( n6048 , n6042 , n6047 );
and ( n6049 , n6038 , n6047 );
or ( n6050 , n6043 , n6048 , n6049 );
and ( n6051 , n6034 , n6050 );
xor ( n6052 , n5889 , n5893 );
xor ( n6053 , n6052 , n5898 );
and ( n6054 , n6050 , n6053 );
and ( n6055 , n6034 , n6053 );
or ( n6056 , n6051 , n6054 , n6055 );
and ( n6057 , n2181 , n4392 );
and ( n6058 , n2080 , n4389 );
nor ( n6059 , n6057 , n6058 );
xnor ( n6060 , n6059 , n3867 );
and ( n6061 , n4402 , n2111 );
not ( n6062 , n6061 );
and ( n6063 , n6062 , n2091 );
and ( n6064 , n6060 , n6063 );
and ( n6065 , n3052 , n2887 );
and ( n6066 , n2897 , n2885 );
nor ( n6067 , n6065 , n6066 );
xnor ( n6068 , n6067 , n2801 );
and ( n6069 , n6064 , n6068 );
and ( n6070 , n3414 , n2654 );
and ( n6071 , n3136 , n2652 );
nor ( n6072 , n6070 , n6071 );
xnor ( n6073 , n6072 , n2570 );
and ( n6074 , n6068 , n6073 );
and ( n6075 , n6064 , n6073 );
or ( n6076 , n6069 , n6074 , n6075 );
xor ( n6077 , n5925 , n5929 );
xor ( n6078 , n6077 , n5934 );
and ( n6079 , n6076 , n6078 );
xor ( n6080 , n5873 , n5877 );
xor ( n6081 , n6080 , n5882 );
and ( n6082 , n6078 , n6081 );
and ( n6083 , n6076 , n6081 );
or ( n6084 , n6079 , n6082 , n6083 );
and ( n6085 , n6056 , n6084 );
xor ( n6086 , n5885 , n5901 );
xor ( n6087 , n6086 , n5910 );
and ( n6088 , n6084 , n6087 );
and ( n6089 , n6056 , n6087 );
or ( n6090 , n6085 , n6088 , n6089 );
and ( n6091 , n2295 , n4107 );
and ( n6092 , n2258 , n4105 );
nor ( n6093 , n6091 , n6092 );
xnor ( n6094 , n6093 , n3870 );
and ( n6095 , n2897 , n3093 );
and ( n6096 , n2773 , n3091 );
nor ( n6097 , n6095 , n6096 );
xnor ( n6098 , n6097 , n3027 );
and ( n6099 , n6094 , n6098 );
and ( n6100 , n4402 , n2113 );
and ( n6101 , n4236 , n2111 );
nor ( n6102 , n6100 , n6101 );
xnor ( n6103 , n6102 , n2091 );
and ( n6104 , n6098 , n6103 );
and ( n6105 , n6094 , n6103 );
or ( n6106 , n6099 , n6104 , n6105 );
and ( n6107 , n2506 , n3742 );
and ( n6108 , n2390 , n3740 );
nor ( n6109 , n6107 , n6108 );
xnor ( n6110 , n6109 , n3538 );
and ( n6111 , n3136 , n2887 );
and ( n6112 , n3052 , n2885 );
nor ( n6113 , n6111 , n6112 );
xnor ( n6114 , n6113 , n2801 );
and ( n6115 , n6110 , n6114 );
and ( n6116 , n3466 , n2654 );
and ( n6117 , n3414 , n2652 );
nor ( n6118 , n6116 , n6117 );
xnor ( n6119 , n6118 , n2570 );
and ( n6120 , n6114 , n6119 );
and ( n6121 , n6110 , n6119 );
or ( n6122 , n6115 , n6120 , n6121 );
and ( n6123 , n6106 , n6122 );
and ( n6124 , n2697 , n3367 );
and ( n6125 , n2615 , n3365 );
nor ( n6126 , n6124 , n6125 );
xnor ( n6127 , n6126 , n3306 );
and ( n6128 , n3911 , n2483 );
and ( n6129 , n3813 , n2481 );
nor ( n6130 , n6128 , n6129 );
xnor ( n6131 , n6130 , n2418 );
and ( n6132 , n6127 , n6131 );
and ( n6133 , n4099 , n2320 );
and ( n6134 , n3859 , n2318 );
nor ( n6135 , n6133 , n6134 );
xnor ( n6136 , n6135 , n2217 );
and ( n6137 , n6131 , n6136 );
and ( n6138 , n6127 , n6136 );
or ( n6139 , n6132 , n6137 , n6138 );
and ( n6140 , n6122 , n6139 );
and ( n6141 , n6106 , n6139 );
or ( n6142 , n6123 , n6140 , n6141 );
xor ( n6143 , n5971 , n5987 );
xor ( n6144 , n6143 , n5992 );
and ( n6145 , n6142 , n6144 );
xor ( n6146 , n6034 , n6050 );
xor ( n6147 , n6146 , n6053 );
and ( n6148 , n6144 , n6147 );
and ( n6149 , n6142 , n6147 );
or ( n6150 , n6145 , n6148 , n6149 );
xor ( n6151 , n5937 , n5939 );
xor ( n6152 , n6151 , n5942 );
and ( n6153 , n6150 , n6152 );
xor ( n6154 , n5995 , n5997 );
xor ( n6155 , n6154 , n6000 );
and ( n6156 , n6152 , n6155 );
and ( n6157 , n6150 , n6155 );
or ( n6158 , n6153 , n6156 , n6157 );
and ( n6159 , n6090 , n6158 );
xor ( n6160 , n6003 , n6005 );
xor ( n6161 , n6160 , n6008 );
and ( n6162 , n6158 , n6161 );
and ( n6163 , n6090 , n6161 );
or ( n6164 , n6159 , n6162 , n6163 );
and ( n6165 , n6022 , n6164 );
xor ( n6166 , n6090 , n6158 );
xor ( n6167 , n6166 , n6161 );
xor ( n6168 , n6026 , n6030 );
xor ( n6169 , n6168 , n5907 );
xor ( n6170 , n6038 , n6042 );
xor ( n6171 , n6170 , n6047 );
and ( n6172 , n6169 , n6171 );
xor ( n6173 , n5975 , n5979 );
xor ( n6174 , n6173 , n5984 );
and ( n6175 , n6171 , n6174 );
and ( n6176 , n6169 , n6174 );
or ( n6177 , n6172 , n6175 , n6176 );
xor ( n6178 , n6076 , n6078 );
xor ( n6179 , n6178 , n6081 );
and ( n6180 , n6177 , n6179 );
xor ( n6181 , n6142 , n6144 );
xor ( n6182 , n6181 , n6147 );
and ( n6183 , n6179 , n6182 );
and ( n6184 , n6177 , n6182 );
or ( n6185 , n6180 , n6183 , n6184 );
xor ( n6186 , n6056 , n6084 );
xor ( n6187 , n6186 , n6087 );
and ( n6188 , n6185 , n6187 );
xor ( n6189 , n6150 , n6152 );
xor ( n6190 , n6189 , n6155 );
and ( n6191 , n6187 , n6190 );
and ( n6192 , n6185 , n6190 );
or ( n6193 , n6188 , n6191 , n6192 );
and ( n6194 , n6167 , n6193 );
xor ( n6195 , n6185 , n6187 );
xor ( n6196 , n6195 , n6190 );
xor ( n6197 , n6106 , n6122 );
xor ( n6198 , n6197 , n6139 );
xor ( n6199 , n6169 , n6171 );
xor ( n6200 , n6199 , n6174 );
and ( n6201 , n6198 , n6200 );
xor ( n6202 , n6064 , n6068 );
xor ( n6203 , n6202 , n6073 );
and ( n6204 , n2615 , n3742 );
and ( n6205 , n2506 , n3740 );
nor ( n6206 , n6204 , n6205 );
xnor ( n6207 , n6206 , n3538 );
and ( n6208 , n3052 , n3093 );
and ( n6209 , n2897 , n3091 );
nor ( n6210 , n6208 , n6209 );
xnor ( n6211 , n6210 , n3027 );
and ( n6212 , n6207 , n6211 );
and ( n6213 , n3414 , n2887 );
and ( n6214 , n3136 , n2885 );
nor ( n6215 , n6213 , n6214 );
xnor ( n6216 , n6215 , n2801 );
and ( n6217 , n6211 , n6216 );
and ( n6218 , n6207 , n6216 );
or ( n6219 , n6212 , n6217 , n6218 );
xor ( n6220 , n6110 , n6114 );
xor ( n6221 , n6220 , n6119 );
and ( n6222 , n6219 , n6221 );
xor ( n6223 , n6127 , n6131 );
xor ( n6224 , n6223 , n6136 );
and ( n6225 , n6221 , n6224 );
and ( n6226 , n6219 , n6224 );
or ( n6227 , n6222 , n6225 , n6226 );
and ( n6228 , n6203 , n6227 );
and ( n6229 , n2258 , n4392 );
and ( n6230 , n2181 , n4389 );
nor ( n6231 , n6229 , n6230 );
xnor ( n6232 , n6231 , n3867 );
and ( n6233 , n2773 , n3367 );
and ( n6234 , n2697 , n3365 );
nor ( n6235 , n6233 , n6234 );
xnor ( n6236 , n6235 , n3306 );
and ( n6237 , n6232 , n6236 );
and ( n6238 , n6236 , n6061 );
and ( n6239 , n6232 , n6061 );
or ( n6240 , n6237 , n6238 , n6239 );
xor ( n6241 , n6060 , n6063 );
and ( n6242 , n6240 , n6241 );
and ( n6243 , n6227 , n6242 );
and ( n6244 , n6203 , n6242 );
or ( n6245 , n6228 , n6243 , n6244 );
and ( n6246 , n6201 , n6245 );
xor ( n6247 , n6177 , n6179 );
xor ( n6248 , n6247 , n6182 );
and ( n6249 , n6245 , n6248 );
and ( n6250 , n6201 , n6248 );
or ( n6251 , n6246 , n6249 , n6250 );
and ( n6252 , n6196 , n6251 );
xor ( n6253 , n6198 , n6200 );
xor ( n6254 , n6094 , n6098 );
xor ( n6255 , n6254 , n6103 );
and ( n6256 , n2390 , n4107 );
and ( n6257 , n2295 , n4105 );
nor ( n6258 , n6256 , n6257 );
xnor ( n6259 , n6258 , n3870 );
and ( n6260 , n3859 , n2483 );
and ( n6261 , n3911 , n2481 );
nor ( n6262 , n6260 , n6261 );
xnor ( n6263 , n6262 , n2418 );
and ( n6264 , n6259 , n6263 );
and ( n6265 , n4236 , n2320 );
and ( n6266 , n4099 , n2318 );
nor ( n6267 , n6265 , n6266 );
xnor ( n6268 , n6267 , n2217 );
and ( n6269 , n6263 , n6268 );
and ( n6270 , n6259 , n6268 );
or ( n6271 , n6264 , n6269 , n6270 );
and ( n6272 , n6255 , n6271 );
xor ( n6273 , n6219 , n6221 );
xor ( n6274 , n6273 , n6224 );
and ( n6275 , n6271 , n6274 );
and ( n6276 , n6255 , n6274 );
or ( n6277 , n6272 , n6275 , n6276 );
and ( n6278 , n6253 , n6277 );
xor ( n6279 , n6240 , n6241 );
and ( n6280 , n2897 , n3367 );
and ( n6281 , n2773 , n3365 );
nor ( n6282 , n6280 , n6281 );
xnor ( n6283 , n6282 , n3306 );
and ( n6284 , n4099 , n2483 );
and ( n6285 , n3859 , n2481 );
nor ( n6286 , n6284 , n6285 );
xnor ( n6287 , n6286 , n2418 );
and ( n6288 , n6283 , n6287 );
and ( n6289 , n4402 , n2320 );
and ( n6290 , n4236 , n2318 );
nor ( n6291 , n6289 , n6290 );
xnor ( n6292 , n6291 , n2217 );
and ( n6293 , n6287 , n6292 );
and ( n6294 , n6283 , n6292 );
or ( n6295 , n6288 , n6293 , n6294 );
and ( n6296 , n2295 , n4392 );
and ( n6297 , n2258 , n4389 );
nor ( n6298 , n6296 , n6297 );
xnor ( n6299 , n6298 , n3867 );
and ( n6300 , n4402 , n2318 );
not ( n6301 , n6300 );
and ( n6302 , n6301 , n2217 );
and ( n6303 , n6299 , n6302 );
and ( n6304 , n6295 , n6303 );
and ( n6305 , n3813 , n2654 );
and ( n6306 , n3466 , n2652 );
nor ( n6307 , n6305 , n6306 );
xnor ( n6308 , n6307 , n2570 );
and ( n6309 , n6303 , n6308 );
and ( n6310 , n6295 , n6308 );
or ( n6311 , n6304 , n6309 , n6310 );
and ( n6312 , n6279 , n6311 );
and ( n6313 , n2506 , n4107 );
and ( n6314 , n2390 , n4105 );
nor ( n6315 , n6313 , n6314 );
xnor ( n6316 , n6315 , n3870 );
and ( n6317 , n2697 , n3742 );
and ( n6318 , n2615 , n3740 );
nor ( n6319 , n6317 , n6318 );
xnor ( n6320 , n6319 , n3538 );
and ( n6321 , n6316 , n6320 );
and ( n6322 , n3136 , n3093 );
and ( n6323 , n3052 , n3091 );
nor ( n6324 , n6322 , n6323 );
xnor ( n6325 , n6324 , n3027 );
and ( n6326 , n6320 , n6325 );
and ( n6327 , n6316 , n6325 );
or ( n6328 , n6321 , n6326 , n6327 );
xor ( n6329 , n6232 , n6236 );
xor ( n6330 , n6329 , n6061 );
and ( n6331 , n6328 , n6330 );
xor ( n6332 , n6207 , n6211 );
xor ( n6333 , n6332 , n6216 );
and ( n6334 , n6330 , n6333 );
and ( n6335 , n6328 , n6333 );
or ( n6336 , n6331 , n6334 , n6335 );
and ( n6337 , n6311 , n6336 );
and ( n6338 , n6279 , n6336 );
or ( n6339 , n6312 , n6337 , n6338 );
and ( n6340 , n6277 , n6339 );
and ( n6341 , n6253 , n6339 );
or ( n6342 , n6278 , n6340 , n6341 );
xor ( n6343 , n6203 , n6227 );
xor ( n6344 , n6343 , n6242 );
xor ( n6345 , n6259 , n6263 );
xor ( n6346 , n6345 , n6268 );
xor ( n6347 , n6295 , n6303 );
xor ( n6348 , n6347 , n6308 );
and ( n6349 , n6346 , n6348 );
xor ( n6350 , n6328 , n6330 );
xor ( n6351 , n6350 , n6333 );
and ( n6352 , n6348 , n6351 );
and ( n6353 , n6346 , n6351 );
or ( n6354 , n6349 , n6352 , n6353 );
xor ( n6355 , n6255 , n6271 );
xor ( n6356 , n6355 , n6274 );
and ( n6357 , n6354 , n6356 );
xor ( n6358 , n6279 , n6311 );
xor ( n6359 , n6358 , n6336 );
and ( n6360 , n6356 , n6359 );
and ( n6361 , n6354 , n6359 );
or ( n6362 , n6357 , n6360 , n6361 );
and ( n6363 , n6344 , n6362 );
xor ( n6364 , n6253 , n6277 );
xor ( n6365 , n6364 , n6339 );
and ( n6366 , n6362 , n6365 );
and ( n6367 , n6344 , n6365 );
or ( n6368 , n6363 , n6366 , n6367 );
and ( n6369 , n6342 , n6368 );
xor ( n6370 , n6201 , n6245 );
xor ( n6371 , n6370 , n6248 );
and ( n6372 , n6368 , n6371 );
and ( n6373 , n6342 , n6371 );
or ( n6374 , n6369 , n6372 , n6373 );
and ( n6375 , n6251 , n6374 );
and ( n6376 , n6196 , n6374 );
or ( n6377 , n6252 , n6375 , n6376 );
and ( n6378 , n6193 , n6377 );
and ( n6379 , n6167 , n6377 );
or ( n6380 , n6194 , n6378 , n6379 );
and ( n6381 , n6164 , n6380 );
and ( n6382 , n6022 , n6380 );
or ( n6383 , n6165 , n6381 , n6382 );
and ( n6384 , n6019 , n6383 );
and ( n6385 , n5970 , n6383 );
or ( n6386 , n6020 , n6384 , n6385 );
and ( n6387 , n5967 , n6386 );
and ( n6388 , n5869 , n6386 );
or ( n6389 , n5968 , n6387 , n6388 );
and ( n6390 , n5866 , n6389 );
and ( n6391 , n5864 , n6389 );
or ( n6392 , n5867 , n6390 , n6391 );
and ( n6393 , n5750 , n6392 );
and ( n6394 , n5642 , n6392 );
or ( n6395 , n5751 , n6393 , n6394 );
and ( n6396 , n5639 , n6395 );
and ( n6397 , n5530 , n6395 );
or ( n6398 , n5640 , n6396 , n6397 );
and ( n6399 , n5527 , n6398 );
and ( n6400 , n5379 , n6398 );
or ( n6401 , n5528 , n6399 , n6400 );
and ( n6402 , n5376 , n6401 );
and ( n6403 , n5358 , n6401 );
or ( n6404 , n5377 , n6402 , n6403 );
and ( n6405 , n5355 , n6404 );
and ( n6406 , n5353 , n6404 );
or ( n6407 , n5356 , n6405 , n6406 );
and ( n6408 , n5233 , n6407 );
and ( n6409 , n4991 , n6407 );
or ( n6410 , n5234 , n6408 , n6409 );
and ( n6411 , n4988 , n6410 );
and ( n6412 , n4970 , n6410 );
or ( n6413 , n4989 , n6411 , n6412 );
and ( n6414 , n4967 , n6413 );
and ( n6415 , n4965 , n6413 );
or ( n6416 , n4968 , n6414 , n6415 );
and ( n6417 , n4799 , n6416 );
and ( n6418 , n4660 , n6416 );
or ( n6419 , n4800 , n6417 , n6418 );
and ( n6420 , n4657 , n6419 );
and ( n6421 , n4495 , n6419 );
or ( n6422 , n4658 , n6420 , n6421 );
and ( n6423 , n4492 , n6422 );
and ( n6424 , n4490 , n6422 );
or ( n6425 , n4493 , n6423 , n6424 );
and ( n6426 , n4334 , n6425 );
and ( n6427 , n4332 , n6425 );
or ( n6428 , n4335 , n6426 , n6427 );
and ( n6429 , n4324 , n6428 );
xor ( n6430 , n4324 , n6428 );
xor ( n6431 , n4332 , n4334 );
xor ( n6432 , n6431 , n6425 );
xor ( n6433 , n4490 , n4492 );
xor ( n6434 , n6433 , n6422 );
xor ( n6435 , n4495 , n4657 );
xor ( n6436 , n6435 , n6419 );
xor ( n6437 , n4660 , n4799 );
xor ( n6438 , n6437 , n6416 );
xor ( n6439 , n4965 , n4967 );
xor ( n6440 , n6439 , n6413 );
xor ( n6441 , n4970 , n4988 );
xor ( n6442 , n6441 , n6410 );
xor ( n6443 , n4991 , n5233 );
xor ( n6444 , n6443 , n6407 );
xor ( n6445 , n5353 , n5355 );
xor ( n6446 , n6445 , n6404 );
xor ( n6447 , n5358 , n5376 );
xor ( n6448 , n6447 , n6401 );
xor ( n6449 , n5379 , n5527 );
xor ( n6450 , n6449 , n6398 );
xor ( n6451 , n5530 , n5639 );
xor ( n6452 , n6451 , n6395 );
xor ( n6453 , n5642 , n5750 );
xor ( n6454 , n6453 , n6392 );
xor ( n6455 , n5864 , n5866 );
xor ( n6456 , n6455 , n6389 );
xor ( n6457 , n5869 , n5967 );
xor ( n6458 , n6457 , n6386 );
xor ( n6459 , n5970 , n6019 );
xor ( n6460 , n6459 , n6383 );
xor ( n6461 , n6022 , n6164 );
xor ( n6462 , n6461 , n6380 );
xor ( n6463 , n6167 , n6193 );
xor ( n6464 , n6463 , n6377 );
xor ( n6465 , n6196 , n6251 );
xor ( n6466 , n6465 , n6374 );
xor ( n6467 , n6342 , n6368 );
xor ( n6468 , n6467 , n6371 );
and ( n6469 , n2390 , n4392 );
and ( n6470 , n2295 , n4389 );
nor ( n6471 , n6469 , n6470 );
xnor ( n6472 , n6471 , n3867 );
and ( n6473 , n2615 , n4107 );
and ( n6474 , n2506 , n4105 );
nor ( n6475 , n6473 , n6474 );
xnor ( n6476 , n6475 , n3870 );
and ( n6477 , n6472 , n6476 );
and ( n6478 , n6476 , n6300 );
and ( n6479 , n6472 , n6300 );
or ( n6480 , n6477 , n6478 , n6479 );
and ( n6481 , n2773 , n3742 );
and ( n6482 , n2697 , n3740 );
nor ( n6483 , n6481 , n6482 );
xnor ( n6484 , n6483 , n3538 );
and ( n6485 , n3813 , n2887 );
and ( n6486 , n3466 , n2885 );
nor ( n6487 , n6485 , n6486 );
xnor ( n6488 , n6487 , n2801 );
and ( n6489 , n6484 , n6488 );
and ( n6490 , n3859 , n2654 );
and ( n6491 , n3911 , n2652 );
nor ( n6492 , n6490 , n6491 );
xnor ( n6493 , n6492 , n2570 );
and ( n6494 , n6488 , n6493 );
and ( n6495 , n6484 , n6493 );
or ( n6496 , n6489 , n6494 , n6495 );
and ( n6497 , n6480 , n6496 );
and ( n6498 , n3052 , n3367 );
and ( n6499 , n2897 , n3365 );
nor ( n6500 , n6498 , n6499 );
xnor ( n6501 , n6500 , n3306 );
and ( n6502 , n3414 , n3093 );
and ( n6503 , n3136 , n3091 );
nor ( n6504 , n6502 , n6503 );
xnor ( n6505 , n6504 , n3027 );
and ( n6506 , n6501 , n6505 );
and ( n6507 , n4236 , n2483 );
and ( n6508 , n4099 , n2481 );
nor ( n6509 , n6507 , n6508 );
xnor ( n6510 , n6509 , n2418 );
and ( n6511 , n6505 , n6510 );
and ( n6512 , n6501 , n6510 );
or ( n6513 , n6506 , n6511 , n6512 );
and ( n6514 , n6496 , n6513 );
and ( n6515 , n6480 , n6513 );
or ( n6516 , n6497 , n6514 , n6515 );
xor ( n6517 , n6283 , n6287 );
xor ( n6518 , n6517 , n6292 );
xor ( n6519 , n6316 , n6320 );
xor ( n6520 , n6519 , n6325 );
and ( n6521 , n6518 , n6520 );
xor ( n6522 , n6299 , n6302 );
and ( n6523 , n3466 , n2887 );
and ( n6524 , n3414 , n2885 );
nor ( n6525 , n6523 , n6524 );
xnor ( n6526 , n6525 , n2801 );
xor ( n6527 , n6522 , n6526 );
and ( n6528 , n3911 , n2654 );
and ( n6529 , n3813 , n2652 );
nor ( n6530 , n6528 , n6529 );
xnor ( n6531 , n6530 , n2570 );
xor ( n6532 , n6527 , n6531 );
and ( n6533 , n6520 , n6532 );
and ( n6534 , n6518 , n6532 );
or ( n6535 , n6521 , n6533 , n6534 );
and ( n6536 , n6516 , n6535 );
and ( n6537 , n6522 , n6526 );
and ( n6538 , n6526 , n6531 );
and ( n6539 , n6522 , n6531 );
or ( n6540 , n6537 , n6538 , n6539 );
xor ( n6541 , n6480 , n6496 );
xor ( n6542 , n6541 , n6513 );
and ( n6543 , n2897 , n3742 );
and ( n6544 , n2773 , n3740 );
nor ( n6545 , n6543 , n6544 );
xnor ( n6546 , n6545 , n3538 );
and ( n6547 , n3466 , n3093 );
and ( n6548 , n3414 , n3091 );
nor ( n6549 , n6547 , n6548 );
xnor ( n6550 , n6549 , n3027 );
and ( n6551 , n6546 , n6550 );
and ( n6552 , n3911 , n2887 );
and ( n6553 , n3813 , n2885 );
nor ( n6554 , n6552 , n6553 );
xnor ( n6555 , n6554 , n2801 );
and ( n6556 , n6550 , n6555 );
and ( n6557 , n6546 , n6555 );
or ( n6558 , n6551 , n6556 , n6557 );
and ( n6559 , n2697 , n4107 );
and ( n6560 , n2615 , n4105 );
nor ( n6561 , n6559 , n6560 );
xnor ( n6562 , n6561 , n3870 );
and ( n6563 , n3136 , n3367 );
and ( n6564 , n3052 , n3365 );
nor ( n6565 , n6563 , n6564 );
xnor ( n6566 , n6565 , n3306 );
and ( n6567 , n6562 , n6566 );
and ( n6568 , n4402 , n2483 );
and ( n6569 , n4236 , n2481 );
nor ( n6570 , n6568 , n6569 );
xnor ( n6571 , n6570 , n2418 );
and ( n6572 , n6566 , n6571 );
and ( n6573 , n6562 , n6571 );
or ( n6574 , n6567 , n6572 , n6573 );
and ( n6575 , n6558 , n6574 );
and ( n6576 , n2506 , n4392 );
and ( n6577 , n2390 , n4389 );
nor ( n6578 , n6576 , n6577 );
xnor ( n6579 , n6578 , n3867 );
and ( n6580 , n4402 , n2481 );
not ( n6581 , n6580 );
and ( n6582 , n6581 , n2418 );
and ( n6583 , n6579 , n6582 );
and ( n6584 , n6574 , n6583 );
and ( n6585 , n6558 , n6583 );
or ( n6586 , n6575 , n6584 , n6585 );
and ( n6587 , n6542 , n6586 );
xor ( n6588 , n6472 , n6476 );
xor ( n6589 , n6588 , n6300 );
xor ( n6590 , n6484 , n6488 );
xor ( n6591 , n6590 , n6493 );
and ( n6592 , n6589 , n6591 );
xor ( n6593 , n6501 , n6505 );
xor ( n6594 , n6593 , n6510 );
and ( n6595 , n6591 , n6594 );
and ( n6596 , n6589 , n6594 );
or ( n6597 , n6592 , n6595 , n6596 );
and ( n6598 , n6586 , n6597 );
and ( n6599 , n6542 , n6597 );
or ( n6600 , n6587 , n6598 , n6599 );
and ( n6601 , n6540 , n6600 );
xor ( n6602 , n6346 , n6348 );
xor ( n6603 , n6602 , n6351 );
and ( n6604 , n6600 , n6603 );
and ( n6605 , n6540 , n6603 );
or ( n6606 , n6601 , n6604 , n6605 );
and ( n6607 , n6536 , n6606 );
xor ( n6608 , n6354 , n6356 );
xor ( n6609 , n6608 , n6359 );
and ( n6610 , n6606 , n6609 );
and ( n6611 , n6536 , n6609 );
or ( n6612 , n6607 , n6610 , n6611 );
xor ( n6613 , n6344 , n6362 );
xor ( n6614 , n6613 , n6365 );
and ( n6615 , n6612 , n6614 );
xor ( n6616 , n6612 , n6614 );
xor ( n6617 , n6516 , n6535 );
xor ( n6618 , n6518 , n6520 );
xor ( n6619 , n6618 , n6532 );
xor ( n6620 , n6579 , n6582 );
and ( n6621 , n2615 , n4392 );
and ( n6622 , n2506 , n4389 );
nor ( n6623 , n6621 , n6622 );
xnor ( n6624 , n6623 , n3867 );
and ( n6625 , n2773 , n4107 );
and ( n6626 , n2697 , n4105 );
nor ( n6627 , n6625 , n6626 );
xnor ( n6628 , n6627 , n3870 );
and ( n6629 , n6624 , n6628 );
and ( n6630 , n6628 , n6580 );
and ( n6631 , n6624 , n6580 );
or ( n6632 , n6629 , n6630 , n6631 );
and ( n6633 , n6620 , n6632 );
and ( n6634 , n4099 , n2654 );
and ( n6635 , n3859 , n2652 );
nor ( n6636 , n6634 , n6635 );
xnor ( n6637 , n6636 , n2570 );
and ( n6638 , n6632 , n6637 );
and ( n6639 , n6620 , n6637 );
or ( n6640 , n6633 , n6638 , n6639 );
and ( n6641 , n3052 , n3742 );
and ( n6642 , n2897 , n3740 );
nor ( n6643 , n6641 , n6642 );
xnor ( n6644 , n6643 , n3538 );
and ( n6645 , n3414 , n3367 );
and ( n6646 , n3136 , n3365 );
nor ( n6647 , n6645 , n6646 );
xnor ( n6648 , n6647 , n3306 );
and ( n6649 , n6644 , n6648 );
and ( n6650 , n3813 , n3093 );
and ( n6651 , n3466 , n3091 );
nor ( n6652 , n6650 , n6651 );
xnor ( n6653 , n6652 , n3027 );
and ( n6654 , n6648 , n6653 );
and ( n6655 , n6644 , n6653 );
or ( n6656 , n6649 , n6654 , n6655 );
xor ( n6657 , n6546 , n6550 );
xor ( n6658 , n6657 , n6555 );
and ( n6659 , n6656 , n6658 );
xor ( n6660 , n6562 , n6566 );
xor ( n6661 , n6660 , n6571 );
and ( n6662 , n6658 , n6661 );
and ( n6663 , n6656 , n6661 );
or ( n6664 , n6659 , n6662 , n6663 );
and ( n6665 , n6640 , n6664 );
xor ( n6666 , n6558 , n6574 );
xor ( n6667 , n6666 , n6583 );
and ( n6668 , n6664 , n6667 );
and ( n6669 , n6640 , n6667 );
or ( n6670 , n6665 , n6668 , n6669 );
and ( n6671 , n6619 , n6670 );
xor ( n6672 , n6542 , n6586 );
xor ( n6673 , n6672 , n6597 );
and ( n6674 , n6670 , n6673 );
and ( n6675 , n6619 , n6673 );
or ( n6676 , n6671 , n6674 , n6675 );
and ( n6677 , n6617 , n6676 );
xor ( n6678 , n6540 , n6600 );
xor ( n6679 , n6678 , n6603 );
and ( n6680 , n6676 , n6679 );
and ( n6681 , n6617 , n6679 );
or ( n6682 , n6677 , n6680 , n6681 );
xor ( n6683 , n6536 , n6606 );
xor ( n6684 , n6683 , n6609 );
and ( n6685 , n6682 , n6684 );
xor ( n6686 , n6682 , n6684 );
xor ( n6687 , n6617 , n6676 );
xor ( n6688 , n6687 , n6679 );
and ( n6689 , n2697 , n4392 );
and ( n6690 , n2615 , n4389 );
nor ( n6691 , n6689 , n6690 );
xnor ( n6692 , n6691 , n3867 );
and ( n6693 , n4402 , n2652 );
not ( n6694 , n6693 );
and ( n6695 , n6694 , n2570 );
and ( n6696 , n6692 , n6695 );
and ( n6697 , n3859 , n2887 );
and ( n6698 , n3911 , n2885 );
nor ( n6699 , n6697 , n6698 );
xnor ( n6700 , n6699 , n2801 );
and ( n6701 , n6696 , n6700 );
and ( n6702 , n4236 , n2654 );
and ( n6703 , n4099 , n2652 );
nor ( n6704 , n6702 , n6703 );
xnor ( n6705 , n6704 , n2570 );
and ( n6706 , n6700 , n6705 );
and ( n6707 , n6696 , n6705 );
or ( n6708 , n6701 , n6706 , n6707 );
and ( n6709 , n3136 , n3742 );
and ( n6710 , n3052 , n3740 );
nor ( n6711 , n6709 , n6710 );
xnor ( n6712 , n6711 , n3538 );
and ( n6713 , n4099 , n2887 );
and ( n6714 , n3859 , n2885 );
nor ( n6715 , n6713 , n6714 );
xnor ( n6716 , n6715 , n2801 );
and ( n6717 , n6712 , n6716 );
and ( n6718 , n4402 , n2654 );
and ( n6719 , n4236 , n2652 );
nor ( n6720 , n6718 , n6719 );
xnor ( n6721 , n6720 , n2570 );
and ( n6722 , n6716 , n6721 );
and ( n6723 , n6712 , n6721 );
or ( n6724 , n6717 , n6722 , n6723 );
and ( n6725 , n2897 , n4107 );
and ( n6726 , n2773 , n4105 );
nor ( n6727 , n6725 , n6726 );
xnor ( n6728 , n6727 , n3870 );
and ( n6729 , n3466 , n3367 );
and ( n6730 , n3414 , n3365 );
nor ( n6731 , n6729 , n6730 );
xnor ( n6732 , n6731 , n3306 );
and ( n6733 , n6728 , n6732 );
and ( n6734 , n3911 , n3093 );
and ( n6735 , n3813 , n3091 );
nor ( n6736 , n6734 , n6735 );
xnor ( n6737 , n6736 , n3027 );
and ( n6738 , n6732 , n6737 );
and ( n6739 , n6728 , n6737 );
or ( n6740 , n6733 , n6738 , n6739 );
and ( n6741 , n6724 , n6740 );
xor ( n6742 , n6624 , n6628 );
xor ( n6743 , n6742 , n6580 );
and ( n6744 , n6740 , n6743 );
and ( n6745 , n6724 , n6743 );
or ( n6746 , n6741 , n6744 , n6745 );
and ( n6747 , n6708 , n6746 );
xor ( n6748 , n6620 , n6632 );
xor ( n6749 , n6748 , n6637 );
and ( n6750 , n6746 , n6749 );
and ( n6751 , n6708 , n6749 );
or ( n6752 , n6747 , n6750 , n6751 );
xor ( n6753 , n6589 , n6591 );
xor ( n6754 , n6753 , n6594 );
and ( n6755 , n6752 , n6754 );
xor ( n6756 , n6640 , n6664 );
xor ( n6757 , n6756 , n6667 );
and ( n6758 , n6754 , n6757 );
and ( n6759 , n6752 , n6757 );
or ( n6760 , n6755 , n6758 , n6759 );
xor ( n6761 , n6619 , n6670 );
xor ( n6762 , n6761 , n6673 );
and ( n6763 , n6760 , n6762 );
xor ( n6764 , n6752 , n6754 );
xor ( n6765 , n6764 , n6757 );
xor ( n6766 , n6692 , n6695 );
and ( n6767 , n3052 , n4107 );
and ( n6768 , n2897 , n4105 );
nor ( n6769 , n6767 , n6768 );
xnor ( n6770 , n6769 , n3870 );
and ( n6771 , n3813 , n3367 );
and ( n6772 , n3466 , n3365 );
nor ( n6773 , n6771 , n6772 );
xnor ( n6774 , n6773 , n3306 );
and ( n6775 , n6770 , n6774 );
and ( n6776 , n6774 , n6693 );
and ( n6777 , n6770 , n6693 );
or ( n6778 , n6775 , n6776 , n6777 );
and ( n6779 , n6766 , n6778 );
and ( n6780 , n2773 , n4392 );
and ( n6781 , n2697 , n4389 );
nor ( n6782 , n6780 , n6781 );
xnor ( n6783 , n6782 , n3867 );
and ( n6784 , n3859 , n3093 );
and ( n6785 , n3911 , n3091 );
nor ( n6786 , n6784 , n6785 );
xnor ( n6787 , n6786 , n3027 );
and ( n6788 , n6783 , n6787 );
and ( n6789 , n4236 , n2887 );
and ( n6790 , n4099 , n2885 );
nor ( n6791 , n6789 , n6790 );
xnor ( n6792 , n6791 , n2801 );
and ( n6793 , n6787 , n6792 );
and ( n6794 , n6783 , n6792 );
or ( n6795 , n6788 , n6793 , n6794 );
and ( n6796 , n6778 , n6795 );
and ( n6797 , n6766 , n6795 );
or ( n6798 , n6779 , n6796 , n6797 );
xor ( n6799 , n6644 , n6648 );
xor ( n6800 , n6799 , n6653 );
and ( n6801 , n6798 , n6800 );
xor ( n6802 , n6696 , n6700 );
xor ( n6803 , n6802 , n6705 );
and ( n6804 , n6800 , n6803 );
and ( n6805 , n6798 , n6803 );
or ( n6806 , n6801 , n6804 , n6805 );
xor ( n6807 , n6656 , n6658 );
xor ( n6808 , n6807 , n6661 );
and ( n6809 , n6806 , n6808 );
xor ( n6810 , n6708 , n6746 );
xor ( n6811 , n6810 , n6749 );
and ( n6812 , n6808 , n6811 );
and ( n6813 , n6806 , n6811 );
or ( n6814 , n6809 , n6812 , n6813 );
and ( n6815 , n6765 , n6814 );
xor ( n6816 , n6806 , n6808 );
xor ( n6817 , n6816 , n6811 );
and ( n6818 , n2897 , n4392 );
and ( n6819 , n2773 , n4389 );
nor ( n6820 , n6818 , n6819 );
xnor ( n6821 , n6820 , n3867 );
and ( n6822 , n3911 , n3367 );
and ( n6823 , n3813 , n3365 );
nor ( n6824 , n6822 , n6823 );
xnor ( n6825 , n6824 , n3306 );
and ( n6826 , n6821 , n6825 );
and ( n6827 , n4099 , n3093 );
and ( n6828 , n3859 , n3091 );
nor ( n6829 , n6827 , n6828 );
xnor ( n6830 , n6829 , n3027 );
and ( n6831 , n6825 , n6830 );
and ( n6832 , n6821 , n6830 );
or ( n6833 , n6826 , n6831 , n6832 );
and ( n6834 , n3136 , n4107 );
and ( n6835 , n3052 , n4105 );
nor ( n6836 , n6834 , n6835 );
xnor ( n6837 , n6836 , n3870 );
and ( n6838 , n4402 , n2885 );
not ( n6839 , n6838 );
and ( n6840 , n6839 , n2801 );
and ( n6841 , n6837 , n6840 );
and ( n6842 , n6833 , n6841 );
and ( n6843 , n3414 , n3742 );
and ( n6844 , n3136 , n3740 );
nor ( n6845 , n6843 , n6844 );
xnor ( n6846 , n6845 , n3538 );
and ( n6847 , n6841 , n6846 );
and ( n6848 , n6833 , n6846 );
or ( n6849 , n6842 , n6847 , n6848 );
xor ( n6850 , n6712 , n6716 );
xor ( n6851 , n6850 , n6721 );
and ( n6852 , n6849 , n6851 );
xor ( n6853 , n6728 , n6732 );
xor ( n6854 , n6853 , n6737 );
and ( n6855 , n6851 , n6854 );
and ( n6856 , n6849 , n6854 );
or ( n6857 , n6852 , n6855 , n6856 );
xor ( n6858 , n6724 , n6740 );
xor ( n6859 , n6858 , n6743 );
and ( n6860 , n6857 , n6859 );
xor ( n6861 , n6798 , n6800 );
xor ( n6862 , n6861 , n6803 );
and ( n6863 , n6859 , n6862 );
and ( n6864 , n6857 , n6862 );
or ( n6865 , n6860 , n6863 , n6864 );
and ( n6866 , n6817 , n6865 );
xor ( n6867 , n6857 , n6859 );
xor ( n6868 , n6867 , n6862 );
xor ( n6869 , n6837 , n6840 );
and ( n6870 , n3466 , n3742 );
and ( n6871 , n3414 , n3740 );
nor ( n6872 , n6870 , n6871 );
xnor ( n6873 , n6872 , n3538 );
and ( n6874 , n6869 , n6873 );
and ( n6875 , n4402 , n2887 );
and ( n6876 , n4236 , n2885 );
nor ( n6877 , n6875 , n6876 );
xnor ( n6878 , n6877 , n2801 );
and ( n6879 , n6873 , n6878 );
and ( n6880 , n6869 , n6878 );
or ( n6881 , n6874 , n6879 , n6880 );
xor ( n6882 , n6770 , n6774 );
xor ( n6883 , n6882 , n6693 );
and ( n6884 , n6881 , n6883 );
xor ( n6885 , n6783 , n6787 );
xor ( n6886 , n6885 , n6792 );
and ( n6887 , n6883 , n6886 );
and ( n6888 , n6881 , n6886 );
or ( n6889 , n6884 , n6887 , n6888 );
xor ( n6890 , n6766 , n6778 );
xor ( n6891 , n6890 , n6795 );
and ( n6892 , n6889 , n6891 );
xor ( n6893 , n6849 , n6851 );
xor ( n6894 , n6893 , n6854 );
and ( n6895 , n6891 , n6894 );
and ( n6896 , n6889 , n6894 );
or ( n6897 , n6892 , n6895 , n6896 );
and ( n6898 , n6868 , n6897 );
xor ( n6899 , n6889 , n6891 );
xor ( n6900 , n6899 , n6894 );
xor ( n6901 , n6833 , n6841 );
xor ( n6902 , n6901 , n6846 );
xor ( n6903 , n6821 , n6825 );
xor ( n6904 , n6903 , n6830 );
and ( n6905 , n3052 , n4392 );
and ( n6906 , n2897 , n4389 );
nor ( n6907 , n6905 , n6906 );
xnor ( n6908 , n6907 , n3867 );
and ( n6909 , n4236 , n3093 );
and ( n6910 , n4099 , n3091 );
nor ( n6911 , n6909 , n6910 );
xnor ( n6912 , n6911 , n3027 );
and ( n6913 , n6908 , n6912 );
and ( n6914 , n6904 , n6913 );
and ( n6915 , n3414 , n4107 );
and ( n6916 , n3136 , n4105 );
nor ( n6917 , n6915 , n6916 );
xnor ( n6918 , n6917 , n3870 );
and ( n6919 , n3813 , n3742 );
and ( n6920 , n3466 , n3740 );
nor ( n6921 , n6919 , n6920 );
xnor ( n6922 , n6921 , n3538 );
and ( n6923 , n6918 , n6922 );
and ( n6924 , n3859 , n3367 );
and ( n6925 , n3911 , n3365 );
nor ( n6926 , n6924 , n6925 );
xnor ( n6927 , n6926 , n3306 );
and ( n6928 , n6922 , n6927 );
and ( n6929 , n6918 , n6927 );
or ( n6930 , n6923 , n6928 , n6929 );
and ( n6931 , n6913 , n6930 );
and ( n6932 , n6904 , n6930 );
or ( n6933 , n6914 , n6931 , n6932 );
and ( n6934 , n6902 , n6933 );
xor ( n6935 , n6881 , n6883 );
xor ( n6936 , n6935 , n6886 );
and ( n6937 , n6933 , n6936 );
and ( n6938 , n6902 , n6936 );
or ( n6939 , n6934 , n6937 , n6938 );
and ( n6940 , n6900 , n6939 );
xor ( n6941 , n6869 , n6873 );
xor ( n6942 , n6941 , n6878 );
xor ( n6943 , n6908 , n6912 );
and ( n6944 , n6838 , n6943 );
and ( n6945 , n3466 , n4107 );
and ( n6946 , n3414 , n4105 );
nor ( n6947 , n6945 , n6946 );
xnor ( n6948 , n6947 , n3870 );
and ( n6949 , n4402 , n3091 );
not ( n6950 , n6949 );
and ( n6951 , n6950 , n3027 );
and ( n6952 , n6948 , n6951 );
and ( n6953 , n6943 , n6952 );
and ( n6954 , n6838 , n6952 );
or ( n6955 , n6944 , n6953 , n6954 );
and ( n6956 , n6942 , n6955 );
xor ( n6957 , n6904 , n6913 );
xor ( n6958 , n6957 , n6930 );
and ( n6959 , n6955 , n6958 );
and ( n6960 , n6942 , n6958 );
or ( n6961 , n6956 , n6959 , n6960 );
xor ( n6962 , n6902 , n6933 );
xor ( n6963 , n6962 , n6936 );
and ( n6964 , n6961 , n6963 );
and ( n6965 , n3136 , n4392 );
and ( n6966 , n3052 , n4389 );
nor ( n6967 , n6965 , n6966 );
xnor ( n6968 , n6967 , n3867 );
and ( n6969 , n4099 , n3367 );
and ( n6970 , n3859 , n3365 );
nor ( n6971 , n6969 , n6970 );
xnor ( n6972 , n6971 , n3306 );
and ( n6973 , n6968 , n6972 );
and ( n6974 , n4402 , n3093 );
and ( n6975 , n4236 , n3091 );
nor ( n6976 , n6974 , n6975 );
xnor ( n6977 , n6976 , n3027 );
and ( n6978 , n6972 , n6977 );
and ( n6979 , n6968 , n6977 );
or ( n6980 , n6973 , n6978 , n6979 );
xor ( n6981 , n6918 , n6922 );
xor ( n6982 , n6981 , n6927 );
and ( n6983 , n6980 , n6982 );
xor ( n6984 , n6948 , n6951 );
and ( n6985 , n3414 , n4392 );
and ( n6986 , n3136 , n4389 );
nor ( n6987 , n6985 , n6986 );
xnor ( n6988 , n6987 , n3867 );
and ( n6989 , n4236 , n3367 );
and ( n6990 , n4099 , n3365 );
nor ( n6991 , n6989 , n6990 );
xnor ( n6992 , n6991 , n3306 );
and ( n6993 , n6988 , n6992 );
and ( n6994 , n6992 , n6949 );
and ( n6995 , n6988 , n6949 );
or ( n6996 , n6993 , n6994 , n6995 );
and ( n6997 , n6984 , n6996 );
and ( n6998 , n3911 , n3742 );
and ( n6999 , n3813 , n3740 );
nor ( n7000 , n6998 , n6999 );
xnor ( n7001 , n7000 , n3538 );
and ( n7002 , n6996 , n7001 );
and ( n7003 , n6984 , n7001 );
or ( n7004 , n6997 , n7002 , n7003 );
and ( n7005 , n6982 , n7004 );
and ( n7006 , n6980 , n7004 );
or ( n7007 , n6983 , n7005 , n7006 );
xor ( n7008 , n6942 , n6955 );
xor ( n7009 , n7008 , n6958 );
and ( n7010 , n7007 , n7009 );
xor ( n7011 , n6838 , n6943 );
xor ( n7012 , n7011 , n6952 );
xor ( n7013 , n6968 , n6972 );
xor ( n7014 , n7013 , n6977 );
xor ( n7015 , n6984 , n6996 );
xor ( n7016 , n7015 , n7001 );
and ( n7017 , n7014 , n7016 );
and ( n7018 , n3466 , n4392 );
and ( n7019 , n3414 , n4389 );
nor ( n7020 , n7018 , n7019 );
xnor ( n7021 , n7020 , n3867 );
and ( n7022 , n4402 , n3365 );
not ( n7023 , n7022 );
and ( n7024 , n7023 , n3306 );
and ( n7025 , n7021 , n7024 );
and ( n7026 , n3813 , n4107 );
and ( n7027 , n3466 , n4105 );
nor ( n7028 , n7026 , n7027 );
xnor ( n7029 , n7028 , n3870 );
and ( n7030 , n7025 , n7029 );
and ( n7031 , n3859 , n3742 );
and ( n7032 , n3911 , n3740 );
nor ( n7033 , n7031 , n7032 );
xnor ( n7034 , n7033 , n3538 );
and ( n7035 , n7029 , n7034 );
and ( n7036 , n7025 , n7034 );
or ( n7037 , n7030 , n7035 , n7036 );
and ( n7038 , n7016 , n7037 );
and ( n7039 , n7014 , n7037 );
or ( n7040 , n7017 , n7038 , n7039 );
and ( n7041 , n7012 , n7040 );
xor ( n7042 , n6980 , n6982 );
xor ( n7043 , n7042 , n7004 );
and ( n7044 , n7040 , n7043 );
and ( n7045 , n7012 , n7043 );
or ( n7046 , n7041 , n7044 , n7045 );
and ( n7047 , n7009 , n7046 );
and ( n7048 , n7007 , n7046 );
or ( n7049 , n7010 , n7047 , n7048 );
and ( n7050 , n6963 , n7049 );
and ( n7051 , n6961 , n7049 );
or ( n7052 , n6964 , n7050 , n7051 );
and ( n7053 , n6939 , n7052 );
and ( n7054 , n6900 , n7052 );
or ( n7055 , n6940 , n7053 , n7054 );
and ( n7056 , n6897 , n7055 );
and ( n7057 , n6868 , n7055 );
or ( n7058 , n6898 , n7056 , n7057 );
and ( n7059 , n6865 , n7058 );
and ( n7060 , n6817 , n7058 );
or ( n7061 , n6866 , n7059 , n7060 );
and ( n7062 , n6814 , n7061 );
and ( n7063 , n6765 , n7061 );
or ( n7064 , n6815 , n7062 , n7063 );
and ( n7065 , n6762 , n7064 );
and ( n7066 , n6760 , n7064 );
or ( n7067 , n6763 , n7065 , n7066 );
and ( n7068 , n6688 , n7067 );
xor ( n7069 , n6688 , n7067 );
xor ( n7070 , n6760 , n6762 );
xor ( n7071 , n7070 , n7064 );
xor ( n7072 , n6765 , n6814 );
xor ( n7073 , n7072 , n7061 );
xor ( n7074 , n6817 , n6865 );
xor ( n7075 , n7074 , n7058 );
xor ( n7076 , n6868 , n6897 );
xor ( n7077 , n7076 , n7055 );
xor ( n7078 , n6900 , n6939 );
xor ( n7079 , n7078 , n7052 );
xor ( n7080 , n6961 , n6963 );
xor ( n7081 , n7080 , n7049 );
xor ( n7082 , n7007 , n7009 );
xor ( n7083 , n7082 , n7046 );
xor ( n7084 , n7012 , n7040 );
xor ( n7085 , n7084 , n7043 );
and ( n7086 , n3911 , n4107 );
and ( n7087 , n3813 , n4105 );
nor ( n7088 , n7086 , n7087 );
xnor ( n7089 , n7088 , n3870 );
and ( n7090 , n4099 , n3742 );
and ( n7091 , n3859 , n3740 );
nor ( n7092 , n7090 , n7091 );
xnor ( n7093 , n7092 , n3538 );
and ( n7094 , n7089 , n7093 );
and ( n7095 , n4402 , n3367 );
and ( n7096 , n4236 , n3365 );
nor ( n7097 , n7095 , n7096 );
xnor ( n7098 , n7097 , n3306 );
and ( n7099 , n7093 , n7098 );
and ( n7100 , n7089 , n7098 );
or ( n7101 , n7094 , n7099 , n7100 );
xor ( n7102 , n6988 , n6992 );
xor ( n7103 , n7102 , n6949 );
and ( n7104 , n7101 , n7103 );
xor ( n7105 , n7025 , n7029 );
xor ( n7106 , n7105 , n7034 );
and ( n7107 , n7103 , n7106 );
and ( n7108 , n7101 , n7106 );
or ( n7109 , n7104 , n7107 , n7108 );
xor ( n7110 , n7014 , n7016 );
xor ( n7111 , n7110 , n7037 );
and ( n7112 , n7109 , n7111 );
xor ( n7113 , n7109 , n7111 );
xor ( n7114 , n7021 , n7024 );
and ( n7115 , n3813 , n4392 );
and ( n7116 , n3466 , n4389 );
nor ( n7117 , n7115 , n7116 );
xnor ( n7118 , n7117 , n3867 );
and ( n7119 , n3859 , n4107 );
and ( n7120 , n3911 , n4105 );
nor ( n7121 , n7119 , n7120 );
xnor ( n7122 , n7121 , n3870 );
and ( n7123 , n7118 , n7122 );
and ( n7124 , n7122 , n7022 );
and ( n7125 , n7118 , n7022 );
or ( n7126 , n7123 , n7124 , n7125 );
and ( n7127 , n7114 , n7126 );
xor ( n7128 , n7089 , n7093 );
xor ( n7129 , n7128 , n7098 );
and ( n7130 , n7126 , n7129 );
and ( n7131 , n7114 , n7129 );
or ( n7132 , n7127 , n7130 , n7131 );
xor ( n7133 , n7101 , n7103 );
xor ( n7134 , n7133 , n7106 );
and ( n7135 , n7132 , n7134 );
xor ( n7136 , n7132 , n7134 );
xor ( n7137 , n7114 , n7126 );
xor ( n7138 , n7137 , n7129 );
and ( n7139 , n3911 , n4392 );
and ( n7140 , n3813 , n4389 );
nor ( n7141 , n7139 , n7140 );
xnor ( n7142 , n7141 , n3867 );
and ( n7143 , n4402 , n3740 );
not ( n7144 , n7143 );
and ( n7145 , n7144 , n3538 );
and ( n7146 , n7142 , n7145 );
and ( n7147 , n4236 , n3742 );
and ( n7148 , n4099 , n3740 );
nor ( n7149 , n7147 , n7148 );
xnor ( n7150 , n7149 , n3538 );
and ( n7151 , n7146 , n7150 );
xor ( n7152 , n7118 , n7122 );
xor ( n7153 , n7152 , n7022 );
and ( n7154 , n7150 , n7153 );
and ( n7155 , n7146 , n7153 );
or ( n7156 , n7151 , n7154 , n7155 );
and ( n7157 , n7138 , n7156 );
xor ( n7158 , n7138 , n7156 );
xor ( n7159 , n7146 , n7150 );
xor ( n7160 , n7159 , n7153 );
xor ( n7161 , n7142 , n7145 );
and ( n7162 , n4099 , n4107 );
and ( n7163 , n3859 , n4105 );
nor ( n7164 , n7162 , n7163 );
xnor ( n7165 , n7164 , n3870 );
and ( n7166 , n7161 , n7165 );
and ( n7167 , n4402 , n3742 );
and ( n7168 , n4236 , n3740 );
nor ( n7169 , n7167 , n7168 );
xnor ( n7170 , n7169 , n3538 );
and ( n7171 , n7165 , n7170 );
and ( n7172 , n7161 , n7170 );
or ( n7173 , n7166 , n7171 , n7172 );
and ( n7174 , n7160 , n7173 );
xor ( n7175 , n7160 , n7173 );
and ( n7176 , n3859 , n4392 );
and ( n7177 , n3911 , n4389 );
nor ( n7178 , n7176 , n7177 );
xnor ( n7179 , n7178 , n3867 );
and ( n7180 , n4236 , n4107 );
and ( n7181 , n4099 , n4105 );
nor ( n7182 , n7180 , n7181 );
xnor ( n7183 , n7182 , n3870 );
and ( n7184 , n7179 , n7183 );
and ( n7185 , n7183 , n7143 );
and ( n7186 , n7179 , n7143 );
or ( n7187 , n7184 , n7185 , n7186 );
xor ( n7188 , n7161 , n7165 );
xor ( n7189 , n7188 , n7170 );
and ( n7190 , n7187 , n7189 );
xor ( n7191 , n7187 , n7189 );
xor ( n7192 , n7179 , n7183 );
xor ( n7193 , n7192 , n7143 );
and ( n7194 , n4099 , n4392 );
and ( n7195 , n3859 , n4389 );
nor ( n7196 , n7194 , n7195 );
xnor ( n7197 , n7196 , n3867 );
and ( n7198 , n4402 , n4105 );
not ( n7199 , n7198 );
and ( n7200 , n7199 , n3870 );
and ( n7201 , n7197 , n7200 );
and ( n7202 , n7193 , n7201 );
xor ( n7203 , n7193 , n7201 );
and ( n7204 , n4402 , n4107 );
and ( n7205 , n4236 , n4105 );
nor ( n7206 , n7204 , n7205 );
xnor ( n7207 , n7206 , n3870 );
xor ( n7208 , n7197 , n7200 );
and ( n7209 , n7207 , n7208 );
xor ( n7210 , n7207 , n7208 );
and ( n7211 , n4236 , n4392 );
and ( n7212 , n4099 , n4389 );
nor ( n7213 , n7211 , n7212 );
xnor ( n7214 , n7213 , n3867 );
and ( n7215 , n7214 , n7198 );
xor ( n7216 , n7214 , n7198 );
and ( n7217 , n4402 , n4392 );
and ( n7218 , n4236 , n4389 );
nor ( n7219 , n7217 , n7218 );
xnor ( n7220 , n7219 , n3867 );
and ( n7221 , n4402 , n4389 );
not ( n7222 , n7221 );
and ( n7223 , n7222 , n3867 );
and ( n7224 , n7220 , n7223 );
and ( n7225 , n7216 , n7224 );
or ( n7226 , n7215 , n7225 );
and ( n7227 , n7210 , n7226 );
or ( n7228 , n7209 , n7227 );
and ( n7229 , n7203 , n7228 );
or ( n7230 , n7202 , n7229 );
and ( n7231 , n7191 , n7230 );
or ( n7232 , n7190 , n7231 );
and ( n7233 , n7175 , n7232 );
or ( n7234 , n7174 , n7233 );
and ( n7235 , n7158 , n7234 );
or ( n7236 , n7157 , n7235 );
and ( n7237 , n7136 , n7236 );
or ( n7238 , n7135 , n7237 );
and ( n7239 , n7113 , n7238 );
or ( n7240 , n7112 , n7239 );
and ( n7241 , n7085 , n7240 );
and ( n7242 , n7083 , n7241 );
and ( n7243 , n7081 , n7242 );
and ( n7244 , n7079 , n7243 );
and ( n7245 , n7077 , n7244 );
and ( n7246 , n7075 , n7245 );
and ( n7247 , n7073 , n7246 );
and ( n7248 , n7071 , n7247 );
and ( n7249 , n7069 , n7248 );
or ( n7250 , n7068 , n7249 );
and ( n7251 , n6686 , n7250 );
or ( n7252 , n6685 , n7251 );
and ( n7253 , n6616 , n7252 );
or ( n7254 , n6615 , n7253 );
and ( n7255 , n6468 , n7254 );
and ( n7256 , n6466 , n7255 );
and ( n7257 , n6464 , n7256 );
and ( n7258 , n6462 , n7257 );
and ( n7259 , n6460 , n7258 );
and ( n7260 , n6458 , n7259 );
and ( n7261 , n6456 , n7260 );
and ( n7262 , n6454 , n7261 );
and ( n7263 , n6452 , n7262 );
and ( n7264 , n6450 , n7263 );
and ( n7265 , n6448 , n7264 );
and ( n7266 , n6446 , n7265 );
and ( n7267 , n6444 , n7266 );
and ( n7268 , n6442 , n7267 );
and ( n7269 , n6440 , n7268 );
and ( n7270 , n6438 , n7269 );
and ( n7271 , n6436 , n7270 );
and ( n7272 , n6434 , n7271 );
and ( n7273 , n6432 , n7272 );
and ( n7274 , n6430 , n7273 );
or ( n7275 , n6429 , n7274 );
and ( n7276 , n4322 , n7275 );
or ( n7277 , n4321 , n7276 );
and ( n7278 , n4025 , n7277 );
or ( n7279 , n4024 , n7278 );
and ( n7280 , n3695 , n7279 );
and ( n7281 , n3693 , n7280 );
and ( n7282 , n3691 , n7281 );
and ( n7283 , n3689 , n7282 );
and ( n7284 , n3687 , n7283 );
and ( n7285 , n3685 , n7284 );
and ( n7286 , n3683 , n7285 );
and ( n7287 , n3681 , n7286 );
and ( n7288 , n3679 , n7287 );
and ( n7289 , n3677 , n7288 );
and ( n7290 , n3675 , n7289 );
and ( n7291 , n3673 , n7290 );
and ( n7292 , n3671 , n7291 );
and ( n7293 , n3669 , n7292 );
and ( n7294 , n3667 , n7293 );
and ( n7295 , n3665 , n7294 );
and ( n7296 , n3663 , n7295 );
and ( n7297 , n3661 , n7296 );
xor ( n7298 , n3659 , n7297 );
buf ( n7299 , n7298 );
buf ( n7300 , n7299 );
buf ( n7301 , n7300 );
buf ( n7302 , n1147 );
buf ( n7303 , n1120 );
xor ( n7304 , n7302 , n7303 );
buf ( n7305 , n1148 );
buf ( n7306 , n1121 );
and ( n7307 , n7305 , n7306 );
xor ( n7308 , n7304 , n7307 );
buf ( n7309 , n7308 );
buf ( n7310 , n7309 );
buf ( n7311 , n7310 );
xor ( n7312 , n7305 , n7306 );
buf ( n7313 , n7312 );
buf ( n7314 , n7313 );
buf ( n7315 , n7314 );
xor ( n7316 , n7311 , n7315 );
not ( n7317 , n7315 );
and ( n7318 , n7316 , n7317 );
and ( n7319 , n7301 , n7318 );
and ( n7320 , n1682 , n1686 );
and ( n7321 , n1686 , n1688 );
and ( n7322 , n1682 , n1688 );
or ( n7323 , n7320 , n7321 , n7322 );
and ( n7324 , n1636 , n1663 );
not ( n7325 , n7324 );
xnor ( n7326 , n7325 , n1671 );
xor ( n7327 , n7323 , n7326 );
and ( n7328 , n1666 , n1657 );
not ( n7329 , n7328 );
xor ( n7330 , n7327 , n7329 );
and ( n7331 , n1679 , n1680 );
and ( n7332 , n1680 , n1689 );
and ( n7333 , n1679 , n1689 );
or ( n7334 , n7331 , n7332 , n7333 );
xor ( n7335 , n7330 , n7334 );
and ( n7336 , n1690 , n1746 );
and ( n7337 , n1746 , n3658 );
and ( n7338 , n1690 , n3658 );
or ( n7339 , n7336 , n7337 , n7338 );
xor ( n7340 , n7335 , n7339 );
and ( n7341 , n3659 , n7297 );
xor ( n7342 , n7340 , n7341 );
buf ( n7343 , n7342 );
buf ( n7344 , n7343 );
buf ( n7345 , n7344 );
and ( n7346 , n7345 , n7315 );
nor ( n7347 , n7319 , n7346 );
xnor ( n7348 , n7347 , n7311 );
xor ( n7349 , n3669 , n7292 );
buf ( n7350 , n7349 );
buf ( n7351 , n7350 );
buf ( n7352 , n7351 );
buf ( n7353 , n1143 );
buf ( n7354 , n1116 );
xor ( n7355 , n7353 , n7354 );
buf ( n7356 , n1144 );
buf ( n7357 , n1117 );
and ( n7358 , n7356 , n7357 );
buf ( n7359 , n1145 );
buf ( n7360 , n1118 );
and ( n7361 , n7359 , n7360 );
buf ( n7362 , n1146 );
buf ( n7363 , n1119 );
and ( n7364 , n7362 , n7363 );
and ( n7365 , n7302 , n7303 );
and ( n7366 , n7303 , n7307 );
and ( n7367 , n7302 , n7307 );
or ( n7368 , n7365 , n7366 , n7367 );
and ( n7369 , n7363 , n7368 );
and ( n7370 , n7362 , n7368 );
or ( n7371 , n7364 , n7369 , n7370 );
and ( n7372 , n7360 , n7371 );
and ( n7373 , n7359 , n7371 );
or ( n7374 , n7361 , n7372 , n7373 );
and ( n7375 , n7357 , n7374 );
and ( n7376 , n7356 , n7374 );
or ( n7377 , n7358 , n7375 , n7376 );
xor ( n7378 , n7355 , n7377 );
buf ( n7379 , n7378 );
buf ( n7380 , n7379 );
buf ( n7381 , n7380 );
xor ( n7382 , n7356 , n7357 );
xor ( n7383 , n7382 , n7374 );
buf ( n7384 , n7383 );
buf ( n7385 , n7384 );
buf ( n7386 , n7385 );
xor ( n7387 , n7381 , n7386 );
xor ( n7388 , n7359 , n7360 );
xor ( n7389 , n7388 , n7371 );
buf ( n7390 , n7389 );
buf ( n7391 , n7390 );
buf ( n7392 , n7391 );
xor ( n7393 , n7386 , n7392 );
not ( n7394 , n7393 );
and ( n7395 , n7387 , n7394 );
and ( n7396 , n7352 , n7395 );
xor ( n7397 , n3667 , n7293 );
buf ( n7398 , n7397 );
buf ( n7399 , n7398 );
buf ( n7400 , n7399 );
and ( n7401 , n7400 , n7393 );
nor ( n7402 , n7396 , n7401 );
and ( n7403 , n7386 , n7392 );
not ( n7404 , n7403 );
and ( n7405 , n7381 , n7404 );
xnor ( n7406 , n7402 , n7405 );
xor ( n7407 , n3693 , n7280 );
buf ( n7408 , n7407 );
buf ( n7409 , n7408 );
buf ( n7410 , n7409 );
buf ( n7411 , n1131 );
buf ( n7412 , n1104 );
xor ( n7413 , n7411 , n7412 );
buf ( n7414 , n1132 );
buf ( n7415 , n1105 );
and ( n7416 , n7414 , n7415 );
buf ( n7417 , n1133 );
buf ( n7418 , n1106 );
and ( n7419 , n7417 , n7418 );
buf ( n7420 , n1134 );
buf ( n7421 , n1107 );
and ( n7422 , n7420 , n7421 );
buf ( n7423 , n1135 );
buf ( n7424 , n1108 );
and ( n7425 , n7423 , n7424 );
buf ( n7426 , n1136 );
buf ( n7427 , n1109 );
and ( n7428 , n7426 , n7427 );
buf ( n7429 , n1137 );
buf ( n7430 , n1110 );
and ( n7431 , n7429 , n7430 );
buf ( n7432 , n1138 );
buf ( n7433 , n1111 );
and ( n7434 , n7432 , n7433 );
buf ( n7435 , n1139 );
buf ( n7436 , n1112 );
and ( n7437 , n7435 , n7436 );
buf ( n7438 , n1140 );
buf ( n7439 , n1113 );
and ( n7440 , n7438 , n7439 );
buf ( n7441 , n1141 );
buf ( n7442 , n1114 );
and ( n7443 , n7441 , n7442 );
buf ( n7444 , n1142 );
buf ( n7445 , n1115 );
and ( n7446 , n7444 , n7445 );
and ( n7447 , n7353 , n7354 );
and ( n7448 , n7354 , n7377 );
and ( n7449 , n7353 , n7377 );
or ( n7450 , n7447 , n7448 , n7449 );
and ( n7451 , n7445 , n7450 );
and ( n7452 , n7444 , n7450 );
or ( n7453 , n7446 , n7451 , n7452 );
and ( n7454 , n7442 , n7453 );
and ( n7455 , n7441 , n7453 );
or ( n7456 , n7443 , n7454 , n7455 );
and ( n7457 , n7439 , n7456 );
and ( n7458 , n7438 , n7456 );
or ( n7459 , n7440 , n7457 , n7458 );
and ( n7460 , n7436 , n7459 );
and ( n7461 , n7435 , n7459 );
or ( n7462 , n7437 , n7460 , n7461 );
and ( n7463 , n7433 , n7462 );
and ( n7464 , n7432 , n7462 );
or ( n7465 , n7434 , n7463 , n7464 );
and ( n7466 , n7430 , n7465 );
and ( n7467 , n7429 , n7465 );
or ( n7468 , n7431 , n7466 , n7467 );
and ( n7469 , n7427 , n7468 );
and ( n7470 , n7426 , n7468 );
or ( n7471 , n7428 , n7469 , n7470 );
and ( n7472 , n7424 , n7471 );
and ( n7473 , n7423 , n7471 );
or ( n7474 , n7425 , n7472 , n7473 );
and ( n7475 , n7421 , n7474 );
and ( n7476 , n7420 , n7474 );
or ( n7477 , n7422 , n7475 , n7476 );
and ( n7478 , n7418 , n7477 );
and ( n7479 , n7417 , n7477 );
or ( n7480 , n7419 , n7478 , n7479 );
and ( n7481 , n7415 , n7480 );
and ( n7482 , n7414 , n7480 );
or ( n7483 , n7416 , n7481 , n7482 );
xor ( n7484 , n7413 , n7483 );
buf ( n7485 , n7484 );
buf ( n7486 , n7485 );
buf ( n7487 , n7486 );
xor ( n7488 , n7414 , n7415 );
xor ( n7489 , n7488 , n7480 );
buf ( n7490 , n7489 );
buf ( n7491 , n7490 );
buf ( n7492 , n7491 );
xor ( n7493 , n7487 , n7492 );
xor ( n7494 , n7417 , n7418 );
xor ( n7495 , n7494 , n7477 );
buf ( n7496 , n7495 );
buf ( n7497 , n7496 );
buf ( n7498 , n7497 );
xor ( n7499 , n7492 , n7498 );
not ( n7500 , n7499 );
and ( n7501 , n7493 , n7500 );
and ( n7502 , n7410 , n7501 );
xor ( n7503 , n3691 , n7281 );
buf ( n7504 , n7503 );
buf ( n7505 , n7504 );
buf ( n7506 , n7505 );
and ( n7507 , n7506 , n7499 );
nor ( n7508 , n7502 , n7507 );
and ( n7509 , n7492 , n7498 );
not ( n7510 , n7509 );
and ( n7511 , n7487 , n7510 );
xnor ( n7512 , n7508 , n7511 );
xor ( n7513 , n4025 , n7277 );
buf ( n7514 , n7513 );
buf ( n7515 , n7514 );
buf ( n7516 , n7515 );
buf ( n7517 , n1129 );
buf ( n7518 , n1102 );
xor ( n7519 , n7517 , n7518 );
buf ( n7520 , n1130 );
buf ( n7521 , n1103 );
and ( n7522 , n7520 , n7521 );
and ( n7523 , n7411 , n7412 );
and ( n7524 , n7412 , n7483 );
and ( n7525 , n7411 , n7483 );
or ( n7526 , n7523 , n7524 , n7525 );
and ( n7527 , n7521 , n7526 );
and ( n7528 , n7520 , n7526 );
or ( n7529 , n7522 , n7527 , n7528 );
xor ( n7530 , n7519 , n7529 );
buf ( n7531 , n7530 );
buf ( n7532 , n7531 );
buf ( n7533 , n7532 );
xor ( n7534 , n7520 , n7521 );
xor ( n7535 , n7534 , n7526 );
buf ( n7536 , n7535 );
buf ( n7537 , n7536 );
buf ( n7538 , n7537 );
xor ( n7539 , n7533 , n7538 );
xor ( n7540 , n7538 , n7487 );
not ( n7541 , n7540 );
and ( n7542 , n7539 , n7541 );
and ( n7543 , n7516 , n7542 );
xor ( n7544 , n3695 , n7279 );
buf ( n7545 , n7544 );
buf ( n7546 , n7545 );
buf ( n7547 , n7546 );
and ( n7548 , n7547 , n7540 );
nor ( n7549 , n7543 , n7548 );
and ( n7550 , n7538 , n7487 );
not ( n7551 , n7550 );
and ( n7552 , n7533 , n7551 );
xnor ( n7553 , n7549 , n7552 );
xor ( n7554 , n7512 , n7553 );
xor ( n7555 , n6434 , n7271 );
buf ( n7556 , n7555 );
buf ( n7557 , n7556 );
buf ( n7558 , n7557 );
buf ( n7559 , n1125 );
buf ( n7560 , n1098 );
xor ( n7561 , n7559 , n7560 );
buf ( n7562 , n1126 );
buf ( n7563 , n1099 );
and ( n7564 , n7562 , n7563 );
buf ( n7565 , n1127 );
buf ( n7566 , n1100 );
and ( n7567 , n7565 , n7566 );
buf ( n7568 , n1128 );
buf ( n7569 , n1101 );
and ( n7570 , n7568 , n7569 );
and ( n7571 , n7517 , n7518 );
and ( n7572 , n7518 , n7529 );
and ( n7573 , n7517 , n7529 );
or ( n7574 , n7571 , n7572 , n7573 );
and ( n7575 , n7569 , n7574 );
and ( n7576 , n7568 , n7574 );
or ( n7577 , n7570 , n7575 , n7576 );
and ( n7578 , n7566 , n7577 );
and ( n7579 , n7565 , n7577 );
or ( n7580 , n7567 , n7578 , n7579 );
and ( n7581 , n7563 , n7580 );
and ( n7582 , n7562 , n7580 );
or ( n7583 , n7564 , n7581 , n7582 );
xor ( n7584 , n7561 , n7583 );
buf ( n7585 , n7584 );
buf ( n7586 , n7585 );
buf ( n7587 , n7586 );
xor ( n7588 , n7562 , n7563 );
xor ( n7589 , n7588 , n7580 );
buf ( n7590 , n7589 );
buf ( n7591 , n7590 );
buf ( n7592 , n7591 );
xor ( n7593 , n7587 , n7592 );
xor ( n7594 , n7565 , n7566 );
xor ( n7595 , n7594 , n7577 );
buf ( n7596 , n7595 );
buf ( n7597 , n7596 );
buf ( n7598 , n7597 );
xor ( n7599 , n7592 , n7598 );
not ( n7600 , n7599 );
and ( n7601 , n7593 , n7600 );
and ( n7602 , n7558 , n7601 );
xor ( n7603 , n6432 , n7272 );
buf ( n7604 , n7603 );
buf ( n7605 , n7604 );
buf ( n7606 , n7605 );
and ( n7607 , n7606 , n7599 );
nor ( n7608 , n7602 , n7607 );
and ( n7609 , n7592 , n7598 );
not ( n7610 , n7609 );
and ( n7611 , n7587 , n7610 );
xnor ( n7612 , n7608 , n7611 );
xor ( n7613 , n7554 , n7612 );
and ( n7614 , n7406 , n7613 );
xor ( n7615 , n6446 , n7265 );
buf ( n7616 , n7615 );
buf ( n7617 , n7616 );
buf ( n7618 , n7617 );
buf ( n7619 , n1092 );
buf ( n7620 , n1093 );
buf ( n7621 , n1094 );
buf ( n7622 , n1122 );
buf ( n7623 , n1095 );
and ( n7624 , n7622 , n7623 );
buf ( n7625 , n1123 );
buf ( n7626 , n1096 );
and ( n7627 , n7625 , n7626 );
buf ( n7628 , n1124 );
buf ( n7629 , n1097 );
and ( n7630 , n7628 , n7629 );
and ( n7631 , n7559 , n7560 );
and ( n7632 , n7560 , n7583 );
and ( n7633 , n7559 , n7583 );
or ( n7634 , n7631 , n7632 , n7633 );
and ( n7635 , n7629 , n7634 );
and ( n7636 , n7628 , n7634 );
or ( n7637 , n7630 , n7635 , n7636 );
and ( n7638 , n7626 , n7637 );
and ( n7639 , n7625 , n7637 );
or ( n7640 , n7627 , n7638 , n7639 );
and ( n7641 , n7623 , n7640 );
and ( n7642 , n7622 , n7640 );
or ( n7643 , n7624 , n7641 , n7642 );
and ( n7644 , n7621 , n7643 );
and ( n7645 , n7620 , n7644 );
xor ( n7646 , n7619 , n7645 );
buf ( n7647 , n7646 );
buf ( n7648 , n7647 );
buf ( n7649 , n7648 );
xor ( n7650 , n7620 , n7644 );
buf ( n7651 , n7650 );
buf ( n7652 , n7651 );
buf ( n7653 , n7652 );
xor ( n7654 , n7649 , n7653 );
xor ( n7655 , n7621 , n7643 );
buf ( n7656 , n7655 );
buf ( n7657 , n7656 );
buf ( n7658 , n7657 );
xor ( n7659 , n7653 , n7658 );
not ( n7660 , n7659 );
and ( n7661 , n7654 , n7660 );
and ( n7662 , n7618 , n7661 );
xor ( n7663 , n6444 , n7266 );
buf ( n7664 , n7663 );
buf ( n7665 , n7664 );
buf ( n7666 , n7665 );
and ( n7667 , n7666 , n7659 );
nor ( n7668 , n7662 , n7667 );
and ( n7669 , n7653 , n7658 );
not ( n7670 , n7669 );
and ( n7671 , n7649 , n7670 );
xnor ( n7672 , n7668 , n7671 );
xor ( n7673 , n6454 , n7261 );
buf ( n7674 , n7673 );
buf ( n7675 , n7674 );
buf ( n7676 , n7675 );
buf ( n7677 , n1090 );
buf ( n7678 , n1091 );
and ( n7679 , n7619 , n7645 );
and ( n7680 , n7678 , n7679 );
and ( n7681 , n7677 , n7680 );
buf ( n7682 , n7681 );
buf ( n7683 , n7682 );
buf ( n7684 , n7683 );
xor ( n7685 , n7677 , n7680 );
buf ( n7686 , n7685 );
buf ( n7687 , n7686 );
buf ( n7688 , n7687 );
xor ( n7689 , n7684 , n7688 );
not ( n7690 , n7689 );
and ( n7691 , n7684 , n7690 );
and ( n7692 , n7676 , n7691 );
xor ( n7693 , n6452 , n7262 );
buf ( n7694 , n7693 );
buf ( n7695 , n7694 );
buf ( n7696 , n7695 );
and ( n7697 , n7696 , n7689 );
nor ( n7698 , n7692 , n7697 );
not ( n7699 , n7698 );
xor ( n7700 , n7672 , n7699 );
xor ( n7701 , n6430 , n7273 );
buf ( n7702 , n7701 );
buf ( n7703 , n7702 );
buf ( n7704 , n7703 );
xor ( n7705 , n7568 , n7569 );
xor ( n7706 , n7705 , n7574 );
buf ( n7707 , n7706 );
buf ( n7708 , n7707 );
buf ( n7709 , n7708 );
xor ( n7710 , n7598 , n7709 );
xor ( n7711 , n7709 , n7533 );
not ( n7712 , n7711 );
and ( n7713 , n7710 , n7712 );
and ( n7714 , n7704 , n7713 );
xor ( n7715 , n4322 , n7275 );
buf ( n7716 , n7715 );
buf ( n7717 , n7716 );
buf ( n7718 , n7717 );
and ( n7719 , n7718 , n7711 );
nor ( n7720 , n7714 , n7719 );
and ( n7721 , n7709 , n7533 );
not ( n7722 , n7721 );
and ( n7723 , n7598 , n7722 );
xnor ( n7724 , n7720 , n7723 );
xor ( n7725 , n7700 , n7724 );
xor ( n7726 , n6438 , n7269 );
buf ( n7727 , n7726 );
buf ( n7728 , n7727 );
buf ( n7729 , n7728 );
xor ( n7730 , n7625 , n7626 );
xor ( n7731 , n7730 , n7637 );
buf ( n7732 , n7731 );
buf ( n7733 , n7732 );
buf ( n7734 , n7733 );
xor ( n7735 , n7628 , n7629 );
xor ( n7736 , n7735 , n7634 );
buf ( n7737 , n7736 );
buf ( n7738 , n7737 );
buf ( n7739 , n7738 );
xor ( n7740 , n7734 , n7739 );
xor ( n7741 , n7739 , n7587 );
not ( n7742 , n7741 );
and ( n7743 , n7740 , n7742 );
and ( n7744 , n7729 , n7743 );
xor ( n7745 , n6436 , n7270 );
buf ( n7746 , n7745 );
buf ( n7747 , n7746 );
buf ( n7748 , n7747 );
and ( n7749 , n7748 , n7741 );
nor ( n7750 , n7744 , n7749 );
and ( n7751 , n7739 , n7587 );
not ( n7752 , n7751 );
and ( n7753 , n7734 , n7752 );
xnor ( n7754 , n7750 , n7753 );
xor ( n7755 , n7725 , n7754 );
and ( n7756 , n7613 , n7755 );
and ( n7757 , n7406 , n7755 );
or ( n7758 , n7614 , n7756 , n7757 );
xor ( n7759 , n3683 , n7285 );
buf ( n7760 , n7759 );
buf ( n7761 , n7760 );
buf ( n7762 , n7761 );
xor ( n7763 , n7429 , n7430 );
xor ( n7764 , n7763 , n7465 );
buf ( n7765 , n7764 );
buf ( n7766 , n7765 );
buf ( n7767 , n7766 );
xor ( n7768 , n7432 , n7433 );
xor ( n7769 , n7768 , n7462 );
buf ( n7770 , n7769 );
buf ( n7771 , n7770 );
buf ( n7772 , n7771 );
xor ( n7773 , n7767 , n7772 );
xor ( n7774 , n7435 , n7436 );
xor ( n7775 , n7774 , n7459 );
buf ( n7776 , n7775 );
buf ( n7777 , n7776 );
buf ( n7778 , n7777 );
xor ( n7779 , n7772 , n7778 );
not ( n7780 , n7779 );
and ( n7781 , n7773 , n7780 );
and ( n7782 , n7762 , n7781 );
xor ( n7783 , n3681 , n7286 );
buf ( n7784 , n7783 );
buf ( n7785 , n7784 );
buf ( n7786 , n7785 );
and ( n7787 , n7786 , n7779 );
nor ( n7788 , n7782 , n7787 );
and ( n7789 , n7772 , n7778 );
not ( n7790 , n7789 );
and ( n7791 , n7767 , n7790 );
xnor ( n7792 , n7788 , n7791 );
and ( n7793 , n7547 , n7501 );
and ( n7794 , n7410 , n7499 );
nor ( n7795 , n7793 , n7794 );
xnor ( n7796 , n7795 , n7511 );
xor ( n7797 , n6440 , n7268 );
buf ( n7798 , n7797 );
buf ( n7799 , n7798 );
buf ( n7800 , n7799 );
and ( n7801 , n7800 , n7743 );
and ( n7802 , n7729 , n7741 );
nor ( n7803 , n7801 , n7802 );
xnor ( n7804 , n7803 , n7753 );
xor ( n7805 , n7796 , n7804 );
xor ( n7806 , n6448 , n7264 );
buf ( n7807 , n7806 );
buf ( n7808 , n7807 );
buf ( n7809 , n7808 );
and ( n7810 , n7809 , n7661 );
and ( n7811 , n7618 , n7659 );
nor ( n7812 , n7810 , n7811 );
xnor ( n7813 , n7812 , n7671 );
xor ( n7814 , n7805 , n7813 );
and ( n7815 , n7792 , n7814 );
xor ( n7816 , n7678 , n7679 );
buf ( n7817 , n7816 );
buf ( n7818 , n7817 );
buf ( n7819 , n7818 );
xor ( n7820 , n7688 , n7819 );
xor ( n7821 , n7819 , n7649 );
not ( n7822 , n7821 );
and ( n7823 , n7820 , n7822 );
and ( n7824 , n7696 , n7823 );
xor ( n7825 , n6450 , n7263 );
buf ( n7826 , n7825 );
buf ( n7827 , n7826 );
buf ( n7828 , n7827 );
and ( n7829 , n7828 , n7821 );
nor ( n7830 , n7824 , n7829 );
and ( n7831 , n7819 , n7649 );
not ( n7832 , n7831 );
and ( n7833 , n7688 , n7832 );
xnor ( n7834 , n7830 , n7833 );
xor ( n7835 , n6456 , n7260 );
buf ( n7836 , n7835 );
buf ( n7837 , n7836 );
buf ( n7838 , n7837 );
and ( n7839 , n7838 , n7691 );
and ( n7840 , n7676 , n7689 );
nor ( n7841 , n7839 , n7840 );
not ( n7842 , n7841 );
xor ( n7843 , n7834 , n7842 );
and ( n7844 , n7676 , n7823 );
and ( n7845 , n7696 , n7821 );
nor ( n7846 , n7844 , n7845 );
xnor ( n7847 , n7846 , n7833 );
xor ( n7848 , n6458 , n7259 );
buf ( n7849 , n7848 );
buf ( n7850 , n7849 );
buf ( n7851 , n7850 );
and ( n7852 , n7851 , n7691 );
and ( n7853 , n7838 , n7689 );
nor ( n7854 , n7852 , n7853 );
not ( n7855 , n7854 );
and ( n7856 , n7847 , n7855 );
xor ( n7857 , n7843 , n7856 );
xor ( n7858 , n7622 , n7623 );
xor ( n7859 , n7858 , n7640 );
buf ( n7860 , n7859 );
buf ( n7861 , n7860 );
buf ( n7862 , n7861 );
xor ( n7863 , n7658 , n7862 );
xor ( n7864 , n7862 , n7734 );
not ( n7865 , n7864 );
and ( n7866 , n7863 , n7865 );
and ( n7867 , n7666 , n7866 );
xor ( n7868 , n6442 , n7267 );
buf ( n7869 , n7868 );
buf ( n7870 , n7869 );
buf ( n7871 , n7870 );
and ( n7872 , n7871 , n7864 );
nor ( n7873 , n7867 , n7872 );
and ( n7874 , n7862 , n7734 );
not ( n7875 , n7874 );
and ( n7876 , n7658 , n7875 );
xnor ( n7877 , n7873 , n7876 );
xor ( n7878 , n7857 , n7877 );
and ( n7879 , n7814 , n7878 );
and ( n7880 , n7792 , n7878 );
or ( n7881 , n7815 , n7879 , n7880 );
xor ( n7882 , n3673 , n7290 );
buf ( n7883 , n7882 );
buf ( n7884 , n7883 );
buf ( n7885 , n7884 );
xor ( n7886 , n7441 , n7442 );
xor ( n7887 , n7886 , n7453 );
buf ( n7888 , n7887 );
buf ( n7889 , n7888 );
buf ( n7890 , n7889 );
xor ( n7891 , n7444 , n7445 );
xor ( n7892 , n7891 , n7450 );
buf ( n7893 , n7892 );
buf ( n7894 , n7893 );
buf ( n7895 , n7894 );
xor ( n7896 , n7890 , n7895 );
xor ( n7897 , n7895 , n7381 );
not ( n7898 , n7897 );
and ( n7899 , n7896 , n7898 );
and ( n7900 , n7885 , n7899 );
xor ( n7901 , n3671 , n7291 );
buf ( n7902 , n7901 );
buf ( n7903 , n7902 );
buf ( n7904 , n7903 );
and ( n7905 , n7904 , n7897 );
nor ( n7906 , n7900 , n7905 );
and ( n7907 , n7895 , n7381 );
not ( n7908 , n7907 );
and ( n7909 , n7890 , n7908 );
xnor ( n7910 , n7906 , n7909 );
and ( n7911 , n7881 , n7910 );
and ( n7912 , n7843 , n7856 );
and ( n7913 , n7856 , n7877 );
and ( n7914 , n7843 , n7877 );
or ( n7915 , n7912 , n7913 , n7914 );
xor ( n7916 , n3685 , n7284 );
buf ( n7917 , n7916 );
buf ( n7918 , n7917 );
buf ( n7919 , n7918 );
xor ( n7920 , n7423 , n7424 );
xor ( n7921 , n7920 , n7471 );
buf ( n7922 , n7921 );
buf ( n7923 , n7922 );
buf ( n7924 , n7923 );
xor ( n7925 , n7426 , n7427 );
xor ( n7926 , n7925 , n7468 );
buf ( n7927 , n7926 );
buf ( n7928 , n7927 );
buf ( n7929 , n7928 );
xor ( n7930 , n7924 , n7929 );
xor ( n7931 , n7929 , n7767 );
not ( n7932 , n7931 );
and ( n7933 , n7930 , n7932 );
and ( n7934 , n7919 , n7933 );
and ( n7935 , n7762 , n7931 );
nor ( n7936 , n7934 , n7935 );
and ( n7937 , n7929 , n7767 );
not ( n7938 , n7937 );
and ( n7939 , n7924 , n7938 );
xnor ( n7940 , n7936 , n7939 );
xor ( n7941 , n7915 , n7940 );
xor ( n7942 , n3689 , n7282 );
buf ( n7943 , n7942 );
buf ( n7944 , n7943 );
buf ( n7945 , n7944 );
xor ( n7946 , n7420 , n7421 );
xor ( n7947 , n7946 , n7474 );
buf ( n7948 , n7947 );
buf ( n7949 , n7948 );
buf ( n7950 , n7949 );
xor ( n7951 , n7498 , n7950 );
xor ( n7952 , n7950 , n7924 );
not ( n7953 , n7952 );
and ( n7954 , n7951 , n7953 );
and ( n7955 , n7945 , n7954 );
xor ( n7956 , n3687 , n7283 );
buf ( n7957 , n7956 );
buf ( n7958 , n7957 );
buf ( n7959 , n7958 );
and ( n7960 , n7959 , n7952 );
nor ( n7961 , n7955 , n7960 );
and ( n7962 , n7950 , n7924 );
not ( n7963 , n7962 );
and ( n7964 , n7498 , n7963 );
xnor ( n7965 , n7961 , n7964 );
xor ( n7966 , n7941 , n7965 );
and ( n7967 , n7910 , n7966 );
and ( n7968 , n7881 , n7966 );
or ( n7969 , n7911 , n7967 , n7968 );
xor ( n7970 , n7758 , n7969 );
and ( n7971 , n7915 , n7940 );
and ( n7972 , n7940 , n7965 );
and ( n7973 , n7915 , n7965 );
or ( n7974 , n7971 , n7972 , n7973 );
and ( n7975 , n7904 , n7899 );
and ( n7976 , n7352 , n7897 );
nor ( n7977 , n7975 , n7976 );
xnor ( n7978 , n7977 , n7909 );
xor ( n7979 , n7974 , n7978 );
and ( n7980 , n7666 , n7661 );
and ( n7981 , n7871 , n7659 );
nor ( n7982 , n7980 , n7981 );
xnor ( n7983 , n7982 , n7671 );
and ( n7984 , n7696 , n7691 );
and ( n7985 , n7828 , n7689 );
nor ( n7986 , n7984 , n7985 );
not ( n7987 , n7986 );
xor ( n7988 , n7983 , n7987 );
and ( n7989 , n7672 , n7699 );
xor ( n7990 , n7988 , n7989 );
and ( n7991 , n7718 , n7713 );
and ( n7992 , n7516 , n7711 );
nor ( n7993 , n7991 , n7992 );
xnor ( n7994 , n7993 , n7723 );
xor ( n7995 , n7990 , n7994 );
xor ( n7996 , n7979 , n7995 );
xor ( n7997 , n7970 , n7996 );
xor ( n7998 , n7348 , n7997 );
and ( n7999 , n7704 , n7542 );
and ( n8000 , n7718 , n7540 );
nor ( n8001 , n7999 , n8000 );
xnor ( n8002 , n8001 , n7552 );
and ( n8003 , n7871 , n7743 );
and ( n8004 , n7800 , n7741 );
nor ( n8005 , n8003 , n8004 );
xnor ( n8006 , n8005 , n7753 );
and ( n8007 , n8002 , n8006 );
and ( n8008 , n7828 , n7661 );
and ( n8009 , n7809 , n7659 );
nor ( n8010 , n8008 , n8009 );
xnor ( n8011 , n8010 , n7671 );
and ( n8012 , n8006 , n8011 );
and ( n8013 , n8002 , n8011 );
or ( n8014 , n8007 , n8012 , n8013 );
and ( n8015 , n7516 , n7501 );
and ( n8016 , n7547 , n7499 );
nor ( n8017 , n8015 , n8016 );
xnor ( n8018 , n8017 , n7511 );
and ( n8019 , n7558 , n7713 );
and ( n8020 , n7606 , n7711 );
nor ( n8021 , n8019 , n8020 );
xnor ( n8022 , n8021 , n7723 );
and ( n8023 , n8018 , n8022 );
and ( n8024 , n7729 , n7601 );
and ( n8025 , n7748 , n7599 );
nor ( n8026 , n8024 , n8025 );
xnor ( n8027 , n8026 , n7611 );
and ( n8028 , n8022 , n8027 );
and ( n8029 , n8018 , n8027 );
or ( n8030 , n8023 , n8028 , n8029 );
and ( n8031 , n8014 , n8030 );
xor ( n8032 , n3679 , n7287 );
buf ( n8033 , n8032 );
buf ( n8034 , n8033 );
buf ( n8035 , n8034 );
xor ( n8036 , n7438 , n7439 );
xor ( n8037 , n8036 , n7456 );
buf ( n8038 , n8037 );
buf ( n8039 , n8038 );
buf ( n8040 , n8039 );
xor ( n8041 , n7778 , n8040 );
xor ( n8042 , n8040 , n7890 );
not ( n8043 , n8042 );
and ( n8044 , n8041 , n8043 );
and ( n8045 , n8035 , n8044 );
xor ( n8046 , n3677 , n7288 );
buf ( n8047 , n8046 );
buf ( n8048 , n8047 );
buf ( n8049 , n8048 );
and ( n8050 , n8049 , n8042 );
nor ( n8051 , n8045 , n8050 );
and ( n8052 , n8040 , n7890 );
not ( n8053 , n8052 );
and ( n8054 , n7778 , n8053 );
xnor ( n8055 , n8051 , n8054 );
and ( n8056 , n8030 , n8055 );
and ( n8057 , n8014 , n8055 );
or ( n8058 , n8031 , n8056 , n8057 );
and ( n8059 , n7838 , n7823 );
and ( n8060 , n7676 , n7821 );
nor ( n8061 , n8059 , n8060 );
xnor ( n8062 , n8061 , n7833 );
xor ( n8063 , n6460 , n7258 );
buf ( n8064 , n8063 );
buf ( n8065 , n8064 );
buf ( n8066 , n8065 );
and ( n8067 , n8066 , n7691 );
and ( n8068 , n7851 , n7689 );
nor ( n8069 , n8067 , n8068 );
not ( n8070 , n8069 );
xor ( n8071 , n8062 , n8070 );
and ( n8072 , n7676 , n7661 );
and ( n8073 , n7696 , n7659 );
nor ( n8074 , n8072 , n8073 );
xnor ( n8075 , n8074 , n7671 );
xor ( n8076 , n6462 , n7257 );
buf ( n8077 , n8076 );
buf ( n8078 , n8077 );
buf ( n8079 , n8078 );
and ( n8080 , n8079 , n7691 );
and ( n8081 , n8066 , n7689 );
nor ( n8082 , n8080 , n8081 );
not ( n8083 , n8082 );
and ( n8084 , n8075 , n8083 );
and ( n8085 , n8071 , n8084 );
and ( n8086 , n7696 , n7661 );
and ( n8087 , n7828 , n7659 );
nor ( n8088 , n8086 , n8087 );
xnor ( n8089 , n8088 , n7671 );
and ( n8090 , n8084 , n8089 );
and ( n8091 , n8071 , n8089 );
or ( n8092 , n8085 , n8090 , n8091 );
and ( n8093 , n7919 , n7781 );
and ( n8094 , n7762 , n7779 );
nor ( n8095 , n8093 , n8094 );
xnor ( n8096 , n8095 , n7791 );
and ( n8097 , n8092 , n8096 );
and ( n8098 , n7410 , n7954 );
and ( n8099 , n7506 , n7952 );
nor ( n8100 , n8098 , n8099 );
xnor ( n8101 , n8100 , n7964 );
and ( n8102 , n8096 , n8101 );
and ( n8103 , n8092 , n8101 );
or ( n8104 , n8097 , n8102 , n8103 );
xor ( n8105 , n3675 , n7289 );
buf ( n8106 , n8105 );
buf ( n8107 , n8106 );
buf ( n8108 , n8107 );
and ( n8109 , n8108 , n7899 );
and ( n8110 , n7885 , n7897 );
nor ( n8111 , n8109 , n8110 );
xnor ( n8112 , n8111 , n7909 );
and ( n8113 , n8104 , n8112 );
and ( n8114 , n7718 , n7542 );
and ( n8115 , n7516 , n7540 );
nor ( n8116 , n8114 , n8115 );
xnor ( n8117 , n8116 , n7552 );
and ( n8118 , n7606 , n7713 );
and ( n8119 , n7704 , n7711 );
nor ( n8120 , n8118 , n8119 );
xnor ( n8121 , n8120 , n7723 );
xor ( n8122 , n8117 , n8121 );
and ( n8123 , n7748 , n7601 );
and ( n8124 , n7558 , n7599 );
nor ( n8125 , n8123 , n8124 );
xnor ( n8126 , n8125 , n7611 );
xor ( n8127 , n8122 , n8126 );
and ( n8128 , n8112 , n8127 );
and ( n8129 , n8104 , n8127 );
or ( n8130 , n8113 , n8128 , n8129 );
and ( n8131 , n8058 , n8130 );
and ( n8132 , n8117 , n8121 );
and ( n8133 , n8121 , n8126 );
and ( n8134 , n8117 , n8126 );
or ( n8135 , n8132 , n8133 , n8134 );
and ( n8136 , n7796 , n7804 );
and ( n8137 , n7804 , n7813 );
and ( n8138 , n7796 , n7813 );
or ( n8139 , n8136 , n8137 , n8138 );
xor ( n8140 , n8135 , n8139 );
and ( n8141 , n7834 , n7842 );
and ( n8142 , n7871 , n7866 );
and ( n8143 , n7800 , n7864 );
nor ( n8144 , n8142 , n8143 );
xnor ( n8145 , n8144 , n7876 );
xor ( n8146 , n8141 , n8145 );
and ( n8147 , n7828 , n7823 );
and ( n8148 , n7809 , n7821 );
nor ( n8149 , n8147 , n8148 );
xnor ( n8150 , n8149 , n7833 );
xor ( n8151 , n8146 , n8150 );
xor ( n8152 , n8140 , n8151 );
and ( n8153 , n8130 , n8152 );
and ( n8154 , n8058 , n8152 );
or ( n8155 , n8131 , n8153 , n8154 );
xor ( n8156 , n3663 , n7295 );
buf ( n8157 , n8156 );
buf ( n8158 , n8157 );
buf ( n8159 , n8158 );
xor ( n8160 , n7362 , n7363 );
xor ( n8161 , n8160 , n7368 );
buf ( n8162 , n8161 );
buf ( n8163 , n8162 );
buf ( n8164 , n8163 );
xor ( n8165 , n7392 , n8164 );
xor ( n8166 , n8164 , n7311 );
not ( n8167 , n8166 );
and ( n8168 , n8165 , n8167 );
and ( n8169 , n8159 , n8168 );
xor ( n8170 , n3661 , n7296 );
buf ( n8171 , n8170 );
buf ( n8172 , n8171 );
buf ( n8173 , n8172 );
and ( n8174 , n8173 , n8166 );
nor ( n8175 , n8169 , n8174 );
and ( n8176 , n8164 , n7311 );
not ( n8177 , n8176 );
and ( n8178 , n7392 , n8177 );
xnor ( n8179 , n8175 , n8178 );
xor ( n8180 , n8155 , n8179 );
and ( n8181 , n8135 , n8139 );
and ( n8182 , n8139 , n8151 );
and ( n8183 , n8135 , n8151 );
or ( n8184 , n8181 , n8182 , n8183 );
and ( n8185 , n8141 , n8145 );
and ( n8186 , n8145 , n8150 );
and ( n8187 , n8141 , n8150 );
or ( n8188 , n8185 , n8186 , n8187 );
and ( n8189 , n7762 , n7933 );
and ( n8190 , n7786 , n7931 );
nor ( n8191 , n8189 , n8190 );
xnor ( n8192 , n8191 , n7939 );
xor ( n8193 , n8188 , n8192 );
and ( n8194 , n7506 , n7501 );
and ( n8195 , n7945 , n7499 );
nor ( n8196 , n8194 , n8195 );
xnor ( n8197 , n8196 , n7511 );
xor ( n8198 , n8193 , n8197 );
xor ( n8199 , n8184 , n8198 );
and ( n8200 , n7700 , n7724 );
and ( n8201 , n7724 , n7754 );
and ( n8202 , n7700 , n7754 );
or ( n8203 , n8200 , n8201 , n8202 );
and ( n8204 , n8108 , n8044 );
and ( n8205 , n7885 , n8042 );
nor ( n8206 , n8204 , n8205 );
xnor ( n8207 , n8206 , n8054 );
xor ( n8208 , n8203 , n8207 );
and ( n8209 , n7547 , n7542 );
and ( n8210 , n7410 , n7540 );
nor ( n8211 , n8209 , n8210 );
xnor ( n8212 , n8211 , n7552 );
and ( n8213 , n7800 , n7866 );
and ( n8214 , n7729 , n7864 );
nor ( n8215 , n8213 , n8214 );
xnor ( n8216 , n8215 , n7876 );
xor ( n8217 , n8212 , n8216 );
and ( n8218 , n7809 , n7823 );
and ( n8219 , n7618 , n7821 );
nor ( n8220 , n8218 , n8219 );
xnor ( n8221 , n8220 , n7833 );
xor ( n8222 , n8217 , n8221 );
xor ( n8223 , n8208 , n8222 );
xor ( n8224 , n8199 , n8223 );
xor ( n8225 , n8180 , n8224 );
xor ( n8226 , n7998 , n8225 );
and ( n8227 , n7547 , n7954 );
and ( n8228 , n7410 , n7952 );
nor ( n8229 , n8227 , n8228 );
xnor ( n8230 , n8229 , n7964 );
and ( n8231 , n7718 , n7501 );
and ( n8232 , n7516 , n7499 );
nor ( n8233 , n8231 , n8232 );
xnor ( n8234 , n8233 , n7511 );
and ( n8235 , n8230 , n8234 );
and ( n8236 , n7606 , n7542 );
and ( n8237 , n7704 , n7540 );
nor ( n8238 , n8236 , n8237 );
xnor ( n8239 , n8238 , n7552 );
and ( n8240 , n8234 , n8239 );
and ( n8241 , n8230 , n8239 );
or ( n8242 , n8235 , n8240 , n8241 );
and ( n8243 , n8049 , n7899 );
and ( n8244 , n8108 , n7897 );
nor ( n8245 , n8243 , n8244 );
xnor ( n8246 , n8245 , n7909 );
and ( n8247 , n8242 , n8246 );
and ( n8248 , n7786 , n8044 );
and ( n8249 , n8035 , n8042 );
nor ( n8250 , n8248 , n8249 );
xnor ( n8251 , n8250 , n8054 );
and ( n8252 , n8246 , n8251 );
and ( n8253 , n8242 , n8251 );
or ( n8254 , n8247 , n8252 , n8253 );
xor ( n8255 , n8075 , n8083 );
and ( n8256 , n8066 , n7823 );
and ( n8257 , n7851 , n7821 );
nor ( n8258 , n8256 , n8257 );
xnor ( n8259 , n8258 , n7833 );
xor ( n8260 , n6464 , n7256 );
buf ( n8261 , n8260 );
buf ( n8262 , n8261 );
buf ( n8263 , n8262 );
and ( n8264 , n8263 , n7691 );
and ( n8265 , n8079 , n7689 );
nor ( n8266 , n8264 , n8265 );
not ( n8267 , n8266 );
and ( n8268 , n8259 , n8267 );
and ( n8269 , n8255 , n8268 );
and ( n8270 , n7851 , n7823 );
and ( n8271 , n7838 , n7821 );
nor ( n8272 , n8270 , n8271 );
xnor ( n8273 , n8272 , n7833 );
and ( n8274 , n8268 , n8273 );
and ( n8275 , n8255 , n8273 );
or ( n8276 , n8269 , n8274 , n8275 );
and ( n8277 , n7959 , n7781 );
and ( n8278 , n7919 , n7779 );
nor ( n8279 , n8277 , n8278 );
xnor ( n8280 , n8279 , n7791 );
and ( n8281 , n8276 , n8280 );
and ( n8282 , n7748 , n7713 );
and ( n8283 , n7558 , n7711 );
nor ( n8284 , n8282 , n8283 );
xnor ( n8285 , n8284 , n7723 );
and ( n8286 , n8280 , n8285 );
and ( n8287 , n8276 , n8285 );
or ( n8288 , n8281 , n8286 , n8287 );
xor ( n8289 , n8002 , n8006 );
xor ( n8290 , n8289 , n8011 );
and ( n8291 , n8288 , n8290 );
xor ( n8292 , n8018 , n8022 );
xor ( n8293 , n8292 , n8027 );
and ( n8294 , n8290 , n8293 );
and ( n8295 , n8288 , n8293 );
or ( n8296 , n8291 , n8294 , n8295 );
and ( n8297 , n8254 , n8296 );
xor ( n8298 , n7792 , n7814 );
xor ( n8299 , n8298 , n7878 );
and ( n8300 , n8296 , n8299 );
and ( n8301 , n8254 , n8299 );
or ( n8302 , n8297 , n8300 , n8301 );
xor ( n8303 , n3665 , n7294 );
buf ( n8304 , n8303 );
buf ( n8305 , n8304 );
buf ( n8306 , n8305 );
and ( n8307 , n8306 , n8168 );
and ( n8308 , n8159 , n8166 );
nor ( n8309 , n8307 , n8308 );
xnor ( n8310 , n8309 , n8178 );
xor ( n8311 , n8302 , n8310 );
xor ( n8312 , n7881 , n7910 );
xor ( n8313 , n8312 , n7966 );
xor ( n8314 , n8311 , n8313 );
and ( n8315 , n7352 , n8168 );
and ( n8316 , n7400 , n8166 );
nor ( n8317 , n8315 , n8316 );
xnor ( n8318 , n8317 , n8178 );
and ( n8319 , n7885 , n7395 );
and ( n8320 , n7904 , n7393 );
nor ( n8321 , n8319 , n8320 );
xnor ( n8322 , n8321 , n7405 );
and ( n8323 , n8318 , n8322 );
xor ( n8324 , n8092 , n8096 );
xor ( n8325 , n8324 , n8101 );
and ( n8326 , n8322 , n8325 );
and ( n8327 , n8318 , n8325 );
or ( n8328 , n8323 , n8326 , n8327 );
and ( n8329 , n7400 , n8168 );
and ( n8330 , n8306 , n8166 );
nor ( n8331 , n8329 , n8330 );
xnor ( n8332 , n8331 , n8178 );
and ( n8333 , n8328 , n8332 );
xor ( n8334 , n8014 , n8030 );
xor ( n8335 , n8334 , n8055 );
and ( n8336 , n8332 , n8335 );
and ( n8337 , n8328 , n8335 );
or ( n8338 , n8333 , n8336 , n8337 );
xor ( n8339 , n8058 , n8130 );
xor ( n8340 , n8339 , n8152 );
xor ( n8341 , n8338 , n8340 );
and ( n8342 , n7800 , n7601 );
and ( n8343 , n7729 , n7599 );
nor ( n8344 , n8342 , n8343 );
xnor ( n8345 , n8344 , n7611 );
and ( n8346 , n7666 , n7743 );
and ( n8347 , n7871 , n7741 );
nor ( n8348 , n8346 , n8347 );
xnor ( n8349 , n8348 , n7753 );
and ( n8350 , n8345 , n8349 );
and ( n8351 , n7809 , n7866 );
and ( n8352 , n7618 , n7864 );
nor ( n8353 , n8351 , n8352 );
xnor ( n8354 , n8353 , n7876 );
and ( n8355 , n8349 , n8354 );
and ( n8356 , n8345 , n8354 );
or ( n8357 , n8350 , n8355 , n8356 );
and ( n8358 , n7945 , n7933 );
and ( n8359 , n7959 , n7931 );
nor ( n8360 , n8358 , n8359 );
xnor ( n8361 , n8360 , n7939 );
and ( n8362 , n8357 , n8361 );
xor ( n8363 , n7847 , n7855 );
and ( n8364 , n8062 , n8070 );
xor ( n8365 , n8363 , n8364 );
and ( n8366 , n7618 , n7866 );
and ( n8367 , n7666 , n7864 );
nor ( n8368 , n8366 , n8367 );
xnor ( n8369 , n8368 , n7876 );
xor ( n8370 , n8365 , n8369 );
and ( n8371 , n8361 , n8370 );
and ( n8372 , n8357 , n8370 );
or ( n8373 , n8362 , n8371 , n8372 );
and ( n8374 , n7904 , n7395 );
and ( n8375 , n7352 , n7393 );
nor ( n8376 , n8374 , n8375 );
xnor ( n8377 , n8376 , n7405 );
and ( n8378 , n8373 , n8377 );
and ( n8379 , n8363 , n8364 );
and ( n8380 , n8364 , n8369 );
and ( n8381 , n8363 , n8369 );
or ( n8382 , n8379 , n8380 , n8381 );
and ( n8383 , n7959 , n7933 );
and ( n8384 , n7919 , n7931 );
nor ( n8385 , n8383 , n8384 );
xnor ( n8386 , n8385 , n7939 );
xor ( n8387 , n8382 , n8386 );
and ( n8388 , n7506 , n7954 );
and ( n8389 , n7945 , n7952 );
nor ( n8390 , n8388 , n8389 );
xnor ( n8391 , n8390 , n7964 );
xor ( n8392 , n8387 , n8391 );
and ( n8393 , n8377 , n8392 );
and ( n8394 , n8373 , n8392 );
or ( n8395 , n8378 , n8393 , n8394 );
and ( n8396 , n8382 , n8386 );
and ( n8397 , n8386 , n8391 );
and ( n8398 , n8382 , n8391 );
or ( n8399 , n8396 , n8397 , n8398 );
and ( n8400 , n8049 , n8044 );
and ( n8401 , n8108 , n8042 );
nor ( n8402 , n8400 , n8401 );
xnor ( n8403 , n8402 , n8054 );
xor ( n8404 , n8399 , n8403 );
and ( n8405 , n7786 , n7781 );
and ( n8406 , n8035 , n7779 );
nor ( n8407 , n8405 , n8406 );
xnor ( n8408 , n8407 , n7791 );
xor ( n8409 , n8404 , n8408 );
xor ( n8410 , n8395 , n8409 );
xor ( n8411 , n7406 , n7613 );
xor ( n8412 , n8411 , n7755 );
xor ( n8413 , n8410 , n8412 );
xor ( n8414 , n8341 , n8413 );
and ( n8415 , n8314 , n8414 );
and ( n8416 , n8226 , n8415 );
and ( n8417 , n8173 , n7318 );
and ( n8418 , n7301 , n7315 );
nor ( n8419 , n8417 , n8418 );
xnor ( n8420 , n8419 , n7311 );
xor ( n8421 , n8259 , n8267 );
and ( n8422 , n8079 , n7823 );
and ( n8423 , n8066 , n7821 );
nor ( n8424 , n8422 , n8423 );
xnor ( n8425 , n8424 , n7833 );
xor ( n8426 , n6466 , n7255 );
buf ( n8427 , n8426 );
buf ( n8428 , n8427 );
buf ( n8429 , n8428 );
and ( n8430 , n8429 , n7691 );
and ( n8431 , n8263 , n7689 );
nor ( n8432 , n8430 , n8431 );
not ( n8433 , n8432 );
and ( n8434 , n8425 , n8433 );
and ( n8435 , n8421 , n8434 );
and ( n8436 , n7838 , n7661 );
and ( n8437 , n7676 , n7659 );
nor ( n8438 , n8436 , n8437 );
xnor ( n8439 , n8438 , n7671 );
and ( n8440 , n8434 , n8439 );
and ( n8441 , n8421 , n8439 );
or ( n8442 , n8435 , n8440 , n8441 );
and ( n8443 , n7871 , n7601 );
and ( n8444 , n7800 , n7599 );
nor ( n8445 , n8443 , n8444 );
xnor ( n8446 , n8445 , n7611 );
and ( n8447 , n8442 , n8446 );
and ( n8448 , n7618 , n7743 );
and ( n8449 , n7666 , n7741 );
nor ( n8450 , n8448 , n8449 );
xnor ( n8451 , n8450 , n7753 );
and ( n8452 , n8446 , n8451 );
and ( n8453 , n8442 , n8451 );
or ( n8454 , n8447 , n8452 , n8453 );
and ( n8455 , n7762 , n8044 );
and ( n8456 , n7786 , n8042 );
nor ( n8457 , n8455 , n8456 );
xnor ( n8458 , n8457 , n8054 );
and ( n8459 , n8454 , n8458 );
and ( n8460 , n7506 , n7933 );
and ( n8461 , n7945 , n7931 );
nor ( n8462 , n8460 , n8461 );
xnor ( n8463 , n8462 , n7939 );
and ( n8464 , n8458 , n8463 );
and ( n8465 , n8454 , n8463 );
or ( n8466 , n8459 , n8464 , n8465 );
and ( n8467 , n8108 , n7395 );
and ( n8468 , n7885 , n7393 );
nor ( n8469 , n8467 , n8468 );
xnor ( n8470 , n8469 , n7405 );
and ( n8471 , n8035 , n7899 );
and ( n8472 , n8049 , n7897 );
nor ( n8473 , n8471 , n8472 );
xnor ( n8474 , n8473 , n7909 );
and ( n8475 , n8470 , n8474 );
xor ( n8476 , n8071 , n8084 );
xor ( n8477 , n8476 , n8089 );
and ( n8478 , n8474 , n8477 );
and ( n8479 , n8470 , n8477 );
or ( n8480 , n8475 , n8478 , n8479 );
and ( n8481 , n8466 , n8480 );
xor ( n8482 , n8357 , n8361 );
xor ( n8483 , n8482 , n8370 );
and ( n8484 , n8480 , n8483 );
and ( n8485 , n8466 , n8483 );
or ( n8486 , n8481 , n8484 , n8485 );
xor ( n8487 , n8104 , n8112 );
xor ( n8488 , n8487 , n8127 );
and ( n8489 , n8486 , n8488 );
xor ( n8490 , n8373 , n8377 );
xor ( n8491 , n8490 , n8392 );
and ( n8492 , n8488 , n8491 );
and ( n8493 , n8486 , n8491 );
or ( n8494 , n8489 , n8492 , n8493 );
and ( n8495 , n8420 , n8494 );
and ( n8496 , n8159 , n7318 );
and ( n8497 , n8173 , n7315 );
nor ( n8498 , n8496 , n8497 );
xnor ( n8499 , n8498 , n7311 );
xor ( n8500 , n8254 , n8296 );
xor ( n8501 , n8500 , n8299 );
and ( n8502 , n8499 , n8501 );
and ( n8503 , n7704 , n7501 );
and ( n8504 , n7718 , n7499 );
nor ( n8505 , n8503 , n8504 );
xnor ( n8506 , n8505 , n7511 );
and ( n8507 , n7558 , n7542 );
and ( n8508 , n7606 , n7540 );
nor ( n8509 , n8507 , n8508 );
xnor ( n8510 , n8509 , n7552 );
and ( n8511 , n8506 , n8510 );
and ( n8512 , n7828 , n7866 );
and ( n8513 , n7809 , n7864 );
nor ( n8514 , n8512 , n8513 );
xnor ( n8515 , n8514 , n7876 );
and ( n8516 , n8510 , n8515 );
and ( n8517 , n8506 , n8515 );
or ( n8518 , n8511 , n8516 , n8517 );
and ( n8519 , n7945 , n7781 );
and ( n8520 , n7959 , n7779 );
nor ( n8521 , n8519 , n8520 );
xnor ( n8522 , n8521 , n7791 );
and ( n8523 , n7410 , n7933 );
and ( n8524 , n7506 , n7931 );
nor ( n8525 , n8523 , n8524 );
xnor ( n8526 , n8525 , n7939 );
and ( n8527 , n8522 , n8526 );
xor ( n8528 , n8255 , n8268 );
xor ( n8529 , n8528 , n8273 );
and ( n8530 , n8526 , n8529 );
and ( n8531 , n8522 , n8529 );
or ( n8532 , n8527 , n8530 , n8531 );
and ( n8533 , n8518 , n8532 );
xor ( n8534 , n8345 , n8349 );
xor ( n8535 , n8534 , n8354 );
and ( n8536 , n8532 , n8535 );
and ( n8537 , n8518 , n8535 );
or ( n8538 , n8533 , n8536 , n8537 );
and ( n8539 , n7919 , n8044 );
and ( n8540 , n7762 , n8042 );
nor ( n8541 , n8539 , n8540 );
xnor ( n8542 , n8541 , n8054 );
and ( n8543 , n7516 , n7954 );
and ( n8544 , n7547 , n7952 );
nor ( n8545 , n8543 , n8544 );
xnor ( n8546 , n8545 , n7964 );
and ( n8547 , n8542 , n8546 );
and ( n8548 , n7729 , n7713 );
and ( n8549 , n7748 , n7711 );
nor ( n8550 , n8548 , n8549 );
xnor ( n8551 , n8550 , n7723 );
and ( n8552 , n8546 , n8551 );
and ( n8553 , n8542 , n8551 );
or ( n8554 , n8547 , n8552 , n8553 );
xor ( n8555 , n8230 , n8234 );
xor ( n8556 , n8555 , n8239 );
and ( n8557 , n8554 , n8556 );
xor ( n8558 , n8276 , n8280 );
xor ( n8559 , n8558 , n8285 );
and ( n8560 , n8556 , n8559 );
and ( n8561 , n8554 , n8559 );
or ( n8562 , n8557 , n8560 , n8561 );
and ( n8563 , n8538 , n8562 );
xor ( n8564 , n8242 , n8246 );
xor ( n8565 , n8564 , n8251 );
and ( n8566 , n8562 , n8565 );
and ( n8567 , n8538 , n8565 );
or ( n8568 , n8563 , n8566 , n8567 );
and ( n8569 , n8501 , n8568 );
and ( n8570 , n8499 , n8568 );
or ( n8571 , n8502 , n8569 , n8570 );
and ( n8572 , n8494 , n8571 );
and ( n8573 , n8420 , n8571 );
or ( n8574 , n8495 , n8572 , n8573 );
and ( n8575 , n8415 , n8574 );
and ( n8576 , n8226 , n8574 );
or ( n8577 , n8416 , n8575 , n8576 );
and ( n8578 , n8338 , n8340 );
and ( n8579 , n8340 , n8413 );
and ( n8580 , n8338 , n8413 );
or ( n8581 , n8578 , n8579 , n8580 );
and ( n8582 , n8395 , n8409 );
and ( n8583 , n8409 , n8412 );
and ( n8584 , n8395 , n8412 );
or ( n8585 , n8582 , n8583 , n8584 );
and ( n8586 , n8302 , n8310 );
and ( n8587 , n8310 , n8313 );
and ( n8588 , n8302 , n8313 );
or ( n8589 , n8586 , n8587 , n8588 );
xor ( n8590 , n8585 , n8589 );
and ( n8591 , n8399 , n8403 );
and ( n8592 , n8403 , n8408 );
and ( n8593 , n8399 , n8408 );
or ( n8594 , n8591 , n8592 , n8593 );
and ( n8595 , n7400 , n7395 );
and ( n8596 , n8306 , n7393 );
nor ( n8597 , n8595 , n8596 );
xnor ( n8598 , n8597 , n7405 );
xor ( n8599 , n8594 , n8598 );
and ( n8600 , n7512 , n7553 );
and ( n8601 , n7553 , n7612 );
and ( n8602 , n7512 , n7612 );
or ( n8603 , n8600 , n8601 , n8602 );
and ( n8604 , n8035 , n7781 );
and ( n8605 , n8049 , n7779 );
nor ( n8606 , n8604 , n8605 );
xnor ( n8607 , n8606 , n7791 );
xor ( n8608 , n8603 , n8607 );
and ( n8609 , n7959 , n7954 );
and ( n8610 , n7919 , n7952 );
nor ( n8611 , n8609 , n8610 );
xnor ( n8612 , n8611 , n7964 );
and ( n8613 , n7606 , n7601 );
and ( n8614 , n7704 , n7599 );
nor ( n8615 , n8613 , n8614 );
xnor ( n8616 , n8615 , n7611 );
xor ( n8617 , n8612 , n8616 );
and ( n8618 , n7748 , n7743 );
and ( n8619 , n7558 , n7741 );
nor ( n8620 , n8618 , n8619 );
xnor ( n8621 , n8620 , n7753 );
xor ( n8622 , n8617 , n8621 );
xor ( n8623 , n8608 , n8622 );
xor ( n8624 , n8599 , n8623 );
xor ( n8625 , n8590 , n8624 );
xor ( n8626 , n8581 , n8625 );
xor ( n8627 , n8314 , n8414 );
and ( n8628 , n8306 , n7318 );
and ( n8629 , n8159 , n7315 );
nor ( n8630 , n8628 , n8629 );
xnor ( n8631 , n8630 , n7311 );
xor ( n8632 , n8288 , n8290 );
xor ( n8633 , n8632 , n8293 );
and ( n8634 , n8631 , n8633 );
xor ( n8635 , n8318 , n8322 );
xor ( n8636 , n8635 , n8325 );
and ( n8637 , n8633 , n8636 );
and ( n8638 , n8631 , n8636 );
or ( n8639 , n8634 , n8637 , n8638 );
and ( n8640 , n7959 , n8044 );
and ( n8641 , n7919 , n8042 );
nor ( n8642 , n8640 , n8641 );
xnor ( n8643 , n8642 , n8054 );
and ( n8644 , n7800 , n7713 );
and ( n8645 , n7729 , n7711 );
nor ( n8646 , n8644 , n8645 );
xnor ( n8647 , n8646 , n7723 );
and ( n8648 , n8643 , n8647 );
and ( n8649 , n7809 , n7743 );
and ( n8650 , n7618 , n7741 );
nor ( n8651 , n8649 , n8650 );
xnor ( n8652 , n8651 , n7753 );
and ( n8653 , n8647 , n8652 );
and ( n8654 , n8643 , n8652 );
or ( n8655 , n8648 , n8653 , n8654 );
and ( n8656 , n7718 , n7954 );
and ( n8657 , n7516 , n7952 );
nor ( n8658 , n8656 , n8657 );
xnor ( n8659 , n8658 , n7964 );
and ( n8660 , n7606 , n7501 );
and ( n8661 , n7704 , n7499 );
nor ( n8662 , n8660 , n8661 );
xnor ( n8663 , n8662 , n7511 );
and ( n8664 , n8659 , n8663 );
and ( n8665 , n7748 , n7542 );
and ( n8666 , n7558 , n7540 );
nor ( n8667 , n8665 , n8666 );
xnor ( n8668 , n8667 , n7552 );
and ( n8669 , n8663 , n8668 );
and ( n8670 , n8659 , n8668 );
or ( n8671 , n8664 , n8669 , n8670 );
and ( n8672 , n8655 , n8671 );
xor ( n8673 , n8442 , n8446 );
xor ( n8674 , n8673 , n8451 );
and ( n8675 , n8671 , n8674 );
and ( n8676 , n8655 , n8674 );
or ( n8677 , n8672 , n8675 , n8676 );
and ( n8678 , n7904 , n8168 );
and ( n8679 , n7352 , n8166 );
nor ( n8680 , n8678 , n8679 );
xnor ( n8681 , n8680 , n8178 );
and ( n8682 , n8677 , n8681 );
xor ( n8683 , n8454 , n8458 );
xor ( n8684 , n8683 , n8463 );
and ( n8685 , n8681 , n8684 );
and ( n8686 , n8677 , n8684 );
or ( n8687 , n8682 , n8685 , n8686 );
xor ( n8688 , n8425 , n8433 );
and ( n8689 , n8066 , n7661 );
and ( n8690 , n7851 , n7659 );
nor ( n8691 , n8689 , n8690 );
xnor ( n8692 , n8691 , n7671 );
xor ( n8693 , n6468 , n7254 );
buf ( n8694 , n8693 );
buf ( n8695 , n8694 );
buf ( n8696 , n8695 );
and ( n8697 , n8696 , n7691 );
and ( n8698 , n8429 , n7689 );
nor ( n8699 , n8697 , n8698 );
not ( n8700 , n8699 );
and ( n8701 , n8692 , n8700 );
and ( n8702 , n8688 , n8701 );
and ( n8703 , n7676 , n7866 );
and ( n8704 , n7696 , n7864 );
nor ( n8705 , n8703 , n8704 );
xnor ( n8706 , n8705 , n7876 );
and ( n8707 , n8701 , n8706 );
and ( n8708 , n8688 , n8706 );
or ( n8709 , n8702 , n8707 , n8708 );
and ( n8710 , n7666 , n7601 );
and ( n8711 , n7871 , n7599 );
nor ( n8712 , n8710 , n8711 );
xnor ( n8713 , n8712 , n7611 );
and ( n8714 , n8709 , n8713 );
and ( n8715 , n7696 , n7866 );
and ( n8716 , n7828 , n7864 );
nor ( n8717 , n8715 , n8716 );
xnor ( n8718 , n8717 , n7876 );
and ( n8719 , n8713 , n8718 );
and ( n8720 , n8709 , n8718 );
or ( n8721 , n8714 , n8719 , n8720 );
and ( n8722 , n8049 , n7395 );
and ( n8723 , n8108 , n7393 );
nor ( n8724 , n8722 , n8723 );
xnor ( n8725 , n8724 , n7405 );
and ( n8726 , n8721 , n8725 );
and ( n8727 , n7786 , n7899 );
and ( n8728 , n8035 , n7897 );
nor ( n8729 , n8727 , n8728 );
xnor ( n8730 , n8729 , n7909 );
and ( n8731 , n8725 , n8730 );
and ( n8732 , n8721 , n8730 );
or ( n8733 , n8726 , n8731 , n8732 );
and ( n8734 , n7400 , n7318 );
and ( n8735 , n8306 , n7315 );
nor ( n8736 , n8734 , n8735 );
xnor ( n8737 , n8736 , n7311 );
and ( n8738 , n8733 , n8737 );
xor ( n8739 , n8518 , n8532 );
xor ( n8740 , n8739 , n8535 );
and ( n8741 , n8737 , n8740 );
and ( n8742 , n8733 , n8740 );
or ( n8743 , n8738 , n8741 , n8742 );
and ( n8744 , n8687 , n8743 );
xor ( n8745 , n8466 , n8480 );
xor ( n8746 , n8745 , n8483 );
and ( n8747 , n8743 , n8746 );
and ( n8748 , n8687 , n8746 );
or ( n8749 , n8744 , n8747 , n8748 );
and ( n8750 , n8639 , n8749 );
xor ( n8751 , n8328 , n8332 );
xor ( n8752 , n8751 , n8335 );
and ( n8753 , n8749 , n8752 );
and ( n8754 , n8639 , n8752 );
or ( n8755 , n8750 , n8753 , n8754 );
and ( n8756 , n8627 , n8755 );
xor ( n8757 , n8486 , n8488 );
xor ( n8758 , n8757 , n8491 );
and ( n8759 , n7762 , n7899 );
and ( n8760 , n7786 , n7897 );
nor ( n8761 , n8759 , n8760 );
xnor ( n8762 , n8761 , n7909 );
and ( n8763 , n7547 , n7933 );
and ( n8764 , n7410 , n7931 );
nor ( n8765 , n8763 , n8764 );
xnor ( n8766 , n8765 , n7939 );
and ( n8767 , n8762 , n8766 );
xor ( n8768 , n8421 , n8434 );
xor ( n8769 , n8768 , n8439 );
and ( n8770 , n8766 , n8769 );
and ( n8771 , n8762 , n8769 );
or ( n8772 , n8767 , n8770 , n8771 );
xor ( n8773 , n8506 , n8510 );
xor ( n8774 , n8773 , n8515 );
and ( n8775 , n8772 , n8774 );
xor ( n8776 , n8542 , n8546 );
xor ( n8777 , n8776 , n8551 );
and ( n8778 , n8774 , n8777 );
and ( n8779 , n8772 , n8777 );
or ( n8780 , n8775 , n8778 , n8779 );
and ( n8781 , n7352 , n7318 );
and ( n8782 , n7400 , n7315 );
nor ( n8783 , n8781 , n8782 );
xnor ( n8784 , n8783 , n7311 );
and ( n8785 , n7885 , n8168 );
and ( n8786 , n7904 , n8166 );
nor ( n8787 , n8785 , n8786 );
xnor ( n8788 , n8787 , n8178 );
and ( n8789 , n8784 , n8788 );
xor ( n8790 , n8522 , n8526 );
xor ( n8791 , n8790 , n8529 );
and ( n8792 , n8788 , n8791 );
and ( n8793 , n8784 , n8791 );
or ( n8794 , n8789 , n8792 , n8793 );
and ( n8795 , n8780 , n8794 );
xor ( n8796 , n8470 , n8474 );
xor ( n8797 , n8796 , n8477 );
and ( n8798 , n8794 , n8797 );
and ( n8799 , n8780 , n8797 );
or ( n8800 , n8795 , n8798 , n8799 );
xor ( n8801 , n8538 , n8562 );
xor ( n8802 , n8801 , n8565 );
and ( n8803 , n8800 , n8802 );
xor ( n8804 , n8631 , n8633 );
xor ( n8805 , n8804 , n8636 );
and ( n8806 , n8802 , n8805 );
and ( n8807 , n8800 , n8805 );
or ( n8808 , n8803 , n8806 , n8807 );
and ( n8809 , n8758 , n8808 );
xor ( n8810 , n8499 , n8501 );
xor ( n8811 , n8810 , n8568 );
and ( n8812 , n8808 , n8811 );
and ( n8813 , n8758 , n8811 );
or ( n8814 , n8809 , n8812 , n8813 );
and ( n8815 , n8755 , n8814 );
and ( n8816 , n8627 , n8814 );
or ( n8817 , n8756 , n8815 , n8816 );
and ( n8818 , n8626 , n8817 );
xor ( n8819 , n8226 , n8415 );
xor ( n8820 , n8819 , n8574 );
and ( n8821 , n8817 , n8820 );
and ( n8822 , n8626 , n8820 );
or ( n8823 , n8818 , n8821 , n8822 );
xor ( n8824 , n8577 , n8823 );
and ( n8825 , n8585 , n8589 );
and ( n8826 , n8589 , n8624 );
and ( n8827 , n8585 , n8624 );
or ( n8828 , n8825 , n8826 , n8827 );
and ( n8829 , n7348 , n7997 );
and ( n8830 , n7997 , n8225 );
and ( n8831 , n7348 , n8225 );
or ( n8832 , n8829 , n8830 , n8831 );
xor ( n8833 , n8828 , n8832 );
and ( n8834 , n7345 , n7318 );
and ( n8835 , n7323 , n7326 );
and ( n8836 , n7326 , n7329 );
and ( n8837 , n7323 , n7329 );
or ( n8838 , n8835 , n8836 , n8837 );
buf ( n8839 , n7328 );
not ( n8840 , n1671 );
xor ( n8841 , n8839 , n8840 );
and ( n8842 , n1636 , n1657 );
xor ( n8843 , n8841 , n8842 );
xor ( n8844 , n8838 , n8843 );
and ( n8845 , n7330 , n7334 );
and ( n8846 , n7334 , n7339 );
and ( n8847 , n7330 , n7339 );
or ( n8848 , n8845 , n8846 , n8847 );
xor ( n8849 , n8844 , n8848 );
and ( n8850 , n7340 , n7341 );
xor ( n8851 , n8849 , n8850 );
buf ( n8852 , n8851 );
buf ( n8853 , n8852 );
buf ( n8854 , n8853 );
and ( n8855 , n8854 , n7315 );
nor ( n8856 , n8834 , n8855 );
xnor ( n8857 , n8856 , n7311 );
xor ( n8858 , n8833 , n8857 );
and ( n8859 , n8155 , n8179 );
and ( n8860 , n8179 , n8224 );
and ( n8861 , n8155 , n8224 );
or ( n8862 , n8859 , n8860 , n8861 );
and ( n8863 , n8594 , n8598 );
and ( n8864 , n8598 , n8623 );
and ( n8865 , n8594 , n8623 );
or ( n8866 , n8863 , n8864 , n8865 );
and ( n8867 , n7758 , n7969 );
and ( n8868 , n7969 , n7996 );
and ( n8869 , n7758 , n7996 );
or ( n8870 , n8867 , n8868 , n8869 );
xor ( n8871 , n8866 , n8870 );
and ( n8872 , n8203 , n8207 );
and ( n8873 , n8207 , n8222 );
and ( n8874 , n8203 , n8222 );
or ( n8875 , n8872 , n8873 , n8874 );
and ( n8876 , n8212 , n8216 );
and ( n8877 , n8216 , n8221 );
and ( n8878 , n8212 , n8221 );
or ( n8879 , n8876 , n8877 , n8878 );
and ( n8880 , n8049 , n7781 );
and ( n8881 , n8108 , n7779 );
nor ( n8882 , n8880 , n8881 );
xnor ( n8883 , n8882 , n7791 );
xor ( n8884 , n8879 , n8883 );
and ( n8885 , n7410 , n7542 );
and ( n8886 , n7506 , n7540 );
nor ( n8887 , n8885 , n8886 );
xnor ( n8888 , n8887 , n7552 );
xor ( n8889 , n8884 , n8888 );
xor ( n8890 , n8875 , n8889 );
and ( n8891 , n8612 , n8616 );
and ( n8892 , n8616 , n8621 );
and ( n8893 , n8612 , n8621 );
or ( n8894 , n8891 , n8892 , n8893 );
and ( n8895 , n7988 , n7989 );
and ( n8896 , n7989 , n7994 );
and ( n8897 , n7988 , n7994 );
or ( n8898 , n8895 , n8896 , n8897 );
xor ( n8899 , n8894 , n8898 );
and ( n8900 , n7786 , n7933 );
and ( n8901 , n8035 , n7931 );
nor ( n8902 , n8900 , n8901 );
xnor ( n8903 , n8902 , n7939 );
xor ( n8904 , n8899 , n8903 );
xor ( n8905 , n8890 , n8904 );
xor ( n8906 , n8871 , n8905 );
xor ( n8907 , n8862 , n8906 );
and ( n8908 , n8173 , n8168 );
and ( n8909 , n7301 , n8166 );
nor ( n8910 , n8908 , n8909 );
xnor ( n8911 , n8910 , n8178 );
and ( n8912 , n8603 , n8607 );
and ( n8913 , n8607 , n8622 );
and ( n8914 , n8603 , n8622 );
or ( n8915 , n8912 , n8913 , n8914 );
and ( n8916 , n7974 , n7978 );
and ( n8917 , n7978 , n7995 );
and ( n8918 , n7974 , n7995 );
or ( n8919 , n8916 , n8917 , n8918 );
xor ( n8920 , n8915 , n8919 );
and ( n8921 , n8306 , n7395 );
and ( n8922 , n8159 , n7393 );
nor ( n8923 , n8921 , n8922 );
xnor ( n8924 , n8923 , n7405 );
xor ( n8925 , n8920 , n8924 );
xor ( n8926 , n8911 , n8925 );
and ( n8927 , n8184 , n8198 );
and ( n8928 , n8198 , n8223 );
and ( n8929 , n8184 , n8223 );
or ( n8930 , n8927 , n8928 , n8929 );
and ( n8931 , n7885 , n8044 );
and ( n8932 , n7904 , n8042 );
nor ( n8933 , n8931 , n8932 );
xnor ( n8934 , n8933 , n8054 );
and ( n8935 , n7704 , n7601 );
and ( n8936 , n7718 , n7599 );
nor ( n8937 , n8935 , n8936 );
xnor ( n8938 , n8937 , n7611 );
and ( n8939 , n7558 , n7743 );
and ( n8940 , n7606 , n7741 );
nor ( n8941 , n8939 , n8940 );
xnor ( n8942 , n8941 , n7753 );
xor ( n8943 , n8938 , n8942 );
and ( n8944 , n7729 , n7866 );
and ( n8945 , n7748 , n7864 );
nor ( n8946 , n8944 , n8945 );
xnor ( n8947 , n8946 , n7876 );
xor ( n8948 , n8943 , n8947 );
xor ( n8949 , n8934 , n8948 );
and ( n8950 , n7983 , n7987 );
and ( n8951 , n7516 , n7713 );
and ( n8952 , n7547 , n7711 );
nor ( n8953 , n8951 , n8952 );
xnor ( n8954 , n8953 , n7723 );
xor ( n8955 , n8950 , n8954 );
and ( n8956 , n7828 , n7691 );
and ( n8957 , n7809 , n7689 );
nor ( n8958 , n8956 , n8957 );
not ( n8959 , n8958 );
xor ( n8960 , n8955 , n8959 );
xor ( n8961 , n8949 , n8960 );
xor ( n8962 , n8930 , n8961 );
and ( n8963 , n8188 , n8192 );
and ( n8964 , n8192 , n8197 );
and ( n8965 , n8188 , n8197 );
or ( n8966 , n8963 , n8964 , n8965 );
and ( n8967 , n7352 , n7899 );
and ( n8968 , n7400 , n7897 );
nor ( n8969 , n8967 , n8968 );
xnor ( n8970 , n8969 , n7909 );
xor ( n8971 , n8966 , n8970 );
and ( n8972 , n7945 , n7501 );
and ( n8973 , n7959 , n7499 );
nor ( n8974 , n8972 , n8973 );
xnor ( n8975 , n8974 , n7511 );
xor ( n8976 , n8971 , n8975 );
and ( n8977 , n7919 , n7954 );
and ( n8978 , n7762 , n7952 );
nor ( n8979 , n8977 , n8978 );
xnor ( n8980 , n8979 , n7964 );
and ( n8981 , n7871 , n7661 );
and ( n8982 , n7800 , n7659 );
nor ( n8983 , n8981 , n8982 );
xnor ( n8984 , n8983 , n7671 );
xor ( n8985 , n8980 , n8984 );
and ( n8986 , n7618 , n7823 );
and ( n8987 , n7666 , n7821 );
nor ( n8988 , n8986 , n8987 );
xnor ( n8989 , n8988 , n7833 );
xor ( n8990 , n8985 , n8989 );
xor ( n8991 , n8976 , n8990 );
xor ( n8992 , n8962 , n8991 );
xor ( n8993 , n8926 , n8992 );
xor ( n8994 , n8907 , n8993 );
xor ( n8995 , n8858 , n8994 );
and ( n8996 , n8581 , n8625 );
xor ( n8997 , n8995 , n8996 );
xor ( n8998 , n8824 , n8997 );
xor ( n8999 , n8420 , n8494 );
xor ( n9000 , n8999 , n8571 );
and ( n9001 , n7516 , n7933 );
and ( n9002 , n7547 , n7931 );
nor ( n9003 , n9001 , n9002 );
xnor ( n9004 , n9003 , n7939 );
and ( n9005 , n7871 , n7713 );
and ( n9006 , n7800 , n7711 );
nor ( n9007 , n9005 , n9006 );
xnor ( n9008 , n9007 , n7723 );
and ( n9009 , n9004 , n9008 );
and ( n9010 , n7828 , n7743 );
and ( n9011 , n7809 , n7741 );
nor ( n9012 , n9010 , n9011 );
xnor ( n9013 , n9012 , n7753 );
and ( n9014 , n9008 , n9013 );
and ( n9015 , n9004 , n9013 );
or ( n9016 , n9009 , n9014 , n9015 );
and ( n9017 , n7704 , n7954 );
and ( n9018 , n7718 , n7952 );
nor ( n9019 , n9017 , n9018 );
xnor ( n9020 , n9019 , n7964 );
and ( n9021 , n7558 , n7501 );
and ( n9022 , n7606 , n7499 );
nor ( n9023 , n9021 , n9022 );
xnor ( n9024 , n9023 , n7511 );
and ( n9025 , n9020 , n9024 );
and ( n9026 , n7729 , n7542 );
and ( n9027 , n7748 , n7540 );
nor ( n9028 , n9026 , n9027 );
xnor ( n9029 , n9028 , n7552 );
and ( n9030 , n9024 , n9029 );
and ( n9031 , n9020 , n9029 );
or ( n9032 , n9025 , n9030 , n9031 );
and ( n9033 , n9016 , n9032 );
and ( n9034 , n8108 , n8168 );
and ( n9035 , n7885 , n8166 );
nor ( n9036 , n9034 , n9035 );
xnor ( n9037 , n9036 , n8178 );
and ( n9038 , n9032 , n9037 );
and ( n9039 , n9016 , n9037 );
or ( n9040 , n9033 , n9038 , n9039 );
xor ( n9041 , n8692 , n8700 );
and ( n9042 , n8079 , n7661 );
and ( n9043 , n8066 , n7659 );
nor ( n9044 , n9042 , n9043 );
xnor ( n9045 , n9044 , n7671 );
xor ( n9046 , n6616 , n7252 );
buf ( n9047 , n9046 );
buf ( n9048 , n9047 );
buf ( n9049 , n9048 );
and ( n9050 , n9049 , n7691 );
and ( n9051 , n8696 , n7689 );
nor ( n9052 , n9050 , n9051 );
not ( n9053 , n9052 );
and ( n9054 , n9045 , n9053 );
and ( n9055 , n9041 , n9054 );
and ( n9056 , n8263 , n7823 );
and ( n9057 , n8079 , n7821 );
nor ( n9058 , n9056 , n9057 );
xnor ( n9059 , n9058 , n7833 );
and ( n9060 , n9054 , n9059 );
and ( n9061 , n9041 , n9059 );
or ( n9062 , n9055 , n9060 , n9061 );
and ( n9063 , n7618 , n7601 );
and ( n9064 , n7666 , n7599 );
nor ( n9065 , n9063 , n9064 );
xnor ( n9066 , n9065 , n7611 );
and ( n9067 , n9062 , n9066 );
and ( n9068 , n7851 , n7661 );
and ( n9069 , n7838 , n7659 );
nor ( n9070 , n9068 , n9069 );
xnor ( n9071 , n9070 , n7671 );
and ( n9072 , n9066 , n9071 );
and ( n9073 , n9062 , n9071 );
or ( n9074 , n9067 , n9072 , n9073 );
and ( n9075 , n7506 , n7781 );
and ( n9076 , n7945 , n7779 );
nor ( n9077 , n9075 , n9076 );
xnor ( n9078 , n9077 , n7791 );
and ( n9079 , n9074 , n9078 );
xor ( n9080 , n8709 , n8713 );
xor ( n9081 , n9080 , n8718 );
and ( n9082 , n9078 , n9081 );
and ( n9083 , n9074 , n9081 );
or ( n9084 , n9079 , n9082 , n9083 );
and ( n9085 , n9040 , n9084 );
xor ( n9086 , n8655 , n8671 );
xor ( n9087 , n9086 , n8674 );
and ( n9088 , n9084 , n9087 );
and ( n9089 , n9040 , n9087 );
or ( n9090 , n9085 , n9088 , n9089 );
xor ( n9091 , n8554 , n8556 );
xor ( n9092 , n9091 , n8559 );
and ( n9093 , n9090 , n9092 );
xor ( n9094 , n8677 , n8681 );
xor ( n9095 , n9094 , n8684 );
and ( n9096 , n9092 , n9095 );
and ( n9097 , n9090 , n9095 );
or ( n9098 , n9093 , n9096 , n9097 );
and ( n9099 , n8035 , n7395 );
and ( n9100 , n8049 , n7393 );
nor ( n9101 , n9099 , n9100 );
xnor ( n9102 , n9101 , n7405 );
xor ( n9103 , n8643 , n8647 );
xor ( n9104 , n9103 , n8652 );
and ( n9105 , n9102 , n9104 );
xor ( n9106 , n8762 , n8766 );
xor ( n9107 , n9106 , n8769 );
and ( n9108 , n9104 , n9107 );
and ( n9109 , n9102 , n9107 );
or ( n9110 , n9105 , n9108 , n9109 );
xor ( n9111 , n8721 , n8725 );
xor ( n9112 , n9111 , n8730 );
and ( n9113 , n9110 , n9112 );
xor ( n9114 , n8772 , n8774 );
xor ( n9115 , n9114 , n8777 );
and ( n9116 , n9112 , n9115 );
and ( n9117 , n9110 , n9115 );
or ( n9118 , n9113 , n9116 , n9117 );
xor ( n9119 , n8780 , n8794 );
xor ( n9120 , n9119 , n8797 );
and ( n9121 , n9118 , n9120 );
xor ( n9122 , n8733 , n8737 );
xor ( n9123 , n9122 , n8740 );
and ( n9124 , n9120 , n9123 );
and ( n9125 , n9118 , n9123 );
or ( n9126 , n9121 , n9124 , n9125 );
and ( n9127 , n9098 , n9126 );
xor ( n9128 , n8687 , n8743 );
xor ( n9129 , n9128 , n8746 );
and ( n9130 , n9126 , n9129 );
and ( n9131 , n9098 , n9129 );
or ( n9132 , n9127 , n9130 , n9131 );
xor ( n9133 , n8639 , n8749 );
xor ( n9134 , n9133 , n8752 );
and ( n9135 , n9132 , n9134 );
and ( n9136 , n9000 , n9135 );
xor ( n9137 , n8627 , n8755 );
xor ( n9138 , n9137 , n8814 );
and ( n9139 , n9135 , n9138 );
and ( n9140 , n9000 , n9138 );
or ( n9141 , n9136 , n9139 , n9140 );
xor ( n9142 , n8626 , n8817 );
xor ( n9143 , n9142 , n8820 );
and ( n9144 , n9141 , n9143 );
xor ( n9145 , n9141 , n9143 );
xor ( n9146 , n9000 , n9135 );
xor ( n9147 , n9146 , n9138 );
xor ( n9148 , n8758 , n8808 );
xor ( n9149 , n9148 , n8811 );
xor ( n9150 , n9132 , n9134 );
and ( n9151 , n9149 , n9150 );
and ( n9152 , n7666 , n7713 );
and ( n9153 , n7871 , n7711 );
nor ( n9154 , n9152 , n9153 );
xnor ( n9155 , n9154 , n7723 );
and ( n9156 , n7696 , n7743 );
and ( n9157 , n7828 , n7741 );
nor ( n9158 , n9156 , n9157 );
xnor ( n9159 , n9158 , n7753 );
and ( n9160 , n9155 , n9159 );
and ( n9161 , n7838 , n7866 );
and ( n9162 , n7676 , n7864 );
nor ( n9163 , n9161 , n9162 );
xnor ( n9164 , n9163 , n7876 );
and ( n9165 , n9159 , n9164 );
and ( n9166 , n9155 , n9164 );
or ( n9167 , n9160 , n9165 , n9166 );
and ( n9168 , n7945 , n8044 );
and ( n9169 , n7959 , n8042 );
nor ( n9170 , n9168 , n9169 );
xnor ( n9171 , n9170 , n8054 );
and ( n9172 , n9167 , n9171 );
xor ( n9173 , n8688 , n8701 );
xor ( n9174 , n9173 , n8706 );
and ( n9175 , n9171 , n9174 );
and ( n9176 , n9167 , n9174 );
or ( n9177 , n9172 , n9175 , n9176 );
and ( n9178 , n7904 , n7318 );
and ( n9179 , n7352 , n7315 );
nor ( n9180 , n9178 , n9179 );
xnor ( n9181 , n9180 , n7311 );
and ( n9182 , n9177 , n9181 );
xor ( n9183 , n8659 , n8663 );
xor ( n9184 , n9183 , n8668 );
and ( n9185 , n9181 , n9184 );
and ( n9186 , n9177 , n9184 );
or ( n9187 , n9182 , n9185 , n9186 );
xor ( n9188 , n9045 , n9053 );
and ( n9189 , n8696 , n7823 );
and ( n9190 , n8429 , n7821 );
nor ( n9191 , n9189 , n9190 );
xnor ( n9192 , n9191 , n7833 );
xor ( n9193 , n6686 , n7250 );
buf ( n9194 , n9193 );
buf ( n9195 , n9194 );
buf ( n9196 , n9195 );
and ( n9197 , n9196 , n7691 );
and ( n9198 , n9049 , n7689 );
nor ( n9199 , n9197 , n9198 );
not ( n9200 , n9199 );
and ( n9201 , n9192 , n9200 );
and ( n9202 , n9188 , n9201 );
and ( n9203 , n8429 , n7823 );
and ( n9204 , n8263 , n7821 );
nor ( n9205 , n9203 , n9204 );
xnor ( n9206 , n9205 , n7833 );
and ( n9207 , n9201 , n9206 );
and ( n9208 , n9188 , n9206 );
or ( n9209 , n9202 , n9207 , n9208 );
and ( n9210 , n7800 , n7542 );
and ( n9211 , n7729 , n7540 );
nor ( n9212 , n9210 , n9211 );
xnor ( n9213 , n9212 , n7552 );
and ( n9214 , n9209 , n9213 );
and ( n9215 , n7809 , n7601 );
and ( n9216 , n7618 , n7599 );
nor ( n9217 , n9215 , n9216 );
xnor ( n9218 , n9217 , n7611 );
and ( n9219 , n9213 , n9218 );
and ( n9220 , n9209 , n9218 );
or ( n9221 , n9214 , n9219 , n9220 );
and ( n9222 , n7919 , n7899 );
and ( n9223 , n7762 , n7897 );
nor ( n9224 , n9222 , n9223 );
xnor ( n9225 , n9224 , n7909 );
and ( n9226 , n9221 , n9225 );
and ( n9227 , n7410 , n7781 );
and ( n9228 , n7506 , n7779 );
nor ( n9229 , n9227 , n9228 );
xnor ( n9230 , n9229 , n7791 );
and ( n9231 , n9225 , n9230 );
and ( n9232 , n9221 , n9230 );
or ( n9233 , n9226 , n9231 , n9232 );
and ( n9234 , n7547 , n7781 );
and ( n9235 , n7410 , n7779 );
nor ( n9236 , n9234 , n9235 );
xnor ( n9237 , n9236 , n7791 );
and ( n9238 , n7718 , n7933 );
and ( n9239 , n7516 , n7931 );
nor ( n9240 , n9238 , n9239 );
xnor ( n9241 , n9240 , n7939 );
and ( n9242 , n9237 , n9241 );
and ( n9243 , n7606 , n7954 );
and ( n9244 , n7704 , n7952 );
nor ( n9245 , n9243 , n9244 );
xnor ( n9246 , n9245 , n7964 );
and ( n9247 , n9241 , n9246 );
and ( n9248 , n9237 , n9246 );
or ( n9249 , n9242 , n9247 , n9248 );
and ( n9250 , n8049 , n8168 );
and ( n9251 , n8108 , n8166 );
nor ( n9252 , n9250 , n9251 );
xnor ( n9253 , n9252 , n8178 );
and ( n9254 , n9249 , n9253 );
xor ( n9255 , n9062 , n9066 );
xor ( n9256 , n9255 , n9071 );
and ( n9257 , n9253 , n9256 );
and ( n9258 , n9249 , n9256 );
or ( n9259 , n9254 , n9257 , n9258 );
and ( n9260 , n9233 , n9259 );
xor ( n9261 , n9074 , n9078 );
xor ( n9262 , n9261 , n9081 );
and ( n9263 , n9259 , n9262 );
and ( n9264 , n9233 , n9262 );
or ( n9265 , n9260 , n9263 , n9264 );
and ( n9266 , n9187 , n9265 );
xor ( n9267 , n8784 , n8788 );
xor ( n9268 , n9267 , n8791 );
and ( n9269 , n9265 , n9268 );
and ( n9270 , n9187 , n9268 );
or ( n9271 , n9266 , n9269 , n9270 );
xor ( n9272 , n9192 , n9200 );
and ( n9273 , n9049 , n7823 );
and ( n9274 , n8696 , n7821 );
nor ( n9275 , n9273 , n9274 );
xnor ( n9276 , n9275 , n7833 );
xor ( n9277 , n7069 , n7248 );
buf ( n9278 , n9277 );
buf ( n9279 , n9278 );
buf ( n9280 , n9279 );
and ( n9281 , n9280 , n7691 );
and ( n9282 , n9196 , n7689 );
nor ( n9283 , n9281 , n9282 );
not ( n9284 , n9283 );
and ( n9285 , n9276 , n9284 );
and ( n9286 , n9272 , n9285 );
and ( n9287 , n8066 , n7866 );
and ( n9288 , n7851 , n7864 );
nor ( n9289 , n9287 , n9288 );
xnor ( n9290 , n9289 , n7876 );
and ( n9291 , n9285 , n9290 );
and ( n9292 , n9272 , n9290 );
or ( n9293 , n9286 , n9291 , n9292 );
and ( n9294 , n7676 , n7743 );
and ( n9295 , n7696 , n7741 );
nor ( n9296 , n9294 , n9295 );
xnor ( n9297 , n9296 , n7753 );
and ( n9298 , n9293 , n9297 );
and ( n9299 , n7851 , n7866 );
and ( n9300 , n7838 , n7864 );
nor ( n9301 , n9299 , n9300 );
xnor ( n9302 , n9301 , n7876 );
and ( n9303 , n9297 , n9302 );
and ( n9304 , n9293 , n9302 );
or ( n9305 , n9298 , n9303 , n9304 );
and ( n9306 , n7959 , n7899 );
and ( n9307 , n7919 , n7897 );
nor ( n9308 , n9306 , n9307 );
xnor ( n9309 , n9308 , n7909 );
and ( n9310 , n9305 , n9309 );
and ( n9311 , n7748 , n7501 );
and ( n9312 , n7558 , n7499 );
nor ( n9313 , n9311 , n9312 );
xnor ( n9314 , n9313 , n7511 );
and ( n9315 , n9309 , n9314 );
and ( n9316 , n9305 , n9314 );
or ( n9317 , n9310 , n9315 , n9316 );
and ( n9318 , n7786 , n7395 );
and ( n9319 , n8035 , n7393 );
nor ( n9320 , n9318 , n9319 );
xnor ( n9321 , n9320 , n7405 );
and ( n9322 , n9317 , n9321 );
xor ( n9323 , n9004 , n9008 );
xor ( n9324 , n9323 , n9013 );
and ( n9325 , n9321 , n9324 );
and ( n9326 , n9317 , n9324 );
or ( n9327 , n9322 , n9325 , n9326 );
xor ( n9328 , n9016 , n9032 );
xor ( n9329 , n9328 , n9037 );
and ( n9330 , n9327 , n9329 );
xor ( n9331 , n9102 , n9104 );
xor ( n9332 , n9331 , n9107 );
and ( n9333 , n9329 , n9332 );
and ( n9334 , n9327 , n9332 );
or ( n9335 , n9330 , n9333 , n9334 );
xor ( n9336 , n9040 , n9084 );
xor ( n9337 , n9336 , n9087 );
and ( n9338 , n9335 , n9337 );
xor ( n9339 , n9110 , n9112 );
xor ( n9340 , n9339 , n9115 );
and ( n9341 , n9337 , n9340 );
and ( n9342 , n9335 , n9340 );
or ( n9343 , n9338 , n9341 , n9342 );
and ( n9344 , n9271 , n9343 );
xor ( n9345 , n9090 , n9092 );
xor ( n9346 , n9345 , n9095 );
and ( n9347 , n9343 , n9346 );
and ( n9348 , n9271 , n9346 );
or ( n9349 , n9344 , n9347 , n9348 );
xor ( n9350 , n8800 , n8802 );
xor ( n9351 , n9350 , n8805 );
and ( n9352 , n9349 , n9351 );
xor ( n9353 , n9098 , n9126 );
xor ( n9354 , n9353 , n9129 );
and ( n9355 , n9351 , n9354 );
and ( n9356 , n9349 , n9354 );
or ( n9357 , n9352 , n9355 , n9356 );
and ( n9358 , n9150 , n9357 );
and ( n9359 , n9149 , n9357 );
or ( n9360 , n9151 , n9358 , n9359 );
and ( n9361 , n9147 , n9360 );
xor ( n9362 , n9147 , n9360 );
xor ( n9363 , n9149 , n9150 );
xor ( n9364 , n9363 , n9357 );
xor ( n9365 , n9349 , n9351 );
xor ( n9366 , n9365 , n9354 );
and ( n9367 , n7762 , n7395 );
and ( n9368 , n7786 , n7393 );
nor ( n9369 , n9367 , n9368 );
xnor ( n9370 , n9369 , n7405 );
and ( n9371 , n7506 , n8044 );
and ( n9372 , n7945 , n8042 );
nor ( n9373 , n9371 , n9372 );
xnor ( n9374 , n9373 , n8054 );
and ( n9375 , n9370 , n9374 );
xor ( n9376 , n9041 , n9054 );
xor ( n9377 , n9376 , n9059 );
and ( n9378 , n9374 , n9377 );
and ( n9379 , n9370 , n9377 );
or ( n9380 , n9375 , n9378 , n9379 );
and ( n9381 , n7885 , n7318 );
and ( n9382 , n7904 , n7315 );
nor ( n9383 , n9381 , n9382 );
xnor ( n9384 , n9383 , n7311 );
and ( n9385 , n9380 , n9384 );
xor ( n9386 , n9020 , n9024 );
xor ( n9387 , n9386 , n9029 );
and ( n9388 , n9384 , n9387 );
and ( n9389 , n9380 , n9387 );
or ( n9390 , n9385 , n9388 , n9389 );
and ( n9391 , n7871 , n7542 );
and ( n9392 , n7800 , n7540 );
nor ( n9393 , n9391 , n9392 );
xnor ( n9394 , n9393 , n7552 );
and ( n9395 , n7618 , n7713 );
and ( n9396 , n7666 , n7711 );
nor ( n9397 , n9395 , n9396 );
xnor ( n9398 , n9397 , n7723 );
and ( n9399 , n9394 , n9398 );
and ( n9400 , n7828 , n7601 );
and ( n9401 , n7809 , n7599 );
nor ( n9402 , n9400 , n9401 );
xnor ( n9403 , n9402 , n7611 );
and ( n9404 , n9398 , n9403 );
and ( n9405 , n9394 , n9403 );
or ( n9406 , n9399 , n9404 , n9405 );
and ( n9407 , n8035 , n8168 );
and ( n9408 , n8049 , n8166 );
nor ( n9409 , n9407 , n9408 );
xnor ( n9410 , n9409 , n8178 );
and ( n9411 , n9406 , n9410 );
xor ( n9412 , n9155 , n9159 );
xor ( n9413 , n9412 , n9164 );
and ( n9414 , n9410 , n9413 );
and ( n9415 , n9406 , n9413 );
or ( n9416 , n9411 , n9414 , n9415 );
xor ( n9417 , n9221 , n9225 );
xor ( n9418 , n9417 , n9230 );
and ( n9419 , n9416 , n9418 );
xor ( n9420 , n9167 , n9171 );
xor ( n9421 , n9420 , n9174 );
and ( n9422 , n9418 , n9421 );
and ( n9423 , n9416 , n9421 );
or ( n9424 , n9419 , n9422 , n9423 );
and ( n9425 , n9390 , n9424 );
xor ( n9426 , n9177 , n9181 );
xor ( n9427 , n9426 , n9184 );
and ( n9428 , n9424 , n9427 );
and ( n9429 , n9390 , n9427 );
or ( n9430 , n9425 , n9428 , n9429 );
and ( n9431 , n7516 , n7781 );
and ( n9432 , n7547 , n7779 );
nor ( n9433 , n9431 , n9432 );
xnor ( n9434 , n9433 , n7791 );
and ( n9435 , n7729 , n7501 );
and ( n9436 , n7748 , n7499 );
nor ( n9437 , n9435 , n9436 );
xnor ( n9438 , n9437 , n7511 );
and ( n9439 , n9434 , n9438 );
xor ( n9440 , n9188 , n9201 );
xor ( n9441 , n9440 , n9206 );
and ( n9442 , n9438 , n9441 );
and ( n9443 , n9434 , n9441 );
or ( n9444 , n9439 , n9442 , n9443 );
and ( n9445 , n8108 , n7318 );
and ( n9446 , n7885 , n7315 );
nor ( n9447 , n9445 , n9446 );
xnor ( n9448 , n9447 , n7311 );
and ( n9449 , n9444 , n9448 );
xor ( n9450 , n9209 , n9213 );
xor ( n9451 , n9450 , n9218 );
and ( n9452 , n9448 , n9451 );
and ( n9453 , n9444 , n9451 );
or ( n9454 , n9449 , n9452 , n9453 );
xor ( n9455 , n9276 , n9284 );
and ( n9456 , n8696 , n7661 );
and ( n9457 , n8429 , n7659 );
nor ( n9458 , n9456 , n9457 );
xnor ( n9459 , n9458 , n7671 );
xor ( n9460 , n7071 , n7247 );
buf ( n9461 , n9460 );
buf ( n9462 , n9461 );
buf ( n9463 , n9462 );
and ( n9464 , n9463 , n7691 );
and ( n9465 , n9280 , n7689 );
nor ( n9466 , n9464 , n9465 );
not ( n9467 , n9466 );
and ( n9468 , n9459 , n9467 );
and ( n9469 , n9455 , n9468 );
and ( n9470 , n8079 , n7866 );
and ( n9471 , n8066 , n7864 );
nor ( n9472 , n9470 , n9471 );
xnor ( n9473 , n9472 , n7876 );
and ( n9474 , n9468 , n9473 );
and ( n9475 , n9455 , n9473 );
or ( n9476 , n9469 , n9474 , n9475 );
and ( n9477 , n7838 , n7743 );
and ( n9478 , n7676 , n7741 );
nor ( n9479 , n9477 , n9478 );
xnor ( n9480 , n9479 , n7753 );
and ( n9481 , n9476 , n9480 );
and ( n9482 , n8263 , n7661 );
and ( n9483 , n8079 , n7659 );
nor ( n9484 , n9482 , n9483 );
xnor ( n9485 , n9484 , n7671 );
and ( n9486 , n9480 , n9485 );
and ( n9487 , n9476 , n9485 );
or ( n9488 , n9481 , n9486 , n9487 );
and ( n9489 , n7704 , n7933 );
and ( n9490 , n7718 , n7931 );
nor ( n9491 , n9489 , n9490 );
xnor ( n9492 , n9491 , n7939 );
and ( n9493 , n9488 , n9492 );
and ( n9494 , n7558 , n7954 );
and ( n9495 , n7606 , n7952 );
nor ( n9496 , n9494 , n9495 );
xnor ( n9497 , n9496 , n7964 );
and ( n9498 , n9492 , n9497 );
and ( n9499 , n9488 , n9497 );
or ( n9500 , n9493 , n9498 , n9499 );
and ( n9501 , n7919 , n7395 );
and ( n9502 , n7762 , n7393 );
nor ( n9503 , n9501 , n9502 );
xnor ( n9504 , n9503 , n7405 );
and ( n9505 , n7945 , n7899 );
and ( n9506 , n7959 , n7897 );
nor ( n9507 , n9505 , n9506 );
xnor ( n9508 , n9507 , n7909 );
and ( n9509 , n9504 , n9508 );
xor ( n9510 , n9293 , n9297 );
xor ( n9511 , n9510 , n9302 );
and ( n9512 , n9508 , n9511 );
and ( n9513 , n9504 , n9511 );
or ( n9514 , n9509 , n9512 , n9513 );
and ( n9515 , n9500 , n9514 );
xor ( n9516 , n9237 , n9241 );
xor ( n9517 , n9516 , n9246 );
and ( n9518 , n9514 , n9517 );
and ( n9519 , n9500 , n9517 );
or ( n9520 , n9515 , n9518 , n9519 );
and ( n9521 , n9454 , n9520 );
xor ( n9522 , n9317 , n9321 );
xor ( n9523 , n9522 , n9324 );
and ( n9524 , n9520 , n9523 );
and ( n9525 , n9454 , n9523 );
or ( n9526 , n9521 , n9524 , n9525 );
and ( n9527 , n7676 , n7601 );
and ( n9528 , n7696 , n7599 );
nor ( n9529 , n9527 , n9528 );
xnor ( n9530 , n9529 , n7611 );
and ( n9531 , n7851 , n7743 );
and ( n9532 , n7838 , n7741 );
nor ( n9533 , n9531 , n9532 );
xnor ( n9534 , n9533 , n7753 );
and ( n9535 , n9530 , n9534 );
and ( n9536 , n8429 , n7661 );
and ( n9537 , n8263 , n7659 );
nor ( n9538 , n9536 , n9537 );
xnor ( n9539 , n9538 , n7671 );
and ( n9540 , n9534 , n9539 );
and ( n9541 , n9530 , n9539 );
or ( n9542 , n9535 , n9540 , n9541 );
and ( n9543 , n7800 , n7501 );
and ( n9544 , n7729 , n7499 );
nor ( n9545 , n9543 , n9544 );
xnor ( n9546 , n9545 , n7511 );
and ( n9547 , n9542 , n9546 );
and ( n9548 , n7809 , n7713 );
and ( n9549 , n7618 , n7711 );
nor ( n9550 , n9548 , n9549 );
xnor ( n9551 , n9550 , n7723 );
and ( n9552 , n9546 , n9551 );
and ( n9553 , n9542 , n9551 );
or ( n9554 , n9547 , n9552 , n9553 );
and ( n9555 , n7666 , n7542 );
and ( n9556 , n7871 , n7540 );
nor ( n9557 , n9555 , n9556 );
xnor ( n9558 , n9557 , n7552 );
and ( n9559 , n7696 , n7601 );
and ( n9560 , n7828 , n7599 );
nor ( n9561 , n9559 , n9560 );
xnor ( n9562 , n9561 , n7611 );
and ( n9563 , n9558 , n9562 );
xor ( n9564 , n9272 , n9285 );
xor ( n9565 , n9564 , n9290 );
and ( n9566 , n9562 , n9565 );
and ( n9567 , n9558 , n9565 );
or ( n9568 , n9563 , n9566 , n9567 );
and ( n9569 , n9554 , n9568 );
and ( n9570 , n7410 , n8044 );
and ( n9571 , n7506 , n8042 );
nor ( n9572 , n9570 , n9571 );
xnor ( n9573 , n9572 , n8054 );
and ( n9574 , n9568 , n9573 );
and ( n9575 , n9554 , n9573 );
or ( n9576 , n9569 , n9574 , n9575 );
xor ( n9577 , n9305 , n9309 );
xor ( n9578 , n9577 , n9314 );
and ( n9579 , n9576 , n9578 );
xor ( n9580 , n9370 , n9374 );
xor ( n9581 , n9580 , n9377 );
and ( n9582 , n9578 , n9581 );
and ( n9583 , n9576 , n9581 );
or ( n9584 , n9579 , n9582 , n9583 );
xor ( n9585 , n9249 , n9253 );
xor ( n9586 , n9585 , n9256 );
and ( n9587 , n9584 , n9586 );
xor ( n9588 , n9380 , n9384 );
xor ( n9589 , n9588 , n9387 );
and ( n9590 , n9586 , n9589 );
and ( n9591 , n9584 , n9589 );
or ( n9592 , n9587 , n9590 , n9591 );
and ( n9593 , n9526 , n9592 );
xor ( n9594 , n9233 , n9259 );
xor ( n9595 , n9594 , n9262 );
and ( n9596 , n9592 , n9595 );
and ( n9597 , n9526 , n9595 );
or ( n9598 , n9593 , n9596 , n9597 );
and ( n9599 , n9430 , n9598 );
xor ( n9600 , n9187 , n9265 );
xor ( n9601 , n9600 , n9268 );
and ( n9602 , n9598 , n9601 );
and ( n9603 , n9430 , n9601 );
or ( n9604 , n9599 , n9602 , n9603 );
xor ( n9605 , n9118 , n9120 );
xor ( n9606 , n9605 , n9123 );
and ( n9607 , n9604 , n9606 );
xor ( n9608 , n9271 , n9343 );
xor ( n9609 , n9608 , n9346 );
and ( n9610 , n9606 , n9609 );
and ( n9611 , n9604 , n9609 );
or ( n9612 , n9607 , n9610 , n9611 );
and ( n9613 , n9366 , n9612 );
xor ( n9614 , n9604 , n9606 );
xor ( n9615 , n9614 , n9609 );
xor ( n9616 , n9390 , n9424 );
xor ( n9617 , n9616 , n9427 );
xor ( n9618 , n9327 , n9329 );
xor ( n9619 , n9618 , n9332 );
and ( n9620 , n9617 , n9619 );
xor ( n9621 , n9526 , n9592 );
xor ( n9622 , n9621 , n9595 );
and ( n9623 , n9619 , n9622 );
and ( n9624 , n9617 , n9622 );
or ( n9625 , n9620 , n9623 , n9624 );
xor ( n9626 , n9335 , n9337 );
xor ( n9627 , n9626 , n9340 );
and ( n9628 , n9625 , n9627 );
xor ( n9629 , n9430 , n9598 );
xor ( n9630 , n9629 , n9601 );
and ( n9631 , n9627 , n9630 );
and ( n9632 , n9625 , n9630 );
or ( n9633 , n9628 , n9631 , n9632 );
and ( n9634 , n9615 , n9633 );
xor ( n9635 , n9625 , n9627 );
xor ( n9636 , n9635 , n9630 );
and ( n9637 , n7718 , n7781 );
and ( n9638 , n7516 , n7779 );
nor ( n9639 , n9637 , n9638 );
xnor ( n9640 , n9639 , n7791 );
and ( n9641 , n7606 , n7933 );
and ( n9642 , n7704 , n7931 );
nor ( n9643 , n9641 , n9642 );
xnor ( n9644 , n9643 , n7939 );
and ( n9645 , n9640 , n9644 );
xor ( n9646 , n9476 , n9480 );
xor ( n9647 , n9646 , n9485 );
and ( n9648 , n9644 , n9647 );
and ( n9649 , n9640 , n9647 );
or ( n9650 , n9645 , n9648 , n9649 );
and ( n9651 , n8049 , n7318 );
and ( n9652 , n8108 , n7315 );
nor ( n9653 , n9651 , n9652 );
xnor ( n9654 , n9653 , n7311 );
and ( n9655 , n9650 , n9654 );
and ( n9656 , n7786 , n8168 );
and ( n9657 , n8035 , n8166 );
nor ( n9658 , n9656 , n9657 );
xnor ( n9659 , n9658 , n8178 );
and ( n9660 , n9654 , n9659 );
and ( n9661 , n9650 , n9659 );
or ( n9662 , n9655 , n9660 , n9661 );
and ( n9663 , n7959 , n7395 );
and ( n9664 , n7919 , n7393 );
nor ( n9665 , n9663 , n9664 );
xnor ( n9666 , n9665 , n7405 );
and ( n9667 , n7547 , n8044 );
and ( n9668 , n7410 , n8042 );
nor ( n9669 , n9667 , n9668 );
xnor ( n9670 , n9669 , n8054 );
and ( n9671 , n9666 , n9670 );
and ( n9672 , n7748 , n7954 );
and ( n9673 , n7558 , n7952 );
nor ( n9674 , n9672 , n9673 );
xnor ( n9675 , n9674 , n7964 );
and ( n9676 , n9670 , n9675 );
and ( n9677 , n9666 , n9675 );
or ( n9678 , n9671 , n9676 , n9677 );
xor ( n9679 , n9394 , n9398 );
xor ( n9680 , n9679 , n9403 );
and ( n9681 , n9678 , n9680 );
xor ( n9682 , n9488 , n9492 );
xor ( n9683 , n9682 , n9497 );
and ( n9684 , n9680 , n9683 );
and ( n9685 , n9678 , n9683 );
or ( n9686 , n9681 , n9684 , n9685 );
and ( n9687 , n9662 , n9686 );
xor ( n9688 , n9406 , n9410 );
xor ( n9689 , n9688 , n9413 );
and ( n9690 , n9686 , n9689 );
and ( n9691 , n9662 , n9689 );
or ( n9692 , n9687 , n9690 , n9691 );
xor ( n9693 , n9459 , n9467 );
and ( n9694 , n9049 , n7661 );
and ( n9695 , n8696 , n7659 );
nor ( n9696 , n9694 , n9695 );
xnor ( n9697 , n9696 , n7671 );
xor ( n9698 , n7073 , n7246 );
buf ( n9699 , n9698 );
buf ( n9700 , n9699 );
buf ( n9701 , n9700 );
and ( n9702 , n9701 , n7691 );
and ( n9703 , n9463 , n7689 );
nor ( n9704 , n9702 , n9703 );
not ( n9705 , n9704 );
and ( n9706 , n9697 , n9705 );
and ( n9707 , n9693 , n9706 );
and ( n9708 , n9196 , n7823 );
and ( n9709 , n9049 , n7821 );
nor ( n9710 , n9708 , n9709 );
xnor ( n9711 , n9710 , n7833 );
and ( n9712 , n9706 , n9711 );
and ( n9713 , n9693 , n9711 );
or ( n9714 , n9707 , n9712 , n9713 );
and ( n9715 , n7618 , n7542 );
and ( n9716 , n7666 , n7540 );
nor ( n9717 , n9715 , n9716 );
xnor ( n9718 , n9717 , n7552 );
and ( n9719 , n9714 , n9718 );
xor ( n9720 , n9455 , n9468 );
xor ( n9721 , n9720 , n9473 );
and ( n9722 , n9718 , n9721 );
and ( n9723 , n9714 , n9721 );
or ( n9724 , n9719 , n9722 , n9723 );
and ( n9725 , n7762 , n8168 );
and ( n9726 , n7786 , n8166 );
nor ( n9727 , n9725 , n9726 );
xnor ( n9728 , n9727 , n8178 );
and ( n9729 , n9724 , n9728 );
and ( n9730 , n7506 , n7899 );
and ( n9731 , n7945 , n7897 );
nor ( n9732 , n9730 , n9731 );
xnor ( n9733 , n9732 , n7909 );
and ( n9734 , n9728 , n9733 );
and ( n9735 , n9724 , n9733 );
or ( n9736 , n9729 , n9734 , n9735 );
xor ( n9737 , n9554 , n9568 );
xor ( n9738 , n9737 , n9573 );
and ( n9739 , n9736 , n9738 );
xor ( n9740 , n9434 , n9438 );
xor ( n9741 , n9740 , n9441 );
and ( n9742 , n9738 , n9741 );
and ( n9743 , n9736 , n9741 );
or ( n9744 , n9739 , n9742 , n9743 );
xor ( n9745 , n9444 , n9448 );
xor ( n9746 , n9745 , n9451 );
and ( n9747 , n9744 , n9746 );
xor ( n9748 , n9500 , n9514 );
xor ( n9749 , n9748 , n9517 );
and ( n9750 , n9746 , n9749 );
and ( n9751 , n9744 , n9749 );
or ( n9752 , n9747 , n9750 , n9751 );
and ( n9753 , n9692 , n9752 );
xor ( n9754 , n9416 , n9418 );
xor ( n9755 , n9754 , n9421 );
and ( n9756 , n9752 , n9755 );
and ( n9757 , n9692 , n9755 );
or ( n9758 , n9753 , n9756 , n9757 );
and ( n9759 , n7838 , n7601 );
and ( n9760 , n7676 , n7599 );
nor ( n9761 , n9759 , n9760 );
xnor ( n9762 , n9761 , n7611 );
and ( n9763 , n8066 , n7743 );
and ( n9764 , n7851 , n7741 );
nor ( n9765 , n9763 , n9764 );
xnor ( n9766 , n9765 , n7753 );
and ( n9767 , n9762 , n9766 );
and ( n9768 , n8263 , n7866 );
and ( n9769 , n8079 , n7864 );
nor ( n9770 , n9768 , n9769 );
xnor ( n9771 , n9770 , n7876 );
and ( n9772 , n9766 , n9771 );
and ( n9773 , n9762 , n9771 );
or ( n9774 , n9767 , n9772 , n9773 );
and ( n9775 , n7871 , n7501 );
and ( n9776 , n7800 , n7499 );
nor ( n9777 , n9775 , n9776 );
xnor ( n9778 , n9777 , n7511 );
and ( n9779 , n9774 , n9778 );
and ( n9780 , n7828 , n7713 );
and ( n9781 , n7809 , n7711 );
nor ( n9782 , n9780 , n9781 );
xnor ( n9783 , n9782 , n7723 );
and ( n9784 , n9778 , n9783 );
and ( n9785 , n9774 , n9783 );
or ( n9786 , n9779 , n9784 , n9785 );
and ( n9787 , n8035 , n7318 );
and ( n9788 , n8049 , n7315 );
nor ( n9789 , n9787 , n9788 );
xnor ( n9790 , n9789 , n7311 );
and ( n9791 , n9786 , n9790 );
xor ( n9792 , n9558 , n9562 );
xor ( n9793 , n9792 , n9565 );
and ( n9794 , n9790 , n9793 );
and ( n9795 , n9786 , n9793 );
or ( n9796 , n9791 , n9794 , n9795 );
xor ( n9797 , n9650 , n9654 );
xor ( n9798 , n9797 , n9659 );
and ( n9799 , n9796 , n9798 );
xor ( n9800 , n9504 , n9508 );
xor ( n9801 , n9800 , n9511 );
and ( n9802 , n9798 , n9801 );
and ( n9803 , n9796 , n9801 );
or ( n9804 , n9799 , n9802 , n9803 );
and ( n9805 , n7516 , n8044 );
and ( n9806 , n7547 , n8042 );
nor ( n9807 , n9805 , n9806 );
xnor ( n9808 , n9807 , n8054 );
and ( n9809 , n7704 , n7781 );
and ( n9810 , n7718 , n7779 );
nor ( n9811 , n9809 , n9810 );
xnor ( n9812 , n9811 , n7791 );
and ( n9813 , n9808 , n9812 );
and ( n9814 , n7729 , n7954 );
and ( n9815 , n7748 , n7952 );
nor ( n9816 , n9814 , n9815 );
xnor ( n9817 , n9816 , n7964 );
and ( n9818 , n9812 , n9817 );
and ( n9819 , n9808 , n9817 );
or ( n9820 , n9813 , n9818 , n9819 );
xor ( n9821 , n9697 , n9705 );
and ( n9822 , n9463 , n7823 );
and ( n9823 , n9280 , n7821 );
nor ( n9824 , n9822 , n9823 );
xnor ( n9825 , n9824 , n7833 );
xor ( n9826 , n7075 , n7245 );
buf ( n9827 , n9826 );
buf ( n9828 , n9827 );
buf ( n9829 , n9828 );
and ( n9830 , n9829 , n7691 );
and ( n9831 , n9701 , n7689 );
nor ( n9832 , n9830 , n9831 );
not ( n9833 , n9832 );
and ( n9834 , n9825 , n9833 );
and ( n9835 , n9821 , n9834 );
and ( n9836 , n9280 , n7823 );
and ( n9837 , n9196 , n7821 );
nor ( n9838 , n9836 , n9837 );
xnor ( n9839 , n9838 , n7833 );
and ( n9840 , n9834 , n9839 );
and ( n9841 , n9821 , n9839 );
or ( n9842 , n9835 , n9840 , n9841 );
and ( n9843 , n7666 , n7501 );
and ( n9844 , n7871 , n7499 );
nor ( n9845 , n9843 , n9844 );
xnor ( n9846 , n9845 , n7511 );
and ( n9847 , n9842 , n9846 );
and ( n9848 , n7696 , n7713 );
and ( n9849 , n7828 , n7711 );
nor ( n9850 , n9848 , n9849 );
xnor ( n9851 , n9850 , n7723 );
and ( n9852 , n9846 , n9851 );
and ( n9853 , n9842 , n9851 );
or ( n9854 , n9847 , n9852 , n9853 );
and ( n9855 , n7945 , n7395 );
and ( n9856 , n7959 , n7393 );
nor ( n9857 , n9855 , n9856 );
xnor ( n9858 , n9857 , n7405 );
and ( n9859 , n9854 , n9858 );
and ( n9860 , n7410 , n7899 );
and ( n9861 , n7506 , n7897 );
nor ( n9862 , n9860 , n9861 );
xnor ( n9863 , n9862 , n7909 );
and ( n9864 , n9858 , n9863 );
and ( n9865 , n9854 , n9863 );
or ( n9866 , n9859 , n9864 , n9865 );
and ( n9867 , n9820 , n9866 );
xor ( n9868 , n9542 , n9546 );
xor ( n9869 , n9868 , n9551 );
and ( n9870 , n9866 , n9869 );
and ( n9871 , n9820 , n9869 );
or ( n9872 , n9867 , n9870 , n9871 );
and ( n9873 , n7919 , n8168 );
and ( n9874 , n7762 , n8166 );
nor ( n9875 , n9873 , n9874 );
xnor ( n9876 , n9875 , n8178 );
and ( n9877 , n7558 , n7933 );
and ( n9878 , n7606 , n7931 );
nor ( n9879 , n9877 , n9878 );
xnor ( n9880 , n9879 , n7939 );
and ( n9881 , n9876 , n9880 );
xor ( n9882 , n9530 , n9534 );
xor ( n9883 , n9882 , n9539 );
and ( n9884 , n9880 , n9883 );
and ( n9885 , n9876 , n9883 );
or ( n9886 , n9881 , n9884 , n9885 );
xor ( n9887 , n9666 , n9670 );
xor ( n9888 , n9887 , n9675 );
and ( n9889 , n9886 , n9888 );
xor ( n9890 , n9640 , n9644 );
xor ( n9891 , n9890 , n9647 );
and ( n9892 , n9888 , n9891 );
and ( n9893 , n9886 , n9891 );
or ( n9894 , n9889 , n9892 , n9893 );
and ( n9895 , n9872 , n9894 );
xor ( n9896 , n9678 , n9680 );
xor ( n9897 , n9896 , n9683 );
and ( n9898 , n9894 , n9897 );
and ( n9899 , n9872 , n9897 );
or ( n9900 , n9895 , n9898 , n9899 );
and ( n9901 , n9804 , n9900 );
xor ( n9902 , n9576 , n9578 );
xor ( n9903 , n9902 , n9581 );
and ( n9904 , n9900 , n9903 );
and ( n9905 , n9804 , n9903 );
or ( n9906 , n9901 , n9904 , n9905 );
xor ( n9907 , n9454 , n9520 );
xor ( n9908 , n9907 , n9523 );
and ( n9909 , n9906 , n9908 );
xor ( n9910 , n9584 , n9586 );
xor ( n9911 , n9910 , n9589 );
and ( n9912 , n9908 , n9911 );
and ( n9913 , n9906 , n9911 );
or ( n9914 , n9909 , n9912 , n9913 );
and ( n9915 , n9758 , n9914 );
xor ( n9916 , n9617 , n9619 );
xor ( n9917 , n9916 , n9622 );
and ( n9918 , n9914 , n9917 );
and ( n9919 , n9758 , n9917 );
or ( n9920 , n9915 , n9918 , n9919 );
and ( n9921 , n9636 , n9920 );
xor ( n9922 , n9758 , n9914 );
xor ( n9923 , n9922 , n9917 );
xor ( n9924 , n9692 , n9752 );
xor ( n9925 , n9924 , n9755 );
xor ( n9926 , n9906 , n9908 );
xor ( n9927 , n9926 , n9911 );
and ( n9928 , n9925 , n9927 );
and ( n9929 , n9923 , n9928 );
xor ( n9930 , n9662 , n9686 );
xor ( n9931 , n9930 , n9689 );
xor ( n9932 , n9744 , n9746 );
xor ( n9933 , n9932 , n9749 );
and ( n9934 , n9931 , n9933 );
xor ( n9935 , n9804 , n9900 );
xor ( n9936 , n9935 , n9903 );
xor ( n9937 , n9931 , n9933 );
and ( n9938 , n9936 , n9937 );
xor ( n9939 , n9796 , n9798 );
xor ( n9940 , n9939 , n9801 );
xor ( n9941 , n9872 , n9894 );
xor ( n9942 , n9941 , n9897 );
and ( n9943 , n9940 , n9942 );
and ( n9944 , n9937 , n9943 );
and ( n9945 , n9936 , n9943 );
or ( n9946 , n9938 , n9944 , n9945 );
and ( n9947 , n9934 , n9946 );
xor ( n9948 , n9925 , n9927 );
and ( n9949 , n9946 , n9948 );
and ( n9950 , n9934 , n9948 );
or ( n9951 , n9947 , n9949 , n9950 );
and ( n9952 , n9928 , n9951 );
and ( n9953 , n9923 , n9951 );
or ( n9954 , n9929 , n9952 , n9953 );
and ( n9955 , n9920 , n9954 );
and ( n9956 , n9636 , n9954 );
or ( n9957 , n9921 , n9955 , n9956 );
and ( n9958 , n9633 , n9957 );
and ( n9959 , n9615 , n9957 );
or ( n9960 , n9634 , n9958 , n9959 );
and ( n9961 , n9612 , n9960 );
and ( n9962 , n9366 , n9960 );
or ( n9963 , n9613 , n9961 , n9962 );
and ( n9964 , n9364 , n9963 );
xor ( n9965 , n9364 , n9963 );
xor ( n9966 , n9366 , n9612 );
xor ( n9967 , n9966 , n9960 );
xor ( n9968 , n9615 , n9633 );
xor ( n9969 , n9968 , n9957 );
xor ( n9970 , n9636 , n9920 );
xor ( n9971 , n9970 , n9954 );
xor ( n9972 , n9923 , n9928 );
xor ( n9973 , n9972 , n9951 );
xor ( n9974 , n9736 , n9738 );
xor ( n9975 , n9974 , n9741 );
and ( n9976 , n7786 , n7318 );
and ( n9977 , n8035 , n7315 );
nor ( n9978 , n9976 , n9977 );
xnor ( n9979 , n9978 , n7311 );
xor ( n9980 , n9808 , n9812 );
xor ( n9981 , n9980 , n9817 );
and ( n9982 , n9979 , n9981 );
and ( n9983 , n7606 , n7781 );
and ( n9984 , n7704 , n7779 );
nor ( n9985 , n9983 , n9984 );
xnor ( n9986 , n9985 , n7791 );
and ( n9987 , n7748 , n7933 );
and ( n9988 , n7558 , n7931 );
nor ( n9989 , n9987 , n9988 );
xnor ( n9990 , n9989 , n7939 );
and ( n9991 , n9986 , n9990 );
and ( n9992 , n9981 , n9991 );
and ( n9993 , n9979 , n9991 );
or ( n9994 , n9982 , n9992 , n9993 );
xor ( n9995 , n9876 , n9880 );
xor ( n9996 , n9995 , n9883 );
and ( n9997 , n7959 , n8168 );
and ( n9998 , n7919 , n8166 );
nor ( n9999 , n9997 , n9998 );
xnor ( n10000 , n9999 , n8178 );
and ( n10001 , n7809 , n7542 );
and ( n10002 , n7618 , n7540 );
nor ( n10003 , n10001 , n10002 );
xnor ( n10004 , n10003 , n7552 );
and ( n10005 , n10000 , n10004 );
xor ( n10006 , n9762 , n9766 );
xor ( n10007 , n10006 , n9771 );
and ( n10008 , n10004 , n10007 );
and ( n10009 , n10000 , n10007 );
or ( n10010 , n10005 , n10008 , n10009 );
and ( n10011 , n9996 , n10010 );
xor ( n10012 , n9979 , n9981 );
xor ( n10013 , n10012 , n9991 );
and ( n10014 , n10010 , n10013 );
and ( n10015 , n9996 , n10013 );
or ( n10016 , n10011 , n10014 , n10015 );
and ( n10017 , n9994 , n10016 );
xor ( n10018 , n9786 , n9790 );
xor ( n10019 , n10018 , n9793 );
and ( n10020 , n10016 , n10019 );
and ( n10021 , n9994 , n10019 );
or ( n10022 , n10017 , n10020 , n10021 );
and ( n10023 , n9975 , n10022 );
xor ( n10024 , n9825 , n9833 );
and ( n10025 , n9701 , n7823 );
and ( n10026 , n9463 , n7821 );
nor ( n10027 , n10025 , n10026 );
xnor ( n10028 , n10027 , n7833 );
xor ( n10029 , n7077 , n7244 );
buf ( n10030 , n10029 );
buf ( n10031 , n10030 );
buf ( n10032 , n10031 );
and ( n10033 , n10032 , n7691 );
and ( n10034 , n9829 , n7689 );
nor ( n10035 , n10033 , n10034 );
not ( n10036 , n10035 );
and ( n10037 , n10028 , n10036 );
and ( n10038 , n10024 , n10037 );
and ( n10039 , n8696 , n7866 );
and ( n10040 , n8429 , n7864 );
nor ( n10041 , n10039 , n10040 );
xnor ( n10042 , n10041 , n7876 );
and ( n10043 , n10037 , n10042 );
and ( n10044 , n10024 , n10042 );
or ( n10045 , n10038 , n10043 , n10044 );
and ( n10046 , n8079 , n7743 );
and ( n10047 , n8066 , n7741 );
nor ( n10048 , n10046 , n10047 );
xnor ( n10049 , n10048 , n7753 );
and ( n10050 , n10045 , n10049 );
and ( n10051 , n8429 , n7866 );
and ( n10052 , n8263 , n7864 );
nor ( n10053 , n10051 , n10052 );
xnor ( n10054 , n10053 , n7876 );
and ( n10055 , n10049 , n10054 );
and ( n10056 , n10045 , n10054 );
or ( n10057 , n10050 , n10055 , n10056 );
and ( n10058 , n7800 , n7954 );
and ( n10059 , n7729 , n7952 );
nor ( n10060 , n10058 , n10059 );
xnor ( n10061 , n10060 , n7964 );
and ( n10062 , n10057 , n10061 );
xor ( n10063 , n9693 , n9706 );
xor ( n10064 , n10063 , n9711 );
and ( n10065 , n10061 , n10064 );
and ( n10066 , n10057 , n10064 );
or ( n10067 , n10062 , n10065 , n10066 );
xor ( n10068 , n9774 , n9778 );
xor ( n10069 , n10068 , n9783 );
and ( n10070 , n10067 , n10069 );
xor ( n10071 , n9714 , n9718 );
xor ( n10072 , n10071 , n9721 );
and ( n10073 , n10069 , n10072 );
and ( n10074 , n10067 , n10072 );
or ( n10075 , n10070 , n10073 , n10074 );
xor ( n10076 , n9724 , n9728 );
xor ( n10077 , n10076 , n9733 );
and ( n10078 , n10075 , n10077 );
and ( n10079 , n10022 , n10078 );
and ( n10080 , n9975 , n10078 );
or ( n10081 , n10023 , n10079 , n10080 );
and ( n10082 , n8066 , n7601 );
and ( n10083 , n7851 , n7599 );
nor ( n10084 , n10082 , n10083 );
xnor ( n10085 , n10084 , n7611 );
and ( n10086 , n8263 , n7743 );
and ( n10087 , n8079 , n7741 );
nor ( n10088 , n10086 , n10087 );
xnor ( n10089 , n10088 , n7753 );
and ( n10090 , n10085 , n10089 );
and ( n10091 , n9196 , n7661 );
and ( n10092 , n9049 , n7659 );
nor ( n10093 , n10091 , n10092 );
xnor ( n10094 , n10093 , n7671 );
and ( n10095 , n10089 , n10094 );
and ( n10096 , n10085 , n10094 );
or ( n10097 , n10090 , n10095 , n10096 );
and ( n10098 , n7676 , n7713 );
and ( n10099 , n7696 , n7711 );
nor ( n10100 , n10098 , n10099 );
xnor ( n10101 , n10100 , n7723 );
and ( n10102 , n10097 , n10101 );
and ( n10103 , n7851 , n7601 );
and ( n10104 , n7838 , n7599 );
nor ( n10105 , n10103 , n10104 );
xnor ( n10106 , n10105 , n7611 );
and ( n10107 , n10101 , n10106 );
and ( n10108 , n10097 , n10106 );
or ( n10109 , n10102 , n10107 , n10108 );
and ( n10110 , n7547 , n7899 );
and ( n10111 , n7410 , n7897 );
nor ( n10112 , n10110 , n10111 );
xnor ( n10113 , n10112 , n7909 );
and ( n10114 , n10109 , n10113 );
and ( n10115 , n7718 , n8044 );
and ( n10116 , n7516 , n8042 );
nor ( n10117 , n10115 , n10116 );
xnor ( n10118 , n10117 , n8054 );
and ( n10119 , n10113 , n10118 );
and ( n10120 , n10109 , n10118 );
or ( n10121 , n10114 , n10119 , n10120 );
and ( n10122 , n7762 , n7318 );
and ( n10123 , n7786 , n7315 );
nor ( n10124 , n10122 , n10123 );
xnor ( n10125 , n10124 , n7311 );
xor ( n10126 , n9986 , n9990 );
and ( n10127 , n10125 , n10126 );
xor ( n10128 , n10000 , n10004 );
xor ( n10129 , n10128 , n10007 );
and ( n10130 , n10126 , n10129 );
and ( n10131 , n10125 , n10129 );
or ( n10132 , n10127 , n10130 , n10131 );
and ( n10133 , n10121 , n10132 );
xor ( n10134 , n9996 , n10010 );
xor ( n10135 , n10134 , n10013 );
and ( n10136 , n10132 , n10135 );
and ( n10137 , n10121 , n10135 );
or ( n10138 , n10133 , n10136 , n10137 );
xor ( n10139 , n9820 , n9866 );
xor ( n10140 , n10139 , n9869 );
and ( n10141 , n10138 , n10140 );
xor ( n10142 , n9994 , n10016 );
xor ( n10143 , n10142 , n10019 );
and ( n10144 , n10140 , n10143 );
and ( n10145 , n10138 , n10143 );
or ( n10146 , n10141 , n10144 , n10145 );
xor ( n10147 , n9940 , n9942 );
and ( n10148 , n10146 , n10147 );
and ( n10149 , n7618 , n7501 );
and ( n10150 , n7666 , n7499 );
nor ( n10151 , n10149 , n10150 );
xnor ( n10152 , n10151 , n7511 );
xor ( n10153 , n10045 , n10049 );
xor ( n10154 , n10153 , n10054 );
and ( n10155 , n10152 , n10154 );
xor ( n10156 , n9821 , n9834 );
xor ( n10157 , n10156 , n9839 );
and ( n10158 , n10154 , n10157 );
and ( n10159 , n10152 , n10157 );
or ( n10160 , n10155 , n10158 , n10159 );
and ( n10161 , n7506 , n7395 );
and ( n10162 , n7945 , n7393 );
nor ( n10163 , n10161 , n10162 );
xnor ( n10164 , n10163 , n7405 );
and ( n10165 , n10160 , n10164 );
xor ( n10166 , n9842 , n9846 );
xor ( n10167 , n10166 , n9851 );
and ( n10168 , n10164 , n10167 );
and ( n10169 , n10160 , n10167 );
or ( n10170 , n10165 , n10168 , n10169 );
xor ( n10171 , n9854 , n9858 );
xor ( n10172 , n10171 , n9863 );
and ( n10173 , n10170 , n10172 );
xor ( n10174 , n10067 , n10069 );
xor ( n10175 , n10174 , n10072 );
and ( n10176 , n10172 , n10175 );
and ( n10177 , n10170 , n10175 );
or ( n10178 , n10173 , n10176 , n10177 );
xor ( n10179 , n9886 , n9888 );
xor ( n10180 , n10179 , n9891 );
and ( n10181 , n10178 , n10180 );
and ( n10182 , n10147 , n10181 );
and ( n10183 , n10146 , n10181 );
or ( n10184 , n10148 , n10182 , n10183 );
and ( n10185 , n10081 , n10184 );
xor ( n10186 , n9936 , n9937 );
xor ( n10187 , n10186 , n9943 );
and ( n10188 , n10184 , n10187 );
and ( n10189 , n10081 , n10187 );
or ( n10190 , n10185 , n10188 , n10189 );
xor ( n10191 , n9934 , n9946 );
xor ( n10192 , n10191 , n9948 );
and ( n10193 , n10190 , n10192 );
xor ( n10194 , n9975 , n10022 );
xor ( n10195 , n10194 , n10078 );
xor ( n10196 , n10075 , n10077 );
xor ( n10197 , n10138 , n10140 );
xor ( n10198 , n10197 , n10143 );
and ( n10199 , n10196 , n10198 );
xor ( n10200 , n10178 , n10180 );
and ( n10201 , n10198 , n10200 );
and ( n10202 , n10196 , n10200 );
or ( n10203 , n10199 , n10201 , n10202 );
and ( n10204 , n10195 , n10203 );
xor ( n10205 , n10146 , n10147 );
xor ( n10206 , n10205 , n10181 );
and ( n10207 , n10203 , n10206 );
and ( n10208 , n10195 , n10206 );
or ( n10209 , n10204 , n10207 , n10208 );
xor ( n10210 , n10081 , n10184 );
xor ( n10211 , n10210 , n10187 );
and ( n10212 , n10209 , n10211 );
xor ( n10213 , n10121 , n10132 );
xor ( n10214 , n10213 , n10135 );
and ( n10215 , n7516 , n7899 );
and ( n10216 , n7547 , n7897 );
nor ( n10217 , n10215 , n10216 );
xnor ( n10218 , n10217 , n7909 );
and ( n10219 , n7704 , n8044 );
and ( n10220 , n7718 , n8042 );
nor ( n10221 , n10219 , n10220 );
xnor ( n10222 , n10221 , n8054 );
and ( n10223 , n10218 , n10222 );
and ( n10224 , n7558 , n7781 );
and ( n10225 , n7606 , n7779 );
nor ( n10226 , n10224 , n10225 );
xnor ( n10227 , n10226 , n7791 );
and ( n10228 , n10222 , n10227 );
and ( n10229 , n10218 , n10227 );
or ( n10230 , n10223 , n10228 , n10229 );
xor ( n10231 , n10028 , n10036 );
and ( n10232 , n9463 , n7661 );
and ( n10233 , n9280 , n7659 );
nor ( n10234 , n10232 , n10233 );
xnor ( n10235 , n10234 , n7671 );
xor ( n10236 , n7079 , n7243 );
buf ( n10237 , n10236 );
buf ( n10238 , n10237 );
buf ( n10239 , n10238 );
and ( n10240 , n10239 , n7691 );
and ( n10241 , n10032 , n7689 );
nor ( n10242 , n10240 , n10241 );
not ( n10243 , n10242 );
and ( n10244 , n10235 , n10243 );
and ( n10245 , n10231 , n10244 );
and ( n10246 , n9049 , n7866 );
and ( n10247 , n8696 , n7864 );
nor ( n10248 , n10246 , n10247 );
xnor ( n10249 , n10248 , n7876 );
and ( n10250 , n10244 , n10249 );
and ( n10251 , n10231 , n10249 );
or ( n10252 , n10245 , n10250 , n10251 );
and ( n10253 , n7838 , n7713 );
and ( n10254 , n7676 , n7711 );
nor ( n10255 , n10253 , n10254 );
xnor ( n10256 , n10255 , n7723 );
and ( n10257 , n10252 , n10256 );
xor ( n10258 , n10024 , n10037 );
xor ( n10259 , n10258 , n10042 );
and ( n10260 , n10256 , n10259 );
and ( n10261 , n10252 , n10259 );
or ( n10262 , n10257 , n10260 , n10261 );
and ( n10263 , n7871 , n7954 );
and ( n10264 , n7800 , n7952 );
nor ( n10265 , n10263 , n10264 );
xnor ( n10266 , n10265 , n7964 );
and ( n10267 , n10262 , n10266 );
and ( n10268 , n7828 , n7542 );
and ( n10269 , n7809 , n7540 );
nor ( n10270 , n10268 , n10269 );
xnor ( n10271 , n10270 , n7552 );
and ( n10272 , n10266 , n10271 );
and ( n10273 , n10262 , n10271 );
or ( n10274 , n10267 , n10272 , n10273 );
and ( n10275 , n10230 , n10274 );
xor ( n10276 , n10057 , n10061 );
xor ( n10277 , n10276 , n10064 );
and ( n10278 , n10274 , n10277 );
and ( n10279 , n10230 , n10277 );
or ( n10280 , n10275 , n10278 , n10279 );
and ( n10281 , n10214 , n10280 );
xor ( n10282 , n10170 , n10172 );
xor ( n10283 , n10282 , n10175 );
and ( n10284 , n10280 , n10283 );
and ( n10285 , n10214 , n10283 );
or ( n10286 , n10281 , n10284 , n10285 );
and ( n10287 , n8079 , n7601 );
and ( n10288 , n8066 , n7599 );
nor ( n10289 , n10287 , n10288 );
xnor ( n10290 , n10289 , n7611 );
and ( n10291 , n8429 , n7743 );
and ( n10292 , n8263 , n7741 );
nor ( n10293 , n10291 , n10292 );
xnor ( n10294 , n10293 , n7753 );
and ( n10295 , n10290 , n10294 );
and ( n10296 , n9280 , n7661 );
and ( n10297 , n9196 , n7659 );
nor ( n10298 , n10296 , n10297 );
xnor ( n10299 , n10298 , n7671 );
and ( n10300 , n10294 , n10299 );
and ( n10301 , n10290 , n10299 );
or ( n10302 , n10295 , n10300 , n10301 );
and ( n10303 , n7666 , n7954 );
and ( n10304 , n7871 , n7952 );
nor ( n10305 , n10303 , n10304 );
xnor ( n10306 , n10305 , n7964 );
and ( n10307 , n10302 , n10306 );
and ( n10308 , n7696 , n7542 );
and ( n10309 , n7828 , n7540 );
nor ( n10310 , n10308 , n10309 );
xnor ( n10311 , n10310 , n7552 );
and ( n10312 , n10306 , n10311 );
and ( n10313 , n10302 , n10311 );
or ( n10314 , n10307 , n10312 , n10313 );
and ( n10315 , n7919 , n7318 );
and ( n10316 , n7762 , n7315 );
nor ( n10317 , n10315 , n10316 );
xnor ( n10318 , n10317 , n7311 );
and ( n10319 , n10314 , n10318 );
and ( n10320 , n7410 , n7395 );
and ( n10321 , n7506 , n7393 );
nor ( n10322 , n10320 , n10321 );
xnor ( n10323 , n10322 , n7405 );
and ( n10324 , n10318 , n10323 );
and ( n10325 , n10314 , n10323 );
or ( n10326 , n10319 , n10324 , n10325 );
xor ( n10327 , n10109 , n10113 );
xor ( n10328 , n10327 , n10118 );
and ( n10329 , n10326 , n10328 );
xor ( n10330 , n10160 , n10164 );
xor ( n10331 , n10330 , n10167 );
and ( n10332 , n10328 , n10331 );
and ( n10333 , n10326 , n10331 );
or ( n10334 , n10329 , n10332 , n10333 );
and ( n10335 , n7959 , n7318 );
and ( n10336 , n7919 , n7315 );
nor ( n10337 , n10335 , n10336 );
xnor ( n10338 , n10337 , n7311 );
and ( n10339 , n7606 , n8044 );
and ( n10340 , n7704 , n8042 );
nor ( n10341 , n10339 , n10340 );
xnor ( n10342 , n10341 , n8054 );
and ( n10343 , n10338 , n10342 );
and ( n10344 , n7748 , n7781 );
and ( n10345 , n7558 , n7779 );
nor ( n10346 , n10344 , n10345 );
xnor ( n10347 , n10346 , n7791 );
and ( n10348 , n10342 , n10347 );
and ( n10349 , n10338 , n10347 );
or ( n10350 , n10343 , n10348 , n10349 );
xor ( n10351 , n10262 , n10266 );
xor ( n10352 , n10351 , n10271 );
and ( n10353 , n10350 , n10352 );
and ( n10354 , n7945 , n8168 );
and ( n10355 , n7959 , n8166 );
nor ( n10356 , n10354 , n10355 );
xnor ( n10357 , n10356 , n8178 );
and ( n10358 , n7729 , n7933 );
and ( n10359 , n7748 , n7931 );
nor ( n10360 , n10358 , n10359 );
xnor ( n10361 , n10360 , n7939 );
xor ( n10362 , n10357 , n10361 );
xor ( n10363 , n10097 , n10101 );
xor ( n10364 , n10363 , n10106 );
xor ( n10365 , n10362 , n10364 );
and ( n10366 , n10352 , n10365 );
and ( n10367 , n10350 , n10365 );
or ( n10368 , n10353 , n10366 , n10367 );
xor ( n10369 , n10235 , n10243 );
and ( n10370 , n9701 , n7661 );
and ( n10371 , n9463 , n7659 );
nor ( n10372 , n10370 , n10371 );
xnor ( n10373 , n10372 , n7671 );
xor ( n10374 , n7081 , n7242 );
buf ( n10375 , n10374 );
buf ( n10376 , n10375 );
buf ( n10377 , n10376 );
and ( n10378 , n10377 , n7691 );
and ( n10379 , n10239 , n7689 );
nor ( n10380 , n10378 , n10379 );
not ( n10381 , n10380 );
and ( n10382 , n10373 , n10381 );
and ( n10383 , n10369 , n10382 );
and ( n10384 , n9829 , n7823 );
and ( n10385 , n9701 , n7821 );
nor ( n10386 , n10384 , n10385 );
xnor ( n10387 , n10386 , n7833 );
and ( n10388 , n10382 , n10387 );
and ( n10389 , n10369 , n10387 );
or ( n10390 , n10383 , n10388 , n10389 );
and ( n10391 , n7676 , n7542 );
and ( n10392 , n7696 , n7540 );
nor ( n10393 , n10391 , n10392 );
xnor ( n10394 , n10393 , n7552 );
and ( n10395 , n10390 , n10394 );
and ( n10396 , n7851 , n7713 );
and ( n10397 , n7838 , n7711 );
nor ( n10398 , n10396 , n10397 );
xnor ( n10399 , n10398 , n7723 );
and ( n10400 , n10394 , n10399 );
and ( n10401 , n10390 , n10399 );
or ( n10402 , n10395 , n10400 , n10401 );
and ( n10403 , n7809 , n7501 );
and ( n10404 , n7618 , n7499 );
nor ( n10405 , n10403 , n10404 );
xnor ( n10406 , n10405 , n7511 );
and ( n10407 , n10402 , n10406 );
xor ( n10408 , n10085 , n10089 );
xor ( n10409 , n10408 , n10094 );
and ( n10410 , n10406 , n10409 );
and ( n10411 , n10402 , n10409 );
or ( n10412 , n10407 , n10410 , n10411 );
and ( n10413 , n7718 , n7899 );
and ( n10414 , n7516 , n7897 );
nor ( n10415 , n10413 , n10414 );
xnor ( n10416 , n10415 , n7909 );
and ( n10417 , n7800 , n7933 );
and ( n10418 , n7729 , n7931 );
nor ( n10419 , n10417 , n10418 );
xnor ( n10420 , n10419 , n7939 );
and ( n10421 , n10416 , n10420 );
xor ( n10422 , n10252 , n10256 );
xor ( n10423 , n10422 , n10259 );
and ( n10424 , n10420 , n10423 );
and ( n10425 , n10416 , n10423 );
or ( n10426 , n10421 , n10424 , n10425 );
and ( n10427 , n10412 , n10426 );
xor ( n10428 , n10152 , n10154 );
xor ( n10429 , n10428 , n10157 );
and ( n10430 , n10426 , n10429 );
and ( n10431 , n10412 , n10429 );
or ( n10432 , n10427 , n10430 , n10431 );
and ( n10433 , n10368 , n10432 );
xor ( n10434 , n10230 , n10274 );
xor ( n10435 , n10434 , n10277 );
and ( n10436 , n10432 , n10435 );
and ( n10437 , n10368 , n10435 );
or ( n10438 , n10433 , n10436 , n10437 );
and ( n10439 , n10334 , n10438 );
and ( n10440 , n8263 , n7601 );
and ( n10441 , n8079 , n7599 );
nor ( n10442 , n10440 , n10441 );
xnor ( n10443 , n10442 , n7611 );
and ( n10444 , n8696 , n7743 );
and ( n10445 , n8429 , n7741 );
nor ( n10446 , n10444 , n10445 );
xnor ( n10447 , n10446 , n7753 );
and ( n10448 , n10443 , n10447 );
and ( n10449 , n9196 , n7866 );
and ( n10450 , n9049 , n7864 );
nor ( n10451 , n10449 , n10450 );
xnor ( n10452 , n10451 , n7876 );
and ( n10453 , n10447 , n10452 );
and ( n10454 , n10443 , n10452 );
or ( n10455 , n10448 , n10453 , n10454 );
and ( n10456 , n7618 , n7954 );
and ( n10457 , n7666 , n7952 );
nor ( n10458 , n10456 , n10457 );
xnor ( n10459 , n10458 , n7964 );
and ( n10460 , n10455 , n10459 );
xor ( n10461 , n10231 , n10244 );
xor ( n10462 , n10461 , n10249 );
and ( n10463 , n10459 , n10462 );
and ( n10464 , n10455 , n10462 );
or ( n10465 , n10460 , n10463 , n10464 );
and ( n10466 , n7506 , n8168 );
and ( n10467 , n7945 , n8166 );
nor ( n10468 , n10466 , n10467 );
xnor ( n10469 , n10468 , n8178 );
and ( n10470 , n10465 , n10469 );
and ( n10471 , n7547 , n7395 );
and ( n10472 , n7410 , n7393 );
nor ( n10473 , n10471 , n10472 );
xnor ( n10474 , n10473 , n7405 );
and ( n10475 , n10469 , n10474 );
and ( n10476 , n10465 , n10474 );
or ( n10477 , n10470 , n10475 , n10476 );
xor ( n10478 , n10218 , n10222 );
xor ( n10479 , n10478 , n10227 );
and ( n10480 , n10477 , n10479 );
xor ( n10481 , n10314 , n10318 );
xor ( n10482 , n10481 , n10323 );
and ( n10483 , n10479 , n10482 );
and ( n10484 , n10477 , n10482 );
or ( n10485 , n10480 , n10483 , n10484 );
xor ( n10486 , n10326 , n10328 );
xor ( n10487 , n10486 , n10331 );
and ( n10488 , n10485 , n10487 );
and ( n10489 , n10438 , n10488 );
and ( n10490 , n10334 , n10488 );
or ( n10491 , n10439 , n10489 , n10490 );
and ( n10492 , n10286 , n10491 );
xor ( n10493 , n10196 , n10198 );
xor ( n10494 , n10493 , n10200 );
and ( n10495 , n10491 , n10494 );
and ( n10496 , n10286 , n10494 );
or ( n10497 , n10492 , n10495 , n10496 );
xor ( n10498 , n10195 , n10203 );
xor ( n10499 , n10498 , n10206 );
and ( n10500 , n10497 , n10499 );
xor ( n10501 , n10214 , n10280 );
xor ( n10502 , n10501 , n10283 );
and ( n10503 , n7410 , n8168 );
and ( n10504 , n7506 , n8166 );
nor ( n10505 , n10503 , n10504 );
xnor ( n10506 , n10505 , n8178 );
xor ( n10507 , n10390 , n10394 );
xor ( n10508 , n10507 , n10399 );
and ( n10509 , n10506 , n10508 );
xor ( n10510 , n10455 , n10459 );
xor ( n10511 , n10510 , n10462 );
and ( n10512 , n10508 , n10511 );
and ( n10513 , n10506 , n10511 );
or ( n10514 , n10509 , n10512 , n10513 );
xor ( n10515 , n10465 , n10469 );
xor ( n10516 , n10515 , n10474 );
and ( n10517 , n10514 , n10516 );
xor ( n10518 , n10416 , n10420 );
xor ( n10519 , n10518 , n10423 );
and ( n10520 , n10516 , n10519 );
and ( n10521 , n10514 , n10519 );
or ( n10522 , n10517 , n10520 , n10521 );
xor ( n10523 , n10477 , n10479 );
xor ( n10524 , n10523 , n10482 );
and ( n10525 , n10522 , n10524 );
xor ( n10526 , n10350 , n10352 );
xor ( n10527 , n10526 , n10365 );
and ( n10528 , n10524 , n10527 );
and ( n10529 , n10522 , n10527 );
or ( n10530 , n10525 , n10528 , n10529 );
and ( n10531 , n7704 , n7899 );
and ( n10532 , n7718 , n7897 );
nor ( n10533 , n10531 , n10532 );
xnor ( n10534 , n10533 , n7909 );
and ( n10535 , n7558 , n8044 );
and ( n10536 , n7606 , n8042 );
nor ( n10537 , n10535 , n10536 );
xnor ( n10538 , n10537 , n8054 );
and ( n10539 , n10534 , n10538 );
and ( n10540 , n7871 , n7933 );
and ( n10541 , n7800 , n7931 );
nor ( n10542 , n10540 , n10541 );
xnor ( n10543 , n10542 , n7939 );
and ( n10544 , n10538 , n10543 );
and ( n10545 , n10534 , n10543 );
or ( n10546 , n10539 , n10544 , n10545 );
and ( n10547 , n10377 , n7823 );
and ( n10548 , n10239 , n7821 );
nor ( n10549 , n10547 , n10548 );
xnor ( n10550 , n10549 , n7833 );
xor ( n10551 , n7085 , n7240 );
buf ( n10552 , n10551 );
buf ( n10553 , n10552 );
buf ( n10554 , n10553 );
and ( n10555 , n10554 , n7691 );
xor ( n10556 , n7083 , n7241 );
buf ( n10557 , n10556 );
buf ( n10558 , n10557 );
buf ( n10559 , n10558 );
and ( n10560 , n10559 , n7689 );
nor ( n10561 , n10555 , n10560 );
not ( n10562 , n10561 );
and ( n10563 , n10550 , n10562 );
and ( n10564 , n9463 , n7866 );
and ( n10565 , n9280 , n7864 );
nor ( n10566 , n10564 , n10565 );
xnor ( n10567 , n10566 , n7876 );
and ( n10568 , n10563 , n10567 );
and ( n10569 , n9829 , n7661 );
and ( n10570 , n9701 , n7659 );
nor ( n10571 , n10569 , n10570 );
xnor ( n10572 , n10571 , n7671 );
and ( n10573 , n10567 , n10572 );
and ( n10574 , n10563 , n10572 );
or ( n10575 , n10568 , n10573 , n10574 );
and ( n10576 , n9049 , n7743 );
and ( n10577 , n8696 , n7741 );
nor ( n10578 , n10576 , n10577 );
xnor ( n10579 , n10578 , n7753 );
and ( n10580 , n10575 , n10579 );
and ( n10581 , n9280 , n7866 );
and ( n10582 , n9196 , n7864 );
nor ( n10583 , n10581 , n10582 );
xnor ( n10584 , n10583 , n7876 );
and ( n10585 , n10579 , n10584 );
and ( n10586 , n10575 , n10584 );
or ( n10587 , n10580 , n10585 , n10586 );
and ( n10588 , n7696 , n7501 );
and ( n10589 , n7828 , n7499 );
nor ( n10590 , n10588 , n10589 );
xnor ( n10591 , n10590 , n7511 );
and ( n10592 , n10587 , n10591 );
xor ( n10593 , n10369 , n10382 );
xor ( n10594 , n10593 , n10387 );
and ( n10595 , n10591 , n10594 );
and ( n10596 , n10587 , n10594 );
or ( n10597 , n10592 , n10595 , n10596 );
and ( n10598 , n7516 , n7395 );
and ( n10599 , n7547 , n7393 );
nor ( n10600 , n10598 , n10599 );
xnor ( n10601 , n10600 , n7405 );
and ( n10602 , n10597 , n10601 );
and ( n10603 , n7729 , n7781 );
and ( n10604 , n7748 , n7779 );
nor ( n10605 , n10603 , n10604 );
xnor ( n10606 , n10605 , n7791 );
and ( n10607 , n10601 , n10606 );
and ( n10608 , n10597 , n10606 );
or ( n10609 , n10602 , n10607 , n10608 );
and ( n10610 , n10546 , n10609 );
xor ( n10611 , n10338 , n10342 );
xor ( n10612 , n10611 , n10347 );
and ( n10613 , n10609 , n10612 );
and ( n10614 , n10546 , n10612 );
or ( n10615 , n10610 , n10613 , n10614 );
xor ( n10616 , n10373 , n10381 );
and ( n10617 , n10239 , n7823 );
and ( n10618 , n10032 , n7821 );
nor ( n10619 , n10617 , n10618 );
xnor ( n10620 , n10619 , n7833 );
and ( n10621 , n10559 , n7691 );
and ( n10622 , n10377 , n7689 );
nor ( n10623 , n10621 , n10622 );
not ( n10624 , n10623 );
and ( n10625 , n10620 , n10624 );
and ( n10626 , n10616 , n10625 );
and ( n10627 , n10032 , n7823 );
and ( n10628 , n9829 , n7821 );
nor ( n10629 , n10627 , n10628 );
xnor ( n10630 , n10629 , n7833 );
and ( n10631 , n10625 , n10630 );
and ( n10632 , n10616 , n10630 );
or ( n10633 , n10626 , n10631 , n10632 );
and ( n10634 , n7838 , n7542 );
and ( n10635 , n7676 , n7540 );
nor ( n10636 , n10634 , n10635 );
xnor ( n10637 , n10636 , n7552 );
and ( n10638 , n10633 , n10637 );
and ( n10639 , n8066 , n7713 );
and ( n10640 , n7851 , n7711 );
nor ( n10641 , n10639 , n10640 );
xnor ( n10642 , n10641 , n7723 );
and ( n10643 , n10637 , n10642 );
and ( n10644 , n10633 , n10642 );
or ( n10645 , n10638 , n10643 , n10644 );
and ( n10646 , n7828 , n7501 );
and ( n10647 , n7809 , n7499 );
nor ( n10648 , n10646 , n10647 );
xnor ( n10649 , n10648 , n7511 );
and ( n10650 , n10645 , n10649 );
xor ( n10651 , n10290 , n10294 );
xor ( n10652 , n10651 , n10299 );
and ( n10653 , n10649 , n10652 );
and ( n10654 , n10645 , n10652 );
or ( n10655 , n10650 , n10653 , n10654 );
xor ( n10656 , n10302 , n10306 );
xor ( n10657 , n10656 , n10311 );
and ( n10658 , n10655 , n10657 );
xor ( n10659 , n10402 , n10406 );
xor ( n10660 , n10659 , n10409 );
and ( n10661 , n10657 , n10660 );
and ( n10662 , n10655 , n10660 );
or ( n10663 , n10658 , n10661 , n10662 );
and ( n10664 , n10615 , n10663 );
xor ( n10665 , n10412 , n10426 );
xor ( n10666 , n10665 , n10429 );
and ( n10667 , n10663 , n10666 );
and ( n10668 , n10615 , n10666 );
or ( n10669 , n10664 , n10667 , n10668 );
and ( n10670 , n10530 , n10669 );
xor ( n10671 , n10368 , n10432 );
xor ( n10672 , n10671 , n10435 );
and ( n10673 , n10669 , n10672 );
and ( n10674 , n10530 , n10672 );
or ( n10675 , n10670 , n10673 , n10674 );
and ( n10676 , n10502 , n10675 );
and ( n10677 , n10357 , n10361 );
and ( n10678 , n10361 , n10364 );
and ( n10679 , n10357 , n10364 );
or ( n10680 , n10677 , n10678 , n10679 );
xor ( n10681 , n10125 , n10126 );
xor ( n10682 , n10681 , n10129 );
and ( n10683 , n10680 , n10682 );
xor ( n10684 , n10485 , n10487 );
and ( n10685 , n10682 , n10684 );
and ( n10686 , n10680 , n10684 );
or ( n10687 , n10683 , n10685 , n10686 );
and ( n10688 , n10675 , n10687 );
and ( n10689 , n10502 , n10687 );
or ( n10690 , n10676 , n10688 , n10689 );
xor ( n10691 , n10286 , n10491 );
xor ( n10692 , n10691 , n10494 );
and ( n10693 , n10690 , n10692 );
xor ( n10694 , n10334 , n10438 );
xor ( n10695 , n10694 , n10488 );
xor ( n10696 , n10530 , n10669 );
xor ( n10697 , n10696 , n10672 );
and ( n10698 , n7676 , n7501 );
and ( n10699 , n7696 , n7499 );
nor ( n10700 , n10698 , n10699 );
xnor ( n10701 , n10700 , n7511 );
and ( n10702 , n7851 , n7542 );
and ( n10703 , n7838 , n7540 );
nor ( n10704 , n10702 , n10703 );
xnor ( n10705 , n10704 , n7552 );
and ( n10706 , n10701 , n10705 );
xor ( n10707 , n10616 , n10625 );
xor ( n10708 , n10707 , n10630 );
and ( n10709 , n10705 , n10708 );
and ( n10710 , n10701 , n10708 );
or ( n10711 , n10706 , n10709 , n10710 );
and ( n10712 , n7800 , n7781 );
and ( n10713 , n7729 , n7779 );
nor ( n10714 , n10712 , n10713 );
xnor ( n10715 , n10714 , n7791 );
and ( n10716 , n10711 , n10715 );
and ( n10717 , n7809 , n7954 );
and ( n10718 , n7618 , n7952 );
nor ( n10719 , n10717 , n10718 );
xnor ( n10720 , n10719 , n7964 );
and ( n10721 , n10715 , n10720 );
and ( n10722 , n10711 , n10720 );
or ( n10723 , n10716 , n10721 , n10722 );
xor ( n10724 , n10620 , n10624 );
and ( n10725 , n8696 , n7601 );
and ( n10726 , n8429 , n7599 );
nor ( n10727 , n10725 , n10726 );
xnor ( n10728 , n10727 , n7611 );
and ( n10729 , n10724 , n10728 );
and ( n10730 , n9196 , n7743 );
and ( n10731 , n9049 , n7741 );
nor ( n10732 , n10730 , n10731 );
xnor ( n10733 , n10732 , n7753 );
and ( n10734 , n10728 , n10733 );
and ( n10735 , n10724 , n10733 );
or ( n10736 , n10729 , n10734 , n10735 );
and ( n10737 , n8079 , n7713 );
and ( n10738 , n8066 , n7711 );
nor ( n10739 , n10737 , n10738 );
xnor ( n10740 , n10739 , n7723 );
and ( n10741 , n10736 , n10740 );
and ( n10742 , n8429 , n7601 );
and ( n10743 , n8263 , n7599 );
nor ( n10744 , n10742 , n10743 );
xnor ( n10745 , n10744 , n7611 );
and ( n10746 , n10740 , n10745 );
and ( n10747 , n10736 , n10745 );
or ( n10748 , n10741 , n10746 , n10747 );
and ( n10749 , n7666 , n7933 );
and ( n10750 , n7871 , n7931 );
nor ( n10751 , n10749 , n10750 );
xnor ( n10752 , n10751 , n7939 );
and ( n10753 , n10748 , n10752 );
xor ( n10754 , n10443 , n10447 );
xor ( n10755 , n10754 , n10452 );
and ( n10756 , n10752 , n10755 );
and ( n10757 , n10748 , n10755 );
or ( n10758 , n10753 , n10756 , n10757 );
and ( n10759 , n10723 , n10758 );
and ( n10760 , n7945 , n7318 );
and ( n10761 , n7959 , n7315 );
nor ( n10762 , n10760 , n10761 );
xnor ( n10763 , n10762 , n7311 );
and ( n10764 , n10758 , n10763 );
and ( n10765 , n10723 , n10763 );
or ( n10766 , n10759 , n10764 , n10765 );
and ( n10767 , n7606 , n7899 );
and ( n10768 , n7704 , n7897 );
nor ( n10769 , n10767 , n10768 );
xnor ( n10770 , n10769 , n7909 );
and ( n10771 , n7748 , n8044 );
and ( n10772 , n7558 , n8042 );
nor ( n10773 , n10771 , n10772 );
xnor ( n10774 , n10773 , n8054 );
and ( n10775 , n10770 , n10774 );
xor ( n10776 , n10633 , n10637 );
xor ( n10777 , n10776 , n10642 );
and ( n10778 , n10774 , n10777 );
and ( n10779 , n10770 , n10777 );
or ( n10780 , n10775 , n10778 , n10779 );
xor ( n10781 , n10534 , n10538 );
xor ( n10782 , n10781 , n10543 );
and ( n10783 , n10780 , n10782 );
xor ( n10784 , n10645 , n10649 );
xor ( n10785 , n10784 , n10652 );
and ( n10786 , n10782 , n10785 );
and ( n10787 , n10780 , n10785 );
or ( n10788 , n10783 , n10786 , n10787 );
and ( n10789 , n10766 , n10788 );
xor ( n10790 , n10655 , n10657 );
xor ( n10791 , n10790 , n10660 );
and ( n10792 , n10788 , n10791 );
and ( n10793 , n10766 , n10791 );
or ( n10794 , n10789 , n10792 , n10793 );
and ( n10795 , n7506 , n7318 );
and ( n10796 , n7945 , n7315 );
nor ( n10797 , n10795 , n10796 );
xnor ( n10798 , n10797 , n7311 );
and ( n10799 , n7547 , n8168 );
and ( n10800 , n7410 , n8166 );
nor ( n10801 , n10799 , n10800 );
xnor ( n10802 , n10801 , n8178 );
and ( n10803 , n10798 , n10802 );
and ( n10804 , n7718 , n7395 );
and ( n10805 , n7516 , n7393 );
nor ( n10806 , n10804 , n10805 );
xnor ( n10807 , n10806 , n7405 );
and ( n10808 , n10802 , n10807 );
and ( n10809 , n10798 , n10807 );
or ( n10810 , n10803 , n10808 , n10809 );
xor ( n10811 , n10597 , n10601 );
xor ( n10812 , n10811 , n10606 );
and ( n10813 , n10810 , n10812 );
xor ( n10814 , n10506 , n10508 );
xor ( n10815 , n10814 , n10511 );
and ( n10816 , n10812 , n10815 );
and ( n10817 , n10810 , n10815 );
or ( n10818 , n10813 , n10816 , n10817 );
xor ( n10819 , n10546 , n10609 );
xor ( n10820 , n10819 , n10612 );
and ( n10821 , n10818 , n10820 );
xor ( n10822 , n10514 , n10516 );
xor ( n10823 , n10822 , n10519 );
and ( n10824 , n10820 , n10823 );
and ( n10825 , n10818 , n10823 );
or ( n10826 , n10821 , n10824 , n10825 );
and ( n10827 , n10794 , n10826 );
xor ( n10828 , n10615 , n10663 );
xor ( n10829 , n10828 , n10666 );
and ( n10830 , n10826 , n10829 );
and ( n10831 , n10794 , n10829 );
or ( n10832 , n10827 , n10830 , n10831 );
and ( n10833 , n10697 , n10832 );
xor ( n10834 , n10680 , n10682 );
xor ( n10835 , n10834 , n10684 );
and ( n10836 , n10832 , n10835 );
and ( n10837 , n10697 , n10835 );
or ( n10838 , n10833 , n10836 , n10837 );
and ( n10839 , n10695 , n10838 );
xor ( n10840 , n10502 , n10675 );
xor ( n10841 , n10840 , n10687 );
and ( n10842 , n10838 , n10841 );
and ( n10843 , n10695 , n10841 );
or ( n10844 , n10839 , n10842 , n10843 );
and ( n10845 , n10692 , n10844 );
and ( n10846 , n10690 , n10844 );
or ( n10847 , n10693 , n10845 , n10846 );
and ( n10848 , n10499 , n10847 );
and ( n10849 , n10497 , n10847 );
or ( n10850 , n10500 , n10848 , n10849 );
and ( n10851 , n10211 , n10850 );
and ( n10852 , n10209 , n10850 );
or ( n10853 , n10212 , n10851 , n10852 );
and ( n10854 , n10192 , n10853 );
and ( n10855 , n10190 , n10853 );
or ( n10856 , n10193 , n10854 , n10855 );
and ( n10857 , n9973 , n10856 );
xor ( n10858 , n9973 , n10856 );
xor ( n10859 , n10190 , n10192 );
xor ( n10860 , n10859 , n10853 );
xor ( n10861 , n10209 , n10211 );
xor ( n10862 , n10861 , n10850 );
xor ( n10863 , n10497 , n10499 );
xor ( n10864 , n10863 , n10847 );
xor ( n10865 , n10690 , n10692 );
xor ( n10866 , n10865 , n10844 );
xor ( n10867 , n10695 , n10838 );
xor ( n10868 , n10867 , n10841 );
xor ( n10869 , n10522 , n10524 );
xor ( n10870 , n10869 , n10527 );
xor ( n10871 , n10794 , n10826 );
xor ( n10872 , n10871 , n10829 );
and ( n10873 , n10870 , n10872 );
xor ( n10874 , n10766 , n10788 );
xor ( n10875 , n10874 , n10791 );
and ( n10876 , n7558 , n7899 );
and ( n10877 , n7606 , n7897 );
nor ( n10878 , n10876 , n10877 );
xnor ( n10879 , n10878 , n7909 );
and ( n10880 , n7729 , n8044 );
and ( n10881 , n7748 , n8042 );
nor ( n10882 , n10880 , n10881 );
xnor ( n10883 , n10882 , n8054 );
and ( n10884 , n10879 , n10883 );
and ( n10885 , n7871 , n7781 );
and ( n10886 , n7800 , n7779 );
nor ( n10887 , n10885 , n10886 );
xnor ( n10888 , n10887 , n7791 );
and ( n10889 , n10883 , n10888 );
and ( n10890 , n10879 , n10888 );
or ( n10891 , n10884 , n10889 , n10890 );
and ( n10892 , n7410 , n7318 );
and ( n10893 , n7506 , n7315 );
nor ( n10894 , n10892 , n10893 );
xnor ( n10895 , n10894 , n7311 );
and ( n10896 , n7516 , n8168 );
and ( n10897 , n7547 , n8166 );
nor ( n10898 , n10896 , n10897 );
xnor ( n10899 , n10898 , n8178 );
and ( n10900 , n10895 , n10899 );
and ( n10901 , n10891 , n10900 );
and ( n10902 , n7618 , n7933 );
and ( n10903 , n7666 , n7931 );
nor ( n10904 , n10902 , n10903 );
xnor ( n10905 , n10904 , n7939 );
xor ( n10906 , n10879 , n10883 );
xor ( n10907 , n10906 , n10888 );
and ( n10908 , n10905 , n10907 );
xor ( n10909 , n10895 , n10899 );
and ( n10910 , n10907 , n10909 );
and ( n10911 , n10905 , n10909 );
or ( n10912 , n10908 , n10910 , n10911 );
and ( n10913 , n10900 , n10912 );
and ( n10914 , n10891 , n10912 );
or ( n10915 , n10901 , n10913 , n10914 );
xor ( n10916 , n10723 , n10758 );
xor ( n10917 , n10916 , n10763 );
and ( n10918 , n10915 , n10917 );
and ( n10919 , n7547 , n7318 );
and ( n10920 , n7410 , n7315 );
nor ( n10921 , n10919 , n10920 );
xnor ( n10922 , n10921 , n7311 );
and ( n10923 , n7718 , n8168 );
and ( n10924 , n7516 , n8166 );
nor ( n10925 , n10923 , n10924 );
xnor ( n10926 , n10925 , n8178 );
and ( n10927 , n10922 , n10926 );
and ( n10928 , n7800 , n8044 );
and ( n10929 , n7729 , n8042 );
nor ( n10930 , n10928 , n10929 );
xnor ( n10931 , n10930 , n8054 );
and ( n10932 , n10926 , n10931 );
and ( n10933 , n10922 , n10931 );
or ( n10934 , n10927 , n10932 , n10933 );
and ( n10935 , n7666 , n7781 );
and ( n10936 , n7871 , n7779 );
nor ( n10937 , n10935 , n10936 );
xnor ( n10938 , n10937 , n7791 );
and ( n10939 , n7809 , n7933 );
and ( n10940 , n7618 , n7931 );
nor ( n10941 , n10939 , n10940 );
xnor ( n10942 , n10941 , n7939 );
and ( n10943 , n10938 , n10942 );
and ( n10944 , n7838 , n7501 );
and ( n10945 , n7676 , n7499 );
nor ( n10946 , n10944 , n10945 );
xnor ( n10947 , n10946 , n7511 );
and ( n10948 , n10942 , n10947 );
and ( n10949 , n10938 , n10947 );
or ( n10950 , n10943 , n10948 , n10949 );
and ( n10951 , n10934 , n10950 );
and ( n10952 , n8066 , n7542 );
and ( n10953 , n7851 , n7540 );
nor ( n10954 , n10952 , n10953 );
xnor ( n10955 , n10954 , n7552 );
and ( n10956 , n8263 , n7713 );
and ( n10957 , n8079 , n7711 );
nor ( n10958 , n10956 , n10957 );
xnor ( n10959 , n10958 , n7723 );
and ( n10960 , n10955 , n10959 );
and ( n10961 , n7516 , n7318 );
and ( n10962 , n7547 , n7315 );
nor ( n10963 , n10961 , n10962 );
xnor ( n10964 , n10963 , n7311 );
and ( n10965 , n7729 , n7899 );
and ( n10966 , n7748 , n7897 );
nor ( n10967 , n10965 , n10966 );
xnor ( n10968 , n10967 , n7909 );
and ( n10969 , n10964 , n10968 );
and ( n10970 , n7871 , n8044 );
and ( n10971 , n7800 , n8042 );
nor ( n10972 , n10970 , n10971 );
xnor ( n10973 , n10972 , n8054 );
and ( n10974 , n10968 , n10973 );
and ( n10975 , n10964 , n10973 );
or ( n10976 , n10969 , n10974 , n10975 );
and ( n10977 , n10959 , n10976 );
and ( n10978 , n10955 , n10976 );
or ( n10979 , n10960 , n10977 , n10978 );
and ( n10980 , n10950 , n10979 );
and ( n10981 , n10934 , n10979 );
or ( n10982 , n10951 , n10980 , n10981 );
xor ( n10983 , n10891 , n10900 );
xor ( n10984 , n10983 , n10912 );
and ( n10985 , n10982 , n10984 );
xor ( n10986 , n10711 , n10715 );
xor ( n10987 , n10986 , n10720 );
and ( n10988 , n10984 , n10987 );
and ( n10989 , n10982 , n10987 );
or ( n10990 , n10985 , n10988 , n10989 );
and ( n10991 , n10917 , n10990 );
and ( n10992 , n10915 , n10990 );
or ( n10993 , n10918 , n10991 , n10992 );
and ( n10994 , n10875 , n10993 );
xor ( n10995 , n10818 , n10820 );
xor ( n10996 , n10995 , n10823 );
and ( n10997 , n10993 , n10996 );
and ( n10998 , n10875 , n10996 );
or ( n10999 , n10994 , n10997 , n10998 );
and ( n11000 , n10872 , n10999 );
and ( n11001 , n10870 , n10999 );
or ( n11002 , n10873 , n11000 , n11001 );
xor ( n11003 , n10697 , n10832 );
xor ( n11004 , n11003 , n10835 );
and ( n11005 , n11002 , n11004 );
and ( n11006 , n8079 , n7542 );
and ( n11007 , n8066 , n7540 );
nor ( n11008 , n11006 , n11007 );
xnor ( n11009 , n11008 , n7552 );
and ( n11010 , n8429 , n7713 );
and ( n11011 , n8263 , n7711 );
nor ( n11012 , n11010 , n11011 );
xnor ( n11013 , n11012 , n7723 );
and ( n11014 , n11009 , n11013 );
and ( n11015 , n9280 , n7743 );
and ( n11016 , n9196 , n7741 );
nor ( n11017 , n11015 , n11016 );
xnor ( n11018 , n11017 , n7753 );
and ( n11019 , n11013 , n11018 );
and ( n11020 , n11009 , n11018 );
or ( n11021 , n11014 , n11019 , n11020 );
and ( n11022 , n7696 , n7954 );
and ( n11023 , n7828 , n7952 );
nor ( n11024 , n11022 , n11023 );
xnor ( n11025 , n11024 , n7964 );
and ( n11026 , n11021 , n11025 );
xor ( n11027 , n10724 , n10728 );
xor ( n11028 , n11027 , n10733 );
and ( n11029 , n11025 , n11028 );
and ( n11030 , n11021 , n11028 );
or ( n11031 , n11026 , n11029 , n11030 );
and ( n11032 , n7704 , n7395 );
and ( n11033 , n7718 , n7393 );
nor ( n11034 , n11032 , n11033 );
xnor ( n11035 , n11034 , n7405 );
and ( n11036 , n11031 , n11035 );
xor ( n11037 , n10701 , n10705 );
xor ( n11038 , n11037 , n10708 );
and ( n11039 , n11035 , n11038 );
and ( n11040 , n11031 , n11038 );
or ( n11041 , n11036 , n11039 , n11040 );
xor ( n11042 , n10798 , n10802 );
xor ( n11043 , n11042 , n10807 );
and ( n11044 , n11041 , n11043 );
xor ( n11045 , n10770 , n10774 );
xor ( n11046 , n11045 , n10777 );
and ( n11047 , n11043 , n11046 );
and ( n11048 , n11041 , n11046 );
or ( n11049 , n11044 , n11047 , n11048 );
xor ( n11050 , n10780 , n10782 );
xor ( n11051 , n11050 , n10785 );
and ( n11052 , n11049 , n11051 );
xor ( n11053 , n10810 , n10812 );
xor ( n11054 , n11053 , n10815 );
and ( n11055 , n11051 , n11054 );
and ( n11056 , n11049 , n11054 );
or ( n11057 , n11052 , n11055 , n11056 );
xor ( n11058 , n10587 , n10591 );
xor ( n11059 , n11058 , n10594 );
xor ( n11060 , n10748 , n10752 );
xor ( n11061 , n11060 , n10755 );
and ( n11062 , n11059 , n11061 );
and ( n11063 , n7828 , n7954 );
and ( n11064 , n7809 , n7952 );
nor ( n11065 , n11063 , n11064 );
xnor ( n11066 , n11065 , n7964 );
xor ( n11067 , n10736 , n10740 );
xor ( n11068 , n11067 , n10745 );
and ( n11069 , n11066 , n11068 );
and ( n11070 , n11061 , n11069 );
and ( n11071 , n11059 , n11069 );
or ( n11072 , n11062 , n11070 , n11071 );
and ( n11073 , n7704 , n8168 );
and ( n11074 , n7718 , n8166 );
nor ( n11075 , n11073 , n11074 );
xnor ( n11076 , n11075 , n8178 );
and ( n11077 , n7558 , n7395 );
and ( n11078 , n7606 , n7393 );
nor ( n11079 , n11077 , n11078 );
xnor ( n11080 , n11079 , n7405 );
and ( n11081 , n11076 , n11080 );
and ( n11082 , n7618 , n7781 );
and ( n11083 , n7666 , n7779 );
nor ( n11084 , n11082 , n11083 );
xnor ( n11085 , n11084 , n7791 );
and ( n11086 , n7676 , n7954 );
and ( n11087 , n7696 , n7952 );
nor ( n11088 , n11086 , n11087 );
xnor ( n11089 , n11088 , n7964 );
and ( n11090 , n11085 , n11089 );
and ( n11091 , n9049 , n7601 );
and ( n11092 , n8696 , n7599 );
nor ( n11093 , n11091 , n11092 );
xnor ( n11094 , n11093 , n7611 );
and ( n11095 , n11089 , n11094 );
and ( n11096 , n11085 , n11094 );
or ( n11097 , n11090 , n11095 , n11096 );
and ( n11098 , n11081 , n11097 );
xor ( n11099 , n10922 , n10926 );
xor ( n11100 , n11099 , n10931 );
and ( n11101 , n11097 , n11100 );
and ( n11102 , n11081 , n11100 );
or ( n11103 , n11098 , n11101 , n11102 );
xor ( n11104 , n10905 , n10907 );
xor ( n11105 , n11104 , n10909 );
and ( n11106 , n11103 , n11105 );
xor ( n11107 , n10575 , n10579 );
xor ( n11108 , n11107 , n10584 );
and ( n11109 , n11105 , n11108 );
and ( n11110 , n11103 , n11108 );
or ( n11111 , n11106 , n11109 , n11110 );
xor ( n11112 , n10938 , n10942 );
xor ( n11113 , n11112 , n10947 );
xor ( n11114 , n10563 , n10567 );
xor ( n11115 , n11114 , n10572 );
and ( n11116 , n11113 , n11115 );
and ( n11117 , n9701 , n7866 );
and ( n11118 , n9463 , n7864 );
nor ( n11119 , n11117 , n11118 );
xnor ( n11120 , n11119 , n7876 );
and ( n11121 , n10032 , n7661 );
and ( n11122 , n9829 , n7659 );
nor ( n11123 , n11121 , n11122 );
xnor ( n11124 , n11123 , n7671 );
and ( n11125 , n11120 , n11124 );
xor ( n11126 , n11009 , n11013 );
xor ( n11127 , n11126 , n11018 );
and ( n11128 , n11124 , n11127 );
and ( n11129 , n11120 , n11127 );
or ( n11130 , n11125 , n11128 , n11129 );
and ( n11131 , n11115 , n11130 );
and ( n11132 , n11113 , n11130 );
or ( n11133 , n11116 , n11131 , n11132 );
xor ( n11134 , n10964 , n10968 );
xor ( n11135 , n11134 , n10973 );
xor ( n11136 , n10550 , n10562 );
and ( n11137 , n11135 , n11136 );
xor ( n11138 , n11076 , n11080 );
and ( n11139 , n11136 , n11138 );
and ( n11140 , n11135 , n11138 );
or ( n11141 , n11137 , n11139 , n11140 );
and ( n11142 , n7606 , n8168 );
and ( n11143 , n7704 , n8166 );
nor ( n11144 , n11142 , n11143 );
xnor ( n11145 , n11144 , n8178 );
and ( n11146 , n7748 , n7395 );
and ( n11147 , n7558 , n7393 );
nor ( n11148 , n11146 , n11147 );
xnor ( n11149 , n11148 , n7405 );
and ( n11150 , n11145 , n11149 );
and ( n11151 , n7809 , n7781 );
and ( n11152 , n7618 , n7779 );
nor ( n11153 , n11151 , n11152 );
xnor ( n11154 , n11153 , n7791 );
and ( n11155 , n11149 , n11154 );
and ( n11156 , n11145 , n11154 );
or ( n11157 , n11150 , n11155 , n11156 );
and ( n11158 , n7800 , n7899 );
and ( n11159 , n7729 , n7897 );
nor ( n11160 , n11158 , n11159 );
xnor ( n11161 , n11160 , n7909 );
and ( n11162 , n7666 , n8044 );
and ( n11163 , n7871 , n8042 );
nor ( n11164 , n11162 , n11163 );
xnor ( n11165 , n11164 , n8054 );
and ( n11166 , n11161 , n11165 );
and ( n11167 , n8066 , n7501 );
and ( n11168 , n7851 , n7499 );
nor ( n11169 , n11167 , n11168 );
xnor ( n11170 , n11169 , n7511 );
and ( n11171 , n11165 , n11170 );
and ( n11172 , n11161 , n11170 );
or ( n11173 , n11166 , n11171 , n11172 );
and ( n11174 , n11157 , n11173 );
and ( n11175 , n8263 , n7542 );
and ( n11176 , n8079 , n7540 );
nor ( n11177 , n11175 , n11176 );
xnor ( n11178 , n11177 , n7552 );
and ( n11179 , n10559 , n7823 );
and ( n11180 , n10377 , n7821 );
nor ( n11181 , n11179 , n11180 );
xnor ( n11182 , n11181 , n7833 );
and ( n11183 , n11178 , n11182 );
xor ( n11184 , n7113 , n7238 );
buf ( n11185 , n11184 );
buf ( n11186 , n11185 );
buf ( n11187 , n11186 );
and ( n11188 , n11187 , n7691 );
and ( n11189 , n10554 , n7689 );
nor ( n11190 , n11188 , n11189 );
not ( n11191 , n11190 );
and ( n11192 , n11182 , n11191 );
and ( n11193 , n11178 , n11191 );
or ( n11194 , n11183 , n11192 , n11193 );
and ( n11195 , n11173 , n11194 );
and ( n11196 , n11157 , n11194 );
or ( n11197 , n11174 , n11195 , n11196 );
and ( n11198 , n11141 , n11197 );
xor ( n11199 , n10955 , n10959 );
xor ( n11200 , n11199 , n10976 );
and ( n11201 , n11197 , n11200 );
and ( n11202 , n11141 , n11200 );
or ( n11203 , n11198 , n11201 , n11202 );
and ( n11204 , n11133 , n11203 );
xor ( n11205 , n10934 , n10950 );
xor ( n11206 , n11205 , n10979 );
and ( n11207 , n11203 , n11206 );
and ( n11208 , n11133 , n11206 );
or ( n11209 , n11204 , n11207 , n11208 );
and ( n11210 , n11111 , n11209 );
xor ( n11211 , n11041 , n11043 );
xor ( n11212 , n11211 , n11046 );
and ( n11213 , n11209 , n11212 );
and ( n11214 , n11111 , n11212 );
or ( n11215 , n11210 , n11213 , n11214 );
and ( n11216 , n11072 , n11215 );
xor ( n11217 , n11031 , n11035 );
xor ( n11218 , n11217 , n11038 );
xor ( n11219 , n11066 , n11068 );
and ( n11220 , n11218 , n11219 );
and ( n11221 , n7606 , n7395 );
and ( n11222 , n7704 , n7393 );
nor ( n11223 , n11221 , n11222 );
xnor ( n11224 , n11223 , n7405 );
and ( n11225 , n7748 , n7899 );
and ( n11226 , n7558 , n7897 );
nor ( n11227 , n11225 , n11226 );
xnor ( n11228 , n11227 , n7909 );
and ( n11229 , n11224 , n11228 );
xor ( n11230 , n11021 , n11025 );
xor ( n11231 , n11230 , n11028 );
and ( n11232 , n11228 , n11231 );
and ( n11233 , n11224 , n11231 );
or ( n11234 , n11229 , n11232 , n11233 );
and ( n11235 , n11219 , n11234 );
and ( n11236 , n11218 , n11234 );
or ( n11237 , n11220 , n11235 , n11236 );
xor ( n11238 , n11081 , n11097 );
xor ( n11239 , n11238 , n11100 );
xor ( n11240 , n11085 , n11089 );
xor ( n11241 , n11240 , n11094 );
and ( n11242 , n10554 , n7823 );
and ( n11243 , n10559 , n7821 );
nor ( n11244 , n11242 , n11243 );
xnor ( n11245 , n11244 , n7833 );
xor ( n11246 , n7136 , n7236 );
buf ( n11247 , n11246 );
buf ( n11248 , n11247 );
buf ( n11249 , n11248 );
and ( n11250 , n11249 , n7691 );
and ( n11251 , n11187 , n7689 );
nor ( n11252 , n11250 , n11251 );
not ( n11253 , n11252 );
and ( n11254 , n11245 , n11253 );
and ( n11255 , n10239 , n7661 );
and ( n11256 , n10032 , n7659 );
nor ( n11257 , n11255 , n11256 );
xnor ( n11258 , n11257 , n7671 );
and ( n11259 , n11254 , n11258 );
and ( n11260 , n11241 , n11259 );
xor ( n11261 , n11145 , n11149 );
xor ( n11262 , n11261 , n11154 );
and ( n11263 , n7704 , n7318 );
and ( n11264 , n7718 , n7315 );
nor ( n11265 , n11263 , n11264 );
xnor ( n11266 , n11265 , n7311 );
and ( n11267 , n7558 , n8168 );
and ( n11268 , n7606 , n8166 );
nor ( n11269 , n11267 , n11268 );
xnor ( n11270 , n11269 , n8178 );
and ( n11271 , n11266 , n11270 );
and ( n11272 , n7828 , n7781 );
and ( n11273 , n7809 , n7779 );
nor ( n11274 , n11272 , n11273 );
xnor ( n11275 , n11274 , n7791 );
and ( n11276 , n11270 , n11275 );
and ( n11277 , n11266 , n11275 );
or ( n11278 , n11271 , n11276 , n11277 );
and ( n11279 , n11262 , n11278 );
xor ( n11280 , n11161 , n11165 );
xor ( n11281 , n11280 , n11170 );
and ( n11282 , n11278 , n11281 );
and ( n11283 , n11262 , n11281 );
or ( n11284 , n11279 , n11282 , n11283 );
and ( n11285 , n11259 , n11284 );
and ( n11286 , n11241 , n11284 );
or ( n11287 , n11260 , n11285 , n11286 );
and ( n11288 , n11239 , n11287 );
xor ( n11289 , n11120 , n11124 );
xor ( n11290 , n11289 , n11127 );
xor ( n11291 , n11135 , n11136 );
xor ( n11292 , n11291 , n11138 );
and ( n11293 , n11290 , n11292 );
xor ( n11294 , n11157 , n11173 );
xor ( n11295 , n11294 , n11194 );
and ( n11296 , n11292 , n11295 );
and ( n11297 , n11290 , n11295 );
or ( n11298 , n11293 , n11296 , n11297 );
and ( n11299 , n11287 , n11298 );
and ( n11300 , n11239 , n11298 );
or ( n11301 , n11288 , n11299 , n11300 );
xor ( n11302 , n11103 , n11105 );
xor ( n11303 , n11302 , n11108 );
and ( n11304 , n11301 , n11303 );
xor ( n11305 , n11133 , n11203 );
xor ( n11306 , n11305 , n11206 );
and ( n11307 , n11303 , n11306 );
and ( n11308 , n11301 , n11306 );
or ( n11309 , n11304 , n11307 , n11308 );
and ( n11310 , n11237 , n11309 );
xor ( n11311 , n10982 , n10984 );
xor ( n11312 , n11311 , n10987 );
and ( n11313 , n11309 , n11312 );
and ( n11314 , n11237 , n11312 );
or ( n11315 , n11310 , n11313 , n11314 );
and ( n11316 , n11215 , n11315 );
and ( n11317 , n11072 , n11315 );
or ( n11318 , n11216 , n11316 , n11317 );
and ( n11319 , n11057 , n11318 );
xor ( n11320 , n10915 , n10917 );
xor ( n11321 , n11320 , n10990 );
xor ( n11322 , n11049 , n11051 );
xor ( n11323 , n11322 , n11054 );
and ( n11324 , n11321 , n11323 );
xor ( n11325 , n11059 , n11061 );
xor ( n11326 , n11325 , n11069 );
xor ( n11327 , n11113 , n11115 );
xor ( n11328 , n11327 , n11130 );
xor ( n11329 , n11141 , n11197 );
xor ( n11330 , n11329 , n11200 );
and ( n11331 , n11328 , n11330 );
xor ( n11332 , n11224 , n11228 );
xor ( n11333 , n11332 , n11231 );
and ( n11334 , n11330 , n11333 );
and ( n11335 , n11328 , n11333 );
or ( n11336 , n11331 , n11334 , n11335 );
xor ( n11337 , n11218 , n11219 );
xor ( n11338 , n11337 , n11234 );
and ( n11339 , n11336 , n11338 );
xor ( n11340 , n11301 , n11303 );
xor ( n11341 , n11340 , n11306 );
and ( n11342 , n11338 , n11341 );
and ( n11343 , n11336 , n11341 );
or ( n11344 , n11339 , n11342 , n11343 );
and ( n11345 , n11326 , n11344 );
xor ( n11346 , n11111 , n11209 );
xor ( n11347 , n11346 , n11212 );
and ( n11348 , n11344 , n11347 );
and ( n11349 , n11326 , n11347 );
or ( n11350 , n11345 , n11348 , n11349 );
and ( n11351 , n11323 , n11350 );
and ( n11352 , n11321 , n11350 );
or ( n11353 , n11324 , n11351 , n11352 );
and ( n11354 , n11318 , n11353 );
and ( n11355 , n11057 , n11353 );
or ( n11356 , n11319 , n11354 , n11355 );
xor ( n11357 , n10870 , n10872 );
xor ( n11358 , n11357 , n10999 );
and ( n11359 , n11356 , n11358 );
xor ( n11360 , n10875 , n10993 );
xor ( n11361 , n11360 , n10996 );
xor ( n11362 , n11057 , n11318 );
xor ( n11363 , n11362 , n11353 );
and ( n11364 , n11361 , n11363 );
xor ( n11365 , n11072 , n11215 );
xor ( n11366 , n11365 , n11315 );
xor ( n11367 , n11321 , n11323 );
xor ( n11368 , n11367 , n11350 );
and ( n11369 , n11366 , n11368 );
xor ( n11370 , n11237 , n11309 );
xor ( n11371 , n11370 , n11312 );
xor ( n11372 , n11326 , n11344 );
xor ( n11373 , n11372 , n11347 );
and ( n11374 , n11371 , n11373 );
xor ( n11375 , n11245 , n11253 );
and ( n11376 , n11187 , n7823 );
and ( n11377 , n10554 , n7821 );
nor ( n11378 , n11376 , n11377 );
xnor ( n11379 , n11378 , n7833 );
xor ( n11380 , n7158 , n7234 );
buf ( n11381 , n11380 );
buf ( n11382 , n11381 );
buf ( n11383 , n11382 );
and ( n11384 , n11383 , n7691 );
and ( n11385 , n11249 , n7689 );
nor ( n11386 , n11384 , n11385 );
not ( n11387 , n11386 );
and ( n11388 , n11379 , n11387 );
and ( n11389 , n11375 , n11388 );
and ( n11390 , n10377 , n7661 );
and ( n11391 , n10239 , n7659 );
nor ( n11392 , n11390 , n11391 );
xnor ( n11393 , n11392 , n7671 );
and ( n11394 , n11388 , n11393 );
and ( n11395 , n11375 , n11393 );
or ( n11396 , n11389 , n11394 , n11395 );
and ( n11397 , n9463 , n7743 );
and ( n11398 , n9280 , n7741 );
nor ( n11399 , n11397 , n11398 );
xnor ( n11400 , n11399 , n7753 );
and ( n11401 , n11396 , n11400 );
and ( n11402 , n9829 , n7866 );
and ( n11403 , n9701 , n7864 );
nor ( n11404 , n11402 , n11403 );
xnor ( n11405 , n11404 , n7876 );
and ( n11406 , n11400 , n11405 );
and ( n11407 , n11396 , n11405 );
or ( n11408 , n11401 , n11406 , n11407 );
xor ( n11409 , n11178 , n11182 );
xor ( n11410 , n11409 , n11191 );
xor ( n11411 , n11254 , n11258 );
and ( n11412 , n11410 , n11411 );
xor ( n11413 , n11262 , n11278 );
xor ( n11414 , n11413 , n11281 );
and ( n11415 , n11411 , n11414 );
and ( n11416 , n11410 , n11414 );
or ( n11417 , n11412 , n11415 , n11416 );
and ( n11418 , n11408 , n11417 );
xor ( n11419 , n11241 , n11259 );
xor ( n11420 , n11419 , n11284 );
and ( n11421 , n11417 , n11420 );
and ( n11422 , n11408 , n11420 );
or ( n11423 , n11418 , n11421 , n11422 );
xor ( n11424 , n11239 , n11287 );
xor ( n11425 , n11424 , n11298 );
and ( n11426 , n11423 , n11425 );
xor ( n11427 , n11379 , n11387 );
and ( n11428 , n11249 , n7823 );
and ( n11429 , n11187 , n7821 );
nor ( n11430 , n11428 , n11429 );
xnor ( n11431 , n11430 , n7833 );
xor ( n11432 , n7175 , n7232 );
buf ( n11433 , n11432 );
buf ( n11434 , n11433 );
buf ( n11435 , n11434 );
and ( n11436 , n11435 , n7691 );
and ( n11437 , n11383 , n7689 );
nor ( n11438 , n11436 , n11437 );
not ( n11439 , n11438 );
and ( n11440 , n11431 , n11439 );
and ( n11441 , n11427 , n11440 );
and ( n11442 , n10559 , n7661 );
and ( n11443 , n10377 , n7659 );
nor ( n11444 , n11442 , n11443 );
xnor ( n11445 , n11444 , n7671 );
and ( n11446 , n11440 , n11445 );
and ( n11447 , n11427 , n11445 );
or ( n11448 , n11441 , n11446 , n11447 );
and ( n11449 , n9701 , n7743 );
and ( n11450 , n9463 , n7741 );
nor ( n11451 , n11449 , n11450 );
xnor ( n11452 , n11451 , n7753 );
and ( n11453 , n11448 , n11452 );
and ( n11454 , n10032 , n7866 );
and ( n11455 , n9829 , n7864 );
nor ( n11456 , n11454 , n11455 );
xnor ( n11457 , n11456 , n7876 );
and ( n11458 , n11452 , n11457 );
and ( n11459 , n11448 , n11457 );
or ( n11460 , n11453 , n11458 , n11459 );
and ( n11461 , n8696 , n7713 );
and ( n11462 , n8429 , n7711 );
nor ( n11463 , n11461 , n11462 );
xnor ( n11464 , n11463 , n7723 );
and ( n11465 , n11460 , n11464 );
and ( n11466 , n9196 , n7601 );
and ( n11467 , n9049 , n7599 );
nor ( n11468 , n11466 , n11467 );
xnor ( n11469 , n11468 , n7611 );
and ( n11470 , n11464 , n11469 );
and ( n11471 , n11460 , n11469 );
or ( n11472 , n11465 , n11470 , n11471 );
and ( n11473 , n7851 , n7501 );
and ( n11474 , n7838 , n7499 );
nor ( n11475 , n11473 , n11474 );
xnor ( n11476 , n11475 , n7511 );
and ( n11477 , n11472 , n11476 );
and ( n11478 , n11425 , n11477 );
and ( n11479 , n11423 , n11477 );
or ( n11480 , n11426 , n11478 , n11479 );
xor ( n11481 , n11336 , n11338 );
xor ( n11482 , n11481 , n11341 );
and ( n11483 , n11480 , n11482 );
and ( n11484 , n9049 , n7713 );
and ( n11485 , n8696 , n7711 );
nor ( n11486 , n11484 , n11485 );
xnor ( n11487 , n11486 , n7723 );
and ( n11488 , n9280 , n7601 );
and ( n11489 , n9196 , n7599 );
nor ( n11490 , n11488 , n11489 );
xnor ( n11491 , n11490 , n7611 );
and ( n11492 , n11487 , n11491 );
xor ( n11493 , n11375 , n11388 );
xor ( n11494 , n11493 , n11393 );
and ( n11495 , n11491 , n11494 );
and ( n11496 , n11487 , n11494 );
or ( n11497 , n11492 , n11495 , n11496 );
and ( n11498 , n7838 , n7954 );
and ( n11499 , n7676 , n7952 );
nor ( n11500 , n11498 , n11499 );
xnor ( n11501 , n11500 , n7964 );
and ( n11502 , n11497 , n11501 );
xor ( n11503 , n11396 , n11400 );
xor ( n11504 , n11503 , n11405 );
and ( n11505 , n11501 , n11504 );
and ( n11506 , n11497 , n11504 );
or ( n11507 , n11502 , n11505 , n11506 );
and ( n11508 , n7828 , n7933 );
and ( n11509 , n7809 , n7931 );
nor ( n11510 , n11508 , n11509 );
xnor ( n11511 , n11510 , n7939 );
and ( n11512 , n11507 , n11511 );
xor ( n11513 , n11328 , n11330 );
xor ( n11514 , n11513 , n11333 );
and ( n11515 , n11512 , n11514 );
xor ( n11516 , n11290 , n11292 );
xor ( n11517 , n11516 , n11295 );
xor ( n11518 , n11408 , n11417 );
xor ( n11519 , n11518 , n11420 );
and ( n11520 , n11517 , n11519 );
xor ( n11521 , n11472 , n11476 );
and ( n11522 , n11519 , n11521 );
and ( n11523 , n11517 , n11521 );
or ( n11524 , n11520 , n11522 , n11523 );
and ( n11525 , n11514 , n11524 );
and ( n11526 , n11512 , n11524 );
or ( n11527 , n11515 , n11525 , n11526 );
and ( n11528 , n11482 , n11527 );
and ( n11529 , n11480 , n11527 );
or ( n11530 , n11483 , n11528 , n11529 );
and ( n11531 , n11373 , n11530 );
and ( n11532 , n11371 , n11530 );
or ( n11533 , n11374 , n11531 , n11532 );
and ( n11534 , n11368 , n11533 );
and ( n11535 , n11366 , n11533 );
or ( n11536 , n11369 , n11534 , n11535 );
and ( n11537 , n11363 , n11536 );
and ( n11538 , n11361 , n11536 );
or ( n11539 , n11364 , n11537 , n11538 );
and ( n11540 , n11358 , n11539 );
and ( n11541 , n11356 , n11539 );
or ( n11542 , n11359 , n11540 , n11541 );
and ( n11543 , n11004 , n11542 );
and ( n11544 , n11002 , n11542 );
or ( n11545 , n11005 , n11543 , n11544 );
and ( n11546 , n10868 , n11545 );
xor ( n11547 , n10868 , n11545 );
xor ( n11548 , n11002 , n11004 );
xor ( n11549 , n11548 , n11542 );
xor ( n11550 , n11356 , n11358 );
xor ( n11551 , n11550 , n11539 );
xor ( n11552 , n11361 , n11363 );
xor ( n11553 , n11552 , n11536 );
xor ( n11554 , n11366 , n11368 );
xor ( n11555 , n11554 , n11533 );
xor ( n11556 , n11371 , n11373 );
xor ( n11557 , n11556 , n11530 );
xor ( n11558 , n11423 , n11425 );
xor ( n11559 , n11558 , n11477 );
xor ( n11560 , n11507 , n11511 );
xor ( n11561 , n11431 , n11439 );
and ( n11562 , n11383 , n7823 );
and ( n11563 , n11249 , n7821 );
nor ( n11564 , n11562 , n11563 );
xnor ( n11565 , n11564 , n7833 );
xor ( n11566 , n7191 , n7230 );
buf ( n11567 , n11566 );
buf ( n11568 , n11567 );
buf ( n11569 , n11568 );
and ( n11570 , n11569 , n7691 );
and ( n11571 , n11435 , n7689 );
nor ( n11572 , n11570 , n11571 );
not ( n11573 , n11572 );
and ( n11574 , n11565 , n11573 );
and ( n11575 , n11561 , n11574 );
and ( n11576 , n10554 , n7661 );
and ( n11577 , n10559 , n7659 );
nor ( n11578 , n11576 , n11577 );
xnor ( n11579 , n11578 , n7671 );
and ( n11580 , n11574 , n11579 );
and ( n11581 , n11561 , n11579 );
or ( n11582 , n11575 , n11580 , n11581 );
and ( n11583 , n10239 , n7866 );
and ( n11584 , n10032 , n7864 );
nor ( n11585 , n11583 , n11584 );
xnor ( n11586 , n11585 , n7876 );
and ( n11587 , n11582 , n11586 );
xor ( n11588 , n11427 , n11440 );
xor ( n11589 , n11588 , n11445 );
and ( n11590 , n11586 , n11589 );
and ( n11591 , n11582 , n11589 );
or ( n11592 , n11587 , n11590 , n11591 );
and ( n11593 , n8079 , n7501 );
and ( n11594 , n8066 , n7499 );
nor ( n11595 , n11593 , n11594 );
xnor ( n11596 , n11595 , n7511 );
and ( n11597 , n11592 , n11596 );
and ( n11598 , n8429 , n7542 );
and ( n11599 , n8263 , n7540 );
nor ( n11600 , n11598 , n11599 );
xnor ( n11601 , n11600 , n7552 );
and ( n11602 , n11596 , n11601 );
and ( n11603 , n11592 , n11601 );
or ( n11604 , n11597 , n11602 , n11603 );
and ( n11605 , n7696 , n7933 );
and ( n11606 , n7828 , n7931 );
nor ( n11607 , n11605 , n11606 );
xnor ( n11608 , n11607 , n7939 );
and ( n11609 , n11604 , n11608 );
xor ( n11610 , n11460 , n11464 );
xor ( n11611 , n11610 , n11469 );
and ( n11612 , n11608 , n11611 );
and ( n11613 , n11604 , n11611 );
or ( n11614 , n11609 , n11612 , n11613 );
and ( n11615 , n11560 , n11614 );
and ( n11616 , n8066 , n7954 );
and ( n11617 , n7851 , n7952 );
nor ( n11618 , n11616 , n11617 );
xnor ( n11619 , n11618 , n7964 );
and ( n11620 , n8263 , n7501 );
and ( n11621 , n8079 , n7499 );
nor ( n11622 , n11620 , n11621 );
xnor ( n11623 , n11622 , n7511 );
and ( n11624 , n11619 , n11623 );
xor ( n11625 , n11582 , n11586 );
xor ( n11626 , n11625 , n11589 );
and ( n11627 , n11623 , n11626 );
and ( n11628 , n11619 , n11626 );
or ( n11629 , n11624 , n11627 , n11628 );
and ( n11630 , n7618 , n8044 );
and ( n11631 , n7666 , n8042 );
nor ( n11632 , n11630 , n11631 );
xnor ( n11633 , n11632 , n8054 );
and ( n11634 , n11629 , n11633 );
xor ( n11635 , n11592 , n11596 );
xor ( n11636 , n11635 , n11601 );
and ( n11637 , n11633 , n11636 );
and ( n11638 , n11629 , n11636 );
or ( n11639 , n11634 , n11637 , n11638 );
and ( n11640 , n7718 , n7318 );
and ( n11641 , n7516 , n7315 );
nor ( n11642 , n11640 , n11641 );
xnor ( n11643 , n11642 , n7311 );
and ( n11644 , n11639 , n11643 );
xor ( n11645 , n11604 , n11608 );
xor ( n11646 , n11645 , n11611 );
and ( n11647 , n11643 , n11646 );
and ( n11648 , n11639 , n11646 );
or ( n11649 , n11644 , n11647 , n11648 );
and ( n11650 , n11614 , n11649 );
and ( n11651 , n11560 , n11649 );
or ( n11652 , n11615 , n11650 , n11651 );
and ( n11653 , n11559 , n11652 );
xor ( n11654 , n11512 , n11514 );
xor ( n11655 , n11654 , n11524 );
and ( n11656 , n11652 , n11655 );
and ( n11657 , n11559 , n11655 );
or ( n11658 , n11653 , n11656 , n11657 );
xor ( n11659 , n11480 , n11482 );
xor ( n11660 , n11659 , n11527 );
and ( n11661 , n11658 , n11660 );
xor ( n11662 , n11517 , n11519 );
xor ( n11663 , n11662 , n11521 );
and ( n11664 , n9196 , n7713 );
and ( n11665 , n9049 , n7711 );
nor ( n11666 , n11664 , n11665 );
xnor ( n11667 , n11666 , n7723 );
and ( n11668 , n9463 , n7601 );
and ( n11669 , n9280 , n7599 );
nor ( n11670 , n11668 , n11669 );
xnor ( n11671 , n11670 , n7611 );
and ( n11672 , n11667 , n11671 );
and ( n11673 , n9829 , n7743 );
and ( n11674 , n9701 , n7741 );
nor ( n11675 , n11673 , n11674 );
xnor ( n11676 , n11675 , n7753 );
and ( n11677 , n11671 , n11676 );
and ( n11678 , n11667 , n11676 );
or ( n11679 , n11672 , n11677 , n11678 );
and ( n11680 , n7851 , n7954 );
and ( n11681 , n7838 , n7952 );
nor ( n11682 , n11680 , n11681 );
xnor ( n11683 , n11682 , n7964 );
and ( n11684 , n11679 , n11683 );
xor ( n11685 , n11448 , n11452 );
xor ( n11686 , n11685 , n11457 );
and ( n11687 , n11683 , n11686 );
and ( n11688 , n11679 , n11686 );
or ( n11689 , n11684 , n11687 , n11688 );
and ( n11690 , n11435 , n7823 );
and ( n11691 , n11383 , n7821 );
nor ( n11692 , n11690 , n11691 );
xnor ( n11693 , n11692 , n7833 );
xor ( n11694 , n7203 , n7228 );
buf ( n11695 , n11694 );
buf ( n11696 , n11695 );
buf ( n11697 , n11696 );
and ( n11698 , n11697 , n7691 );
and ( n11699 , n11569 , n7689 );
nor ( n11700 , n11698 , n11699 );
not ( n11701 , n11700 );
xor ( n11702 , n11693 , n11701 );
and ( n11703 , n11569 , n7823 );
and ( n11704 , n11435 , n7821 );
nor ( n11705 , n11703 , n11704 );
xnor ( n11706 , n11705 , n7833 );
xor ( n11707 , n7210 , n7226 );
buf ( n11708 , n11707 );
buf ( n11709 , n11708 );
buf ( n11710 , n11709 );
and ( n11711 , n11710 , n7691 );
and ( n11712 , n11697 , n7689 );
nor ( n11713 , n11711 , n11712 );
not ( n11714 , n11713 );
and ( n11715 , n11706 , n11714 );
and ( n11716 , n11702 , n11715 );
and ( n11717 , n11249 , n7661 );
and ( n11718 , n11187 , n7659 );
nor ( n11719 , n11717 , n11718 );
xnor ( n11720 , n11719 , n7671 );
and ( n11721 , n11715 , n11720 );
and ( n11722 , n11702 , n11720 );
or ( n11723 , n11716 , n11721 , n11722 );
and ( n11724 , n10559 , n7866 );
and ( n11725 , n10377 , n7864 );
nor ( n11726 , n11724 , n11725 );
xnor ( n11727 , n11726 , n7876 );
and ( n11728 , n11723 , n11727 );
xor ( n11729 , n11565 , n11573 );
and ( n11730 , n11693 , n11701 );
xor ( n11731 , n11729 , n11730 );
and ( n11732 , n11187 , n7661 );
and ( n11733 , n10554 , n7659 );
nor ( n11734 , n11732 , n11733 );
xnor ( n11735 , n11734 , n7671 );
xor ( n11736 , n11731 , n11735 );
and ( n11737 , n11727 , n11736 );
and ( n11738 , n11723 , n11736 );
or ( n11739 , n11728 , n11737 , n11738 );
and ( n11740 , n9701 , n7601 );
and ( n11741 , n9463 , n7599 );
nor ( n11742 , n11740 , n11741 );
xnor ( n11743 , n11742 , n7611 );
and ( n11744 , n11739 , n11743 );
and ( n11745 , n10032 , n7743 );
and ( n11746 , n9829 , n7741 );
nor ( n11747 , n11745 , n11746 );
xnor ( n11748 , n11747 , n7753 );
and ( n11749 , n11743 , n11748 );
and ( n11750 , n11739 , n11748 );
or ( n11751 , n11744 , n11749 , n11750 );
and ( n11752 , n11729 , n11730 );
and ( n11753 , n11730 , n11735 );
and ( n11754 , n11729 , n11735 );
or ( n11755 , n11752 , n11753 , n11754 );
and ( n11756 , n10377 , n7866 );
and ( n11757 , n10239 , n7864 );
nor ( n11758 , n11756 , n11757 );
xnor ( n11759 , n11758 , n7876 );
and ( n11760 , n11755 , n11759 );
xor ( n11761 , n11561 , n11574 );
xor ( n11762 , n11761 , n11579 );
and ( n11763 , n11759 , n11762 );
and ( n11764 , n11755 , n11762 );
or ( n11765 , n11760 , n11763 , n11764 );
and ( n11766 , n11751 , n11765 );
and ( n11767 , n8696 , n7542 );
and ( n11768 , n8429 , n7540 );
nor ( n11769 , n11767 , n11768 );
xnor ( n11770 , n11769 , n7552 );
and ( n11771 , n11765 , n11770 );
and ( n11772 , n11751 , n11770 );
or ( n11773 , n11766 , n11771 , n11772 );
and ( n11774 , n7676 , n7933 );
and ( n11775 , n7696 , n7931 );
nor ( n11776 , n11774 , n11775 );
xnor ( n11777 , n11776 , n7939 );
and ( n11778 , n11773 , n11777 );
xor ( n11779 , n11487 , n11491 );
xor ( n11780 , n11779 , n11494 );
and ( n11781 , n11777 , n11780 );
and ( n11782 , n11773 , n11780 );
or ( n11783 , n11778 , n11781 , n11782 );
and ( n11784 , n11689 , n11783 );
xor ( n11785 , n11497 , n11501 );
xor ( n11786 , n11785 , n11504 );
and ( n11787 , n11783 , n11786 );
and ( n11788 , n11689 , n11786 );
or ( n11789 , n11784 , n11787 , n11788 );
and ( n11790 , n11663 , n11789 );
xor ( n11791 , n11560 , n11614 );
xor ( n11792 , n11791 , n11649 );
and ( n11793 , n11789 , n11792 );
and ( n11794 , n11663 , n11792 );
or ( n11795 , n11790 , n11793 , n11794 );
xor ( n11796 , n11559 , n11652 );
xor ( n11797 , n11796 , n11655 );
and ( n11798 , n11795 , n11797 );
xor ( n11799 , n11410 , n11411 );
xor ( n11800 , n11799 , n11414 );
xor ( n11801 , n11639 , n11643 );
xor ( n11802 , n11801 , n11646 );
and ( n11803 , n11800 , n11802 );
xor ( n11804 , n11689 , n11783 );
xor ( n11805 , n11804 , n11786 );
and ( n11806 , n11802 , n11805 );
and ( n11807 , n11800 , n11805 );
or ( n11808 , n11803 , n11806 , n11807 );
xor ( n11809 , n11706 , n11714 );
and ( n11810 , n11697 , n7823 );
and ( n11811 , n11569 , n7821 );
nor ( n11812 , n11810 , n11811 );
xnor ( n11813 , n11812 , n7833 );
xor ( n11814 , n7216 , n7224 );
buf ( n11815 , n11814 );
buf ( n11816 , n11815 );
buf ( n11817 , n11816 );
and ( n11818 , n11817 , n7691 );
and ( n11819 , n11710 , n7689 );
nor ( n11820 , n11818 , n11819 );
not ( n11821 , n11820 );
and ( n11822 , n11813 , n11821 );
and ( n11823 , n11809 , n11822 );
and ( n11824 , n11383 , n7661 );
and ( n11825 , n11249 , n7659 );
nor ( n11826 , n11824 , n11825 );
xnor ( n11827 , n11826 , n7671 );
and ( n11828 , n11822 , n11827 );
and ( n11829 , n11809 , n11827 );
or ( n11830 , n11823 , n11828 , n11829 );
and ( n11831 , n10554 , n7866 );
and ( n11832 , n10559 , n7864 );
nor ( n11833 , n11831 , n11832 );
xnor ( n11834 , n11833 , n7876 );
and ( n11835 , n11830 , n11834 );
xor ( n11836 , n11702 , n11715 );
xor ( n11837 , n11836 , n11720 );
and ( n11838 , n11834 , n11837 );
and ( n11839 , n11830 , n11837 );
or ( n11840 , n11835 , n11838 , n11839 );
and ( n11841 , n9829 , n7601 );
and ( n11842 , n9701 , n7599 );
nor ( n11843 , n11841 , n11842 );
xnor ( n11844 , n11843 , n7611 );
and ( n11845 , n11840 , n11844 );
and ( n11846 , n10239 , n7743 );
and ( n11847 , n10032 , n7741 );
nor ( n11848 , n11846 , n11847 );
xnor ( n11849 , n11848 , n7753 );
and ( n11850 , n11844 , n11849 );
and ( n11851 , n11840 , n11849 );
or ( n11852 , n11845 , n11850 , n11851 );
and ( n11853 , n9049 , n7542 );
and ( n11854 , n8696 , n7540 );
nor ( n11855 , n11853 , n11854 );
xnor ( n11856 , n11855 , n7552 );
and ( n11857 , n11852 , n11856 );
and ( n11858 , n9280 , n7713 );
and ( n11859 , n9196 , n7711 );
nor ( n11860 , n11858 , n11859 );
xnor ( n11861 , n11860 , n7723 );
and ( n11862 , n11856 , n11861 );
and ( n11863 , n11852 , n11861 );
or ( n11864 , n11857 , n11862 , n11863 );
and ( n11865 , n7838 , n7933 );
and ( n11866 , n7676 , n7931 );
nor ( n11867 , n11865 , n11866 );
xnor ( n11868 , n11867 , n7939 );
and ( n11869 , n11864 , n11868 );
xor ( n11870 , n11667 , n11671 );
xor ( n11871 , n11870 , n11676 );
and ( n11872 , n11868 , n11871 );
and ( n11873 , n11864 , n11871 );
or ( n11874 , n11869 , n11872 , n11873 );
and ( n11875 , n7871 , n7899 );
and ( n11876 , n7800 , n7897 );
nor ( n11877 , n11875 , n11876 );
xnor ( n11878 , n11877 , n7909 );
and ( n11879 , n11874 , n11878 );
xor ( n11880 , n11679 , n11683 );
xor ( n11881 , n11880 , n11686 );
and ( n11882 , n11878 , n11881 );
and ( n11883 , n11874 , n11881 );
or ( n11884 , n11879 , n11882 , n11883 );
and ( n11885 , n8079 , n7954 );
and ( n11886 , n8066 , n7952 );
nor ( n11887 , n11885 , n11886 );
xnor ( n11888 , n11887 , n7964 );
and ( n11889 , n8429 , n7501 );
and ( n11890 , n8263 , n7499 );
nor ( n11891 , n11889 , n11890 );
xnor ( n11892 , n11891 , n7511 );
and ( n11893 , n11888 , n11892 );
xor ( n11894 , n11755 , n11759 );
xor ( n11895 , n11894 , n11762 );
and ( n11896 , n11892 , n11895 );
and ( n11897 , n11888 , n11895 );
or ( n11898 , n11893 , n11896 , n11897 );
and ( n11899 , n7696 , n7781 );
and ( n11900 , n7828 , n7779 );
nor ( n11901 , n11899 , n11900 );
xnor ( n11902 , n11901 , n7791 );
and ( n11903 , n11898 , n11902 );
xor ( n11904 , n11751 , n11765 );
xor ( n11905 , n11904 , n11770 );
and ( n11906 , n11902 , n11905 );
and ( n11907 , n11898 , n11905 );
or ( n11908 , n11903 , n11906 , n11907 );
xor ( n11909 , n11773 , n11777 );
xor ( n11910 , n11909 , n11780 );
and ( n11911 , n11908 , n11910 );
and ( n11912 , n11884 , n11911 );
and ( n11913 , n8696 , n7501 );
and ( n11914 , n8429 , n7499 );
nor ( n11915 , n11913 , n11914 );
xnor ( n11916 , n11915 , n7511 );
and ( n11917 , n9463 , n7713 );
and ( n11918 , n9280 , n7711 );
nor ( n11919 , n11917 , n11918 );
xnor ( n11920 , n11919 , n7723 );
and ( n11921 , n11916 , n11920 );
xor ( n11922 , n11723 , n11727 );
xor ( n11923 , n11922 , n11736 );
and ( n11924 , n11920 , n11923 );
and ( n11925 , n11916 , n11923 );
or ( n11926 , n11921 , n11924 , n11925 );
and ( n11927 , n7676 , n7781 );
and ( n11928 , n7696 , n7779 );
nor ( n11929 , n11927 , n11928 );
xnor ( n11930 , n11929 , n7791 );
and ( n11931 , n11926 , n11930 );
xor ( n11932 , n11739 , n11743 );
xor ( n11933 , n11932 , n11748 );
and ( n11934 , n11930 , n11933 );
and ( n11935 , n11926 , n11933 );
or ( n11936 , n11931 , n11934 , n11935 );
and ( n11937 , n7666 , n7899 );
and ( n11938 , n7871 , n7897 );
nor ( n11939 , n11937 , n11938 );
xnor ( n11940 , n11939 , n7909 );
and ( n11941 , n11936 , n11940 );
xor ( n11942 , n11619 , n11623 );
xor ( n11943 , n11942 , n11626 );
and ( n11944 , n11940 , n11943 );
and ( n11945 , n11936 , n11943 );
or ( n11946 , n11941 , n11944 , n11945 );
xor ( n11947 , n11629 , n11633 );
xor ( n11948 , n11947 , n11636 );
and ( n11949 , n11946 , n11948 );
and ( n11950 , n11911 , n11949 );
and ( n11951 , n11884 , n11949 );
or ( n11952 , n11912 , n11950 , n11951 );
and ( n11953 , n11808 , n11952 );
xor ( n11954 , n11663 , n11789 );
xor ( n11955 , n11954 , n11792 );
and ( n11956 , n11952 , n11955 );
and ( n11957 , n11808 , n11955 );
or ( n11958 , n11953 , n11956 , n11957 );
and ( n11959 , n11797 , n11958 );
and ( n11960 , n11795 , n11958 );
or ( n11961 , n11798 , n11959 , n11960 );
and ( n11962 , n11660 , n11961 );
and ( n11963 , n11658 , n11961 );
or ( n11964 , n11661 , n11962 , n11963 );
and ( n11965 , n11557 , n11964 );
xor ( n11966 , n11557 , n11964 );
xor ( n11967 , n11658 , n11660 );
xor ( n11968 , n11967 , n11961 );
xor ( n11969 , n11795 , n11797 );
xor ( n11970 , n11969 , n11958 );
and ( n11971 , n7606 , n7318 );
and ( n11972 , n7704 , n7315 );
nor ( n11973 , n11971 , n11972 );
xnor ( n11974 , n11973 , n7311 );
and ( n11975 , n7748 , n8168 );
and ( n11976 , n7558 , n8166 );
nor ( n11977 , n11975 , n11976 );
xnor ( n11978 , n11977 , n8178 );
and ( n11979 , n11974 , n11978 );
xor ( n11980 , n11864 , n11868 );
xor ( n11981 , n11980 , n11871 );
and ( n11982 , n11978 , n11981 );
and ( n11983 , n11974 , n11981 );
or ( n11984 , n11979 , n11982 , n11983 );
xor ( n11985 , n11874 , n11878 );
xor ( n11986 , n11985 , n11881 );
and ( n11987 , n11984 , n11986 );
and ( n11988 , n7729 , n7395 );
and ( n11989 , n7748 , n7393 );
nor ( n11990 , n11988 , n11989 );
xnor ( n11991 , n11990 , n7405 );
xor ( n11992 , n11908 , n11910 );
and ( n11993 , n11991 , n11992 );
xor ( n11994 , n11946 , n11948 );
and ( n11995 , n11992 , n11994 );
and ( n11996 , n11991 , n11994 );
or ( n11997 , n11993 , n11995 , n11996 );
and ( n11998 , n11987 , n11997 );
xor ( n11999 , n11800 , n11802 );
xor ( n12000 , n11999 , n11805 );
and ( n12001 , n11997 , n12000 );
and ( n12002 , n11987 , n12000 );
or ( n12003 , n11998 , n12001 , n12002 );
xor ( n12004 , n11808 , n11952 );
xor ( n12005 , n12004 , n11955 );
and ( n12006 , n12003 , n12005 );
xor ( n12007 , n11884 , n11911 );
xor ( n12008 , n12007 , n11949 );
xor ( n12009 , n7220 , n7223 );
buf ( n12010 , n12009 );
buf ( n12011 , n12010 );
buf ( n12012 , n12011 );
and ( n12013 , n12012 , n7691 );
and ( n12014 , n11817 , n7689 );
nor ( n12015 , n12013 , n12014 );
not ( n12016 , n12015 );
and ( n12017 , n11569 , n7661 );
and ( n12018 , n11435 , n7659 );
nor ( n12019 , n12017 , n12018 );
xnor ( n12020 , n12019 , n7671 );
and ( n12021 , n11710 , n7823 );
and ( n12022 , n11697 , n7821 );
nor ( n12023 , n12021 , n12022 );
xnor ( n12024 , n12023 , n7833 );
xor ( n12025 , n12020 , n12024 );
and ( n12026 , n12016 , n12025 );
and ( n12027 , n11249 , n7866 );
and ( n12028 , n11187 , n7864 );
nor ( n12029 , n12027 , n12028 );
xnor ( n12030 , n12029 , n7876 );
and ( n12031 , n12026 , n12030 );
xor ( n12032 , n11813 , n11821 );
and ( n12033 , n12020 , n12024 );
xor ( n12034 , n12032 , n12033 );
and ( n12035 , n11435 , n7661 );
and ( n12036 , n11383 , n7659 );
nor ( n12037 , n12035 , n12036 );
xnor ( n12038 , n12037 , n7671 );
xor ( n12039 , n12034 , n12038 );
and ( n12040 , n12030 , n12039 );
and ( n12041 , n12026 , n12039 );
or ( n12042 , n12031 , n12040 , n12041 );
and ( n12043 , n10559 , n7743 );
and ( n12044 , n10377 , n7741 );
nor ( n12045 , n12043 , n12044 );
xnor ( n12046 , n12045 , n7753 );
and ( n12047 , n12042 , n12046 );
and ( n12048 , n12032 , n12033 );
and ( n12049 , n12033 , n12038 );
and ( n12050 , n12032 , n12038 );
or ( n12051 , n12048 , n12049 , n12050 );
and ( n12052 , n11187 , n7866 );
and ( n12053 , n10554 , n7864 );
nor ( n12054 , n12052 , n12053 );
xnor ( n12055 , n12054 , n7876 );
xor ( n12056 , n12051 , n12055 );
xor ( n12057 , n11809 , n11822 );
xor ( n12058 , n12057 , n11827 );
xor ( n12059 , n12056 , n12058 );
and ( n12060 , n12046 , n12059 );
and ( n12061 , n12042 , n12059 );
or ( n12062 , n12047 , n12060 , n12061 );
and ( n12063 , n9701 , n7713 );
and ( n12064 , n9463 , n7711 );
nor ( n12065 , n12063 , n12064 );
xnor ( n12066 , n12065 , n7723 );
and ( n12067 , n12062 , n12066 );
and ( n12068 , n10032 , n7601 );
and ( n12069 , n9829 , n7599 );
nor ( n12070 , n12068 , n12069 );
xnor ( n12071 , n12070 , n7611 );
and ( n12072 , n12066 , n12071 );
and ( n12073 , n12062 , n12071 );
or ( n12074 , n12067 , n12072 , n12073 );
and ( n12075 , n8066 , n7933 );
and ( n12076 , n7851 , n7931 );
nor ( n12077 , n12075 , n12076 );
xnor ( n12078 , n12077 , n7939 );
and ( n12079 , n12074 , n12078 );
and ( n12080 , n8263 , n7954 );
and ( n12081 , n8079 , n7952 );
nor ( n12082 , n12080 , n12081 );
xnor ( n12083 , n12082 , n7964 );
and ( n12084 , n12078 , n12083 );
and ( n12085 , n12074 , n12083 );
or ( n12086 , n12079 , n12084 , n12085 );
and ( n12087 , n7618 , n7899 );
and ( n12088 , n7666 , n7897 );
nor ( n12089 , n12087 , n12088 );
xnor ( n12090 , n12089 , n7909 );
and ( n12091 , n12086 , n12090 );
xor ( n12092 , n11888 , n11892 );
xor ( n12093 , n12092 , n11895 );
and ( n12094 , n12090 , n12093 );
and ( n12095 , n12086 , n12093 );
or ( n12096 , n12091 , n12094 , n12095 );
xor ( n12097 , n11898 , n11902 );
xor ( n12098 , n12097 , n11905 );
and ( n12099 , n12096 , n12098 );
xor ( n12100 , n11936 , n11940 );
xor ( n12101 , n12100 , n11943 );
and ( n12102 , n12098 , n12101 );
and ( n12103 , n12096 , n12101 );
or ( n12104 , n12099 , n12102 , n12103 );
xor ( n12105 , n11266 , n11270 );
xor ( n12106 , n12105 , n11275 );
and ( n12107 , n12104 , n12106 );
and ( n12108 , n12008 , n12107 );
and ( n12109 , n7800 , n7395 );
and ( n12110 , n7729 , n7393 );
nor ( n12111 , n12109 , n12110 );
xnor ( n12112 , n12111 , n7405 );
and ( n12113 , n7809 , n8044 );
and ( n12114 , n7618 , n8042 );
nor ( n12115 , n12113 , n12114 );
xnor ( n12116 , n12115 , n8054 );
and ( n12117 , n12112 , n12116 );
and ( n12118 , n12051 , n12055 );
and ( n12119 , n12055 , n12058 );
and ( n12120 , n12051 , n12058 );
or ( n12121 , n12118 , n12119 , n12120 );
and ( n12122 , n10377 , n7743 );
and ( n12123 , n10239 , n7741 );
nor ( n12124 , n12122 , n12123 );
xnor ( n12125 , n12124 , n7753 );
and ( n12126 , n12121 , n12125 );
xor ( n12127 , n11830 , n11834 );
xor ( n12128 , n12127 , n11837 );
and ( n12129 , n12125 , n12128 );
and ( n12130 , n12121 , n12128 );
or ( n12131 , n12126 , n12129 , n12130 );
and ( n12132 , n9196 , n7542 );
and ( n12133 , n9049 , n7540 );
nor ( n12134 , n12132 , n12133 );
xnor ( n12135 , n12134 , n7552 );
and ( n12136 , n12131 , n12135 );
xor ( n12137 , n11840 , n11844 );
xor ( n12138 , n12137 , n11849 );
and ( n12139 , n12135 , n12138 );
and ( n12140 , n12131 , n12138 );
or ( n12141 , n12136 , n12139 , n12140 );
and ( n12142 , n7851 , n7933 );
and ( n12143 , n7838 , n7931 );
nor ( n12144 , n12142 , n12143 );
xnor ( n12145 , n12144 , n7939 );
and ( n12146 , n12141 , n12145 );
xor ( n12147 , n11852 , n11856 );
xor ( n12148 , n12147 , n11861 );
and ( n12149 , n12145 , n12148 );
and ( n12150 , n12141 , n12148 );
or ( n12151 , n12146 , n12149 , n12150 );
and ( n12152 , n12116 , n12151 );
and ( n12153 , n12112 , n12151 );
or ( n12154 , n12117 , n12152 , n12153 );
xor ( n12155 , n11984 , n11986 );
and ( n12156 , n12154 , n12155 );
xor ( n12157 , n11991 , n11992 );
xor ( n12158 , n12157 , n11994 );
and ( n12159 , n12155 , n12158 );
and ( n12160 , n12154 , n12158 );
or ( n12161 , n12156 , n12159 , n12160 );
and ( n12162 , n12107 , n12161 );
and ( n12163 , n12008 , n12161 );
or ( n12164 , n12108 , n12162 , n12163 );
and ( n12165 , n12005 , n12164 );
and ( n12166 , n12003 , n12164 );
or ( n12167 , n12006 , n12165 , n12166 );
and ( n12168 , n11970 , n12167 );
xor ( n12169 , n11987 , n11997 );
xor ( n12170 , n12169 , n12000 );
xor ( n12171 , n12104 , n12106 );
and ( n12172 , n8079 , n7933 );
and ( n12173 , n8066 , n7931 );
nor ( n12174 , n12172 , n12173 );
xnor ( n12175 , n12174 , n7939 );
and ( n12176 , n8429 , n7954 );
and ( n12177 , n8263 , n7952 );
nor ( n12178 , n12176 , n12177 );
xnor ( n12179 , n12178 , n7964 );
and ( n12180 , n12175 , n12179 );
xor ( n12181 , n12121 , n12125 );
xor ( n12182 , n12181 , n12128 );
and ( n12183 , n12179 , n12182 );
and ( n12184 , n12175 , n12182 );
or ( n12185 , n12180 , n12183 , n12184 );
and ( n12186 , n7696 , n8044 );
and ( n12187 , n7828 , n8042 );
nor ( n12188 , n12186 , n12187 );
xnor ( n12189 , n12188 , n8054 );
and ( n12190 , n12185 , n12189 );
and ( n12191 , n7838 , n7781 );
and ( n12192 , n7676 , n7779 );
nor ( n12193 , n12191 , n12192 );
xnor ( n12194 , n12193 , n7791 );
and ( n12195 , n12189 , n12194 );
and ( n12196 , n12185 , n12194 );
or ( n12197 , n12190 , n12195 , n12196 );
and ( n12198 , n7558 , n7318 );
and ( n12199 , n7606 , n7315 );
nor ( n12200 , n12198 , n12199 );
xnor ( n12201 , n12200 , n7311 );
and ( n12202 , n12197 , n12201 );
xor ( n12203 , n12086 , n12090 );
xor ( n12204 , n12203 , n12093 );
and ( n12205 , n12201 , n12204 );
and ( n12206 , n12197 , n12204 );
or ( n12207 , n12202 , n12205 , n12206 );
xor ( n12208 , n11974 , n11978 );
xor ( n12209 , n12208 , n11981 );
and ( n12210 , n12207 , n12209 );
xor ( n12211 , n12096 , n12098 );
xor ( n12212 , n12211 , n12101 );
and ( n12213 , n12209 , n12212 );
and ( n12214 , n12207 , n12212 );
or ( n12215 , n12210 , n12213 , n12214 );
and ( n12216 , n12171 , n12215 );
and ( n12217 , n7871 , n7395 );
and ( n12218 , n7800 , n7393 );
nor ( n12219 , n12217 , n12218 );
xnor ( n12220 , n12219 , n7405 );
and ( n12221 , n7828 , n8044 );
and ( n12222 , n7809 , n8042 );
nor ( n12223 , n12221 , n12222 );
xnor ( n12224 , n12223 , n8054 );
and ( n12225 , n12220 , n12224 );
xor ( n12226 , n11926 , n11930 );
xor ( n12227 , n12226 , n11933 );
and ( n12228 , n12224 , n12227 );
and ( n12229 , n12220 , n12227 );
or ( n12230 , n12225 , n12228 , n12229 );
xor ( n12231 , n12112 , n12116 );
xor ( n12232 , n12231 , n12151 );
and ( n12233 , n12230 , n12232 );
and ( n12234 , n11697 , n7661 );
and ( n12235 , n11569 , n7659 );
nor ( n12236 , n12234 , n12235 );
xnor ( n12237 , n12236 , n7671 );
and ( n12238 , n11817 , n7823 );
and ( n12239 , n11710 , n7821 );
nor ( n12240 , n12238 , n12239 );
xnor ( n12241 , n12240 , n7833 );
and ( n12242 , n12237 , n12241 );
buf ( n12243 , n7221 );
buf ( n12244 , n12243 );
buf ( n12245 , n12244 );
buf ( n12246 , n12245 );
and ( n12247 , n12246 , n7691 );
and ( n12248 , n12012 , n7689 );
nor ( n12249 , n12247 , n12248 );
not ( n12250 , n12249 );
and ( n12251 , n12241 , n12250 );
and ( n12252 , n12237 , n12250 );
or ( n12253 , n12242 , n12251 , n12252 );
and ( n12254 , n11187 , n7743 );
and ( n12255 , n10554 , n7741 );
nor ( n12256 , n12254 , n12255 );
xnor ( n12257 , n12256 , n7753 );
and ( n12258 , n12253 , n12257 );
and ( n12259 , n11383 , n7866 );
and ( n12260 , n11249 , n7864 );
nor ( n12261 , n12259 , n12260 );
xnor ( n12262 , n12261 , n7876 );
and ( n12263 , n12257 , n12262 );
and ( n12264 , n12253 , n12262 );
or ( n12265 , n12258 , n12263 , n12264 );
and ( n12266 , n10554 , n7743 );
and ( n12267 , n10559 , n7741 );
nor ( n12268 , n12266 , n12267 );
xnor ( n12269 , n12268 , n7753 );
and ( n12270 , n12265 , n12269 );
xor ( n12271 , n12026 , n12030 );
xor ( n12272 , n12271 , n12039 );
and ( n12273 , n12269 , n12272 );
and ( n12274 , n12265 , n12272 );
or ( n12275 , n12270 , n12273 , n12274 );
and ( n12276 , n9829 , n7713 );
and ( n12277 , n9701 , n7711 );
nor ( n12278 , n12276 , n12277 );
xnor ( n12279 , n12278 , n7723 );
and ( n12280 , n12275 , n12279 );
and ( n12281 , n10239 , n7601 );
and ( n12282 , n10032 , n7599 );
nor ( n12283 , n12281 , n12282 );
xnor ( n12284 , n12283 , n7611 );
and ( n12285 , n12279 , n12284 );
and ( n12286 , n12275 , n12284 );
or ( n12287 , n12280 , n12285 , n12286 );
and ( n12288 , n9049 , n7501 );
and ( n12289 , n8696 , n7499 );
nor ( n12290 , n12288 , n12289 );
xnor ( n12291 , n12290 , n7511 );
and ( n12292 , n12287 , n12291 );
and ( n12293 , n9280 , n7542 );
and ( n12294 , n9196 , n7540 );
nor ( n12295 , n12293 , n12294 );
xnor ( n12296 , n12295 , n7552 );
and ( n12297 , n12291 , n12296 );
and ( n12298 , n12287 , n12296 );
or ( n12299 , n12292 , n12297 , n12298 );
xor ( n12300 , n12131 , n12135 );
xor ( n12301 , n12300 , n12138 );
and ( n12302 , n12299 , n12301 );
xor ( n12303 , n11916 , n11920 );
xor ( n12304 , n12303 , n11923 );
and ( n12305 , n12301 , n12304 );
and ( n12306 , n12299 , n12304 );
or ( n12307 , n12302 , n12305 , n12306 );
and ( n12308 , n7729 , n8168 );
and ( n12309 , n7748 , n8166 );
nor ( n12310 , n12308 , n12309 );
xnor ( n12311 , n12310 , n8178 );
and ( n12312 , n12307 , n12311 );
xor ( n12313 , n12141 , n12145 );
xor ( n12314 , n12313 , n12148 );
and ( n12315 , n12311 , n12314 );
and ( n12316 , n12307 , n12314 );
or ( n12317 , n12312 , n12315 , n12316 );
and ( n12318 , n12232 , n12317 );
and ( n12319 , n12230 , n12317 );
or ( n12320 , n12233 , n12318 , n12319 );
and ( n12321 , n12215 , n12320 );
and ( n12322 , n12171 , n12320 );
or ( n12323 , n12216 , n12321 , n12322 );
and ( n12324 , n12170 , n12323 );
xor ( n12325 , n12008 , n12107 );
xor ( n12326 , n12325 , n12161 );
and ( n12327 , n12323 , n12326 );
and ( n12328 , n12170 , n12326 );
or ( n12329 , n12324 , n12327 , n12328 );
xor ( n12330 , n12003 , n12005 );
xor ( n12331 , n12330 , n12164 );
and ( n12332 , n12329 , n12331 );
xor ( n12333 , n12170 , n12323 );
xor ( n12334 , n12333 , n12326 );
xor ( n12335 , n12154 , n12155 );
xor ( n12336 , n12335 , n12158 );
xor ( n12337 , n12171 , n12215 );
xor ( n12338 , n12337 , n12320 );
and ( n12339 , n12336 , n12338 );
and ( n12340 , n11697 , n7866 );
and ( n12341 , n11569 , n7864 );
nor ( n12342 , n12340 , n12341 );
xnor ( n12343 , n12342 , n7876 );
and ( n12344 , n12246 , n7821 );
not ( n12345 , n12344 );
and ( n12346 , n12345 , n7833 );
and ( n12347 , n12343 , n12346 );
and ( n12348 , n11383 , n7743 );
and ( n12349 , n11249 , n7741 );
nor ( n12350 , n12348 , n12349 );
xnor ( n12351 , n12350 , n7753 );
and ( n12352 , n12347 , n12351 );
and ( n12353 , n11710 , n7661 );
and ( n12354 , n11697 , n7659 );
nor ( n12355 , n12353 , n12354 );
xnor ( n12356 , n12355 , n7671 );
and ( n12357 , n12351 , n12356 );
and ( n12358 , n12347 , n12356 );
or ( n12359 , n12352 , n12357 , n12358 );
and ( n12360 , n10554 , n7601 );
and ( n12361 , n10559 , n7599 );
nor ( n12362 , n12360 , n12361 );
xnor ( n12363 , n12362 , n7611 );
and ( n12364 , n12359 , n12363 );
xor ( n12365 , n12237 , n12241 );
xor ( n12366 , n12365 , n12250 );
and ( n12367 , n12363 , n12366 );
and ( n12368 , n12359 , n12366 );
or ( n12369 , n12364 , n12367 , n12368 );
and ( n12370 , n10239 , n7713 );
and ( n12371 , n10032 , n7711 );
nor ( n12372 , n12370 , n12371 );
xnor ( n12373 , n12372 , n7723 );
and ( n12374 , n12369 , n12373 );
xor ( n12375 , n12253 , n12257 );
xor ( n12376 , n12375 , n12262 );
and ( n12377 , n12373 , n12376 );
and ( n12378 , n12369 , n12376 );
or ( n12379 , n12374 , n12377 , n12378 );
and ( n12380 , n9463 , n7501 );
and ( n12381 , n9280 , n7499 );
nor ( n12382 , n12380 , n12381 );
xnor ( n12383 , n12382 , n7511 );
and ( n12384 , n9829 , n7542 );
and ( n12385 , n9701 , n7540 );
nor ( n12386 , n12384 , n12385 );
xnor ( n12387 , n12386 , n7552 );
and ( n12388 , n12383 , n12387 );
xor ( n12389 , n12016 , n12025 );
and ( n12390 , n11569 , n7866 );
and ( n12391 , n11435 , n7864 );
nor ( n12392 , n12390 , n12391 );
xnor ( n12393 , n12392 , n7876 );
and ( n12394 , n12012 , n7823 );
and ( n12395 , n11817 , n7821 );
nor ( n12396 , n12394 , n12395 );
xnor ( n12397 , n12396 , n7833 );
and ( n12398 , n12393 , n12397 );
and ( n12399 , n12246 , n7689 );
and ( n12400 , n12397 , n12399 );
and ( n12401 , n12393 , n12399 );
or ( n12402 , n12398 , n12400 , n12401 );
and ( n12403 , n11249 , n7743 );
and ( n12404 , n11187 , n7741 );
nor ( n12405 , n12403 , n12404 );
xnor ( n12406 , n12405 , n7753 );
and ( n12407 , n12402 , n12406 );
and ( n12408 , n11435 , n7866 );
and ( n12409 , n11383 , n7864 );
nor ( n12410 , n12408 , n12409 );
xnor ( n12411 , n12410 , n7876 );
and ( n12412 , n12406 , n12411 );
and ( n12413 , n12402 , n12411 );
or ( n12414 , n12407 , n12412 , n12413 );
xor ( n12415 , n12389 , n12414 );
and ( n12416 , n10559 , n7601 );
and ( n12417 , n10377 , n7599 );
nor ( n12418 , n12416 , n12417 );
xnor ( n12419 , n12418 , n7611 );
xor ( n12420 , n12415 , n12419 );
and ( n12421 , n12387 , n12420 );
and ( n12422 , n12383 , n12420 );
or ( n12423 , n12388 , n12421 , n12422 );
and ( n12424 , n12379 , n12423 );
and ( n12425 , n9280 , n7501 );
and ( n12426 , n9196 , n7499 );
nor ( n12427 , n12425 , n12426 );
xnor ( n12428 , n12427 , n7511 );
and ( n12429 , n12423 , n12428 );
and ( n12430 , n12379 , n12428 );
or ( n12431 , n12424 , n12429 , n12430 );
and ( n12432 , n7838 , n8044 );
and ( n12433 , n7676 , n8042 );
nor ( n12434 , n12432 , n12433 );
xnor ( n12435 , n12434 , n8054 );
and ( n12436 , n12431 , n12435 );
and ( n12437 , n8696 , n7954 );
and ( n12438 , n8429 , n7952 );
nor ( n12439 , n12437 , n12438 );
xnor ( n12440 , n12439 , n7964 );
and ( n12441 , n9463 , n7542 );
and ( n12442 , n9280 , n7540 );
nor ( n12443 , n12441 , n12442 );
xnor ( n12444 , n12443 , n7552 );
xor ( n12445 , n12440 , n12444 );
xor ( n12446 , n12042 , n12046 );
xor ( n12447 , n12446 , n12059 );
xor ( n12448 , n12445 , n12447 );
and ( n12449 , n12435 , n12448 );
and ( n12450 , n12431 , n12448 );
or ( n12451 , n12436 , n12449 , n12450 );
and ( n12452 , n7729 , n7318 );
and ( n12453 , n7748 , n7315 );
nor ( n12454 , n12452 , n12453 );
xnor ( n12455 , n12454 , n7311 );
and ( n12456 , n12451 , n12455 );
and ( n12457 , n12389 , n12414 );
and ( n12458 , n12414 , n12419 );
and ( n12459 , n12389 , n12419 );
or ( n12460 , n12457 , n12458 , n12459 );
and ( n12461 , n10032 , n7713 );
and ( n12462 , n9829 , n7711 );
nor ( n12463 , n12461 , n12462 );
xnor ( n12464 , n12463 , n7723 );
and ( n12465 , n12460 , n12464 );
and ( n12466 , n10377 , n7601 );
and ( n12467 , n10239 , n7599 );
nor ( n12468 , n12466 , n12467 );
xnor ( n12469 , n12468 , n7611 );
and ( n12470 , n12464 , n12469 );
and ( n12471 , n12460 , n12469 );
or ( n12472 , n12465 , n12470 , n12471 );
and ( n12473 , n8066 , n7781 );
and ( n12474 , n7851 , n7779 );
nor ( n12475 , n12473 , n12474 );
xnor ( n12476 , n12475 , n7791 );
and ( n12477 , n12472 , n12476 );
and ( n12478 , n9196 , n7501 );
and ( n12479 , n9049 , n7499 );
nor ( n12480 , n12478 , n12479 );
xnor ( n12481 , n12480 , n7511 );
and ( n12482 , n12476 , n12481 );
and ( n12483 , n12472 , n12481 );
or ( n12484 , n12477 , n12482 , n12483 );
and ( n12485 , n7676 , n8044 );
and ( n12486 , n7696 , n8042 );
nor ( n12487 , n12485 , n12486 );
xnor ( n12488 , n12487 , n8054 );
xor ( n12489 , n12484 , n12488 );
and ( n12490 , n7851 , n7781 );
and ( n12491 , n7838 , n7779 );
nor ( n12492 , n12490 , n12491 );
xnor ( n12493 , n12492 , n7791 );
xor ( n12494 , n12489 , n12493 );
and ( n12495 , n12455 , n12494 );
and ( n12496 , n12451 , n12494 );
or ( n12497 , n12456 , n12495 , n12496 );
and ( n12498 , n12440 , n12444 );
and ( n12499 , n12444 , n12447 );
and ( n12500 , n12440 , n12447 );
or ( n12501 , n12498 , n12499 , n12500 );
xor ( n12502 , n12062 , n12066 );
xor ( n12503 , n12502 , n12071 );
and ( n12504 , n12501 , n12503 );
xor ( n12505 , n12287 , n12291 );
xor ( n12506 , n12505 , n12296 );
and ( n12507 , n12503 , n12506 );
and ( n12508 , n12501 , n12506 );
or ( n12509 , n12504 , n12507 , n12508 );
and ( n12510 , n7748 , n7318 );
and ( n12511 , n7558 , n7315 );
nor ( n12512 , n12510 , n12511 );
xnor ( n12513 , n12512 , n7311 );
xor ( n12514 , n12509 , n12513 );
and ( n12515 , n7800 , n8168 );
and ( n12516 , n7729 , n8166 );
nor ( n12517 , n12515 , n12516 );
xnor ( n12518 , n12517 , n8178 );
xor ( n12519 , n12514 , n12518 );
and ( n12520 , n12497 , n12519 );
and ( n12521 , n12484 , n12488 );
and ( n12522 , n12488 , n12493 );
and ( n12523 , n12484 , n12493 );
or ( n12524 , n12521 , n12522 , n12523 );
xor ( n12525 , n12185 , n12189 );
xor ( n12526 , n12525 , n12194 );
xor ( n12527 , n12524 , n12526 );
xor ( n12528 , n12299 , n12301 );
xor ( n12529 , n12528 , n12304 );
xor ( n12530 , n12527 , n12529 );
and ( n12531 , n12519 , n12530 );
and ( n12532 , n12497 , n12530 );
or ( n12533 , n12520 , n12531 , n12532 );
and ( n12534 , n12509 , n12513 );
and ( n12535 , n12513 , n12518 );
and ( n12536 , n12509 , n12518 );
or ( n12537 , n12534 , n12535 , n12536 );
and ( n12538 , n7666 , n7395 );
and ( n12539 , n7871 , n7393 );
nor ( n12540 , n12538 , n12539 );
xnor ( n12541 , n12540 , n7405 );
and ( n12542 , n7809 , n7899 );
and ( n12543 , n7618 , n7897 );
nor ( n12544 , n12542 , n12543 );
xnor ( n12545 , n12544 , n7909 );
and ( n12546 , n12541 , n12545 );
xor ( n12547 , n12074 , n12078 );
xor ( n12548 , n12547 , n12083 );
and ( n12549 , n12545 , n12548 );
and ( n12550 , n12541 , n12548 );
or ( n12551 , n12546 , n12549 , n12550 );
xor ( n12552 , n12537 , n12551 );
xor ( n12553 , n12220 , n12224 );
xor ( n12554 , n12553 , n12227 );
xor ( n12555 , n12552 , n12554 );
and ( n12556 , n12533 , n12555 );
xor ( n12557 , n12197 , n12201 );
xor ( n12558 , n12557 , n12204 );
and ( n12559 , n12555 , n12558 );
and ( n12560 , n12533 , n12558 );
or ( n12561 , n12556 , n12559 , n12560 );
xor ( n12562 , n12207 , n12209 );
xor ( n12563 , n12562 , n12212 );
and ( n12564 , n12561 , n12563 );
and ( n12565 , n12338 , n12564 );
and ( n12566 , n12336 , n12564 );
or ( n12567 , n12339 , n12565 , n12566 );
and ( n12568 , n12334 , n12567 );
and ( n12569 , n12537 , n12551 );
and ( n12570 , n12551 , n12554 );
and ( n12571 , n12537 , n12554 );
or ( n12572 , n12569 , n12570 , n12571 );
xor ( n12573 , n12230 , n12232 );
xor ( n12574 , n12573 , n12317 );
and ( n12575 , n12572 , n12574 );
and ( n12576 , n7871 , n8168 );
and ( n12577 , n7800 , n8166 );
nor ( n12578 , n12576 , n12577 );
xnor ( n12579 , n12578 , n8178 );
and ( n12580 , n7828 , n7899 );
and ( n12581 , n7809 , n7897 );
nor ( n12582 , n12580 , n12581 );
xnor ( n12583 , n12582 , n7909 );
and ( n12584 , n12579 , n12583 );
xor ( n12585 , n12501 , n12503 );
xor ( n12586 , n12585 , n12506 );
and ( n12587 , n12583 , n12586 );
and ( n12588 , n12579 , n12586 );
or ( n12589 , n12584 , n12587 , n12588 );
and ( n12590 , n9049 , n7954 );
and ( n12591 , n8696 , n7952 );
nor ( n12592 , n12590 , n12591 );
xnor ( n12593 , n12592 , n7964 );
and ( n12594 , n9701 , n7542 );
and ( n12595 , n9463 , n7540 );
nor ( n12596 , n12594 , n12595 );
xnor ( n12597 , n12596 , n7552 );
and ( n12598 , n12593 , n12597 );
xor ( n12599 , n12265 , n12269 );
xor ( n12600 , n12599 , n12272 );
and ( n12601 , n12597 , n12600 );
and ( n12602 , n12593 , n12600 );
or ( n12603 , n12598 , n12601 , n12602 );
and ( n12604 , n8263 , n7933 );
and ( n12605 , n8079 , n7931 );
nor ( n12606 , n12604 , n12605 );
xnor ( n12607 , n12606 , n7939 );
and ( n12608 , n12603 , n12607 );
xor ( n12609 , n12275 , n12279 );
xor ( n12610 , n12609 , n12284 );
and ( n12611 , n12607 , n12610 );
and ( n12612 , n12603 , n12610 );
or ( n12613 , n12608 , n12611 , n12612 );
and ( n12614 , n7618 , n7395 );
and ( n12615 , n7666 , n7393 );
nor ( n12616 , n12614 , n12615 );
xnor ( n12617 , n12616 , n7405 );
and ( n12618 , n12613 , n12617 );
xor ( n12619 , n12175 , n12179 );
xor ( n12620 , n12619 , n12182 );
and ( n12621 , n12617 , n12620 );
and ( n12622 , n12613 , n12620 );
or ( n12623 , n12618 , n12621 , n12622 );
and ( n12624 , n12589 , n12623 );
xor ( n12625 , n12541 , n12545 );
xor ( n12626 , n12625 , n12548 );
and ( n12627 , n12623 , n12626 );
and ( n12628 , n12589 , n12626 );
or ( n12629 , n12624 , n12627 , n12628 );
and ( n12630 , n12524 , n12526 );
and ( n12631 , n12526 , n12529 );
and ( n12632 , n12524 , n12529 );
or ( n12633 , n12630 , n12631 , n12632 );
and ( n12634 , n12629 , n12633 );
xor ( n12635 , n12307 , n12311 );
xor ( n12636 , n12635 , n12314 );
and ( n12637 , n12633 , n12636 );
and ( n12638 , n12629 , n12636 );
or ( n12639 , n12634 , n12637 , n12638 );
and ( n12640 , n12574 , n12639 );
and ( n12641 , n12572 , n12639 );
or ( n12642 , n12575 , n12640 , n12641 );
xor ( n12643 , n12561 , n12563 );
and ( n12644 , n8079 , n7781 );
and ( n12645 , n8066 , n7779 );
nor ( n12646 , n12644 , n12645 );
xnor ( n12647 , n12646 , n7791 );
and ( n12648 , n8429 , n7933 );
and ( n12649 , n8263 , n7931 );
nor ( n12650 , n12648 , n12649 );
xnor ( n12651 , n12650 , n7939 );
and ( n12652 , n12647 , n12651 );
xor ( n12653 , n12460 , n12464 );
xor ( n12654 , n12653 , n12469 );
and ( n12655 , n12651 , n12654 );
and ( n12656 , n12647 , n12654 );
or ( n12657 , n12652 , n12655 , n12656 );
and ( n12658 , n7696 , n7899 );
and ( n12659 , n7828 , n7897 );
nor ( n12660 , n12658 , n12659 );
xnor ( n12661 , n12660 , n7909 );
and ( n12662 , n12657 , n12661 );
xor ( n12663 , n12472 , n12476 );
xor ( n12664 , n12663 , n12481 );
and ( n12665 , n12661 , n12664 );
and ( n12666 , n12657 , n12664 );
or ( n12667 , n12662 , n12665 , n12666 );
and ( n12668 , n7800 , n7318 );
and ( n12669 , n7729 , n7315 );
nor ( n12670 , n12668 , n12669 );
xnor ( n12671 , n12670 , n7311 );
and ( n12672 , n7666 , n8168 );
and ( n12673 , n7871 , n8166 );
nor ( n12674 , n12672 , n12673 );
xnor ( n12675 , n12674 , n8178 );
and ( n12676 , n12671 , n12675 );
xor ( n12677 , n12603 , n12607 );
xor ( n12678 , n12677 , n12610 );
and ( n12679 , n12675 , n12678 );
and ( n12680 , n12671 , n12678 );
or ( n12681 , n12676 , n12679 , n12680 );
and ( n12682 , n12667 , n12681 );
xor ( n12683 , n12613 , n12617 );
xor ( n12684 , n12683 , n12620 );
and ( n12685 , n12681 , n12684 );
and ( n12686 , n12667 , n12684 );
or ( n12687 , n12682 , n12685 , n12686 );
xor ( n12688 , n12589 , n12623 );
xor ( n12689 , n12688 , n12626 );
and ( n12690 , n12687 , n12689 );
xor ( n12691 , n12497 , n12519 );
xor ( n12692 , n12691 , n12530 );
and ( n12693 , n12689 , n12692 );
and ( n12694 , n12687 , n12692 );
or ( n12695 , n12690 , n12693 , n12694 );
xor ( n12696 , n12629 , n12633 );
xor ( n12697 , n12696 , n12636 );
and ( n12698 , n12695 , n12697 );
xor ( n12699 , n12533 , n12555 );
xor ( n12700 , n12699 , n12558 );
and ( n12701 , n12697 , n12700 );
and ( n12702 , n12695 , n12700 );
or ( n12703 , n12698 , n12701 , n12702 );
and ( n12704 , n12643 , n12703 );
xor ( n12705 , n12572 , n12574 );
xor ( n12706 , n12705 , n12639 );
and ( n12707 , n12703 , n12706 );
and ( n12708 , n12643 , n12706 );
or ( n12709 , n12704 , n12707 , n12708 );
and ( n12710 , n12642 , n12709 );
xor ( n12711 , n12336 , n12338 );
xor ( n12712 , n12711 , n12564 );
and ( n12713 , n12709 , n12712 );
and ( n12714 , n12642 , n12712 );
or ( n12715 , n12710 , n12713 , n12714 );
and ( n12716 , n12567 , n12715 );
and ( n12717 , n12334 , n12715 );
or ( n12718 , n12568 , n12716 , n12717 );
and ( n12719 , n12331 , n12718 );
and ( n12720 , n12329 , n12718 );
or ( n12721 , n12332 , n12719 , n12720 );
and ( n12722 , n12167 , n12721 );
and ( n12723 , n11970 , n12721 );
or ( n12724 , n12168 , n12722 , n12723 );
and ( n12725 , n11968 , n12724 );
xor ( n12726 , n11968 , n12724 );
xor ( n12727 , n11970 , n12167 );
xor ( n12728 , n12727 , n12721 );
xor ( n12729 , n12329 , n12331 );
xor ( n12730 , n12729 , n12718 );
xor ( n12731 , n12334 , n12567 );
xor ( n12732 , n12731 , n12715 );
xor ( n12733 , n12642 , n12709 );
xor ( n12734 , n12733 , n12712 );
xor ( n12735 , n12643 , n12703 );
xor ( n12736 , n12735 , n12706 );
xor ( n12737 , n12695 , n12697 );
xor ( n12738 , n12737 , n12700 );
and ( n12739 , n9701 , n7501 );
and ( n12740 , n9463 , n7499 );
nor ( n12741 , n12739 , n12740 );
xnor ( n12742 , n12741 , n7511 );
and ( n12743 , n10032 , n7542 );
and ( n12744 , n9829 , n7540 );
nor ( n12745 , n12743 , n12744 );
xnor ( n12746 , n12745 , n7552 );
and ( n12747 , n12742 , n12746 );
xor ( n12748 , n12359 , n12363 );
xor ( n12749 , n12748 , n12366 );
and ( n12750 , n12746 , n12749 );
and ( n12751 , n12742 , n12749 );
or ( n12752 , n12747 , n12750 , n12751 );
xor ( n12753 , n12369 , n12373 );
xor ( n12754 , n12753 , n12376 );
and ( n12755 , n12752 , n12754 );
xor ( n12756 , n12383 , n12387 );
xor ( n12757 , n12756 , n12420 );
and ( n12758 , n12754 , n12757 );
and ( n12759 , n12752 , n12757 );
or ( n12760 , n12755 , n12758 , n12759 );
and ( n12761 , n7676 , n7899 );
and ( n12762 , n7696 , n7897 );
nor ( n12763 , n12761 , n12762 );
xnor ( n12764 , n12763 , n7909 );
and ( n12765 , n12760 , n12764 );
xor ( n12766 , n12379 , n12423 );
xor ( n12767 , n12766 , n12428 );
and ( n12768 , n12764 , n12767 );
and ( n12769 , n12760 , n12767 );
or ( n12770 , n12765 , n12768 , n12769 );
xor ( n12771 , n12343 , n12346 );
and ( n12772 , n11569 , n7743 );
and ( n12773 , n11435 , n7741 );
nor ( n12774 , n12772 , n12773 );
xnor ( n12775 , n12774 , n7753 );
and ( n12776 , n11710 , n7866 );
and ( n12777 , n11697 , n7864 );
nor ( n12778 , n12776 , n12777 );
xnor ( n12779 , n12778 , n7876 );
and ( n12780 , n12775 , n12779 );
and ( n12781 , n12779 , n12344 );
and ( n12782 , n12775 , n12344 );
or ( n12783 , n12780 , n12781 , n12782 );
and ( n12784 , n12771 , n12783 );
and ( n12785 , n11249 , n7601 );
and ( n12786 , n11187 , n7599 );
nor ( n12787 , n12785 , n12786 );
xnor ( n12788 , n12787 , n7611 );
and ( n12789 , n12783 , n12788 );
and ( n12790 , n12771 , n12788 );
or ( n12791 , n12784 , n12789 , n12790 );
and ( n12792 , n10559 , n7713 );
and ( n12793 , n10377 , n7711 );
nor ( n12794 , n12792 , n12793 );
xnor ( n12795 , n12794 , n7723 );
and ( n12796 , n12791 , n12795 );
xor ( n12797 , n12347 , n12351 );
xor ( n12798 , n12797 , n12356 );
and ( n12799 , n12795 , n12798 );
and ( n12800 , n12791 , n12798 );
or ( n12801 , n12796 , n12799 , n12800 );
and ( n12802 , n11697 , n7743 );
and ( n12803 , n11569 , n7741 );
nor ( n12804 , n12802 , n12803 );
xnor ( n12805 , n12804 , n7753 );
and ( n12806 , n12246 , n7659 );
not ( n12807 , n12806 );
and ( n12808 , n12807 , n7671 );
and ( n12809 , n12805 , n12808 );
and ( n12810 , n11383 , n7601 );
and ( n12811 , n11249 , n7599 );
nor ( n12812 , n12810 , n12811 );
xnor ( n12813 , n12812 , n7611 );
and ( n12814 , n12809 , n12813 );
and ( n12815 , n12012 , n7661 );
and ( n12816 , n11817 , n7659 );
nor ( n12817 , n12815 , n12816 );
xnor ( n12818 , n12817 , n7671 );
and ( n12819 , n12813 , n12818 );
and ( n12820 , n12809 , n12818 );
or ( n12821 , n12814 , n12819 , n12820 );
and ( n12822 , n10554 , n7713 );
and ( n12823 , n10559 , n7711 );
nor ( n12824 , n12822 , n12823 );
xnor ( n12825 , n12824 , n7723 );
and ( n12826 , n12821 , n12825 );
and ( n12827 , n11435 , n7743 );
and ( n12828 , n11383 , n7741 );
nor ( n12829 , n12827 , n12828 );
xnor ( n12830 , n12829 , n7753 );
and ( n12831 , n11817 , n7661 );
and ( n12832 , n11710 , n7659 );
nor ( n12833 , n12831 , n12832 );
xnor ( n12834 , n12833 , n7671 );
xor ( n12835 , n12830 , n12834 );
and ( n12836 , n12246 , n7823 );
and ( n12837 , n12012 , n7821 );
nor ( n12838 , n12836 , n12837 );
xnor ( n12839 , n12838 , n7833 );
xor ( n12840 , n12835 , n12839 );
and ( n12841 , n12825 , n12840 );
and ( n12842 , n12821 , n12840 );
or ( n12843 , n12826 , n12841 , n12842 );
and ( n12844 , n10239 , n7542 );
and ( n12845 , n10032 , n7540 );
nor ( n12846 , n12844 , n12845 );
xnor ( n12847 , n12846 , n7552 );
and ( n12848 , n12843 , n12847 );
and ( n12849 , n12830 , n12834 );
and ( n12850 , n12834 , n12839 );
and ( n12851 , n12830 , n12839 );
or ( n12852 , n12849 , n12850 , n12851 );
and ( n12853 , n11187 , n7601 );
and ( n12854 , n10554 , n7599 );
nor ( n12855 , n12853 , n12854 );
xnor ( n12856 , n12855 , n7611 );
xor ( n12857 , n12852 , n12856 );
xor ( n12858 , n12393 , n12397 );
xor ( n12859 , n12858 , n12399 );
xor ( n12860 , n12857 , n12859 );
and ( n12861 , n12847 , n12860 );
and ( n12862 , n12843 , n12860 );
or ( n12863 , n12848 , n12861 , n12862 );
and ( n12864 , n12801 , n12863 );
and ( n12865 , n9280 , n7954 );
and ( n12866 , n9196 , n7952 );
nor ( n12867 , n12865 , n12866 );
xnor ( n12868 , n12867 , n7964 );
and ( n12869 , n12863 , n12868 );
and ( n12870 , n12801 , n12868 );
or ( n12871 , n12864 , n12869 , n12870 );
and ( n12872 , n8066 , n8044 );
and ( n12873 , n7851 , n8042 );
nor ( n12874 , n12872 , n12873 );
xnor ( n12875 , n12874 , n8054 );
and ( n12876 , n12871 , n12875 );
and ( n12877 , n8263 , n7781 );
and ( n12878 , n8079 , n7779 );
nor ( n12879 , n12877 , n12878 );
xnor ( n12880 , n12879 , n7791 );
and ( n12881 , n12875 , n12880 );
and ( n12882 , n12871 , n12880 );
or ( n12883 , n12876 , n12881 , n12882 );
and ( n12884 , n7618 , n8168 );
and ( n12885 , n7666 , n8166 );
nor ( n12886 , n12884 , n12885 );
xnor ( n12887 , n12886 , n8178 );
and ( n12888 , n12883 , n12887 );
xor ( n12889 , n12647 , n12651 );
xor ( n12890 , n12889 , n12654 );
and ( n12891 , n12887 , n12890 );
and ( n12892 , n12883 , n12890 );
or ( n12893 , n12888 , n12891 , n12892 );
and ( n12894 , n12770 , n12893 );
xor ( n12895 , n12657 , n12661 );
xor ( n12896 , n12895 , n12664 );
and ( n12897 , n12893 , n12896 );
and ( n12898 , n12770 , n12896 );
or ( n12899 , n12894 , n12897 , n12898 );
and ( n12900 , n12852 , n12856 );
and ( n12901 , n12856 , n12859 );
and ( n12902 , n12852 , n12859 );
or ( n12903 , n12900 , n12901 , n12902 );
and ( n12904 , n10377 , n7713 );
and ( n12905 , n10239 , n7711 );
nor ( n12906 , n12904 , n12905 );
xnor ( n12907 , n12906 , n7723 );
and ( n12908 , n12903 , n12907 );
xor ( n12909 , n12402 , n12406 );
xor ( n12910 , n12909 , n12411 );
and ( n12911 , n12907 , n12910 );
and ( n12912 , n12903 , n12910 );
or ( n12913 , n12908 , n12911 , n12912 );
and ( n12914 , n8696 , n7933 );
and ( n12915 , n8429 , n7931 );
nor ( n12916 , n12914 , n12915 );
xnor ( n12917 , n12916 , n7939 );
and ( n12918 , n12913 , n12917 );
and ( n12919 , n9196 , n7954 );
and ( n12920 , n9049 , n7952 );
nor ( n12921 , n12919 , n12920 );
xnor ( n12922 , n12921 , n7964 );
and ( n12923 , n12917 , n12922 );
and ( n12924 , n12913 , n12922 );
or ( n12925 , n12918 , n12923 , n12924 );
and ( n12926 , n7851 , n8044 );
and ( n12927 , n7838 , n8042 );
nor ( n12928 , n12926 , n12927 );
xnor ( n12929 , n12928 , n8054 );
and ( n12930 , n12925 , n12929 );
xor ( n12931 , n12593 , n12597 );
xor ( n12932 , n12931 , n12600 );
and ( n12933 , n12929 , n12932 );
and ( n12934 , n12925 , n12932 );
or ( n12935 , n12930 , n12933 , n12934 );
and ( n12936 , n7809 , n7395 );
and ( n12937 , n7618 , n7393 );
nor ( n12938 , n12936 , n12937 );
xnor ( n12939 , n12938 , n7405 );
and ( n12940 , n12935 , n12939 );
xor ( n12941 , n12431 , n12435 );
xor ( n12942 , n12941 , n12448 );
and ( n12943 , n12939 , n12942 );
and ( n12944 , n12935 , n12942 );
or ( n12945 , n12940 , n12943 , n12944 );
and ( n12946 , n12899 , n12945 );
xor ( n12947 , n12579 , n12583 );
xor ( n12948 , n12947 , n12586 );
and ( n12949 , n12945 , n12948 );
and ( n12950 , n12899 , n12948 );
or ( n12951 , n12946 , n12949 , n12950 );
and ( n12952 , n9463 , n7954 );
and ( n12953 , n9280 , n7952 );
nor ( n12954 , n12952 , n12953 );
xnor ( n12955 , n12954 , n7964 );
and ( n12956 , n9829 , n7501 );
and ( n12957 , n9701 , n7499 );
nor ( n12958 , n12956 , n12957 );
xnor ( n12959 , n12958 , n7511 );
and ( n12960 , n12955 , n12959 );
xor ( n12961 , n12791 , n12795 );
xor ( n12962 , n12961 , n12798 );
and ( n12963 , n12959 , n12962 );
and ( n12964 , n12955 , n12962 );
or ( n12965 , n12960 , n12963 , n12964 );
and ( n12966 , n9049 , n7933 );
and ( n12967 , n8696 , n7931 );
nor ( n12968 , n12966 , n12967 );
xnor ( n12969 , n12968 , n7939 );
and ( n12970 , n12965 , n12969 );
xor ( n12971 , n12903 , n12907 );
xor ( n12972 , n12971 , n12910 );
and ( n12973 , n12969 , n12972 );
and ( n12974 , n12965 , n12972 );
or ( n12975 , n12970 , n12973 , n12974 );
and ( n12976 , n7838 , n7899 );
and ( n12977 , n7676 , n7897 );
nor ( n12978 , n12976 , n12977 );
xnor ( n12979 , n12978 , n7909 );
and ( n12980 , n12975 , n12979 );
xor ( n12981 , n12913 , n12917 );
xor ( n12982 , n12981 , n12922 );
and ( n12983 , n12979 , n12982 );
and ( n12984 , n12975 , n12982 );
or ( n12985 , n12980 , n12983 , n12984 );
and ( n12986 , n8079 , n8044 );
and ( n12987 , n8066 , n8042 );
nor ( n12988 , n12986 , n12987 );
xnor ( n12989 , n12988 , n8054 );
and ( n12990 , n8429 , n7781 );
and ( n12991 , n8263 , n7779 );
nor ( n12992 , n12990 , n12991 );
xnor ( n12993 , n12992 , n7791 );
and ( n12994 , n12989 , n12993 );
xor ( n12995 , n12742 , n12746 );
xor ( n12996 , n12995 , n12749 );
and ( n12997 , n12993 , n12996 );
and ( n12998 , n12989 , n12996 );
or ( n12999 , n12994 , n12997 , n12998 );
and ( n13000 , n7696 , n7395 );
and ( n13001 , n7828 , n7393 );
nor ( n13002 , n13000 , n13001 );
xnor ( n13003 , n13002 , n7405 );
and ( n13004 , n12999 , n13003 );
xor ( n13005 , n12752 , n12754 );
xor ( n13006 , n13005 , n12757 );
and ( n13007 , n13003 , n13006 );
and ( n13008 , n12999 , n13006 );
or ( n13009 , n13004 , n13007 , n13008 );
and ( n13010 , n12985 , n13009 );
xor ( n13011 , n12760 , n12764 );
xor ( n13012 , n13011 , n12767 );
and ( n13013 , n13009 , n13012 );
and ( n13014 , n12985 , n13012 );
or ( n13015 , n13010 , n13013 , n13014 );
and ( n13016 , n7871 , n7318 );
and ( n13017 , n7800 , n7315 );
nor ( n13018 , n13016 , n13017 );
xnor ( n13019 , n13018 , n7311 );
and ( n13020 , n7828 , n7395 );
and ( n13021 , n7809 , n7393 );
nor ( n13022 , n13020 , n13021 );
xnor ( n13023 , n13022 , n7405 );
and ( n13024 , n13019 , n13023 );
xor ( n13025 , n12925 , n12929 );
xor ( n13026 , n13025 , n12932 );
and ( n13027 , n13023 , n13026 );
and ( n13028 , n13019 , n13026 );
or ( n13029 , n13024 , n13027 , n13028 );
and ( n13030 , n13015 , n13029 );
xor ( n13031 , n12671 , n12675 );
xor ( n13032 , n13031 , n12678 );
and ( n13033 , n13029 , n13032 );
and ( n13034 , n13015 , n13032 );
or ( n13035 , n13030 , n13033 , n13034 );
xor ( n13036 , n12451 , n12455 );
xor ( n13037 , n13036 , n12494 );
and ( n13038 , n13035 , n13037 );
xor ( n13039 , n12667 , n12681 );
xor ( n13040 , n13039 , n12684 );
and ( n13041 , n13037 , n13040 );
and ( n13042 , n13035 , n13040 );
or ( n13043 , n13038 , n13041 , n13042 );
and ( n13044 , n12951 , n13043 );
xor ( n13045 , n12687 , n12689 );
xor ( n13046 , n13045 , n12692 );
and ( n13047 , n13043 , n13046 );
and ( n13048 , n12951 , n13046 );
or ( n13049 , n13044 , n13047 , n13048 );
and ( n13050 , n12738 , n13049 );
xor ( n13051 , n12738 , n13049 );
xor ( n13052 , n12770 , n12893 );
xor ( n13053 , n13052 , n12896 );
xor ( n13054 , n13015 , n13029 );
xor ( n13055 , n13054 , n13032 );
and ( n13056 , n13053 , n13055 );
xor ( n13057 , n12935 , n12939 );
xor ( n13058 , n13057 , n12942 );
and ( n13059 , n13055 , n13058 );
and ( n13060 , n13053 , n13058 );
or ( n13061 , n13056 , n13059 , n13060 );
xor ( n13062 , n12899 , n12945 );
xor ( n13063 , n13062 , n12948 );
and ( n13064 , n13061 , n13063 );
xor ( n13065 , n13035 , n13037 );
xor ( n13066 , n13065 , n13040 );
and ( n13067 , n13063 , n13066 );
and ( n13068 , n13061 , n13066 );
or ( n13069 , n13064 , n13067 , n13068 );
xor ( n13070 , n12951 , n13043 );
xor ( n13071 , n13070 , n13046 );
and ( n13072 , n13069 , n13071 );
xor ( n13073 , n13069 , n13071 );
xor ( n13074 , n13061 , n13063 );
xor ( n13075 , n13074 , n13066 );
xor ( n13076 , n12805 , n12808 );
and ( n13077 , n11569 , n7601 );
and ( n13078 , n11435 , n7599 );
nor ( n13079 , n13077 , n13078 );
xnor ( n13080 , n13079 , n7611 );
and ( n13081 , n11710 , n7743 );
and ( n13082 , n11697 , n7741 );
nor ( n13083 , n13081 , n13082 );
xnor ( n13084 , n13083 , n7753 );
and ( n13085 , n13080 , n13084 );
and ( n13086 , n13084 , n12806 );
and ( n13087 , n13080 , n12806 );
or ( n13088 , n13085 , n13086 , n13087 );
and ( n13089 , n13076 , n13088 );
and ( n13090 , n11249 , n7713 );
and ( n13091 , n11187 , n7711 );
nor ( n13092 , n13090 , n13091 );
xnor ( n13093 , n13092 , n7723 );
and ( n13094 , n13088 , n13093 );
and ( n13095 , n13076 , n13093 );
or ( n13096 , n13089 , n13094 , n13095 );
and ( n13097 , n10559 , n7542 );
and ( n13098 , n10377 , n7540 );
nor ( n13099 , n13097 , n13098 );
xnor ( n13100 , n13099 , n7552 );
and ( n13101 , n13096 , n13100 );
xor ( n13102 , n12809 , n12813 );
xor ( n13103 , n13102 , n12818 );
and ( n13104 , n13100 , n13103 );
and ( n13105 , n13096 , n13103 );
or ( n13106 , n13101 , n13104 , n13105 );
and ( n13107 , n9701 , n7954 );
and ( n13108 , n9463 , n7952 );
nor ( n13109 , n13107 , n13108 );
xnor ( n13110 , n13109 , n7964 );
and ( n13111 , n13106 , n13110 );
xor ( n13112 , n12821 , n12825 );
xor ( n13113 , n13112 , n12840 );
and ( n13114 , n13110 , n13113 );
and ( n13115 , n13106 , n13113 );
or ( n13116 , n13111 , n13114 , n13115 );
and ( n13117 , n8263 , n8044 );
and ( n13118 , n8079 , n8042 );
nor ( n13119 , n13117 , n13118 );
xnor ( n13120 , n13119 , n8054 );
and ( n13121 , n13116 , n13120 );
and ( n13122 , n9196 , n7933 );
and ( n13123 , n9049 , n7931 );
nor ( n13124 , n13122 , n13123 );
xnor ( n13125 , n13124 , n7939 );
and ( n13126 , n13120 , n13125 );
and ( n13127 , n13116 , n13125 );
or ( n13128 , n13121 , n13126 , n13127 );
and ( n13129 , n7851 , n7899 );
and ( n13130 , n7838 , n7897 );
nor ( n13131 , n13129 , n13130 );
xnor ( n13132 , n13131 , n7909 );
and ( n13133 , n13128 , n13132 );
xor ( n13134 , n12801 , n12863 );
xor ( n13135 , n13134 , n12868 );
and ( n13136 , n13132 , n13135 );
and ( n13137 , n13128 , n13135 );
or ( n13138 , n13133 , n13136 , n13137 );
and ( n13139 , n11435 , n7601 );
and ( n13140 , n11383 , n7599 );
nor ( n13141 , n13139 , n13140 );
xnor ( n13142 , n13141 , n7611 );
and ( n13143 , n11817 , n7866 );
and ( n13144 , n11710 , n7864 );
nor ( n13145 , n13143 , n13144 );
xnor ( n13146 , n13145 , n7876 );
and ( n13147 , n13142 , n13146 );
and ( n13148 , n12246 , n7661 );
and ( n13149 , n12012 , n7659 );
nor ( n13150 , n13148 , n13149 );
xnor ( n13151 , n13150 , n7671 );
and ( n13152 , n13146 , n13151 );
and ( n13153 , n13142 , n13151 );
or ( n13154 , n13147 , n13152 , n13153 );
and ( n13155 , n11187 , n7713 );
and ( n13156 , n10554 , n7711 );
nor ( n13157 , n13155 , n13156 );
xnor ( n13158 , n13157 , n7723 );
and ( n13159 , n13154 , n13158 );
xor ( n13160 , n12775 , n12779 );
xor ( n13161 , n13160 , n12344 );
and ( n13162 , n13158 , n13161 );
and ( n13163 , n13154 , n13161 );
or ( n13164 , n13159 , n13162 , n13163 );
and ( n13165 , n10377 , n7542 );
and ( n13166 , n10239 , n7540 );
nor ( n13167 , n13165 , n13166 );
xnor ( n13168 , n13167 , n7552 );
and ( n13169 , n13164 , n13168 );
xor ( n13170 , n12771 , n12783 );
xor ( n13171 , n13170 , n12788 );
and ( n13172 , n13168 , n13171 );
and ( n13173 , n13164 , n13171 );
or ( n13174 , n13169 , n13172 , n13173 );
and ( n13175 , n8696 , n7781 );
and ( n13176 , n8429 , n7779 );
nor ( n13177 , n13175 , n13176 );
xnor ( n13178 , n13177 , n7791 );
and ( n13179 , n13174 , n13178 );
xor ( n13180 , n12843 , n12847 );
xor ( n13181 , n13180 , n12860 );
and ( n13182 , n13178 , n13181 );
and ( n13183 , n13174 , n13181 );
or ( n13184 , n13179 , n13182 , n13183 );
and ( n13185 , n7676 , n7395 );
and ( n13186 , n7696 , n7393 );
nor ( n13187 , n13185 , n13186 );
xnor ( n13188 , n13187 , n7405 );
and ( n13189 , n13184 , n13188 );
xor ( n13190 , n12965 , n12969 );
xor ( n13191 , n13190 , n12972 );
and ( n13192 , n13188 , n13191 );
and ( n13193 , n13184 , n13191 );
or ( n13194 , n13189 , n13192 , n13193 );
and ( n13195 , n13138 , n13194 );
xor ( n13196 , n12975 , n12979 );
xor ( n13197 , n13196 , n12982 );
and ( n13198 , n13194 , n13197 );
and ( n13199 , n13138 , n13197 );
or ( n13200 , n13195 , n13198 , n13199 );
and ( n13201 , n9049 , n7781 );
and ( n13202 , n8696 , n7779 );
nor ( n13203 , n13201 , n13202 );
xnor ( n13204 , n13203 , n7791 );
and ( n13205 , n10032 , n7501 );
and ( n13206 , n9829 , n7499 );
nor ( n13207 , n13205 , n13206 );
xnor ( n13208 , n13207 , n7511 );
and ( n13209 , n13204 , n13208 );
xor ( n13210 , n13164 , n13168 );
xor ( n13211 , n13210 , n13171 );
and ( n13212 , n13208 , n13211 );
and ( n13213 , n13204 , n13211 );
or ( n13214 , n13209 , n13212 , n13213 );
and ( n13215 , n8066 , n7899 );
and ( n13216 , n7851 , n7897 );
nor ( n13217 , n13215 , n13216 );
xnor ( n13218 , n13217 , n7909 );
and ( n13219 , n13214 , n13218 );
xor ( n13220 , n12955 , n12959 );
xor ( n13221 , n13220 , n12962 );
and ( n13222 , n13218 , n13221 );
and ( n13223 , n13214 , n13221 );
or ( n13224 , n13219 , n13222 , n13223 );
and ( n13225 , n7618 , n7318 );
and ( n13226 , n7666 , n7315 );
nor ( n13227 , n13225 , n13226 );
xnor ( n13228 , n13227 , n7311 );
and ( n13229 , n13224 , n13228 );
xor ( n13230 , n12989 , n12993 );
xor ( n13231 , n13230 , n12996 );
and ( n13232 , n13228 , n13231 );
and ( n13233 , n13224 , n13231 );
or ( n13234 , n13229 , n13232 , n13233 );
and ( n13235 , n7666 , n7318 );
and ( n13236 , n7871 , n7315 );
nor ( n13237 , n13235 , n13236 );
xnor ( n13238 , n13237 , n7311 );
and ( n13239 , n7809 , n8168 );
and ( n13240 , n7618 , n8166 );
nor ( n13241 , n13239 , n13240 );
xnor ( n13242 , n13241 , n8178 );
xor ( n13243 , n13238 , n13242 );
xor ( n13244 , n12871 , n12875 );
xor ( n13245 , n13244 , n12880 );
xor ( n13246 , n13243 , n13245 );
and ( n13247 , n13234 , n13246 );
xor ( n13248 , n12999 , n13003 );
xor ( n13249 , n13248 , n13006 );
and ( n13250 , n13246 , n13249 );
and ( n13251 , n13234 , n13249 );
or ( n13252 , n13247 , n13250 , n13251 );
and ( n13253 , n13200 , n13252 );
xor ( n13254 , n12985 , n13009 );
xor ( n13255 , n13254 , n13012 );
and ( n13256 , n13252 , n13255 );
and ( n13257 , n13200 , n13255 );
or ( n13258 , n13253 , n13256 , n13257 );
and ( n13259 , n13238 , n13242 );
and ( n13260 , n13242 , n13245 );
and ( n13261 , n13238 , n13245 );
or ( n13262 , n13259 , n13260 , n13261 );
xor ( n13263 , n12883 , n12887 );
xor ( n13264 , n13263 , n12890 );
and ( n13265 , n13262 , n13264 );
xor ( n13266 , n13019 , n13023 );
xor ( n13267 , n13266 , n13026 );
and ( n13268 , n13264 , n13267 );
and ( n13269 , n13262 , n13267 );
or ( n13270 , n13265 , n13268 , n13269 );
and ( n13271 , n13258 , n13270 );
xor ( n13272 , n13053 , n13055 );
xor ( n13273 , n13272 , n13058 );
and ( n13274 , n13270 , n13273 );
and ( n13275 , n13258 , n13273 );
or ( n13276 , n13271 , n13274 , n13275 );
and ( n13277 , n13075 , n13276 );
xor ( n13278 , n13075 , n13276 );
xor ( n13279 , n13258 , n13270 );
xor ( n13280 , n13279 , n13273 );
and ( n13281 , n11697 , n7601 );
and ( n13282 , n11569 , n7599 );
nor ( n13283 , n13281 , n13282 );
xnor ( n13284 , n13283 , n7611 );
and ( n13285 , n12246 , n7864 );
not ( n13286 , n13285 );
and ( n13287 , n13286 , n7876 );
and ( n13288 , n13284 , n13287 );
and ( n13289 , n11383 , n7713 );
and ( n13290 , n11249 , n7711 );
nor ( n13291 , n13289 , n13290 );
xnor ( n13292 , n13291 , n7723 );
and ( n13293 , n13288 , n13292 );
and ( n13294 , n12012 , n7866 );
and ( n13295 , n11817 , n7864 );
nor ( n13296 , n13294 , n13295 );
xnor ( n13297 , n13296 , n7876 );
and ( n13298 , n13292 , n13297 );
and ( n13299 , n13288 , n13297 );
or ( n13300 , n13293 , n13298 , n13299 );
and ( n13301 , n10554 , n7542 );
and ( n13302 , n10559 , n7540 );
nor ( n13303 , n13301 , n13302 );
xnor ( n13304 , n13303 , n7552 );
and ( n13305 , n13300 , n13304 );
xor ( n13306 , n13142 , n13146 );
xor ( n13307 , n13306 , n13151 );
and ( n13308 , n13304 , n13307 );
and ( n13309 , n13300 , n13307 );
or ( n13310 , n13305 , n13308 , n13309 );
and ( n13311 , n10239 , n7501 );
and ( n13312 , n10032 , n7499 );
nor ( n13313 , n13311 , n13312 );
xnor ( n13314 , n13313 , n7511 );
and ( n13315 , n13310 , n13314 );
xor ( n13316 , n13154 , n13158 );
xor ( n13317 , n13316 , n13161 );
and ( n13318 , n13314 , n13317 );
and ( n13319 , n13310 , n13317 );
or ( n13320 , n13315 , n13318 , n13319 );
and ( n13321 , n9463 , n7933 );
and ( n13322 , n9280 , n7931 );
nor ( n13323 , n13321 , n13322 );
xnor ( n13324 , n13323 , n7939 );
and ( n13325 , n9829 , n7954 );
and ( n13326 , n9701 , n7952 );
nor ( n13327 , n13325 , n13326 );
xnor ( n13328 , n13327 , n7964 );
and ( n13329 , n13324 , n13328 );
xor ( n13330 , n13096 , n13100 );
xor ( n13331 , n13330 , n13103 );
and ( n13332 , n13328 , n13331 );
and ( n13333 , n13324 , n13331 );
or ( n13334 , n13329 , n13332 , n13333 );
and ( n13335 , n13320 , n13334 );
and ( n13336 , n9280 , n7933 );
and ( n13337 , n9196 , n7931 );
nor ( n13338 , n13336 , n13337 );
xnor ( n13339 , n13338 , n7939 );
and ( n13340 , n13334 , n13339 );
and ( n13341 , n13320 , n13339 );
or ( n13342 , n13335 , n13340 , n13341 );
and ( n13343 , n7838 , n7395 );
and ( n13344 , n7676 , n7393 );
nor ( n13345 , n13343 , n13344 );
xnor ( n13346 , n13345 , n7405 );
and ( n13347 , n13342 , n13346 );
xor ( n13348 , n13174 , n13178 );
xor ( n13349 , n13348 , n13181 );
and ( n13350 , n13346 , n13349 );
and ( n13351 , n13342 , n13349 );
or ( n13352 , n13347 , n13350 , n13351 );
and ( n13353 , n7828 , n8168 );
and ( n13354 , n7809 , n8166 );
nor ( n13355 , n13353 , n13354 );
xnor ( n13356 , n13355 , n8178 );
and ( n13357 , n13352 , n13356 );
xor ( n13358 , n13184 , n13188 );
xor ( n13359 , n13358 , n13191 );
and ( n13360 , n13356 , n13359 );
and ( n13361 , n13352 , n13359 );
or ( n13362 , n13357 , n13360 , n13361 );
xor ( n13363 , n13138 , n13194 );
xor ( n13364 , n13363 , n13197 );
and ( n13365 , n13362 , n13364 );
xor ( n13366 , n13234 , n13246 );
xor ( n13367 , n13366 , n13249 );
and ( n13368 , n13364 , n13367 );
and ( n13369 , n13362 , n13367 );
or ( n13370 , n13365 , n13368 , n13369 );
xor ( n13371 , n13200 , n13252 );
xor ( n13372 , n13371 , n13255 );
and ( n13373 , n13370 , n13372 );
xor ( n13374 , n13262 , n13264 );
xor ( n13375 , n13374 , n13267 );
and ( n13376 , n13372 , n13375 );
and ( n13377 , n13370 , n13375 );
or ( n13378 , n13373 , n13376 , n13377 );
and ( n13379 , n13280 , n13378 );
xor ( n13380 , n13280 , n13378 );
xor ( n13381 , n13370 , n13372 );
xor ( n13382 , n13381 , n13375 );
and ( n13383 , n8079 , n7899 );
and ( n13384 , n8066 , n7897 );
nor ( n13385 , n13383 , n13384 );
xnor ( n13386 , n13385 , n7909 );
and ( n13387 , n8429 , n8044 );
and ( n13388 , n8263 , n8042 );
nor ( n13389 , n13387 , n13388 );
xnor ( n13390 , n13389 , n8054 );
and ( n13391 , n13386 , n13390 );
xor ( n13392 , n13106 , n13110 );
xor ( n13393 , n13392 , n13113 );
and ( n13394 , n13390 , n13393 );
and ( n13395 , n13386 , n13393 );
or ( n13396 , n13391 , n13394 , n13395 );
and ( n13397 , n7696 , n8168 );
and ( n13398 , n7828 , n8166 );
nor ( n13399 , n13397 , n13398 );
xnor ( n13400 , n13399 , n8178 );
and ( n13401 , n13396 , n13400 );
xor ( n13402 , n13116 , n13120 );
xor ( n13403 , n13402 , n13125 );
and ( n13404 , n13400 , n13403 );
and ( n13405 , n13396 , n13403 );
or ( n13406 , n13401 , n13404 , n13405 );
xor ( n13407 , n13128 , n13132 );
xor ( n13408 , n13407 , n13135 );
and ( n13409 , n13406 , n13408 );
xor ( n13410 , n13224 , n13228 );
xor ( n13411 , n13410 , n13231 );
and ( n13412 , n13408 , n13411 );
and ( n13413 , n13406 , n13411 );
or ( n13414 , n13409 , n13412 , n13413 );
and ( n13415 , n11435 , n7713 );
and ( n13416 , n11383 , n7711 );
nor ( n13417 , n13415 , n13416 );
xnor ( n13418 , n13417 , n7723 );
and ( n13419 , n11817 , n7743 );
and ( n13420 , n11710 , n7741 );
nor ( n13421 , n13419 , n13420 );
xnor ( n13422 , n13421 , n7753 );
and ( n13423 , n13418 , n13422 );
and ( n13424 , n12246 , n7866 );
and ( n13425 , n12012 , n7864 );
nor ( n13426 , n13424 , n13425 );
xnor ( n13427 , n13426 , n7876 );
and ( n13428 , n13422 , n13427 );
and ( n13429 , n13418 , n13427 );
or ( n13430 , n13423 , n13428 , n13429 );
and ( n13431 , n11187 , n7542 );
and ( n13432 , n10554 , n7540 );
nor ( n13433 , n13431 , n13432 );
xnor ( n13434 , n13433 , n7552 );
and ( n13435 , n13430 , n13434 );
xor ( n13436 , n13080 , n13084 );
xor ( n13437 , n13436 , n12806 );
and ( n13438 , n13434 , n13437 );
and ( n13439 , n13430 , n13437 );
or ( n13440 , n13435 , n13438 , n13439 );
and ( n13441 , n10377 , n7501 );
and ( n13442 , n10239 , n7499 );
nor ( n13443 , n13441 , n13442 );
xnor ( n13444 , n13443 , n7511 );
and ( n13445 , n13440 , n13444 );
xor ( n13446 , n13076 , n13088 );
xor ( n13447 , n13446 , n13093 );
and ( n13448 , n13444 , n13447 );
and ( n13449 , n13440 , n13447 );
or ( n13450 , n13445 , n13448 , n13449 );
and ( n13451 , n8696 , n8044 );
and ( n13452 , n8429 , n8042 );
nor ( n13453 , n13451 , n13452 );
xnor ( n13454 , n13453 , n8054 );
and ( n13455 , n13450 , n13454 );
xor ( n13456 , n13310 , n13314 );
xor ( n13457 , n13456 , n13317 );
and ( n13458 , n13454 , n13457 );
and ( n13459 , n13450 , n13457 );
or ( n13460 , n13455 , n13458 , n13459 );
and ( n13461 , n7851 , n7395 );
and ( n13462 , n7838 , n7393 );
nor ( n13463 , n13461 , n13462 );
xnor ( n13464 , n13463 , n7405 );
and ( n13465 , n13460 , n13464 );
xor ( n13466 , n13320 , n13334 );
xor ( n13467 , n13466 , n13339 );
and ( n13468 , n13464 , n13467 );
and ( n13469 , n13460 , n13467 );
or ( n13470 , n13465 , n13468 , n13469 );
and ( n13471 , n7809 , n7318 );
and ( n13472 , n7618 , n7315 );
nor ( n13473 , n13471 , n13472 );
xnor ( n13474 , n13473 , n7311 );
and ( n13475 , n13470 , n13474 );
xor ( n13476 , n13214 , n13218 );
xor ( n13477 , n13476 , n13221 );
and ( n13478 , n13474 , n13477 );
and ( n13479 , n13470 , n13477 );
or ( n13480 , n13475 , n13478 , n13479 );
xor ( n13481 , n13284 , n13287 );
and ( n13482 , n11569 , n7713 );
and ( n13483 , n11435 , n7711 );
nor ( n13484 , n13482 , n13483 );
xnor ( n13485 , n13484 , n7723 );
and ( n13486 , n12012 , n7743 );
and ( n13487 , n11817 , n7741 );
nor ( n13488 , n13486 , n13487 );
xnor ( n13489 , n13488 , n7753 );
and ( n13490 , n13485 , n13489 );
and ( n13491 , n13489 , n13285 );
and ( n13492 , n13485 , n13285 );
or ( n13493 , n13490 , n13491 , n13492 );
and ( n13494 , n13481 , n13493 );
and ( n13495 , n11249 , n7542 );
and ( n13496 , n11187 , n7540 );
nor ( n13497 , n13495 , n13496 );
xnor ( n13498 , n13497 , n7552 );
and ( n13499 , n13493 , n13498 );
and ( n13500 , n13481 , n13498 );
or ( n13501 , n13494 , n13499 , n13500 );
and ( n13502 , n10559 , n7501 );
and ( n13503 , n10377 , n7499 );
nor ( n13504 , n13502 , n13503 );
xnor ( n13505 , n13504 , n7511 );
and ( n13506 , n13501 , n13505 );
xor ( n13507 , n13288 , n13292 );
xor ( n13508 , n13507 , n13297 );
and ( n13509 , n13505 , n13508 );
and ( n13510 , n13501 , n13508 );
or ( n13511 , n13506 , n13509 , n13510 );
and ( n13512 , n10032 , n7954 );
and ( n13513 , n9829 , n7952 );
nor ( n13514 , n13512 , n13513 );
xnor ( n13515 , n13514 , n7964 );
and ( n13516 , n13511 , n13515 );
xor ( n13517 , n13300 , n13304 );
xor ( n13518 , n13517 , n13307 );
and ( n13519 , n13515 , n13518 );
and ( n13520 , n13511 , n13518 );
or ( n13521 , n13516 , n13519 , n13520 );
and ( n13522 , n8066 , n7395 );
and ( n13523 , n7851 , n7393 );
nor ( n13524 , n13522 , n13523 );
xnor ( n13525 , n13524 , n7405 );
and ( n13526 , n13521 , n13525 );
and ( n13527 , n9196 , n7781 );
and ( n13528 , n9049 , n7779 );
nor ( n13529 , n13527 , n13528 );
xnor ( n13530 , n13529 , n7791 );
and ( n13531 , n13525 , n13530 );
and ( n13532 , n13521 , n13530 );
or ( n13533 , n13526 , n13531 , n13532 );
and ( n13534 , n7676 , n8168 );
and ( n13535 , n7696 , n8166 );
nor ( n13536 , n13534 , n13535 );
xnor ( n13537 , n13536 , n8178 );
and ( n13538 , n13533 , n13537 );
xor ( n13539 , n13204 , n13208 );
xor ( n13540 , n13539 , n13211 );
and ( n13541 , n13537 , n13540 );
and ( n13542 , n13533 , n13540 );
or ( n13543 , n13538 , n13541 , n13542 );
xor ( n13544 , n13396 , n13400 );
xor ( n13545 , n13544 , n13403 );
and ( n13546 , n13543 , n13545 );
xor ( n13547 , n13342 , n13346 );
xor ( n13548 , n13547 , n13349 );
and ( n13549 , n13545 , n13548 );
and ( n13550 , n13543 , n13548 );
or ( n13551 , n13546 , n13549 , n13550 );
and ( n13552 , n13480 , n13551 );
xor ( n13553 , n13352 , n13356 );
xor ( n13554 , n13553 , n13359 );
and ( n13555 , n13551 , n13554 );
and ( n13556 , n13480 , n13554 );
or ( n13557 , n13552 , n13555 , n13556 );
and ( n13558 , n13414 , n13557 );
xor ( n13559 , n13362 , n13364 );
xor ( n13560 , n13559 , n13367 );
and ( n13561 , n13557 , n13560 );
and ( n13562 , n13414 , n13560 );
or ( n13563 , n13558 , n13561 , n13562 );
and ( n13564 , n13382 , n13563 );
xor ( n13565 , n13382 , n13563 );
and ( n13566 , n8079 , n7395 );
and ( n13567 , n8066 , n7393 );
nor ( n13568 , n13566 , n13567 );
xnor ( n13569 , n13568 , n7405 );
and ( n13570 , n8429 , n7899 );
and ( n13571 , n8263 , n7897 );
nor ( n13572 , n13570 , n13571 );
xnor ( n13573 , n13572 , n7909 );
and ( n13574 , n13569 , n13573 );
xor ( n13575 , n13511 , n13515 );
xor ( n13576 , n13575 , n13518 );
and ( n13577 , n13573 , n13576 );
and ( n13578 , n13569 , n13576 );
or ( n13579 , n13574 , n13577 , n13578 );
and ( n13580 , n7696 , n7318 );
and ( n13581 , n7828 , n7315 );
nor ( n13582 , n13580 , n13581 );
xnor ( n13583 , n13582 , n7311 );
and ( n13584 , n13579 , n13583 );
xor ( n13585 , n13521 , n13525 );
xor ( n13586 , n13585 , n13530 );
and ( n13587 , n13583 , n13586 );
and ( n13588 , n13579 , n13586 );
or ( n13589 , n13584 , n13587 , n13588 );
and ( n13590 , n9463 , n7781 );
and ( n13591 , n9280 , n7779 );
nor ( n13592 , n13590 , n13591 );
xnor ( n13593 , n13592 , n7791 );
and ( n13594 , n9829 , n7933 );
and ( n13595 , n9701 , n7931 );
nor ( n13596 , n13594 , n13595 );
xnor ( n13597 , n13596 , n7939 );
and ( n13598 , n13593 , n13597 );
xor ( n13599 , n13501 , n13505 );
xor ( n13600 , n13599 , n13508 );
and ( n13601 , n13597 , n13600 );
and ( n13602 , n13593 , n13600 );
or ( n13603 , n13598 , n13601 , n13602 );
and ( n13604 , n9049 , n8044 );
and ( n13605 , n8696 , n8042 );
nor ( n13606 , n13604 , n13605 );
xnor ( n13607 , n13606 , n8054 );
and ( n13608 , n13603 , n13607 );
and ( n13609 , n9280 , n7781 );
and ( n13610 , n9196 , n7779 );
nor ( n13611 , n13609 , n13610 );
xnor ( n13612 , n13611 , n7791 );
and ( n13613 , n13607 , n13612 );
and ( n13614 , n13603 , n13612 );
or ( n13615 , n13608 , n13613 , n13614 );
and ( n13616 , n7838 , n8168 );
and ( n13617 , n7676 , n8166 );
nor ( n13618 , n13616 , n13617 );
xnor ( n13619 , n13618 , n8178 );
and ( n13620 , n13615 , n13619 );
xor ( n13621 , n13450 , n13454 );
xor ( n13622 , n13621 , n13457 );
and ( n13623 , n13619 , n13622 );
and ( n13624 , n13615 , n13622 );
or ( n13625 , n13620 , n13623 , n13624 );
and ( n13626 , n13589 , n13625 );
xor ( n13627 , n13533 , n13537 );
xor ( n13628 , n13627 , n13540 );
and ( n13629 , n13625 , n13628 );
and ( n13630 , n13589 , n13628 );
or ( n13631 , n13626 , n13629 , n13630 );
and ( n13632 , n11697 , n7713 );
and ( n13633 , n11569 , n7711 );
nor ( n13634 , n13632 , n13633 );
xnor ( n13635 , n13634 , n7723 );
and ( n13636 , n12246 , n7741 );
not ( n13637 , n13636 );
and ( n13638 , n13637 , n7753 );
and ( n13639 , n13635 , n13638 );
and ( n13640 , n11383 , n7542 );
and ( n13641 , n11249 , n7540 );
nor ( n13642 , n13640 , n13641 );
xnor ( n13643 , n13642 , n7552 );
and ( n13644 , n13639 , n13643 );
and ( n13645 , n11710 , n7601 );
and ( n13646 , n11697 , n7599 );
nor ( n13647 , n13645 , n13646 );
xnor ( n13648 , n13647 , n7611 );
and ( n13649 , n13643 , n13648 );
and ( n13650 , n13639 , n13648 );
or ( n13651 , n13644 , n13649 , n13650 );
and ( n13652 , n10554 , n7501 );
and ( n13653 , n10559 , n7499 );
nor ( n13654 , n13652 , n13653 );
xnor ( n13655 , n13654 , n7511 );
and ( n13656 , n13651 , n13655 );
xor ( n13657 , n13418 , n13422 );
xor ( n13658 , n13657 , n13427 );
and ( n13659 , n13655 , n13658 );
and ( n13660 , n13651 , n13658 );
or ( n13661 , n13656 , n13659 , n13660 );
and ( n13662 , n10239 , n7954 );
and ( n13663 , n10032 , n7952 );
nor ( n13664 , n13662 , n13663 );
xnor ( n13665 , n13664 , n7964 );
and ( n13666 , n13661 , n13665 );
xor ( n13667 , n13430 , n13434 );
xor ( n13668 , n13667 , n13437 );
and ( n13669 , n13665 , n13668 );
and ( n13670 , n13661 , n13668 );
or ( n13671 , n13666 , n13669 , n13670 );
and ( n13672 , n9701 , n7933 );
and ( n13673 , n9463 , n7931 );
nor ( n13674 , n13672 , n13673 );
xnor ( n13675 , n13674 , n7939 );
and ( n13676 , n13671 , n13675 );
xor ( n13677 , n13440 , n13444 );
xor ( n13678 , n13677 , n13447 );
and ( n13679 , n13675 , n13678 );
and ( n13680 , n13671 , n13678 );
or ( n13681 , n13676 , n13679 , n13680 );
and ( n13682 , n8263 , n7899 );
and ( n13683 , n8079 , n7897 );
nor ( n13684 , n13682 , n13683 );
xnor ( n13685 , n13684 , n7909 );
and ( n13686 , n13681 , n13685 );
xor ( n13687 , n13324 , n13328 );
xor ( n13688 , n13687 , n13331 );
and ( n13689 , n13685 , n13688 );
and ( n13690 , n13681 , n13688 );
or ( n13691 , n13686 , n13689 , n13690 );
and ( n13692 , n7828 , n7318 );
and ( n13693 , n7809 , n7315 );
nor ( n13694 , n13692 , n13693 );
xnor ( n13695 , n13694 , n7311 );
and ( n13696 , n13691 , n13695 );
xor ( n13697 , n13386 , n13390 );
xor ( n13698 , n13697 , n13393 );
and ( n13699 , n13695 , n13698 );
and ( n13700 , n13691 , n13698 );
or ( n13701 , n13696 , n13699 , n13700 );
and ( n13702 , n13631 , n13701 );
xor ( n13703 , n13470 , n13474 );
xor ( n13704 , n13703 , n13477 );
and ( n13705 , n13701 , n13704 );
and ( n13706 , n13631 , n13704 );
or ( n13707 , n13702 , n13705 , n13706 );
xor ( n13708 , n13406 , n13408 );
xor ( n13709 , n13708 , n13411 );
and ( n13710 , n13707 , n13709 );
xor ( n13711 , n13480 , n13551 );
xor ( n13712 , n13711 , n13554 );
and ( n13713 , n13709 , n13712 );
and ( n13714 , n13707 , n13712 );
or ( n13715 , n13710 , n13713 , n13714 );
xor ( n13716 , n13414 , n13557 );
xor ( n13717 , n13716 , n13560 );
and ( n13718 , n13715 , n13717 );
xor ( n13719 , n13715 , n13717 );
xor ( n13720 , n13707 , n13709 );
xor ( n13721 , n13720 , n13712 );
and ( n13722 , n11435 , n7542 );
and ( n13723 , n11383 , n7540 );
nor ( n13724 , n13722 , n13723 );
xnor ( n13725 , n13724 , n7552 );
and ( n13726 , n11817 , n7601 );
and ( n13727 , n11710 , n7599 );
nor ( n13728 , n13726 , n13727 );
xnor ( n13729 , n13728 , n7611 );
and ( n13730 , n13725 , n13729 );
and ( n13731 , n12246 , n7743 );
and ( n13732 , n12012 , n7741 );
nor ( n13733 , n13731 , n13732 );
xnor ( n13734 , n13733 , n7753 );
and ( n13735 , n13729 , n13734 );
and ( n13736 , n13725 , n13734 );
or ( n13737 , n13730 , n13735 , n13736 );
and ( n13738 , n11187 , n7501 );
and ( n13739 , n10554 , n7499 );
nor ( n13740 , n13738 , n13739 );
xnor ( n13741 , n13740 , n7511 );
and ( n13742 , n13737 , n13741 );
xor ( n13743 , n13485 , n13489 );
xor ( n13744 , n13743 , n13285 );
and ( n13745 , n13741 , n13744 );
and ( n13746 , n13737 , n13744 );
or ( n13747 , n13742 , n13745 , n13746 );
and ( n13748 , n10377 , n7954 );
and ( n13749 , n10239 , n7952 );
nor ( n13750 , n13748 , n13749 );
xnor ( n13751 , n13750 , n7964 );
and ( n13752 , n13747 , n13751 );
xor ( n13753 , n13481 , n13493 );
xor ( n13754 , n13753 , n13498 );
and ( n13755 , n13751 , n13754 );
and ( n13756 , n13747 , n13754 );
or ( n13757 , n13752 , n13755 , n13756 );
and ( n13758 , n9196 , n8044 );
and ( n13759 , n9049 , n8042 );
nor ( n13760 , n13758 , n13759 );
xnor ( n13761 , n13760 , n8054 );
and ( n13762 , n13757 , n13761 );
xor ( n13763 , n13661 , n13665 );
xor ( n13764 , n13763 , n13668 );
and ( n13765 , n13761 , n13764 );
and ( n13766 , n13757 , n13764 );
or ( n13767 , n13762 , n13765 , n13766 );
xor ( n13768 , n13603 , n13607 );
xor ( n13769 , n13768 , n13612 );
and ( n13770 , n13767 , n13769 );
xor ( n13771 , n13671 , n13675 );
xor ( n13772 , n13771 , n13678 );
and ( n13773 , n13769 , n13772 );
and ( n13774 , n13767 , n13772 );
or ( n13775 , n13770 , n13773 , n13774 );
xor ( n13776 , n13681 , n13685 );
xor ( n13777 , n13776 , n13688 );
and ( n13778 , n13775 , n13777 );
xor ( n13779 , n13615 , n13619 );
xor ( n13780 , n13779 , n13622 );
and ( n13781 , n13777 , n13780 );
and ( n13782 , n13775 , n13780 );
or ( n13783 , n13778 , n13781 , n13782 );
xor ( n13784 , n13460 , n13464 );
xor ( n13785 , n13784 , n13467 );
and ( n13786 , n13783 , n13785 );
xor ( n13787 , n13691 , n13695 );
xor ( n13788 , n13787 , n13698 );
and ( n13789 , n13785 , n13788 );
and ( n13790 , n13783 , n13788 );
or ( n13791 , n13786 , n13789 , n13790 );
xor ( n13792 , n13543 , n13545 );
xor ( n13793 , n13792 , n13548 );
and ( n13794 , n13791 , n13793 );
xor ( n13795 , n13631 , n13701 );
xor ( n13796 , n13795 , n13704 );
and ( n13797 , n13793 , n13796 );
and ( n13798 , n13791 , n13796 );
or ( n13799 , n13794 , n13797 , n13798 );
and ( n13800 , n13721 , n13799 );
xor ( n13801 , n13721 , n13799 );
xor ( n13802 , n13791 , n13793 );
xor ( n13803 , n13802 , n13796 );
xor ( n13804 , n13635 , n13638 );
and ( n13805 , n11569 , n7542 );
and ( n13806 , n11435 , n7540 );
nor ( n13807 , n13805 , n13806 );
xnor ( n13808 , n13807 , n7552 );
and ( n13809 , n11710 , n7713 );
and ( n13810 , n11697 , n7711 );
nor ( n13811 , n13809 , n13810 );
xnor ( n13812 , n13811 , n7723 );
and ( n13813 , n13808 , n13812 );
and ( n13814 , n13812 , n13636 );
and ( n13815 , n13808 , n13636 );
or ( n13816 , n13813 , n13814 , n13815 );
and ( n13817 , n13804 , n13816 );
and ( n13818 , n11249 , n7501 );
and ( n13819 , n11187 , n7499 );
nor ( n13820 , n13818 , n13819 );
xnor ( n13821 , n13820 , n7511 );
and ( n13822 , n13816 , n13821 );
and ( n13823 , n13804 , n13821 );
or ( n13824 , n13817 , n13822 , n13823 );
and ( n13825 , n10559 , n7954 );
and ( n13826 , n10377 , n7952 );
nor ( n13827 , n13825 , n13826 );
xnor ( n13828 , n13827 , n7964 );
and ( n13829 , n13824 , n13828 );
xor ( n13830 , n13639 , n13643 );
xor ( n13831 , n13830 , n13648 );
and ( n13832 , n13828 , n13831 );
and ( n13833 , n13824 , n13831 );
or ( n13834 , n13829 , n13832 , n13833 );
and ( n13835 , n9701 , n7781 );
and ( n13836 , n9463 , n7779 );
nor ( n13837 , n13835 , n13836 );
xnor ( n13838 , n13837 , n7791 );
and ( n13839 , n13834 , n13838 );
xor ( n13840 , n13651 , n13655 );
xor ( n13841 , n13840 , n13658 );
and ( n13842 , n13838 , n13841 );
and ( n13843 , n13834 , n13841 );
or ( n13844 , n13839 , n13842 , n13843 );
and ( n13845 , n8066 , n8168 );
and ( n13846 , n7851 , n8166 );
nor ( n13847 , n13845 , n13846 );
xnor ( n13848 , n13847 , n8178 );
and ( n13849 , n13844 , n13848 );
and ( n13850 , n8696 , n7899 );
and ( n13851 , n8429 , n7897 );
nor ( n13852 , n13850 , n13851 );
xnor ( n13853 , n13852 , n7909 );
and ( n13854 , n13848 , n13853 );
and ( n13855 , n13844 , n13853 );
or ( n13856 , n13849 , n13854 , n13855 );
and ( n13857 , n7676 , n7318 );
and ( n13858 , n7696 , n7315 );
nor ( n13859 , n13857 , n13858 );
xnor ( n13860 , n13859 , n7311 );
and ( n13861 , n13856 , n13860 );
and ( n13862 , n7851 , n8168 );
and ( n13863 , n7838 , n8166 );
nor ( n13864 , n13862 , n13863 );
xnor ( n13865 , n13864 , n8178 );
and ( n13866 , n13860 , n13865 );
and ( n13867 , n13856 , n13865 );
or ( n13868 , n13861 , n13866 , n13867 );
and ( n13869 , n9280 , n8044 );
and ( n13870 , n9196 , n8042 );
nor ( n13871 , n13869 , n13870 );
xnor ( n13872 , n13871 , n8054 );
and ( n13873 , n10032 , n7933 );
and ( n13874 , n9829 , n7931 );
nor ( n13875 , n13873 , n13874 );
xnor ( n13876 , n13875 , n7939 );
and ( n13877 , n13872 , n13876 );
xor ( n13878 , n13747 , n13751 );
xor ( n13879 , n13878 , n13754 );
and ( n13880 , n13876 , n13879 );
and ( n13881 , n13872 , n13879 );
or ( n13882 , n13877 , n13880 , n13881 );
and ( n13883 , n8263 , n7395 );
and ( n13884 , n8079 , n7393 );
nor ( n13885 , n13883 , n13884 );
xnor ( n13886 , n13885 , n7405 );
and ( n13887 , n13882 , n13886 );
xor ( n13888 , n13593 , n13597 );
xor ( n13889 , n13888 , n13600 );
and ( n13890 , n13886 , n13889 );
and ( n13891 , n13882 , n13889 );
or ( n13892 , n13887 , n13890 , n13891 );
and ( n13893 , n11817 , n7713 );
and ( n13894 , n11710 , n7711 );
nor ( n13895 , n13893 , n13894 );
xnor ( n13896 , n13895 , n7723 );
and ( n13897 , n12246 , n7599 );
not ( n13898 , n13897 );
and ( n13899 , n13898 , n7611 );
and ( n13900 , n13896 , n13899 );
and ( n13901 , n11383 , n7501 );
and ( n13902 , n11249 , n7499 );
nor ( n13903 , n13901 , n13902 );
xnor ( n13904 , n13903 , n7511 );
and ( n13905 , n13900 , n13904 );
and ( n13906 , n12012 , n7601 );
and ( n13907 , n11817 , n7599 );
nor ( n13908 , n13906 , n13907 );
xnor ( n13909 , n13908 , n7611 );
and ( n13910 , n13904 , n13909 );
and ( n13911 , n13900 , n13909 );
or ( n13912 , n13905 , n13910 , n13911 );
and ( n13913 , n10554 , n7954 );
and ( n13914 , n10559 , n7952 );
nor ( n13915 , n13913 , n13914 );
xnor ( n13916 , n13915 , n7964 );
and ( n13917 , n13912 , n13916 );
xor ( n13918 , n13725 , n13729 );
xor ( n13919 , n13918 , n13734 );
and ( n13920 , n13916 , n13919 );
and ( n13921 , n13912 , n13919 );
or ( n13922 , n13917 , n13920 , n13921 );
and ( n13923 , n10239 , n7933 );
and ( n13924 , n10032 , n7931 );
nor ( n13925 , n13923 , n13924 );
xnor ( n13926 , n13925 , n7939 );
and ( n13927 , n13922 , n13926 );
xor ( n13928 , n13737 , n13741 );
xor ( n13929 , n13928 , n13744 );
and ( n13930 , n13926 , n13929 );
and ( n13931 , n13922 , n13929 );
or ( n13932 , n13927 , n13930 , n13931 );
and ( n13933 , n9463 , n8044 );
and ( n13934 , n9280 , n8042 );
nor ( n13935 , n13933 , n13934 );
xnor ( n13936 , n13935 , n8054 );
and ( n13937 , n9829 , n7781 );
and ( n13938 , n9701 , n7779 );
nor ( n13939 , n13937 , n13938 );
xnor ( n13940 , n13939 , n7791 );
and ( n13941 , n13936 , n13940 );
xor ( n13942 , n13824 , n13828 );
xor ( n13943 , n13942 , n13831 );
and ( n13944 , n13940 , n13943 );
and ( n13945 , n13936 , n13943 );
or ( n13946 , n13941 , n13944 , n13945 );
and ( n13947 , n13932 , n13946 );
and ( n13948 , n9049 , n7899 );
and ( n13949 , n8696 , n7897 );
nor ( n13950 , n13948 , n13949 );
xnor ( n13951 , n13950 , n7909 );
and ( n13952 , n13946 , n13951 );
and ( n13953 , n13932 , n13951 );
or ( n13954 , n13947 , n13952 , n13953 );
and ( n13955 , n7838 , n7318 );
and ( n13956 , n7676 , n7315 );
nor ( n13957 , n13955 , n13956 );
xnor ( n13958 , n13957 , n7311 );
and ( n13959 , n13954 , n13958 );
xor ( n13960 , n13757 , n13761 );
xor ( n13961 , n13960 , n13764 );
and ( n13962 , n13958 , n13961 );
and ( n13963 , n13954 , n13961 );
or ( n13964 , n13959 , n13962 , n13963 );
and ( n13965 , n13892 , n13964 );
xor ( n13966 , n13569 , n13573 );
xor ( n13967 , n13966 , n13576 );
and ( n13968 , n13964 , n13967 );
and ( n13969 , n13892 , n13967 );
or ( n13970 , n13965 , n13968 , n13969 );
and ( n13971 , n13868 , n13970 );
xor ( n13972 , n13579 , n13583 );
xor ( n13973 , n13972 , n13586 );
and ( n13974 , n13970 , n13973 );
and ( n13975 , n13868 , n13973 );
or ( n13976 , n13971 , n13974 , n13975 );
xor ( n13977 , n13589 , n13625 );
xor ( n13978 , n13977 , n13628 );
and ( n13979 , n13976 , n13978 );
xor ( n13980 , n13783 , n13785 );
xor ( n13981 , n13980 , n13788 );
and ( n13982 , n13978 , n13981 );
and ( n13983 , n13976 , n13981 );
or ( n13984 , n13979 , n13982 , n13983 );
and ( n13985 , n13803 , n13984 );
xor ( n13986 , n13803 , n13984 );
xor ( n13987 , n13976 , n13978 );
xor ( n13988 , n13987 , n13981 );
and ( n13989 , n8079 , n8168 );
and ( n13990 , n8066 , n8166 );
nor ( n13991 , n13989 , n13990 );
xnor ( n13992 , n13991 , n8178 );
and ( n13993 , n8429 , n7395 );
and ( n13994 , n8263 , n7393 );
nor ( n13995 , n13993 , n13994 );
xnor ( n13996 , n13995 , n7405 );
and ( n13997 , n13992 , n13996 );
xor ( n13998 , n13834 , n13838 );
xor ( n13999 , n13998 , n13841 );
and ( n14000 , n13996 , n13999 );
and ( n14001 , n13992 , n13999 );
or ( n14002 , n13997 , n14000 , n14001 );
xor ( n14003 , n13844 , n13848 );
xor ( n14004 , n14003 , n13853 );
and ( n14005 , n14002 , n14004 );
xor ( n14006 , n13882 , n13886 );
xor ( n14007 , n14006 , n13889 );
and ( n14008 , n14004 , n14007 );
and ( n14009 , n14002 , n14007 );
or ( n14010 , n14005 , n14008 , n14009 );
xor ( n14011 , n13856 , n13860 );
xor ( n14012 , n14011 , n13865 );
and ( n14013 , n14010 , n14012 );
xor ( n14014 , n13767 , n13769 );
xor ( n14015 , n14014 , n13772 );
and ( n14016 , n14012 , n14015 );
and ( n14017 , n14010 , n14015 );
or ( n14018 , n14013 , n14016 , n14017 );
xor ( n14019 , n13868 , n13970 );
xor ( n14020 , n14019 , n13973 );
and ( n14021 , n14018 , n14020 );
xor ( n14022 , n13775 , n13777 );
xor ( n14023 , n14022 , n13780 );
and ( n14024 , n14020 , n14023 );
and ( n14025 , n14018 , n14023 );
or ( n14026 , n14021 , n14024 , n14025 );
and ( n14027 , n13988 , n14026 );
xor ( n14028 , n13988 , n14026 );
xor ( n14029 , n14018 , n14020 );
xor ( n14030 , n14029 , n14023 );
and ( n14031 , n11697 , n7501 );
and ( n14032 , n11569 , n7499 );
nor ( n14033 , n14031 , n14032 );
xnor ( n14034 , n14033 , n7511 );
and ( n14035 , n12246 , n7711 );
not ( n14036 , n14035 );
and ( n14037 , n14036 , n7723 );
and ( n14038 , n14034 , n14037 );
and ( n14039 , n11383 , n7954 );
and ( n14040 , n11249 , n7952 );
nor ( n14041 , n14039 , n14040 );
xnor ( n14042 , n14041 , n7964 );
and ( n14043 , n14038 , n14042 );
and ( n14044 , n11569 , n7501 );
and ( n14045 , n11435 , n7499 );
nor ( n14046 , n14044 , n14045 );
xnor ( n14047 , n14046 , n7511 );
and ( n14048 , n14042 , n14047 );
and ( n14049 , n14038 , n14047 );
or ( n14050 , n14043 , n14048 , n14049 );
and ( n14051 , n10554 , n7933 );
and ( n14052 , n10559 , n7931 );
nor ( n14053 , n14051 , n14052 );
xnor ( n14054 , n14053 , n7939 );
and ( n14055 , n14050 , n14054 );
and ( n14056 , n11435 , n7501 );
and ( n14057 , n11383 , n7499 );
nor ( n14058 , n14056 , n14057 );
xnor ( n14059 , n14058 , n7511 );
and ( n14060 , n11697 , n7542 );
and ( n14061 , n11569 , n7540 );
nor ( n14062 , n14060 , n14061 );
xnor ( n14063 , n14062 , n7552 );
xor ( n14064 , n14059 , n14063 );
and ( n14065 , n12246 , n7601 );
and ( n14066 , n12012 , n7599 );
nor ( n14067 , n14065 , n14066 );
xnor ( n14068 , n14067 , n7611 );
xor ( n14069 , n14064 , n14068 );
and ( n14070 , n14054 , n14069 );
and ( n14071 , n14050 , n14069 );
or ( n14072 , n14055 , n14070 , n14071 );
and ( n14073 , n10239 , n7781 );
and ( n14074 , n10032 , n7779 );
nor ( n14075 , n14073 , n14074 );
xnor ( n14076 , n14075 , n7791 );
and ( n14077 , n14072 , n14076 );
and ( n14078 , n14059 , n14063 );
and ( n14079 , n14063 , n14068 );
and ( n14080 , n14059 , n14068 );
or ( n14081 , n14078 , n14079 , n14080 );
and ( n14082 , n11187 , n7954 );
and ( n14083 , n10554 , n7952 );
nor ( n14084 , n14082 , n14083 );
xnor ( n14085 , n14084 , n7964 );
xor ( n14086 , n14081 , n14085 );
xor ( n14087 , n13808 , n13812 );
xor ( n14088 , n14087 , n13636 );
xor ( n14089 , n14086 , n14088 );
and ( n14090 , n14076 , n14089 );
and ( n14091 , n14072 , n14089 );
or ( n14092 , n14077 , n14090 , n14091 );
and ( n14093 , n10032 , n7781 );
and ( n14094 , n9829 , n7779 );
nor ( n14095 , n14093 , n14094 );
xnor ( n14096 , n14095 , n7791 );
and ( n14097 , n14092 , n14096 );
and ( n14098 , n14081 , n14085 );
and ( n14099 , n14085 , n14088 );
and ( n14100 , n14081 , n14088 );
or ( n14101 , n14098 , n14099 , n14100 );
and ( n14102 , n10377 , n7933 );
and ( n14103 , n10239 , n7931 );
nor ( n14104 , n14102 , n14103 );
xnor ( n14105 , n14104 , n7939 );
xor ( n14106 , n14101 , n14105 );
xor ( n14107 , n13804 , n13816 );
xor ( n14108 , n14107 , n13821 );
xor ( n14109 , n14106 , n14108 );
and ( n14110 , n14096 , n14109 );
and ( n14111 , n14092 , n14109 );
or ( n14112 , n14097 , n14110 , n14111 );
and ( n14113 , n8066 , n7318 );
and ( n14114 , n7851 , n7315 );
nor ( n14115 , n14113 , n14114 );
xnor ( n14116 , n14115 , n7311 );
and ( n14117 , n14112 , n14116 );
and ( n14118 , n8263 , n8168 );
and ( n14119 , n8079 , n8166 );
nor ( n14120 , n14118 , n14119 );
xnor ( n14121 , n14120 , n8178 );
and ( n14122 , n14116 , n14121 );
and ( n14123 , n14112 , n14121 );
or ( n14124 , n14117 , n14122 , n14123 );
xor ( n14125 , n13896 , n13899 );
and ( n14126 , n11710 , n7542 );
and ( n14127 , n11697 , n7540 );
nor ( n14128 , n14126 , n14127 );
xnor ( n14129 , n14128 , n7552 );
and ( n14130 , n12012 , n7713 );
and ( n14131 , n11817 , n7711 );
nor ( n14132 , n14130 , n14131 );
xnor ( n14133 , n14132 , n7723 );
and ( n14134 , n14129 , n14133 );
and ( n14135 , n14133 , n13897 );
and ( n14136 , n14129 , n13897 );
or ( n14137 , n14134 , n14135 , n14136 );
and ( n14138 , n14125 , n14137 );
and ( n14139 , n11249 , n7954 );
and ( n14140 , n11187 , n7952 );
nor ( n14141 , n14139 , n14140 );
xnor ( n14142 , n14141 , n7964 );
and ( n14143 , n14137 , n14142 );
and ( n14144 , n14125 , n14142 );
or ( n14145 , n14138 , n14143 , n14144 );
and ( n14146 , n10559 , n7933 );
and ( n14147 , n10377 , n7931 );
nor ( n14148 , n14146 , n14147 );
xnor ( n14149 , n14148 , n7939 );
and ( n14150 , n14145 , n14149 );
xor ( n14151 , n13900 , n13904 );
xor ( n14152 , n14151 , n13909 );
and ( n14153 , n14149 , n14152 );
and ( n14154 , n14145 , n14152 );
or ( n14155 , n14150 , n14153 , n14154 );
and ( n14156 , n9701 , n8044 );
and ( n14157 , n9463 , n8042 );
nor ( n14158 , n14156 , n14157 );
xnor ( n14159 , n14158 , n8054 );
and ( n14160 , n14155 , n14159 );
xor ( n14161 , n13912 , n13916 );
xor ( n14162 , n14161 , n13919 );
and ( n14163 , n14159 , n14162 );
and ( n14164 , n14155 , n14162 );
or ( n14165 , n14160 , n14163 , n14164 );
and ( n14166 , n9196 , n7899 );
and ( n14167 , n9049 , n7897 );
nor ( n14168 , n14166 , n14167 );
xnor ( n14169 , n14168 , n7909 );
and ( n14170 , n14165 , n14169 );
xor ( n14171 , n13936 , n13940 );
xor ( n14172 , n14171 , n13943 );
and ( n14173 , n14169 , n14172 );
and ( n14174 , n14165 , n14172 );
or ( n14175 , n14170 , n14173 , n14174 );
and ( n14176 , n14124 , n14175 );
and ( n14177 , n7851 , n7318 );
and ( n14178 , n7838 , n7315 );
nor ( n14179 , n14177 , n14178 );
xnor ( n14180 , n14179 , n7311 );
and ( n14181 , n14175 , n14180 );
and ( n14182 , n14124 , n14180 );
or ( n14183 , n14176 , n14181 , n14182 );
and ( n14184 , n14101 , n14105 );
and ( n14185 , n14105 , n14108 );
and ( n14186 , n14101 , n14108 );
or ( n14187 , n14184 , n14185 , n14186 );
and ( n14188 , n8696 , n7395 );
and ( n14189 , n8429 , n7393 );
nor ( n14190 , n14188 , n14189 );
xnor ( n14191 , n14190 , n7405 );
and ( n14192 , n14187 , n14191 );
xor ( n14193 , n13922 , n13926 );
xor ( n14194 , n14193 , n13929 );
and ( n14195 , n14191 , n14194 );
and ( n14196 , n14187 , n14194 );
or ( n14197 , n14192 , n14195 , n14196 );
xor ( n14198 , n13932 , n13946 );
xor ( n14199 , n14198 , n13951 );
and ( n14200 , n14197 , n14199 );
xor ( n14201 , n13872 , n13876 );
xor ( n14202 , n14201 , n13879 );
and ( n14203 , n14199 , n14202 );
and ( n14204 , n14197 , n14202 );
or ( n14205 , n14200 , n14203 , n14204 );
and ( n14206 , n14183 , n14205 );
xor ( n14207 , n13954 , n13958 );
xor ( n14208 , n14207 , n13961 );
and ( n14209 , n14205 , n14208 );
and ( n14210 , n14183 , n14208 );
or ( n14211 , n14206 , n14209 , n14210 );
xor ( n14212 , n13892 , n13964 );
xor ( n14213 , n14212 , n13967 );
and ( n14214 , n14211 , n14213 );
xor ( n14215 , n14010 , n14012 );
xor ( n14216 , n14215 , n14015 );
and ( n14217 , n14213 , n14216 );
and ( n14218 , n14211 , n14216 );
or ( n14219 , n14214 , n14217 , n14218 );
and ( n14220 , n14030 , n14219 );
xor ( n14221 , n14030 , n14219 );
xor ( n14222 , n14211 , n14213 );
xor ( n14223 , n14222 , n14216 );
and ( n14224 , n9463 , n7899 );
and ( n14225 , n9280 , n7897 );
nor ( n14226 , n14224 , n14225 );
xnor ( n14227 , n14226 , n7909 );
and ( n14228 , n9829 , n8044 );
and ( n14229 , n9701 , n8042 );
nor ( n14230 , n14228 , n14229 );
xnor ( n14231 , n14230 , n8054 );
and ( n14232 , n14227 , n14231 );
xor ( n14233 , n14145 , n14149 );
xor ( n14234 , n14233 , n14152 );
and ( n14235 , n14231 , n14234 );
and ( n14236 , n14227 , n14234 );
or ( n14237 , n14232 , n14235 , n14236 );
and ( n14238 , n9049 , n7395 );
and ( n14239 , n8696 , n7393 );
nor ( n14240 , n14238 , n14239 );
xnor ( n14241 , n14240 , n7405 );
and ( n14242 , n14237 , n14241 );
and ( n14243 , n9280 , n7899 );
and ( n14244 , n9196 , n7897 );
nor ( n14245 , n14243 , n14244 );
xnor ( n14246 , n14245 , n7909 );
and ( n14247 , n14241 , n14246 );
and ( n14248 , n14237 , n14246 );
or ( n14249 , n14242 , n14247 , n14248 );
and ( n14250 , n8079 , n7318 );
and ( n14251 , n8066 , n7315 );
nor ( n14252 , n14250 , n14251 );
xnor ( n14253 , n14252 , n7311 );
and ( n14254 , n8429 , n8168 );
and ( n14255 , n8263 , n8166 );
nor ( n14256 , n14254 , n14255 );
xnor ( n14257 , n14256 , n8178 );
and ( n14258 , n14253 , n14257 );
xor ( n14259 , n14155 , n14159 );
xor ( n14260 , n14259 , n14162 );
and ( n14261 , n14257 , n14260 );
and ( n14262 , n14253 , n14260 );
or ( n14263 , n14258 , n14261 , n14262 );
and ( n14264 , n14249 , n14263 );
xor ( n14265 , n14187 , n14191 );
xor ( n14266 , n14265 , n14194 );
and ( n14267 , n14263 , n14266 );
and ( n14268 , n14249 , n14266 );
or ( n14269 , n14264 , n14267 , n14268 );
xor ( n14270 , n13992 , n13996 );
xor ( n14271 , n14270 , n13999 );
and ( n14272 , n14269 , n14271 );
xor ( n14273 , n14197 , n14199 );
xor ( n14274 , n14273 , n14202 );
and ( n14275 , n14271 , n14274 );
and ( n14276 , n14269 , n14274 );
or ( n14277 , n14272 , n14275 , n14276 );
xor ( n14278 , n14002 , n14004 );
xor ( n14279 , n14278 , n14007 );
and ( n14280 , n14277 , n14279 );
xor ( n14281 , n14183 , n14205 );
xor ( n14282 , n14281 , n14208 );
and ( n14283 , n14279 , n14282 );
and ( n14284 , n14277 , n14282 );
or ( n14285 , n14280 , n14283 , n14284 );
and ( n14286 , n14223 , n14285 );
xor ( n14287 , n14223 , n14285 );
xor ( n14288 , n14277 , n14279 );
xor ( n14289 , n14288 , n14282 );
xor ( n14290 , n14034 , n14037 );
and ( n14291 , n11817 , n7542 );
and ( n14292 , n11710 , n7540 );
nor ( n14293 , n14291 , n14292 );
xnor ( n14294 , n14293 , n7552 );
and ( n14295 , n14290 , n14294 );
and ( n14296 , n12246 , n7713 );
and ( n14297 , n12012 , n7711 );
nor ( n14298 , n14296 , n14297 );
xnor ( n14299 , n14298 , n7723 );
and ( n14300 , n14294 , n14299 );
and ( n14301 , n14290 , n14299 );
or ( n14302 , n14295 , n14300 , n14301 );
and ( n14303 , n11187 , n7933 );
and ( n14304 , n10554 , n7931 );
nor ( n14305 , n14303 , n14304 );
xnor ( n14306 , n14305 , n7939 );
and ( n14307 , n14302 , n14306 );
xor ( n14308 , n14129 , n14133 );
xor ( n14309 , n14308 , n13897 );
and ( n14310 , n14306 , n14309 );
and ( n14311 , n14302 , n14309 );
or ( n14312 , n14307 , n14310 , n14311 );
and ( n14313 , n11569 , n7954 );
and ( n14314 , n11435 , n7952 );
nor ( n14315 , n14313 , n14314 );
xnor ( n14316 , n14315 , n7964 );
and ( n14317 , n11710 , n7501 );
and ( n14318 , n11697 , n7499 );
nor ( n14319 , n14317 , n14318 );
xnor ( n14320 , n14319 , n7511 );
and ( n14321 , n14316 , n14320 );
and ( n14322 , n14320 , n14035 );
and ( n14323 , n14316 , n14035 );
or ( n14324 , n14321 , n14322 , n14323 );
and ( n14325 , n11435 , n7954 );
and ( n14326 , n11383 , n7952 );
nor ( n14327 , n14325 , n14326 );
xnor ( n14328 , n14327 , n7964 );
and ( n14329 , n14324 , n14328 );
xor ( n14330 , n14290 , n14294 );
xor ( n14331 , n14330 , n14299 );
and ( n14332 , n14328 , n14331 );
and ( n14333 , n14324 , n14331 );
or ( n14334 , n14329 , n14332 , n14333 );
xor ( n14335 , n14038 , n14042 );
xor ( n14336 , n14335 , n14047 );
and ( n14337 , n14334 , n14336 );
xor ( n14338 , n14302 , n14306 );
xor ( n14339 , n14338 , n14309 );
and ( n14340 , n14336 , n14339 );
and ( n14341 , n14334 , n14339 );
or ( n14342 , n14337 , n14340 , n14341 );
and ( n14343 , n14312 , n14342 );
xor ( n14344 , n14125 , n14137 );
xor ( n14345 , n14344 , n14142 );
and ( n14346 , n14342 , n14345 );
and ( n14347 , n14312 , n14345 );
or ( n14348 , n14343 , n14346 , n14347 );
and ( n14349 , n8696 , n8168 );
and ( n14350 , n8429 , n8166 );
nor ( n14351 , n14349 , n14350 );
xnor ( n14352 , n14351 , n8178 );
and ( n14353 , n14348 , n14352 );
and ( n14354 , n9196 , n7395 );
and ( n14355 , n9049 , n7393 );
nor ( n14356 , n14354 , n14355 );
xnor ( n14357 , n14356 , n7405 );
and ( n14358 , n14352 , n14357 );
and ( n14359 , n14348 , n14357 );
or ( n14360 , n14353 , n14358 , n14359 );
xor ( n14361 , n14237 , n14241 );
xor ( n14362 , n14361 , n14246 );
and ( n14363 , n14360 , n14362 );
xor ( n14364 , n14092 , n14096 );
xor ( n14365 , n14364 , n14109 );
and ( n14366 , n14362 , n14365 );
and ( n14367 , n14360 , n14365 );
or ( n14368 , n14363 , n14366 , n14367 );
xor ( n14369 , n14112 , n14116 );
xor ( n14370 , n14369 , n14121 );
and ( n14371 , n14368 , n14370 );
xor ( n14372 , n14165 , n14169 );
xor ( n14373 , n14372 , n14172 );
and ( n14374 , n14370 , n14373 );
and ( n14375 , n14368 , n14373 );
or ( n14376 , n14371 , n14374 , n14375 );
xor ( n14377 , n14124 , n14175 );
xor ( n14378 , n14377 , n14180 );
and ( n14379 , n14376 , n14378 );
xor ( n14380 , n14269 , n14271 );
xor ( n14381 , n14380 , n14274 );
and ( n14382 , n14378 , n14381 );
and ( n14383 , n14376 , n14381 );
or ( n14384 , n14379 , n14382 , n14383 );
and ( n14385 , n14289 , n14384 );
xor ( n14386 , n14289 , n14384 );
xor ( n14387 , n14376 , n14378 );
xor ( n14388 , n14387 , n14381 );
and ( n14389 , n9049 , n8168 );
and ( n14390 , n8696 , n8166 );
nor ( n14391 , n14389 , n14390 );
xnor ( n14392 , n14391 , n8178 );
and ( n14393 , n9280 , n7395 );
and ( n14394 , n9196 , n7393 );
nor ( n14395 , n14393 , n14394 );
xnor ( n14396 , n14395 , n7405 );
and ( n14397 , n14392 , n14396 );
and ( n14398 , n9701 , n7899 );
and ( n14399 , n9463 , n7897 );
nor ( n14400 , n14398 , n14399 );
xnor ( n14401 , n14400 , n7909 );
and ( n14402 , n14396 , n14401 );
and ( n14403 , n14392 , n14401 );
or ( n14404 , n14397 , n14402 , n14403 );
and ( n14405 , n11697 , n7954 );
and ( n14406 , n11569 , n7952 );
nor ( n14407 , n14405 , n14406 );
xnor ( n14408 , n14407 , n7964 );
and ( n14409 , n12246 , n7540 );
not ( n14410 , n14409 );
and ( n14411 , n14410 , n7552 );
and ( n14412 , n14408 , n14411 );
and ( n14413 , n12012 , n7542 );
and ( n14414 , n11817 , n7540 );
nor ( n14415 , n14413 , n14414 );
xnor ( n14416 , n14415 , n7552 );
and ( n14417 , n14412 , n14416 );
xor ( n14418 , n14316 , n14320 );
xor ( n14419 , n14418 , n14035 );
and ( n14420 , n14416 , n14419 );
and ( n14421 , n14412 , n14419 );
or ( n14422 , n14417 , n14420 , n14421 );
and ( n14423 , n11249 , n7933 );
and ( n14424 , n11187 , n7931 );
nor ( n14425 , n14423 , n14424 );
xnor ( n14426 , n14425 , n7939 );
and ( n14427 , n14422 , n14426 );
xor ( n14428 , n14324 , n14328 );
xor ( n14429 , n14428 , n14331 );
and ( n14430 , n14426 , n14429 );
and ( n14431 , n14422 , n14429 );
or ( n14432 , n14427 , n14430 , n14431 );
and ( n14433 , n10239 , n8044 );
and ( n14434 , n10032 , n8042 );
nor ( n14435 , n14433 , n14434 );
xnor ( n14436 , n14435 , n8054 );
and ( n14437 , n14432 , n14436 );
and ( n14438 , n10559 , n7781 );
and ( n14439 , n10377 , n7779 );
nor ( n14440 , n14438 , n14439 );
xnor ( n14441 , n14440 , n7791 );
and ( n14442 , n14436 , n14441 );
and ( n14443 , n14432 , n14441 );
or ( n14444 , n14437 , n14442 , n14443 );
xor ( n14445 , n14312 , n14342 );
xor ( n14446 , n14445 , n14345 );
and ( n14447 , n14444 , n14446 );
and ( n14448 , n10032 , n8044 );
and ( n14449 , n9829 , n8042 );
nor ( n14450 , n14448 , n14449 );
xnor ( n14451 , n14450 , n8054 );
and ( n14452 , n10377 , n7781 );
and ( n14453 , n10239 , n7779 );
nor ( n14454 , n14452 , n14453 );
xnor ( n14455 , n14454 , n7791 );
xor ( n14456 , n14451 , n14455 );
xor ( n14457 , n14050 , n14054 );
xor ( n14458 , n14457 , n14069 );
xor ( n14459 , n14456 , n14458 );
and ( n14460 , n14446 , n14459 );
and ( n14461 , n14444 , n14459 );
or ( n14462 , n14447 , n14460 , n14461 );
and ( n14463 , n14404 , n14462 );
and ( n14464 , n8263 , n7318 );
and ( n14465 , n8079 , n7315 );
nor ( n14466 , n14464 , n14465 );
xnor ( n14467 , n14466 , n7311 );
and ( n14468 , n14462 , n14467 );
and ( n14469 , n14404 , n14467 );
or ( n14470 , n14463 , n14468 , n14469 );
and ( n14471 , n14451 , n14455 );
and ( n14472 , n14455 , n14458 );
and ( n14473 , n14451 , n14458 );
or ( n14474 , n14471 , n14472 , n14473 );
xor ( n14475 , n14072 , n14076 );
xor ( n14476 , n14475 , n14089 );
and ( n14477 , n14474 , n14476 );
xor ( n14478 , n14227 , n14231 );
xor ( n14479 , n14478 , n14234 );
and ( n14480 , n14476 , n14479 );
and ( n14481 , n14474 , n14479 );
or ( n14482 , n14477 , n14480 , n14481 );
and ( n14483 , n14470 , n14482 );
xor ( n14484 , n14253 , n14257 );
xor ( n14485 , n14484 , n14260 );
and ( n14486 , n14482 , n14485 );
and ( n14487 , n14470 , n14485 );
or ( n14488 , n14483 , n14486 , n14487 );
xor ( n14489 , n14249 , n14263 );
xor ( n14490 , n14489 , n14266 );
and ( n14491 , n14488 , n14490 );
xor ( n14492 , n14368 , n14370 );
xor ( n14493 , n14492 , n14373 );
and ( n14494 , n14490 , n14493 );
and ( n14495 , n14488 , n14493 );
or ( n14496 , n14491 , n14494 , n14495 );
and ( n14497 , n14388 , n14496 );
xor ( n14498 , n14388 , n14496 );
xor ( n14499 , n14488 , n14490 );
xor ( n14500 , n14499 , n14493 );
xor ( n14501 , n14408 , n14411 );
and ( n14502 , n11817 , n7501 );
and ( n14503 , n11710 , n7499 );
nor ( n14504 , n14502 , n14503 );
xnor ( n14505 , n14504 , n7511 );
and ( n14506 , n14501 , n14505 );
and ( n14507 , n12246 , n7542 );
and ( n14508 , n12012 , n7540 );
nor ( n14509 , n14507 , n14508 );
xnor ( n14510 , n14509 , n7552 );
and ( n14511 , n14505 , n14510 );
and ( n14512 , n14501 , n14510 );
or ( n14513 , n14506 , n14511 , n14512 );
and ( n14514 , n11187 , n7781 );
and ( n14515 , n10554 , n7779 );
nor ( n14516 , n14514 , n14515 );
xnor ( n14517 , n14516 , n7791 );
and ( n14518 , n14513 , n14517 );
and ( n14519 , n11383 , n7933 );
and ( n14520 , n11249 , n7931 );
nor ( n14521 , n14519 , n14520 );
xnor ( n14522 , n14521 , n7939 );
and ( n14523 , n14517 , n14522 );
and ( n14524 , n14513 , n14522 );
or ( n14525 , n14518 , n14523 , n14524 );
and ( n14526 , n10554 , n7781 );
and ( n14527 , n10559 , n7779 );
nor ( n14528 , n14526 , n14527 );
xnor ( n14529 , n14528 , n7791 );
and ( n14530 , n14525 , n14529 );
xor ( n14531 , n14422 , n14426 );
xor ( n14532 , n14531 , n14429 );
and ( n14533 , n14529 , n14532 );
and ( n14534 , n14525 , n14532 );
or ( n14535 , n14530 , n14533 , n14534 );
and ( n14536 , n8696 , n7318 );
and ( n14537 , n8429 , n7315 );
nor ( n14538 , n14536 , n14537 );
xnor ( n14539 , n14538 , n7311 );
and ( n14540 , n14535 , n14539 );
xor ( n14541 , n14432 , n14436 );
xor ( n14542 , n14541 , n14441 );
and ( n14543 , n14539 , n14542 );
and ( n14544 , n14535 , n14542 );
or ( n14545 , n14540 , n14543 , n14544 );
and ( n14546 , n9463 , n7395 );
and ( n14547 , n9280 , n7393 );
nor ( n14548 , n14546 , n14547 );
xnor ( n14549 , n14548 , n7405 );
and ( n14550 , n9829 , n7899 );
and ( n14551 , n9701 , n7897 );
nor ( n14552 , n14550 , n14551 );
xnor ( n14553 , n14552 , n7909 );
and ( n14554 , n14549 , n14553 );
xor ( n14555 , n14334 , n14336 );
xor ( n14556 , n14555 , n14339 );
and ( n14557 , n14553 , n14556 );
and ( n14558 , n14549 , n14556 );
or ( n14559 , n14554 , n14557 , n14558 );
and ( n14560 , n14545 , n14559 );
and ( n14561 , n8429 , n7318 );
and ( n14562 , n8263 , n7315 );
nor ( n14563 , n14561 , n14562 );
xnor ( n14564 , n14563 , n7311 );
and ( n14565 , n14559 , n14564 );
and ( n14566 , n14545 , n14564 );
or ( n14567 , n14560 , n14565 , n14566 );
xor ( n14568 , n14348 , n14352 );
xor ( n14569 , n14568 , n14357 );
and ( n14570 , n14567 , n14569 );
xor ( n14571 , n14474 , n14476 );
xor ( n14572 , n14571 , n14479 );
and ( n14573 , n14569 , n14572 );
and ( n14574 , n14567 , n14572 );
or ( n14575 , n14570 , n14573 , n14574 );
xor ( n14576 , n14360 , n14362 );
xor ( n14577 , n14576 , n14365 );
and ( n14578 , n14575 , n14577 );
xor ( n14579 , n14470 , n14482 );
xor ( n14580 , n14579 , n14485 );
and ( n14581 , n14577 , n14580 );
and ( n14582 , n14575 , n14580 );
or ( n14583 , n14578 , n14581 , n14582 );
and ( n14584 , n14500 , n14583 );
xor ( n14585 , n14500 , n14583 );
xor ( n14586 , n14575 , n14577 );
xor ( n14587 , n14586 , n14580 );
and ( n14588 , n11710 , n7954 );
and ( n14589 , n11697 , n7952 );
nor ( n14590 , n14588 , n14589 );
xnor ( n14591 , n14590 , n7964 );
and ( n14592 , n12012 , n7501 );
and ( n14593 , n11817 , n7499 );
nor ( n14594 , n14592 , n14593 );
xnor ( n14595 , n14594 , n7511 );
and ( n14596 , n14591 , n14595 );
and ( n14597 , n14595 , n14409 );
and ( n14598 , n14591 , n14409 );
or ( n14599 , n14596 , n14597 , n14598 );
and ( n14600 , n11435 , n7933 );
and ( n14601 , n11383 , n7931 );
nor ( n14602 , n14600 , n14601 );
xnor ( n14603 , n14602 , n7939 );
and ( n14604 , n14599 , n14603 );
xor ( n14605 , n14501 , n14505 );
xor ( n14606 , n14605 , n14510 );
and ( n14607 , n14603 , n14606 );
and ( n14608 , n14599 , n14606 );
or ( n14609 , n14604 , n14607 , n14608 );
xor ( n14610 , n14513 , n14517 );
xor ( n14611 , n14610 , n14522 );
and ( n14612 , n14609 , n14611 );
xor ( n14613 , n14412 , n14416 );
xor ( n14614 , n14613 , n14419 );
and ( n14615 , n14611 , n14614 );
and ( n14616 , n14609 , n14614 );
or ( n14617 , n14612 , n14615 , n14616 );
and ( n14618 , n9701 , n7395 );
and ( n14619 , n9463 , n7393 );
nor ( n14620 , n14618 , n14619 );
xnor ( n14621 , n14620 , n7405 );
and ( n14622 , n14617 , n14621 );
and ( n14623 , n10377 , n8044 );
and ( n14624 , n10239 , n8042 );
nor ( n14625 , n14623 , n14624 );
xnor ( n14626 , n14625 , n8054 );
and ( n14627 , n14621 , n14626 );
and ( n14628 , n14617 , n14626 );
or ( n14629 , n14622 , n14627 , n14628 );
and ( n14630 , n9196 , n8168 );
and ( n14631 , n9049 , n8166 );
nor ( n14632 , n14630 , n14631 );
xnor ( n14633 , n14632 , n8178 );
and ( n14634 , n14629 , n14633 );
xor ( n14635 , n14549 , n14553 );
xor ( n14636 , n14635 , n14556 );
and ( n14637 , n14633 , n14636 );
and ( n14638 , n14629 , n14636 );
or ( n14639 , n14634 , n14637 , n14638 );
xor ( n14640 , n14392 , n14396 );
xor ( n14641 , n14640 , n14401 );
and ( n14642 , n14639 , n14641 );
xor ( n14643 , n14444 , n14446 );
xor ( n14644 , n14643 , n14459 );
and ( n14645 , n14641 , n14644 );
and ( n14646 , n14639 , n14644 );
or ( n14647 , n14642 , n14645 , n14646 );
xor ( n14648 , n14404 , n14462 );
xor ( n14649 , n14648 , n14467 );
and ( n14650 , n14647 , n14649 );
xor ( n14651 , n14567 , n14569 );
xor ( n14652 , n14651 , n14572 );
and ( n14653 , n14649 , n14652 );
and ( n14654 , n14647 , n14652 );
or ( n14655 , n14650 , n14653 , n14654 );
and ( n14656 , n14587 , n14655 );
xor ( n14657 , n14587 , n14655 );
and ( n14658 , n11817 , n7954 );
and ( n14659 , n11710 , n7952 );
nor ( n14660 , n14658 , n14659 );
xnor ( n14661 , n14660 , n7964 );
and ( n14662 , n12246 , n7499 );
not ( n14663 , n14662 );
and ( n14664 , n14663 , n7511 );
and ( n14665 , n14661 , n14664 );
and ( n14666 , n11569 , n7933 );
and ( n14667 , n11435 , n7931 );
nor ( n14668 , n14666 , n14667 );
xnor ( n14669 , n14668 , n7939 );
and ( n14670 , n14665 , n14669 );
xor ( n14671 , n14591 , n14595 );
xor ( n14672 , n14671 , n14409 );
and ( n14673 , n14669 , n14672 );
and ( n14674 , n14665 , n14672 );
or ( n14675 , n14670 , n14673 , n14674 );
and ( n14676 , n11249 , n7781 );
and ( n14677 , n11187 , n7779 );
nor ( n14678 , n14676 , n14677 );
xnor ( n14679 , n14678 , n7791 );
and ( n14680 , n14675 , n14679 );
xor ( n14681 , n14599 , n14603 );
xor ( n14682 , n14681 , n14606 );
and ( n14683 , n14679 , n14682 );
and ( n14684 , n14675 , n14682 );
or ( n14685 , n14680 , n14683 , n14684 );
and ( n14686 , n10239 , n7899 );
and ( n14687 , n10032 , n7897 );
nor ( n14688 , n14686 , n14687 );
xnor ( n14689 , n14688 , n7909 );
and ( n14690 , n14685 , n14689 );
and ( n14691 , n10559 , n8044 );
and ( n14692 , n10377 , n8042 );
nor ( n14693 , n14691 , n14692 );
xnor ( n14694 , n14693 , n8054 );
and ( n14695 , n14689 , n14694 );
and ( n14696 , n14685 , n14694 );
or ( n14697 , n14690 , n14695 , n14696 );
and ( n14698 , n9463 , n8168 );
and ( n14699 , n9280 , n8166 );
nor ( n14700 , n14698 , n14699 );
xnor ( n14701 , n14700 , n8178 );
and ( n14702 , n9829 , n7395 );
and ( n14703 , n9701 , n7393 );
nor ( n14704 , n14702 , n14703 );
xnor ( n14705 , n14704 , n7405 );
and ( n14706 , n14701 , n14705 );
xor ( n14707 , n14609 , n14611 );
xor ( n14708 , n14707 , n14614 );
and ( n14709 , n14705 , n14708 );
and ( n14710 , n14701 , n14708 );
or ( n14711 , n14706 , n14709 , n14710 );
and ( n14712 , n14697 , n14711 );
and ( n14713 , n9049 , n7318 );
and ( n14714 , n8696 , n7315 );
nor ( n14715 , n14713 , n14714 );
xnor ( n14716 , n14715 , n7311 );
and ( n14717 , n14711 , n14716 );
and ( n14718 , n14697 , n14716 );
or ( n14719 , n14712 , n14717 , n14718 );
and ( n14720 , n9280 , n8168 );
and ( n14721 , n9196 , n8166 );
nor ( n14722 , n14720 , n14721 );
xnor ( n14723 , n14722 , n8178 );
and ( n14724 , n10032 , n7899 );
and ( n14725 , n9829 , n7897 );
nor ( n14726 , n14724 , n14725 );
xnor ( n14727 , n14726 , n7909 );
and ( n14728 , n14723 , n14727 );
xor ( n14729 , n14525 , n14529 );
xor ( n14730 , n14729 , n14532 );
and ( n14731 , n14727 , n14730 );
and ( n14732 , n14723 , n14730 );
or ( n14733 , n14728 , n14731 , n14732 );
and ( n14734 , n14719 , n14733 );
xor ( n14735 , n14535 , n14539 );
xor ( n14736 , n14735 , n14542 );
and ( n14737 , n14733 , n14736 );
and ( n14738 , n14719 , n14736 );
or ( n14739 , n14734 , n14737 , n14738 );
xor ( n14740 , n14545 , n14559 );
xor ( n14741 , n14740 , n14564 );
and ( n14742 , n14739 , n14741 );
xor ( n14743 , n14639 , n14641 );
xor ( n14744 , n14743 , n14644 );
and ( n14745 , n14741 , n14744 );
and ( n14746 , n14739 , n14744 );
or ( n14747 , n14742 , n14745 , n14746 );
xor ( n14748 , n14647 , n14649 );
xor ( n14749 , n14748 , n14652 );
and ( n14750 , n14747 , n14749 );
xor ( n14751 , n14747 , n14749 );
xor ( n14752 , n14739 , n14741 );
xor ( n14753 , n14752 , n14744 );
xor ( n14754 , n14661 , n14664 );
and ( n14755 , n11697 , n7933 );
and ( n14756 , n11569 , n7931 );
nor ( n14757 , n14755 , n14756 );
xnor ( n14758 , n14757 , n7939 );
and ( n14759 , n14754 , n14758 );
and ( n14760 , n12246 , n7501 );
and ( n14761 , n12012 , n7499 );
nor ( n14762 , n14760 , n14761 );
xnor ( n14763 , n14762 , n7511 );
and ( n14764 , n14758 , n14763 );
and ( n14765 , n14754 , n14763 );
or ( n14766 , n14759 , n14764 , n14765 );
and ( n14767 , n11383 , n7781 );
and ( n14768 , n11249 , n7779 );
nor ( n14769 , n14767 , n14768 );
xnor ( n14770 , n14769 , n7791 );
and ( n14771 , n14766 , n14770 );
xor ( n14772 , n14665 , n14669 );
xor ( n14773 , n14772 , n14672 );
and ( n14774 , n14770 , n14773 );
and ( n14775 , n14766 , n14773 );
or ( n14776 , n14771 , n14774 , n14775 );
and ( n14777 , n10554 , n8044 );
and ( n14778 , n10559 , n8042 );
nor ( n14779 , n14777 , n14778 );
xnor ( n14780 , n14779 , n8054 );
and ( n14781 , n14776 , n14780 );
xor ( n14782 , n14675 , n14679 );
xor ( n14783 , n14782 , n14682 );
and ( n14784 , n14780 , n14783 );
and ( n14785 , n14776 , n14783 );
or ( n14786 , n14781 , n14784 , n14785 );
and ( n14787 , n9196 , n7318 );
and ( n14788 , n9049 , n7315 );
nor ( n14789 , n14787 , n14788 );
xnor ( n14790 , n14789 , n7311 );
and ( n14791 , n14786 , n14790 );
xor ( n14792 , n14685 , n14689 );
xor ( n14793 , n14792 , n14694 );
and ( n14794 , n14790 , n14793 );
and ( n14795 , n14786 , n14793 );
or ( n14796 , n14791 , n14794 , n14795 );
xor ( n14797 , n14617 , n14621 );
xor ( n14798 , n14797 , n14626 );
and ( n14799 , n14796 , n14798 );
xor ( n14800 , n14723 , n14727 );
xor ( n14801 , n14800 , n14730 );
and ( n14802 , n14798 , n14801 );
and ( n14803 , n14796 , n14801 );
or ( n14804 , n14799 , n14802 , n14803 );
xor ( n14805 , n14719 , n14733 );
xor ( n14806 , n14805 , n14736 );
and ( n14807 , n14804 , n14806 );
xor ( n14808 , n14629 , n14633 );
xor ( n14809 , n14808 , n14636 );
and ( n14810 , n14806 , n14809 );
and ( n14811 , n14804 , n14809 );
or ( n14812 , n14807 , n14810 , n14811 );
and ( n14813 , n14753 , n14812 );
xor ( n14814 , n14753 , n14812 );
xor ( n14815 , n14804 , n14806 );
xor ( n14816 , n14815 , n14809 );
and ( n14817 , n11710 , n7933 );
and ( n14818 , n11697 , n7931 );
nor ( n14819 , n14817 , n14818 );
xnor ( n14820 , n14819 , n7939 );
and ( n14821 , n12012 , n7954 );
and ( n14822 , n11817 , n7952 );
nor ( n14823 , n14821 , n14822 );
xnor ( n14824 , n14823 , n7964 );
and ( n14825 , n14820 , n14824 );
and ( n14826 , n14824 , n14662 );
and ( n14827 , n14820 , n14662 );
or ( n14828 , n14825 , n14826 , n14827 );
and ( n14829 , n11435 , n7781 );
and ( n14830 , n11383 , n7779 );
nor ( n14831 , n14829 , n14830 );
xnor ( n14832 , n14831 , n7791 );
and ( n14833 , n14828 , n14832 );
xor ( n14834 , n14754 , n14758 );
xor ( n14835 , n14834 , n14763 );
and ( n14836 , n14832 , n14835 );
and ( n14837 , n14828 , n14835 );
or ( n14838 , n14833 , n14836 , n14837 );
and ( n14839 , n11187 , n8044 );
and ( n14840 , n10554 , n8042 );
nor ( n14841 , n14839 , n14840 );
xnor ( n14842 , n14841 , n8054 );
and ( n14843 , n14838 , n14842 );
xor ( n14844 , n14766 , n14770 );
xor ( n14845 , n14844 , n14773 );
and ( n14846 , n14842 , n14845 );
and ( n14847 , n14838 , n14845 );
or ( n14848 , n14843 , n14846 , n14847 );
and ( n14849 , n9701 , n8168 );
and ( n14850 , n9463 , n8166 );
nor ( n14851 , n14849 , n14850 );
xnor ( n14852 , n14851 , n8178 );
and ( n14853 , n14848 , n14852 );
and ( n14854 , n10377 , n7899 );
and ( n14855 , n10239 , n7897 );
nor ( n14856 , n14854 , n14855 );
xnor ( n14857 , n14856 , n7909 );
and ( n14858 , n14852 , n14857 );
and ( n14859 , n14848 , n14857 );
or ( n14860 , n14853 , n14858 , n14859 );
and ( n14861 , n11817 , n7933 );
and ( n14862 , n11710 , n7931 );
nor ( n14863 , n14861 , n14862 );
xnor ( n14864 , n14863 , n7939 );
and ( n14865 , n12246 , n7952 );
not ( n14866 , n14865 );
and ( n14867 , n14866 , n7964 );
and ( n14868 , n14864 , n14867 );
and ( n14869 , n11569 , n7781 );
and ( n14870 , n11435 , n7779 );
nor ( n14871 , n14869 , n14870 );
xnor ( n14872 , n14871 , n7791 );
and ( n14873 , n14868 , n14872 );
xor ( n14874 , n14820 , n14824 );
xor ( n14875 , n14874 , n14662 );
and ( n14876 , n14872 , n14875 );
and ( n14877 , n14868 , n14875 );
or ( n14878 , n14873 , n14876 , n14877 );
and ( n14879 , n11249 , n8044 );
and ( n14880 , n11187 , n8042 );
nor ( n14881 , n14879 , n14880 );
xnor ( n14882 , n14881 , n8054 );
and ( n14883 , n14878 , n14882 );
xor ( n14884 , n14828 , n14832 );
xor ( n14885 , n14884 , n14835 );
and ( n14886 , n14882 , n14885 );
and ( n14887 , n14878 , n14885 );
or ( n14888 , n14883 , n14886 , n14887 );
and ( n14889 , n10239 , n7395 );
and ( n14890 , n10032 , n7393 );
nor ( n14891 , n14889 , n14890 );
xnor ( n14892 , n14891 , n7405 );
and ( n14893 , n14888 , n14892 );
and ( n14894 , n10559 , n7899 );
and ( n14895 , n10377 , n7897 );
nor ( n14896 , n14894 , n14895 );
xnor ( n14897 , n14896 , n7909 );
and ( n14898 , n14892 , n14897 );
and ( n14899 , n14888 , n14897 );
or ( n14900 , n14893 , n14898 , n14899 );
and ( n14901 , n10032 , n7395 );
and ( n14902 , n9829 , n7393 );
nor ( n14903 , n14901 , n14902 );
xnor ( n14904 , n14903 , n7405 );
and ( n14905 , n14900 , n14904 );
xor ( n14906 , n14776 , n14780 );
xor ( n14907 , n14906 , n14783 );
and ( n14908 , n14904 , n14907 );
and ( n14909 , n14900 , n14907 );
or ( n14910 , n14905 , n14908 , n14909 );
and ( n14911 , n14860 , n14910 );
xor ( n14912 , n14701 , n14705 );
xor ( n14913 , n14912 , n14708 );
and ( n14914 , n14910 , n14913 );
and ( n14915 , n14860 , n14913 );
or ( n14916 , n14911 , n14914 , n14915 );
xor ( n14917 , n14697 , n14711 );
xor ( n14918 , n14917 , n14716 );
and ( n14919 , n14916 , n14918 );
xor ( n14920 , n14796 , n14798 );
xor ( n14921 , n14920 , n14801 );
and ( n14922 , n14918 , n14921 );
and ( n14923 , n14916 , n14921 );
or ( n14924 , n14919 , n14922 , n14923 );
and ( n14925 , n14816 , n14924 );
xor ( n14926 , n14816 , n14924 );
xor ( n14927 , n14916 , n14918 );
xor ( n14928 , n14927 , n14921 );
xor ( n14929 , n14864 , n14867 );
and ( n14930 , n11697 , n7781 );
and ( n14931 , n11569 , n7779 );
nor ( n14932 , n14930 , n14931 );
xnor ( n14933 , n14932 , n7791 );
and ( n14934 , n14929 , n14933 );
and ( n14935 , n12246 , n7954 );
and ( n14936 , n12012 , n7952 );
nor ( n14937 , n14935 , n14936 );
xnor ( n14938 , n14937 , n7964 );
and ( n14939 , n14933 , n14938 );
and ( n14940 , n14929 , n14938 );
or ( n14941 , n14934 , n14939 , n14940 );
and ( n14942 , n11187 , n7899 );
and ( n14943 , n10554 , n7897 );
nor ( n14944 , n14942 , n14943 );
xnor ( n14945 , n14944 , n7909 );
and ( n14946 , n14941 , n14945 );
and ( n14947 , n11383 , n8044 );
and ( n14948 , n11249 , n8042 );
nor ( n14949 , n14947 , n14948 );
xnor ( n14950 , n14949 , n8054 );
and ( n14951 , n14945 , n14950 );
and ( n14952 , n14941 , n14950 );
or ( n14953 , n14946 , n14951 , n14952 );
and ( n14954 , n10554 , n7899 );
and ( n14955 , n10559 , n7897 );
nor ( n14956 , n14954 , n14955 );
xnor ( n14957 , n14956 , n7909 );
and ( n14958 , n14953 , n14957 );
xor ( n14959 , n14878 , n14882 );
xor ( n14960 , n14959 , n14885 );
and ( n14961 , n14957 , n14960 );
and ( n14962 , n14953 , n14960 );
or ( n14963 , n14958 , n14961 , n14962 );
and ( n14964 , n9829 , n8168 );
and ( n14965 , n9701 , n8166 );
nor ( n14966 , n14964 , n14965 );
xnor ( n14967 , n14966 , n8178 );
and ( n14968 , n14963 , n14967 );
xor ( n14969 , n14838 , n14842 );
xor ( n14970 , n14969 , n14845 );
and ( n14971 , n14967 , n14970 );
and ( n14972 , n14963 , n14970 );
or ( n14973 , n14968 , n14971 , n14972 );
and ( n14974 , n9280 , n7318 );
and ( n14975 , n9196 , n7315 );
nor ( n14976 , n14974 , n14975 );
xnor ( n14977 , n14976 , n7311 );
and ( n14978 , n14973 , n14977 );
xor ( n14979 , n14848 , n14852 );
xor ( n14980 , n14979 , n14857 );
and ( n14981 , n14977 , n14980 );
and ( n14982 , n14973 , n14980 );
or ( n14983 , n14978 , n14981 , n14982 );
xor ( n14984 , n14786 , n14790 );
xor ( n14985 , n14984 , n14793 );
and ( n14986 , n14983 , n14985 );
xor ( n14987 , n14860 , n14910 );
xor ( n14988 , n14987 , n14913 );
and ( n14989 , n14985 , n14988 );
and ( n14990 , n14983 , n14988 );
or ( n14991 , n14986 , n14989 , n14990 );
and ( n14992 , n14928 , n14991 );
xor ( n14993 , n14928 , n14991 );
xor ( n14994 , n14983 , n14985 );
xor ( n14995 , n14994 , n14988 );
and ( n14996 , n11710 , n7781 );
and ( n14997 , n11697 , n7779 );
nor ( n14998 , n14996 , n14997 );
xnor ( n14999 , n14998 , n7791 );
and ( n15000 , n12012 , n7933 );
and ( n15001 , n11817 , n7931 );
nor ( n15002 , n15000 , n15001 );
xnor ( n15003 , n15002 , n7939 );
and ( n15004 , n14999 , n15003 );
and ( n15005 , n15003 , n14865 );
and ( n15006 , n14999 , n14865 );
or ( n15007 , n15004 , n15005 , n15006 );
and ( n15008 , n11435 , n8044 );
and ( n15009 , n11383 , n8042 );
nor ( n15010 , n15008 , n15009 );
xnor ( n15011 , n15010 , n8054 );
and ( n15012 , n15007 , n15011 );
xor ( n15013 , n14929 , n14933 );
xor ( n15014 , n15013 , n14938 );
and ( n15015 , n15011 , n15014 );
and ( n15016 , n15007 , n15014 );
or ( n15017 , n15012 , n15015 , n15016 );
xor ( n15018 , n14941 , n14945 );
xor ( n15019 , n15018 , n14950 );
and ( n15020 , n15017 , n15019 );
xor ( n15021 , n14868 , n14872 );
xor ( n15022 , n15021 , n14875 );
and ( n15023 , n15019 , n15022 );
and ( n15024 , n15017 , n15022 );
or ( n15025 , n15020 , n15023 , n15024 );
and ( n15026 , n10032 , n8168 );
and ( n15027 , n9829 , n8166 );
nor ( n15028 , n15026 , n15027 );
xnor ( n15029 , n15028 , n8178 );
and ( n15030 , n15025 , n15029 );
and ( n15031 , n10377 , n7395 );
and ( n15032 , n10239 , n7393 );
nor ( n15033 , n15031 , n15032 );
xnor ( n15034 , n15033 , n7405 );
and ( n15035 , n15029 , n15034 );
and ( n15036 , n15025 , n15034 );
or ( n15037 , n15030 , n15035 , n15036 );
and ( n15038 , n9463 , n7318 );
and ( n15039 , n9280 , n7315 );
nor ( n15040 , n15038 , n15039 );
xnor ( n15041 , n15040 , n7311 );
and ( n15042 , n15037 , n15041 );
xor ( n15043 , n14888 , n14892 );
xor ( n15044 , n15043 , n14897 );
and ( n15045 , n15041 , n15044 );
and ( n15046 , n15037 , n15044 );
or ( n15047 , n15042 , n15045 , n15046 );
xor ( n15048 , n14973 , n14977 );
xor ( n15049 , n15048 , n14980 );
and ( n15050 , n15047 , n15049 );
xor ( n15051 , n14900 , n14904 );
xor ( n15052 , n15051 , n14907 );
and ( n15053 , n15049 , n15052 );
and ( n15054 , n15047 , n15052 );
or ( n15055 , n15050 , n15053 , n15054 );
and ( n15056 , n14995 , n15055 );
xor ( n15057 , n14995 , n15055 );
and ( n15058 , n11817 , n7781 );
and ( n15059 , n11710 , n7779 );
nor ( n15060 , n15058 , n15059 );
xnor ( n15061 , n15060 , n7791 );
and ( n15062 , n12246 , n7931 );
not ( n15063 , n15062 );
and ( n15064 , n15063 , n7939 );
and ( n15065 , n15061 , n15064 );
and ( n15066 , n11569 , n8044 );
and ( n15067 , n11435 , n8042 );
nor ( n15068 , n15066 , n15067 );
xnor ( n15069 , n15068 , n8054 );
and ( n15070 , n15065 , n15069 );
xor ( n15071 , n14999 , n15003 );
xor ( n15072 , n15071 , n14865 );
and ( n15073 , n15069 , n15072 );
and ( n15074 , n15065 , n15072 );
or ( n15075 , n15070 , n15073 , n15074 );
and ( n15076 , n11249 , n7899 );
and ( n15077 , n11187 , n7897 );
nor ( n15078 , n15076 , n15077 );
xnor ( n15079 , n15078 , n7909 );
and ( n15080 , n15075 , n15079 );
xor ( n15081 , n15007 , n15011 );
xor ( n15082 , n15081 , n15014 );
and ( n15083 , n15079 , n15082 );
and ( n15084 , n15075 , n15082 );
or ( n15085 , n15080 , n15083 , n15084 );
and ( n15086 , n10239 , n8168 );
and ( n15087 , n10032 , n8166 );
nor ( n15088 , n15086 , n15087 );
xnor ( n15089 , n15088 , n8178 );
and ( n15090 , n15085 , n15089 );
and ( n15091 , n10559 , n7395 );
and ( n15092 , n10377 , n7393 );
nor ( n15093 , n15091 , n15092 );
xnor ( n15094 , n15093 , n7405 );
and ( n15095 , n15089 , n15094 );
and ( n15096 , n15085 , n15094 );
or ( n15097 , n15090 , n15095 , n15096 );
and ( n15098 , n9701 , n7318 );
and ( n15099 , n9463 , n7315 );
nor ( n15100 , n15098 , n15099 );
xnor ( n15101 , n15100 , n7311 );
and ( n15102 , n15097 , n15101 );
xor ( n15103 , n14953 , n14957 );
xor ( n15104 , n15103 , n14960 );
and ( n15105 , n15101 , n15104 );
and ( n15106 , n15097 , n15104 );
or ( n15107 , n15102 , n15105 , n15106 );
xor ( n15108 , n15037 , n15041 );
xor ( n15109 , n15108 , n15044 );
and ( n15110 , n15107 , n15109 );
xor ( n15111 , n14963 , n14967 );
xor ( n15112 , n15111 , n14970 );
and ( n15113 , n15109 , n15112 );
and ( n15114 , n15107 , n15112 );
or ( n15115 , n15110 , n15113 , n15114 );
xor ( n15116 , n15047 , n15049 );
xor ( n15117 , n15116 , n15052 );
and ( n15118 , n15115 , n15117 );
xor ( n15119 , n15115 , n15117 );
xor ( n15120 , n15107 , n15109 );
xor ( n15121 , n15120 , n15112 );
xor ( n15122 , n15061 , n15064 );
and ( n15123 , n11697 , n8044 );
and ( n15124 , n11569 , n8042 );
nor ( n15125 , n15123 , n15124 );
xnor ( n15126 , n15125 , n8054 );
and ( n15127 , n15122 , n15126 );
and ( n15128 , n12246 , n7933 );
and ( n15129 , n12012 , n7931 );
nor ( n15130 , n15128 , n15129 );
xnor ( n15131 , n15130 , n7939 );
and ( n15132 , n15126 , n15131 );
and ( n15133 , n15122 , n15131 );
or ( n15134 , n15127 , n15132 , n15133 );
and ( n15135 , n11383 , n7899 );
and ( n15136 , n11249 , n7897 );
nor ( n15137 , n15135 , n15136 );
xnor ( n15138 , n15137 , n7909 );
and ( n15139 , n15134 , n15138 );
xor ( n15140 , n15065 , n15069 );
xor ( n15141 , n15140 , n15072 );
and ( n15142 , n15138 , n15141 );
and ( n15143 , n15134 , n15141 );
or ( n15144 , n15139 , n15142 , n15143 );
and ( n15145 , n10554 , n7395 );
and ( n15146 , n10559 , n7393 );
nor ( n15147 , n15145 , n15146 );
xnor ( n15148 , n15147 , n7405 );
and ( n15149 , n15144 , n15148 );
xor ( n15150 , n15075 , n15079 );
xor ( n15151 , n15150 , n15082 );
and ( n15152 , n15148 , n15151 );
and ( n15153 , n15144 , n15151 );
or ( n15154 , n15149 , n15152 , n15153 );
and ( n15155 , n9829 , n7318 );
and ( n15156 , n9701 , n7315 );
nor ( n15157 , n15155 , n15156 );
xnor ( n15158 , n15157 , n7311 );
and ( n15159 , n15154 , n15158 );
xor ( n15160 , n15017 , n15019 );
xor ( n15161 , n15160 , n15022 );
and ( n15162 , n15158 , n15161 );
and ( n15163 , n15154 , n15161 );
or ( n15164 , n15159 , n15162 , n15163 );
xor ( n15165 , n15025 , n15029 );
xor ( n15166 , n15165 , n15034 );
and ( n15167 , n15164 , n15166 );
xor ( n15168 , n15097 , n15101 );
xor ( n15169 , n15168 , n15104 );
and ( n15170 , n15166 , n15169 );
and ( n15171 , n15164 , n15169 );
or ( n15172 , n15167 , n15170 , n15171 );
and ( n15173 , n15121 , n15172 );
xor ( n15174 , n15121 , n15172 );
xor ( n15175 , n15164 , n15166 );
xor ( n15176 , n15175 , n15169 );
and ( n15177 , n11710 , n8044 );
and ( n15178 , n11697 , n8042 );
nor ( n15179 , n15177 , n15178 );
xnor ( n15180 , n15179 , n8054 );
and ( n15181 , n12012 , n7781 );
and ( n15182 , n11817 , n7779 );
nor ( n15183 , n15181 , n15182 );
xnor ( n15184 , n15183 , n7791 );
and ( n15185 , n15180 , n15184 );
and ( n15186 , n15184 , n15062 );
and ( n15187 , n15180 , n15062 );
or ( n15188 , n15185 , n15186 , n15187 );
and ( n15189 , n11435 , n7899 );
and ( n15190 , n11383 , n7897 );
nor ( n15191 , n15189 , n15190 );
xnor ( n15192 , n15191 , n7909 );
and ( n15193 , n15188 , n15192 );
xor ( n15194 , n15122 , n15126 );
xor ( n15195 , n15194 , n15131 );
and ( n15196 , n15192 , n15195 );
and ( n15197 , n15188 , n15195 );
or ( n15198 , n15193 , n15196 , n15197 );
and ( n15199 , n11187 , n7395 );
and ( n15200 , n10554 , n7393 );
nor ( n15201 , n15199 , n15200 );
xnor ( n15202 , n15201 , n7405 );
and ( n15203 , n15198 , n15202 );
xor ( n15204 , n15134 , n15138 );
xor ( n15205 , n15204 , n15141 );
and ( n15206 , n15202 , n15205 );
and ( n15207 , n15198 , n15205 );
or ( n15208 , n15203 , n15206 , n15207 );
and ( n15209 , n10032 , n7318 );
and ( n15210 , n9829 , n7315 );
nor ( n15211 , n15209 , n15210 );
xnor ( n15212 , n15211 , n7311 );
and ( n15213 , n15208 , n15212 );
and ( n15214 , n10377 , n8168 );
and ( n15215 , n10239 , n8166 );
nor ( n15216 , n15214 , n15215 );
xnor ( n15217 , n15216 , n8178 );
and ( n15218 , n15212 , n15217 );
and ( n15219 , n15208 , n15217 );
or ( n15220 , n15213 , n15218 , n15219 );
xor ( n15221 , n15085 , n15089 );
xor ( n15222 , n15221 , n15094 );
and ( n15223 , n15220 , n15222 );
xor ( n15224 , n15154 , n15158 );
xor ( n15225 , n15224 , n15161 );
and ( n15226 , n15222 , n15225 );
and ( n15227 , n15220 , n15225 );
or ( n15228 , n15223 , n15226 , n15227 );
and ( n15229 , n15176 , n15228 );
xor ( n15230 , n15176 , n15228 );
and ( n15231 , n11817 , n8044 );
and ( n15232 , n11710 , n8042 );
nor ( n15233 , n15231 , n15232 );
xnor ( n15234 , n15233 , n8054 );
and ( n15235 , n12246 , n7779 );
not ( n15236 , n15235 );
and ( n15237 , n15236 , n7791 );
and ( n15238 , n15234 , n15237 );
and ( n15239 , n11569 , n7899 );
and ( n15240 , n11435 , n7897 );
nor ( n15241 , n15239 , n15240 );
xnor ( n15242 , n15241 , n7909 );
and ( n15243 , n15238 , n15242 );
xor ( n15244 , n15180 , n15184 );
xor ( n15245 , n15244 , n15062 );
and ( n15246 , n15242 , n15245 );
and ( n15247 , n15238 , n15245 );
or ( n15248 , n15243 , n15246 , n15247 );
and ( n15249 , n11249 , n7395 );
and ( n15250 , n11187 , n7393 );
nor ( n15251 , n15249 , n15250 );
xnor ( n15252 , n15251 , n7405 );
and ( n15253 , n15248 , n15252 );
xor ( n15254 , n15188 , n15192 );
xor ( n15255 , n15254 , n15195 );
and ( n15256 , n15252 , n15255 );
and ( n15257 , n15248 , n15255 );
or ( n15258 , n15253 , n15256 , n15257 );
and ( n15259 , n10239 , n7318 );
and ( n15260 , n10032 , n7315 );
nor ( n15261 , n15259 , n15260 );
xnor ( n15262 , n15261 , n7311 );
and ( n15263 , n15258 , n15262 );
and ( n15264 , n10559 , n8168 );
and ( n15265 , n10377 , n8166 );
nor ( n15266 , n15264 , n15265 );
xnor ( n15267 , n15266 , n8178 );
and ( n15268 , n15262 , n15267 );
and ( n15269 , n15258 , n15267 );
or ( n15270 , n15263 , n15268 , n15269 );
xor ( n15271 , n15208 , n15212 );
xor ( n15272 , n15271 , n15217 );
and ( n15273 , n15270 , n15272 );
xor ( n15274 , n15144 , n15148 );
xor ( n15275 , n15274 , n15151 );
and ( n15276 , n15272 , n15275 );
and ( n15277 , n15270 , n15275 );
or ( n15278 , n15273 , n15276 , n15277 );
xor ( n15279 , n15220 , n15222 );
xor ( n15280 , n15279 , n15225 );
and ( n15281 , n15278 , n15280 );
xor ( n15282 , n15278 , n15280 );
xor ( n15283 , n15270 , n15272 );
xor ( n15284 , n15283 , n15275 );
xor ( n15285 , n15234 , n15237 );
and ( n15286 , n11697 , n7899 );
and ( n15287 , n11569 , n7897 );
nor ( n15288 , n15286 , n15287 );
xnor ( n15289 , n15288 , n7909 );
and ( n15290 , n15285 , n15289 );
and ( n15291 , n12246 , n7781 );
and ( n15292 , n12012 , n7779 );
nor ( n15293 , n15291 , n15292 );
xnor ( n15294 , n15293 , n7791 );
and ( n15295 , n15289 , n15294 );
and ( n15296 , n15285 , n15294 );
or ( n15297 , n15290 , n15295 , n15296 );
and ( n15298 , n11383 , n7395 );
and ( n15299 , n11249 , n7393 );
nor ( n15300 , n15298 , n15299 );
xnor ( n15301 , n15300 , n7405 );
and ( n15302 , n15297 , n15301 );
xor ( n15303 , n15238 , n15242 );
xor ( n15304 , n15303 , n15245 );
and ( n15305 , n15301 , n15304 );
and ( n15306 , n15297 , n15304 );
or ( n15307 , n15302 , n15305 , n15306 );
and ( n15308 , n10554 , n8168 );
and ( n15309 , n10559 , n8166 );
nor ( n15310 , n15308 , n15309 );
xnor ( n15311 , n15310 , n8178 );
and ( n15312 , n15307 , n15311 );
xor ( n15313 , n15248 , n15252 );
xor ( n15314 , n15313 , n15255 );
and ( n15315 , n15311 , n15314 );
and ( n15316 , n15307 , n15314 );
or ( n15317 , n15312 , n15315 , n15316 );
xor ( n15318 , n15258 , n15262 );
xor ( n15319 , n15318 , n15267 );
and ( n15320 , n15317 , n15319 );
xor ( n15321 , n15198 , n15202 );
xor ( n15322 , n15321 , n15205 );
and ( n15323 , n15319 , n15322 );
and ( n15324 , n15317 , n15322 );
or ( n15325 , n15320 , n15323 , n15324 );
and ( n15326 , n15284 , n15325 );
xor ( n15327 , n15284 , n15325 );
xor ( n15328 , n15317 , n15319 );
xor ( n15329 , n15328 , n15322 );
and ( n15330 , n11710 , n7899 );
and ( n15331 , n11697 , n7897 );
nor ( n15332 , n15330 , n15331 );
xnor ( n15333 , n15332 , n7909 );
and ( n15334 , n12012 , n8044 );
and ( n15335 , n11817 , n8042 );
nor ( n15336 , n15334 , n15335 );
xnor ( n15337 , n15336 , n8054 );
and ( n15338 , n15333 , n15337 );
and ( n15339 , n15337 , n15235 );
and ( n15340 , n15333 , n15235 );
or ( n15341 , n15338 , n15339 , n15340 );
and ( n15342 , n11435 , n7395 );
and ( n15343 , n11383 , n7393 );
nor ( n15344 , n15342 , n15343 );
xnor ( n15345 , n15344 , n7405 );
and ( n15346 , n15341 , n15345 );
xor ( n15347 , n15285 , n15289 );
xor ( n15348 , n15347 , n15294 );
and ( n15349 , n15345 , n15348 );
and ( n15350 , n15341 , n15348 );
or ( n15351 , n15346 , n15349 , n15350 );
and ( n15352 , n11187 , n8168 );
and ( n15353 , n10554 , n8166 );
nor ( n15354 , n15352 , n15353 );
xnor ( n15355 , n15354 , n8178 );
and ( n15356 , n15351 , n15355 );
xor ( n15357 , n15297 , n15301 );
xor ( n15358 , n15357 , n15304 );
and ( n15359 , n15355 , n15358 );
and ( n15360 , n15351 , n15358 );
or ( n15361 , n15356 , n15359 , n15360 );
and ( n15362 , n10377 , n7318 );
and ( n15363 , n10239 , n7315 );
nor ( n15364 , n15362 , n15363 );
xnor ( n15365 , n15364 , n7311 );
and ( n15366 , n15361 , n15365 );
xor ( n15367 , n15307 , n15311 );
xor ( n15368 , n15367 , n15314 );
and ( n15369 , n15365 , n15368 );
and ( n15370 , n15361 , n15368 );
or ( n15371 , n15366 , n15369 , n15370 );
and ( n15372 , n15329 , n15371 );
xor ( n15373 , n15329 , n15371 );
and ( n15374 , n11817 , n7899 );
and ( n15375 , n11710 , n7897 );
nor ( n15376 , n15374 , n15375 );
xnor ( n15377 , n15376 , n7909 );
and ( n15378 , n12246 , n8042 );
not ( n15379 , n15378 );
and ( n15380 , n15379 , n8054 );
and ( n15381 , n15377 , n15380 );
and ( n15382 , n11569 , n7395 );
and ( n15383 , n11435 , n7393 );
nor ( n15384 , n15382 , n15383 );
xnor ( n15385 , n15384 , n7405 );
and ( n15386 , n15381 , n15385 );
xor ( n15387 , n15333 , n15337 );
xor ( n15388 , n15387 , n15235 );
and ( n15389 , n15385 , n15388 );
and ( n15390 , n15381 , n15388 );
or ( n15391 , n15386 , n15389 , n15390 );
and ( n15392 , n11249 , n8168 );
and ( n15393 , n11187 , n8166 );
nor ( n15394 , n15392 , n15393 );
xnor ( n15395 , n15394 , n8178 );
and ( n15396 , n15391 , n15395 );
xor ( n15397 , n15341 , n15345 );
xor ( n15398 , n15397 , n15348 );
and ( n15399 , n15395 , n15398 );
and ( n15400 , n15391 , n15398 );
or ( n15401 , n15396 , n15399 , n15400 );
and ( n15402 , n10559 , n7318 );
and ( n15403 , n10377 , n7315 );
nor ( n15404 , n15402 , n15403 );
xnor ( n15405 , n15404 , n7311 );
and ( n15406 , n15401 , n15405 );
xor ( n15407 , n15351 , n15355 );
xor ( n15408 , n15407 , n15358 );
and ( n15409 , n15405 , n15408 );
and ( n15410 , n15401 , n15408 );
or ( n15411 , n15406 , n15409 , n15410 );
xor ( n15412 , n15361 , n15365 );
xor ( n15413 , n15412 , n15368 );
and ( n15414 , n15411 , n15413 );
xor ( n15415 , n15411 , n15413 );
xor ( n15416 , n15401 , n15405 );
xor ( n15417 , n15416 , n15408 );
xor ( n15418 , n15377 , n15380 );
and ( n15419 , n11697 , n7395 );
and ( n15420 , n11569 , n7393 );
nor ( n15421 , n15419 , n15420 );
xnor ( n15422 , n15421 , n7405 );
and ( n15423 , n15418 , n15422 );
and ( n15424 , n12246 , n8044 );
and ( n15425 , n12012 , n8042 );
nor ( n15426 , n15424 , n15425 );
xnor ( n15427 , n15426 , n8054 );
and ( n15428 , n15422 , n15427 );
and ( n15429 , n15418 , n15427 );
or ( n15430 , n15423 , n15428 , n15429 );
and ( n15431 , n11383 , n8168 );
and ( n15432 , n11249 , n8166 );
nor ( n15433 , n15431 , n15432 );
xnor ( n15434 , n15433 , n8178 );
and ( n15435 , n15430 , n15434 );
xor ( n15436 , n15381 , n15385 );
xor ( n15437 , n15436 , n15388 );
and ( n15438 , n15434 , n15437 );
and ( n15439 , n15430 , n15437 );
or ( n15440 , n15435 , n15438 , n15439 );
and ( n15441 , n10554 , n7318 );
and ( n15442 , n10559 , n7315 );
nor ( n15443 , n15441 , n15442 );
xnor ( n15444 , n15443 , n7311 );
and ( n15445 , n15440 , n15444 );
xor ( n15446 , n15391 , n15395 );
xor ( n15447 , n15446 , n15398 );
and ( n15448 , n15444 , n15447 );
and ( n15449 , n15440 , n15447 );
or ( n15450 , n15445 , n15448 , n15449 );
and ( n15451 , n15417 , n15450 );
xor ( n15452 , n15417 , n15450 );
and ( n15453 , n11710 , n7395 );
and ( n15454 , n11697 , n7393 );
nor ( n15455 , n15453 , n15454 );
xnor ( n15456 , n15455 , n7405 );
and ( n15457 , n12012 , n7899 );
and ( n15458 , n11817 , n7897 );
nor ( n15459 , n15457 , n15458 );
xnor ( n15460 , n15459 , n7909 );
and ( n15461 , n15456 , n15460 );
and ( n15462 , n15460 , n15378 );
and ( n15463 , n15456 , n15378 );
or ( n15464 , n15461 , n15462 , n15463 );
and ( n15465 , n11435 , n8168 );
and ( n15466 , n11383 , n8166 );
nor ( n15467 , n15465 , n15466 );
xnor ( n15468 , n15467 , n8178 );
and ( n15469 , n15464 , n15468 );
xor ( n15470 , n15418 , n15422 );
xor ( n15471 , n15470 , n15427 );
and ( n15472 , n15468 , n15471 );
and ( n15473 , n15464 , n15471 );
or ( n15474 , n15469 , n15472 , n15473 );
and ( n15475 , n11187 , n7318 );
and ( n15476 , n10554 , n7315 );
nor ( n15477 , n15475 , n15476 );
xnor ( n15478 , n15477 , n7311 );
and ( n15479 , n15474 , n15478 );
xor ( n15480 , n15430 , n15434 );
xor ( n15481 , n15480 , n15437 );
and ( n15482 , n15478 , n15481 );
and ( n15483 , n15474 , n15481 );
or ( n15484 , n15479 , n15482 , n15483 );
xor ( n15485 , n15440 , n15444 );
xor ( n15486 , n15485 , n15447 );
and ( n15487 , n15484 , n15486 );
xor ( n15488 , n15484 , n15486 );
xor ( n15489 , n15474 , n15478 );
xor ( n15490 , n15489 , n15481 );
and ( n15491 , n11817 , n7395 );
and ( n15492 , n11710 , n7393 );
nor ( n15493 , n15491 , n15492 );
xnor ( n15494 , n15493 , n7405 );
and ( n15495 , n12246 , n7897 );
not ( n15496 , n15495 );
and ( n15497 , n15496 , n7909 );
and ( n15498 , n15494 , n15497 );
and ( n15499 , n11569 , n8168 );
and ( n15500 , n11435 , n8166 );
nor ( n15501 , n15499 , n15500 );
xnor ( n15502 , n15501 , n8178 );
and ( n15503 , n15498 , n15502 );
xor ( n15504 , n15456 , n15460 );
xor ( n15505 , n15504 , n15378 );
and ( n15506 , n15502 , n15505 );
and ( n15507 , n15498 , n15505 );
or ( n15508 , n15503 , n15506 , n15507 );
and ( n15509 , n11249 , n7318 );
and ( n15510 , n11187 , n7315 );
nor ( n15511 , n15509 , n15510 );
xnor ( n15512 , n15511 , n7311 );
and ( n15513 , n15508 , n15512 );
xor ( n15514 , n15464 , n15468 );
xor ( n15515 , n15514 , n15471 );
and ( n15516 , n15512 , n15515 );
and ( n15517 , n15508 , n15515 );
or ( n15518 , n15513 , n15516 , n15517 );
and ( n15519 , n15490 , n15518 );
xor ( n15520 , n15490 , n15518 );
xor ( n15521 , n15494 , n15497 );
and ( n15522 , n11697 , n8168 );
and ( n15523 , n11569 , n8166 );
nor ( n15524 , n15522 , n15523 );
xnor ( n15525 , n15524 , n8178 );
and ( n15526 , n15521 , n15525 );
and ( n15527 , n12246 , n7899 );
and ( n15528 , n12012 , n7897 );
nor ( n15529 , n15527 , n15528 );
xnor ( n15530 , n15529 , n7909 );
and ( n15531 , n15525 , n15530 );
and ( n15532 , n15521 , n15530 );
or ( n15533 , n15526 , n15531 , n15532 );
and ( n15534 , n11383 , n7318 );
and ( n15535 , n11249 , n7315 );
nor ( n15536 , n15534 , n15535 );
xnor ( n15537 , n15536 , n7311 );
and ( n15538 , n15533 , n15537 );
xor ( n15539 , n15498 , n15502 );
xor ( n15540 , n15539 , n15505 );
and ( n15541 , n15537 , n15540 );
and ( n15542 , n15533 , n15540 );
or ( n15543 , n15538 , n15541 , n15542 );
xor ( n15544 , n15508 , n15512 );
xor ( n15545 , n15544 , n15515 );
and ( n15546 , n15543 , n15545 );
xor ( n15547 , n15543 , n15545 );
xor ( n15548 , n15533 , n15537 );
xor ( n15549 , n15548 , n15540 );
and ( n15550 , n12246 , n7393 );
not ( n15551 , n15550 );
and ( n15552 , n15551 , n7405 );
and ( n15553 , n12246 , n7395 );
and ( n15554 , n12012 , n7393 );
nor ( n15555 , n15553 , n15554 );
xnor ( n15556 , n15555 , n7405 );
and ( n15557 , n15552 , n15556 );
and ( n15558 , n12012 , n7395 );
and ( n15559 , n11817 , n7393 );
nor ( n15560 , n15558 , n15559 );
xnor ( n15561 , n15560 , n7405 );
and ( n15562 , n15557 , n15561 );
and ( n15563 , n15561 , n15495 );
and ( n15564 , n15557 , n15495 );
or ( n15565 , n15562 , n15563 , n15564 );
and ( n15566 , n11435 , n7318 );
and ( n15567 , n11383 , n7315 );
nor ( n15568 , n15566 , n15567 );
xnor ( n15569 , n15568 , n7311 );
and ( n15570 , n15565 , n15569 );
xor ( n15571 , n15521 , n15525 );
xor ( n15572 , n15571 , n15530 );
and ( n15573 , n15569 , n15572 );
and ( n15574 , n15565 , n15572 );
or ( n15575 , n15570 , n15573 , n15574 );
and ( n15576 , n15549 , n15575 );
xor ( n15577 , n15549 , n15575 );
xor ( n15578 , n15565 , n15569 );
xor ( n15579 , n15578 , n15572 );
and ( n15580 , n11569 , n7318 );
and ( n15581 , n11435 , n7315 );
nor ( n15582 , n15580 , n15581 );
xnor ( n15583 , n15582 , n7311 );
and ( n15584 , n11710 , n8168 );
and ( n15585 , n11697 , n8166 );
nor ( n15586 , n15584 , n15585 );
xnor ( n15587 , n15586 , n8178 );
and ( n15588 , n15583 , n15587 );
xor ( n15589 , n15557 , n15561 );
xor ( n15590 , n15589 , n15495 );
and ( n15591 , n15587 , n15590 );
and ( n15592 , n15583 , n15590 );
or ( n15593 , n15588 , n15591 , n15592 );
and ( n15594 , n15579 , n15593 );
xor ( n15595 , n15579 , n15593 );
xor ( n15596 , n15583 , n15587 );
xor ( n15597 , n15596 , n15590 );
xor ( n15598 , n15552 , n15556 );
and ( n15599 , n12246 , n8166 );
not ( n15600 , n15599 );
and ( n15601 , n15600 , n8178 );
and ( n15602 , n12246 , n8168 );
and ( n15603 , n12012 , n8166 );
nor ( n15604 , n15602 , n15603 );
xnor ( n15605 , n15604 , n8178 );
and ( n15606 , n15601 , n15605 );
and ( n15607 , n12012 , n8168 );
and ( n15608 , n11817 , n8166 );
nor ( n15609 , n15607 , n15608 );
xnor ( n15610 , n15609 , n8178 );
and ( n15611 , n15606 , n15610 );
and ( n15612 , n15610 , n15550 );
and ( n15613 , n15606 , n15550 );
or ( n15614 , n15611 , n15612 , n15613 );
and ( n15615 , n15598 , n15614 );
and ( n15616 , n11817 , n8168 );
and ( n15617 , n11710 , n8166 );
nor ( n15618 , n15616 , n15617 );
xnor ( n15619 , n15618 , n8178 );
and ( n15620 , n15614 , n15619 );
and ( n15621 , n15598 , n15619 );
or ( n15622 , n15615 , n15620 , n15621 );
and ( n15623 , n15597 , n15622 );
xor ( n15624 , n15597 , n15622 );
and ( n15625 , n11697 , n7318 );
and ( n15626 , n11569 , n7315 );
nor ( n15627 , n15625 , n15626 );
xnor ( n15628 , n15627 , n7311 );
xor ( n15629 , n15598 , n15614 );
xor ( n15630 , n15629 , n15619 );
and ( n15631 , n15628 , n15630 );
xor ( n15632 , n15628 , n15630 );
and ( n15633 , n11710 , n7318 );
and ( n15634 , n11697 , n7315 );
nor ( n15635 , n15633 , n15634 );
xnor ( n15636 , n15635 , n7311 );
xor ( n15637 , n15606 , n15610 );
xor ( n15638 , n15637 , n15550 );
and ( n15639 , n15636 , n15638 );
xor ( n15640 , n15636 , n15638 );
and ( n15641 , n11817 , n7318 );
and ( n15642 , n11710 , n7315 );
nor ( n15643 , n15641 , n15642 );
xnor ( n15644 , n15643 , n7311 );
xor ( n15645 , n15601 , n15605 );
and ( n15646 , n15644 , n15645 );
xor ( n15647 , n15644 , n15645 );
and ( n15648 , n12012 , n7318 );
and ( n15649 , n11817 , n7315 );
nor ( n15650 , n15648 , n15649 );
xnor ( n15651 , n15650 , n7311 );
and ( n15652 , n15651 , n15599 );
xor ( n15653 , n15651 , n15599 );
and ( n15654 , n12246 , n7318 );
and ( n15655 , n12012 , n7315 );
nor ( n15656 , n15654 , n15655 );
xnor ( n15657 , n15656 , n7311 );
and ( n15658 , n12246 , n7315 );
not ( n15659 , n15658 );
and ( n15660 , n15659 , n7311 );
and ( n15661 , n15657 , n15660 );
and ( n15662 , n15653 , n15661 );
or ( n15663 , n15652 , n15662 );
and ( n15664 , n15647 , n15663 );
or ( n15665 , n15646 , n15664 );
and ( n15666 , n15640 , n15665 );
or ( n15667 , n15639 , n15666 );
and ( n15668 , n15632 , n15667 );
or ( n15669 , n15631 , n15668 );
and ( n15670 , n15624 , n15669 );
or ( n15671 , n15623 , n15670 );
and ( n15672 , n15595 , n15671 );
or ( n15673 , n15594 , n15672 );
and ( n15674 , n15577 , n15673 );
or ( n15675 , n15576 , n15674 );
and ( n15676 , n15547 , n15675 );
or ( n15677 , n15546 , n15676 );
and ( n15678 , n15520 , n15677 );
or ( n15679 , n15519 , n15678 );
and ( n15680 , n15488 , n15679 );
or ( n15681 , n15487 , n15680 );
and ( n15682 , n15452 , n15681 );
or ( n15683 , n15451 , n15682 );
and ( n15684 , n15415 , n15683 );
or ( n15685 , n15414 , n15684 );
and ( n15686 , n15373 , n15685 );
or ( n15687 , n15372 , n15686 );
and ( n15688 , n15327 , n15687 );
or ( n15689 , n15326 , n15688 );
and ( n15690 , n15282 , n15689 );
or ( n15691 , n15281 , n15690 );
and ( n15692 , n15230 , n15691 );
or ( n15693 , n15229 , n15692 );
and ( n15694 , n15174 , n15693 );
or ( n15695 , n15173 , n15694 );
and ( n15696 , n15119 , n15695 );
or ( n15697 , n15118 , n15696 );
and ( n15698 , n15057 , n15697 );
or ( n15699 , n15056 , n15698 );
and ( n15700 , n14993 , n15699 );
or ( n15701 , n14992 , n15700 );
and ( n15702 , n14926 , n15701 );
or ( n15703 , n14925 , n15702 );
and ( n15704 , n14814 , n15703 );
or ( n15705 , n14813 , n15704 );
and ( n15706 , n14751 , n15705 );
or ( n15707 , n14750 , n15706 );
and ( n15708 , n14657 , n15707 );
or ( n15709 , n14656 , n15708 );
and ( n15710 , n14585 , n15709 );
or ( n15711 , n14584 , n15710 );
and ( n15712 , n14498 , n15711 );
or ( n15713 , n14497 , n15712 );
and ( n15714 , n14386 , n15713 );
or ( n15715 , n14385 , n15714 );
and ( n15716 , n14287 , n15715 );
or ( n15717 , n14286 , n15716 );
and ( n15718 , n14221 , n15717 );
or ( n15719 , n14220 , n15718 );
and ( n15720 , n14028 , n15719 );
or ( n15721 , n14027 , n15720 );
and ( n15722 , n13986 , n15721 );
or ( n15723 , n13985 , n15722 );
and ( n15724 , n13801 , n15723 );
or ( n15725 , n13800 , n15724 );
and ( n15726 , n13719 , n15725 );
or ( n15727 , n13718 , n15726 );
and ( n15728 , n13565 , n15727 );
or ( n15729 , n13564 , n15728 );
and ( n15730 , n13380 , n15729 );
or ( n15731 , n13379 , n15730 );
and ( n15732 , n13278 , n15731 );
or ( n15733 , n13277 , n15732 );
and ( n15734 , n13073 , n15733 );
or ( n15735 , n13072 , n15734 );
and ( n15736 , n13051 , n15735 );
or ( n15737 , n13050 , n15736 );
and ( n15738 , n12736 , n15737 );
and ( n15739 , n12734 , n15738 );
and ( n15740 , n12732 , n15739 );
and ( n15741 , n12730 , n15740 );
and ( n15742 , n12728 , n15741 );
and ( n15743 , n12726 , n15742 );
or ( n15744 , n12725 , n15743 );
and ( n15745 , n11966 , n15744 );
or ( n15746 , n11965 , n15745 );
and ( n15747 , n11555 , n15746 );
and ( n15748 , n11553 , n15747 );
and ( n15749 , n11551 , n15748 );
and ( n15750 , n11549 , n15749 );
and ( n15751 , n11547 , n15750 );
or ( n15752 , n11546 , n15751 );
and ( n15753 , n10866 , n15752 );
and ( n15754 , n10864 , n15753 );
and ( n15755 , n10862 , n15754 );
and ( n15756 , n10860 , n15755 );
and ( n15757 , n10858 , n15756 );
or ( n15758 , n10857 , n15757 );
and ( n15759 , n9971 , n15758 );
and ( n15760 , n9969 , n15759 );
and ( n15761 , n9967 , n15760 );
and ( n15762 , n9965 , n15761 );
or ( n15763 , n9964 , n15762 );
and ( n15764 , n9362 , n15763 );
or ( n15765 , n9361 , n15764 );
and ( n15766 , n9145 , n15765 );
or ( n15767 , n9144 , n15766 );
xor ( n15768 , n8998 , n15767 );
buf ( n15769 , n15768 );
buf ( n15770 , n15769 );
xor ( n15771 , n9145 , n15765 );
buf ( n15772 , n15771 );
buf ( n15773 , n15772 );
xor ( n15774 , n9362 , n15763 );
buf ( n15775 , n15774 );
buf ( n15776 , n15775 );
xor ( n15777 , n9965 , n15761 );
buf ( n15778 , n15777 );
buf ( n15779 , n15778 );
xor ( n15780 , n9967 , n15760 );
buf ( n15781 , n15780 );
buf ( n15782 , n15781 );
xor ( n15783 , n9969 , n15759 );
buf ( n15784 , n15783 );
buf ( n15785 , n15784 );
xor ( n15786 , n9971 , n15758 );
buf ( n15787 , n15786 );
buf ( n15788 , n15787 );
xor ( n15789 , n10858 , n15756 );
buf ( n15790 , n15789 );
buf ( n15791 , n15790 );
xor ( n15792 , n10860 , n15755 );
buf ( n15793 , n15792 );
buf ( n15794 , n15793 );
xor ( n15795 , n10862 , n15754 );
buf ( n15796 , n15795 );
buf ( n15797 , n15796 );
xor ( n15798 , n10864 , n15753 );
buf ( n15799 , n15798 );
buf ( n15800 , n15799 );
xor ( n15801 , n10866 , n15752 );
buf ( n15802 , n15801 );
buf ( n15803 , n15802 );
xor ( n15804 , n11547 , n15750 );
buf ( n15805 , n15804 );
buf ( n15806 , n15805 );
xor ( n15807 , n11549 , n15749 );
buf ( n15808 , n15807 );
buf ( n15809 , n15808 );
xor ( n15810 , n11551 , n15748 );
buf ( n15811 , n15810 );
buf ( n15812 , n15811 );
xor ( n15813 , n11553 , n15747 );
buf ( n15814 , n15813 );
buf ( n15815 , n15814 );
xor ( n15816 , n11555 , n15746 );
buf ( n15817 , n15816 );
buf ( n15818 , n15817 );
xor ( n15819 , n11966 , n15744 );
buf ( n15820 , n15819 );
buf ( n15821 , n15820 );
xor ( n15822 , n12726 , n15742 );
buf ( n15823 , n15822 );
buf ( n15824 , n15823 );
xor ( n15825 , n12728 , n15741 );
buf ( n15826 , n15825 );
buf ( n15827 , n15826 );
xor ( n15828 , n12730 , n15740 );
buf ( n15829 , n15828 );
buf ( n15830 , n15829 );
xor ( n15831 , n12732 , n15739 );
buf ( n15832 , n15831 );
buf ( n15833 , n15832 );
xor ( n15834 , n12734 , n15738 );
buf ( n15835 , n15834 );
buf ( n15836 , n15835 );
xor ( n15837 , n12736 , n15737 );
buf ( n15838 , n15837 );
buf ( n15839 , n15838 );
xor ( n15840 , n13051 , n15735 );
buf ( n15841 , n15840 );
buf ( n15842 , n15841 );
xor ( n15843 , n13073 , n15733 );
buf ( n15844 , n15843 );
buf ( n15845 , n15844 );
xor ( n15846 , n13278 , n15731 );
buf ( n15847 , n15846 );
buf ( n15848 , n15847 );
xor ( n15849 , n13380 , n15729 );
buf ( n15850 , n15849 );
buf ( n15851 , n15850 );
xor ( n15852 , n13565 , n15727 );
buf ( n15853 , n15852 );
buf ( n15854 , n15853 );
xor ( n15855 , n13719 , n15725 );
buf ( n15856 , n15855 );
buf ( n15857 , n15856 );
xor ( n15858 , n13801 , n15723 );
buf ( n15859 , n15858 );
buf ( n15860 , n15859 );
xor ( n15861 , n13986 , n15721 );
buf ( n15862 , n15861 );
buf ( n15863 , n15862 );
xor ( n15864 , n14028 , n15719 );
buf ( n15865 , n15864 );
buf ( n15866 , n15865 );
xor ( n15867 , n14221 , n15717 );
buf ( n15868 , n15867 );
buf ( n15869 , n15868 );
xor ( n15870 , n14287 , n15715 );
buf ( n15871 , n15870 );
buf ( n15872 , n15871 );
xor ( n15873 , n14386 , n15713 );
buf ( n15874 , n15873 );
buf ( n15875 , n15874 );
xor ( n15876 , n14498 , n15711 );
buf ( n15877 , n15876 );
buf ( n15878 , n15877 );
xor ( n15879 , n14585 , n15709 );
buf ( n15880 , n15879 );
buf ( n15881 , n15880 );
xor ( n15882 , n14657 , n15707 );
buf ( n15883 , n15882 );
buf ( n15884 , n15883 );
xor ( n15885 , n14751 , n15705 );
buf ( n15886 , n15885 );
buf ( n15887 , n15886 );
xor ( n15888 , n14814 , n15703 );
buf ( n15889 , n15888 );
buf ( n15890 , n15889 );
xor ( n15891 , n14926 , n15701 );
buf ( n15892 , n15891 );
buf ( n15893 , n15892 );
xor ( n15894 , n14993 , n15699 );
buf ( n15895 , n15894 );
buf ( n15896 , n15895 );
xor ( n15897 , n15057 , n15697 );
buf ( n15898 , n15897 );
buf ( n15899 , n15898 );
xor ( n15900 , n15119 , n15695 );
buf ( n15901 , n15900 );
buf ( n15902 , n15901 );
xor ( n15903 , n15174 , n15693 );
buf ( n15904 , n15903 );
buf ( n15905 , n15904 );
xor ( n15906 , n15230 , n15691 );
buf ( n15907 , n15906 );
buf ( n15908 , n15907 );
xor ( n15909 , n15282 , n15689 );
buf ( n15910 , n15909 );
buf ( n15911 , n15910 );
xor ( n15912 , n15327 , n15687 );
buf ( n15913 , n15912 );
buf ( n15914 , n15913 );
xor ( n15915 , n15373 , n15685 );
buf ( n15916 , n15915 );
buf ( n15917 , n15916 );
xor ( n15918 , n15415 , n15683 );
buf ( n15919 , n15918 );
buf ( n15920 , n15919 );
xor ( n15921 , n15452 , n15681 );
buf ( n15922 , n15921 );
buf ( n15923 , n15922 );
xor ( n15924 , n15488 , n15679 );
buf ( n15925 , n15924 );
buf ( n15926 , n15925 );
xor ( n15927 , n15520 , n15677 );
buf ( n15928 , n15927 );
buf ( n15929 , n15928 );
xor ( n15930 , n15547 , n15675 );
buf ( n15931 , n15930 );
buf ( n15932 , n15931 );
xor ( n15933 , n15577 , n15673 );
buf ( n15934 , n15933 );
buf ( n15935 , n15934 );
xor ( n15936 , n15595 , n15671 );
buf ( n15937 , n15936 );
buf ( n15938 , n15937 );
xor ( n15939 , n15624 , n15669 );
buf ( n15940 , n15939 );
buf ( n15941 , n15940 );
xor ( n15942 , n15632 , n15667 );
buf ( n15943 , n15942 );
buf ( n15944 , n15943 );
xor ( n15945 , n15640 , n15665 );
buf ( n15946 , n15945 );
buf ( n15947 , n15946 );
xor ( n15948 , n15647 , n15663 );
buf ( n15949 , n15948 );
buf ( n15950 , n15949 );
xor ( n15951 , n15653 , n15661 );
buf ( n15952 , n15951 );
buf ( n15953 , n15952 );
xor ( n15954 , n15657 , n15660 );
buf ( n15955 , n15954 );
buf ( n15956 , n15955 );
buf ( n15957 , n15658 );
buf ( n15958 , n15957 );
buf ( n15959 , n15958 );
buf ( n15960 , n1097 );
buf ( n15961 , n15960 );
buf ( n15962 , n1160 );
buf ( n15963 , n15962 );
buf ( n15964 , n1161 );
buf ( n15965 , n15964 );
xor ( n15966 , n15963 , n15965 );
buf ( n15967 , n1162 );
buf ( n15968 , n15967 );
xor ( n15969 , n15965 , n15968 );
not ( n15970 , n15969 );
and ( n15971 , n15966 , n15970 );
and ( n15972 , n15961 , n15971 );
buf ( n15973 , n1096 );
buf ( n15974 , n15973 );
and ( n15975 , n15974 , n15969 );
nor ( n15976 , n15972 , n15975 );
and ( n15977 , n15965 , n15968 );
not ( n15978 , n15977 );
and ( n15979 , n15963 , n15978 );
xnor ( n15980 , n15976 , n15979 );
buf ( n15981 , n1103 );
buf ( n15982 , n15981 );
buf ( n15983 , n1154 );
buf ( n15984 , n15983 );
buf ( n15985 , n1155 );
buf ( n15986 , n15985 );
xor ( n15987 , n15984 , n15986 );
buf ( n15988 , n1156 );
buf ( n15989 , n15988 );
xor ( n15990 , n15986 , n15989 );
not ( n15991 , n15990 );
and ( n15992 , n15987 , n15991 );
and ( n15993 , n15982 , n15992 );
buf ( n15994 , n1102 );
buf ( n15995 , n15994 );
and ( n15996 , n15995 , n15990 );
nor ( n15997 , n15993 , n15996 );
and ( n15998 , n15986 , n15989 );
not ( n15999 , n15998 );
and ( n16000 , n15984 , n15999 );
xnor ( n16001 , n15997 , n16000 );
xor ( n16002 , n15980 , n16001 );
buf ( n16003 , n1104 );
buf ( n16004 , n16003 );
and ( n16005 , n16004 , n15984 );
xor ( n16006 , n16002 , n16005 );
buf ( n16007 , n1093 );
buf ( n16008 , n16007 );
buf ( n16009 , n1164 );
buf ( n16010 , n16009 );
buf ( n16011 , n1165 );
buf ( n16012 , n16011 );
xor ( n16013 , n16010 , n16012 );
buf ( n16014 , n1166 );
buf ( n16015 , n16014 );
xor ( n16016 , n16012 , n16015 );
not ( n16017 , n16016 );
and ( n16018 , n16013 , n16017 );
and ( n16019 , n16008 , n16018 );
buf ( n16020 , n1092 );
buf ( n16021 , n16020 );
and ( n16022 , n16021 , n16016 );
nor ( n16023 , n16019 , n16022 );
and ( n16024 , n16012 , n16015 );
not ( n16025 , n16024 );
and ( n16026 , n16010 , n16025 );
xnor ( n16027 , n16023 , n16026 );
buf ( n16028 , n1099 );
buf ( n16029 , n16028 );
buf ( n16030 , n1158 );
buf ( n16031 , n16030 );
buf ( n16032 , n1159 );
buf ( n16033 , n16032 );
xor ( n16034 , n16031 , n16033 );
xor ( n16035 , n16033 , n15963 );
not ( n16036 , n16035 );
and ( n16037 , n16034 , n16036 );
and ( n16038 , n16029 , n16037 );
buf ( n16039 , n1098 );
buf ( n16040 , n16039 );
and ( n16041 , n16040 , n16035 );
nor ( n16042 , n16038 , n16041 );
and ( n16043 , n16033 , n15963 );
not ( n16044 , n16043 );
and ( n16045 , n16031 , n16044 );
xnor ( n16046 , n16042 , n16045 );
xor ( n16047 , n16027 , n16046 );
buf ( n16048 , n1101 );
buf ( n16049 , n16048 );
buf ( n16050 , n1157 );
buf ( n16051 , n16050 );
xor ( n16052 , n15989 , n16051 );
xor ( n16053 , n16051 , n16031 );
not ( n16054 , n16053 );
and ( n16055 , n16052 , n16054 );
and ( n16056 , n16049 , n16055 );
buf ( n16057 , n1100 );
buf ( n16058 , n16057 );
and ( n16059 , n16058 , n16053 );
nor ( n16060 , n16056 , n16059 );
and ( n16061 , n16051 , n16031 );
not ( n16062 , n16061 );
and ( n16063 , n15989 , n16062 );
xnor ( n16064 , n16060 , n16063 );
xor ( n16065 , n16047 , n16064 );
and ( n16066 , n16006 , n16065 );
buf ( n16067 , n1168 );
buf ( n16068 , n16067 );
buf ( n16069 , n1169 );
buf ( n16070 , n16069 );
buf ( n16071 , n1170 );
buf ( n16072 , n16071 );
and ( n16073 , n16070 , n16072 );
not ( n16074 , n16073 );
and ( n16075 , n16068 , n16074 );
not ( n16076 , n16075 );
buf ( n16077 , n1091 );
buf ( n16078 , n16077 );
buf ( n16079 , n1167 );
buf ( n16080 , n16079 );
xor ( n16081 , n16015 , n16080 );
xor ( n16082 , n16080 , n16068 );
not ( n16083 , n16082 );
and ( n16084 , n16081 , n16083 );
and ( n16085 , n16078 , n16084 );
buf ( n16086 , n1090 );
buf ( n16087 , n16086 );
and ( n16088 , n16087 , n16082 );
nor ( n16089 , n16085 , n16088 );
and ( n16090 , n16080 , n16068 );
not ( n16091 , n16090 );
and ( n16092 , n16015 , n16091 );
xnor ( n16093 , n16089 , n16092 );
xor ( n16094 , n16076 , n16093 );
buf ( n16095 , n1095 );
buf ( n16096 , n16095 );
buf ( n16097 , n1163 );
buf ( n16098 , n16097 );
xor ( n16099 , n15968 , n16098 );
xor ( n16100 , n16098 , n16010 );
not ( n16101 , n16100 );
and ( n16102 , n16099 , n16101 );
and ( n16103 , n16096 , n16102 );
buf ( n16104 , n1094 );
buf ( n16105 , n16104 );
and ( n16106 , n16105 , n16100 );
nor ( n16107 , n16103 , n16106 );
and ( n16108 , n16098 , n16010 );
not ( n16109 , n16108 );
and ( n16110 , n15968 , n16109 );
xnor ( n16111 , n16107 , n16110 );
xor ( n16112 , n16094 , n16111 );
and ( n16113 , n16065 , n16112 );
and ( n16114 , n16006 , n16112 );
or ( n16115 , n16066 , n16113 , n16114 );
and ( n16116 , n15980 , n16001 );
and ( n16117 , n16001 , n16005 );
and ( n16118 , n15980 , n16005 );
or ( n16119 , n16116 , n16117 , n16118 );
and ( n16120 , n16027 , n16046 );
and ( n16121 , n16046 , n16064 );
and ( n16122 , n16027 , n16064 );
or ( n16123 , n16120 , n16121 , n16122 );
xor ( n16124 , n16119 , n16123 );
and ( n16125 , n16105 , n16102 );
and ( n16126 , n16008 , n16100 );
nor ( n16127 , n16125 , n16126 );
xnor ( n16128 , n16127 , n16110 );
and ( n16129 , n16040 , n16037 );
and ( n16130 , n15961 , n16035 );
nor ( n16131 , n16129 , n16130 );
xnor ( n16132 , n16131 , n16045 );
xor ( n16133 , n16128 , n16132 );
and ( n16134 , n16058 , n16055 );
and ( n16135 , n16029 , n16053 );
nor ( n16136 , n16134 , n16135 );
xnor ( n16137 , n16136 , n16063 );
xor ( n16138 , n16133 , n16137 );
xor ( n16139 , n16124 , n16138 );
and ( n16140 , n16115 , n16139 );
and ( n16141 , n15974 , n16102 );
and ( n16142 , n16096 , n16100 );
nor ( n16143 , n16141 , n16142 );
xnor ( n16144 , n16143 , n16110 );
and ( n16145 , n16004 , n15992 );
and ( n16146 , n15982 , n15990 );
nor ( n16147 , n16145 , n16146 );
xnor ( n16148 , n16147 , n16000 );
and ( n16149 , n16144 , n16148 );
buf ( n16150 , n1105 );
buf ( n16151 , n16150 );
and ( n16152 , n16151 , n15984 );
and ( n16153 , n16148 , n16152 );
and ( n16154 , n16144 , n16152 );
or ( n16155 , n16149 , n16153 , n16154 );
and ( n16156 , n16021 , n16084 );
and ( n16157 , n16078 , n16082 );
nor ( n16158 , n16156 , n16157 );
xnor ( n16159 , n16158 , n16092 );
and ( n16160 , n16105 , n16018 );
and ( n16161 , n16008 , n16016 );
nor ( n16162 , n16160 , n16161 );
xnor ( n16163 , n16162 , n16026 );
and ( n16164 , n16159 , n16163 );
and ( n16165 , n16040 , n15971 );
and ( n16166 , n15961 , n15969 );
nor ( n16167 , n16165 , n16166 );
xnor ( n16168 , n16167 , n15979 );
and ( n16169 , n16163 , n16168 );
and ( n16170 , n16159 , n16168 );
or ( n16171 , n16164 , n16169 , n16170 );
and ( n16172 , n16155 , n16171 );
xor ( n16173 , n16068 , n16070 );
xor ( n16174 , n16070 , n16072 );
not ( n16175 , n16174 );
and ( n16176 , n16173 , n16175 );
and ( n16177 , n16087 , n16176 );
not ( n16178 , n16177 );
xnor ( n16179 , n16178 , n16075 );
buf ( n16180 , n16179 );
and ( n16181 , n16171 , n16180 );
and ( n16182 , n16155 , n16180 );
or ( n16183 , n16172 , n16181 , n16182 );
and ( n16184 , n16021 , n16018 );
and ( n16185 , n16078 , n16016 );
nor ( n16186 , n16184 , n16185 );
xnor ( n16187 , n16186 , n16026 );
and ( n16188 , n15974 , n15971 );
and ( n16189 , n16096 , n15969 );
nor ( n16190 , n16188 , n16189 );
xnor ( n16191 , n16190 , n15979 );
xor ( n16192 , n16187 , n16191 );
and ( n16193 , n15982 , n15984 );
xor ( n16194 , n16192 , n16193 );
xor ( n16195 , n16183 , n16194 );
and ( n16196 , n16076 , n16093 );
and ( n16197 , n16093 , n16111 );
and ( n16198 , n16076 , n16111 );
or ( n16199 , n16196 , n16197 , n16198 );
and ( n16200 , n16087 , n16084 );
not ( n16201 , n16200 );
xnor ( n16202 , n16201 , n16092 );
not ( n16203 , n16202 );
xor ( n16204 , n16199 , n16203 );
and ( n16205 , n15995 , n15992 );
and ( n16206 , n16049 , n15990 );
nor ( n16207 , n16205 , n16206 );
xnor ( n16208 , n16207 , n16000 );
xor ( n16209 , n16204 , n16208 );
xor ( n16210 , n16195 , n16209 );
and ( n16211 , n16139 , n16210 );
and ( n16212 , n16115 , n16210 );
or ( n16213 , n16140 , n16211 , n16212 );
and ( n16214 , n16199 , n16203 );
and ( n16215 , n16203 , n16208 );
and ( n16216 , n16199 , n16208 );
or ( n16217 , n16214 , n16215 , n16216 );
and ( n16218 , n16008 , n16102 );
and ( n16219 , n16021 , n16100 );
nor ( n16220 , n16218 , n16219 );
xnor ( n16221 , n16220 , n16110 );
and ( n16222 , n15961 , n16037 );
and ( n16223 , n15974 , n16035 );
nor ( n16224 , n16222 , n16223 );
xnor ( n16225 , n16224 , n16045 );
xor ( n16226 , n16221 , n16225 );
and ( n16227 , n15995 , n15984 );
xor ( n16228 , n16226 , n16227 );
xor ( n16229 , n16217 , n16228 );
buf ( n16230 , n16202 );
and ( n16231 , n16029 , n16055 );
and ( n16232 , n16040 , n16053 );
nor ( n16233 , n16231 , n16232 );
xnor ( n16234 , n16233 , n16063 );
xor ( n16235 , n16230 , n16234 );
and ( n16236 , n16049 , n15992 );
and ( n16237 , n16058 , n15990 );
nor ( n16238 , n16236 , n16237 );
xnor ( n16239 , n16238 , n16000 );
xor ( n16240 , n16235 , n16239 );
xor ( n16241 , n16229 , n16240 );
xor ( n16242 , n16213 , n16241 );
and ( n16243 , n16119 , n16123 );
and ( n16244 , n16123 , n16138 );
and ( n16245 , n16119 , n16138 );
or ( n16246 , n16243 , n16244 , n16245 );
and ( n16247 , n16183 , n16194 );
and ( n16248 , n16194 , n16209 );
and ( n16249 , n16183 , n16209 );
or ( n16250 , n16247 , n16248 , n16249 );
xor ( n16251 , n16246 , n16250 );
and ( n16252 , n16128 , n16132 );
and ( n16253 , n16132 , n16137 );
and ( n16254 , n16128 , n16137 );
or ( n16255 , n16252 , n16253 , n16254 );
and ( n16256 , n16187 , n16191 );
and ( n16257 , n16191 , n16193 );
and ( n16258 , n16187 , n16193 );
or ( n16259 , n16256 , n16257 , n16258 );
xor ( n16260 , n16255 , n16259 );
not ( n16261 , n16092 );
and ( n16262 , n16078 , n16018 );
and ( n16263 , n16087 , n16016 );
nor ( n16264 , n16262 , n16263 );
xnor ( n16265 , n16264 , n16026 );
xor ( n16266 , n16261 , n16265 );
and ( n16267 , n16096 , n15971 );
and ( n16268 , n16105 , n15969 );
nor ( n16269 , n16267 , n16268 );
xnor ( n16270 , n16269 , n15979 );
xor ( n16271 , n16266 , n16270 );
xor ( n16272 , n16260 , n16271 );
xor ( n16273 , n16251 , n16272 );
xor ( n16274 , n16242 , n16273 );
and ( n16275 , n16008 , n16084 );
and ( n16276 , n16021 , n16082 );
nor ( n16277 , n16275 , n16276 );
xnor ( n16278 , n16277 , n16092 );
and ( n16279 , n16029 , n15971 );
and ( n16280 , n16040 , n15969 );
nor ( n16281 , n16279 , n16280 );
xnor ( n16282 , n16281 , n15979 );
and ( n16283 , n16278 , n16282 );
buf ( n16284 , n1106 );
buf ( n16285 , n16284 );
and ( n16286 , n16285 , n15984 );
and ( n16287 , n16282 , n16286 );
and ( n16288 , n16278 , n16286 );
or ( n16289 , n16283 , n16287 , n16288 );
and ( n16290 , n15961 , n16102 );
and ( n16291 , n15974 , n16100 );
nor ( n16292 , n16290 , n16291 );
xnor ( n16293 , n16292 , n16110 );
and ( n16294 , n15982 , n16055 );
and ( n16295 , n15995 , n16053 );
nor ( n16296 , n16294 , n16295 );
xnor ( n16297 , n16296 , n16063 );
and ( n16298 , n16293 , n16297 );
and ( n16299 , n16151 , n15992 );
and ( n16300 , n16004 , n15990 );
nor ( n16301 , n16299 , n16300 );
xnor ( n16302 , n16301 , n16000 );
and ( n16303 , n16297 , n16302 );
and ( n16304 , n16293 , n16302 );
or ( n16305 , n16298 , n16303 , n16304 );
and ( n16306 , n16289 , n16305 );
buf ( n16307 , n1171 );
buf ( n16308 , n16307 );
buf ( n16309 , n1172 );
buf ( n16310 , n16309 );
and ( n16311 , n16308 , n16310 );
not ( n16312 , n16311 );
and ( n16313 , n16072 , n16312 );
not ( n16314 , n16313 );
and ( n16315 , n16078 , n16176 );
and ( n16316 , n16087 , n16174 );
nor ( n16317 , n16315 , n16316 );
xnor ( n16318 , n16317 , n16075 );
and ( n16319 , n16314 , n16318 );
and ( n16320 , n16096 , n16018 );
and ( n16321 , n16105 , n16016 );
nor ( n16322 , n16320 , n16321 );
xnor ( n16323 , n16322 , n16026 );
and ( n16324 , n16318 , n16323 );
and ( n16325 , n16314 , n16323 );
or ( n16326 , n16319 , n16324 , n16325 );
and ( n16327 , n16305 , n16326 );
and ( n16328 , n16289 , n16326 );
or ( n16329 , n16306 , n16327 , n16328 );
not ( n16330 , n16179 );
and ( n16331 , n16058 , n16037 );
and ( n16332 , n16029 , n16035 );
nor ( n16333 , n16331 , n16332 );
xnor ( n16334 , n16333 , n16045 );
and ( n16335 , n16330 , n16334 );
and ( n16336 , n15995 , n16055 );
and ( n16337 , n16049 , n16053 );
nor ( n16338 , n16336 , n16337 );
xnor ( n16339 , n16338 , n16063 );
and ( n16340 , n16334 , n16339 );
and ( n16341 , n16330 , n16339 );
or ( n16342 , n16335 , n16340 , n16341 );
and ( n16343 , n16329 , n16342 );
xor ( n16344 , n16155 , n16171 );
xor ( n16345 , n16344 , n16180 );
and ( n16346 , n16342 , n16345 );
and ( n16347 , n16329 , n16345 );
or ( n16348 , n16343 , n16346 , n16347 );
xor ( n16349 , n16144 , n16148 );
xor ( n16350 , n16349 , n16152 );
xor ( n16351 , n16159 , n16163 );
xor ( n16352 , n16351 , n16168 );
and ( n16353 , n16350 , n16352 );
xor ( n16354 , n16330 , n16334 );
xor ( n16355 , n16354 , n16339 );
and ( n16356 , n16352 , n16355 );
and ( n16357 , n16350 , n16355 );
or ( n16358 , n16353 , n16356 , n16357 );
and ( n16359 , n15974 , n16018 );
and ( n16360 , n16096 , n16016 );
nor ( n16361 , n16359 , n16360 );
xnor ( n16362 , n16361 , n16026 );
and ( n16363 , n16004 , n16055 );
and ( n16364 , n15982 , n16053 );
nor ( n16365 , n16363 , n16364 );
xnor ( n16366 , n16365 , n16063 );
and ( n16367 , n16362 , n16366 );
and ( n16368 , n16285 , n15992 );
and ( n16369 , n16151 , n15990 );
nor ( n16370 , n16368 , n16369 );
xnor ( n16371 , n16370 , n16000 );
and ( n16372 , n16366 , n16371 );
and ( n16373 , n16362 , n16371 );
or ( n16374 , n16367 , n16372 , n16373 );
xor ( n16375 , n16072 , n16308 );
xor ( n16376 , n16308 , n16310 );
not ( n16377 , n16376 );
and ( n16378 , n16375 , n16377 );
and ( n16379 , n16087 , n16378 );
not ( n16380 , n16379 );
xnor ( n16381 , n16380 , n16313 );
buf ( n16382 , n16381 );
and ( n16383 , n16374 , n16382 );
and ( n16384 , n16049 , n16037 );
and ( n16385 , n16058 , n16035 );
nor ( n16386 , n16384 , n16385 );
xnor ( n16387 , n16386 , n16045 );
and ( n16388 , n16382 , n16387 );
and ( n16389 , n16374 , n16387 );
or ( n16390 , n16383 , n16388 , n16389 );
and ( n16391 , n16021 , n16176 );
and ( n16392 , n16078 , n16174 );
nor ( n16393 , n16391 , n16392 );
xnor ( n16394 , n16393 , n16075 );
and ( n16395 , n16040 , n16102 );
and ( n16396 , n15961 , n16100 );
nor ( n16397 , n16395 , n16396 );
xnor ( n16398 , n16397 , n16110 );
and ( n16399 , n16394 , n16398 );
buf ( n16400 , n1107 );
buf ( n16401 , n16400 );
and ( n16402 , n16401 , n15984 );
and ( n16403 , n16398 , n16402 );
and ( n16404 , n16394 , n16402 );
or ( n16405 , n16399 , n16403 , n16404 );
and ( n16406 , n16105 , n16084 );
and ( n16407 , n16008 , n16082 );
nor ( n16408 , n16406 , n16407 );
xnor ( n16409 , n16408 , n16092 );
and ( n16410 , n16058 , n15971 );
and ( n16411 , n16029 , n15969 );
nor ( n16412 , n16410 , n16411 );
xnor ( n16413 , n16412 , n15979 );
and ( n16414 , n16409 , n16413 );
and ( n16415 , n15995 , n16037 );
and ( n16416 , n16049 , n16035 );
nor ( n16417 , n16415 , n16416 );
xnor ( n16418 , n16417 , n16045 );
and ( n16419 , n16413 , n16418 );
and ( n16420 , n16409 , n16418 );
or ( n16421 , n16414 , n16419 , n16420 );
and ( n16422 , n16405 , n16421 );
xor ( n16423 , n16278 , n16282 );
xor ( n16424 , n16423 , n16286 );
and ( n16425 , n16421 , n16424 );
and ( n16426 , n16405 , n16424 );
or ( n16427 , n16422 , n16425 , n16426 );
and ( n16428 , n16390 , n16427 );
xor ( n16429 , n16289 , n16305 );
xor ( n16430 , n16429 , n16326 );
and ( n16431 , n16427 , n16430 );
and ( n16432 , n16390 , n16430 );
or ( n16433 , n16428 , n16431 , n16432 );
and ( n16434 , n16358 , n16433 );
xor ( n16435 , n16006 , n16065 );
xor ( n16436 , n16435 , n16112 );
and ( n16437 , n16433 , n16436 );
and ( n16438 , n16358 , n16436 );
or ( n16439 , n16434 , n16437 , n16438 );
and ( n16440 , n16348 , n16439 );
xor ( n16441 , n16115 , n16139 );
xor ( n16442 , n16441 , n16210 );
and ( n16443 , n16439 , n16442 );
and ( n16444 , n16348 , n16442 );
or ( n16445 , n16440 , n16443 , n16444 );
xor ( n16446 , n16274 , n16445 );
xor ( n16447 , n16348 , n16439 );
xor ( n16448 , n16447 , n16442 );
xor ( n16449 , n16293 , n16297 );
xor ( n16450 , n16449 , n16302 );
xor ( n16451 , n16314 , n16318 );
xor ( n16452 , n16451 , n16323 );
and ( n16453 , n16450 , n16452 );
xor ( n16454 , n16374 , n16382 );
xor ( n16455 , n16454 , n16387 );
and ( n16456 , n16452 , n16455 );
and ( n16457 , n16450 , n16455 );
or ( n16458 , n16453 , n16456 , n16457 );
and ( n16459 , n15961 , n16018 );
and ( n16460 , n15974 , n16016 );
nor ( n16461 , n16459 , n16460 );
xnor ( n16462 , n16461 , n16026 );
and ( n16463 , n15982 , n16037 );
and ( n16464 , n15995 , n16035 );
nor ( n16465 , n16463 , n16464 );
xnor ( n16466 , n16465 , n16045 );
and ( n16467 , n16462 , n16466 );
and ( n16468 , n16151 , n16055 );
and ( n16469 , n16004 , n16053 );
nor ( n16470 , n16468 , n16469 );
xnor ( n16471 , n16470 , n16063 );
and ( n16472 , n16466 , n16471 );
and ( n16473 , n16462 , n16471 );
or ( n16474 , n16467 , n16472 , n16473 );
buf ( n16475 , n1173 );
buf ( n16476 , n16475 );
buf ( n16477 , n1174 );
buf ( n16478 , n16477 );
and ( n16479 , n16476 , n16478 );
not ( n16480 , n16479 );
and ( n16481 , n16310 , n16480 );
not ( n16482 , n16481 );
and ( n16483 , n16078 , n16378 );
and ( n16484 , n16087 , n16376 );
nor ( n16485 , n16483 , n16484 );
xnor ( n16486 , n16485 , n16313 );
and ( n16487 , n16482 , n16486 );
and ( n16488 , n16096 , n16084 );
and ( n16489 , n16105 , n16082 );
nor ( n16490 , n16488 , n16489 );
xnor ( n16491 , n16490 , n16092 );
and ( n16492 , n16486 , n16491 );
and ( n16493 , n16482 , n16491 );
or ( n16494 , n16487 , n16492 , n16493 );
and ( n16495 , n16474 , n16494 );
not ( n16496 , n16381 );
and ( n16497 , n16494 , n16496 );
and ( n16498 , n16474 , n16496 );
or ( n16499 , n16495 , n16497 , n16498 );
and ( n16500 , n16008 , n16176 );
and ( n16501 , n16021 , n16174 );
nor ( n16502 , n16500 , n16501 );
xnor ( n16503 , n16502 , n16075 );
and ( n16504 , n16401 , n15992 );
and ( n16505 , n16285 , n15990 );
nor ( n16506 , n16504 , n16505 );
xnor ( n16507 , n16506 , n16000 );
and ( n16508 , n16503 , n16507 );
buf ( n16509 , n1108 );
buf ( n16510 , n16509 );
and ( n16511 , n16510 , n15984 );
and ( n16512 , n16507 , n16511 );
and ( n16513 , n16503 , n16511 );
or ( n16514 , n16508 , n16512 , n16513 );
xor ( n16515 , n16394 , n16398 );
xor ( n16516 , n16515 , n16402 );
and ( n16517 , n16514 , n16516 );
xor ( n16518 , n16362 , n16366 );
xor ( n16519 , n16518 , n16371 );
and ( n16520 , n16516 , n16519 );
and ( n16521 , n16514 , n16519 );
or ( n16522 , n16517 , n16520 , n16521 );
and ( n16523 , n16499 , n16522 );
xor ( n16524 , n16405 , n16421 );
xor ( n16525 , n16524 , n16424 );
and ( n16526 , n16522 , n16525 );
and ( n16527 , n16499 , n16525 );
or ( n16528 , n16523 , n16526 , n16527 );
and ( n16529 , n16458 , n16528 );
xor ( n16530 , n16350 , n16352 );
xor ( n16531 , n16530 , n16355 );
and ( n16532 , n16528 , n16531 );
and ( n16533 , n16458 , n16531 );
or ( n16534 , n16529 , n16532 , n16533 );
xor ( n16535 , n16329 , n16342 );
xor ( n16536 , n16535 , n16345 );
and ( n16537 , n16534 , n16536 );
xor ( n16538 , n16358 , n16433 );
xor ( n16539 , n16538 , n16436 );
and ( n16540 , n16536 , n16539 );
and ( n16541 , n16534 , n16539 );
or ( n16542 , n16537 , n16540 , n16541 );
and ( n16543 , n16448 , n16542 );
xor ( n16544 , n16534 , n16536 );
xor ( n16545 , n16544 , n16539 );
and ( n16546 , n15974 , n16084 );
and ( n16547 , n16096 , n16082 );
nor ( n16548 , n16546 , n16547 );
xnor ( n16549 , n16548 , n16092 );
and ( n16550 , n16004 , n16037 );
and ( n16551 , n15982 , n16035 );
nor ( n16552 , n16550 , n16551 );
xnor ( n16553 , n16552 , n16045 );
and ( n16554 , n16549 , n16553 );
and ( n16555 , n16285 , n16055 );
and ( n16556 , n16151 , n16053 );
nor ( n16557 , n16555 , n16556 );
xnor ( n16558 , n16557 , n16063 );
and ( n16559 , n16553 , n16558 );
and ( n16560 , n16549 , n16558 );
or ( n16561 , n16554 , n16559 , n16560 );
xor ( n16562 , n16310 , n16476 );
xor ( n16563 , n16476 , n16478 );
not ( n16564 , n16563 );
and ( n16565 , n16562 , n16564 );
and ( n16566 , n16087 , n16565 );
not ( n16567 , n16566 );
xnor ( n16568 , n16567 , n16481 );
and ( n16569 , n16105 , n16176 );
and ( n16570 , n16008 , n16174 );
nor ( n16571 , n16569 , n16570 );
xnor ( n16572 , n16571 , n16075 );
and ( n16573 , n16568 , n16572 );
and ( n16574 , n16058 , n16102 );
and ( n16575 , n16029 , n16100 );
nor ( n16576 , n16574 , n16575 );
xnor ( n16577 , n16576 , n16110 );
and ( n16578 , n16572 , n16577 );
and ( n16579 , n16568 , n16577 );
or ( n16580 , n16573 , n16578 , n16579 );
and ( n16581 , n16561 , n16580 );
and ( n16582 , n16040 , n16018 );
and ( n16583 , n15961 , n16016 );
nor ( n16584 , n16582 , n16583 );
xnor ( n16585 , n16584 , n16026 );
and ( n16586 , n16510 , n15992 );
and ( n16587 , n16401 , n15990 );
nor ( n16588 , n16586 , n16587 );
xnor ( n16589 , n16588 , n16000 );
and ( n16590 , n16585 , n16589 );
buf ( n16591 , n1109 );
buf ( n16592 , n16591 );
and ( n16593 , n16592 , n15984 );
and ( n16594 , n16589 , n16593 );
and ( n16595 , n16585 , n16593 );
or ( n16596 , n16590 , n16594 , n16595 );
and ( n16597 , n16580 , n16596 );
and ( n16598 , n16561 , n16596 );
or ( n16599 , n16581 , n16597 , n16598 );
and ( n16600 , n16021 , n16378 );
and ( n16601 , n16078 , n16376 );
nor ( n16602 , n16600 , n16601 );
xnor ( n16603 , n16602 , n16313 );
buf ( n16604 , n16603 );
and ( n16605 , n16029 , n16102 );
and ( n16606 , n16040 , n16100 );
nor ( n16607 , n16605 , n16606 );
xnor ( n16608 , n16607 , n16110 );
and ( n16609 , n16604 , n16608 );
and ( n16610 , n16049 , n15971 );
and ( n16611 , n16058 , n15969 );
nor ( n16612 , n16610 , n16611 );
xnor ( n16613 , n16612 , n15979 );
and ( n16614 , n16608 , n16613 );
and ( n16615 , n16604 , n16613 );
or ( n16616 , n16609 , n16614 , n16615 );
and ( n16617 , n16599 , n16616 );
xor ( n16618 , n16409 , n16413 );
xor ( n16619 , n16618 , n16418 );
and ( n16620 , n16616 , n16619 );
and ( n16621 , n16599 , n16619 );
or ( n16622 , n16617 , n16620 , n16621 );
xor ( n16623 , n16462 , n16466 );
xor ( n16624 , n16623 , n16471 );
xor ( n16625 , n16482 , n16486 );
xor ( n16626 , n16625 , n16491 );
and ( n16627 , n16624 , n16626 );
xor ( n16628 , n16503 , n16507 );
xor ( n16629 , n16628 , n16511 );
and ( n16630 , n16626 , n16629 );
and ( n16631 , n16624 , n16629 );
or ( n16632 , n16627 , n16630 , n16631 );
xor ( n16633 , n16474 , n16494 );
xor ( n16634 , n16633 , n16496 );
and ( n16635 , n16632 , n16634 );
xor ( n16636 , n16514 , n16516 );
xor ( n16637 , n16636 , n16519 );
and ( n16638 , n16634 , n16637 );
and ( n16639 , n16632 , n16637 );
or ( n16640 , n16635 , n16638 , n16639 );
and ( n16641 , n16622 , n16640 );
xor ( n16642 , n16450 , n16452 );
xor ( n16643 , n16642 , n16455 );
and ( n16644 , n16640 , n16643 );
and ( n16645 , n16622 , n16643 );
or ( n16646 , n16641 , n16644 , n16645 );
xor ( n16647 , n16390 , n16427 );
xor ( n16648 , n16647 , n16430 );
and ( n16649 , n16646 , n16648 );
xor ( n16650 , n16458 , n16528 );
xor ( n16651 , n16650 , n16531 );
and ( n16652 , n16648 , n16651 );
and ( n16653 , n16646 , n16651 );
or ( n16654 , n16649 , n16652 , n16653 );
and ( n16655 , n16545 , n16654 );
xor ( n16656 , n16646 , n16648 );
xor ( n16657 , n16656 , n16651 );
and ( n16658 , n16029 , n16018 );
and ( n16659 , n16040 , n16016 );
nor ( n16660 , n16658 , n16659 );
xnor ( n16661 , n16660 , n16026 );
and ( n16662 , n16049 , n16102 );
and ( n16663 , n16058 , n16100 );
nor ( n16664 , n16662 , n16663 );
xnor ( n16665 , n16664 , n16110 );
and ( n16666 , n16661 , n16665 );
buf ( n16667 , n1110 );
buf ( n16668 , n16667 );
and ( n16669 , n16668 , n15984 );
and ( n16670 , n16665 , n16669 );
and ( n16671 , n16661 , n16669 );
or ( n16672 , n16666 , n16670 , n16671 );
and ( n16673 , n15961 , n16084 );
and ( n16674 , n15974 , n16082 );
nor ( n16675 , n16673 , n16674 );
xnor ( n16676 , n16675 , n16092 );
and ( n16677 , n15982 , n15971 );
and ( n16678 , n15995 , n15969 );
nor ( n16679 , n16677 , n16678 );
xnor ( n16680 , n16679 , n15979 );
and ( n16681 , n16676 , n16680 );
and ( n16682 , n16151 , n16037 );
and ( n16683 , n16004 , n16035 );
nor ( n16684 , n16682 , n16683 );
xnor ( n16685 , n16684 , n16045 );
and ( n16686 , n16680 , n16685 );
and ( n16687 , n16676 , n16685 );
or ( n16688 , n16681 , n16686 , n16687 );
and ( n16689 , n16672 , n16688 );
buf ( n16690 , n1175 );
buf ( n16691 , n16690 );
buf ( n16692 , n1176 );
buf ( n16693 , n16692 );
and ( n16694 , n16691 , n16693 );
not ( n16695 , n16694 );
and ( n16696 , n16478 , n16695 );
not ( n16697 , n16696 );
and ( n16698 , n16078 , n16565 );
and ( n16699 , n16087 , n16563 );
nor ( n16700 , n16698 , n16699 );
xnor ( n16701 , n16700 , n16481 );
and ( n16702 , n16697 , n16701 );
and ( n16703 , n16096 , n16176 );
and ( n16704 , n16105 , n16174 );
nor ( n16705 , n16703 , n16704 );
xnor ( n16706 , n16705 , n16075 );
and ( n16707 , n16701 , n16706 );
and ( n16708 , n16697 , n16706 );
or ( n16709 , n16702 , n16707 , n16708 );
and ( n16710 , n16688 , n16709 );
and ( n16711 , n16672 , n16709 );
or ( n16712 , n16689 , n16710 , n16711 );
and ( n16713 , n16008 , n16378 );
and ( n16714 , n16021 , n16376 );
nor ( n16715 , n16713 , n16714 );
xnor ( n16716 , n16715 , n16313 );
and ( n16717 , n16401 , n16055 );
and ( n16718 , n16285 , n16053 );
nor ( n16719 , n16717 , n16718 );
xnor ( n16720 , n16719 , n16063 );
and ( n16721 , n16716 , n16720 );
and ( n16722 , n16592 , n15992 );
and ( n16723 , n16510 , n15990 );
nor ( n16724 , n16722 , n16723 );
xnor ( n16725 , n16724 , n16000 );
and ( n16726 , n16720 , n16725 );
and ( n16727 , n16716 , n16725 );
or ( n16728 , n16721 , n16726 , n16727 );
not ( n16729 , n16603 );
and ( n16730 , n16728 , n16729 );
and ( n16731 , n15995 , n15971 );
and ( n16732 , n16049 , n15969 );
nor ( n16733 , n16731 , n16732 );
xnor ( n16734 , n16733 , n15979 );
and ( n16735 , n16729 , n16734 );
and ( n16736 , n16728 , n16734 );
or ( n16737 , n16730 , n16735 , n16736 );
and ( n16738 , n16712 , n16737 );
xor ( n16739 , n16604 , n16608 );
xor ( n16740 , n16739 , n16613 );
and ( n16741 , n16737 , n16740 );
and ( n16742 , n16712 , n16740 );
or ( n16743 , n16738 , n16741 , n16742 );
xor ( n16744 , n16549 , n16553 );
xor ( n16745 , n16744 , n16558 );
xor ( n16746 , n16568 , n16572 );
xor ( n16747 , n16746 , n16577 );
and ( n16748 , n16745 , n16747 );
xor ( n16749 , n16585 , n16589 );
xor ( n16750 , n16749 , n16593 );
and ( n16751 , n16747 , n16750 );
and ( n16752 , n16745 , n16750 );
or ( n16753 , n16748 , n16751 , n16752 );
xor ( n16754 , n16561 , n16580 );
xor ( n16755 , n16754 , n16596 );
and ( n16756 , n16753 , n16755 );
xor ( n16757 , n16624 , n16626 );
xor ( n16758 , n16757 , n16629 );
and ( n16759 , n16755 , n16758 );
and ( n16760 , n16753 , n16758 );
or ( n16761 , n16756 , n16759 , n16760 );
and ( n16762 , n16743 , n16761 );
xor ( n16763 , n16599 , n16616 );
xor ( n16764 , n16763 , n16619 );
and ( n16765 , n16761 , n16764 );
and ( n16766 , n16743 , n16764 );
or ( n16767 , n16762 , n16765 , n16766 );
xor ( n16768 , n16499 , n16522 );
xor ( n16769 , n16768 , n16525 );
and ( n16770 , n16767 , n16769 );
xor ( n16771 , n16622 , n16640 );
xor ( n16772 , n16771 , n16643 );
and ( n16773 , n16769 , n16772 );
and ( n16774 , n16767 , n16772 );
or ( n16775 , n16770 , n16773 , n16774 );
and ( n16776 , n16657 , n16775 );
xor ( n16777 , n16767 , n16769 );
xor ( n16778 , n16777 , n16772 );
xor ( n16779 , n16478 , n16691 );
xor ( n16780 , n16691 , n16693 );
not ( n16781 , n16780 );
and ( n16782 , n16779 , n16781 );
and ( n16783 , n16087 , n16782 );
not ( n16784 , n16783 );
xnor ( n16785 , n16784 , n16696 );
and ( n16786 , n16105 , n16378 );
and ( n16787 , n16008 , n16376 );
nor ( n16788 , n16786 , n16787 );
xnor ( n16789 , n16788 , n16313 );
and ( n16790 , n16785 , n16789 );
buf ( n16791 , n1111 );
buf ( n16792 , n16791 );
and ( n16793 , n16792 , n15984 );
and ( n16794 , n16789 , n16793 );
and ( n16795 , n16785 , n16793 );
or ( n16796 , n16790 , n16794 , n16795 );
and ( n16797 , n15974 , n16176 );
and ( n16798 , n16096 , n16174 );
nor ( n16799 , n16797 , n16798 );
xnor ( n16800 , n16799 , n16075 );
and ( n16801 , n16004 , n15971 );
and ( n16802 , n15982 , n15969 );
nor ( n16803 , n16801 , n16802 );
xnor ( n16804 , n16803 , n15979 );
and ( n16805 , n16800 , n16804 );
and ( n16806 , n16285 , n16037 );
and ( n16807 , n16151 , n16035 );
nor ( n16808 , n16806 , n16807 );
xnor ( n16809 , n16808 , n16045 );
and ( n16810 , n16804 , n16809 );
and ( n16811 , n16800 , n16809 );
or ( n16812 , n16805 , n16810 , n16811 );
and ( n16813 , n16796 , n16812 );
and ( n16814 , n16021 , n16565 );
and ( n16815 , n16078 , n16563 );
nor ( n16816 , n16814 , n16815 );
xnor ( n16817 , n16816 , n16481 );
buf ( n16818 , n16817 );
and ( n16819 , n16812 , n16818 );
and ( n16820 , n16796 , n16818 );
or ( n16821 , n16813 , n16819 , n16820 );
xor ( n16822 , n16672 , n16688 );
xor ( n16823 , n16822 , n16709 );
and ( n16824 , n16821 , n16823 );
xor ( n16825 , n16728 , n16729 );
xor ( n16826 , n16825 , n16734 );
and ( n16827 , n16823 , n16826 );
and ( n16828 , n16821 , n16826 );
or ( n16829 , n16824 , n16827 , n16828 );
xor ( n16830 , n16712 , n16737 );
xor ( n16831 , n16830 , n16740 );
and ( n16832 , n16829 , n16831 );
xor ( n16833 , n16753 , n16755 );
xor ( n16834 , n16833 , n16758 );
and ( n16835 , n16831 , n16834 );
and ( n16836 , n16829 , n16834 );
or ( n16837 , n16832 , n16835 , n16836 );
xor ( n16838 , n16632 , n16634 );
xor ( n16839 , n16838 , n16637 );
and ( n16840 , n16837 , n16839 );
xor ( n16841 , n16743 , n16761 );
xor ( n16842 , n16841 , n16764 );
and ( n16843 , n16839 , n16842 );
and ( n16844 , n16837 , n16842 );
or ( n16845 , n16840 , n16843 , n16844 );
and ( n16846 , n16778 , n16845 );
xor ( n16847 , n16837 , n16839 );
xor ( n16848 , n16847 , n16842 );
and ( n16849 , n16040 , n16084 );
and ( n16850 , n15961 , n16082 );
nor ( n16851 , n16849 , n16850 );
xnor ( n16852 , n16851 , n16092 );
and ( n16853 , n16510 , n16055 );
and ( n16854 , n16401 , n16053 );
nor ( n16855 , n16853 , n16854 );
xnor ( n16856 , n16855 , n16063 );
and ( n16857 , n16852 , n16856 );
and ( n16858 , n16668 , n15992 );
and ( n16859 , n16592 , n15990 );
nor ( n16860 , n16858 , n16859 );
xnor ( n16861 , n16860 , n16000 );
and ( n16862 , n16856 , n16861 );
and ( n16863 , n16852 , n16861 );
or ( n16864 , n16857 , n16862 , n16863 );
xor ( n16865 , n16661 , n16665 );
xor ( n16866 , n16865 , n16669 );
and ( n16867 , n16864 , n16866 );
xor ( n16868 , n16716 , n16720 );
xor ( n16869 , n16868 , n16725 );
and ( n16870 , n16866 , n16869 );
and ( n16871 , n16864 , n16869 );
or ( n16872 , n16867 , n16870 , n16871 );
not ( n16873 , n16817 );
and ( n16874 , n16058 , n16018 );
and ( n16875 , n16029 , n16016 );
nor ( n16876 , n16874 , n16875 );
xnor ( n16877 , n16876 , n16026 );
and ( n16878 , n16873 , n16877 );
and ( n16879 , n15995 , n16102 );
and ( n16880 , n16049 , n16100 );
nor ( n16881 , n16879 , n16880 );
xnor ( n16882 , n16881 , n16110 );
and ( n16883 , n16877 , n16882 );
and ( n16884 , n16873 , n16882 );
or ( n16885 , n16878 , n16883 , n16884 );
xor ( n16886 , n16676 , n16680 );
xor ( n16887 , n16886 , n16685 );
and ( n16888 , n16885 , n16887 );
xor ( n16889 , n16697 , n16701 );
xor ( n16890 , n16889 , n16706 );
and ( n16891 , n16887 , n16890 );
and ( n16892 , n16885 , n16890 );
or ( n16893 , n16888 , n16891 , n16892 );
and ( n16894 , n16872 , n16893 );
xor ( n16895 , n16745 , n16747 );
xor ( n16896 , n16895 , n16750 );
and ( n16897 , n16893 , n16896 );
and ( n16898 , n16872 , n16896 );
or ( n16899 , n16894 , n16897 , n16898 );
and ( n16900 , n16029 , n16084 );
and ( n16901 , n16040 , n16082 );
nor ( n16902 , n16900 , n16901 );
xnor ( n16903 , n16902 , n16092 );
and ( n16904 , n16792 , n15992 );
and ( n16905 , n16668 , n15990 );
nor ( n16906 , n16904 , n16905 );
xnor ( n16907 , n16906 , n16000 );
and ( n16908 , n16903 , n16907 );
buf ( n16909 , n1112 );
buf ( n16910 , n16909 );
and ( n16911 , n16910 , n15984 );
and ( n16912 , n16907 , n16911 );
and ( n16913 , n16903 , n16911 );
or ( n16914 , n16908 , n16912 , n16913 );
and ( n16915 , n16008 , n16565 );
and ( n16916 , n16021 , n16563 );
nor ( n16917 , n16915 , n16916 );
xnor ( n16918 , n16917 , n16481 );
and ( n16919 , n16401 , n16037 );
and ( n16920 , n16285 , n16035 );
nor ( n16921 , n16919 , n16920 );
xnor ( n16922 , n16921 , n16045 );
and ( n16923 , n16918 , n16922 );
and ( n16924 , n16592 , n16055 );
and ( n16925 , n16510 , n16053 );
nor ( n16926 , n16924 , n16925 );
xnor ( n16927 , n16926 , n16063 );
and ( n16928 , n16922 , n16927 );
and ( n16929 , n16918 , n16927 );
or ( n16930 , n16923 , n16928 , n16929 );
and ( n16931 , n16914 , n16930 );
buf ( n16932 , n1177 );
buf ( n16933 , n16932 );
buf ( n16934 , n1178 );
buf ( n16935 , n16934 );
and ( n16936 , n16933 , n16935 );
not ( n16937 , n16936 );
and ( n16938 , n16693 , n16937 );
not ( n16939 , n16938 );
and ( n16940 , n16078 , n16782 );
and ( n16941 , n16087 , n16780 );
nor ( n16942 , n16940 , n16941 );
xnor ( n16943 , n16942 , n16696 );
and ( n16944 , n16939 , n16943 );
and ( n16945 , n16096 , n16378 );
and ( n16946 , n16105 , n16376 );
nor ( n16947 , n16945 , n16946 );
xnor ( n16948 , n16947 , n16313 );
and ( n16949 , n16943 , n16948 );
and ( n16950 , n16939 , n16948 );
or ( n16951 , n16944 , n16949 , n16950 );
and ( n16952 , n16930 , n16951 );
and ( n16953 , n16914 , n16951 );
or ( n16954 , n16931 , n16952 , n16953 );
and ( n16955 , n15961 , n16176 );
and ( n16956 , n15974 , n16174 );
nor ( n16957 , n16955 , n16956 );
xnor ( n16958 , n16957 , n16075 );
and ( n16959 , n15982 , n16102 );
and ( n16960 , n15995 , n16100 );
nor ( n16961 , n16959 , n16960 );
xnor ( n16962 , n16961 , n16110 );
and ( n16963 , n16958 , n16962 );
and ( n16964 , n16151 , n15971 );
and ( n16965 , n16004 , n15969 );
nor ( n16966 , n16964 , n16965 );
xnor ( n16967 , n16966 , n15979 );
and ( n16968 , n16962 , n16967 );
and ( n16969 , n16958 , n16967 );
or ( n16970 , n16963 , n16968 , n16969 );
xor ( n16971 , n16785 , n16789 );
xor ( n16972 , n16971 , n16793 );
and ( n16973 , n16970 , n16972 );
xor ( n16974 , n16800 , n16804 );
xor ( n16975 , n16974 , n16809 );
and ( n16976 , n16972 , n16975 );
and ( n16977 , n16970 , n16975 );
or ( n16978 , n16973 , n16976 , n16977 );
and ( n16979 , n16954 , n16978 );
xor ( n16980 , n16796 , n16812 );
xor ( n16981 , n16980 , n16818 );
and ( n16982 , n16978 , n16981 );
and ( n16983 , n16954 , n16981 );
or ( n16984 , n16979 , n16982 , n16983 );
and ( n16985 , n16105 , n16565 );
and ( n16986 , n16008 , n16563 );
nor ( n16987 , n16985 , n16986 );
xnor ( n16988 , n16987 , n16481 );
and ( n16989 , n15995 , n16018 );
and ( n16990 , n16049 , n16016 );
nor ( n16991 , n16989 , n16990 );
xnor ( n16992 , n16991 , n16026 );
and ( n16993 , n16988 , n16992 );
buf ( n16994 , n1113 );
buf ( n16995 , n16994 );
and ( n16996 , n16995 , n15984 );
and ( n16997 , n16992 , n16996 );
and ( n16998 , n16988 , n16996 );
or ( n16999 , n16993 , n16997 , n16998 );
and ( n17000 , n15974 , n16378 );
and ( n17001 , n16096 , n16376 );
nor ( n17002 , n17000 , n17001 );
xnor ( n17003 , n17002 , n16313 );
and ( n17004 , n16004 , n16102 );
and ( n17005 , n15982 , n16100 );
nor ( n17006 , n17004 , n17005 );
xnor ( n17007 , n17006 , n16110 );
and ( n17008 , n17003 , n17007 );
and ( n17009 , n16285 , n15971 );
and ( n17010 , n16151 , n15969 );
nor ( n17011 , n17009 , n17010 );
xnor ( n17012 , n17011 , n15979 );
and ( n17013 , n17007 , n17012 );
and ( n17014 , n17003 , n17012 );
or ( n17015 , n17008 , n17013 , n17014 );
and ( n17016 , n16999 , n17015 );
xor ( n17017 , n16693 , n16933 );
xor ( n17018 , n16933 , n16935 );
not ( n17019 , n17018 );
and ( n17020 , n17017 , n17019 );
and ( n17021 , n16087 , n17020 );
not ( n17022 , n17021 );
xnor ( n17023 , n17022 , n16938 );
and ( n17024 , n16058 , n16084 );
and ( n17025 , n16029 , n16082 );
nor ( n17026 , n17024 , n17025 );
xnor ( n17027 , n17026 , n16092 );
and ( n17028 , n17023 , n17027 );
and ( n17029 , n16910 , n15992 );
and ( n17030 , n16792 , n15990 );
nor ( n17031 , n17029 , n17030 );
xnor ( n17032 , n17031 , n16000 );
and ( n17033 , n17027 , n17032 );
and ( n17034 , n17023 , n17032 );
or ( n17035 , n17028 , n17033 , n17034 );
and ( n17036 , n17015 , n17035 );
and ( n17037 , n16999 , n17035 );
or ( n17038 , n17016 , n17036 , n17037 );
xor ( n17039 , n16852 , n16856 );
xor ( n17040 , n17039 , n16861 );
and ( n17041 , n17038 , n17040 );
xor ( n17042 , n16873 , n16877 );
xor ( n17043 , n17042 , n16882 );
and ( n17044 , n17040 , n17043 );
and ( n17045 , n17038 , n17043 );
or ( n17046 , n17041 , n17044 , n17045 );
xor ( n17047 , n16864 , n16866 );
xor ( n17048 , n17047 , n16869 );
and ( n17049 , n17046 , n17048 );
xor ( n17050 , n16885 , n16887 );
xor ( n17051 , n17050 , n16890 );
and ( n17052 , n17048 , n17051 );
and ( n17053 , n17046 , n17051 );
or ( n17054 , n17049 , n17052 , n17053 );
and ( n17055 , n16984 , n17054 );
xor ( n17056 , n16821 , n16823 );
xor ( n17057 , n17056 , n16826 );
and ( n17058 , n17054 , n17057 );
and ( n17059 , n16984 , n17057 );
or ( n17060 , n17055 , n17058 , n17059 );
and ( n17061 , n16899 , n17060 );
xor ( n17062 , n16829 , n16831 );
xor ( n17063 , n17062 , n16834 );
and ( n17064 , n17060 , n17063 );
and ( n17065 , n16899 , n17063 );
or ( n17066 , n17061 , n17064 , n17065 );
and ( n17067 , n16848 , n17066 );
xor ( n17068 , n16899 , n17060 );
xor ( n17069 , n17068 , n17063 );
and ( n17070 , n16040 , n16176 );
and ( n17071 , n15961 , n16174 );
nor ( n17072 , n17070 , n17071 );
xnor ( n17073 , n17072 , n16075 );
and ( n17074 , n16510 , n16037 );
and ( n17075 , n16401 , n16035 );
nor ( n17076 , n17074 , n17075 );
xnor ( n17077 , n17076 , n16045 );
and ( n17078 , n17073 , n17077 );
and ( n17079 , n16668 , n16055 );
and ( n17080 , n16592 , n16053 );
nor ( n17081 , n17079 , n17080 );
xnor ( n17082 , n17081 , n16063 );
and ( n17083 , n17077 , n17082 );
and ( n17084 , n17073 , n17082 );
or ( n17085 , n17078 , n17083 , n17084 );
and ( n17086 , n16021 , n16782 );
and ( n17087 , n16078 , n16780 );
nor ( n17088 , n17086 , n17087 );
xnor ( n17089 , n17088 , n16696 );
buf ( n17090 , n17089 );
and ( n17091 , n17085 , n17090 );
and ( n17092 , n16049 , n16018 );
and ( n17093 , n16058 , n16016 );
nor ( n17094 , n17092 , n17093 );
xnor ( n17095 , n17094 , n16026 );
and ( n17096 , n17090 , n17095 );
and ( n17097 , n17085 , n17095 );
or ( n17098 , n17091 , n17096 , n17097 );
xor ( n17099 , n16958 , n16962 );
xor ( n17100 , n17099 , n16967 );
xor ( n17101 , n16918 , n16922 );
xor ( n17102 , n17101 , n16927 );
and ( n17103 , n17100 , n17102 );
xor ( n17104 , n16939 , n16943 );
xor ( n17105 , n17104 , n16948 );
and ( n17106 , n17102 , n17105 );
and ( n17107 , n17100 , n17105 );
or ( n17108 , n17103 , n17106 , n17107 );
and ( n17109 , n17098 , n17108 );
xor ( n17110 , n16914 , n16930 );
xor ( n17111 , n17110 , n16951 );
and ( n17112 , n17108 , n17111 );
and ( n17113 , n17098 , n17111 );
or ( n17114 , n17109 , n17112 , n17113 );
and ( n17115 , n15961 , n16378 );
and ( n17116 , n15974 , n16376 );
nor ( n17117 , n17115 , n17116 );
xnor ( n17118 , n17117 , n16313 );
and ( n17119 , n15982 , n16018 );
and ( n17120 , n15995 , n16016 );
nor ( n17121 , n17119 , n17120 );
xnor ( n17122 , n17121 , n16026 );
and ( n17123 , n17118 , n17122 );
and ( n17124 , n16151 , n16102 );
and ( n17125 , n16004 , n16100 );
nor ( n17126 , n17124 , n17125 );
xnor ( n17127 , n17126 , n16110 );
and ( n17128 , n17122 , n17127 );
and ( n17129 , n17118 , n17127 );
or ( n17130 , n17123 , n17128 , n17129 );
and ( n17131 , n16008 , n16782 );
and ( n17132 , n16021 , n16780 );
nor ( n17133 , n17131 , n17132 );
xnor ( n17134 , n17133 , n16696 );
and ( n17135 , n16401 , n15971 );
and ( n17136 , n16285 , n15969 );
nor ( n17137 , n17135 , n17136 );
xnor ( n17138 , n17137 , n15979 );
and ( n17139 , n17134 , n17138 );
and ( n17140 , n16592 , n16037 );
and ( n17141 , n16510 , n16035 );
nor ( n17142 , n17140 , n17141 );
xnor ( n17143 , n17142 , n16045 );
and ( n17144 , n17138 , n17143 );
and ( n17145 , n17134 , n17143 );
or ( n17146 , n17139 , n17144 , n17145 );
and ( n17147 , n17130 , n17146 );
not ( n17148 , n17089 );
and ( n17149 , n17146 , n17148 );
and ( n17150 , n17130 , n17148 );
or ( n17151 , n17147 , n17149 , n17150 );
xor ( n17152 , n16903 , n16907 );
xor ( n17153 , n17152 , n16911 );
and ( n17154 , n17151 , n17153 );
xor ( n17155 , n17085 , n17090 );
xor ( n17156 , n17155 , n17095 );
and ( n17157 , n17153 , n17156 );
and ( n17158 , n17151 , n17156 );
or ( n17159 , n17154 , n17157 , n17158 );
xor ( n17160 , n16970 , n16972 );
xor ( n17161 , n17160 , n16975 );
and ( n17162 , n17159 , n17161 );
xor ( n17163 , n17038 , n17040 );
xor ( n17164 , n17163 , n17043 );
and ( n17165 , n17161 , n17164 );
and ( n17166 , n17159 , n17164 );
or ( n17167 , n17162 , n17165 , n17166 );
and ( n17168 , n17114 , n17167 );
xor ( n17169 , n16954 , n16978 );
xor ( n17170 , n17169 , n16981 );
and ( n17171 , n17167 , n17170 );
and ( n17172 , n17114 , n17170 );
or ( n17173 , n17168 , n17171 , n17172 );
xor ( n17174 , n16872 , n16893 );
xor ( n17175 , n17174 , n16896 );
and ( n17176 , n17173 , n17175 );
xor ( n17177 , n16984 , n17054 );
xor ( n17178 , n17177 , n17057 );
and ( n17179 , n17175 , n17178 );
and ( n17180 , n17173 , n17178 );
or ( n17181 , n17176 , n17179 , n17180 );
and ( n17182 , n17069 , n17181 );
xor ( n17183 , n17173 , n17175 );
xor ( n17184 , n17183 , n17178 );
buf ( n17185 , n1179 );
buf ( n17186 , n17185 );
buf ( n17187 , n1180 );
buf ( n17188 , n17187 );
and ( n17189 , n17186 , n17188 );
not ( n17190 , n17189 );
and ( n17191 , n16935 , n17190 );
not ( n17192 , n17191 );
and ( n17193 , n16078 , n17020 );
and ( n17194 , n16087 , n17018 );
nor ( n17195 , n17193 , n17194 );
xnor ( n17196 , n17195 , n16938 );
and ( n17197 , n17192 , n17196 );
and ( n17198 , n16096 , n16565 );
and ( n17199 , n16105 , n16563 );
nor ( n17200 , n17198 , n17199 );
xnor ( n17201 , n17200 , n16481 );
and ( n17202 , n17196 , n17201 );
and ( n17203 , n17192 , n17201 );
or ( n17204 , n17197 , n17202 , n17203 );
and ( n17205 , n16029 , n16176 );
and ( n17206 , n16040 , n16174 );
nor ( n17207 , n17205 , n17206 );
xnor ( n17208 , n17207 , n16075 );
and ( n17209 , n16792 , n16055 );
and ( n17210 , n16668 , n16053 );
nor ( n17211 , n17209 , n17210 );
xnor ( n17212 , n17211 , n16063 );
and ( n17213 , n17208 , n17212 );
and ( n17214 , n16995 , n15992 );
and ( n17215 , n16910 , n15990 );
nor ( n17216 , n17214 , n17215 );
xnor ( n17217 , n17216 , n16000 );
and ( n17218 , n17212 , n17217 );
and ( n17219 , n17208 , n17217 );
or ( n17220 , n17213 , n17218 , n17219 );
and ( n17221 , n17204 , n17220 );
xor ( n17222 , n16988 , n16992 );
xor ( n17223 , n17222 , n16996 );
and ( n17224 , n17220 , n17223 );
and ( n17225 , n17204 , n17223 );
or ( n17226 , n17221 , n17224 , n17225 );
xor ( n17227 , n17003 , n17007 );
xor ( n17228 , n17227 , n17012 );
xor ( n17229 , n17023 , n17027 );
xor ( n17230 , n17229 , n17032 );
and ( n17231 , n17228 , n17230 );
xor ( n17232 , n17073 , n17077 );
xor ( n17233 , n17232 , n17082 );
and ( n17234 , n17230 , n17233 );
and ( n17235 , n17228 , n17233 );
or ( n17236 , n17231 , n17234 , n17235 );
and ( n17237 , n17226 , n17236 );
xor ( n17238 , n16999 , n17015 );
xor ( n17239 , n17238 , n17035 );
and ( n17240 , n17236 , n17239 );
and ( n17241 , n17226 , n17239 );
or ( n17242 , n17237 , n17240 , n17241 );
xor ( n17243 , n16935 , n17186 );
xor ( n17244 , n17186 , n17188 );
not ( n17245 , n17244 );
and ( n17246 , n17243 , n17245 );
and ( n17247 , n16087 , n17246 );
not ( n17248 , n17247 );
xnor ( n17249 , n17248 , n17191 );
and ( n17250 , n16058 , n16176 );
and ( n17251 , n16029 , n16174 );
nor ( n17252 , n17250 , n17251 );
xnor ( n17253 , n17252 , n16075 );
and ( n17254 , n17249 , n17253 );
and ( n17255 , n16910 , n16055 );
and ( n17256 , n16792 , n16053 );
nor ( n17257 , n17255 , n17256 );
xnor ( n17258 , n17257 , n16063 );
and ( n17259 , n17253 , n17258 );
and ( n17260 , n17249 , n17258 );
or ( n17261 , n17254 , n17259 , n17260 );
and ( n17262 , n16040 , n16378 );
and ( n17263 , n15961 , n16376 );
nor ( n17264 , n17262 , n17263 );
xnor ( n17265 , n17264 , n16313 );
and ( n17266 , n16510 , n15971 );
and ( n17267 , n16401 , n15969 );
nor ( n17268 , n17266 , n17267 );
xnor ( n17269 , n17268 , n15979 );
and ( n17270 , n17265 , n17269 );
and ( n17271 , n16668 , n16037 );
and ( n17272 , n16592 , n16035 );
nor ( n17273 , n17271 , n17272 );
xnor ( n17274 , n17273 , n16045 );
and ( n17275 , n17269 , n17274 );
and ( n17276 , n17265 , n17274 );
or ( n17277 , n17270 , n17275 , n17276 );
and ( n17278 , n17261 , n17277 );
and ( n17279 , n15974 , n16565 );
and ( n17280 , n16096 , n16563 );
nor ( n17281 , n17279 , n17280 );
xnor ( n17282 , n17281 , n16481 );
and ( n17283 , n16004 , n16018 );
and ( n17284 , n15982 , n16016 );
nor ( n17285 , n17283 , n17284 );
xnor ( n17286 , n17285 , n16026 );
and ( n17287 , n17282 , n17286 );
and ( n17288 , n16285 , n16102 );
and ( n17289 , n16151 , n16100 );
nor ( n17290 , n17288 , n17289 );
xnor ( n17291 , n17290 , n16110 );
and ( n17292 , n17286 , n17291 );
and ( n17293 , n17282 , n17291 );
or ( n17294 , n17287 , n17292 , n17293 );
and ( n17295 , n17277 , n17294 );
and ( n17296 , n17261 , n17294 );
or ( n17297 , n17278 , n17295 , n17296 );
and ( n17298 , n16021 , n17020 );
and ( n17299 , n16078 , n17018 );
nor ( n17300 , n17298 , n17299 );
xnor ( n17301 , n17300 , n16938 );
buf ( n17302 , n17301 );
and ( n17303 , n16049 , n16084 );
and ( n17304 , n16058 , n16082 );
nor ( n17305 , n17303 , n17304 );
xnor ( n17306 , n17305 , n16092 );
and ( n17307 , n17302 , n17306 );
buf ( n17308 , n1114 );
buf ( n17309 , n17308 );
and ( n17310 , n17309 , n15984 );
and ( n17311 , n17306 , n17310 );
and ( n17312 , n17302 , n17310 );
or ( n17313 , n17307 , n17311 , n17312 );
and ( n17314 , n17297 , n17313 );
xor ( n17315 , n17130 , n17146 );
xor ( n17316 , n17315 , n17148 );
and ( n17317 , n17313 , n17316 );
and ( n17318 , n17297 , n17316 );
or ( n17319 , n17314 , n17317 , n17318 );
xor ( n17320 , n17100 , n17102 );
xor ( n17321 , n17320 , n17105 );
and ( n17322 , n17319 , n17321 );
xor ( n17323 , n17151 , n17153 );
xor ( n17324 , n17323 , n17156 );
and ( n17325 , n17321 , n17324 );
and ( n17326 , n17319 , n17324 );
or ( n17327 , n17322 , n17325 , n17326 );
and ( n17328 , n17242 , n17327 );
xor ( n17329 , n17098 , n17108 );
xor ( n17330 , n17329 , n17111 );
and ( n17331 , n17327 , n17330 );
and ( n17332 , n17242 , n17330 );
or ( n17333 , n17328 , n17331 , n17332 );
xor ( n17334 , n17046 , n17048 );
xor ( n17335 , n17334 , n17051 );
and ( n17336 , n17333 , n17335 );
xor ( n17337 , n17114 , n17167 );
xor ( n17338 , n17337 , n17170 );
and ( n17339 , n17335 , n17338 );
and ( n17340 , n17333 , n17338 );
or ( n17341 , n17336 , n17339 , n17340 );
and ( n17342 , n17184 , n17341 );
xor ( n17343 , n17333 , n17335 );
xor ( n17344 , n17343 , n17338 );
and ( n17345 , n16105 , n16782 );
and ( n17346 , n16008 , n16780 );
nor ( n17347 , n17345 , n17346 );
xnor ( n17348 , n17347 , n16696 );
and ( n17349 , n17309 , n15992 );
and ( n17350 , n16995 , n15990 );
nor ( n17351 , n17349 , n17350 );
xnor ( n17352 , n17351 , n16000 );
and ( n17353 , n17348 , n17352 );
buf ( n17354 , n1115 );
buf ( n17355 , n17354 );
and ( n17356 , n17355 , n15984 );
and ( n17357 , n17352 , n17356 );
and ( n17358 , n17348 , n17356 );
or ( n17359 , n17353 , n17357 , n17358 );
xor ( n17360 , n17118 , n17122 );
xor ( n17361 , n17360 , n17127 );
and ( n17362 , n17359 , n17361 );
xor ( n17363 , n17192 , n17196 );
xor ( n17364 , n17363 , n17201 );
and ( n17365 , n17361 , n17364 );
and ( n17366 , n17359 , n17364 );
or ( n17367 , n17362 , n17365 , n17366 );
xor ( n17368 , n17134 , n17138 );
xor ( n17369 , n17368 , n17143 );
xor ( n17370 , n17208 , n17212 );
xor ( n17371 , n17370 , n17217 );
and ( n17372 , n17369 , n17371 );
xor ( n17373 , n17302 , n17306 );
xor ( n17374 , n17373 , n17310 );
and ( n17375 , n17371 , n17374 );
and ( n17376 , n17369 , n17374 );
or ( n17377 , n17372 , n17375 , n17376 );
and ( n17378 , n17367 , n17377 );
xor ( n17379 , n17204 , n17220 );
xor ( n17380 , n17379 , n17223 );
and ( n17381 , n17377 , n17380 );
and ( n17382 , n17367 , n17380 );
or ( n17383 , n17378 , n17381 , n17382 );
and ( n17384 , n15961 , n16565 );
and ( n17385 , n15974 , n16563 );
nor ( n17386 , n17384 , n17385 );
xnor ( n17387 , n17386 , n16481 );
and ( n17388 , n15982 , n16084 );
and ( n17389 , n15995 , n16082 );
nor ( n17390 , n17388 , n17389 );
xnor ( n17391 , n17390 , n16092 );
and ( n17392 , n17387 , n17391 );
and ( n17393 , n16151 , n16018 );
and ( n17394 , n16004 , n16016 );
nor ( n17395 , n17393 , n17394 );
xnor ( n17396 , n17395 , n16026 );
and ( n17397 , n17391 , n17396 );
and ( n17398 , n17387 , n17396 );
or ( n17399 , n17392 , n17397 , n17398 );
buf ( n17400 , n1181 );
buf ( n17401 , n17400 );
buf ( n17402 , n1182 );
buf ( n17403 , n17402 );
and ( n17404 , n17401 , n17403 );
not ( n17405 , n17404 );
and ( n17406 , n17188 , n17405 );
not ( n17407 , n17406 );
and ( n17408 , n16078 , n17246 );
and ( n17409 , n16087 , n17244 );
nor ( n17410 , n17408 , n17409 );
xnor ( n17411 , n17410 , n17191 );
and ( n17412 , n17407 , n17411 );
and ( n17413 , n16096 , n16782 );
and ( n17414 , n16105 , n16780 );
nor ( n17415 , n17413 , n17414 );
xnor ( n17416 , n17415 , n16696 );
and ( n17417 , n17411 , n17416 );
and ( n17418 , n17407 , n17416 );
or ( n17419 , n17412 , n17417 , n17418 );
and ( n17420 , n17399 , n17419 );
and ( n17421 , n16008 , n17020 );
and ( n17422 , n16021 , n17018 );
nor ( n17423 , n17421 , n17422 );
xnor ( n17424 , n17423 , n16938 );
and ( n17425 , n16401 , n16102 );
and ( n17426 , n16285 , n16100 );
nor ( n17427 , n17425 , n17426 );
xnor ( n17428 , n17427 , n16110 );
and ( n17429 , n17424 , n17428 );
and ( n17430 , n16592 , n15971 );
and ( n17431 , n16510 , n15969 );
nor ( n17432 , n17430 , n17431 );
xnor ( n17433 , n17432 , n15979 );
and ( n17434 , n17428 , n17433 );
and ( n17435 , n17424 , n17433 );
or ( n17436 , n17429 , n17434 , n17435 );
and ( n17437 , n17419 , n17436 );
and ( n17438 , n17399 , n17436 );
or ( n17439 , n17420 , n17437 , n17438 );
and ( n17440 , n16029 , n16378 );
and ( n17441 , n16040 , n16376 );
nor ( n17442 , n17440 , n17441 );
xnor ( n17443 , n17442 , n16313 );
and ( n17444 , n16792 , n16037 );
and ( n17445 , n16668 , n16035 );
nor ( n17446 , n17444 , n17445 );
xnor ( n17447 , n17446 , n16045 );
and ( n17448 , n17443 , n17447 );
and ( n17449 , n16995 , n16055 );
and ( n17450 , n16910 , n16053 );
nor ( n17451 , n17449 , n17450 );
xnor ( n17452 , n17451 , n16063 );
and ( n17453 , n17447 , n17452 );
and ( n17454 , n17443 , n17452 );
or ( n17455 , n17448 , n17453 , n17454 );
not ( n17456 , n17301 );
and ( n17457 , n17455 , n17456 );
and ( n17458 , n15995 , n16084 );
and ( n17459 , n16049 , n16082 );
nor ( n17460 , n17458 , n17459 );
xnor ( n17461 , n17460 , n16092 );
and ( n17462 , n17456 , n17461 );
and ( n17463 , n17455 , n17461 );
or ( n17464 , n17457 , n17462 , n17463 );
and ( n17465 , n17439 , n17464 );
xor ( n17466 , n17261 , n17277 );
xor ( n17467 , n17466 , n17294 );
and ( n17468 , n17464 , n17467 );
and ( n17469 , n17439 , n17467 );
or ( n17470 , n17465 , n17468 , n17469 );
xor ( n17471 , n17228 , n17230 );
xor ( n17472 , n17471 , n17233 );
and ( n17473 , n17470 , n17472 );
xor ( n17474 , n17297 , n17313 );
xor ( n17475 , n17474 , n17316 );
and ( n17476 , n17472 , n17475 );
and ( n17477 , n17470 , n17475 );
or ( n17478 , n17473 , n17476 , n17477 );
and ( n17479 , n17383 , n17478 );
xor ( n17480 , n17226 , n17236 );
xor ( n17481 , n17480 , n17239 );
and ( n17482 , n17478 , n17481 );
and ( n17483 , n17383 , n17481 );
or ( n17484 , n17479 , n17482 , n17483 );
xor ( n17485 , n17159 , n17161 );
xor ( n17486 , n17485 , n17164 );
and ( n17487 , n17484 , n17486 );
xor ( n17488 , n17242 , n17327 );
xor ( n17489 , n17488 , n17330 );
and ( n17490 , n17486 , n17489 );
and ( n17491 , n17484 , n17489 );
or ( n17492 , n17487 , n17490 , n17491 );
and ( n17493 , n17344 , n17492 );
xor ( n17494 , n17484 , n17486 );
xor ( n17495 , n17494 , n17489 );
xor ( n17496 , n17249 , n17253 );
xor ( n17497 , n17496 , n17258 );
xor ( n17498 , n17265 , n17269 );
xor ( n17499 , n17498 , n17274 );
and ( n17500 , n17497 , n17499 );
xor ( n17501 , n17455 , n17456 );
xor ( n17502 , n17501 , n17461 );
and ( n17503 , n17499 , n17502 );
and ( n17504 , n17497 , n17502 );
or ( n17505 , n17500 , n17503 , n17504 );
and ( n17506 , n16021 , n17246 );
and ( n17507 , n16078 , n17244 );
nor ( n17508 , n17506 , n17507 );
xnor ( n17509 , n17508 , n17191 );
and ( n17510 , n15974 , n16782 );
and ( n17511 , n16096 , n16780 );
nor ( n17512 , n17510 , n17511 );
xnor ( n17513 , n17512 , n16696 );
and ( n17514 , n17509 , n17513 );
and ( n17515 , n16004 , n16084 );
and ( n17516 , n15982 , n16082 );
nor ( n17517 , n17515 , n17516 );
xnor ( n17518 , n17517 , n16092 );
and ( n17519 , n17513 , n17518 );
and ( n17520 , n17509 , n17518 );
or ( n17521 , n17514 , n17519 , n17520 );
and ( n17522 , n16040 , n16565 );
and ( n17523 , n15961 , n16563 );
nor ( n17524 , n17522 , n17523 );
xnor ( n17525 , n17524 , n16481 );
and ( n17526 , n16285 , n16018 );
and ( n17527 , n16151 , n16016 );
nor ( n17528 , n17526 , n17527 );
xnor ( n17529 , n17528 , n16026 );
and ( n17530 , n17525 , n17529 );
and ( n17531 , n16510 , n16102 );
and ( n17532 , n16401 , n16100 );
nor ( n17533 , n17531 , n17532 );
xnor ( n17534 , n17533 , n16110 );
and ( n17535 , n17529 , n17534 );
and ( n17536 , n17525 , n17534 );
or ( n17537 , n17530 , n17535 , n17536 );
and ( n17538 , n17521 , n17537 );
xor ( n17539 , n17188 , n17401 );
xor ( n17540 , n17401 , n17403 );
not ( n17541 , n17540 );
and ( n17542 , n17539 , n17541 );
and ( n17543 , n16087 , n17542 );
not ( n17544 , n17543 );
xnor ( n17545 , n17544 , n17406 );
buf ( n17546 , n17545 );
and ( n17547 , n17537 , n17546 );
and ( n17548 , n17521 , n17546 );
or ( n17549 , n17538 , n17547 , n17548 );
and ( n17550 , n15995 , n16176 );
and ( n17551 , n16049 , n16174 );
nor ( n17552 , n17550 , n17551 );
xnor ( n17553 , n17552 , n16075 );
and ( n17554 , n16910 , n16037 );
and ( n17555 , n16792 , n16035 );
nor ( n17556 , n17554 , n17555 );
xnor ( n17557 , n17556 , n16045 );
and ( n17558 , n17553 , n17557 );
and ( n17559 , n17309 , n16055 );
and ( n17560 , n16995 , n16053 );
nor ( n17561 , n17559 , n17560 );
xnor ( n17562 , n17561 , n16063 );
and ( n17563 , n17557 , n17562 );
and ( n17564 , n17553 , n17562 );
or ( n17565 , n17558 , n17563 , n17564 );
and ( n17566 , n16105 , n17020 );
and ( n17567 , n16008 , n17018 );
nor ( n17568 , n17566 , n17567 );
xnor ( n17569 , n17568 , n16938 );
and ( n17570 , n16058 , n16378 );
and ( n17571 , n16029 , n16376 );
nor ( n17572 , n17570 , n17571 );
xnor ( n17573 , n17572 , n16313 );
and ( n17574 , n17569 , n17573 );
and ( n17575 , n16668 , n15971 );
and ( n17576 , n16592 , n15969 );
nor ( n17577 , n17575 , n17576 );
xnor ( n17578 , n17577 , n15979 );
and ( n17579 , n17573 , n17578 );
and ( n17580 , n17569 , n17578 );
or ( n17581 , n17574 , n17579 , n17580 );
and ( n17582 , n17565 , n17581 );
xor ( n17583 , n17387 , n17391 );
xor ( n17584 , n17583 , n17396 );
and ( n17585 , n17581 , n17584 );
and ( n17586 , n17565 , n17584 );
or ( n17587 , n17582 , n17585 , n17586 );
and ( n17588 , n17549 , n17587 );
xor ( n17589 , n17399 , n17419 );
xor ( n17590 , n17589 , n17436 );
and ( n17591 , n17587 , n17590 );
and ( n17592 , n17549 , n17590 );
or ( n17593 , n17588 , n17591 , n17592 );
and ( n17594 , n17505 , n17593 );
xor ( n17595 , n17439 , n17464 );
xor ( n17596 , n17595 , n17467 );
and ( n17597 , n17593 , n17596 );
and ( n17598 , n17505 , n17596 );
or ( n17599 , n17594 , n17597 , n17598 );
and ( n17600 , n16049 , n16176 );
and ( n17601 , n16058 , n16174 );
nor ( n17602 , n17600 , n17601 );
xnor ( n17603 , n17602 , n16075 );
and ( n17604 , n17355 , n15992 );
and ( n17605 , n17309 , n15990 );
nor ( n17606 , n17604 , n17605 );
xnor ( n17607 , n17606 , n16000 );
and ( n17608 , n17603 , n17607 );
buf ( n17609 , n1116 );
buf ( n17610 , n17609 );
and ( n17611 , n17610 , n15984 );
and ( n17612 , n17607 , n17611 );
and ( n17613 , n17603 , n17611 );
or ( n17614 , n17608 , n17612 , n17613 );
xor ( n17615 , n17348 , n17352 );
xor ( n17616 , n17615 , n17356 );
and ( n17617 , n17614 , n17616 );
xor ( n17618 , n17282 , n17286 );
xor ( n17619 , n17618 , n17291 );
and ( n17620 , n17616 , n17619 );
and ( n17621 , n17614 , n17619 );
or ( n17622 , n17617 , n17620 , n17621 );
xor ( n17623 , n17359 , n17361 );
xor ( n17624 , n17623 , n17364 );
and ( n17625 , n17622 , n17624 );
xor ( n17626 , n17369 , n17371 );
xor ( n17627 , n17626 , n17374 );
and ( n17628 , n17624 , n17627 );
and ( n17629 , n17622 , n17627 );
or ( n17630 , n17625 , n17628 , n17629 );
and ( n17631 , n17599 , n17630 );
xor ( n17632 , n17367 , n17377 );
xor ( n17633 , n17632 , n17380 );
and ( n17634 , n17630 , n17633 );
and ( n17635 , n17599 , n17633 );
or ( n17636 , n17631 , n17634 , n17635 );
xor ( n17637 , n17319 , n17321 );
xor ( n17638 , n17637 , n17324 );
and ( n17639 , n17636 , n17638 );
xor ( n17640 , n17383 , n17478 );
xor ( n17641 , n17640 , n17481 );
and ( n17642 , n17638 , n17641 );
and ( n17643 , n17636 , n17641 );
or ( n17644 , n17639 , n17642 , n17643 );
and ( n17645 , n17495 , n17644 );
xor ( n17646 , n17636 , n17638 );
xor ( n17647 , n17646 , n17641 );
xor ( n17648 , n17603 , n17607 );
xor ( n17649 , n17648 , n17611 );
xor ( n17650 , n17407 , n17411 );
xor ( n17651 , n17650 , n17416 );
and ( n17652 , n17649 , n17651 );
xor ( n17653 , n17443 , n17447 );
xor ( n17654 , n17653 , n17452 );
and ( n17655 , n17651 , n17654 );
and ( n17656 , n17649 , n17654 );
or ( n17657 , n17652 , n17655 , n17656 );
buf ( n17658 , n1183 );
buf ( n17659 , n17658 );
buf ( n17660 , n1184 );
buf ( n17661 , n17660 );
and ( n17662 , n17659 , n17661 );
not ( n17663 , n17662 );
and ( n17664 , n17403 , n17663 );
not ( n17665 , n17664 );
and ( n17666 , n16078 , n17542 );
and ( n17667 , n16087 , n17540 );
nor ( n17668 , n17666 , n17667 );
xnor ( n17669 , n17668 , n17406 );
and ( n17670 , n17665 , n17669 );
and ( n17671 , n16096 , n17020 );
and ( n17672 , n16105 , n17018 );
nor ( n17673 , n17671 , n17672 );
xnor ( n17674 , n17673 , n16938 );
and ( n17675 , n17669 , n17674 );
and ( n17676 , n17665 , n17674 );
or ( n17677 , n17670 , n17675 , n17676 );
and ( n17678 , n15982 , n16176 );
and ( n17679 , n15995 , n16174 );
nor ( n17680 , n17678 , n17679 );
xnor ( n17681 , n17680 , n16075 );
and ( n17682 , n16151 , n16084 );
and ( n17683 , n16004 , n16082 );
nor ( n17684 , n17682 , n17683 );
xnor ( n17685 , n17684 , n16092 );
and ( n17686 , n17681 , n17685 );
buf ( n17687 , n1118 );
buf ( n17688 , n17687 );
and ( n17689 , n17688 , n15984 );
and ( n17690 , n17685 , n17689 );
and ( n17691 , n17681 , n17689 );
or ( n17692 , n17686 , n17690 , n17691 );
and ( n17693 , n17677 , n17692 );
and ( n17694 , n15961 , n16782 );
and ( n17695 , n15974 , n16780 );
nor ( n17696 , n17694 , n17695 );
xnor ( n17697 , n17696 , n16696 );
and ( n17698 , n16401 , n16018 );
and ( n17699 , n16285 , n16016 );
nor ( n17700 , n17698 , n17699 );
xnor ( n17701 , n17700 , n16026 );
and ( n17702 , n17697 , n17701 );
and ( n17703 , n16592 , n16102 );
and ( n17704 , n16510 , n16100 );
nor ( n17705 , n17703 , n17704 );
xnor ( n17706 , n17705 , n16110 );
and ( n17707 , n17701 , n17706 );
and ( n17708 , n17697 , n17706 );
or ( n17709 , n17702 , n17707 , n17708 );
and ( n17710 , n17692 , n17709 );
and ( n17711 , n17677 , n17709 );
or ( n17712 , n17693 , n17710 , n17711 );
not ( n17713 , n17545 );
and ( n17714 , n17610 , n15992 );
and ( n17715 , n17355 , n15990 );
nor ( n17716 , n17714 , n17715 );
xnor ( n17717 , n17716 , n16000 );
and ( n17718 , n17713 , n17717 );
buf ( n17719 , n1117 );
buf ( n17720 , n17719 );
and ( n17721 , n17720 , n15984 );
and ( n17722 , n17717 , n17721 );
and ( n17723 , n17713 , n17721 );
or ( n17724 , n17718 , n17722 , n17723 );
and ( n17725 , n17712 , n17724 );
xor ( n17726 , n17424 , n17428 );
xor ( n17727 , n17726 , n17433 );
and ( n17728 , n17724 , n17727 );
and ( n17729 , n17712 , n17727 );
or ( n17730 , n17725 , n17728 , n17729 );
and ( n17731 , n17657 , n17730 );
xor ( n17732 , n17614 , n17616 );
xor ( n17733 , n17732 , n17619 );
and ( n17734 , n17730 , n17733 );
and ( n17735 , n17657 , n17733 );
or ( n17736 , n17731 , n17734 , n17735 );
xor ( n17737 , n17505 , n17593 );
xor ( n17738 , n17737 , n17596 );
and ( n17739 , n17736 , n17738 );
xor ( n17740 , n17622 , n17624 );
xor ( n17741 , n17740 , n17627 );
and ( n17742 , n17738 , n17741 );
and ( n17743 , n17736 , n17741 );
or ( n17744 , n17739 , n17742 , n17743 );
xor ( n17745 , n17470 , n17472 );
xor ( n17746 , n17745 , n17475 );
and ( n17747 , n17744 , n17746 );
xor ( n17748 , n17599 , n17630 );
xor ( n17749 , n17748 , n17633 );
and ( n17750 , n17746 , n17749 );
and ( n17751 , n17744 , n17749 );
or ( n17752 , n17747 , n17750 , n17751 );
and ( n17753 , n17647 , n17752 );
xor ( n17754 , n17744 , n17746 );
xor ( n17755 , n17754 , n17749 );
and ( n17756 , n16049 , n16378 );
and ( n17757 , n16058 , n16376 );
nor ( n17758 , n17756 , n17757 );
xnor ( n17759 , n17758 , n16313 );
and ( n17760 , n16995 , n16037 );
and ( n17761 , n16910 , n16035 );
nor ( n17762 , n17760 , n17761 );
xnor ( n17763 , n17762 , n16045 );
and ( n17764 , n17759 , n17763 );
and ( n17765 , n17355 , n16055 );
and ( n17766 , n17309 , n16053 );
nor ( n17767 , n17765 , n17766 );
xnor ( n17768 , n17767 , n16063 );
and ( n17769 , n17763 , n17768 );
and ( n17770 , n17759 , n17768 );
or ( n17771 , n17764 , n17769 , n17770 );
and ( n17772 , n16008 , n17246 );
and ( n17773 , n16021 , n17244 );
nor ( n17774 , n17772 , n17773 );
xnor ( n17775 , n17774 , n17191 );
and ( n17776 , n16029 , n16565 );
and ( n17777 , n16040 , n16563 );
nor ( n17778 , n17776 , n17777 );
xnor ( n17779 , n17778 , n16481 );
and ( n17780 , n17775 , n17779 );
and ( n17781 , n16792 , n15971 );
and ( n17782 , n16668 , n15969 );
nor ( n17783 , n17781 , n17782 );
xnor ( n17784 , n17783 , n15979 );
and ( n17785 , n17779 , n17784 );
and ( n17786 , n17775 , n17784 );
or ( n17787 , n17780 , n17785 , n17786 );
and ( n17788 , n17771 , n17787 );
xor ( n17789 , n17509 , n17513 );
xor ( n17790 , n17789 , n17518 );
and ( n17791 , n17787 , n17790 );
and ( n17792 , n17771 , n17790 );
or ( n17793 , n17788 , n17791 , n17792 );
xor ( n17794 , n17521 , n17537 );
xor ( n17795 , n17794 , n17546 );
and ( n17796 , n17793 , n17795 );
xor ( n17797 , n17565 , n17581 );
xor ( n17798 , n17797 , n17584 );
and ( n17799 , n17795 , n17798 );
and ( n17800 , n17793 , n17798 );
or ( n17801 , n17796 , n17799 , n17800 );
xor ( n17802 , n17497 , n17499 );
xor ( n17803 , n17802 , n17502 );
and ( n17804 , n17801 , n17803 );
xor ( n17805 , n17549 , n17587 );
xor ( n17806 , n17805 , n17590 );
and ( n17807 , n17803 , n17806 );
and ( n17808 , n17801 , n17806 );
or ( n17809 , n17804 , n17807 , n17808 );
xor ( n17810 , n17525 , n17529 );
xor ( n17811 , n17810 , n17534 );
xor ( n17812 , n17553 , n17557 );
xor ( n17813 , n17812 , n17562 );
and ( n17814 , n17811 , n17813 );
xor ( n17815 , n17569 , n17573 );
xor ( n17816 , n17815 , n17578 );
and ( n17817 , n17813 , n17816 );
and ( n17818 , n17811 , n17816 );
or ( n17819 , n17814 , n17817 , n17818 );
xor ( n17820 , n17649 , n17651 );
xor ( n17821 , n17820 , n17654 );
and ( n17822 , n17819 , n17821 );
xor ( n17823 , n17712 , n17724 );
xor ( n17824 , n17823 , n17727 );
and ( n17825 , n17821 , n17824 );
and ( n17826 , n17819 , n17824 );
or ( n17827 , n17822 , n17825 , n17826 );
xor ( n17828 , n17801 , n17803 );
xor ( n17829 , n17828 , n17806 );
and ( n17830 , n17827 , n17829 );
xor ( n17831 , n17657 , n17730 );
xor ( n17832 , n17831 , n17733 );
and ( n17833 , n17829 , n17832 );
and ( n17834 , n17827 , n17832 );
or ( n17835 , n17830 , n17833 , n17834 );
and ( n17836 , n17809 , n17835 );
xor ( n17837 , n17736 , n17738 );
xor ( n17838 , n17837 , n17741 );
and ( n17839 , n17835 , n17838 );
and ( n17840 , n17809 , n17838 );
or ( n17841 , n17836 , n17839 , n17840 );
and ( n17842 , n17755 , n17841 );
xor ( n17843 , n17809 , n17835 );
xor ( n17844 , n17843 , n17838 );
and ( n17845 , n16105 , n17246 );
and ( n17846 , n16008 , n17244 );
nor ( n17847 , n17845 , n17846 );
xnor ( n17848 , n17847 , n17191 );
and ( n17849 , n16510 , n16018 );
and ( n17850 , n16401 , n16016 );
nor ( n17851 , n17849 , n17850 );
xnor ( n17852 , n17851 , n16026 );
and ( n17853 , n17848 , n17852 );
and ( n17854 , n16668 , n16102 );
and ( n17855 , n16592 , n16100 );
nor ( n17856 , n17854 , n17855 );
xnor ( n17857 , n17856 , n16110 );
and ( n17858 , n17852 , n17857 );
and ( n17859 , n17848 , n17857 );
or ( n17860 , n17853 , n17858 , n17859 );
and ( n17861 , n16058 , n16565 );
and ( n17862 , n16029 , n16563 );
nor ( n17863 , n17861 , n17862 );
xnor ( n17864 , n17863 , n16481 );
and ( n17865 , n16910 , n15971 );
and ( n17866 , n16792 , n15969 );
nor ( n17867 , n17865 , n17866 );
xnor ( n17868 , n17867 , n15979 );
and ( n17869 , n17864 , n17868 );
and ( n17870 , n17309 , n16037 );
and ( n17871 , n16995 , n16035 );
nor ( n17872 , n17870 , n17871 );
xnor ( n17873 , n17872 , n16045 );
and ( n17874 , n17868 , n17873 );
and ( n17875 , n17864 , n17873 );
or ( n17876 , n17869 , n17874 , n17875 );
and ( n17877 , n17860 , n17876 );
and ( n17878 , n16040 , n16782 );
and ( n17879 , n15961 , n16780 );
nor ( n17880 , n17878 , n17879 );
xnor ( n17881 , n17880 , n16696 );
and ( n17882 , n16004 , n16176 );
and ( n17883 , n15982 , n16174 );
nor ( n17884 , n17882 , n17883 );
xnor ( n17885 , n17884 , n16075 );
and ( n17886 , n17881 , n17885 );
and ( n17887 , n16285 , n16084 );
and ( n17888 , n16151 , n16082 );
nor ( n17889 , n17887 , n17888 );
xnor ( n17890 , n17889 , n16092 );
and ( n17891 , n17885 , n17890 );
and ( n17892 , n17881 , n17890 );
or ( n17893 , n17886 , n17891 , n17892 );
and ( n17894 , n17876 , n17893 );
and ( n17895 , n17860 , n17893 );
or ( n17896 , n17877 , n17894 , n17895 );
and ( n17897 , n16021 , n17542 );
and ( n17898 , n16078 , n17540 );
nor ( n17899 , n17897 , n17898 );
xnor ( n17900 , n17899 , n17406 );
and ( n17901 , n15974 , n17020 );
and ( n17902 , n16096 , n17018 );
nor ( n17903 , n17901 , n17902 );
xnor ( n17904 , n17903 , n16938 );
and ( n17905 , n17900 , n17904 );
buf ( n17906 , n1119 );
buf ( n17907 , n17906 );
and ( n17908 , n17907 , n15984 );
and ( n17909 , n17904 , n17908 );
and ( n17910 , n17900 , n17908 );
or ( n17911 , n17905 , n17909 , n17910 );
xor ( n17912 , n17403 , n17659 );
xor ( n17913 , n17659 , n17661 );
not ( n17914 , n17913 );
and ( n17915 , n17912 , n17914 );
and ( n17916 , n16087 , n17915 );
not ( n17917 , n17916 );
xnor ( n17918 , n17917 , n17664 );
buf ( n17919 , n17918 );
and ( n17920 , n17911 , n17919 );
and ( n17921 , n17720 , n15992 );
and ( n17922 , n17610 , n15990 );
nor ( n17923 , n17921 , n17922 );
xnor ( n17924 , n17923 , n16000 );
and ( n17925 , n17919 , n17924 );
and ( n17926 , n17911 , n17924 );
or ( n17927 , n17920 , n17925 , n17926 );
and ( n17928 , n17896 , n17927 );
xor ( n17929 , n17713 , n17717 );
xor ( n17930 , n17929 , n17721 );
and ( n17931 , n17927 , n17930 );
and ( n17932 , n17896 , n17930 );
or ( n17933 , n17928 , n17931 , n17932 );
and ( n17934 , n15995 , n16378 );
and ( n17935 , n16049 , n16376 );
nor ( n17936 , n17934 , n17935 );
xnor ( n17937 , n17936 , n16313 );
and ( n17938 , n17610 , n16055 );
and ( n17939 , n17355 , n16053 );
nor ( n17940 , n17938 , n17939 );
xnor ( n17941 , n17940 , n16063 );
and ( n17942 , n17937 , n17941 );
and ( n17943 , n17688 , n15992 );
and ( n17944 , n17720 , n15990 );
nor ( n17945 , n17943 , n17944 );
xnor ( n17946 , n17945 , n16000 );
and ( n17947 , n17941 , n17946 );
and ( n17948 , n17937 , n17946 );
or ( n17949 , n17942 , n17947 , n17948 );
xor ( n17950 , n17665 , n17669 );
xor ( n17951 , n17950 , n17674 );
and ( n17952 , n17949 , n17951 );
xor ( n17953 , n17681 , n17685 );
xor ( n17954 , n17953 , n17689 );
and ( n17955 , n17951 , n17954 );
and ( n17956 , n17949 , n17954 );
or ( n17957 , n17952 , n17955 , n17956 );
xor ( n17958 , n17677 , n17692 );
xor ( n17959 , n17958 , n17709 );
and ( n17960 , n17957 , n17959 );
xor ( n17961 , n17771 , n17787 );
xor ( n17962 , n17961 , n17790 );
and ( n17963 , n17959 , n17962 );
and ( n17964 , n17957 , n17962 );
or ( n17965 , n17960 , n17963 , n17964 );
and ( n17966 , n17933 , n17965 );
xor ( n17967 , n17793 , n17795 );
xor ( n17968 , n17967 , n17798 );
and ( n17969 , n17965 , n17968 );
and ( n17970 , n17933 , n17968 );
or ( n17971 , n17966 , n17969 , n17970 );
xor ( n17972 , n17759 , n17763 );
xor ( n17973 , n17972 , n17768 );
xor ( n17974 , n17697 , n17701 );
xor ( n17975 , n17974 , n17706 );
and ( n17976 , n17973 , n17975 );
xor ( n17977 , n17775 , n17779 );
xor ( n17978 , n17977 , n17784 );
and ( n17979 , n17975 , n17978 );
and ( n17980 , n17973 , n17978 );
or ( n17981 , n17976 , n17979 , n17980 );
and ( n17982 , n15961 , n17020 );
and ( n17983 , n15974 , n17018 );
nor ( n17984 , n17982 , n17983 );
xnor ( n17985 , n17984 , n16938 );
and ( n17986 , n16401 , n16084 );
and ( n17987 , n16285 , n16082 );
nor ( n17988 , n17986 , n17987 );
xnor ( n17989 , n17988 , n16092 );
and ( n17990 , n17985 , n17989 );
and ( n17991 , n16592 , n16018 );
and ( n17992 , n16510 , n16016 );
nor ( n17993 , n17991 , n17992 );
xnor ( n17994 , n17993 , n16026 );
and ( n17995 , n17989 , n17994 );
and ( n17996 , n17985 , n17994 );
or ( n17997 , n17990 , n17995 , n17996 );
and ( n17998 , n16008 , n17542 );
and ( n17999 , n16021 , n17540 );
nor ( n18000 , n17998 , n17999 );
xnor ( n18001 , n18000 , n17406 );
and ( n18002 , n16029 , n16782 );
and ( n18003 , n16040 , n16780 );
nor ( n18004 , n18002 , n18003 );
xnor ( n18005 , n18004 , n16696 );
and ( n18006 , n18001 , n18005 );
and ( n18007 , n16792 , n16102 );
and ( n18008 , n16668 , n16100 );
nor ( n18009 , n18007 , n18008 );
xnor ( n18010 , n18009 , n16110 );
and ( n18011 , n18005 , n18010 );
and ( n18012 , n18001 , n18010 );
or ( n18013 , n18006 , n18011 , n18012 );
and ( n18014 , n17997 , n18013 );
and ( n18015 , n16078 , n17915 );
and ( n18016 , n16087 , n17913 );
nor ( n18017 , n18015 , n18016 );
xnor ( n18018 , n18017 , n17664 );
and ( n18019 , n16096 , n17246 );
and ( n18020 , n16105 , n17244 );
nor ( n18021 , n18019 , n18020 );
xnor ( n18022 , n18021 , n17191 );
and ( n18023 , n18018 , n18022 );
and ( n18024 , n16151 , n16176 );
and ( n18025 , n16004 , n16174 );
nor ( n18026 , n18024 , n18025 );
xnor ( n18027 , n18026 , n16075 );
and ( n18028 , n18022 , n18027 );
and ( n18029 , n18018 , n18027 );
or ( n18030 , n18023 , n18028 , n18029 );
and ( n18031 , n18013 , n18030 );
and ( n18032 , n17997 , n18030 );
or ( n18033 , n18014 , n18031 , n18032 );
and ( n18034 , n15982 , n16378 );
and ( n18035 , n15995 , n16376 );
nor ( n18036 , n18034 , n18035 );
xnor ( n18037 , n18036 , n16313 );
and ( n18038 , n17907 , n15992 );
and ( n18039 , n17688 , n15990 );
nor ( n18040 , n18038 , n18039 );
xnor ( n18041 , n18040 , n16000 );
and ( n18042 , n18037 , n18041 );
buf ( n18043 , n1120 );
buf ( n18044 , n18043 );
and ( n18045 , n18044 , n15984 );
and ( n18046 , n18041 , n18045 );
and ( n18047 , n18037 , n18045 );
or ( n18048 , n18042 , n18046 , n18047 );
not ( n18049 , n17661 );
buf ( n18050 , n18049 );
and ( n18051 , n18048 , n18050 );
not ( n18052 , n17918 );
and ( n18053 , n18050 , n18052 );
and ( n18054 , n18048 , n18052 );
or ( n18055 , n18051 , n18053 , n18054 );
and ( n18056 , n18033 , n18055 );
xor ( n18057 , n17911 , n17919 );
xor ( n18058 , n18057 , n17924 );
and ( n18059 , n18055 , n18058 );
and ( n18060 , n18033 , n18058 );
or ( n18061 , n18056 , n18059 , n18060 );
and ( n18062 , n17981 , n18061 );
xor ( n18063 , n17811 , n17813 );
xor ( n18064 , n18063 , n17816 );
and ( n18065 , n18061 , n18064 );
and ( n18066 , n17981 , n18064 );
or ( n18067 , n18062 , n18065 , n18066 );
xor ( n18068 , n17900 , n17904 );
xor ( n18069 , n18068 , n17908 );
xor ( n18070 , n17848 , n17852 );
xor ( n18071 , n18070 , n17857 );
and ( n18072 , n18069 , n18071 );
xor ( n18073 , n17864 , n17868 );
xor ( n18074 , n18073 , n17873 );
and ( n18075 , n18071 , n18074 );
and ( n18076 , n18069 , n18074 );
or ( n18077 , n18072 , n18075 , n18076 );
and ( n18078 , n16049 , n16565 );
and ( n18079 , n16058 , n16563 );
nor ( n18080 , n18078 , n18079 );
xnor ( n18081 , n18080 , n16481 );
and ( n18082 , n16995 , n15971 );
and ( n18083 , n16910 , n15969 );
nor ( n18084 , n18082 , n18083 );
xnor ( n18085 , n18084 , n15979 );
and ( n18086 , n18081 , n18085 );
and ( n18087 , n17355 , n16037 );
and ( n18088 , n17309 , n16035 );
nor ( n18089 , n18087 , n18088 );
xnor ( n18090 , n18089 , n16045 );
and ( n18091 , n18085 , n18090 );
and ( n18092 , n18081 , n18090 );
or ( n18093 , n18086 , n18091 , n18092 );
xor ( n18094 , n17881 , n17885 );
xor ( n18095 , n18094 , n17890 );
and ( n18096 , n18093 , n18095 );
xor ( n18097 , n17937 , n17941 );
xor ( n18098 , n18097 , n17946 );
and ( n18099 , n18095 , n18098 );
and ( n18100 , n18093 , n18098 );
or ( n18101 , n18096 , n18099 , n18100 );
and ( n18102 , n18077 , n18101 );
xor ( n18103 , n17860 , n17876 );
xor ( n18104 , n18103 , n17893 );
and ( n18105 , n18101 , n18104 );
and ( n18106 , n18077 , n18104 );
or ( n18107 , n18102 , n18105 , n18106 );
xor ( n18108 , n17896 , n17927 );
xor ( n18109 , n18108 , n17930 );
and ( n18110 , n18107 , n18109 );
xor ( n18111 , n17957 , n17959 );
xor ( n18112 , n18111 , n17962 );
and ( n18113 , n18109 , n18112 );
and ( n18114 , n18107 , n18112 );
or ( n18115 , n18110 , n18113 , n18114 );
and ( n18116 , n18067 , n18115 );
xor ( n18117 , n17819 , n17821 );
xor ( n18118 , n18117 , n17824 );
and ( n18119 , n18115 , n18118 );
and ( n18120 , n18067 , n18118 );
or ( n18121 , n18116 , n18119 , n18120 );
and ( n18122 , n17971 , n18121 );
xor ( n18123 , n17827 , n17829 );
xor ( n18124 , n18123 , n17832 );
and ( n18125 , n18121 , n18124 );
and ( n18126 , n17971 , n18124 );
or ( n18127 , n18122 , n18125 , n18126 );
and ( n18128 , n17844 , n18127 );
xor ( n18129 , n17971 , n18121 );
xor ( n18130 , n18129 , n18124 );
and ( n18131 , n15995 , n16565 );
and ( n18132 , n16049 , n16563 );
nor ( n18133 , n18131 , n18132 );
xnor ( n18134 , n18133 , n16481 );
and ( n18135 , n16910 , n16102 );
and ( n18136 , n16792 , n16100 );
nor ( n18137 , n18135 , n18136 );
xnor ( n18138 , n18137 , n16110 );
and ( n18139 , n18134 , n18138 );
and ( n18140 , n17309 , n15971 );
and ( n18141 , n16995 , n15969 );
nor ( n18142 , n18140 , n18141 );
xnor ( n18143 , n18142 , n15979 );
and ( n18144 , n18138 , n18143 );
and ( n18145 , n18134 , n18143 );
or ( n18146 , n18139 , n18144 , n18145 );
and ( n18147 , n16040 , n17020 );
and ( n18148 , n15961 , n17018 );
nor ( n18149 , n18147 , n18148 );
xnor ( n18150 , n18149 , n16938 );
and ( n18151 , n16285 , n16176 );
and ( n18152 , n16151 , n16174 );
nor ( n18153 , n18151 , n18152 );
xnor ( n18154 , n18153 , n16075 );
and ( n18155 , n18150 , n18154 );
and ( n18156 , n16510 , n16084 );
and ( n18157 , n16401 , n16082 );
nor ( n18158 , n18156 , n18157 );
xnor ( n18159 , n18158 , n16092 );
and ( n18160 , n18154 , n18159 );
and ( n18161 , n18150 , n18159 );
or ( n18162 , n18155 , n18160 , n18161 );
and ( n18163 , n18146 , n18162 );
and ( n18164 , n15974 , n17246 );
and ( n18165 , n16096 , n17244 );
nor ( n18166 , n18164 , n18165 );
xnor ( n18167 , n18166 , n17191 );
and ( n18168 , n16004 , n16378 );
and ( n18169 , n15982 , n16376 );
nor ( n18170 , n18168 , n18169 );
xnor ( n18171 , n18170 , n16313 );
and ( n18172 , n18167 , n18171 );
and ( n18173 , n18044 , n15992 );
and ( n18174 , n17907 , n15990 );
nor ( n18175 , n18173 , n18174 );
xnor ( n18176 , n18175 , n16000 );
and ( n18177 , n18171 , n18176 );
and ( n18178 , n18167 , n18176 );
or ( n18179 , n18172 , n18177 , n18178 );
and ( n18180 , n18162 , n18179 );
and ( n18181 , n18146 , n18179 );
or ( n18182 , n18163 , n18180 , n18181 );
buf ( n18183 , n1185 );
buf ( n18184 , n18183 );
xor ( n18185 , n17661 , n18184 );
not ( n18186 , n18184 );
and ( n18187 , n18185 , n18186 );
and ( n18188 , n16087 , n18187 );
not ( n18189 , n18188 );
xnor ( n18190 , n18189 , n17661 );
and ( n18191 , n16021 , n17915 );
and ( n18192 , n16078 , n17913 );
nor ( n18193 , n18191 , n18192 );
xnor ( n18194 , n18193 , n17664 );
and ( n18195 , n18190 , n18194 );
buf ( n18196 , n1121 );
buf ( n18197 , n18196 );
and ( n18198 , n18197 , n15984 );
and ( n18199 , n18194 , n18198 );
and ( n18200 , n18190 , n18198 );
or ( n18201 , n18195 , n18199 , n18200 );
and ( n18202 , n18201 , n17661 );
and ( n18203 , n17720 , n16055 );
and ( n18204 , n17610 , n16053 );
nor ( n18205 , n18203 , n18204 );
xnor ( n18206 , n18205 , n16063 );
and ( n18207 , n17661 , n18206 );
and ( n18208 , n18201 , n18206 );
or ( n18209 , n18202 , n18207 , n18208 );
and ( n18210 , n18182 , n18209 );
xor ( n18211 , n17997 , n18013 );
xor ( n18212 , n18211 , n18030 );
and ( n18213 , n18209 , n18212 );
and ( n18214 , n18182 , n18212 );
or ( n18215 , n18210 , n18213 , n18214 );
and ( n18216 , n16105 , n17542 );
and ( n18217 , n16008 , n17540 );
nor ( n18218 , n18216 , n18217 );
xnor ( n18219 , n18218 , n17406 );
and ( n18220 , n16058 , n16782 );
and ( n18221 , n16029 , n16780 );
nor ( n18222 , n18220 , n18221 );
xnor ( n18223 , n18222 , n16696 );
and ( n18224 , n18219 , n18223 );
and ( n18225 , n16668 , n16018 );
and ( n18226 , n16592 , n16016 );
nor ( n18227 , n18225 , n18226 );
xnor ( n18228 , n18227 , n16026 );
and ( n18229 , n18223 , n18228 );
and ( n18230 , n18219 , n18228 );
or ( n18231 , n18224 , n18229 , n18230 );
xor ( n18232 , n18037 , n18041 );
xor ( n18233 , n18232 , n18045 );
and ( n18234 , n18231 , n18233 );
xor ( n18235 , n18081 , n18085 );
xor ( n18236 , n18235 , n18090 );
and ( n18237 , n18233 , n18236 );
and ( n18238 , n18231 , n18236 );
or ( n18239 , n18234 , n18237 , n18238 );
xor ( n18240 , n17985 , n17989 );
xor ( n18241 , n18240 , n17994 );
xor ( n18242 , n18001 , n18005 );
xor ( n18243 , n18242 , n18010 );
and ( n18244 , n18241 , n18243 );
xor ( n18245 , n18018 , n18022 );
xor ( n18246 , n18245 , n18027 );
and ( n18247 , n18243 , n18246 );
and ( n18248 , n18241 , n18246 );
or ( n18249 , n18244 , n18247 , n18248 );
and ( n18250 , n18239 , n18249 );
xor ( n18251 , n18048 , n18050 );
xor ( n18252 , n18251 , n18052 );
and ( n18253 , n18249 , n18252 );
and ( n18254 , n18239 , n18252 );
or ( n18255 , n18250 , n18253 , n18254 );
and ( n18256 , n18215 , n18255 );
xor ( n18257 , n18077 , n18101 );
xor ( n18258 , n18257 , n18104 );
and ( n18259 , n18255 , n18258 );
and ( n18260 , n18215 , n18258 );
or ( n18261 , n18256 , n18259 , n18260 );
xor ( n18262 , n17949 , n17951 );
xor ( n18263 , n18262 , n17954 );
xor ( n18264 , n17973 , n17975 );
xor ( n18265 , n18264 , n17978 );
and ( n18266 , n18263 , n18265 );
xor ( n18267 , n18033 , n18055 );
xor ( n18268 , n18267 , n18058 );
and ( n18269 , n18265 , n18268 );
and ( n18270 , n18263 , n18268 );
or ( n18271 , n18266 , n18269 , n18270 );
and ( n18272 , n18261 , n18271 );
xor ( n18273 , n17981 , n18061 );
xor ( n18274 , n18273 , n18064 );
and ( n18275 , n18271 , n18274 );
and ( n18276 , n18261 , n18274 );
or ( n18277 , n18272 , n18275 , n18276 );
xor ( n18278 , n17933 , n17965 );
xor ( n18279 , n18278 , n17968 );
and ( n18280 , n18277 , n18279 );
xor ( n18281 , n18067 , n18115 );
xor ( n18282 , n18281 , n18118 );
and ( n18283 , n18279 , n18282 );
and ( n18284 , n18277 , n18282 );
or ( n18285 , n18280 , n18283 , n18284 );
and ( n18286 , n18130 , n18285 );
xor ( n18287 , n18277 , n18279 );
xor ( n18288 , n18287 , n18282 );
xor ( n18289 , n18134 , n18138 );
xor ( n18290 , n18289 , n18143 );
xor ( n18291 , n18219 , n18223 );
xor ( n18292 , n18291 , n18228 );
and ( n18293 , n18290 , n18292 );
xor ( n18294 , n18150 , n18154 );
xor ( n18295 , n18294 , n18159 );
and ( n18296 , n18292 , n18295 );
and ( n18297 , n18290 , n18295 );
or ( n18298 , n18293 , n18296 , n18297 );
xor ( n18299 , n18146 , n18162 );
xor ( n18300 , n18299 , n18179 );
and ( n18301 , n18298 , n18300 );
xor ( n18302 , n18201 , n17661 );
xor ( n18303 , n18302 , n18206 );
and ( n18304 , n18300 , n18303 );
and ( n18305 , n18298 , n18303 );
or ( n18306 , n18301 , n18304 , n18305 );
xor ( n18307 , n18069 , n18071 );
xor ( n18308 , n18307 , n18074 );
and ( n18309 , n18306 , n18308 );
xor ( n18310 , n18093 , n18095 );
xor ( n18311 , n18310 , n18098 );
and ( n18312 , n18308 , n18311 );
and ( n18313 , n18306 , n18311 );
or ( n18314 , n18309 , n18312 , n18313 );
and ( n18315 , n16096 , n17542 );
and ( n18316 , n16105 , n17540 );
nor ( n18317 , n18315 , n18316 );
xnor ( n18318 , n18317 , n17406 );
and ( n18319 , n16592 , n16084 );
and ( n18320 , n16510 , n16082 );
nor ( n18321 , n18319 , n18320 );
xnor ( n18322 , n18321 , n16092 );
and ( n18323 , n18318 , n18322 );
and ( n18324 , n16792 , n16018 );
and ( n18325 , n16668 , n16016 );
nor ( n18326 , n18324 , n18325 );
xnor ( n18327 , n18326 , n16026 );
and ( n18328 , n18322 , n18327 );
and ( n18329 , n18318 , n18327 );
or ( n18330 , n18323 , n18328 , n18329 );
and ( n18331 , n16008 , n17915 );
and ( n18332 , n16021 , n17913 );
nor ( n18333 , n18331 , n18332 );
xnor ( n18334 , n18333 , n17664 );
and ( n18335 , n15961 , n17246 );
and ( n18336 , n15974 , n17244 );
nor ( n18337 , n18335 , n18336 );
xnor ( n18338 , n18337 , n17191 );
and ( n18339 , n18334 , n18338 );
and ( n18340 , n18197 , n15992 );
and ( n18341 , n18044 , n15990 );
nor ( n18342 , n18340 , n18341 );
xnor ( n18343 , n18342 , n16000 );
and ( n18344 , n18338 , n18343 );
and ( n18345 , n18334 , n18343 );
or ( n18346 , n18339 , n18344 , n18345 );
and ( n18347 , n18330 , n18346 );
and ( n18348 , n16029 , n17020 );
and ( n18349 , n16040 , n17018 );
nor ( n18350 , n18348 , n18349 );
xnor ( n18351 , n18350 , n16938 );
and ( n18352 , n16151 , n16378 );
and ( n18353 , n16004 , n16376 );
nor ( n18354 , n18352 , n18353 );
xnor ( n18355 , n18354 , n16313 );
and ( n18356 , n18351 , n18355 );
and ( n18357 , n16401 , n16176 );
and ( n18358 , n16285 , n16174 );
nor ( n18359 , n18357 , n18358 );
xnor ( n18360 , n18359 , n16075 );
and ( n18361 , n18355 , n18360 );
and ( n18362 , n18351 , n18360 );
or ( n18363 , n18356 , n18361 , n18362 );
and ( n18364 , n18346 , n18363 );
and ( n18365 , n18330 , n18363 );
or ( n18366 , n18347 , n18364 , n18365 );
and ( n18367 , n16078 , n18187 );
and ( n18368 , n16087 , n18184 );
nor ( n18369 , n18367 , n18368 );
xnor ( n18370 , n18369 , n17661 );
and ( n18371 , n18197 , n15990 );
not ( n18372 , n18371 );
and ( n18373 , n18372 , n16000 );
and ( n18374 , n18370 , n18373 );
and ( n18375 , n17610 , n16037 );
and ( n18376 , n17355 , n16035 );
nor ( n18377 , n18375 , n18376 );
xnor ( n18378 , n18377 , n16045 );
and ( n18379 , n18374 , n18378 );
and ( n18380 , n17688 , n16055 );
and ( n18381 , n17720 , n16053 );
nor ( n18382 , n18380 , n18381 );
xnor ( n18383 , n18382 , n16063 );
and ( n18384 , n18378 , n18383 );
and ( n18385 , n18374 , n18383 );
or ( n18386 , n18379 , n18384 , n18385 );
and ( n18387 , n18366 , n18386 );
and ( n18388 , n16049 , n16782 );
and ( n18389 , n16058 , n16780 );
nor ( n18390 , n18388 , n18389 );
xnor ( n18391 , n18390 , n16696 );
and ( n18392 , n16995 , n16102 );
and ( n18393 , n16910 , n16100 );
nor ( n18394 , n18392 , n18393 );
xnor ( n18395 , n18394 , n16110 );
and ( n18396 , n18391 , n18395 );
and ( n18397 , n17355 , n15971 );
and ( n18398 , n17309 , n15969 );
nor ( n18399 , n18397 , n18398 );
xnor ( n18400 , n18399 , n15979 );
and ( n18401 , n18395 , n18400 );
and ( n18402 , n18391 , n18400 );
or ( n18403 , n18396 , n18401 , n18402 );
and ( n18404 , n15982 , n16565 );
and ( n18405 , n15995 , n16563 );
nor ( n18406 , n18404 , n18405 );
xnor ( n18407 , n18406 , n16481 );
and ( n18408 , n17720 , n16037 );
and ( n18409 , n17610 , n16035 );
nor ( n18410 , n18408 , n18409 );
xnor ( n18411 , n18410 , n16045 );
and ( n18412 , n18407 , n18411 );
and ( n18413 , n17907 , n16055 );
and ( n18414 , n17688 , n16053 );
nor ( n18415 , n18413 , n18414 );
xnor ( n18416 , n18415 , n16063 );
and ( n18417 , n18411 , n18416 );
and ( n18418 , n18407 , n18416 );
or ( n18419 , n18412 , n18417 , n18418 );
and ( n18420 , n18403 , n18419 );
xor ( n18421 , n18190 , n18194 );
xor ( n18422 , n18421 , n18198 );
and ( n18423 , n18419 , n18422 );
and ( n18424 , n18403 , n18422 );
or ( n18425 , n18420 , n18423 , n18424 );
and ( n18426 , n18386 , n18425 );
and ( n18427 , n18366 , n18425 );
or ( n18428 , n18387 , n18426 , n18427 );
xor ( n18429 , n18182 , n18209 );
xor ( n18430 , n18429 , n18212 );
and ( n18431 , n18428 , n18430 );
xor ( n18432 , n18239 , n18249 );
xor ( n18433 , n18432 , n18252 );
and ( n18434 , n18430 , n18433 );
and ( n18435 , n18428 , n18433 );
or ( n18436 , n18431 , n18434 , n18435 );
and ( n18437 , n18314 , n18436 );
xor ( n18438 , n18263 , n18265 );
xor ( n18439 , n18438 , n18268 );
and ( n18440 , n18436 , n18439 );
and ( n18441 , n18314 , n18439 );
or ( n18442 , n18437 , n18440 , n18441 );
xor ( n18443 , n18107 , n18109 );
xor ( n18444 , n18443 , n18112 );
and ( n18445 , n18442 , n18444 );
xor ( n18446 , n18261 , n18271 );
xor ( n18447 , n18446 , n18274 );
and ( n18448 , n18444 , n18447 );
and ( n18449 , n18442 , n18447 );
or ( n18450 , n18445 , n18448 , n18449 );
and ( n18451 , n18288 , n18450 );
xor ( n18452 , n18442 , n18444 );
xor ( n18453 , n18452 , n18447 );
and ( n18454 , n16058 , n17020 );
and ( n18455 , n16029 , n17018 );
nor ( n18456 , n18454 , n18455 );
xnor ( n18457 , n18456 , n16938 );
and ( n18458 , n16668 , n16084 );
and ( n18459 , n16592 , n16082 );
nor ( n18460 , n18458 , n18459 );
xnor ( n18461 , n18460 , n16092 );
and ( n18462 , n18457 , n18461 );
and ( n18463 , n16910 , n16018 );
and ( n18464 , n16792 , n16016 );
nor ( n18465 , n18463 , n18464 );
xnor ( n18466 , n18465 , n16026 );
and ( n18467 , n18461 , n18466 );
and ( n18468 , n18457 , n18466 );
or ( n18469 , n18462 , n18467 , n18468 );
and ( n18470 , n16004 , n16565 );
and ( n18471 , n15982 , n16563 );
nor ( n18472 , n18470 , n18471 );
xnor ( n18473 , n18472 , n16481 );
and ( n18474 , n17610 , n15971 );
and ( n18475 , n17355 , n15969 );
nor ( n18476 , n18474 , n18475 );
xnor ( n18477 , n18476 , n15979 );
and ( n18478 , n18473 , n18477 );
and ( n18479 , n17688 , n16037 );
and ( n18480 , n17720 , n16035 );
nor ( n18481 , n18479 , n18480 );
xnor ( n18482 , n18481 , n16045 );
and ( n18483 , n18477 , n18482 );
and ( n18484 , n18473 , n18482 );
or ( n18485 , n18478 , n18483 , n18484 );
and ( n18486 , n18469 , n18485 );
and ( n18487 , n15974 , n17542 );
and ( n18488 , n16096 , n17540 );
nor ( n18489 , n18487 , n18488 );
xnor ( n18490 , n18489 , n17406 );
and ( n18491 , n15995 , n16782 );
and ( n18492 , n16049 , n16780 );
nor ( n18493 , n18491 , n18492 );
xnor ( n18494 , n18493 , n16696 );
and ( n18495 , n18490 , n18494 );
and ( n18496 , n17309 , n16102 );
and ( n18497 , n16995 , n16100 );
nor ( n18498 , n18496 , n18497 );
xnor ( n18499 , n18498 , n16110 );
and ( n18500 , n18494 , n18499 );
and ( n18501 , n18490 , n18499 );
or ( n18502 , n18495 , n18500 , n18501 );
and ( n18503 , n18485 , n18502 );
and ( n18504 , n18469 , n18502 );
or ( n18505 , n18486 , n18503 , n18504 );
xor ( n18506 , n18167 , n18171 );
xor ( n18507 , n18506 , n18176 );
and ( n18508 , n18505 , n18507 );
xor ( n18509 , n18374 , n18378 );
xor ( n18510 , n18509 , n18383 );
and ( n18511 , n18507 , n18510 );
and ( n18512 , n18505 , n18510 );
or ( n18513 , n18508 , n18511 , n18512 );
xor ( n18514 , n18231 , n18233 );
xor ( n18515 , n18514 , n18236 );
and ( n18516 , n18513 , n18515 );
xor ( n18517 , n18241 , n18243 );
xor ( n18518 , n18517 , n18246 );
and ( n18519 , n18515 , n18518 );
and ( n18520 , n18513 , n18518 );
or ( n18521 , n18516 , n18519 , n18520 );
xor ( n18522 , n18370 , n18373 );
and ( n18523 , n16040 , n17246 );
and ( n18524 , n15961 , n17244 );
nor ( n18525 , n18523 , n18524 );
xnor ( n18526 , n18525 , n17191 );
and ( n18527 , n16285 , n16378 );
and ( n18528 , n16151 , n16376 );
nor ( n18529 , n18527 , n18528 );
xnor ( n18530 , n18529 , n16313 );
and ( n18531 , n18526 , n18530 );
and ( n18532 , n16510 , n16176 );
and ( n18533 , n16401 , n16174 );
nor ( n18534 , n18532 , n18533 );
xnor ( n18535 , n18534 , n16075 );
and ( n18536 , n18530 , n18535 );
and ( n18537 , n18526 , n18535 );
or ( n18538 , n18531 , n18536 , n18537 );
and ( n18539 , n18522 , n18538 );
and ( n18540 , n16021 , n18187 );
and ( n18541 , n16078 , n18184 );
nor ( n18542 , n18540 , n18541 );
xnor ( n18543 , n18542 , n17661 );
and ( n18544 , n16105 , n17915 );
and ( n18545 , n16008 , n17913 );
nor ( n18546 , n18544 , n18545 );
xnor ( n18547 , n18546 , n17664 );
and ( n18548 , n18543 , n18547 );
and ( n18549 , n18547 , n18371 );
and ( n18550 , n18543 , n18371 );
or ( n18551 , n18548 , n18549 , n18550 );
and ( n18552 , n18538 , n18551 );
and ( n18553 , n18522 , n18551 );
or ( n18554 , n18539 , n18552 , n18553 );
xor ( n18555 , n18334 , n18338 );
xor ( n18556 , n18555 , n18343 );
xor ( n18557 , n18407 , n18411 );
xor ( n18558 , n18557 , n18416 );
and ( n18559 , n18556 , n18558 );
xor ( n18560 , n18351 , n18355 );
xor ( n18561 , n18560 , n18360 );
and ( n18562 , n18558 , n18561 );
and ( n18563 , n18556 , n18561 );
or ( n18564 , n18559 , n18562 , n18563 );
and ( n18565 , n18554 , n18564 );
xor ( n18566 , n18403 , n18419 );
xor ( n18567 , n18566 , n18422 );
and ( n18568 , n18564 , n18567 );
and ( n18569 , n18554 , n18567 );
or ( n18570 , n18565 , n18568 , n18569 );
xor ( n18571 , n18366 , n18386 );
xor ( n18572 , n18571 , n18425 );
and ( n18573 , n18570 , n18572 );
xor ( n18574 , n18298 , n18300 );
xor ( n18575 , n18574 , n18303 );
and ( n18576 , n18572 , n18575 );
and ( n18577 , n18570 , n18575 );
or ( n18578 , n18573 , n18576 , n18577 );
and ( n18579 , n18521 , n18578 );
xor ( n18580 , n18306 , n18308 );
xor ( n18581 , n18580 , n18311 );
and ( n18582 , n18578 , n18581 );
and ( n18583 , n18521 , n18581 );
or ( n18584 , n18579 , n18582 , n18583 );
xor ( n18585 , n18215 , n18255 );
xor ( n18586 , n18585 , n18258 );
and ( n18587 , n18584 , n18586 );
xor ( n18588 , n18314 , n18436 );
xor ( n18589 , n18588 , n18439 );
and ( n18590 , n18586 , n18589 );
and ( n18591 , n18584 , n18589 );
or ( n18592 , n18587 , n18590 , n18591 );
and ( n18593 , n18453 , n18592 );
and ( n18594 , n15961 , n17542 );
and ( n18595 , n15974 , n17540 );
nor ( n18596 , n18594 , n18595 );
xnor ( n18597 , n18596 , n17406 );
and ( n18598 , n15982 , n16782 );
and ( n18599 , n15995 , n16780 );
nor ( n18600 , n18598 , n18599 );
xnor ( n18601 , n18600 , n16696 );
and ( n18602 , n18597 , n18601 );
and ( n18603 , n16995 , n16018 );
and ( n18604 , n16910 , n16016 );
nor ( n18605 , n18603 , n18604 );
xnor ( n18606 , n18605 , n16026 );
and ( n18607 , n18601 , n18606 );
and ( n18608 , n18597 , n18606 );
or ( n18609 , n18602 , n18607 , n18608 );
and ( n18610 , n16151 , n16565 );
and ( n18611 , n16004 , n16563 );
nor ( n18612 , n18610 , n18611 );
xnor ( n18613 , n18612 , n16481 );
and ( n18614 , n17355 , n16102 );
and ( n18615 , n17309 , n16100 );
nor ( n18616 , n18614 , n18615 );
xnor ( n18617 , n18616 , n16110 );
and ( n18618 , n18613 , n18617 );
and ( n18619 , n17720 , n15971 );
and ( n18620 , n17610 , n15969 );
nor ( n18621 , n18619 , n18620 );
xnor ( n18622 , n18621 , n15979 );
and ( n18623 , n18617 , n18622 );
and ( n18624 , n18613 , n18622 );
or ( n18625 , n18618 , n18623 , n18624 );
and ( n18626 , n18609 , n18625 );
and ( n18627 , n16049 , n17020 );
and ( n18628 , n16058 , n17018 );
nor ( n18629 , n18627 , n18628 );
xnor ( n18630 , n18629 , n16938 );
and ( n18631 , n16592 , n16176 );
and ( n18632 , n16510 , n16174 );
nor ( n18633 , n18631 , n18632 );
xnor ( n18634 , n18633 , n16075 );
and ( n18635 , n18630 , n18634 );
and ( n18636 , n16792 , n16084 );
and ( n18637 , n16668 , n16082 );
nor ( n18638 , n18636 , n18637 );
xnor ( n18639 , n18638 , n16092 );
and ( n18640 , n18634 , n18639 );
and ( n18641 , n18630 , n18639 );
or ( n18642 , n18635 , n18640 , n18641 );
and ( n18643 , n18625 , n18642 );
and ( n18644 , n18609 , n18642 );
or ( n18645 , n18626 , n18643 , n18644 );
xor ( n18646 , n18318 , n18322 );
xor ( n18647 , n18646 , n18327 );
and ( n18648 , n18645 , n18647 );
xor ( n18649 , n18391 , n18395 );
xor ( n18650 , n18649 , n18400 );
and ( n18651 , n18647 , n18650 );
and ( n18652 , n18645 , n18650 );
or ( n18653 , n18648 , n18651 , n18652 );
xor ( n18654 , n18330 , n18346 );
xor ( n18655 , n18654 , n18363 );
and ( n18656 , n18653 , n18655 );
xor ( n18657 , n18290 , n18292 );
xor ( n18658 , n18657 , n18295 );
and ( n18659 , n18655 , n18658 );
and ( n18660 , n18653 , n18658 );
or ( n18661 , n18656 , n18659 , n18660 );
and ( n18662 , n16096 , n17915 );
and ( n18663 , n16105 , n17913 );
nor ( n18664 , n18662 , n18663 );
xnor ( n18665 , n18664 , n17664 );
and ( n18666 , n16029 , n17246 );
and ( n18667 , n16040 , n17244 );
nor ( n18668 , n18666 , n18667 );
xnor ( n18669 , n18668 , n17191 );
and ( n18670 , n18665 , n18669 );
and ( n18671 , n16401 , n16378 );
and ( n18672 , n16285 , n16376 );
nor ( n18673 , n18671 , n18672 );
xnor ( n18674 , n18673 , n16313 );
and ( n18675 , n18669 , n18674 );
and ( n18676 , n18665 , n18674 );
or ( n18677 , n18670 , n18675 , n18676 );
and ( n18678 , n16008 , n18187 );
and ( n18679 , n16021 , n18184 );
nor ( n18680 , n18678 , n18679 );
xnor ( n18681 , n18680 , n17661 );
and ( n18682 , n18197 , n16053 );
not ( n18683 , n18682 );
and ( n18684 , n18683 , n16063 );
and ( n18685 , n18681 , n18684 );
and ( n18686 , n18677 , n18685 );
and ( n18687 , n18044 , n16055 );
and ( n18688 , n17907 , n16053 );
nor ( n18689 , n18687 , n18688 );
xnor ( n18690 , n18689 , n16063 );
and ( n18691 , n18685 , n18690 );
and ( n18692 , n18677 , n18690 );
or ( n18693 , n18686 , n18691 , n18692 );
xor ( n18694 , n18469 , n18485 );
xor ( n18695 , n18694 , n18502 );
and ( n18696 , n18693 , n18695 );
xor ( n18697 , n18522 , n18538 );
xor ( n18698 , n18697 , n18551 );
and ( n18699 , n18695 , n18698 );
and ( n18700 , n18693 , n18698 );
or ( n18701 , n18696 , n18699 , n18700 );
xor ( n18702 , n18473 , n18477 );
xor ( n18703 , n18702 , n18482 );
xor ( n18704 , n18543 , n18547 );
xor ( n18705 , n18704 , n18371 );
and ( n18706 , n18703 , n18705 );
xor ( n18707 , n18490 , n18494 );
xor ( n18708 , n18707 , n18499 );
and ( n18709 , n18705 , n18708 );
and ( n18710 , n18703 , n18708 );
or ( n18711 , n18706 , n18709 , n18710 );
xor ( n18712 , n18681 , n18684 );
and ( n18713 , n17907 , n16037 );
and ( n18714 , n17688 , n16035 );
nor ( n18715 , n18713 , n18714 );
xnor ( n18716 , n18715 , n16045 );
and ( n18717 , n18712 , n18716 );
and ( n18718 , n18197 , n16055 );
and ( n18719 , n18044 , n16053 );
nor ( n18720 , n18718 , n18719 );
xnor ( n18721 , n18720 , n16063 );
and ( n18722 , n18716 , n18721 );
and ( n18723 , n18712 , n18721 );
or ( n18724 , n18717 , n18722 , n18723 );
xor ( n18725 , n18457 , n18461 );
xor ( n18726 , n18725 , n18466 );
and ( n18727 , n18724 , n18726 );
xor ( n18728 , n18526 , n18530 );
xor ( n18729 , n18728 , n18535 );
and ( n18730 , n18726 , n18729 );
and ( n18731 , n18724 , n18729 );
or ( n18732 , n18727 , n18730 , n18731 );
and ( n18733 , n18711 , n18732 );
xor ( n18734 , n18556 , n18558 );
xor ( n18735 , n18734 , n18561 );
and ( n18736 , n18732 , n18735 );
and ( n18737 , n18711 , n18735 );
or ( n18738 , n18733 , n18736 , n18737 );
and ( n18739 , n18701 , n18738 );
xor ( n18740 , n18505 , n18507 );
xor ( n18741 , n18740 , n18510 );
and ( n18742 , n18738 , n18741 );
and ( n18743 , n18701 , n18741 );
or ( n18744 , n18739 , n18742 , n18743 );
and ( n18745 , n18661 , n18744 );
xor ( n18746 , n18513 , n18515 );
xor ( n18747 , n18746 , n18518 );
and ( n18748 , n18744 , n18747 );
and ( n18749 , n18661 , n18747 );
or ( n18750 , n18745 , n18748 , n18749 );
xor ( n18751 , n18428 , n18430 );
xor ( n18752 , n18751 , n18433 );
and ( n18753 , n18750 , n18752 );
xor ( n18754 , n18521 , n18578 );
xor ( n18755 , n18754 , n18581 );
and ( n18756 , n18752 , n18755 );
and ( n18757 , n18750 , n18755 );
or ( n18758 , n18753 , n18756 , n18757 );
xor ( n18759 , n18584 , n18586 );
xor ( n18760 , n18759 , n18589 );
and ( n18761 , n18758 , n18760 );
xor ( n18762 , n18750 , n18752 );
xor ( n18763 , n18762 , n18755 );
xor ( n18764 , n18554 , n18564 );
xor ( n18765 , n18764 , n18567 );
xor ( n18766 , n18653 , n18655 );
xor ( n18767 , n18766 , n18658 );
and ( n18768 , n18765 , n18767 );
xor ( n18769 , n18701 , n18738 );
xor ( n18770 , n18769 , n18741 );
and ( n18771 , n18767 , n18770 );
and ( n18772 , n18765 , n18770 );
or ( n18773 , n18768 , n18771 , n18772 );
xor ( n18774 , n18570 , n18572 );
xor ( n18775 , n18774 , n18575 );
and ( n18776 , n18773 , n18775 );
xor ( n18777 , n18661 , n18744 );
xor ( n18778 , n18777 , n18747 );
and ( n18779 , n18775 , n18778 );
and ( n18780 , n18773 , n18778 );
or ( n18781 , n18776 , n18779 , n18780 );
and ( n18782 , n18763 , n18781 );
xor ( n18783 , n18773 , n18775 );
xor ( n18784 , n18783 , n18778 );
xor ( n18785 , n18693 , n18695 );
xor ( n18786 , n18785 , n18698 );
xor ( n18787 , n18711 , n18732 );
xor ( n18788 , n18787 , n18735 );
and ( n18789 , n18786 , n18788 );
xor ( n18790 , n18645 , n18647 );
xor ( n18791 , n18790 , n18650 );
xor ( n18792 , n18677 , n18685 );
xor ( n18793 , n18792 , n18690 );
xor ( n18794 , n18597 , n18601 );
xor ( n18795 , n18794 , n18606 );
xor ( n18796 , n18613 , n18617 );
xor ( n18797 , n18796 , n18622 );
and ( n18798 , n18795 , n18797 );
xor ( n18799 , n18630 , n18634 );
xor ( n18800 , n18799 , n18639 );
and ( n18801 , n18797 , n18800 );
and ( n18802 , n18795 , n18800 );
or ( n18803 , n18798 , n18801 , n18802 );
and ( n18804 , n18793 , n18803 );
and ( n18805 , n15974 , n17915 );
and ( n18806 , n16096 , n17913 );
nor ( n18807 , n18805 , n18806 );
xnor ( n18808 , n18807 , n17664 );
and ( n18809 , n16058 , n17246 );
and ( n18810 , n16029 , n17244 );
nor ( n18811 , n18809 , n18810 );
xnor ( n18812 , n18811 , n17191 );
and ( n18813 , n18808 , n18812 );
and ( n18814 , n18812 , n18682 );
and ( n18815 , n18808 , n18682 );
or ( n18816 , n18813 , n18814 , n18815 );
and ( n18817 , n16105 , n18187 );
and ( n18818 , n16008 , n18184 );
nor ( n18819 , n18817 , n18818 );
xnor ( n18820 , n18819 , n17661 );
and ( n18821 , n16910 , n16084 );
and ( n18822 , n16792 , n16082 );
nor ( n18823 , n18821 , n18822 );
xnor ( n18824 , n18823 , n16092 );
and ( n18825 , n18820 , n18824 );
and ( n18826 , n17309 , n16018 );
and ( n18827 , n16995 , n16016 );
nor ( n18828 , n18826 , n18827 );
xnor ( n18829 , n18828 , n16026 );
and ( n18830 , n18824 , n18829 );
and ( n18831 , n18820 , n18829 );
or ( n18832 , n18825 , n18830 , n18831 );
and ( n18833 , n18816 , n18832 );
and ( n18834 , n15995 , n17020 );
and ( n18835 , n16049 , n17018 );
nor ( n18836 , n18834 , n18835 );
xnor ( n18837 , n18836 , n16938 );
and ( n18838 , n16510 , n16378 );
and ( n18839 , n16401 , n16376 );
nor ( n18840 , n18838 , n18839 );
xnor ( n18841 , n18840 , n16313 );
and ( n18842 , n18837 , n18841 );
and ( n18843 , n16668 , n16176 );
and ( n18844 , n16592 , n16174 );
nor ( n18845 , n18843 , n18844 );
xnor ( n18846 , n18845 , n16075 );
and ( n18847 , n18841 , n18846 );
and ( n18848 , n18837 , n18846 );
or ( n18849 , n18842 , n18847 , n18848 );
and ( n18850 , n18832 , n18849 );
and ( n18851 , n18816 , n18849 );
or ( n18852 , n18833 , n18850 , n18851 );
and ( n18853 , n18803 , n18852 );
and ( n18854 , n18793 , n18852 );
or ( n18855 , n18804 , n18853 , n18854 );
and ( n18856 , n18791 , n18855 );
and ( n18857 , n16040 , n17542 );
and ( n18858 , n15961 , n17540 );
nor ( n18859 , n18857 , n18858 );
xnor ( n18860 , n18859 , n17406 );
and ( n18861 , n16285 , n16565 );
and ( n18862 , n16151 , n16563 );
nor ( n18863 , n18861 , n18862 );
xnor ( n18864 , n18863 , n16481 );
and ( n18865 , n18860 , n18864 );
and ( n18866 , n18044 , n16037 );
and ( n18867 , n17907 , n16035 );
nor ( n18868 , n18866 , n18867 );
xnor ( n18869 , n18868 , n16045 );
and ( n18870 , n18864 , n18869 );
and ( n18871 , n18860 , n18869 );
or ( n18872 , n18865 , n18870 , n18871 );
and ( n18873 , n16004 , n16782 );
and ( n18874 , n15982 , n16780 );
nor ( n18875 , n18873 , n18874 );
xnor ( n18876 , n18875 , n16696 );
and ( n18877 , n17610 , n16102 );
and ( n18878 , n17355 , n16100 );
nor ( n18879 , n18877 , n18878 );
xnor ( n18880 , n18879 , n16110 );
and ( n18881 , n18876 , n18880 );
and ( n18882 , n17688 , n15971 );
and ( n18883 , n17720 , n15969 );
nor ( n18884 , n18882 , n18883 );
xnor ( n18885 , n18884 , n15979 );
and ( n18886 , n18880 , n18885 );
and ( n18887 , n18876 , n18885 );
or ( n18888 , n18881 , n18886 , n18887 );
and ( n18889 , n18872 , n18888 );
xor ( n18890 , n18665 , n18669 );
xor ( n18891 , n18890 , n18674 );
and ( n18892 , n18888 , n18891 );
and ( n18893 , n18872 , n18891 );
or ( n18894 , n18889 , n18892 , n18893 );
xor ( n18895 , n18609 , n18625 );
xor ( n18896 , n18895 , n18642 );
and ( n18897 , n18894 , n18896 );
xor ( n18898 , n18724 , n18726 );
xor ( n18899 , n18898 , n18729 );
and ( n18900 , n18896 , n18899 );
and ( n18901 , n18894 , n18899 );
or ( n18902 , n18897 , n18900 , n18901 );
and ( n18903 , n18855 , n18902 );
and ( n18904 , n18791 , n18902 );
or ( n18905 , n18856 , n18903 , n18904 );
and ( n18906 , n18789 , n18905 );
xor ( n18907 , n18765 , n18767 );
xor ( n18908 , n18907 , n18770 );
and ( n18909 , n18905 , n18908 );
and ( n18910 , n18789 , n18908 );
or ( n18911 , n18906 , n18909 , n18910 );
and ( n18912 , n18784 , n18911 );
and ( n18913 , n16049 , n17246 );
and ( n18914 , n16058 , n17244 );
nor ( n18915 , n18913 , n18914 );
xnor ( n18916 , n18915 , n17191 );
and ( n18917 , n16592 , n16378 );
and ( n18918 , n16510 , n16376 );
nor ( n18919 , n18917 , n18918 );
xnor ( n18920 , n18919 , n16313 );
and ( n18921 , n18916 , n18920 );
and ( n18922 , n16792 , n16176 );
and ( n18923 , n16668 , n16174 );
nor ( n18924 , n18922 , n18923 );
xnor ( n18925 , n18924 , n16075 );
and ( n18926 , n18920 , n18925 );
and ( n18927 , n18916 , n18925 );
or ( n18928 , n18921 , n18926 , n18927 );
and ( n18929 , n15982 , n17020 );
and ( n18930 , n15995 , n17018 );
nor ( n18931 , n18929 , n18930 );
xnor ( n18932 , n18931 , n16938 );
and ( n18933 , n16995 , n16084 );
and ( n18934 , n16910 , n16082 );
nor ( n18935 , n18933 , n18934 );
xnor ( n18936 , n18935 , n16092 );
and ( n18937 , n18932 , n18936 );
and ( n18938 , n17355 , n16018 );
and ( n18939 , n17309 , n16016 );
nor ( n18940 , n18938 , n18939 );
xnor ( n18941 , n18940 , n16026 );
and ( n18942 , n18936 , n18941 );
and ( n18943 , n18932 , n18941 );
or ( n18944 , n18937 , n18942 , n18943 );
and ( n18945 , n18928 , n18944 );
and ( n18946 , n15961 , n17915 );
and ( n18947 , n15974 , n17913 );
nor ( n18948 , n18946 , n18947 );
xnor ( n18949 , n18948 , n17664 );
and ( n18950 , n18197 , n16035 );
not ( n18951 , n18950 );
and ( n18952 , n18951 , n16045 );
and ( n18953 , n18949 , n18952 );
and ( n18954 , n18944 , n18953 );
and ( n18955 , n18928 , n18953 );
or ( n18956 , n18945 , n18954 , n18955 );
xor ( n18957 , n18808 , n18812 );
xor ( n18958 , n18957 , n18682 );
xor ( n18959 , n18860 , n18864 );
xor ( n18960 , n18959 , n18869 );
and ( n18961 , n18958 , n18960 );
xor ( n18962 , n18820 , n18824 );
xor ( n18963 , n18962 , n18829 );
and ( n18964 , n18960 , n18963 );
and ( n18965 , n18958 , n18963 );
or ( n18966 , n18961 , n18964 , n18965 );
and ( n18967 , n18956 , n18966 );
xor ( n18968 , n18712 , n18716 );
xor ( n18969 , n18968 , n18721 );
and ( n18970 , n18966 , n18969 );
and ( n18971 , n18956 , n18969 );
or ( n18972 , n18967 , n18970 , n18971 );
xor ( n18973 , n18703 , n18705 );
xor ( n18974 , n18973 , n18708 );
and ( n18975 , n18972 , n18974 );
xor ( n18976 , n18786 , n18788 );
and ( n18977 , n18975 , n18976 );
xor ( n18978 , n18872 , n18888 );
xor ( n18979 , n18978 , n18891 );
and ( n18980 , n16029 , n17542 );
and ( n18981 , n16040 , n17540 );
nor ( n18982 , n18980 , n18981 );
xnor ( n18983 , n18982 , n17406 );
and ( n18984 , n17907 , n15971 );
and ( n18985 , n17688 , n15969 );
nor ( n18986 , n18984 , n18985 );
xnor ( n18987 , n18986 , n15979 );
and ( n18988 , n18983 , n18987 );
and ( n18989 , n18197 , n16037 );
and ( n18990 , n18044 , n16035 );
nor ( n18991 , n18989 , n18990 );
xnor ( n18992 , n18991 , n16045 );
and ( n18993 , n18987 , n18992 );
and ( n18994 , n18983 , n18992 );
or ( n18995 , n18988 , n18993 , n18994 );
and ( n18996 , n16096 , n18187 );
and ( n18997 , n16105 , n18184 );
nor ( n18998 , n18996 , n18997 );
xnor ( n18999 , n18998 , n17661 );
and ( n19000 , n16151 , n16782 );
and ( n19001 , n16004 , n16780 );
nor ( n19002 , n19000 , n19001 );
xnor ( n19003 , n19002 , n16696 );
and ( n19004 , n18999 , n19003 );
and ( n19005 , n17720 , n16102 );
and ( n19006 , n17610 , n16100 );
nor ( n19007 , n19005 , n19006 );
xnor ( n19008 , n19007 , n16110 );
and ( n19009 , n19003 , n19008 );
and ( n19010 , n18999 , n19008 );
or ( n19011 , n19004 , n19009 , n19010 );
and ( n19012 , n18995 , n19011 );
xor ( n19013 , n18837 , n18841 );
xor ( n19014 , n19013 , n18846 );
and ( n19015 , n19011 , n19014 );
and ( n19016 , n18995 , n19014 );
or ( n19017 , n19012 , n19015 , n19016 );
and ( n19018 , n18979 , n19017 );
xor ( n19019 , n18816 , n18832 );
xor ( n19020 , n19019 , n18849 );
and ( n19021 , n19017 , n19020 );
and ( n19022 , n18979 , n19020 );
or ( n19023 , n19018 , n19021 , n19022 );
xor ( n19024 , n18793 , n18803 );
xor ( n19025 , n19024 , n18852 );
and ( n19026 , n19023 , n19025 );
xor ( n19027 , n18894 , n18896 );
xor ( n19028 , n19027 , n18899 );
and ( n19029 , n19025 , n19028 );
and ( n19030 , n19023 , n19028 );
or ( n19031 , n19026 , n19029 , n19030 );
and ( n19032 , n18976 , n19031 );
and ( n19033 , n18975 , n19031 );
or ( n19034 , n18977 , n19032 , n19033 );
xor ( n19035 , n18791 , n18855 );
xor ( n19036 , n19035 , n18902 );
xor ( n19037 , n18972 , n18974 );
and ( n19038 , n15974 , n18187 );
and ( n19039 , n16096 , n18184 );
nor ( n19040 , n19038 , n19039 );
xnor ( n19041 , n19040 , n17661 );
and ( n19042 , n17309 , n16084 );
and ( n19043 , n16995 , n16082 );
nor ( n19044 , n19042 , n19043 );
xnor ( n19045 , n19044 , n16092 );
and ( n19046 , n19041 , n19045 );
and ( n19047 , n17610 , n16018 );
and ( n19048 , n17355 , n16016 );
nor ( n19049 , n19047 , n19048 );
xnor ( n19050 , n19049 , n16026 );
and ( n19051 , n19045 , n19050 );
and ( n19052 , n19041 , n19050 );
or ( n19053 , n19046 , n19051 , n19052 );
and ( n19054 , n16285 , n16782 );
and ( n19055 , n16151 , n16780 );
nor ( n19056 , n19054 , n19055 );
xnor ( n19057 , n19056 , n16696 );
and ( n19058 , n17688 , n16102 );
and ( n19059 , n17720 , n16100 );
nor ( n19060 , n19058 , n19059 );
xnor ( n19061 , n19060 , n16110 );
and ( n19062 , n19057 , n19061 );
and ( n19063 , n18044 , n15971 );
and ( n19064 , n17907 , n15969 );
nor ( n19065 , n19063 , n19064 );
xnor ( n19066 , n19065 , n15979 );
and ( n19067 , n19061 , n19066 );
and ( n19068 , n19057 , n19066 );
or ( n19069 , n19062 , n19067 , n19068 );
and ( n19070 , n19053 , n19069 );
and ( n19071 , n16004 , n17020 );
and ( n19072 , n15982 , n17018 );
nor ( n19073 , n19071 , n19072 );
xnor ( n19074 , n19073 , n16938 );
and ( n19075 , n16668 , n16378 );
and ( n19076 , n16592 , n16376 );
nor ( n19077 , n19075 , n19076 );
xnor ( n19078 , n19077 , n16313 );
and ( n19079 , n19074 , n19078 );
and ( n19080 , n16910 , n16176 );
and ( n19081 , n16792 , n16174 );
nor ( n19082 , n19080 , n19081 );
xnor ( n19083 , n19082 , n16075 );
and ( n19084 , n19078 , n19083 );
and ( n19085 , n19074 , n19083 );
or ( n19086 , n19079 , n19084 , n19085 );
and ( n19087 , n19069 , n19086 );
and ( n19088 , n19053 , n19086 );
or ( n19089 , n19070 , n19087 , n19088 );
xor ( n19090 , n18949 , n18952 );
and ( n19091 , n16040 , n17915 );
and ( n19092 , n15961 , n17913 );
nor ( n19093 , n19091 , n19092 );
xnor ( n19094 , n19093 , n17664 );
and ( n19095 , n15995 , n17246 );
and ( n19096 , n16049 , n17244 );
nor ( n19097 , n19095 , n19096 );
xnor ( n19098 , n19097 , n17191 );
and ( n19099 , n19094 , n19098 );
and ( n19100 , n19098 , n18950 );
and ( n19101 , n19094 , n18950 );
or ( n19102 , n19099 , n19100 , n19101 );
and ( n19103 , n19090 , n19102 );
and ( n19104 , n16401 , n16565 );
and ( n19105 , n16285 , n16563 );
nor ( n19106 , n19104 , n19105 );
xnor ( n19107 , n19106 , n16481 );
and ( n19108 , n19102 , n19107 );
and ( n19109 , n19090 , n19107 );
or ( n19110 , n19103 , n19108 , n19109 );
and ( n19111 , n19089 , n19110 );
xor ( n19112 , n18876 , n18880 );
xor ( n19113 , n19112 , n18885 );
and ( n19114 , n19110 , n19113 );
and ( n19115 , n19089 , n19113 );
or ( n19116 , n19111 , n19114 , n19115 );
xor ( n19117 , n18983 , n18987 );
xor ( n19118 , n19117 , n18992 );
xor ( n19119 , n18999 , n19003 );
xor ( n19120 , n19119 , n19008 );
and ( n19121 , n19118 , n19120 );
xor ( n19122 , n18916 , n18920 );
xor ( n19123 , n19122 , n18925 );
and ( n19124 , n19120 , n19123 );
and ( n19125 , n19118 , n19123 );
or ( n19126 , n19121 , n19124 , n19125 );
xor ( n19127 , n18928 , n18944 );
xor ( n19128 , n19127 , n18953 );
and ( n19129 , n19126 , n19128 );
xor ( n19130 , n18995 , n19011 );
xor ( n19131 , n19130 , n19014 );
and ( n19132 , n19128 , n19131 );
and ( n19133 , n19126 , n19131 );
or ( n19134 , n19129 , n19132 , n19133 );
and ( n19135 , n19116 , n19134 );
xor ( n19136 , n18795 , n18797 );
xor ( n19137 , n19136 , n18800 );
and ( n19138 , n19134 , n19137 );
and ( n19139 , n19116 , n19137 );
or ( n19140 , n19135 , n19138 , n19139 );
and ( n19141 , n19037 , n19140 );
xor ( n19142 , n18956 , n18966 );
xor ( n19143 , n19142 , n18969 );
xor ( n19144 , n18979 , n19017 );
xor ( n19145 , n19144 , n19020 );
and ( n19146 , n19143 , n19145 );
xor ( n19147 , n19116 , n19134 );
xor ( n19148 , n19147 , n19137 );
and ( n19149 , n19145 , n19148 );
and ( n19150 , n19143 , n19148 );
or ( n19151 , n19146 , n19149 , n19150 );
and ( n19152 , n19140 , n19151 );
and ( n19153 , n19037 , n19151 );
or ( n19154 , n19141 , n19152 , n19153 );
and ( n19155 , n19036 , n19154 );
xor ( n19156 , n18975 , n18976 );
xor ( n19157 , n19156 , n19031 );
and ( n19158 , n19154 , n19157 );
and ( n19159 , n19036 , n19157 );
or ( n19160 , n19155 , n19158 , n19159 );
and ( n19161 , n19034 , n19160 );
xor ( n19162 , n18789 , n18905 );
xor ( n19163 , n19162 , n18908 );
and ( n19164 , n19160 , n19163 );
and ( n19165 , n19034 , n19163 );
or ( n19166 , n19161 , n19164 , n19165 );
and ( n19167 , n18911 , n19166 );
and ( n19168 , n18784 , n19166 );
or ( n19169 , n18912 , n19167 , n19168 );
and ( n19170 , n18781 , n19169 );
and ( n19171 , n18763 , n19169 );
or ( n19172 , n18782 , n19170 , n19171 );
and ( n19173 , n18760 , n19172 );
and ( n19174 , n18758 , n19172 );
or ( n19175 , n18761 , n19173 , n19174 );
and ( n19176 , n18592 , n19175 );
and ( n19177 , n18453 , n19175 );
or ( n19178 , n18593 , n19176 , n19177 );
and ( n19179 , n18450 , n19178 );
and ( n19180 , n18288 , n19178 );
or ( n19181 , n18451 , n19179 , n19180 );
and ( n19182 , n18285 , n19181 );
and ( n19183 , n18130 , n19181 );
or ( n19184 , n18286 , n19182 , n19183 );
and ( n19185 , n18127 , n19184 );
and ( n19186 , n17844 , n19184 );
or ( n19187 , n18128 , n19185 , n19186 );
and ( n19188 , n17841 , n19187 );
and ( n19189 , n17755 , n19187 );
or ( n19190 , n17842 , n19188 , n19189 );
and ( n19191 , n17752 , n19190 );
and ( n19192 , n17647 , n19190 );
or ( n19193 , n17753 , n19191 , n19192 );
and ( n19194 , n17644 , n19193 );
and ( n19195 , n17495 , n19193 );
or ( n19196 , n17645 , n19194 , n19195 );
and ( n19197 , n17492 , n19196 );
and ( n19198 , n17344 , n19196 );
or ( n19199 , n17493 , n19197 , n19198 );
and ( n19200 , n17341 , n19199 );
and ( n19201 , n17184 , n19199 );
or ( n19202 , n17342 , n19200 , n19201 );
and ( n19203 , n17181 , n19202 );
and ( n19204 , n17069 , n19202 );
or ( n19205 , n17182 , n19203 , n19204 );
and ( n19206 , n17066 , n19205 );
and ( n19207 , n16848 , n19205 );
or ( n19208 , n17067 , n19206 , n19207 );
and ( n19209 , n16845 , n19208 );
and ( n19210 , n16778 , n19208 );
or ( n19211 , n16846 , n19209 , n19210 );
and ( n19212 , n16775 , n19211 );
and ( n19213 , n16657 , n19211 );
or ( n19214 , n16776 , n19212 , n19213 );
and ( n19215 , n16654 , n19214 );
and ( n19216 , n16545 , n19214 );
or ( n19217 , n16655 , n19215 , n19216 );
and ( n19218 , n16542 , n19217 );
and ( n19219 , n16448 , n19217 );
or ( n19220 , n16543 , n19218 , n19219 );
xor ( n19221 , n16446 , n19220 );
xor ( n19222 , n16448 , n16542 );
xor ( n19223 , n19222 , n19217 );
xor ( n19224 , n16545 , n16654 );
xor ( n19225 , n19224 , n19214 );
xor ( n19226 , n16657 , n16775 );
xor ( n19227 , n19226 , n19211 );
xor ( n19228 , n16778 , n16845 );
xor ( n19229 , n19228 , n19208 );
xor ( n19230 , n16848 , n17066 );
xor ( n19231 , n19230 , n19205 );
xor ( n19232 , n17069 , n17181 );
xor ( n19233 , n19232 , n19202 );
xor ( n19234 , n17184 , n17341 );
xor ( n19235 , n19234 , n19199 );
xor ( n19236 , n17344 , n17492 );
xor ( n19237 , n19236 , n19196 );
xor ( n19238 , n17495 , n17644 );
xor ( n19239 , n19238 , n19193 );
xor ( n19240 , n17647 , n17752 );
xor ( n19241 , n19240 , n19190 );
xor ( n19242 , n17755 , n17841 );
xor ( n19243 , n19242 , n19187 );
xor ( n19244 , n17844 , n18127 );
xor ( n19245 , n19244 , n19184 );
xor ( n19246 , n18130 , n18285 );
xor ( n19247 , n19246 , n19181 );
xor ( n19248 , n18288 , n18450 );
xor ( n19249 , n19248 , n19178 );
xor ( n19250 , n18453 , n18592 );
xor ( n19251 , n19250 , n19175 );
xor ( n19252 , n18758 , n18760 );
xor ( n19253 , n19252 , n19172 );
xor ( n19254 , n18763 , n18781 );
xor ( n19255 , n19254 , n19169 );
xor ( n19256 , n18784 , n18911 );
xor ( n19257 , n19256 , n19166 );
xor ( n19258 , n19034 , n19160 );
xor ( n19259 , n19258 , n19163 );
xor ( n19260 , n19023 , n19025 );
xor ( n19261 , n19260 , n19028 );
and ( n19262 , n15982 , n17246 );
and ( n19263 , n15995 , n17244 );
nor ( n19264 , n19262 , n19263 );
xnor ( n19265 , n19264 , n17191 );
and ( n19266 , n16792 , n16378 );
and ( n19267 , n16668 , n16376 );
nor ( n19268 , n19266 , n19267 );
xnor ( n19269 , n19268 , n16313 );
and ( n19270 , n19265 , n19269 );
and ( n19271 , n16995 , n16176 );
and ( n19272 , n16910 , n16174 );
nor ( n19273 , n19271 , n19272 );
xnor ( n19274 , n19273 , n16075 );
and ( n19275 , n19269 , n19274 );
and ( n19276 , n19265 , n19274 );
or ( n19277 , n19270 , n19275 , n19276 );
and ( n19278 , n15961 , n18187 );
and ( n19279 , n15974 , n18184 );
nor ( n19280 , n19278 , n19279 );
xnor ( n19281 , n19280 , n17661 );
and ( n19282 , n16401 , n16782 );
and ( n19283 , n16285 , n16780 );
nor ( n19284 , n19282 , n19283 );
xnor ( n19285 , n19284 , n16696 );
and ( n19286 , n19281 , n19285 );
and ( n19287 , n17907 , n16102 );
and ( n19288 , n17688 , n16100 );
nor ( n19289 , n19287 , n19288 );
xnor ( n19290 , n19289 , n16110 );
and ( n19291 , n19285 , n19290 );
and ( n19292 , n19281 , n19290 );
or ( n19293 , n19286 , n19291 , n19292 );
and ( n19294 , n19277 , n19293 );
and ( n19295 , n16151 , n17020 );
and ( n19296 , n16004 , n17018 );
nor ( n19297 , n19295 , n19296 );
xnor ( n19298 , n19297 , n16938 );
and ( n19299 , n17355 , n16084 );
and ( n19300 , n17309 , n16082 );
nor ( n19301 , n19299 , n19300 );
xnor ( n19302 , n19301 , n16092 );
and ( n19303 , n19298 , n19302 );
and ( n19304 , n17720 , n16018 );
and ( n19305 , n17610 , n16016 );
nor ( n19306 , n19304 , n19305 );
xnor ( n19307 , n19306 , n16026 );
and ( n19308 , n19302 , n19307 );
and ( n19309 , n19298 , n19307 );
or ( n19310 , n19303 , n19308 , n19309 );
and ( n19311 , n19293 , n19310 );
and ( n19312 , n19277 , n19310 );
or ( n19313 , n19294 , n19311 , n19312 );
and ( n19314 , n16049 , n17542 );
and ( n19315 , n16058 , n17540 );
nor ( n19316 , n19314 , n19315 );
xnor ( n19317 , n19316 , n17406 );
and ( n19318 , n16592 , n16565 );
and ( n19319 , n16510 , n16563 );
nor ( n19320 , n19318 , n19319 );
xnor ( n19321 , n19320 , n16481 );
and ( n19322 , n19317 , n19321 );
and ( n19323 , n18197 , n15971 );
and ( n19324 , n18044 , n15969 );
nor ( n19325 , n19323 , n19324 );
xnor ( n19326 , n19325 , n15979 );
and ( n19327 , n19321 , n19326 );
and ( n19328 , n19317 , n19326 );
or ( n19329 , n19322 , n19327 , n19328 );
xor ( n19330 , n19094 , n19098 );
xor ( n19331 , n19330 , n18950 );
and ( n19332 , n19329 , n19331 );
xor ( n19333 , n19041 , n19045 );
xor ( n19334 , n19333 , n19050 );
and ( n19335 , n19331 , n19334 );
and ( n19336 , n19329 , n19334 );
or ( n19337 , n19332 , n19335 , n19336 );
and ( n19338 , n19313 , n19337 );
xor ( n19339 , n19053 , n19069 );
xor ( n19340 , n19339 , n19086 );
and ( n19341 , n19337 , n19340 );
and ( n19342 , n19313 , n19340 );
or ( n19343 , n19338 , n19341 , n19342 );
and ( n19344 , n16029 , n17915 );
and ( n19345 , n16040 , n17913 );
nor ( n19346 , n19344 , n19345 );
xnor ( n19347 , n19346 , n17664 );
and ( n19348 , n18197 , n15969 );
not ( n19349 , n19348 );
and ( n19350 , n19349 , n15979 );
and ( n19351 , n19347 , n19350 );
and ( n19352 , n16058 , n17542 );
and ( n19353 , n16029 , n17540 );
nor ( n19354 , n19352 , n19353 );
xnor ( n19355 , n19354 , n17406 );
and ( n19356 , n19351 , n19355 );
and ( n19357 , n16510 , n16565 );
and ( n19358 , n16401 , n16563 );
nor ( n19359 , n19357 , n19358 );
xnor ( n19360 , n19359 , n16481 );
and ( n19361 , n19355 , n19360 );
and ( n19362 , n19351 , n19360 );
or ( n19363 , n19356 , n19361 , n19362 );
xor ( n19364 , n18932 , n18936 );
xor ( n19365 , n19364 , n18941 );
and ( n19366 , n19363 , n19365 );
xor ( n19367 , n19090 , n19102 );
xor ( n19368 , n19367 , n19107 );
and ( n19369 , n19365 , n19368 );
and ( n19370 , n19363 , n19368 );
or ( n19371 , n19366 , n19369 , n19370 );
and ( n19372 , n19343 , n19371 );
xor ( n19373 , n18958 , n18960 );
xor ( n19374 , n19373 , n18963 );
and ( n19375 , n19371 , n19374 );
and ( n19376 , n19343 , n19374 );
or ( n19377 , n19372 , n19375 , n19376 );
xor ( n19378 , n19057 , n19061 );
xor ( n19379 , n19378 , n19066 );
xor ( n19380 , n19074 , n19078 );
xor ( n19381 , n19380 , n19083 );
and ( n19382 , n19379 , n19381 );
xor ( n19383 , n19351 , n19355 );
xor ( n19384 , n19383 , n19360 );
and ( n19385 , n19381 , n19384 );
and ( n19386 , n19379 , n19384 );
or ( n19387 , n19382 , n19385 , n19386 );
xor ( n19388 , n19118 , n19120 );
xor ( n19389 , n19388 , n19123 );
and ( n19390 , n19387 , n19389 );
xor ( n19391 , n19363 , n19365 );
xor ( n19392 , n19391 , n19368 );
and ( n19393 , n19389 , n19392 );
and ( n19394 , n19387 , n19392 );
or ( n19395 , n19390 , n19393 , n19394 );
xor ( n19396 , n19089 , n19110 );
xor ( n19397 , n19396 , n19113 );
and ( n19398 , n19395 , n19397 );
xor ( n19399 , n19126 , n19128 );
xor ( n19400 , n19399 , n19131 );
and ( n19401 , n19397 , n19400 );
and ( n19402 , n19395 , n19400 );
or ( n19403 , n19398 , n19401 , n19402 );
and ( n19404 , n19377 , n19403 );
xor ( n19405 , n19143 , n19145 );
xor ( n19406 , n19405 , n19148 );
and ( n19407 , n19403 , n19406 );
and ( n19408 , n19377 , n19406 );
or ( n19409 , n19404 , n19407 , n19408 );
and ( n19410 , n19261 , n19409 );
xor ( n19411 , n19037 , n19140 );
xor ( n19412 , n19411 , n19151 );
and ( n19413 , n19409 , n19412 );
and ( n19414 , n19261 , n19412 );
or ( n19415 , n19410 , n19413 , n19414 );
xor ( n19416 , n19036 , n19154 );
xor ( n19417 , n19416 , n19157 );
and ( n19418 , n19415 , n19417 );
xor ( n19419 , n19415 , n19417 );
xor ( n19420 , n19261 , n19409 );
xor ( n19421 , n19420 , n19412 );
xor ( n19422 , n19347 , n19350 );
and ( n19423 , n16285 , n17020 );
and ( n19424 , n16151 , n17018 );
nor ( n19425 , n19423 , n19424 );
xnor ( n19426 , n19425 , n16938 );
and ( n19427 , n16910 , n16378 );
and ( n19428 , n16792 , n16376 );
nor ( n19429 , n19427 , n19428 );
xnor ( n19430 , n19429 , n16313 );
and ( n19431 , n19426 , n19430 );
and ( n19432 , n17309 , n16176 );
and ( n19433 , n16995 , n16174 );
nor ( n19434 , n19432 , n19433 );
xnor ( n19435 , n19434 , n16075 );
and ( n19436 , n19430 , n19435 );
and ( n19437 , n19426 , n19435 );
or ( n19438 , n19431 , n19436 , n19437 );
and ( n19439 , n19422 , n19438 );
and ( n19440 , n16040 , n18187 );
and ( n19441 , n15961 , n18184 );
nor ( n19442 , n19440 , n19441 );
xnor ( n19443 , n19442 , n17661 );
and ( n19444 , n17610 , n16084 );
and ( n19445 , n17355 , n16082 );
nor ( n19446 , n19444 , n19445 );
xnor ( n19447 , n19446 , n16092 );
and ( n19448 , n19443 , n19447 );
and ( n19449 , n17688 , n16018 );
and ( n19450 , n17720 , n16016 );
nor ( n19451 , n19449 , n19450 );
xnor ( n19452 , n19451 , n16026 );
and ( n19453 , n19447 , n19452 );
and ( n19454 , n19443 , n19452 );
or ( n19455 , n19448 , n19453 , n19454 );
and ( n19456 , n19438 , n19455 );
and ( n19457 , n19422 , n19455 );
or ( n19458 , n19439 , n19456 , n19457 );
xor ( n19459 , n19265 , n19269 );
xor ( n19460 , n19459 , n19274 );
xor ( n19461 , n19281 , n19285 );
xor ( n19462 , n19461 , n19290 );
and ( n19463 , n19460 , n19462 );
xor ( n19464 , n19298 , n19302 );
xor ( n19465 , n19464 , n19307 );
and ( n19466 , n19462 , n19465 );
and ( n19467 , n19460 , n19465 );
or ( n19468 , n19463 , n19466 , n19467 );
and ( n19469 , n19458 , n19468 );
and ( n19470 , n15995 , n17542 );
and ( n19471 , n16049 , n17540 );
nor ( n19472 , n19470 , n19471 );
xnor ( n19473 , n19472 , n17406 );
and ( n19474 , n16510 , n16782 );
and ( n19475 , n16401 , n16780 );
nor ( n19476 , n19474 , n19475 );
xnor ( n19477 , n19476 , n16696 );
and ( n19478 , n19473 , n19477 );
and ( n19479 , n18044 , n16102 );
and ( n19480 , n17907 , n16100 );
nor ( n19481 , n19479 , n19480 );
xnor ( n19482 , n19481 , n16110 );
and ( n19483 , n19477 , n19482 );
and ( n19484 , n19473 , n19482 );
or ( n19485 , n19478 , n19483 , n19484 );
and ( n19486 , n16058 , n17915 );
and ( n19487 , n16029 , n17913 );
nor ( n19488 , n19486 , n19487 );
xnor ( n19489 , n19488 , n17664 );
and ( n19490 , n16004 , n17246 );
and ( n19491 , n15982 , n17244 );
nor ( n19492 , n19490 , n19491 );
xnor ( n19493 , n19492 , n17191 );
and ( n19494 , n19489 , n19493 );
and ( n19495 , n19493 , n19348 );
and ( n19496 , n19489 , n19348 );
or ( n19497 , n19494 , n19495 , n19496 );
and ( n19498 , n19485 , n19497 );
xor ( n19499 , n19317 , n19321 );
xor ( n19500 , n19499 , n19326 );
and ( n19501 , n19497 , n19500 );
and ( n19502 , n19485 , n19500 );
or ( n19503 , n19498 , n19501 , n19502 );
and ( n19504 , n19468 , n19503 );
and ( n19505 , n19458 , n19503 );
or ( n19506 , n19469 , n19504 , n19505 );
xor ( n19507 , n19277 , n19293 );
xor ( n19508 , n19507 , n19310 );
xor ( n19509 , n19329 , n19331 );
xor ( n19510 , n19509 , n19334 );
and ( n19511 , n19508 , n19510 );
xor ( n19512 , n19379 , n19381 );
xor ( n19513 , n19512 , n19384 );
and ( n19514 , n19510 , n19513 );
and ( n19515 , n19508 , n19513 );
or ( n19516 , n19511 , n19514 , n19515 );
and ( n19517 , n19506 , n19516 );
xor ( n19518 , n19313 , n19337 );
xor ( n19519 , n19518 , n19340 );
and ( n19520 , n19516 , n19519 );
and ( n19521 , n19506 , n19519 );
or ( n19522 , n19517 , n19520 , n19521 );
xor ( n19523 , n19343 , n19371 );
xor ( n19524 , n19523 , n19374 );
and ( n19525 , n19522 , n19524 );
xor ( n19526 , n19395 , n19397 );
xor ( n19527 , n19526 , n19400 );
and ( n19528 , n19524 , n19527 );
and ( n19529 , n19522 , n19527 );
or ( n19530 , n19525 , n19528 , n19529 );
xor ( n19531 , n19377 , n19403 );
xor ( n19532 , n19531 , n19406 );
and ( n19533 , n19530 , n19532 );
xor ( n19534 , n19522 , n19524 );
xor ( n19535 , n19534 , n19527 );
and ( n19536 , n16029 , n18187 );
and ( n19537 , n16040 , n18184 );
nor ( n19538 , n19536 , n19537 );
xnor ( n19539 , n19538 , n17661 );
and ( n19540 , n15982 , n17542 );
and ( n19541 , n15995 , n17540 );
nor ( n19542 , n19540 , n19541 );
xnor ( n19543 , n19542 , n17406 );
and ( n19544 , n19539 , n19543 );
and ( n19545 , n18197 , n16102 );
and ( n19546 , n18044 , n16100 );
nor ( n19547 , n19545 , n19546 );
xnor ( n19548 , n19547 , n16110 );
and ( n19549 , n19543 , n19548 );
and ( n19550 , n19539 , n19548 );
or ( n19551 , n19544 , n19549 , n19550 );
and ( n19552 , n16151 , n17246 );
and ( n19553 , n16004 , n17244 );
nor ( n19554 , n19552 , n19553 );
xnor ( n19555 , n19554 , n17191 );
and ( n19556 , n16995 , n16378 );
and ( n19557 , n16910 , n16376 );
nor ( n19558 , n19556 , n19557 );
xnor ( n19559 , n19558 , n16313 );
and ( n19560 , n19555 , n19559 );
and ( n19561 , n17355 , n16176 );
and ( n19562 , n17309 , n16174 );
nor ( n19563 , n19561 , n19562 );
xnor ( n19564 , n19563 , n16075 );
and ( n19565 , n19559 , n19564 );
and ( n19566 , n19555 , n19564 );
or ( n19567 , n19560 , n19565 , n19566 );
and ( n19568 , n19551 , n19567 );
xor ( n19569 , n19473 , n19477 );
xor ( n19570 , n19569 , n19482 );
and ( n19571 , n19567 , n19570 );
and ( n19572 , n19551 , n19570 );
or ( n19573 , n19568 , n19571 , n19572 );
xor ( n19574 , n19422 , n19438 );
xor ( n19575 , n19574 , n19455 );
and ( n19576 , n19573 , n19575 );
xor ( n19577 , n19460 , n19462 );
xor ( n19578 , n19577 , n19465 );
and ( n19579 , n19575 , n19578 );
and ( n19580 , n19573 , n19578 );
or ( n19581 , n19576 , n19579 , n19580 );
and ( n19582 , n16401 , n17020 );
and ( n19583 , n16285 , n17018 );
nor ( n19584 , n19582 , n19583 );
xnor ( n19585 , n19584 , n16938 );
and ( n19586 , n17720 , n16084 );
and ( n19587 , n17610 , n16082 );
nor ( n19588 , n19586 , n19587 );
xnor ( n19589 , n19588 , n16092 );
and ( n19590 , n19585 , n19589 );
and ( n19591 , n17907 , n16018 );
and ( n19592 , n17688 , n16016 );
nor ( n19593 , n19591 , n19592 );
xnor ( n19594 , n19593 , n16026 );
and ( n19595 , n19589 , n19594 );
and ( n19596 , n19585 , n19594 );
or ( n19597 , n19590 , n19595 , n19596 );
and ( n19598 , n16049 , n17915 );
and ( n19599 , n16058 , n17913 );
nor ( n19600 , n19598 , n19599 );
xnor ( n19601 , n19600 , n17664 );
and ( n19602 , n18197 , n16100 );
not ( n19603 , n19602 );
and ( n19604 , n19603 , n16110 );
and ( n19605 , n19601 , n19604 );
and ( n19606 , n19597 , n19605 );
and ( n19607 , n16668 , n16565 );
and ( n19608 , n16592 , n16563 );
nor ( n19609 , n19607 , n19608 );
xnor ( n19610 , n19609 , n16481 );
and ( n19611 , n19605 , n19610 );
and ( n19612 , n19597 , n19610 );
or ( n19613 , n19606 , n19611 , n19612 );
xor ( n19614 , n19489 , n19493 );
xor ( n19615 , n19614 , n19348 );
xor ( n19616 , n19426 , n19430 );
xor ( n19617 , n19616 , n19435 );
and ( n19618 , n19615 , n19617 );
xor ( n19619 , n19443 , n19447 );
xor ( n19620 , n19619 , n19452 );
and ( n19621 , n19617 , n19620 );
and ( n19622 , n19615 , n19620 );
or ( n19623 , n19618 , n19621 , n19622 );
and ( n19624 , n19613 , n19623 );
xor ( n19625 , n19485 , n19497 );
xor ( n19626 , n19625 , n19500 );
and ( n19627 , n19623 , n19626 );
and ( n19628 , n19613 , n19626 );
or ( n19629 , n19624 , n19627 , n19628 );
and ( n19630 , n19581 , n19629 );
xor ( n19631 , n19458 , n19468 );
xor ( n19632 , n19631 , n19503 );
and ( n19633 , n19629 , n19632 );
and ( n19634 , n19581 , n19632 );
or ( n19635 , n19630 , n19633 , n19634 );
xor ( n19636 , n19387 , n19389 );
xor ( n19637 , n19636 , n19392 );
and ( n19638 , n19635 , n19637 );
xor ( n19639 , n19506 , n19516 );
xor ( n19640 , n19639 , n19519 );
and ( n19641 , n19637 , n19640 );
and ( n19642 , n19635 , n19640 );
or ( n19643 , n19638 , n19641 , n19642 );
and ( n19644 , n19535 , n19643 );
and ( n19645 , n16004 , n17542 );
and ( n19646 , n15982 , n17540 );
nor ( n19647 , n19645 , n19646 );
xnor ( n19648 , n19647 , n17406 );
and ( n19649 , n16668 , n16782 );
and ( n19650 , n16592 , n16780 );
nor ( n19651 , n19649 , n19650 );
xnor ( n19652 , n19651 , n16696 );
and ( n19653 , n19648 , n19652 );
and ( n19654 , n16910 , n16565 );
and ( n19655 , n16792 , n16563 );
nor ( n19656 , n19654 , n19655 );
xnor ( n19657 , n19656 , n16481 );
and ( n19658 , n19652 , n19657 );
and ( n19659 , n19648 , n19657 );
or ( n19660 , n19653 , n19658 , n19659 );
and ( n19661 , n15995 , n17915 );
and ( n19662 , n16049 , n17913 );
nor ( n19663 , n19661 , n19662 );
xnor ( n19664 , n19663 , n17664 );
and ( n19665 , n16285 , n17246 );
and ( n19666 , n16151 , n17244 );
nor ( n19667 , n19665 , n19666 );
xnor ( n19668 , n19667 , n17191 );
and ( n19669 , n19664 , n19668 );
and ( n19670 , n19668 , n19602 );
and ( n19671 , n19664 , n19602 );
or ( n19672 , n19669 , n19670 , n19671 );
and ( n19673 , n19660 , n19672 );
and ( n19674 , n16058 , n18187 );
and ( n19675 , n16029 , n18184 );
nor ( n19676 , n19674 , n19675 );
xnor ( n19677 , n19676 , n17661 );
and ( n19678 , n17688 , n16084 );
and ( n19679 , n17720 , n16082 );
nor ( n19680 , n19678 , n19679 );
xnor ( n19681 , n19680 , n16092 );
and ( n19682 , n19677 , n19681 );
and ( n19683 , n18044 , n16018 );
and ( n19684 , n17907 , n16016 );
nor ( n19685 , n19683 , n19684 );
xnor ( n19686 , n19685 , n16026 );
and ( n19687 , n19681 , n19686 );
and ( n19688 , n19677 , n19686 );
or ( n19689 , n19682 , n19687 , n19688 );
and ( n19690 , n19672 , n19689 );
and ( n19691 , n19660 , n19689 );
or ( n19692 , n19673 , n19690 , n19691 );
xor ( n19693 , n19601 , n19604 );
and ( n19694 , n16592 , n16782 );
and ( n19695 , n16510 , n16780 );
nor ( n19696 , n19694 , n19695 );
xnor ( n19697 , n19696 , n16696 );
and ( n19698 , n19693 , n19697 );
and ( n19699 , n16792 , n16565 );
and ( n19700 , n16668 , n16563 );
nor ( n19701 , n19699 , n19700 );
xnor ( n19702 , n19701 , n16481 );
and ( n19703 , n19697 , n19702 );
and ( n19704 , n19693 , n19702 );
or ( n19705 , n19698 , n19703 , n19704 );
and ( n19706 , n19692 , n19705 );
xor ( n19707 , n19597 , n19605 );
xor ( n19708 , n19707 , n19610 );
and ( n19709 , n19705 , n19708 );
and ( n19710 , n19692 , n19708 );
or ( n19711 , n19706 , n19709 , n19710 );
and ( n19712 , n16510 , n17020 );
and ( n19713 , n16401 , n17018 );
nor ( n19714 , n19712 , n19713 );
xnor ( n19715 , n19714 , n16938 );
and ( n19716 , n17309 , n16378 );
and ( n19717 , n16995 , n16376 );
nor ( n19718 , n19716 , n19717 );
xnor ( n19719 , n19718 , n16313 );
and ( n19720 , n19715 , n19719 );
and ( n19721 , n17610 , n16176 );
and ( n19722 , n17355 , n16174 );
nor ( n19723 , n19721 , n19722 );
xnor ( n19724 , n19723 , n16075 );
and ( n19725 , n19719 , n19724 );
and ( n19726 , n19715 , n19724 );
or ( n19727 , n19720 , n19725 , n19726 );
xor ( n19728 , n19539 , n19543 );
xor ( n19729 , n19728 , n19548 );
and ( n19730 , n19727 , n19729 );
xor ( n19731 , n19585 , n19589 );
xor ( n19732 , n19731 , n19594 );
and ( n19733 , n19729 , n19732 );
and ( n19734 , n19727 , n19732 );
or ( n19735 , n19730 , n19733 , n19734 );
xor ( n19736 , n19615 , n19617 );
xor ( n19737 , n19736 , n19620 );
and ( n19738 , n19735 , n19737 );
xor ( n19739 , n19551 , n19567 );
xor ( n19740 , n19739 , n19570 );
and ( n19741 , n19737 , n19740 );
and ( n19742 , n19735 , n19740 );
or ( n19743 , n19738 , n19741 , n19742 );
and ( n19744 , n19711 , n19743 );
xor ( n19745 , n19613 , n19623 );
xor ( n19746 , n19745 , n19626 );
and ( n19747 , n19743 , n19746 );
and ( n19748 , n19711 , n19746 );
or ( n19749 , n19744 , n19747 , n19748 );
xor ( n19750 , n19581 , n19629 );
xor ( n19751 , n19750 , n19632 );
and ( n19752 , n19749 , n19751 );
xor ( n19753 , n19508 , n19510 );
xor ( n19754 , n19753 , n19513 );
and ( n19755 , n19751 , n19754 );
and ( n19756 , n19749 , n19754 );
or ( n19757 , n19752 , n19755 , n19756 );
xor ( n19758 , n19635 , n19637 );
xor ( n19759 , n19758 , n19640 );
and ( n19760 , n19757 , n19759 );
xor ( n19761 , n19749 , n19751 );
xor ( n19762 , n19761 , n19754 );
xor ( n19763 , n19573 , n19575 );
xor ( n19764 , n19763 , n19578 );
xor ( n19765 , n19711 , n19743 );
xor ( n19766 , n19765 , n19746 );
and ( n19767 , n19764 , n19766 );
and ( n19768 , n16049 , n18187 );
and ( n19769 , n16058 , n18184 );
nor ( n19770 , n19768 , n19769 );
xnor ( n19771 , n19770 , n17661 );
and ( n19772 , n16151 , n17542 );
and ( n19773 , n16004 , n17540 );
nor ( n19774 , n19772 , n19773 );
xnor ( n19775 , n19774 , n17406 );
and ( n19776 , n19771 , n19775 );
and ( n19777 , n16792 , n16782 );
and ( n19778 , n16668 , n16780 );
nor ( n19779 , n19777 , n19778 );
xnor ( n19780 , n19779 , n16696 );
and ( n19781 , n19775 , n19780 );
and ( n19782 , n19771 , n19780 );
or ( n19783 , n19776 , n19781 , n19782 );
and ( n19784 , n16592 , n17020 );
and ( n19785 , n16510 , n17018 );
nor ( n19786 , n19784 , n19785 );
xnor ( n19787 , n19786 , n16938 );
and ( n19788 , n17907 , n16084 );
and ( n19789 , n17688 , n16082 );
nor ( n19790 , n19788 , n19789 );
xnor ( n19791 , n19790 , n16092 );
and ( n19792 , n19787 , n19791 );
and ( n19793 , n18197 , n16018 );
and ( n19794 , n18044 , n16016 );
nor ( n19795 , n19793 , n19794 );
xnor ( n19796 , n19795 , n16026 );
and ( n19797 , n19791 , n19796 );
and ( n19798 , n19787 , n19796 );
or ( n19799 , n19792 , n19797 , n19798 );
and ( n19800 , n19783 , n19799 );
and ( n19801 , n15982 , n17915 );
and ( n19802 , n15995 , n17913 );
nor ( n19803 , n19801 , n19802 );
xnor ( n19804 , n19803 , n17664 );
and ( n19805 , n18197 , n16016 );
not ( n19806 , n19805 );
and ( n19807 , n19806 , n16026 );
and ( n19808 , n19804 , n19807 );
and ( n19809 , n19799 , n19808 );
and ( n19810 , n19783 , n19808 );
or ( n19811 , n19800 , n19809 , n19810 );
xor ( n19812 , n19555 , n19559 );
xor ( n19813 , n19812 , n19564 );
and ( n19814 , n19811 , n19813 );
xor ( n19815 , n19693 , n19697 );
xor ( n19816 , n19815 , n19702 );
and ( n19817 , n19813 , n19816 );
and ( n19818 , n19811 , n19816 );
or ( n19819 , n19814 , n19817 , n19818 );
xor ( n19820 , n19692 , n19705 );
xor ( n19821 , n19820 , n19708 );
and ( n19822 , n19819 , n19821 );
and ( n19823 , n19766 , n19822 );
and ( n19824 , n19764 , n19822 );
or ( n19825 , n19767 , n19823 , n19824 );
and ( n19826 , n19762 , n19825 );
xor ( n19827 , n19735 , n19737 );
xor ( n19828 , n19827 , n19740 );
and ( n19829 , n16401 , n17246 );
and ( n19830 , n16285 , n17244 );
nor ( n19831 , n19829 , n19830 );
xnor ( n19832 , n19831 , n17191 );
and ( n19833 , n17355 , n16378 );
and ( n19834 , n17309 , n16376 );
nor ( n19835 , n19833 , n19834 );
xnor ( n19836 , n19835 , n16313 );
and ( n19837 , n19832 , n19836 );
and ( n19838 , n17720 , n16176 );
and ( n19839 , n17610 , n16174 );
nor ( n19840 , n19838 , n19839 );
xnor ( n19841 , n19840 , n16075 );
and ( n19842 , n19836 , n19841 );
and ( n19843 , n19832 , n19841 );
or ( n19844 , n19837 , n19842 , n19843 );
xor ( n19845 , n19715 , n19719 );
xor ( n19846 , n19845 , n19724 );
and ( n19847 , n19844 , n19846 );
xor ( n19848 , n19648 , n19652 );
xor ( n19849 , n19848 , n19657 );
and ( n19850 , n19846 , n19849 );
and ( n19851 , n19844 , n19849 );
or ( n19852 , n19847 , n19850 , n19851 );
xor ( n19853 , n19660 , n19672 );
xor ( n19854 , n19853 , n19689 );
and ( n19855 , n19852 , n19854 );
and ( n19856 , n19828 , n19855 );
xor ( n19857 , n19819 , n19821 );
and ( n19858 , n19855 , n19857 );
and ( n19859 , n19828 , n19857 );
or ( n19860 , n19856 , n19858 , n19859 );
xor ( n19861 , n19764 , n19766 );
xor ( n19862 , n19861 , n19822 );
and ( n19863 , n19860 , n19862 );
xor ( n19864 , n19804 , n19807 );
and ( n19865 , n16004 , n17915 );
and ( n19866 , n15982 , n17913 );
nor ( n19867 , n19865 , n19866 );
xnor ( n19868 , n19867 , n17664 );
and ( n19869 , n17610 , n16378 );
and ( n19870 , n17355 , n16376 );
nor ( n19871 , n19869 , n19870 );
xnor ( n19872 , n19871 , n16313 );
and ( n19873 , n19868 , n19872 );
and ( n19874 , n17688 , n16176 );
and ( n19875 , n17720 , n16174 );
nor ( n19876 , n19874 , n19875 );
xnor ( n19877 , n19876 , n16075 );
and ( n19878 , n19872 , n19877 );
and ( n19879 , n19868 , n19877 );
or ( n19880 , n19873 , n19878 , n19879 );
and ( n19881 , n19864 , n19880 );
and ( n19882 , n16995 , n16565 );
and ( n19883 , n16910 , n16563 );
nor ( n19884 , n19882 , n19883 );
xnor ( n19885 , n19884 , n16481 );
and ( n19886 , n19880 , n19885 );
and ( n19887 , n19864 , n19885 );
or ( n19888 , n19881 , n19886 , n19887 );
xor ( n19889 , n19664 , n19668 );
xor ( n19890 , n19889 , n19602 );
and ( n19891 , n19888 , n19890 );
xor ( n19892 , n19677 , n19681 );
xor ( n19893 , n19892 , n19686 );
and ( n19894 , n19890 , n19893 );
and ( n19895 , n19888 , n19893 );
or ( n19896 , n19891 , n19894 , n19895 );
xor ( n19897 , n19811 , n19813 );
xor ( n19898 , n19897 , n19816 );
and ( n19899 , n19896 , n19898 );
and ( n19900 , n15995 , n18187 );
and ( n19901 , n16049 , n18184 );
nor ( n19902 , n19900 , n19901 );
xnor ( n19903 , n19902 , n17661 );
and ( n19904 , n16510 , n17246 );
and ( n19905 , n16401 , n17244 );
nor ( n19906 , n19904 , n19905 );
xnor ( n19907 , n19906 , n17191 );
and ( n19908 , n19903 , n19907 );
and ( n19909 , n19907 , n19805 );
and ( n19910 , n19903 , n19805 );
or ( n19911 , n19908 , n19909 , n19910 );
and ( n19912 , n16285 , n17542 );
and ( n19913 , n16151 , n17540 );
nor ( n19914 , n19912 , n19913 );
xnor ( n19915 , n19914 , n17406 );
and ( n19916 , n16668 , n17020 );
and ( n19917 , n16592 , n17018 );
nor ( n19918 , n19916 , n19917 );
xnor ( n19919 , n19918 , n16938 );
and ( n19920 , n19915 , n19919 );
and ( n19921 , n18044 , n16084 );
and ( n19922 , n17907 , n16082 );
nor ( n19923 , n19921 , n19922 );
xnor ( n19924 , n19923 , n16092 );
and ( n19925 , n19919 , n19924 );
and ( n19926 , n19915 , n19924 );
or ( n19927 , n19920 , n19925 , n19926 );
and ( n19928 , n19911 , n19927 );
xor ( n19929 , n19771 , n19775 );
xor ( n19930 , n19929 , n19780 );
and ( n19931 , n19927 , n19930 );
and ( n19932 , n19911 , n19930 );
or ( n19933 , n19928 , n19931 , n19932 );
and ( n19934 , n15982 , n18187 );
and ( n19935 , n15995 , n18184 );
nor ( n19936 , n19934 , n19935 );
xnor ( n19937 , n19936 , n17661 );
and ( n19938 , n18197 , n16082 );
not ( n19939 , n19938 );
and ( n19940 , n19939 , n16092 );
and ( n19941 , n19937 , n19940 );
and ( n19942 , n16910 , n16782 );
and ( n19943 , n16792 , n16780 );
nor ( n19944 , n19942 , n19943 );
xnor ( n19945 , n19944 , n16696 );
and ( n19946 , n19941 , n19945 );
and ( n19947 , n17309 , n16565 );
and ( n19948 , n16995 , n16563 );
nor ( n19949 , n19947 , n19948 );
xnor ( n19950 , n19949 , n16481 );
and ( n19951 , n19945 , n19950 );
and ( n19952 , n19941 , n19950 );
or ( n19953 , n19946 , n19951 , n19952 );
xor ( n19954 , n19787 , n19791 );
xor ( n19955 , n19954 , n19796 );
and ( n19956 , n19953 , n19955 );
xor ( n19957 , n19832 , n19836 );
xor ( n19958 , n19957 , n19841 );
and ( n19959 , n19955 , n19958 );
and ( n19960 , n19953 , n19958 );
or ( n19961 , n19956 , n19959 , n19960 );
and ( n19962 , n19933 , n19961 );
xor ( n19963 , n19783 , n19799 );
xor ( n19964 , n19963 , n19808 );
and ( n19965 , n19961 , n19964 );
and ( n19966 , n19933 , n19964 );
or ( n19967 , n19962 , n19965 , n19966 );
and ( n19968 , n16151 , n17915 );
and ( n19969 , n16004 , n17913 );
nor ( n19970 , n19968 , n19969 );
xnor ( n19971 , n19970 , n17664 );
and ( n19972 , n16792 , n17020 );
and ( n19973 , n16668 , n17018 );
nor ( n19974 , n19972 , n19973 );
xnor ( n19975 , n19974 , n16938 );
and ( n19976 , n19971 , n19975 );
and ( n19977 , n18197 , n16084 );
and ( n19978 , n18044 , n16082 );
nor ( n19979 , n19977 , n19978 );
xnor ( n19980 , n19979 , n16092 );
and ( n19981 , n19975 , n19980 );
and ( n19982 , n19971 , n19980 );
or ( n19983 , n19976 , n19981 , n19982 );
and ( n19984 , n16592 , n17246 );
and ( n19985 , n16510 , n17244 );
nor ( n19986 , n19984 , n19985 );
xnor ( n19987 , n19986 , n17191 );
and ( n19988 , n17720 , n16378 );
and ( n19989 , n17610 , n16376 );
nor ( n19990 , n19988 , n19989 );
xnor ( n19991 , n19990 , n16313 );
and ( n19992 , n19987 , n19991 );
and ( n19993 , n17907 , n16176 );
and ( n19994 , n17688 , n16174 );
nor ( n19995 , n19993 , n19994 );
xnor ( n19996 , n19995 , n16075 );
and ( n19997 , n19991 , n19996 );
and ( n19998 , n19987 , n19996 );
or ( n19999 , n19992 , n19997 , n19998 );
and ( n20000 , n19983 , n19999 );
and ( n20001 , n16401 , n17542 );
and ( n20002 , n16285 , n17540 );
nor ( n20003 , n20001 , n20002 );
xnor ( n20004 , n20003 , n17406 );
and ( n20005 , n16995 , n16782 );
and ( n20006 , n16910 , n16780 );
nor ( n20007 , n20005 , n20006 );
xnor ( n20008 , n20007 , n16696 );
and ( n20009 , n20004 , n20008 );
and ( n20010 , n17355 , n16565 );
and ( n20011 , n17309 , n16563 );
nor ( n20012 , n20010 , n20011 );
xnor ( n20013 , n20012 , n16481 );
and ( n20014 , n20008 , n20013 );
and ( n20015 , n20004 , n20013 );
or ( n20016 , n20009 , n20014 , n20015 );
and ( n20017 , n19999 , n20016 );
and ( n20018 , n19983 , n20016 );
or ( n20019 , n20000 , n20017 , n20018 );
xor ( n20020 , n19864 , n19880 );
xor ( n20021 , n20020 , n19885 );
and ( n20022 , n20019 , n20021 );
xor ( n20023 , n19911 , n19927 );
xor ( n20024 , n20023 , n19930 );
and ( n20025 , n20021 , n20024 );
and ( n20026 , n20019 , n20024 );
or ( n20027 , n20022 , n20025 , n20026 );
xor ( n20028 , n19844 , n19846 );
xor ( n20029 , n20028 , n19849 );
and ( n20030 , n20027 , n20029 );
xor ( n20031 , n19888 , n19890 );
xor ( n20032 , n20031 , n19893 );
and ( n20033 , n20029 , n20032 );
and ( n20034 , n20027 , n20032 );
or ( n20035 , n20030 , n20033 , n20034 );
and ( n20036 , n19967 , n20035 );
and ( n20037 , n19899 , n20036 );
xor ( n20038 , n19727 , n19729 );
xor ( n20039 , n20038 , n19732 );
xor ( n20040 , n19852 , n19854 );
and ( n20041 , n20039 , n20040 );
xor ( n20042 , n19896 , n19898 );
and ( n20043 , n20040 , n20042 );
and ( n20044 , n20039 , n20042 );
or ( n20045 , n20041 , n20043 , n20044 );
and ( n20046 , n20036 , n20045 );
and ( n20047 , n19899 , n20045 );
or ( n20048 , n20037 , n20046 , n20047 );
and ( n20049 , n19862 , n20048 );
and ( n20050 , n19860 , n20048 );
or ( n20051 , n19863 , n20049 , n20050 );
and ( n20052 , n19825 , n20051 );
and ( n20053 , n19762 , n20051 );
or ( n20054 , n19826 , n20052 , n20053 );
and ( n20055 , n19759 , n20054 );
and ( n20056 , n19757 , n20054 );
or ( n20057 , n19760 , n20055 , n20056 );
and ( n20058 , n19643 , n20057 );
and ( n20059 , n19535 , n20057 );
or ( n20060 , n19644 , n20058 , n20059 );
and ( n20061 , n19532 , n20060 );
and ( n20062 , n19530 , n20060 );
or ( n20063 , n19533 , n20061 , n20062 );
and ( n20064 , n19421 , n20063 );
xor ( n20065 , n19421 , n20063 );
xor ( n20066 , n19530 , n19532 );
xor ( n20067 , n20066 , n20060 );
xor ( n20068 , n19535 , n19643 );
xor ( n20069 , n20068 , n20057 );
xor ( n20070 , n19757 , n19759 );
xor ( n20071 , n20070 , n20054 );
xor ( n20072 , n19762 , n19825 );
xor ( n20073 , n20072 , n20051 );
xor ( n20074 , n19828 , n19855 );
xor ( n20075 , n20074 , n19857 );
xor ( n20076 , n19967 , n20035 );
xor ( n20077 , n19903 , n19907 );
xor ( n20078 , n20077 , n19805 );
xor ( n20079 , n19915 , n19919 );
xor ( n20080 , n20079 , n19924 );
and ( n20081 , n20078 , n20080 );
xor ( n20082 , n19868 , n19872 );
xor ( n20083 , n20082 , n19877 );
and ( n20084 , n20080 , n20083 );
and ( n20085 , n20078 , n20083 );
or ( n20086 , n20081 , n20084 , n20085 );
xor ( n20087 , n19953 , n19955 );
xor ( n20088 , n20087 , n19958 );
and ( n20089 , n20086 , n20088 );
xor ( n20090 , n20019 , n20021 );
xor ( n20091 , n20090 , n20024 );
and ( n20092 , n20088 , n20091 );
and ( n20093 , n20086 , n20091 );
or ( n20094 , n20089 , n20092 , n20093 );
xor ( n20095 , n19933 , n19961 );
xor ( n20096 , n20095 , n19964 );
and ( n20097 , n20094 , n20096 );
xor ( n20098 , n20027 , n20029 );
xor ( n20099 , n20098 , n20032 );
and ( n20100 , n20096 , n20099 );
and ( n20101 , n20094 , n20099 );
or ( n20102 , n20097 , n20100 , n20101 );
and ( n20103 , n20076 , n20102 );
xor ( n20104 , n20039 , n20040 );
xor ( n20105 , n20104 , n20042 );
and ( n20106 , n20102 , n20105 );
and ( n20107 , n20076 , n20105 );
or ( n20108 , n20103 , n20106 , n20107 );
and ( n20109 , n20075 , n20108 );
xor ( n20110 , n19899 , n20036 );
xor ( n20111 , n20110 , n20045 );
and ( n20112 , n20108 , n20111 );
and ( n20113 , n20075 , n20111 );
or ( n20114 , n20109 , n20112 , n20113 );
xor ( n20115 , n19860 , n19862 );
xor ( n20116 , n20115 , n20048 );
and ( n20117 , n20114 , n20116 );
xor ( n20118 , n20114 , n20116 );
xor ( n20119 , n20075 , n20108 );
xor ( n20120 , n20119 , n20111 );
xor ( n20121 , n20076 , n20102 );
xor ( n20122 , n20121 , n20105 );
xor ( n20123 , n20094 , n20096 );
xor ( n20124 , n20123 , n20099 );
xor ( n20125 , n19937 , n19940 );
and ( n20126 , n16004 , n18187 );
and ( n20127 , n15982 , n18184 );
nor ( n20128 , n20126 , n20127 );
xnor ( n20129 , n20128 , n17661 );
and ( n20130 , n16668 , n17246 );
and ( n20131 , n16592 , n17244 );
nor ( n20132 , n20130 , n20131 );
xnor ( n20133 , n20132 , n17191 );
and ( n20134 , n20129 , n20133 );
and ( n20135 , n20133 , n19938 );
and ( n20136 , n20129 , n19938 );
or ( n20137 , n20134 , n20135 , n20136 );
and ( n20138 , n20125 , n20137 );
and ( n20139 , n16285 , n17915 );
and ( n20140 , n16151 , n17913 );
nor ( n20141 , n20139 , n20140 );
xnor ( n20142 , n20141 , n17664 );
and ( n20143 , n17688 , n16378 );
and ( n20144 , n17720 , n16376 );
nor ( n20145 , n20143 , n20144 );
xnor ( n20146 , n20145 , n16313 );
and ( n20147 , n20142 , n20146 );
and ( n20148 , n18044 , n16176 );
and ( n20149 , n17907 , n16174 );
nor ( n20150 , n20148 , n20149 );
xnor ( n20151 , n20150 , n16075 );
and ( n20152 , n20146 , n20151 );
and ( n20153 , n20142 , n20151 );
or ( n20154 , n20147 , n20152 , n20153 );
and ( n20155 , n20137 , n20154 );
and ( n20156 , n20125 , n20154 );
or ( n20157 , n20138 , n20155 , n20156 );
and ( n20158 , n16510 , n17542 );
and ( n20159 , n16401 , n17540 );
nor ( n20160 , n20158 , n20159 );
xnor ( n20161 , n20160 , n17406 );
and ( n20162 , n16910 , n17020 );
and ( n20163 , n16792 , n17018 );
nor ( n20164 , n20162 , n20163 );
xnor ( n20165 , n20164 , n16938 );
and ( n20166 , n20161 , n20165 );
and ( n20167 , n17309 , n16782 );
and ( n20168 , n16995 , n16780 );
nor ( n20169 , n20167 , n20168 );
xnor ( n20170 , n20169 , n16696 );
and ( n20171 , n20165 , n20170 );
and ( n20172 , n20161 , n20170 );
or ( n20173 , n20166 , n20171 , n20172 );
xor ( n20174 , n19987 , n19991 );
xor ( n20175 , n20174 , n19996 );
and ( n20176 , n20173 , n20175 );
xor ( n20177 , n20004 , n20008 );
xor ( n20178 , n20177 , n20013 );
and ( n20179 , n20175 , n20178 );
and ( n20180 , n20173 , n20178 );
or ( n20181 , n20176 , n20179 , n20180 );
and ( n20182 , n20157 , n20181 );
xor ( n20183 , n19941 , n19945 );
xor ( n20184 , n20183 , n19950 );
and ( n20185 , n20181 , n20184 );
and ( n20186 , n20157 , n20184 );
or ( n20187 , n20182 , n20185 , n20186 );
xor ( n20188 , n19983 , n19999 );
xor ( n20189 , n20188 , n20016 );
xor ( n20190 , n20078 , n20080 );
xor ( n20191 , n20190 , n20083 );
and ( n20192 , n20189 , n20191 );
xor ( n20193 , n20157 , n20181 );
xor ( n20194 , n20193 , n20184 );
and ( n20195 , n20191 , n20194 );
and ( n20196 , n20189 , n20194 );
or ( n20197 , n20192 , n20195 , n20196 );
and ( n20198 , n20187 , n20197 );
xor ( n20199 , n20086 , n20088 );
xor ( n20200 , n20199 , n20091 );
and ( n20201 , n20197 , n20200 );
and ( n20202 , n20187 , n20200 );
or ( n20203 , n20198 , n20201 , n20202 );
and ( n20204 , n20124 , n20203 );
xor ( n20205 , n20187 , n20197 );
xor ( n20206 , n20205 , n20200 );
and ( n20207 , n16792 , n17246 );
and ( n20208 , n16668 , n17244 );
nor ( n20209 , n20207 , n20208 );
xnor ( n20210 , n20209 , n17191 );
and ( n20211 , n17907 , n16378 );
and ( n20212 , n17688 , n16376 );
nor ( n20213 , n20211 , n20212 );
xnor ( n20214 , n20213 , n16313 );
and ( n20215 , n20210 , n20214 );
and ( n20216 , n18197 , n16176 );
and ( n20217 , n18044 , n16174 );
nor ( n20218 , n20216 , n20217 );
xnor ( n20219 , n20218 , n16075 );
and ( n20220 , n20214 , n20219 );
and ( n20221 , n20210 , n20219 );
or ( n20222 , n20215 , n20220 , n20221 );
and ( n20223 , n16151 , n18187 );
and ( n20224 , n16004 , n18184 );
nor ( n20225 , n20223 , n20224 );
xnor ( n20226 , n20225 , n17661 );
and ( n20227 , n18197 , n16174 );
not ( n20228 , n20227 );
and ( n20229 , n20228 , n16075 );
and ( n20230 , n20226 , n20229 );
and ( n20231 , n20222 , n20230 );
and ( n20232 , n17610 , n16565 );
and ( n20233 , n17355 , n16563 );
nor ( n20234 , n20232 , n20233 );
xnor ( n20235 , n20234 , n16481 );
and ( n20236 , n20230 , n20235 );
and ( n20237 , n20222 , n20235 );
or ( n20238 , n20231 , n20236 , n20237 );
xor ( n20239 , n19971 , n19975 );
xor ( n20240 , n20239 , n19980 );
and ( n20241 , n20238 , n20240 );
xor ( n20242 , n20125 , n20137 );
xor ( n20243 , n20242 , n20154 );
and ( n20244 , n20240 , n20243 );
and ( n20245 , n20238 , n20243 );
or ( n20246 , n20241 , n20244 , n20245 );
and ( n20247 , n16401 , n17915 );
and ( n20248 , n16285 , n17913 );
nor ( n20249 , n20247 , n20248 );
xnor ( n20250 , n20249 , n17664 );
and ( n20251 , n16592 , n17542 );
and ( n20252 , n16510 , n17540 );
nor ( n20253 , n20251 , n20252 );
xnor ( n20254 , n20253 , n17406 );
and ( n20255 , n20250 , n20254 );
and ( n20256 , n16995 , n17020 );
and ( n20257 , n16910 , n17018 );
nor ( n20258 , n20256 , n20257 );
xnor ( n20259 , n20258 , n16938 );
and ( n20260 , n20254 , n20259 );
and ( n20261 , n20250 , n20259 );
or ( n20262 , n20255 , n20260 , n20261 );
xor ( n20263 , n20129 , n20133 );
xor ( n20264 , n20263 , n19938 );
and ( n20265 , n20262 , n20264 );
xor ( n20266 , n20161 , n20165 );
xor ( n20267 , n20266 , n20170 );
and ( n20268 , n20264 , n20267 );
and ( n20269 , n20262 , n20267 );
or ( n20270 , n20265 , n20268 , n20269 );
xor ( n20271 , n20226 , n20229 );
and ( n20272 , n17355 , n16782 );
and ( n20273 , n17309 , n16780 );
nor ( n20274 , n20272 , n20273 );
xnor ( n20275 , n20274 , n16696 );
and ( n20276 , n20271 , n20275 );
and ( n20277 , n17720 , n16565 );
and ( n20278 , n17610 , n16563 );
nor ( n20279 , n20277 , n20278 );
xnor ( n20280 , n20279 , n16481 );
and ( n20281 , n20275 , n20280 );
and ( n20282 , n20271 , n20280 );
or ( n20283 , n20276 , n20281 , n20282 );
xor ( n20284 , n20142 , n20146 );
xor ( n20285 , n20284 , n20151 );
and ( n20286 , n20283 , n20285 );
xor ( n20287 , n20222 , n20230 );
xor ( n20288 , n20287 , n20235 );
and ( n20289 , n20285 , n20288 );
and ( n20290 , n20283 , n20288 );
or ( n20291 , n20286 , n20289 , n20290 );
and ( n20292 , n20270 , n20291 );
xor ( n20293 , n20173 , n20175 );
xor ( n20294 , n20293 , n20178 );
and ( n20295 , n20291 , n20294 );
and ( n20296 , n20270 , n20294 );
or ( n20297 , n20292 , n20295 , n20296 );
and ( n20298 , n20246 , n20297 );
xor ( n20299 , n20189 , n20191 );
xor ( n20300 , n20299 , n20194 );
and ( n20301 , n20297 , n20300 );
and ( n20302 , n20246 , n20300 );
or ( n20303 , n20298 , n20301 , n20302 );
and ( n20304 , n20206 , n20303 );
xor ( n20305 , n20246 , n20297 );
xor ( n20306 , n20305 , n20300 );
and ( n20307 , n16285 , n18187 );
and ( n20308 , n16151 , n18184 );
nor ( n20309 , n20307 , n20308 );
xnor ( n20310 , n20309 , n17661 );
and ( n20311 , n16510 , n17915 );
and ( n20312 , n16401 , n17913 );
nor ( n20313 , n20311 , n20312 );
xnor ( n20314 , n20313 , n17664 );
and ( n20315 , n20310 , n20314 );
and ( n20316 , n20314 , n20227 );
and ( n20317 , n20310 , n20227 );
or ( n20318 , n20315 , n20316 , n20317 );
and ( n20319 , n16668 , n17542 );
and ( n20320 , n16592 , n17540 );
nor ( n20321 , n20319 , n20320 );
xnor ( n20322 , n20321 , n17406 );
and ( n20323 , n17610 , n16782 );
and ( n20324 , n17355 , n16780 );
nor ( n20325 , n20323 , n20324 );
xnor ( n20326 , n20325 , n16696 );
and ( n20327 , n20322 , n20326 );
and ( n20328 , n17688 , n16565 );
and ( n20329 , n17720 , n16563 );
nor ( n20330 , n20328 , n20329 );
xnor ( n20331 , n20330 , n16481 );
and ( n20332 , n20326 , n20331 );
and ( n20333 , n20322 , n20331 );
or ( n20334 , n20327 , n20332 , n20333 );
and ( n20335 , n20318 , n20334 );
and ( n20336 , n16910 , n17246 );
and ( n20337 , n16792 , n17244 );
nor ( n20338 , n20336 , n20337 );
xnor ( n20339 , n20338 , n17191 );
and ( n20340 , n17309 , n17020 );
and ( n20341 , n16995 , n17018 );
nor ( n20342 , n20340 , n20341 );
xnor ( n20343 , n20342 , n16938 );
and ( n20344 , n20339 , n20343 );
and ( n20345 , n18044 , n16378 );
and ( n20346 , n17907 , n16376 );
nor ( n20347 , n20345 , n20346 );
xnor ( n20348 , n20347 , n16313 );
and ( n20349 , n20343 , n20348 );
and ( n20350 , n20339 , n20348 );
or ( n20351 , n20344 , n20349 , n20350 );
and ( n20352 , n20334 , n20351 );
and ( n20353 , n20318 , n20351 );
or ( n20354 , n20335 , n20352 , n20353 );
xor ( n20355 , n20210 , n20214 );
xor ( n20356 , n20355 , n20219 );
xor ( n20357 , n20250 , n20254 );
xor ( n20358 , n20357 , n20259 );
and ( n20359 , n20356 , n20358 );
xor ( n20360 , n20271 , n20275 );
xor ( n20361 , n20360 , n20280 );
and ( n20362 , n20358 , n20361 );
and ( n20363 , n20356 , n20361 );
or ( n20364 , n20359 , n20362 , n20363 );
and ( n20365 , n20354 , n20364 );
xor ( n20366 , n20262 , n20264 );
xor ( n20367 , n20366 , n20267 );
and ( n20368 , n20364 , n20367 );
and ( n20369 , n20354 , n20367 );
or ( n20370 , n20365 , n20368 , n20369 );
xor ( n20371 , n20238 , n20240 );
xor ( n20372 , n20371 , n20243 );
and ( n20373 , n20370 , n20372 );
xor ( n20374 , n20270 , n20291 );
xor ( n20375 , n20374 , n20294 );
and ( n20376 , n20372 , n20375 );
and ( n20377 , n20370 , n20375 );
or ( n20378 , n20373 , n20376 , n20377 );
and ( n20379 , n20306 , n20378 );
xor ( n20380 , n20370 , n20372 );
xor ( n20381 , n20380 , n20375 );
and ( n20382 , n16592 , n17915 );
and ( n20383 , n16510 , n17913 );
nor ( n20384 , n20382 , n20383 );
xnor ( n20385 , n20384 , n17664 );
and ( n20386 , n16995 , n17246 );
and ( n20387 , n16910 , n17244 );
nor ( n20388 , n20386 , n20387 );
xnor ( n20389 , n20388 , n17191 );
and ( n20390 , n20385 , n20389 );
and ( n20391 , n18197 , n16378 );
and ( n20392 , n18044 , n16376 );
nor ( n20393 , n20391 , n20392 );
xnor ( n20394 , n20393 , n16313 );
and ( n20395 , n20389 , n20394 );
and ( n20396 , n20385 , n20394 );
or ( n20397 , n20390 , n20395 , n20396 );
and ( n20398 , n16792 , n17542 );
and ( n20399 , n16668 , n17540 );
nor ( n20400 , n20398 , n20399 );
xnor ( n20401 , n20400 , n17406 );
and ( n20402 , n17355 , n17020 );
and ( n20403 , n17309 , n17018 );
nor ( n20404 , n20402 , n20403 );
xnor ( n20405 , n20404 , n16938 );
and ( n20406 , n20401 , n20405 );
and ( n20407 , n17720 , n16782 );
and ( n20408 , n17610 , n16780 );
nor ( n20409 , n20407 , n20408 );
xnor ( n20410 , n20409 , n16696 );
and ( n20411 , n20405 , n20410 );
and ( n20412 , n20401 , n20410 );
or ( n20413 , n20406 , n20411 , n20412 );
and ( n20414 , n20397 , n20413 );
and ( n20415 , n16401 , n18187 );
and ( n20416 , n16285 , n18184 );
nor ( n20417 , n20415 , n20416 );
xnor ( n20418 , n20417 , n17661 );
and ( n20419 , n18197 , n16376 );
not ( n20420 , n20419 );
and ( n20421 , n20420 , n16313 );
and ( n20422 , n20418 , n20421 );
and ( n20423 , n20413 , n20422 );
and ( n20424 , n20397 , n20422 );
or ( n20425 , n20414 , n20423 , n20424 );
xor ( n20426 , n20310 , n20314 );
xor ( n20427 , n20426 , n20227 );
xor ( n20428 , n20322 , n20326 );
xor ( n20429 , n20428 , n20331 );
and ( n20430 , n20427 , n20429 );
xor ( n20431 , n20339 , n20343 );
xor ( n20432 , n20431 , n20348 );
and ( n20433 , n20429 , n20432 );
and ( n20434 , n20427 , n20432 );
or ( n20435 , n20430 , n20433 , n20434 );
and ( n20436 , n20425 , n20435 );
xor ( n20437 , n20318 , n20334 );
xor ( n20438 , n20437 , n20351 );
and ( n20439 , n20435 , n20438 );
and ( n20440 , n20425 , n20438 );
or ( n20441 , n20436 , n20439 , n20440 );
xor ( n20442 , n20283 , n20285 );
xor ( n20443 , n20442 , n20288 );
and ( n20444 , n20441 , n20443 );
xor ( n20445 , n20354 , n20364 );
xor ( n20446 , n20445 , n20367 );
and ( n20447 , n20443 , n20446 );
and ( n20448 , n20441 , n20446 );
or ( n20449 , n20444 , n20447 , n20448 );
and ( n20450 , n20381 , n20449 );
xor ( n20451 , n20356 , n20358 );
xor ( n20452 , n20451 , n20361 );
xor ( n20453 , n20425 , n20435 );
xor ( n20454 , n20453 , n20438 );
and ( n20455 , n20452 , n20454 );
xor ( n20456 , n20418 , n20421 );
and ( n20457 , n16510 , n18187 );
and ( n20458 , n16401 , n18184 );
nor ( n20459 , n20457 , n20458 );
xnor ( n20460 , n20459 , n17661 );
and ( n20461 , n16668 , n17915 );
and ( n20462 , n16592 , n17913 );
nor ( n20463 , n20461 , n20462 );
xnor ( n20464 , n20463 , n17664 );
and ( n20465 , n20460 , n20464 );
and ( n20466 , n20464 , n20419 );
and ( n20467 , n20460 , n20419 );
or ( n20468 , n20465 , n20466 , n20467 );
and ( n20469 , n20456 , n20468 );
and ( n20470 , n17907 , n16565 );
and ( n20471 , n17688 , n16563 );
nor ( n20472 , n20470 , n20471 );
xnor ( n20473 , n20472 , n16481 );
and ( n20474 , n20468 , n20473 );
and ( n20475 , n20456 , n20473 );
or ( n20476 , n20469 , n20474 , n20475 );
xor ( n20477 , n20397 , n20413 );
xor ( n20478 , n20477 , n20422 );
and ( n20479 , n20476 , n20478 );
and ( n20480 , n20454 , n20479 );
and ( n20481 , n20452 , n20479 );
or ( n20482 , n20455 , n20480 , n20481 );
xor ( n20483 , n20441 , n20443 );
xor ( n20484 , n20483 , n20446 );
and ( n20485 , n20482 , n20484 );
and ( n20486 , n16592 , n18187 );
and ( n20487 , n16510 , n18184 );
nor ( n20488 , n20486 , n20487 );
xnor ( n20489 , n20488 , n17661 );
and ( n20490 , n18197 , n16563 );
not ( n20491 , n20490 );
and ( n20492 , n20491 , n16481 );
and ( n20493 , n20489 , n20492 );
and ( n20494 , n17688 , n16782 );
and ( n20495 , n17720 , n16780 );
nor ( n20496 , n20494 , n20495 );
xnor ( n20497 , n20496 , n16696 );
and ( n20498 , n20493 , n20497 );
and ( n20499 , n18044 , n16565 );
and ( n20500 , n17907 , n16563 );
nor ( n20501 , n20499 , n20500 );
xnor ( n20502 , n20501 , n16481 );
and ( n20503 , n20497 , n20502 );
and ( n20504 , n20493 , n20502 );
or ( n20505 , n20498 , n20503 , n20504 );
and ( n20506 , n16792 , n17915 );
and ( n20507 , n16668 , n17913 );
nor ( n20508 , n20506 , n20507 );
xnor ( n20509 , n20508 , n17664 );
and ( n20510 , n17355 , n17246 );
and ( n20511 , n17309 , n17244 );
nor ( n20512 , n20510 , n20511 );
xnor ( n20513 , n20512 , n17191 );
and ( n20514 , n20509 , n20513 );
and ( n20515 , n17720 , n17020 );
and ( n20516 , n17610 , n17018 );
nor ( n20517 , n20515 , n20516 );
xnor ( n20518 , n20517 , n16938 );
and ( n20519 , n20513 , n20518 );
and ( n20520 , n20509 , n20518 );
or ( n20521 , n20514 , n20519 , n20520 );
and ( n20522 , n16995 , n17542 );
and ( n20523 , n16910 , n17540 );
nor ( n20524 , n20522 , n20523 );
xnor ( n20525 , n20524 , n17406 );
and ( n20526 , n17907 , n16782 );
and ( n20527 , n17688 , n16780 );
nor ( n20528 , n20526 , n20527 );
xnor ( n20529 , n20528 , n16696 );
and ( n20530 , n20525 , n20529 );
and ( n20531 , n18197 , n16565 );
and ( n20532 , n18044 , n16563 );
nor ( n20533 , n20531 , n20532 );
xnor ( n20534 , n20533 , n16481 );
and ( n20535 , n20529 , n20534 );
and ( n20536 , n20525 , n20534 );
or ( n20537 , n20530 , n20535 , n20536 );
and ( n20538 , n20521 , n20537 );
xor ( n20539 , n20460 , n20464 );
xor ( n20540 , n20539 , n20419 );
and ( n20541 , n20537 , n20540 );
and ( n20542 , n20521 , n20540 );
or ( n20543 , n20538 , n20541 , n20542 );
and ( n20544 , n20505 , n20543 );
xor ( n20545 , n20456 , n20468 );
xor ( n20546 , n20545 , n20473 );
and ( n20547 , n20543 , n20546 );
and ( n20548 , n20505 , n20546 );
or ( n20549 , n20544 , n20547 , n20548 );
xor ( n20550 , n20427 , n20429 );
xor ( n20551 , n20550 , n20432 );
and ( n20552 , n20549 , n20551 );
xor ( n20553 , n20452 , n20454 );
xor ( n20554 , n20553 , n20479 );
and ( n20555 , n20552 , n20554 );
xor ( n20556 , n20385 , n20389 );
xor ( n20557 , n20556 , n20394 );
xor ( n20558 , n20401 , n20405 );
xor ( n20559 , n20558 , n20410 );
and ( n20560 , n20557 , n20559 );
and ( n20561 , n16910 , n17542 );
and ( n20562 , n16792 , n17540 );
nor ( n20563 , n20561 , n20562 );
xnor ( n20564 , n20563 , n17406 );
and ( n20565 , n17309 , n17246 );
and ( n20566 , n16995 , n17244 );
nor ( n20567 , n20565 , n20566 );
xnor ( n20568 , n20567 , n17191 );
and ( n20569 , n20564 , n20568 );
and ( n20570 , n17610 , n17020 );
and ( n20571 , n17355 , n17018 );
nor ( n20572 , n20570 , n20571 );
xnor ( n20573 , n20572 , n16938 );
and ( n20574 , n20568 , n20573 );
and ( n20575 , n20564 , n20573 );
or ( n20576 , n20569 , n20574 , n20575 );
and ( n20577 , n20559 , n20576 );
and ( n20578 , n20557 , n20576 );
or ( n20579 , n20560 , n20577 , n20578 );
xor ( n20580 , n20476 , n20478 );
and ( n20581 , n20579 , n20580 );
xor ( n20582 , n20549 , n20551 );
and ( n20583 , n20580 , n20582 );
and ( n20584 , n20579 , n20582 );
or ( n20585 , n20581 , n20583 , n20584 );
and ( n20586 , n20554 , n20585 );
and ( n20587 , n20552 , n20585 );
or ( n20588 , n20555 , n20586 , n20587 );
and ( n20589 , n20484 , n20588 );
and ( n20590 , n20482 , n20588 );
or ( n20591 , n20485 , n20589 , n20590 );
and ( n20592 , n20449 , n20591 );
and ( n20593 , n20381 , n20591 );
or ( n20594 , n20450 , n20592 , n20593 );
and ( n20595 , n20378 , n20594 );
and ( n20596 , n20306 , n20594 );
or ( n20597 , n20379 , n20595 , n20596 );
and ( n20598 , n20303 , n20597 );
and ( n20599 , n20206 , n20597 );
or ( n20600 , n20304 , n20598 , n20599 );
and ( n20601 , n20203 , n20600 );
and ( n20602 , n20124 , n20600 );
or ( n20603 , n20204 , n20601 , n20602 );
and ( n20604 , n20122 , n20603 );
xor ( n20605 , n20122 , n20603 );
xor ( n20606 , n20124 , n20203 );
xor ( n20607 , n20606 , n20600 );
xor ( n20608 , n20206 , n20303 );
xor ( n20609 , n20608 , n20597 );
xor ( n20610 , n20306 , n20378 );
xor ( n20611 , n20610 , n20594 );
xor ( n20612 , n20381 , n20449 );
xor ( n20613 , n20612 , n20591 );
xor ( n20614 , n20482 , n20484 );
xor ( n20615 , n20614 , n20588 );
xor ( n20616 , n20552 , n20554 );
xor ( n20617 , n20616 , n20585 );
xor ( n20618 , n20557 , n20559 );
xor ( n20619 , n20618 , n20576 );
xor ( n20620 , n20505 , n20543 );
xor ( n20621 , n20620 , n20546 );
and ( n20622 , n20619 , n20621 );
xor ( n20623 , n20564 , n20568 );
xor ( n20624 , n20623 , n20573 );
xor ( n20625 , n20493 , n20497 );
xor ( n20626 , n20625 , n20502 );
and ( n20627 , n20624 , n20626 );
and ( n20628 , n16910 , n17915 );
and ( n20629 , n16792 , n17913 );
nor ( n20630 , n20628 , n20629 );
xnor ( n20631 , n20630 , n17664 );
and ( n20632 , n17610 , n17246 );
and ( n20633 , n17355 , n17244 );
nor ( n20634 , n20632 , n20633 );
xnor ( n20635 , n20634 , n17191 );
and ( n20636 , n20631 , n20635 );
and ( n20637 , n20635 , n20490 );
and ( n20638 , n20631 , n20490 );
or ( n20639 , n20636 , n20637 , n20638 );
xor ( n20640 , n20489 , n20492 );
and ( n20641 , n20639 , n20640 );
and ( n20642 , n20626 , n20641 );
and ( n20643 , n20624 , n20641 );
or ( n20644 , n20627 , n20642 , n20643 );
and ( n20645 , n20621 , n20644 );
and ( n20646 , n20619 , n20644 );
or ( n20647 , n20622 , n20645 , n20646 );
xor ( n20648 , n20579 , n20580 );
xor ( n20649 , n20648 , n20582 );
and ( n20650 , n20647 , n20649 );
and ( n20651 , n16792 , n18187 );
and ( n20652 , n16668 , n18184 );
nor ( n20653 , n20651 , n20652 );
xnor ( n20654 , n20653 , n17661 );
and ( n20655 , n17720 , n17246 );
and ( n20656 , n17610 , n17244 );
nor ( n20657 , n20655 , n20656 );
xnor ( n20658 , n20657 , n17191 );
and ( n20659 , n20654 , n20658 );
and ( n20660 , n17907 , n17020 );
and ( n20661 , n17688 , n17018 );
nor ( n20662 , n20660 , n20661 );
xnor ( n20663 , n20662 , n16938 );
and ( n20664 , n20658 , n20663 );
and ( n20665 , n20654 , n20663 );
or ( n20666 , n20659 , n20664 , n20665 );
and ( n20667 , n16995 , n17915 );
and ( n20668 , n16910 , n17913 );
nor ( n20669 , n20667 , n20668 );
xnor ( n20670 , n20669 , n17664 );
and ( n20671 , n18197 , n16780 );
not ( n20672 , n20671 );
and ( n20673 , n20672 , n16696 );
and ( n20674 , n20670 , n20673 );
and ( n20675 , n20666 , n20674 );
and ( n20676 , n17309 , n17542 );
and ( n20677 , n16995 , n17540 );
nor ( n20678 , n20676 , n20677 );
xnor ( n20679 , n20678 , n17406 );
and ( n20680 , n20674 , n20679 );
and ( n20681 , n20666 , n20679 );
or ( n20682 , n20675 , n20680 , n20681 );
xor ( n20683 , n20509 , n20513 );
xor ( n20684 , n20683 , n20518 );
and ( n20685 , n20682 , n20684 );
xor ( n20686 , n20525 , n20529 );
xor ( n20687 , n20686 , n20534 );
and ( n20688 , n20684 , n20687 );
and ( n20689 , n20682 , n20687 );
or ( n20690 , n20685 , n20688 , n20689 );
xor ( n20691 , n20521 , n20537 );
xor ( n20692 , n20691 , n20540 );
and ( n20693 , n20690 , n20692 );
xor ( n20694 , n20619 , n20621 );
xor ( n20695 , n20694 , n20644 );
and ( n20696 , n20693 , n20695 );
xor ( n20697 , n20624 , n20626 );
xor ( n20698 , n20697 , n20641 );
xor ( n20699 , n20690 , n20692 );
and ( n20700 , n20698 , n20699 );
and ( n20701 , n16668 , n18187 );
and ( n20702 , n16592 , n18184 );
nor ( n20703 , n20701 , n20702 );
xnor ( n20704 , n20703 , n17661 );
and ( n20705 , n17688 , n17020 );
and ( n20706 , n17720 , n17018 );
nor ( n20707 , n20705 , n20706 );
xnor ( n20708 , n20707 , n16938 );
and ( n20709 , n20704 , n20708 );
and ( n20710 , n18044 , n16782 );
and ( n20711 , n17907 , n16780 );
nor ( n20712 , n20710 , n20711 );
xnor ( n20713 , n20712 , n16696 );
and ( n20714 , n20708 , n20713 );
and ( n20715 , n20704 , n20713 );
or ( n20716 , n20709 , n20714 , n20715 );
xor ( n20717 , n20639 , n20640 );
and ( n20718 , n20716 , n20717 );
xor ( n20719 , n20682 , n20684 );
xor ( n20720 , n20719 , n20687 );
and ( n20721 , n20717 , n20720 );
and ( n20722 , n20716 , n20720 );
or ( n20723 , n20718 , n20721 , n20722 );
and ( n20724 , n20699 , n20723 );
and ( n20725 , n20698 , n20723 );
or ( n20726 , n20700 , n20724 , n20725 );
and ( n20727 , n20695 , n20726 );
and ( n20728 , n20693 , n20726 );
or ( n20729 , n20696 , n20727 , n20728 );
and ( n20730 , n20649 , n20729 );
and ( n20731 , n20647 , n20729 );
or ( n20732 , n20650 , n20730 , n20731 );
and ( n20733 , n20617 , n20732 );
xor ( n20734 , n20617 , n20732 );
xor ( n20735 , n20647 , n20649 );
xor ( n20736 , n20735 , n20729 );
xor ( n20737 , n20693 , n20695 );
xor ( n20738 , n20737 , n20726 );
xor ( n20739 , n20670 , n20673 );
and ( n20740 , n17355 , n17542 );
and ( n20741 , n17309 , n17540 );
nor ( n20742 , n20740 , n20741 );
xnor ( n20743 , n20742 , n17406 );
and ( n20744 , n20739 , n20743 );
and ( n20745 , n18197 , n16782 );
and ( n20746 , n18044 , n16780 );
nor ( n20747 , n20745 , n20746 );
xnor ( n20748 , n20747 , n16696 );
and ( n20749 , n20743 , n20748 );
and ( n20750 , n20739 , n20748 );
or ( n20751 , n20744 , n20749 , n20750 );
xor ( n20752 , n20631 , n20635 );
xor ( n20753 , n20752 , n20490 );
and ( n20754 , n20751 , n20753 );
xor ( n20755 , n20704 , n20708 );
xor ( n20756 , n20755 , n20713 );
and ( n20757 , n20753 , n20756 );
and ( n20758 , n20751 , n20756 );
or ( n20759 , n20754 , n20757 , n20758 );
and ( n20760 , n16910 , n18187 );
and ( n20761 , n16792 , n18184 );
nor ( n20762 , n20760 , n20761 );
xnor ( n20763 , n20762 , n17661 );
and ( n20764 , n17610 , n17542 );
and ( n20765 , n17355 , n17540 );
nor ( n20766 , n20764 , n20765 );
xnor ( n20767 , n20766 , n17406 );
and ( n20768 , n20763 , n20767 );
and ( n20769 , n18044 , n17020 );
and ( n20770 , n17907 , n17018 );
nor ( n20771 , n20769 , n20770 );
xnor ( n20772 , n20771 , n16938 );
and ( n20773 , n20767 , n20772 );
and ( n20774 , n20763 , n20772 );
or ( n20775 , n20768 , n20773 , n20774 );
and ( n20776 , n17309 , n17915 );
and ( n20777 , n16995 , n17913 );
nor ( n20778 , n20776 , n20777 );
xnor ( n20779 , n20778 , n17664 );
and ( n20780 , n17688 , n17246 );
and ( n20781 , n17720 , n17244 );
nor ( n20782 , n20780 , n20781 );
xnor ( n20783 , n20782 , n17191 );
and ( n20784 , n20779 , n20783 );
and ( n20785 , n20783 , n20671 );
and ( n20786 , n20779 , n20671 );
or ( n20787 , n20784 , n20785 , n20786 );
and ( n20788 , n20775 , n20787 );
xor ( n20789 , n20654 , n20658 );
xor ( n20790 , n20789 , n20663 );
and ( n20791 , n20787 , n20790 );
and ( n20792 , n20775 , n20790 );
or ( n20793 , n20788 , n20791 , n20792 );
xor ( n20794 , n20666 , n20674 );
xor ( n20795 , n20794 , n20679 );
and ( n20796 , n20793 , n20795 );
xor ( n20797 , n20751 , n20753 );
xor ( n20798 , n20797 , n20756 );
and ( n20799 , n20795 , n20798 );
and ( n20800 , n20793 , n20798 );
or ( n20801 , n20796 , n20799 , n20800 );
and ( n20802 , n20759 , n20801 );
xor ( n20803 , n20716 , n20717 );
xor ( n20804 , n20803 , n20720 );
and ( n20805 , n20801 , n20804 );
and ( n20806 , n20759 , n20804 );
or ( n20807 , n20802 , n20805 , n20806 );
xor ( n20808 , n20698 , n20699 );
xor ( n20809 , n20808 , n20723 );
and ( n20810 , n20807 , n20809 );
xor ( n20811 , n20807 , n20809 );
xor ( n20812 , n20759 , n20801 );
xor ( n20813 , n20812 , n20804 );
and ( n20814 , n16995 , n18187 );
and ( n20815 , n16910 , n18184 );
nor ( n20816 , n20814 , n20815 );
xnor ( n20817 , n20816 , n17661 );
and ( n20818 , n17907 , n17246 );
and ( n20819 , n17688 , n17244 );
nor ( n20820 , n20818 , n20819 );
xnor ( n20821 , n20820 , n17191 );
and ( n20822 , n20817 , n20821 );
and ( n20823 , n18197 , n17020 );
and ( n20824 , n18044 , n17018 );
nor ( n20825 , n20823 , n20824 );
xnor ( n20826 , n20825 , n16938 );
and ( n20827 , n20821 , n20826 );
and ( n20828 , n20817 , n20826 );
or ( n20829 , n20822 , n20827 , n20828 );
and ( n20830 , n17355 , n17915 );
and ( n20831 , n17309 , n17913 );
nor ( n20832 , n20830 , n20831 );
xnor ( n20833 , n20832 , n17664 );
and ( n20834 , n18197 , n17018 );
not ( n20835 , n20834 );
and ( n20836 , n20835 , n16938 );
and ( n20837 , n20833 , n20836 );
and ( n20838 , n20829 , n20837 );
xor ( n20839 , n20779 , n20783 );
xor ( n20840 , n20839 , n20671 );
and ( n20841 , n20837 , n20840 );
and ( n20842 , n20829 , n20840 );
or ( n20843 , n20838 , n20841 , n20842 );
xor ( n20844 , n20739 , n20743 );
xor ( n20845 , n20844 , n20748 );
and ( n20846 , n20843 , n20845 );
xor ( n20847 , n20775 , n20787 );
xor ( n20848 , n20847 , n20790 );
and ( n20849 , n20845 , n20848 );
and ( n20850 , n20843 , n20848 );
or ( n20851 , n20846 , n20849 , n20850 );
xor ( n20852 , n20793 , n20795 );
xor ( n20853 , n20852 , n20798 );
and ( n20854 , n20851 , n20853 );
xor ( n20855 , n20851 , n20853 );
xor ( n20856 , n20843 , n20845 );
xor ( n20857 , n20856 , n20848 );
xor ( n20858 , n20833 , n20836 );
and ( n20859 , n17309 , n18187 );
and ( n20860 , n16995 , n18184 );
nor ( n20861 , n20859 , n20860 );
xnor ( n20862 , n20861 , n17661 );
and ( n20863 , n18044 , n17246 );
and ( n20864 , n17907 , n17244 );
nor ( n20865 , n20863 , n20864 );
xnor ( n20866 , n20865 , n17191 );
and ( n20867 , n20862 , n20866 );
and ( n20868 , n20866 , n20834 );
and ( n20869 , n20862 , n20834 );
or ( n20870 , n20867 , n20868 , n20869 );
and ( n20871 , n20858 , n20870 );
and ( n20872 , n17720 , n17542 );
and ( n20873 , n17610 , n17540 );
nor ( n20874 , n20872 , n20873 );
xnor ( n20875 , n20874 , n17406 );
and ( n20876 , n20870 , n20875 );
and ( n20877 , n20858 , n20875 );
or ( n20878 , n20871 , n20876 , n20877 );
xor ( n20879 , n20763 , n20767 );
xor ( n20880 , n20879 , n20772 );
and ( n20881 , n20878 , n20880 );
xor ( n20882 , n20829 , n20837 );
xor ( n20883 , n20882 , n20840 );
and ( n20884 , n20880 , n20883 );
and ( n20885 , n20878 , n20883 );
or ( n20886 , n20881 , n20884 , n20885 );
and ( n20887 , n20857 , n20886 );
xor ( n20888 , n20857 , n20886 );
xor ( n20889 , n20878 , n20880 );
xor ( n20890 , n20889 , n20883 );
and ( n20891 , n17355 , n18187 );
and ( n20892 , n17309 , n18184 );
nor ( n20893 , n20891 , n20892 );
xnor ( n20894 , n20893 , n17661 );
and ( n20895 , n18197 , n17244 );
not ( n20896 , n20895 );
and ( n20897 , n20896 , n17191 );
and ( n20898 , n20894 , n20897 );
and ( n20899 , n17610 , n17915 );
and ( n20900 , n17355 , n17913 );
nor ( n20901 , n20899 , n20900 );
xnor ( n20902 , n20901 , n17664 );
and ( n20903 , n20898 , n20902 );
and ( n20904 , n17688 , n17542 );
and ( n20905 , n17720 , n17540 );
nor ( n20906 , n20904 , n20905 );
xnor ( n20907 , n20906 , n17406 );
and ( n20908 , n20902 , n20907 );
and ( n20909 , n20898 , n20907 );
or ( n20910 , n20903 , n20908 , n20909 );
xor ( n20911 , n20817 , n20821 );
xor ( n20912 , n20911 , n20826 );
and ( n20913 , n20910 , n20912 );
xor ( n20914 , n20858 , n20870 );
xor ( n20915 , n20914 , n20875 );
and ( n20916 , n20912 , n20915 );
and ( n20917 , n20910 , n20915 );
or ( n20918 , n20913 , n20916 , n20917 );
and ( n20919 , n20890 , n20918 );
xor ( n20920 , n20890 , n20918 );
xor ( n20921 , n20910 , n20912 );
xor ( n20922 , n20921 , n20915 );
and ( n20923 , n17720 , n17915 );
and ( n20924 , n17610 , n17913 );
nor ( n20925 , n20923 , n20924 );
xnor ( n20926 , n20925 , n17664 );
and ( n20927 , n17907 , n17542 );
and ( n20928 , n17688 , n17540 );
nor ( n20929 , n20927 , n20928 );
xnor ( n20930 , n20929 , n17406 );
and ( n20931 , n20926 , n20930 );
and ( n20932 , n18197 , n17246 );
and ( n20933 , n18044 , n17244 );
nor ( n20934 , n20932 , n20933 );
xnor ( n20935 , n20934 , n17191 );
and ( n20936 , n20930 , n20935 );
and ( n20937 , n20926 , n20935 );
or ( n20938 , n20931 , n20936 , n20937 );
xor ( n20939 , n20862 , n20866 );
xor ( n20940 , n20939 , n20834 );
and ( n20941 , n20938 , n20940 );
xor ( n20942 , n20898 , n20902 );
xor ( n20943 , n20942 , n20907 );
and ( n20944 , n20940 , n20943 );
and ( n20945 , n20938 , n20943 );
or ( n20946 , n20941 , n20944 , n20945 );
and ( n20947 , n20922 , n20946 );
xor ( n20948 , n20922 , n20946 );
xor ( n20949 , n20894 , n20897 );
and ( n20950 , n17610 , n18187 );
and ( n20951 , n17355 , n18184 );
nor ( n20952 , n20950 , n20951 );
xnor ( n20953 , n20952 , n17661 );
and ( n20954 , n17688 , n17915 );
and ( n20955 , n17720 , n17913 );
nor ( n20956 , n20954 , n20955 );
xnor ( n20957 , n20956 , n17664 );
and ( n20958 , n20953 , n20957 );
and ( n20959 , n20957 , n20895 );
and ( n20960 , n20953 , n20895 );
or ( n20961 , n20958 , n20959 , n20960 );
and ( n20962 , n20949 , n20961 );
xor ( n20963 , n20926 , n20930 );
xor ( n20964 , n20963 , n20935 );
and ( n20965 , n20961 , n20964 );
and ( n20966 , n20949 , n20964 );
or ( n20967 , n20962 , n20965 , n20966 );
xor ( n20968 , n20938 , n20940 );
xor ( n20969 , n20968 , n20943 );
and ( n20970 , n20967 , n20969 );
xor ( n20971 , n20967 , n20969 );
xor ( n20972 , n20949 , n20961 );
xor ( n20973 , n20972 , n20964 );
and ( n20974 , n17720 , n18187 );
and ( n20975 , n17610 , n18184 );
nor ( n20976 , n20974 , n20975 );
xnor ( n20977 , n20976 , n17661 );
and ( n20978 , n18197 , n17540 );
not ( n20979 , n20978 );
and ( n20980 , n20979 , n17406 );
and ( n20981 , n20977 , n20980 );
and ( n20982 , n18044 , n17542 );
and ( n20983 , n17907 , n17540 );
nor ( n20984 , n20982 , n20983 );
xnor ( n20985 , n20984 , n17406 );
and ( n20986 , n20981 , n20985 );
xor ( n20987 , n20953 , n20957 );
xor ( n20988 , n20987 , n20895 );
and ( n20989 , n20985 , n20988 );
and ( n20990 , n20981 , n20988 );
or ( n20991 , n20986 , n20989 , n20990 );
and ( n20992 , n20973 , n20991 );
xor ( n20993 , n20973 , n20991 );
xor ( n20994 , n20981 , n20985 );
xor ( n20995 , n20994 , n20988 );
xor ( n20996 , n20977 , n20980 );
and ( n20997 , n17907 , n17915 );
and ( n20998 , n17688 , n17913 );
nor ( n20999 , n20997 , n20998 );
xnor ( n21000 , n20999 , n17664 );
and ( n21001 , n20996 , n21000 );
and ( n21002 , n18197 , n17542 );
and ( n21003 , n18044 , n17540 );
nor ( n21004 , n21002 , n21003 );
xnor ( n21005 , n21004 , n17406 );
and ( n21006 , n21000 , n21005 );
and ( n21007 , n20996 , n21005 );
or ( n21008 , n21001 , n21006 , n21007 );
and ( n21009 , n20995 , n21008 );
xor ( n21010 , n20995 , n21008 );
and ( n21011 , n17688 , n18187 );
and ( n21012 , n17720 , n18184 );
nor ( n21013 , n21011 , n21012 );
xnor ( n21014 , n21013 , n17661 );
and ( n21015 , n18044 , n17915 );
and ( n21016 , n17907 , n17913 );
nor ( n21017 , n21015 , n21016 );
xnor ( n21018 , n21017 , n17664 );
and ( n21019 , n21014 , n21018 );
and ( n21020 , n21018 , n20978 );
and ( n21021 , n21014 , n20978 );
or ( n21022 , n21019 , n21020 , n21021 );
xor ( n21023 , n20996 , n21000 );
xor ( n21024 , n21023 , n21005 );
and ( n21025 , n21022 , n21024 );
xor ( n21026 , n21022 , n21024 );
xor ( n21027 , n21014 , n21018 );
xor ( n21028 , n21027 , n20978 );
and ( n21029 , n17907 , n18187 );
and ( n21030 , n17688 , n18184 );
nor ( n21031 , n21029 , n21030 );
xnor ( n21032 , n21031 , n17661 );
and ( n21033 , n18197 , n17913 );
not ( n21034 , n21033 );
and ( n21035 , n21034 , n17664 );
and ( n21036 , n21032 , n21035 );
and ( n21037 , n21028 , n21036 );
xor ( n21038 , n21028 , n21036 );
and ( n21039 , n18197 , n17915 );
and ( n21040 , n18044 , n17913 );
nor ( n21041 , n21039 , n21040 );
xnor ( n21042 , n21041 , n17664 );
xor ( n21043 , n21032 , n21035 );
and ( n21044 , n21042 , n21043 );
xor ( n21045 , n21042 , n21043 );
and ( n21046 , n18044 , n18187 );
and ( n21047 , n17907 , n18184 );
nor ( n21048 , n21046 , n21047 );
xnor ( n21049 , n21048 , n17661 );
and ( n21050 , n21049 , n21033 );
xor ( n21051 , n21049 , n21033 );
and ( n21052 , n18197 , n18187 );
and ( n21053 , n18044 , n18184 );
nor ( n21054 , n21052 , n21053 );
xnor ( n21055 , n21054 , n17661 );
and ( n21056 , n18197 , n18184 );
not ( n21057 , n21056 );
and ( n21058 , n21057 , n17661 );
and ( n21059 , n21055 , n21058 );
and ( n21060 , n21051 , n21059 );
or ( n21061 , n21050 , n21060 );
and ( n21062 , n21045 , n21061 );
or ( n21063 , n21044 , n21062 );
and ( n21064 , n21038 , n21063 );
or ( n21065 , n21037 , n21064 );
and ( n21066 , n21026 , n21065 );
or ( n21067 , n21025 , n21066 );
and ( n21068 , n21010 , n21067 );
or ( n21069 , n21009 , n21068 );
and ( n21070 , n20993 , n21069 );
or ( n21071 , n20992 , n21070 );
and ( n21072 , n20971 , n21071 );
or ( n21073 , n20970 , n21072 );
and ( n21074 , n20948 , n21073 );
or ( n21075 , n20947 , n21074 );
and ( n21076 , n20920 , n21075 );
or ( n21077 , n20919 , n21076 );
and ( n21078 , n20888 , n21077 );
or ( n21079 , n20887 , n21078 );
and ( n21080 , n20855 , n21079 );
or ( n21081 , n20854 , n21080 );
and ( n21082 , n20813 , n21081 );
and ( n21083 , n20811 , n21082 );
or ( n21084 , n20810 , n21083 );
and ( n21085 , n20738 , n21084 );
and ( n21086 , n20736 , n21085 );
and ( n21087 , n20734 , n21086 );
or ( n21088 , n20733 , n21087 );
and ( n21089 , n20615 , n21088 );
and ( n21090 , n20613 , n21089 );
and ( n21091 , n20611 , n21090 );
and ( n21092 , n20609 , n21091 );
and ( n21093 , n20607 , n21092 );
and ( n21094 , n20605 , n21093 );
or ( n21095 , n20604 , n21094 );
and ( n21096 , n20120 , n21095 );
and ( n21097 , n20118 , n21096 );
or ( n21098 , n20117 , n21097 );
and ( n21099 , n20073 , n21098 );
and ( n21100 , n20071 , n21099 );
and ( n21101 , n20069 , n21100 );
and ( n21102 , n20067 , n21101 );
and ( n21103 , n20065 , n21102 );
or ( n21104 , n20064 , n21103 );
and ( n21105 , n19419 , n21104 );
or ( n21106 , n19418 , n21105 );
and ( n21107 , n19259 , n21106 );
and ( n21108 , n19257 , n21107 );
and ( n21109 , n19255 , n21108 );
and ( n21110 , n19253 , n21109 );
and ( n21111 , n19251 , n21110 );
and ( n21112 , n19249 , n21111 );
and ( n21113 , n19247 , n21112 );
and ( n21114 , n19245 , n21113 );
and ( n21115 , n19243 , n21114 );
and ( n21116 , n19241 , n21115 );
and ( n21117 , n19239 , n21116 );
and ( n21118 , n19237 , n21117 );
and ( n21119 , n19235 , n21118 );
and ( n21120 , n19233 , n21119 );
and ( n21121 , n19231 , n21120 );
and ( n21122 , n19229 , n21121 );
and ( n21123 , n19227 , n21122 );
and ( n21124 , n19225 , n21123 );
and ( n21125 , n19223 , n21124 );
xor ( n21126 , n19221 , n21125 );
buf ( n21127 , n21126 );
buf ( n21128 , n21127 );
buf ( n21129 , n21128 );
buf ( n21130 , n1178 );
buf ( n21131 , n21130 );
buf ( n21132 , n1179 );
buf ( n21133 , n21132 );
xor ( n21134 , n21131 , n21133 );
buf ( n21135 , n1180 );
buf ( n21136 , n21135 );
xor ( n21137 , n21133 , n21136 );
not ( n21138 , n21137 );
and ( n21139 , n21134 , n21138 );
and ( n21140 , n21129 , n21139 );
and ( n21141 , n16213 , n16241 );
and ( n21142 , n16241 , n16273 );
and ( n21143 , n16213 , n16273 );
or ( n21144 , n21141 , n21142 , n21143 );
and ( n21145 , n16217 , n16228 );
and ( n21146 , n16228 , n16240 );
and ( n21147 , n16217 , n16240 );
or ( n21148 , n21145 , n21146 , n21147 );
and ( n21149 , n16246 , n16250 );
and ( n21150 , n16250 , n16272 );
and ( n21151 , n16246 , n16272 );
or ( n21152 , n21149 , n21150 , n21151 );
xor ( n21153 , n21148 , n21152 );
and ( n21154 , n16255 , n16259 );
and ( n21155 , n16259 , n16271 );
and ( n21156 , n16255 , n16271 );
or ( n21157 , n21154 , n21155 , n21156 );
and ( n21158 , n16221 , n16225 );
and ( n21159 , n16225 , n16227 );
and ( n21160 , n16221 , n16227 );
or ( n21161 , n21158 , n21159 , n21160 );
and ( n21162 , n16261 , n16265 );
and ( n21163 , n16265 , n16270 );
and ( n21164 , n16261 , n16270 );
or ( n21165 , n21162 , n21163 , n21164 );
xor ( n21166 , n21161 , n21165 );
and ( n21167 , n16087 , n16018 );
not ( n21168 , n21167 );
xnor ( n21169 , n21168 , n16026 );
not ( n21170 , n21169 );
xor ( n21171 , n21166 , n21170 );
xor ( n21172 , n21157 , n21171 );
and ( n21173 , n16230 , n16234 );
and ( n21174 , n16234 , n16239 );
and ( n21175 , n16230 , n16239 );
or ( n21176 , n21173 , n21174 , n21175 );
and ( n21177 , n16105 , n15971 );
and ( n21178 , n16008 , n15969 );
nor ( n21179 , n21177 , n21178 );
xnor ( n21180 , n21179 , n15979 );
and ( n21181 , n16058 , n15992 );
and ( n21182 , n16029 , n15990 );
nor ( n21183 , n21181 , n21182 );
xnor ( n21184 , n21183 , n16000 );
xor ( n21185 , n21180 , n21184 );
and ( n21186 , n16049 , n15984 );
xor ( n21187 , n21185 , n21186 );
xor ( n21188 , n21176 , n21187 );
and ( n21189 , n16021 , n16102 );
and ( n21190 , n16078 , n16100 );
nor ( n21191 , n21189 , n21190 );
xnor ( n21192 , n21191 , n16110 );
and ( n21193 , n15974 , n16037 );
and ( n21194 , n16096 , n16035 );
nor ( n21195 , n21193 , n21194 );
xnor ( n21196 , n21195 , n16045 );
xor ( n21197 , n21192 , n21196 );
and ( n21198 , n16040 , n16055 );
and ( n21199 , n15961 , n16053 );
nor ( n21200 , n21198 , n21199 );
xnor ( n21201 , n21200 , n16063 );
xor ( n21202 , n21197 , n21201 );
xor ( n21203 , n21188 , n21202 );
xor ( n21204 , n21172 , n21203 );
xor ( n21205 , n21153 , n21204 );
xor ( n21206 , n21144 , n21205 );
and ( n21207 , n16274 , n16445 );
and ( n21208 , n16445 , n19220 );
and ( n21209 , n16274 , n19220 );
or ( n21210 , n21207 , n21208 , n21209 );
xor ( n21211 , n21206 , n21210 );
and ( n21212 , n19221 , n21125 );
xor ( n21213 , n21211 , n21212 );
buf ( n21214 , n21213 );
buf ( n21215 , n21214 );
buf ( n21216 , n21215 );
and ( n21217 , n21216 , n21137 );
nor ( n21218 , n21140 , n21217 );
and ( n21219 , n21133 , n21136 );
not ( n21220 , n21219 );
and ( n21221 , n21131 , n21220 );
xnor ( n21222 , n21218 , n21221 );
xor ( n21223 , n19237 , n21117 );
buf ( n21224 , n21223 );
buf ( n21225 , n21224 );
buf ( n21226 , n21225 );
buf ( n21227 , n1170 );
buf ( n21228 , n21227 );
buf ( n21229 , n1171 );
buf ( n21230 , n21229 );
xor ( n21231 , n21228 , n21230 );
buf ( n21232 , n1172 );
buf ( n21233 , n21232 );
xor ( n21234 , n21230 , n21233 );
not ( n21235 , n21234 );
and ( n21236 , n21231 , n21235 );
and ( n21237 , n21226 , n21236 );
xor ( n21238 , n19235 , n21118 );
buf ( n21239 , n21238 );
buf ( n21240 , n21239 );
buf ( n21241 , n21240 );
and ( n21242 , n21241 , n21234 );
nor ( n21243 , n21237 , n21242 );
and ( n21244 , n21230 , n21233 );
not ( n21245 , n21244 );
and ( n21246 , n21228 , n21245 );
xnor ( n21247 , n21243 , n21246 );
and ( n21248 , n21222 , n21247 );
xor ( n21249 , n19241 , n21115 );
buf ( n21250 , n21249 );
buf ( n21251 , n21250 );
buf ( n21252 , n21251 );
buf ( n21253 , n1168 );
buf ( n21254 , n21253 );
buf ( n21255 , n1169 );
buf ( n21256 , n21255 );
xor ( n21257 , n21254 , n21256 );
xor ( n21258 , n21256 , n21228 );
not ( n21259 , n21258 );
and ( n21260 , n21257 , n21259 );
and ( n21261 , n21252 , n21260 );
xor ( n21262 , n19239 , n21116 );
buf ( n21263 , n21262 );
buf ( n21264 , n21263 );
buf ( n21265 , n21264 );
and ( n21266 , n21265 , n21258 );
nor ( n21267 , n21261 , n21266 );
and ( n21268 , n21256 , n21228 );
not ( n21269 , n21268 );
and ( n21270 , n21254 , n21269 );
xnor ( n21271 , n21267 , n21270 );
and ( n21272 , n21247 , n21271 );
and ( n21273 , n21222 , n21271 );
or ( n21274 , n21248 , n21272 , n21273 );
and ( n21275 , n21161 , n21165 );
and ( n21276 , n21165 , n21170 );
and ( n21277 , n21161 , n21170 );
or ( n21278 , n21275 , n21276 , n21277 );
and ( n21279 , n21176 , n21187 );
and ( n21280 , n21187 , n21202 );
and ( n21281 , n21176 , n21202 );
or ( n21282 , n21279 , n21280 , n21281 );
and ( n21283 , n21278 , n21282 );
and ( n21284 , n21192 , n21196 );
and ( n21285 , n21196 , n21201 );
and ( n21286 , n21192 , n21201 );
or ( n21287 , n21284 , n21285 , n21286 );
buf ( n21288 , n21169 );
xor ( n21289 , n21287 , n21288 );
and ( n21290 , n16058 , n15984 );
xor ( n21291 , n21289 , n21290 );
and ( n21292 , n21282 , n21291 );
and ( n21293 , n21278 , n21291 );
or ( n21294 , n21283 , n21292 , n21293 );
not ( n21295 , n16026 );
and ( n21296 , n16078 , n16102 );
and ( n21297 , n16087 , n16100 );
nor ( n21298 , n21296 , n21297 );
xnor ( n21299 , n21298 , n16110 );
and ( n21300 , n21295 , n21299 );
and ( n21301 , n16096 , n16037 );
and ( n21302 , n16105 , n16035 );
nor ( n21303 , n21301 , n21302 );
xnor ( n21304 , n21303 , n16045 );
and ( n21305 , n21299 , n21304 );
and ( n21306 , n21295 , n21304 );
or ( n21307 , n21300 , n21305 , n21306 );
and ( n21308 , n16008 , n15971 );
and ( n21309 , n16021 , n15969 );
nor ( n21310 , n21308 , n21309 );
xnor ( n21311 , n21310 , n15979 );
and ( n21312 , n15961 , n16055 );
and ( n21313 , n15974 , n16053 );
nor ( n21314 , n21312 , n21313 );
xnor ( n21315 , n21314 , n16063 );
and ( n21316 , n21311 , n21315 );
and ( n21317 , n16029 , n15992 );
and ( n21318 , n16040 , n15990 );
nor ( n21319 , n21317 , n21318 );
xnor ( n21320 , n21319 , n16000 );
and ( n21321 , n21315 , n21320 );
and ( n21322 , n21311 , n21320 );
or ( n21323 , n21316 , n21321 , n21322 );
xor ( n21324 , n21307 , n21323 );
and ( n21325 , n16087 , n16102 );
not ( n21326 , n21325 );
xnor ( n21327 , n21326 , n16110 );
and ( n21328 , n15974 , n16055 );
and ( n21329 , n16096 , n16053 );
nor ( n21330 , n21328 , n21329 );
xnor ( n21331 , n21330 , n16063 );
xor ( n21332 , n21327 , n21331 );
and ( n21333 , n16040 , n15992 );
and ( n21334 , n15961 , n15990 );
nor ( n21335 , n21333 , n21334 );
xnor ( n21336 , n21335 , n16000 );
xor ( n21337 , n21332 , n21336 );
xor ( n21338 , n21324 , n21337 );
xor ( n21339 , n21294 , n21338 );
and ( n21340 , n21287 , n21288 );
and ( n21341 , n21288 , n21290 );
and ( n21342 , n21287 , n21290 );
or ( n21343 , n21340 , n21341 , n21342 );
and ( n21344 , n21180 , n21184 );
and ( n21345 , n21184 , n21186 );
and ( n21346 , n21180 , n21186 );
or ( n21347 , n21344 , n21345 , n21346 );
xor ( n21348 , n21295 , n21299 );
xor ( n21349 , n21348 , n21304 );
and ( n21350 , n21347 , n21349 );
xor ( n21351 , n21311 , n21315 );
xor ( n21352 , n21351 , n21320 );
and ( n21353 , n21349 , n21352 );
and ( n21354 , n21347 , n21352 );
or ( n21355 , n21350 , n21353 , n21354 );
xor ( n21356 , n21343 , n21355 );
and ( n21357 , n16021 , n15971 );
and ( n21358 , n16078 , n15969 );
nor ( n21359 , n21357 , n21358 );
xnor ( n21360 , n21359 , n15979 );
not ( n21361 , n21360 );
and ( n21362 , n16105 , n16037 );
and ( n21363 , n16008 , n16035 );
nor ( n21364 , n21362 , n21363 );
xnor ( n21365 , n21364 , n16045 );
xor ( n21366 , n21361 , n21365 );
and ( n21367 , n16029 , n15984 );
xor ( n21368 , n21366 , n21367 );
xor ( n21369 , n21356 , n21368 );
xor ( n21370 , n21339 , n21369 );
and ( n21371 , n21157 , n21171 );
and ( n21372 , n21171 , n21203 );
and ( n21373 , n21157 , n21203 );
or ( n21374 , n21371 , n21372 , n21373 );
xor ( n21375 , n21347 , n21349 );
xor ( n21376 , n21375 , n21352 );
and ( n21377 , n21374 , n21376 );
xor ( n21378 , n21278 , n21282 );
xor ( n21379 , n21378 , n21291 );
and ( n21380 , n21376 , n21379 );
and ( n21381 , n21374 , n21379 );
or ( n21382 , n21377 , n21380 , n21381 );
xor ( n21383 , n21370 , n21382 );
xor ( n21384 , n21374 , n21376 );
xor ( n21385 , n21384 , n21379 );
and ( n21386 , n21148 , n21152 );
and ( n21387 , n21152 , n21204 );
and ( n21388 , n21148 , n21204 );
or ( n21389 , n21386 , n21387 , n21388 );
and ( n21390 , n21385 , n21389 );
and ( n21391 , n21144 , n21205 );
and ( n21392 , n21205 , n21210 );
and ( n21393 , n21144 , n21210 );
or ( n21394 , n21391 , n21392 , n21393 );
and ( n21395 , n21389 , n21394 );
and ( n21396 , n21385 , n21394 );
or ( n21397 , n21390 , n21395 , n21396 );
xor ( n21398 , n21383 , n21397 );
xor ( n21399 , n21385 , n21389 );
xor ( n21400 , n21399 , n21394 );
and ( n21401 , n21211 , n21212 );
and ( n21402 , n21400 , n21401 );
xor ( n21403 , n21398 , n21402 );
buf ( n21404 , n21403 );
buf ( n21405 , n21404 );
buf ( n21406 , n21405 );
buf ( n21407 , n1181 );
buf ( n21408 , n21407 );
xor ( n21409 , n21136 , n21408 );
buf ( n21410 , n1182 );
buf ( n21411 , n21410 );
xor ( n21412 , n21408 , n21411 );
not ( n21413 , n21412 );
and ( n21414 , n21409 , n21413 );
and ( n21415 , n21406 , n21414 );
and ( n21416 , n21307 , n21323 );
and ( n21417 , n21323 , n21337 );
and ( n21418 , n21307 , n21337 );
or ( n21419 , n21416 , n21417 , n21418 );
and ( n21420 , n21343 , n21355 );
and ( n21421 , n21355 , n21368 );
and ( n21422 , n21343 , n21368 );
or ( n21423 , n21420 , n21421 , n21422 );
xor ( n21424 , n21419 , n21423 );
and ( n21425 , n21361 , n21365 );
and ( n21426 , n21365 , n21367 );
and ( n21427 , n21361 , n21367 );
or ( n21428 , n21425 , n21426 , n21427 );
not ( n21429 , n16110 );
and ( n21430 , n16078 , n15971 );
and ( n21431 , n16087 , n15969 );
nor ( n21432 , n21430 , n21431 );
xnor ( n21433 , n21432 , n15979 );
xor ( n21434 , n21429 , n21433 );
and ( n21435 , n16096 , n16055 );
and ( n21436 , n16105 , n16053 );
nor ( n21437 , n21435 , n21436 );
xnor ( n21438 , n21437 , n16063 );
xor ( n21439 , n21434 , n21438 );
xor ( n21440 , n21428 , n21439 );
and ( n21441 , n21327 , n21331 );
and ( n21442 , n21331 , n21336 );
and ( n21443 , n21327 , n21336 );
or ( n21444 , n21441 , n21442 , n21443 );
buf ( n21445 , n21360 );
xor ( n21446 , n21444 , n21445 );
and ( n21447 , n16008 , n16037 );
and ( n21448 , n16021 , n16035 );
nor ( n21449 , n21447 , n21448 );
xnor ( n21450 , n21449 , n16045 );
and ( n21451 , n15961 , n15992 );
and ( n21452 , n15974 , n15990 );
nor ( n21453 , n21451 , n21452 );
xnor ( n21454 , n21453 , n16000 );
xor ( n21455 , n21450 , n21454 );
and ( n21456 , n16040 , n15984 );
xor ( n21457 , n21455 , n21456 );
xor ( n21458 , n21446 , n21457 );
xor ( n21459 , n21440 , n21458 );
xor ( n21460 , n21424 , n21459 );
and ( n21461 , n21294 , n21338 );
and ( n21462 , n21338 , n21369 );
and ( n21463 , n21294 , n21369 );
or ( n21464 , n21461 , n21462 , n21463 );
xor ( n21465 , n21460 , n21464 );
and ( n21466 , n21370 , n21382 );
and ( n21467 , n21382 , n21397 );
and ( n21468 , n21370 , n21397 );
or ( n21469 , n21466 , n21467 , n21468 );
xor ( n21470 , n21465 , n21469 );
and ( n21471 , n21398 , n21402 );
xor ( n21472 , n21470 , n21471 );
buf ( n21473 , n21472 );
buf ( n21474 , n21473 );
buf ( n21475 , n21474 );
and ( n21476 , n21475 , n21412 );
nor ( n21477 , n21415 , n21476 );
and ( n21478 , n21408 , n21411 );
not ( n21479 , n21478 );
and ( n21480 , n21136 , n21479 );
xnor ( n21481 , n21477 , n21480 );
and ( n21482 , n21274 , n21481 );
xor ( n21483 , n20069 , n21100 );
buf ( n21484 , n21483 );
buf ( n21485 , n21484 );
buf ( n21486 , n21485 );
buf ( n21487 , n1156 );
buf ( n21488 , n21487 );
buf ( n21489 , n1157 );
buf ( n21490 , n21489 );
xor ( n21491 , n21488 , n21490 );
buf ( n21492 , n1158 );
buf ( n21493 , n21492 );
xor ( n21494 , n21490 , n21493 );
not ( n21495 , n21494 );
and ( n21496 , n21491 , n21495 );
and ( n21497 , n21486 , n21496 );
xor ( n21498 , n20067 , n21101 );
buf ( n21499 , n21498 );
buf ( n21500 , n21499 );
buf ( n21501 , n21500 );
and ( n21502 , n21501 , n21494 );
nor ( n21503 , n21497 , n21502 );
and ( n21504 , n21490 , n21493 );
not ( n21505 , n21504 );
and ( n21506 , n21488 , n21505 );
xnor ( n21507 , n21503 , n21506 );
xor ( n21508 , n20118 , n21096 );
buf ( n21509 , n21508 );
buf ( n21510 , n21509 );
buf ( n21511 , n21510 );
buf ( n21512 , n1154 );
buf ( n21513 , n21512 );
and ( n21514 , n21511 , n21513 );
and ( n21515 , n21507 , n21514 );
xor ( n21516 , n19257 , n21107 );
buf ( n21517 , n21516 );
buf ( n21518 , n21517 );
buf ( n21519 , n21518 );
buf ( n21520 , n1160 );
buf ( n21521 , n21520 );
buf ( n21522 , n1161 );
buf ( n21523 , n21522 );
xor ( n21524 , n21521 , n21523 );
buf ( n21525 , n1162 );
buf ( n21526 , n21525 );
xor ( n21527 , n21523 , n21526 );
not ( n21528 , n21527 );
and ( n21529 , n21524 , n21528 );
and ( n21530 , n21519 , n21529 );
xor ( n21531 , n19255 , n21108 );
buf ( n21532 , n21531 );
buf ( n21533 , n21532 );
buf ( n21534 , n21533 );
and ( n21535 , n21534 , n21527 );
nor ( n21536 , n21530 , n21535 );
and ( n21537 , n21523 , n21526 );
not ( n21538 , n21537 );
and ( n21539 , n21521 , n21538 );
xnor ( n21540 , n21536 , n21539 );
and ( n21541 , n21515 , n21540 );
xor ( n21542 , n20071 , n21099 );
buf ( n21543 , n21542 );
buf ( n21544 , n21543 );
buf ( n21545 , n21544 );
buf ( n21546 , n1155 );
buf ( n21547 , n21546 );
xor ( n21548 , n21513 , n21547 );
xor ( n21549 , n21547 , n21488 );
not ( n21550 , n21549 );
and ( n21551 , n21548 , n21550 );
and ( n21552 , n21545 , n21551 );
and ( n21553 , n21486 , n21549 );
nor ( n21554 , n21552 , n21553 );
and ( n21555 , n21547 , n21488 );
not ( n21556 , n21555 );
and ( n21557 , n21513 , n21556 );
xnor ( n21558 , n21554 , n21557 );
and ( n21559 , n21540 , n21558 );
and ( n21560 , n21515 , n21558 );
or ( n21561 , n21541 , n21559 , n21560 );
and ( n21562 , n21241 , n21236 );
xor ( n21563 , n19233 , n21119 );
buf ( n21564 , n21563 );
buf ( n21565 , n21564 );
buf ( n21566 , n21565 );
and ( n21567 , n21566 , n21234 );
nor ( n21568 , n21562 , n21567 );
xnor ( n21569 , n21568 , n21246 );
xor ( n21570 , n21561 , n21569 );
xor ( n21571 , n19243 , n21114 );
buf ( n21572 , n21571 );
buf ( n21573 , n21572 );
buf ( n21574 , n21573 );
buf ( n21575 , n1166 );
buf ( n21576 , n21575 );
buf ( n21577 , n1167 );
buf ( n21578 , n21577 );
xor ( n21579 , n21576 , n21578 );
xor ( n21580 , n21578 , n21254 );
not ( n21581 , n21580 );
and ( n21582 , n21579 , n21581 );
and ( n21583 , n21574 , n21582 );
and ( n21584 , n21252 , n21580 );
nor ( n21585 , n21583 , n21584 );
and ( n21586 , n21578 , n21254 );
not ( n21587 , n21586 );
and ( n21588 , n21576 , n21587 );
xnor ( n21589 , n21585 , n21588 );
xor ( n21590 , n21570 , n21589 );
and ( n21591 , n21481 , n21590 );
and ( n21592 , n21274 , n21590 );
or ( n21593 , n21482 , n21591 , n21592 );
xor ( n21594 , n21507 , n21514 );
and ( n21595 , n21511 , n21551 );
xor ( n21596 , n20073 , n21098 );
buf ( n21597 , n21596 );
buf ( n21598 , n21597 );
buf ( n21599 , n21598 );
and ( n21600 , n21599 , n21549 );
nor ( n21601 , n21595 , n21600 );
xnor ( n21602 , n21601 , n21557 );
xor ( n21603 , n20120 , n21095 );
buf ( n21604 , n21603 );
buf ( n21605 , n21604 );
buf ( n21606 , n21605 );
and ( n21607 , n21606 , n21513 );
xor ( n21608 , n21602 , n21607 );
and ( n21609 , n21606 , n21551 );
and ( n21610 , n21511 , n21549 );
nor ( n21611 , n21609 , n21610 );
xnor ( n21612 , n21611 , n21557 );
xor ( n21613 , n20605 , n21093 );
buf ( n21614 , n21613 );
buf ( n21615 , n21614 );
buf ( n21616 , n21615 );
and ( n21617 , n21616 , n21513 );
and ( n21618 , n21612 , n21617 );
and ( n21619 , n21608 , n21618 );
buf ( n21620 , n1159 );
buf ( n21621 , n21620 );
xor ( n21622 , n21493 , n21621 );
xor ( n21623 , n21621 , n21521 );
not ( n21624 , n21623 );
and ( n21625 , n21622 , n21624 );
and ( n21626 , n21501 , n21625 );
xor ( n21627 , n20065 , n21102 );
buf ( n21628 , n21627 );
buf ( n21629 , n21628 );
buf ( n21630 , n21629 );
and ( n21631 , n21630 , n21623 );
nor ( n21632 , n21626 , n21631 );
and ( n21633 , n21621 , n21521 );
not ( n21634 , n21633 );
and ( n21635 , n21493 , n21634 );
xnor ( n21636 , n21632 , n21635 );
and ( n21637 , n21618 , n21636 );
and ( n21638 , n21608 , n21636 );
or ( n21639 , n21619 , n21637 , n21638 );
and ( n21640 , n21594 , n21639 );
and ( n21641 , n21630 , n21625 );
xor ( n21642 , n19419 , n21104 );
buf ( n21643 , n21642 );
buf ( n21644 , n21643 );
buf ( n21645 , n21644 );
and ( n21646 , n21645 , n21623 );
nor ( n21647 , n21641 , n21646 );
xnor ( n21648 , n21647 , n21635 );
and ( n21649 , n21639 , n21648 );
and ( n21650 , n21594 , n21648 );
or ( n21651 , n21640 , n21649 , n21650 );
xor ( n21652 , n19225 , n21123 );
buf ( n21653 , n21652 );
buf ( n21654 , n21653 );
buf ( n21655 , n21654 );
buf ( n21656 , n1176 );
buf ( n21657 , n21656 );
buf ( n21658 , n1177 );
buf ( n21659 , n21658 );
xor ( n21660 , n21657 , n21659 );
xor ( n21661 , n21659 , n21131 );
not ( n21662 , n21661 );
and ( n21663 , n21660 , n21662 );
and ( n21664 , n21655 , n21663 );
xor ( n21665 , n19223 , n21124 );
buf ( n21666 , n21665 );
buf ( n21667 , n21666 );
buf ( n21668 , n21667 );
and ( n21669 , n21668 , n21661 );
nor ( n21670 , n21664 , n21669 );
and ( n21671 , n21659 , n21131 );
not ( n21672 , n21671 );
and ( n21673 , n21657 , n21672 );
xnor ( n21674 , n21670 , n21673 );
and ( n21675 , n21651 , n21674 );
xor ( n21676 , n19229 , n21121 );
buf ( n21677 , n21676 );
buf ( n21678 , n21677 );
buf ( n21679 , n21678 );
buf ( n21680 , n1174 );
buf ( n21681 , n21680 );
buf ( n21682 , n1175 );
buf ( n21683 , n21682 );
xor ( n21684 , n21681 , n21683 );
xor ( n21685 , n21683 , n21657 );
not ( n21686 , n21685 );
and ( n21687 , n21684 , n21686 );
and ( n21688 , n21679 , n21687 );
xor ( n21689 , n19227 , n21122 );
buf ( n21690 , n21689 );
buf ( n21691 , n21690 );
buf ( n21692 , n21691 );
and ( n21693 , n21692 , n21685 );
nor ( n21694 , n21688 , n21693 );
and ( n21695 , n21683 , n21657 );
not ( n21696 , n21695 );
and ( n21697 , n21681 , n21696 );
xnor ( n21698 , n21694 , n21697 );
and ( n21699 , n21674 , n21698 );
and ( n21700 , n21651 , n21698 );
or ( n21701 , n21675 , n21699 , n21700 );
buf ( n21702 , n1173 );
buf ( n21703 , n21702 );
xor ( n21704 , n21233 , n21703 );
xor ( n21705 , n21703 , n21681 );
not ( n21706 , n21705 );
and ( n21707 , n21704 , n21706 );
and ( n21708 , n21566 , n21707 );
xor ( n21709 , n19231 , n21120 );
buf ( n21710 , n21709 );
buf ( n21711 , n21710 );
buf ( n21712 , n21711 );
and ( n21713 , n21712 , n21705 );
nor ( n21714 , n21708 , n21713 );
and ( n21715 , n21703 , n21681 );
not ( n21716 , n21715 );
and ( n21717 , n21233 , n21716 );
xnor ( n21718 , n21714 , n21717 );
xor ( n21719 , n21515 , n21540 );
xor ( n21720 , n21719 , n21558 );
and ( n21721 , n21718 , n21720 );
and ( n21722 , n21501 , n21496 );
and ( n21723 , n21630 , n21494 );
nor ( n21724 , n21722 , n21723 );
xnor ( n21725 , n21724 , n21506 );
and ( n21726 , n21599 , n21513 );
xor ( n21727 , n21725 , n21726 );
xor ( n21728 , n19253 , n21109 );
buf ( n21729 , n21728 );
buf ( n21730 , n21729 );
buf ( n21731 , n21730 );
buf ( n21732 , n1163 );
buf ( n21733 , n21732 );
xor ( n21734 , n21526 , n21733 );
buf ( n21735 , n1164 );
buf ( n21736 , n21735 );
xor ( n21737 , n21733 , n21736 );
not ( n21738 , n21737 );
and ( n21739 , n21734 , n21738 );
and ( n21740 , n21731 , n21739 );
xor ( n21741 , n19251 , n21110 );
buf ( n21742 , n21741 );
buf ( n21743 , n21742 );
buf ( n21744 , n21743 );
and ( n21745 , n21744 , n21737 );
nor ( n21746 , n21740 , n21745 );
and ( n21747 , n21733 , n21736 );
not ( n21748 , n21747 );
and ( n21749 , n21526 , n21748 );
xnor ( n21750 , n21746 , n21749 );
xor ( n21751 , n21727 , n21750 );
and ( n21752 , n21645 , n21625 );
xor ( n21753 , n19259 , n21106 );
buf ( n21754 , n21753 );
buf ( n21755 , n21754 );
buf ( n21756 , n21755 );
and ( n21757 , n21756 , n21623 );
nor ( n21758 , n21752 , n21757 );
xnor ( n21759 , n21758 , n21635 );
xor ( n21760 , n21751 , n21759 );
and ( n21761 , n21720 , n21760 );
and ( n21762 , n21718 , n21760 );
or ( n21763 , n21721 , n21761 , n21762 );
and ( n21764 , n21701 , n21763 );
and ( n21765 , n21692 , n21687 );
and ( n21766 , n21655 , n21685 );
nor ( n21767 , n21765 , n21766 );
xnor ( n21768 , n21767 , n21697 );
and ( n21769 , n21265 , n21260 );
and ( n21770 , n21226 , n21258 );
nor ( n21771 , n21769 , n21770 );
xnor ( n21772 , n21771 , n21270 );
xor ( n21773 , n21768 , n21772 );
xor ( n21774 , n19247 , n21112 );
buf ( n21775 , n21774 );
buf ( n21776 , n21775 );
buf ( n21777 , n21776 );
buf ( n21778 , n1165 );
buf ( n21779 , n21778 );
xor ( n21780 , n21736 , n21779 );
xor ( n21781 , n21779 , n21576 );
not ( n21782 , n21781 );
and ( n21783 , n21780 , n21782 );
and ( n21784 , n21777 , n21783 );
xor ( n21785 , n19245 , n21113 );
buf ( n21786 , n21785 );
buf ( n21787 , n21786 );
buf ( n21788 , n21787 );
and ( n21789 , n21788 , n21781 );
nor ( n21790 , n21784 , n21789 );
and ( n21791 , n21779 , n21576 );
not ( n21792 , n21791 );
and ( n21793 , n21736 , n21792 );
xnor ( n21794 , n21790 , n21793 );
xor ( n21795 , n21773 , n21794 );
and ( n21796 , n21763 , n21795 );
and ( n21797 , n21701 , n21795 );
or ( n21798 , n21764 , n21796 , n21797 );
and ( n21799 , n21593 , n21798 );
and ( n21800 , n21561 , n21569 );
and ( n21801 , n21569 , n21589 );
and ( n21802 , n21561 , n21589 );
or ( n21803 , n21800 , n21801 , n21802 );
and ( n21804 , n21475 , n21414 );
and ( n21805 , n21444 , n21445 );
and ( n21806 , n21445 , n21457 );
and ( n21807 , n21444 , n21457 );
or ( n21808 , n21805 , n21806 , n21807 );
and ( n21809 , n21428 , n21439 );
and ( n21810 , n21439 , n21458 );
and ( n21811 , n21428 , n21458 );
or ( n21812 , n21809 , n21810 , n21811 );
xor ( n21813 , n21808 , n21812 );
and ( n21814 , n21429 , n21433 );
and ( n21815 , n21433 , n21438 );
and ( n21816 , n21429 , n21438 );
or ( n21817 , n21814 , n21815 , n21816 );
and ( n21818 , n16087 , n15971 );
not ( n21819 , n21818 );
xnor ( n21820 , n21819 , n15979 );
and ( n21821 , n15974 , n15992 );
and ( n21822 , n16096 , n15990 );
nor ( n21823 , n21821 , n21822 );
xnor ( n21824 , n21823 , n16000 );
xor ( n21825 , n21820 , n21824 );
and ( n21826 , n15961 , n15984 );
xor ( n21827 , n21825 , n21826 );
xor ( n21828 , n21817 , n21827 );
and ( n21829 , n21450 , n21454 );
and ( n21830 , n21454 , n21456 );
and ( n21831 , n21450 , n21456 );
or ( n21832 , n21829 , n21830 , n21831 );
and ( n21833 , n16021 , n16037 );
and ( n21834 , n16078 , n16035 );
nor ( n21835 , n21833 , n21834 );
xnor ( n21836 , n21835 , n16045 );
not ( n21837 , n21836 );
xor ( n21838 , n21832 , n21837 );
and ( n21839 , n16105 , n16055 );
and ( n21840 , n16008 , n16053 );
nor ( n21841 , n21839 , n21840 );
xnor ( n21842 , n21841 , n16063 );
xor ( n21843 , n21838 , n21842 );
xor ( n21844 , n21828 , n21843 );
xor ( n21845 , n21813 , n21844 );
and ( n21846 , n21419 , n21423 );
and ( n21847 , n21423 , n21459 );
and ( n21848 , n21419 , n21459 );
or ( n21849 , n21846 , n21847 , n21848 );
xor ( n21850 , n21845 , n21849 );
and ( n21851 , n21460 , n21464 );
and ( n21852 , n21464 , n21469 );
and ( n21853 , n21460 , n21469 );
or ( n21854 , n21851 , n21852 , n21853 );
xor ( n21855 , n21850 , n21854 );
and ( n21856 , n21470 , n21471 );
xor ( n21857 , n21855 , n21856 );
buf ( n21858 , n21857 );
buf ( n21859 , n21858 );
buf ( n21860 , n21859 );
and ( n21861 , n21860 , n21412 );
nor ( n21862 , n21804 , n21861 );
xnor ( n21863 , n21862 , n21480 );
xor ( n21864 , n21803 , n21863 );
and ( n21865 , n21486 , n21551 );
and ( n21866 , n21501 , n21549 );
nor ( n21867 , n21865 , n21866 );
xnor ( n21868 , n21867 , n21557 );
and ( n21869 , n21545 , n21513 );
xor ( n21870 , n21868 , n21869 );
and ( n21871 , n21725 , n21726 );
and ( n21872 , n21870 , n21871 );
and ( n21873 , n21756 , n21625 );
and ( n21874 , n21519 , n21623 );
nor ( n21875 , n21873 , n21874 );
xnor ( n21876 , n21875 , n21635 );
and ( n21877 , n21871 , n21876 );
and ( n21878 , n21870 , n21876 );
or ( n21879 , n21872 , n21877 , n21878 );
and ( n21880 , n21566 , n21236 );
and ( n21881 , n21712 , n21234 );
nor ( n21882 , n21880 , n21881 );
xnor ( n21883 , n21882 , n21246 );
xor ( n21884 , n21879 , n21883 );
and ( n21885 , n21252 , n21582 );
and ( n21886 , n21265 , n21580 );
nor ( n21887 , n21885 , n21886 );
xnor ( n21888 , n21887 , n21588 );
xor ( n21889 , n21884 , n21888 );
xor ( n21890 , n21864 , n21889 );
and ( n21891 , n21798 , n21890 );
and ( n21892 , n21593 , n21890 );
or ( n21893 , n21799 , n21891 , n21892 );
and ( n21894 , n21768 , n21772 );
and ( n21895 , n21772 , n21794 );
and ( n21896 , n21768 , n21794 );
or ( n21897 , n21894 , n21895 , n21896 );
not ( n21898 , n15979 );
and ( n21899 , n16078 , n16037 );
and ( n21900 , n16087 , n16035 );
nor ( n21901 , n21899 , n21900 );
xnor ( n21902 , n21901 , n16045 );
and ( n21903 , n21898 , n21902 );
and ( n21904 , n16096 , n15992 );
and ( n21905 , n16105 , n15990 );
nor ( n21906 , n21904 , n21905 );
xnor ( n21907 , n21906 , n16000 );
and ( n21908 , n21902 , n21907 );
and ( n21909 , n21898 , n21907 );
or ( n21910 , n21903 , n21908 , n21909 );
and ( n21911 , n16087 , n16037 );
not ( n21912 , n21911 );
xnor ( n21913 , n21912 , n16045 );
not ( n21914 , n21913 );
and ( n21915 , n21910 , n21914 );
and ( n21916 , n16021 , n16055 );
and ( n21917 , n16078 , n16053 );
nor ( n21918 , n21916 , n21917 );
xnor ( n21919 , n21918 , n16063 );
and ( n21920 , n16105 , n15992 );
and ( n21921 , n16008 , n15990 );
nor ( n21922 , n21920 , n21921 );
xnor ( n21923 , n21922 , n16000 );
xor ( n21924 , n21919 , n21923 );
and ( n21925 , n16096 , n15984 );
xor ( n21926 , n21924 , n21925 );
and ( n21927 , n21914 , n21926 );
and ( n21928 , n21910 , n21926 );
or ( n21929 , n21915 , n21927 , n21928 );
not ( n21930 , n16045 );
and ( n21931 , n16078 , n16055 );
and ( n21932 , n16087 , n16053 );
nor ( n21933 , n21931 , n21932 );
xnor ( n21934 , n21933 , n16063 );
xor ( n21935 , n21930 , n21934 );
and ( n21936 , n16105 , n15984 );
xor ( n21937 , n21935 , n21936 );
xor ( n21938 , n21929 , n21937 );
and ( n21939 , n21919 , n21923 );
and ( n21940 , n21923 , n21925 );
and ( n21941 , n21919 , n21925 );
or ( n21942 , n21939 , n21940 , n21941 );
buf ( n21943 , n21913 );
xor ( n21944 , n21942 , n21943 );
and ( n21945 , n16008 , n15992 );
and ( n21946 , n16021 , n15990 );
nor ( n21947 , n21945 , n21946 );
xnor ( n21948 , n21947 , n16000 );
xor ( n21949 , n21944 , n21948 );
xor ( n21950 , n21938 , n21949 );
buf ( n21951 , n21836 );
and ( n21952 , n16008 , n16055 );
and ( n21953 , n16021 , n16053 );
nor ( n21954 , n21952 , n21953 );
xnor ( n21955 , n21954 , n16063 );
and ( n21956 , n21951 , n21955 );
and ( n21957 , n15974 , n15984 );
and ( n21958 , n21955 , n21957 );
and ( n21959 , n21951 , n21957 );
or ( n21960 , n21956 , n21958 , n21959 );
and ( n21961 , n21820 , n21824 );
and ( n21962 , n21824 , n21826 );
and ( n21963 , n21820 , n21826 );
or ( n21964 , n21961 , n21962 , n21963 );
xor ( n21965 , n21898 , n21902 );
xor ( n21966 , n21965 , n21907 );
and ( n21967 , n21964 , n21966 );
xor ( n21968 , n21951 , n21955 );
xor ( n21969 , n21968 , n21957 );
and ( n21970 , n21966 , n21969 );
and ( n21971 , n21964 , n21969 );
or ( n21972 , n21967 , n21970 , n21971 );
and ( n21973 , n21960 , n21972 );
xor ( n21974 , n21910 , n21914 );
xor ( n21975 , n21974 , n21926 );
and ( n21976 , n21972 , n21975 );
and ( n21977 , n21960 , n21975 );
or ( n21978 , n21973 , n21976 , n21977 );
xor ( n21979 , n21950 , n21978 );
xor ( n21980 , n21960 , n21972 );
xor ( n21981 , n21980 , n21975 );
and ( n21982 , n21832 , n21837 );
and ( n21983 , n21837 , n21842 );
and ( n21984 , n21832 , n21842 );
or ( n21985 , n21982 , n21983 , n21984 );
and ( n21986 , n21817 , n21827 );
and ( n21987 , n21827 , n21843 );
and ( n21988 , n21817 , n21843 );
or ( n21989 , n21986 , n21987 , n21988 );
and ( n21990 , n21985 , n21989 );
xor ( n21991 , n21964 , n21966 );
xor ( n21992 , n21991 , n21969 );
and ( n21993 , n21989 , n21992 );
and ( n21994 , n21985 , n21992 );
or ( n21995 , n21990 , n21993 , n21994 );
and ( n21996 , n21981 , n21995 );
and ( n21997 , n21808 , n21812 );
and ( n21998 , n21812 , n21844 );
and ( n21999 , n21808 , n21844 );
or ( n22000 , n21997 , n21998 , n21999 );
xor ( n22001 , n21985 , n21989 );
xor ( n22002 , n22001 , n21992 );
and ( n22003 , n22000 , n22002 );
and ( n22004 , n21845 , n21849 );
and ( n22005 , n21849 , n21854 );
and ( n22006 , n21845 , n21854 );
or ( n22007 , n22004 , n22005 , n22006 );
and ( n22008 , n22002 , n22007 );
and ( n22009 , n22000 , n22007 );
or ( n22010 , n22003 , n22008 , n22009 );
and ( n22011 , n21995 , n22010 );
and ( n22012 , n21981 , n22010 );
or ( n22013 , n21996 , n22011 , n22012 );
xor ( n22014 , n21979 , n22013 );
xor ( n22015 , n21981 , n21995 );
xor ( n22016 , n22015 , n22010 );
xor ( n22017 , n22000 , n22002 );
xor ( n22018 , n22017 , n22007 );
and ( n22019 , n21855 , n21856 );
and ( n22020 , n22018 , n22019 );
and ( n22021 , n22016 , n22020 );
xor ( n22022 , n22014 , n22021 );
buf ( n22023 , n22022 );
buf ( n22024 , n22023 );
buf ( n22025 , n22024 );
buf ( n22026 , n1184 );
buf ( n22027 , n22026 );
buf ( n22028 , n1185 );
buf ( n22029 , n22028 );
xor ( n22030 , n22027 , n22029 );
not ( n22031 , n22029 );
and ( n22032 , n22030 , n22031 );
and ( n22033 , n22025 , n22032 );
and ( n22034 , n21930 , n21934 );
and ( n22035 , n21934 , n21936 );
and ( n22036 , n21930 , n21936 );
or ( n22037 , n22034 , n22035 , n22036 );
and ( n22038 , n21942 , n21943 );
and ( n22039 , n21943 , n21948 );
and ( n22040 , n21942 , n21948 );
or ( n22041 , n22038 , n22039 , n22040 );
xor ( n22042 , n22037 , n22041 );
and ( n22043 , n16087 , n16055 );
not ( n22044 , n22043 );
xnor ( n22045 , n22044 , n16063 );
not ( n22046 , n22045 );
and ( n22047 , n16021 , n15992 );
and ( n22048 , n16078 , n15990 );
nor ( n22049 , n22047 , n22048 );
xnor ( n22050 , n22049 , n16000 );
xor ( n22051 , n22046 , n22050 );
and ( n22052 , n16008 , n15984 );
xor ( n22053 , n22051 , n22052 );
xor ( n22054 , n22042 , n22053 );
and ( n22055 , n21929 , n21937 );
and ( n22056 , n21937 , n21949 );
and ( n22057 , n21929 , n21949 );
or ( n22058 , n22055 , n22056 , n22057 );
xor ( n22059 , n22054 , n22058 );
and ( n22060 , n21950 , n21978 );
and ( n22061 , n21978 , n22013 );
and ( n22062 , n21950 , n22013 );
or ( n22063 , n22060 , n22061 , n22062 );
xor ( n22064 , n22059 , n22063 );
and ( n22065 , n22014 , n22021 );
xor ( n22066 , n22064 , n22065 );
buf ( n22067 , n22066 );
buf ( n22068 , n22067 );
buf ( n22069 , n22068 );
and ( n22070 , n22069 , n22029 );
nor ( n22071 , n22033 , n22070 );
xnor ( n22072 , n22071 , n22027 );
and ( n22073 , n21897 , n22072 );
xor ( n22074 , n21400 , n21401 );
buf ( n22075 , n22074 );
buf ( n22076 , n22075 );
buf ( n22077 , n22076 );
and ( n22078 , n22077 , n21139 );
and ( n22079 , n21406 , n21137 );
nor ( n22080 , n22078 , n22079 );
xnor ( n22081 , n22080 , n21221 );
and ( n22082 , n22072 , n22081 );
and ( n22083 , n21897 , n22081 );
or ( n22084 , n22073 , n22082 , n22083 );
and ( n22085 , n21744 , n21739 );
xor ( n22086 , n19249 , n21111 );
buf ( n22087 , n22086 );
buf ( n22088 , n22087 );
buf ( n22089 , n22088 );
and ( n22090 , n22089 , n21737 );
nor ( n22091 , n22085 , n22090 );
xnor ( n22092 , n22091 , n21749 );
and ( n22093 , n21534 , n21529 );
and ( n22094 , n21731 , n21527 );
nor ( n22095 , n22093 , n22094 );
xnor ( n22096 , n22095 , n21539 );
and ( n22097 , n22092 , n22096 );
and ( n22098 , n21630 , n21496 );
and ( n22099 , n21645 , n21494 );
nor ( n22100 , n22098 , n22099 );
xnor ( n22101 , n22100 , n21506 );
and ( n22102 , n22096 , n22101 );
and ( n22103 , n22092 , n22101 );
or ( n22104 , n22097 , n22102 , n22103 );
xor ( n22105 , n22018 , n22019 );
buf ( n22106 , n22105 );
buf ( n22107 , n22106 );
buf ( n22108 , n22107 );
buf ( n22109 , n1183 );
buf ( n22110 , n22109 );
xor ( n22111 , n21411 , n22110 );
xor ( n22112 , n22110 , n22027 );
not ( n22113 , n22112 );
and ( n22114 , n22111 , n22113 );
and ( n22115 , n22108 , n22114 );
xor ( n22116 , n22016 , n22020 );
buf ( n22117 , n22116 );
buf ( n22118 , n22117 );
buf ( n22119 , n22118 );
and ( n22120 , n22119 , n22112 );
nor ( n22121 , n22115 , n22120 );
and ( n22122 , n22110 , n22027 );
not ( n22123 , n22122 );
and ( n22124 , n21411 , n22123 );
xnor ( n22125 , n22121 , n22124 );
and ( n22126 , n22104 , n22125 );
and ( n22127 , n22089 , n21739 );
and ( n22128 , n21777 , n21737 );
nor ( n22129 , n22127 , n22128 );
xnor ( n22130 , n22129 , n21749 );
and ( n22131 , n21731 , n21529 );
and ( n22132 , n21744 , n21527 );
nor ( n22133 , n22131 , n22132 );
xnor ( n22134 , n22133 , n21539 );
xor ( n22135 , n22130 , n22134 );
and ( n22136 , n21645 , n21496 );
and ( n22137 , n21756 , n21494 );
nor ( n22138 , n22136 , n22137 );
xnor ( n22139 , n22138 , n21506 );
xor ( n22140 , n22135 , n22139 );
and ( n22141 , n22125 , n22140 );
and ( n22142 , n22104 , n22140 );
or ( n22143 , n22126 , n22141 , n22142 );
xor ( n22144 , n22084 , n22143 );
and ( n22145 , n22130 , n22134 );
and ( n22146 , n22134 , n22139 );
and ( n22147 , n22130 , n22139 );
or ( n22148 , n22145 , n22146 , n22147 );
and ( n22149 , n21406 , n21139 );
and ( n22150 , n21475 , n21137 );
nor ( n22151 , n22149 , n22150 );
xnor ( n22152 , n22151 , n21221 );
xor ( n22153 , n22148 , n22152 );
and ( n22154 , n21216 , n21663 );
and ( n22155 , n22077 , n21661 );
nor ( n22156 , n22154 , n22155 );
xnor ( n22157 , n22156 , n21673 );
xor ( n22158 , n22153 , n22157 );
xor ( n22159 , n22144 , n22158 );
and ( n22160 , n21893 , n22159 );
and ( n22161 , n21803 , n21863 );
and ( n22162 , n21863 , n21889 );
and ( n22163 , n21803 , n21889 );
or ( n22164 , n22161 , n22162 , n22163 );
and ( n22165 , n21727 , n21750 );
and ( n22166 , n21750 , n21759 );
and ( n22167 , n21727 , n21759 );
or ( n22168 , n22165 , n22166 , n22167 );
and ( n22169 , n21860 , n22114 );
and ( n22170 , n22108 , n22112 );
nor ( n22171 , n22169 , n22170 );
xnor ( n22172 , n22171 , n22124 );
and ( n22173 , n22168 , n22172 );
and ( n22174 , n21668 , n21663 );
and ( n22175 , n21129 , n21661 );
nor ( n22176 , n22174 , n22175 );
xnor ( n22177 , n22176 , n21673 );
and ( n22178 , n22172 , n22177 );
and ( n22179 , n22168 , n22177 );
or ( n22180 , n22173 , n22178 , n22179 );
and ( n22181 , n21129 , n21663 );
and ( n22182 , n21216 , n21661 );
nor ( n22183 , n22181 , n22182 );
xnor ( n22184 , n22183 , n21673 );
and ( n22185 , n21226 , n21260 );
and ( n22186 , n21241 , n21258 );
nor ( n22187 , n22185 , n22186 );
xnor ( n22188 , n22187 , n21270 );
xor ( n22189 , n22184 , n22188 );
and ( n22190 , n21788 , n21783 );
and ( n22191 , n21574 , n21781 );
nor ( n22192 , n22190 , n22191 );
xnor ( n22193 , n22192 , n21793 );
xor ( n22194 , n22189 , n22193 );
and ( n22195 , n22180 , n22194 );
and ( n22196 , n21655 , n21687 );
and ( n22197 , n21668 , n21685 );
nor ( n22198 , n22196 , n22197 );
xnor ( n22199 , n22198 , n21697 );
and ( n22200 , n21679 , n21707 );
and ( n22201 , n21692 , n21705 );
nor ( n22202 , n22200 , n22201 );
xnor ( n22203 , n22202 , n21717 );
xor ( n22204 , n22199 , n22203 );
and ( n22205 , n21501 , n21551 );
and ( n22206 , n21630 , n21549 );
nor ( n22207 , n22205 , n22206 );
xnor ( n22208 , n22207 , n21557 );
and ( n22209 , n21486 , n21513 );
xor ( n22210 , n22208 , n22209 );
and ( n22211 , n21868 , n21869 );
xor ( n22212 , n22210 , n22211 );
and ( n22213 , n21519 , n21625 );
and ( n22214 , n21534 , n21623 );
nor ( n22215 , n22213 , n22214 );
xnor ( n22216 , n22215 , n21635 );
xor ( n22217 , n22212 , n22216 );
xor ( n22218 , n22204 , n22217 );
and ( n22219 , n22194 , n22218 );
and ( n22220 , n22180 , n22218 );
or ( n22221 , n22195 , n22219 , n22220 );
xor ( n22222 , n22164 , n22221 );
and ( n22223 , n22184 , n22188 );
and ( n22224 , n22188 , n22193 );
and ( n22225 , n22184 , n22193 );
or ( n22226 , n22223 , n22224 , n22225 );
and ( n22227 , n21879 , n21883 );
and ( n22228 , n21883 , n21888 );
and ( n22229 , n21879 , n21888 );
or ( n22230 , n22227 , n22228 , n22229 );
xor ( n22231 , n22226 , n22230 );
and ( n22232 , n22119 , n22114 );
and ( n22233 , n22025 , n22112 );
nor ( n22234 , n22232 , n22233 );
xnor ( n22235 , n22234 , n22124 );
xor ( n22236 , n22231 , n22235 );
xor ( n22237 , n22222 , n22236 );
and ( n22238 , n22159 , n22237 );
and ( n22239 , n21893 , n22237 );
or ( n22240 , n22160 , n22238 , n22239 );
and ( n22241 , n21216 , n21139 );
and ( n22242 , n22077 , n21137 );
nor ( n22243 , n22241 , n22242 );
xnor ( n22244 , n22243 , n21221 );
and ( n22245 , n21712 , n21707 );
and ( n22246 , n21679 , n21705 );
nor ( n22247 , n22245 , n22246 );
xnor ( n22248 , n22247 , n21717 );
and ( n22249 , n22244 , n22248 );
xor ( n22250 , n21870 , n21871 );
xor ( n22251 , n22250 , n21876 );
and ( n22252 , n22248 , n22251 );
and ( n22253 , n22244 , n22251 );
or ( n22254 , n22249 , n22252 , n22253 );
and ( n22255 , n21602 , n21607 );
and ( n22256 , n21756 , n21529 );
and ( n22257 , n21519 , n21527 );
nor ( n22258 , n22256 , n22257 );
xnor ( n22259 , n22258 , n21539 );
and ( n22260 , n22255 , n22259 );
and ( n22261 , n21599 , n21551 );
and ( n22262 , n21545 , n21549 );
nor ( n22263 , n22261 , n22262 );
xnor ( n22264 , n22263 , n21557 );
and ( n22265 , n22259 , n22264 );
and ( n22266 , n22255 , n22264 );
or ( n22267 , n22260 , n22265 , n22266 );
and ( n22268 , n21788 , n21582 );
and ( n22269 , n21574 , n21580 );
nor ( n22270 , n22268 , n22269 );
xnor ( n22271 , n22270 , n21588 );
and ( n22272 , n22267 , n22271 );
and ( n22273 , n22089 , n21783 );
and ( n22274 , n21777 , n21781 );
nor ( n22275 , n22273 , n22274 );
xnor ( n22276 , n22275 , n21793 );
and ( n22277 , n22271 , n22276 );
and ( n22278 , n22267 , n22276 );
or ( n22279 , n22272 , n22277 , n22278 );
and ( n22280 , n22119 , n22032 );
and ( n22281 , n22025 , n22029 );
nor ( n22282 , n22280 , n22281 );
xnor ( n22283 , n22282 , n22027 );
and ( n22284 , n22279 , n22283 );
xor ( n22285 , n22092 , n22096 );
xor ( n22286 , n22285 , n22101 );
and ( n22287 , n22283 , n22286 );
and ( n22288 , n22279 , n22286 );
or ( n22289 , n22284 , n22287 , n22288 );
and ( n22290 , n22254 , n22289 );
xor ( n22291 , n22104 , n22125 );
xor ( n22292 , n22291 , n22140 );
and ( n22293 , n22289 , n22292 );
and ( n22294 , n22254 , n22292 );
or ( n22295 , n22290 , n22293 , n22294 );
and ( n22296 , n22199 , n22203 );
and ( n22297 , n22203 , n22217 );
and ( n22298 , n22199 , n22217 );
or ( n22299 , n22296 , n22297 , n22298 );
and ( n22300 , n22069 , n22032 );
and ( n22301 , n22046 , n22050 );
and ( n22302 , n22050 , n22052 );
and ( n22303 , n22046 , n22052 );
or ( n22304 , n22301 , n22302 , n22303 );
buf ( n22305 , n22045 );
xor ( n22306 , n22304 , n22305 );
not ( n22307 , n16063 );
and ( n22308 , n16078 , n15992 );
and ( n22309 , n16087 , n15990 );
nor ( n22310 , n22308 , n22309 );
xnor ( n22311 , n22310 , n16000 );
xor ( n22312 , n22307 , n22311 );
and ( n22313 , n16021 , n15984 );
xor ( n22314 , n22312 , n22313 );
xor ( n22315 , n22306 , n22314 );
and ( n22316 , n22037 , n22041 );
and ( n22317 , n22041 , n22053 );
and ( n22318 , n22037 , n22053 );
or ( n22319 , n22316 , n22317 , n22318 );
xor ( n22320 , n22315 , n22319 );
and ( n22321 , n22054 , n22058 );
and ( n22322 , n22058 , n22063 );
and ( n22323 , n22054 , n22063 );
or ( n22324 , n22321 , n22322 , n22323 );
xor ( n22325 , n22320 , n22324 );
and ( n22326 , n22064 , n22065 );
xor ( n22327 , n22325 , n22326 );
buf ( n22328 , n22327 );
buf ( n22329 , n22328 );
buf ( n22330 , n22329 );
and ( n22331 , n22330 , n22029 );
nor ( n22332 , n22300 , n22331 );
xnor ( n22333 , n22332 , n22027 );
xor ( n22334 , n22299 , n22333 );
and ( n22335 , n21777 , n21739 );
and ( n22336 , n21788 , n21737 );
nor ( n22337 , n22335 , n22336 );
xnor ( n22338 , n22337 , n21749 );
and ( n22339 , n21744 , n21529 );
and ( n22340 , n22089 , n21527 );
nor ( n22341 , n22339 , n22340 );
xnor ( n22342 , n22341 , n21539 );
xor ( n22343 , n22338 , n22342 );
and ( n22344 , n21534 , n21625 );
and ( n22345 , n21731 , n21623 );
nor ( n22346 , n22344 , n22345 );
xnor ( n22347 , n22346 , n21635 );
xor ( n22348 , n22343 , n22347 );
xor ( n22349 , n22334 , n22348 );
and ( n22350 , n22295 , n22349 );
and ( n22351 , n21692 , n21707 );
and ( n22352 , n21655 , n21705 );
nor ( n22353 , n22351 , n22352 );
xnor ( n22354 , n22353 , n21717 );
and ( n22355 , n21712 , n21236 );
and ( n22356 , n21679 , n21234 );
nor ( n22357 , n22355 , n22356 );
xnor ( n22358 , n22357 , n21246 );
xor ( n22359 , n22354 , n22358 );
and ( n22360 , n21574 , n21783 );
and ( n22361 , n21252 , n21781 );
nor ( n22362 , n22360 , n22361 );
xnor ( n22363 , n22362 , n21793 );
xor ( n22364 , n22359 , n22363 );
and ( n22365 , n22210 , n22211 );
and ( n22366 , n22211 , n22216 );
and ( n22367 , n22210 , n22216 );
or ( n22368 , n22365 , n22366 , n22367 );
and ( n22369 , n21241 , n21260 );
and ( n22370 , n21566 , n21258 );
nor ( n22371 , n22369 , n22370 );
xnor ( n22372 , n22371 , n21270 );
xor ( n22373 , n22368 , n22372 );
and ( n22374 , n21265 , n21582 );
and ( n22375 , n21226 , n21580 );
nor ( n22376 , n22374 , n22375 );
xnor ( n22377 , n22376 , n21588 );
xor ( n22378 , n22373 , n22377 );
xor ( n22379 , n22364 , n22378 );
and ( n22380 , n21860 , n21414 );
and ( n22381 , n22108 , n21412 );
nor ( n22382 , n22380 , n22381 );
xnor ( n22383 , n22382 , n21480 );
and ( n22384 , n21668 , n21687 );
and ( n22385 , n21129 , n21685 );
nor ( n22386 , n22384 , n22385 );
xnor ( n22387 , n22386 , n21697 );
xor ( n22388 , n22383 , n22387 );
and ( n22389 , n21756 , n21496 );
and ( n22390 , n21519 , n21494 );
nor ( n22391 , n22389 , n22390 );
xnor ( n22392 , n22391 , n21506 );
and ( n22393 , n21501 , n21513 );
xor ( n22394 , n22392 , n22393 );
and ( n22395 , n22208 , n22209 );
xor ( n22396 , n22394 , n22395 );
and ( n22397 , n21630 , n21551 );
and ( n22398 , n21645 , n21549 );
nor ( n22399 , n22397 , n22398 );
xnor ( n22400 , n22399 , n21557 );
xor ( n22401 , n22396 , n22400 );
xor ( n22402 , n22388 , n22401 );
xor ( n22403 , n22379 , n22402 );
and ( n22404 , n22349 , n22403 );
and ( n22405 , n22295 , n22403 );
or ( n22406 , n22350 , n22404 , n22405 );
and ( n22407 , n22240 , n22406 );
and ( n22408 , n22084 , n22143 );
and ( n22409 , n22143 , n22158 );
and ( n22410 , n22084 , n22158 );
or ( n22411 , n22408 , n22409 , n22410 );
and ( n22412 , n22354 , n22358 );
and ( n22413 , n22358 , n22363 );
and ( n22414 , n22354 , n22363 );
or ( n22415 , n22412 , n22413 , n22414 );
and ( n22416 , n22383 , n22387 );
and ( n22417 , n22387 , n22401 );
and ( n22418 , n22383 , n22401 );
or ( n22419 , n22416 , n22417 , n22418 );
xor ( n22420 , n22415 , n22419 );
and ( n22421 , n21566 , n21260 );
and ( n22422 , n21712 , n21258 );
nor ( n22423 , n22421 , n22422 );
xnor ( n22424 , n22423 , n21270 );
and ( n22425 , n21226 , n21582 );
and ( n22426 , n21241 , n21580 );
nor ( n22427 , n22425 , n22426 );
xnor ( n22428 , n22427 , n21588 );
xor ( n22429 , n22424 , n22428 );
and ( n22430 , n21252 , n21783 );
and ( n22431 , n21265 , n21781 );
nor ( n22432 , n22430 , n22431 );
xnor ( n22433 , n22432 , n21793 );
xor ( n22434 , n22429 , n22433 );
xor ( n22435 , n22420 , n22434 );
xor ( n22436 , n22411 , n22435 );
and ( n22437 , n22148 , n22152 );
and ( n22438 , n22152 , n22157 );
and ( n22439 , n22148 , n22157 );
or ( n22440 , n22437 , n22438 , n22439 );
and ( n22441 , n22330 , n22032 );
and ( n22442 , n22307 , n22311 );
and ( n22443 , n22311 , n22313 );
and ( n22444 , n22307 , n22313 );
or ( n22445 , n22442 , n22443 , n22444 );
and ( n22446 , n16087 , n15992 );
not ( n22447 , n22446 );
xnor ( n22448 , n22447 , n16000 );
xor ( n22449 , n22445 , n22448 );
and ( n22450 , n16078 , n15984 );
not ( n22451 , n22450 );
xor ( n22452 , n22449 , n22451 );
and ( n22453 , n22304 , n22305 );
and ( n22454 , n22305 , n22314 );
and ( n22455 , n22304 , n22314 );
or ( n22456 , n22453 , n22454 , n22455 );
xor ( n22457 , n22452 , n22456 );
and ( n22458 , n22315 , n22319 );
and ( n22459 , n22319 , n22324 );
and ( n22460 , n22315 , n22324 );
or ( n22461 , n22458 , n22459 , n22460 );
xor ( n22462 , n22457 , n22461 );
and ( n22463 , n22325 , n22326 );
xor ( n22464 , n22462 , n22463 );
buf ( n22465 , n22464 );
buf ( n22466 , n22465 );
buf ( n22467 , n22466 );
and ( n22468 , n22467 , n22029 );
nor ( n22469 , n22441 , n22468 );
xnor ( n22470 , n22469 , n22027 );
xor ( n22471 , n22440 , n22470 );
and ( n22472 , n22394 , n22395 );
and ( n22473 , n22395 , n22400 );
and ( n22474 , n22394 , n22400 );
or ( n22475 , n22472 , n22473 , n22474 );
and ( n22476 , n21129 , n21687 );
and ( n22477 , n21216 , n21685 );
nor ( n22478 , n22476 , n22477 );
xnor ( n22479 , n22478 , n21697 );
xor ( n22480 , n22475 , n22479 );
and ( n22481 , n21679 , n21236 );
and ( n22482 , n21692 , n21234 );
nor ( n22483 , n22481 , n22482 );
xnor ( n22484 , n22483 , n21246 );
xor ( n22485 , n22480 , n22484 );
xor ( n22486 , n22471 , n22485 );
xor ( n22487 , n22436 , n22486 );
and ( n22488 , n22406 , n22487 );
and ( n22489 , n22240 , n22487 );
or ( n22490 , n22407 , n22488 , n22489 );
and ( n22491 , n22415 , n22419 );
and ( n22492 , n22419 , n22434 );
and ( n22493 , n22415 , n22434 );
or ( n22494 , n22491 , n22492 , n22493 );
and ( n22495 , n22467 , n22032 );
and ( n22496 , n22445 , n22448 );
and ( n22497 , n22448 , n22451 );
and ( n22498 , n22445 , n22451 );
or ( n22499 , n22496 , n22497 , n22498 );
buf ( n22500 , n22450 );
not ( n22501 , n16000 );
xor ( n22502 , n22500 , n22501 );
and ( n22503 , n16087 , n15984 );
xor ( n22504 , n22502 , n22503 );
xor ( n22505 , n22499 , n22504 );
and ( n22506 , n22452 , n22456 );
and ( n22507 , n22456 , n22461 );
and ( n22508 , n22452 , n22461 );
or ( n22509 , n22506 , n22507 , n22508 );
xor ( n22510 , n22505 , n22509 );
and ( n22511 , n22462 , n22463 );
xor ( n22512 , n22510 , n22511 );
buf ( n22513 , n22512 );
buf ( n22514 , n22513 );
buf ( n22515 , n22514 );
and ( n22516 , n22515 , n22029 );
nor ( n22517 , n22495 , n22516 );
xnor ( n22518 , n22517 , n22027 );
and ( n22519 , n22119 , n21414 );
and ( n22520 , n22025 , n21412 );
nor ( n22521 , n22519 , n22520 );
xnor ( n22522 , n22521 , n21480 );
and ( n22523 , n21406 , n21663 );
and ( n22524 , n21475 , n21661 );
nor ( n22525 , n22523 , n22524 );
xnor ( n22526 , n22525 , n21673 );
xor ( n22527 , n22522 , n22526 );
and ( n22528 , n21519 , n21496 );
and ( n22529 , n21534 , n21494 );
nor ( n22530 , n22528 , n22529 );
xnor ( n22531 , n22530 , n21506 );
and ( n22532 , n21630 , n21513 );
and ( n22533 , n22531 , n22532 );
and ( n22534 , n21534 , n21496 );
and ( n22535 , n21731 , n21494 );
nor ( n22536 , n22534 , n22535 );
xnor ( n22537 , n22536 , n21506 );
xor ( n22538 , n22533 , n22537 );
and ( n22539 , n21756 , n21551 );
and ( n22540 , n21519 , n21549 );
nor ( n22541 , n22539 , n22540 );
xnor ( n22542 , n22541 , n21557 );
xor ( n22543 , n22538 , n22542 );
and ( n22544 , n21645 , n21513 );
xor ( n22545 , n22543 , n22544 );
xor ( n22546 , n22527 , n22545 );
xor ( n22547 , n22518 , n22546 );
and ( n22548 , n22069 , n22114 );
and ( n22549 , n22330 , n22112 );
nor ( n22550 , n22548 , n22549 );
xnor ( n22551 , n22550 , n22124 );
and ( n22552 , n21692 , n21236 );
and ( n22553 , n21655 , n21234 );
nor ( n22554 , n22552 , n22553 );
xnor ( n22555 , n22554 , n21246 );
and ( n22556 , n21265 , n21783 );
and ( n22557 , n21226 , n21781 );
nor ( n22558 , n22556 , n22557 );
xnor ( n22559 , n22558 , n21793 );
xor ( n22560 , n22555 , n22559 );
and ( n22561 , n21574 , n21739 );
and ( n22562 , n21252 , n21737 );
nor ( n22563 , n22561 , n22562 );
xnor ( n22564 , n22563 , n21749 );
xor ( n22565 , n22560 , n22564 );
xor ( n22566 , n22551 , n22565 );
xor ( n22567 , n22531 , n22532 );
and ( n22568 , n22392 , n22393 );
and ( n22569 , n22567 , n22568 );
and ( n22570 , n21645 , n21551 );
and ( n22571 , n21756 , n21549 );
nor ( n22572 , n22570 , n22571 );
xnor ( n22573 , n22572 , n21557 );
and ( n22574 , n22568 , n22573 );
and ( n22575 , n22567 , n22573 );
or ( n22576 , n22569 , n22574 , n22575 );
and ( n22577 , n21860 , n21139 );
and ( n22578 , n22108 , n21137 );
nor ( n22579 , n22577 , n22578 );
xnor ( n22580 , n22579 , n21221 );
xor ( n22581 , n22576 , n22580 );
and ( n22582 , n21712 , n21260 );
and ( n22583 , n21679 , n21258 );
nor ( n22584 , n22582 , n22583 );
xnor ( n22585 , n22584 , n21270 );
xor ( n22586 , n22581 , n22585 );
xor ( n22587 , n22566 , n22586 );
xor ( n22588 , n22547 , n22587 );
xor ( n22589 , n22494 , n22588 );
and ( n22590 , n22475 , n22479 );
and ( n22591 , n22479 , n22484 );
and ( n22592 , n22475 , n22484 );
or ( n22593 , n22590 , n22591 , n22592 );
and ( n22594 , n22364 , n22378 );
and ( n22595 , n22378 , n22402 );
and ( n22596 , n22364 , n22402 );
or ( n22597 , n22594 , n22595 , n22596 );
and ( n22598 , n21475 , n21139 );
and ( n22599 , n21860 , n21137 );
nor ( n22600 , n22598 , n22599 );
xnor ( n22601 , n22600 , n21221 );
and ( n22602 , n22077 , n21663 );
and ( n22603 , n21406 , n21661 );
nor ( n22604 , n22602 , n22603 );
xnor ( n22605 , n22604 , n21673 );
xor ( n22606 , n22601 , n22605 );
xor ( n22607 , n22567 , n22568 );
xor ( n22608 , n22607 , n22573 );
xor ( n22609 , n22606 , n22608 );
and ( n22610 , n22597 , n22609 );
and ( n22611 , n22368 , n22372 );
and ( n22612 , n22372 , n22377 );
and ( n22613 , n22368 , n22377 );
or ( n22614 , n22611 , n22612 , n22613 );
and ( n22615 , n22025 , n22114 );
and ( n22616 , n22069 , n22112 );
nor ( n22617 , n22615 , n22616 );
xnor ( n22618 , n22617 , n22124 );
xor ( n22619 , n22614 , n22618 );
and ( n22620 , n21788 , n21739 );
and ( n22621 , n21574 , n21737 );
nor ( n22622 , n22620 , n22621 );
xnor ( n22623 , n22622 , n21749 );
and ( n22624 , n22089 , n21529 );
and ( n22625 , n21777 , n21527 );
nor ( n22626 , n22624 , n22625 );
xnor ( n22627 , n22626 , n21539 );
xor ( n22628 , n22623 , n22627 );
and ( n22629 , n21731 , n21625 );
and ( n22630 , n21744 , n21623 );
nor ( n22631 , n22629 , n22630 );
xnor ( n22632 , n22631 , n21635 );
xor ( n22633 , n22628 , n22632 );
xor ( n22634 , n22619 , n22633 );
and ( n22635 , n22609 , n22634 );
and ( n22636 , n22597 , n22634 );
or ( n22637 , n22610 , n22635 , n22636 );
xor ( n22638 , n22593 , n22637 );
and ( n22639 , n22614 , n22618 );
and ( n22640 , n22618 , n22633 );
and ( n22641 , n22614 , n22633 );
or ( n22642 , n22639 , n22640 , n22641 );
and ( n22643 , n21241 , n21582 );
and ( n22644 , n21566 , n21580 );
nor ( n22645 , n22643 , n22644 );
xnor ( n22646 , n22645 , n21588 );
xor ( n22647 , n22642 , n22646 );
and ( n22648 , n22424 , n22428 );
and ( n22649 , n22428 , n22433 );
and ( n22650 , n22424 , n22433 );
or ( n22651 , n22648 , n22649 , n22650 );
and ( n22652 , n21777 , n21529 );
and ( n22653 , n21788 , n21527 );
nor ( n22654 , n22652 , n22653 );
xnor ( n22655 , n22654 , n21539 );
xor ( n22656 , n22651 , n22655 );
and ( n22657 , n21744 , n21625 );
and ( n22658 , n22089 , n21623 );
nor ( n22659 , n22657 , n22658 );
xnor ( n22660 , n22659 , n21635 );
xor ( n22661 , n22656 , n22660 );
xor ( n22662 , n22647 , n22661 );
xor ( n22663 , n22638 , n22662 );
xor ( n22664 , n22589 , n22663 );
xor ( n22665 , n22490 , n22664 );
and ( n22666 , n22411 , n22435 );
and ( n22667 , n22435 , n22486 );
and ( n22668 , n22411 , n22486 );
or ( n22669 , n22666 , n22667 , n22668 );
and ( n22670 , n22164 , n22221 );
and ( n22671 , n22221 , n22236 );
and ( n22672 , n22164 , n22236 );
or ( n22673 , n22670 , n22671 , n22672 );
and ( n22674 , n22226 , n22230 );
and ( n22675 , n22230 , n22235 );
and ( n22676 , n22226 , n22235 );
or ( n22677 , n22674 , n22675 , n22676 );
and ( n22678 , n22299 , n22333 );
and ( n22679 , n22333 , n22348 );
and ( n22680 , n22299 , n22348 );
or ( n22681 , n22678 , n22679 , n22680 );
xor ( n22682 , n22677 , n22681 );
and ( n22683 , n22338 , n22342 );
and ( n22684 , n22342 , n22347 );
and ( n22685 , n22338 , n22347 );
or ( n22686 , n22683 , n22684 , n22685 );
and ( n22687 , n22108 , n21414 );
and ( n22688 , n22119 , n21412 );
nor ( n22689 , n22687 , n22688 );
xnor ( n22690 , n22689 , n21480 );
xor ( n22691 , n22686 , n22690 );
and ( n22692 , n21655 , n21707 );
and ( n22693 , n21668 , n21705 );
nor ( n22694 , n22692 , n22693 );
xnor ( n22695 , n22694 , n21717 );
xor ( n22696 , n22691 , n22695 );
xor ( n22697 , n22682 , n22696 );
and ( n22698 , n22673 , n22697 );
xor ( n22699 , n22597 , n22609 );
xor ( n22700 , n22699 , n22634 );
and ( n22701 , n22697 , n22700 );
and ( n22702 , n22673 , n22700 );
or ( n22703 , n22698 , n22701 , n22702 );
xor ( n22704 , n22669 , n22703 );
and ( n22705 , n21692 , n21663 );
and ( n22706 , n21655 , n21661 );
nor ( n22707 , n22705 , n22706 );
xnor ( n22708 , n22707 , n21673 );
and ( n22709 , n21574 , n21260 );
and ( n22710 , n21252 , n21258 );
nor ( n22711 , n22709 , n22710 );
xnor ( n22712 , n22711 , n21270 );
and ( n22713 , n22708 , n22712 );
xor ( n22714 , n22255 , n22259 );
xor ( n22715 , n22714 , n22264 );
and ( n22716 , n22712 , n22715 );
and ( n22717 , n22708 , n22715 );
or ( n22718 , n22713 , n22716 , n22717 );
and ( n22719 , n22077 , n21414 );
and ( n22720 , n21406 , n21412 );
nor ( n22721 , n22719 , n22720 );
xnor ( n22722 , n22721 , n21480 );
and ( n22723 , n22718 , n22722 );
xor ( n22724 , n22267 , n22271 );
xor ( n22725 , n22724 , n22276 );
and ( n22726 , n22722 , n22725 );
and ( n22727 , n22718 , n22725 );
or ( n22728 , n22723 , n22726 , n22727 );
xor ( n22729 , n22168 , n22172 );
xor ( n22730 , n22729 , n22177 );
and ( n22731 , n22728 , n22730 );
xor ( n22732 , n22244 , n22248 );
xor ( n22733 , n22732 , n22251 );
and ( n22734 , n22730 , n22733 );
and ( n22735 , n22728 , n22733 );
or ( n22736 , n22731 , n22734 , n22735 );
xor ( n22737 , n21897 , n22072 );
xor ( n22738 , n22737 , n22081 );
and ( n22739 , n22736 , n22738 );
xor ( n22740 , n22180 , n22194 );
xor ( n22741 , n22740 , n22218 );
and ( n22742 , n22738 , n22741 );
and ( n22743 , n22736 , n22741 );
or ( n22744 , n22739 , n22742 , n22743 );
and ( n22745 , n21777 , n21582 );
and ( n22746 , n21788 , n21580 );
nor ( n22747 , n22745 , n22746 );
xnor ( n22748 , n22747 , n21588 );
and ( n22749 , n21744 , n21783 );
and ( n22750 , n22089 , n21781 );
nor ( n22751 , n22749 , n22750 );
xnor ( n22752 , n22751 , n21793 );
and ( n22753 , n22748 , n22752 );
and ( n22754 , n21534 , n21739 );
and ( n22755 , n21731 , n21737 );
nor ( n22756 , n22754 , n22755 );
xnor ( n22757 , n22756 , n21749 );
and ( n22758 , n22752 , n22757 );
and ( n22759 , n22748 , n22757 );
or ( n22760 , n22753 , n22758 , n22759 );
and ( n22761 , n21519 , n21739 );
and ( n22762 , n21534 , n21737 );
nor ( n22763 , n22761 , n22762 );
xnor ( n22764 , n22763 , n21749 );
and ( n22765 , n21645 , n21529 );
and ( n22766 , n21756 , n21527 );
nor ( n22767 , n22765 , n22766 );
xnor ( n22768 , n22767 , n21539 );
and ( n22769 , n22764 , n22768 );
and ( n22770 , n21545 , n21496 );
and ( n22771 , n21486 , n21494 );
nor ( n22772 , n22770 , n22771 );
xnor ( n22773 , n22772 , n21506 );
and ( n22774 , n22768 , n22773 );
and ( n22775 , n22764 , n22773 );
or ( n22776 , n22769 , n22774 , n22775 );
and ( n22777 , n21241 , n21707 );
and ( n22778 , n21566 , n21705 );
nor ( n22779 , n22777 , n22778 );
xnor ( n22780 , n22779 , n21717 );
and ( n22781 , n22776 , n22780 );
and ( n22782 , n21265 , n21236 );
and ( n22783 , n21226 , n21234 );
nor ( n22784 , n22782 , n22783 );
xnor ( n22785 , n22784 , n21246 );
and ( n22786 , n22780 , n22785 );
and ( n22787 , n22776 , n22785 );
or ( n22788 , n22781 , n22786 , n22787 );
and ( n22789 , n22760 , n22788 );
and ( n22790 , n22108 , n22032 );
and ( n22791 , n22119 , n22029 );
nor ( n22792 , n22790 , n22791 );
xnor ( n22793 , n22792 , n22027 );
and ( n22794 , n22788 , n22793 );
and ( n22795 , n22760 , n22793 );
or ( n22796 , n22789 , n22794 , n22795 );
xor ( n22797 , n22279 , n22283 );
xor ( n22798 , n22797 , n22286 );
and ( n22799 , n22796 , n22798 );
xor ( n22800 , n21274 , n21481 );
xor ( n22801 , n22800 , n21590 );
and ( n22802 , n22798 , n22801 );
and ( n22803 , n22796 , n22801 );
or ( n22804 , n22799 , n22802 , n22803 );
xor ( n22805 , n21612 , n21617 );
and ( n22806 , n21511 , n21496 );
and ( n22807 , n21599 , n21494 );
nor ( n22808 , n22806 , n22807 );
xnor ( n22809 , n22808 , n21506 );
xor ( n22810 , n20607 , n21092 );
buf ( n22811 , n22810 );
buf ( n22812 , n22811 );
buf ( n22813 , n22812 );
and ( n22814 , n22813 , n21513 );
and ( n22815 , n22809 , n22814 );
and ( n22816 , n22805 , n22815 );
and ( n22817 , n21486 , n21625 );
and ( n22818 , n21501 , n21623 );
nor ( n22819 , n22817 , n22818 );
xnor ( n22820 , n22819 , n21635 );
and ( n22821 , n22815 , n22820 );
and ( n22822 , n22805 , n22820 );
or ( n22823 , n22816 , n22821 , n22822 );
and ( n22824 , n21788 , n21260 );
and ( n22825 , n21574 , n21258 );
nor ( n22826 , n22824 , n22825 );
xnor ( n22827 , n22826 , n21270 );
and ( n22828 , n22823 , n22827 );
and ( n22829 , n21731 , n21783 );
and ( n22830 , n21744 , n21781 );
nor ( n22831 , n22829 , n22830 );
xnor ( n22832 , n22831 , n21793 );
and ( n22833 , n22827 , n22832 );
and ( n22834 , n22823 , n22832 );
or ( n22835 , n22828 , n22833 , n22834 );
and ( n22836 , n21216 , n21414 );
and ( n22837 , n22077 , n21412 );
nor ( n22838 , n22836 , n22837 );
xnor ( n22839 , n22838 , n21480 );
and ( n22840 , n22835 , n22839 );
and ( n22841 , n21712 , n21687 );
and ( n22842 , n21679 , n21685 );
nor ( n22843 , n22841 , n22842 );
xnor ( n22844 , n22843 , n21697 );
and ( n22845 , n22839 , n22844 );
and ( n22846 , n22835 , n22844 );
or ( n22847 , n22840 , n22845 , n22846 );
xor ( n22848 , n21222 , n21247 );
xor ( n22849 , n22848 , n21271 );
and ( n22850 , n22847 , n22849 );
xor ( n22851 , n21651 , n21674 );
xor ( n22852 , n22851 , n21698 );
and ( n22853 , n22849 , n22852 );
and ( n22854 , n22847 , n22852 );
or ( n22855 , n22850 , n22853 , n22854 );
and ( n22856 , n21860 , n22032 );
and ( n22857 , n22108 , n22029 );
nor ( n22858 , n22856 , n22857 );
xnor ( n22859 , n22858 , n22027 );
and ( n22860 , n21668 , n21139 );
and ( n22861 , n21129 , n21137 );
nor ( n22862 , n22860 , n22861 );
xnor ( n22863 , n22862 , n21221 );
and ( n22864 , n22859 , n22863 );
xor ( n22865 , n21594 , n21639 );
xor ( n22866 , n22865 , n21648 );
and ( n22867 , n22863 , n22866 );
and ( n22868 , n22859 , n22866 );
or ( n22869 , n22864 , n22867 , n22868 );
and ( n22870 , n21475 , n22114 );
and ( n22871 , n21860 , n22112 );
nor ( n22872 , n22870 , n22871 );
xnor ( n22873 , n22872 , n22124 );
and ( n22874 , n22869 , n22873 );
xor ( n22875 , n21718 , n21720 );
xor ( n22876 , n22875 , n21760 );
and ( n22877 , n22873 , n22876 );
and ( n22878 , n22869 , n22876 );
or ( n22879 , n22874 , n22877 , n22878 );
and ( n22880 , n22855 , n22879 );
xor ( n22881 , n21701 , n21763 );
xor ( n22882 , n22881 , n21795 );
and ( n22883 , n22879 , n22882 );
and ( n22884 , n22855 , n22882 );
or ( n22885 , n22880 , n22883 , n22884 );
and ( n22886 , n22804 , n22885 );
xor ( n22887 , n22254 , n22289 );
xor ( n22888 , n22887 , n22292 );
and ( n22889 , n22885 , n22888 );
and ( n22890 , n22804 , n22888 );
or ( n22891 , n22886 , n22889 , n22890 );
and ( n22892 , n22744 , n22891 );
xor ( n22893 , n22295 , n22349 );
xor ( n22894 , n22893 , n22403 );
and ( n22895 , n22891 , n22894 );
and ( n22896 , n22744 , n22894 );
or ( n22897 , n22892 , n22895 , n22896 );
xor ( n22898 , n22673 , n22697 );
xor ( n22899 , n22898 , n22700 );
and ( n22900 , n22897 , n22899 );
xor ( n22901 , n22240 , n22406 );
xor ( n22902 , n22901 , n22487 );
and ( n22903 , n22899 , n22902 );
and ( n22904 , n22897 , n22902 );
or ( n22905 , n22900 , n22903 , n22904 );
xor ( n22906 , n22704 , n22905 );
and ( n22907 , n22440 , n22470 );
and ( n22908 , n22470 , n22485 );
and ( n22909 , n22440 , n22485 );
or ( n22910 , n22907 , n22908 , n22909 );
and ( n22911 , n22677 , n22681 );
and ( n22912 , n22681 , n22696 );
and ( n22913 , n22677 , n22696 );
or ( n22914 , n22911 , n22912 , n22913 );
xor ( n22915 , n22910 , n22914 );
and ( n22916 , n22686 , n22690 );
and ( n22917 , n22690 , n22695 );
and ( n22918 , n22686 , n22695 );
or ( n22919 , n22916 , n22917 , n22918 );
and ( n22920 , n22601 , n22605 );
and ( n22921 , n22605 , n22608 );
and ( n22922 , n22601 , n22608 );
or ( n22923 , n22920 , n22921 , n22922 );
xor ( n22924 , n22919 , n22923 );
and ( n22925 , n22623 , n22627 );
and ( n22926 , n22627 , n22632 );
and ( n22927 , n22623 , n22632 );
or ( n22928 , n22925 , n22926 , n22927 );
and ( n22929 , n21216 , n21687 );
and ( n22930 , n22077 , n21685 );
nor ( n22931 , n22929 , n22930 );
xnor ( n22932 , n22931 , n21697 );
xor ( n22933 , n22928 , n22932 );
and ( n22934 , n21668 , n21707 );
and ( n22935 , n21129 , n21705 );
nor ( n22936 , n22934 , n22935 );
xnor ( n22937 , n22936 , n21717 );
xor ( n22938 , n22933 , n22937 );
xor ( n22939 , n22924 , n22938 );
xor ( n22940 , n22915 , n22939 );
xor ( n22941 , n22906 , n22940 );
xor ( n22942 , n22665 , n22941 );
xor ( n22943 , n22897 , n22899 );
xor ( n22944 , n22943 , n22902 );
and ( n22945 , n21252 , n21236 );
and ( n22946 , n21265 , n21234 );
nor ( n22947 , n22945 , n22946 );
xnor ( n22948 , n22947 , n21246 );
and ( n22949 , n22089 , n21582 );
and ( n22950 , n21777 , n21580 );
nor ( n22951 , n22949 , n22950 );
xnor ( n22952 , n22951 , n21588 );
and ( n22953 , n22948 , n22952 );
xor ( n22954 , n21608 , n21618 );
xor ( n22955 , n22954 , n21636 );
and ( n22956 , n22952 , n22955 );
and ( n22957 , n22948 , n22955 );
or ( n22958 , n22953 , n22956 , n22957 );
and ( n22959 , n21406 , n22114 );
and ( n22960 , n21475 , n22112 );
nor ( n22961 , n22959 , n22960 );
xnor ( n22962 , n22961 , n22124 );
and ( n22963 , n22958 , n22962 );
xor ( n22964 , n22748 , n22752 );
xor ( n22965 , n22964 , n22757 );
and ( n22966 , n22962 , n22965 );
and ( n22967 , n22958 , n22965 );
or ( n22968 , n22963 , n22966 , n22967 );
xor ( n22969 , n22760 , n22788 );
xor ( n22970 , n22969 , n22793 );
and ( n22971 , n22968 , n22970 );
xor ( n22972 , n22718 , n22722 );
xor ( n22973 , n22972 , n22725 );
and ( n22974 , n22970 , n22973 );
and ( n22975 , n22968 , n22973 );
or ( n22976 , n22971 , n22974 , n22975 );
xor ( n22977 , n22728 , n22730 );
xor ( n22978 , n22977 , n22733 );
and ( n22979 , n22976 , n22978 );
xor ( n22980 , n22796 , n22798 );
xor ( n22981 , n22980 , n22801 );
and ( n22982 , n22978 , n22981 );
and ( n22983 , n22976 , n22981 );
or ( n22984 , n22979 , n22982 , n22983 );
xor ( n22985 , n21593 , n21798 );
xor ( n22986 , n22985 , n21890 );
and ( n22987 , n22984 , n22986 );
xor ( n22988 , n22736 , n22738 );
xor ( n22989 , n22988 , n22741 );
and ( n22990 , n22986 , n22989 );
and ( n22991 , n22984 , n22989 );
or ( n22992 , n22987 , n22990 , n22991 );
xor ( n22993 , n21893 , n22159 );
xor ( n22994 , n22993 , n22237 );
and ( n22995 , n22992 , n22994 );
xor ( n22996 , n22744 , n22891 );
xor ( n22997 , n22996 , n22894 );
and ( n22998 , n22994 , n22997 );
and ( n22999 , n22992 , n22997 );
or ( n23000 , n22995 , n22998 , n22999 );
and ( n23001 , n22944 , n23000 );
and ( n23002 , n22077 , n22114 );
and ( n23003 , n21406 , n22112 );
nor ( n23004 , n23002 , n23003 );
xnor ( n23005 , n23004 , n22124 );
xor ( n23006 , n22823 , n22827 );
xor ( n23007 , n23006 , n22832 );
and ( n23008 , n23005 , n23007 );
xor ( n23009 , n22948 , n22952 );
xor ( n23010 , n23009 , n22955 );
and ( n23011 , n23007 , n23010 );
and ( n23012 , n23005 , n23010 );
or ( n23013 , n23008 , n23011 , n23012 );
xor ( n23014 , n22835 , n22839 );
xor ( n23015 , n23014 , n22844 );
and ( n23016 , n23013 , n23015 );
xor ( n23017 , n22958 , n22962 );
xor ( n23018 , n23017 , n22965 );
and ( n23019 , n23015 , n23018 );
and ( n23020 , n23013 , n23018 );
or ( n23021 , n23016 , n23019 , n23020 );
xor ( n23022 , n22847 , n22849 );
xor ( n23023 , n23022 , n22852 );
and ( n23024 , n23021 , n23023 );
xor ( n23025 , n22968 , n22970 );
xor ( n23026 , n23025 , n22973 );
and ( n23027 , n23023 , n23026 );
and ( n23028 , n23021 , n23026 );
or ( n23029 , n23024 , n23027 , n23028 );
and ( n23030 , n21756 , n21739 );
and ( n23031 , n21519 , n21737 );
nor ( n23032 , n23030 , n23031 );
xnor ( n23033 , n23032 , n21749 );
and ( n23034 , n21630 , n21529 );
and ( n23035 , n21645 , n21527 );
nor ( n23036 , n23034 , n23035 );
xnor ( n23037 , n23036 , n21539 );
and ( n23038 , n23033 , n23037 );
and ( n23039 , n21599 , n21496 );
and ( n23040 , n21545 , n21494 );
nor ( n23041 , n23039 , n23040 );
xnor ( n23042 , n23041 , n21506 );
and ( n23043 , n23037 , n23042 );
and ( n23044 , n23033 , n23042 );
or ( n23045 , n23038 , n23043 , n23044 );
and ( n23046 , n21129 , n21414 );
and ( n23047 , n21216 , n21412 );
nor ( n23048 , n23046 , n23047 );
xnor ( n23049 , n23048 , n21480 );
and ( n23050 , n23045 , n23049 );
and ( n23051 , n21566 , n21687 );
and ( n23052 , n21712 , n21685 );
nor ( n23053 , n23051 , n23052 );
xnor ( n23054 , n23053 , n21697 );
and ( n23055 , n23049 , n23054 );
and ( n23056 , n23045 , n23054 );
or ( n23057 , n23050 , n23055 , n23056 );
xor ( n23058 , n22776 , n22780 );
xor ( n23059 , n23058 , n22785 );
and ( n23060 , n23057 , n23059 );
xor ( n23061 , n22708 , n22712 );
xor ( n23062 , n23061 , n22715 );
and ( n23063 , n23059 , n23062 );
and ( n23064 , n23057 , n23062 );
or ( n23065 , n23060 , n23063 , n23064 );
xor ( n23066 , n22809 , n22814 );
and ( n23067 , n21606 , n21496 );
and ( n23068 , n21511 , n21494 );
nor ( n23069 , n23067 , n23068 );
xnor ( n23070 , n23069 , n21506 );
xor ( n23071 , n20609 , n21091 );
buf ( n23072 , n23071 );
buf ( n23073 , n23072 );
buf ( n23074 , n23073 );
and ( n23075 , n23074 , n21513 );
and ( n23076 , n23070 , n23075 );
and ( n23077 , n23066 , n23076 );
and ( n23078 , n21616 , n21551 );
and ( n23079 , n21606 , n21549 );
nor ( n23080 , n23078 , n23079 );
xnor ( n23081 , n23080 , n21557 );
and ( n23082 , n23076 , n23081 );
and ( n23083 , n23066 , n23081 );
or ( n23084 , n23077 , n23082 , n23083 );
and ( n23085 , n21777 , n21260 );
and ( n23086 , n21788 , n21258 );
nor ( n23087 , n23085 , n23086 );
xnor ( n23088 , n23087 , n21270 );
and ( n23089 , n23084 , n23088 );
and ( n23090 , n21534 , n21783 );
and ( n23091 , n21731 , n21781 );
nor ( n23092 , n23090 , n23091 );
xnor ( n23093 , n23092 , n21793 );
and ( n23094 , n23088 , n23093 );
and ( n23095 , n23084 , n23093 );
or ( n23096 , n23089 , n23094 , n23095 );
and ( n23097 , n21519 , n21783 );
and ( n23098 , n21534 , n21781 );
nor ( n23099 , n23097 , n23098 );
xnor ( n23100 , n23099 , n21793 );
and ( n23101 , n21501 , n21529 );
and ( n23102 , n21630 , n21527 );
nor ( n23103 , n23101 , n23102 );
xnor ( n23104 , n23103 , n21539 );
and ( n23105 , n23100 , n23104 );
and ( n23106 , n21545 , n21625 );
and ( n23107 , n21486 , n21623 );
nor ( n23108 , n23106 , n23107 );
xnor ( n23109 , n23108 , n21635 );
and ( n23110 , n23104 , n23109 );
and ( n23111 , n23100 , n23109 );
or ( n23112 , n23105 , n23110 , n23111 );
and ( n23113 , n21744 , n21582 );
and ( n23114 , n22089 , n21580 );
nor ( n23115 , n23113 , n23114 );
xnor ( n23116 , n23115 , n21588 );
and ( n23117 , n23112 , n23116 );
xor ( n23118 , n22805 , n22815 );
xor ( n23119 , n23118 , n22820 );
and ( n23120 , n23116 , n23119 );
and ( n23121 , n23112 , n23119 );
or ( n23122 , n23117 , n23120 , n23121 );
and ( n23123 , n23096 , n23122 );
and ( n23124 , n21679 , n21663 );
and ( n23125 , n21692 , n21661 );
nor ( n23126 , n23124 , n23125 );
xnor ( n23127 , n23126 , n21673 );
and ( n23128 , n23122 , n23127 );
and ( n23129 , n23096 , n23127 );
or ( n23130 , n23123 , n23128 , n23129 );
and ( n23131 , n21655 , n21139 );
and ( n23132 , n21668 , n21137 );
nor ( n23133 , n23131 , n23132 );
xnor ( n23134 , n23133 , n21221 );
and ( n23135 , n21226 , n21707 );
and ( n23136 , n21241 , n21705 );
nor ( n23137 , n23135 , n23136 );
xnor ( n23138 , n23137 , n21717 );
and ( n23139 , n23134 , n23138 );
xor ( n23140 , n22764 , n22768 );
xor ( n23141 , n23140 , n22773 );
and ( n23142 , n23138 , n23141 );
and ( n23143 , n23134 , n23141 );
or ( n23144 , n23139 , n23142 , n23143 );
and ( n23145 , n23130 , n23144 );
xor ( n23146 , n22859 , n22863 );
xor ( n23147 , n23146 , n22866 );
and ( n23148 , n23144 , n23147 );
and ( n23149 , n23130 , n23147 );
or ( n23150 , n23145 , n23148 , n23149 );
and ( n23151 , n23065 , n23150 );
xor ( n23152 , n22869 , n22873 );
xor ( n23153 , n23152 , n22876 );
and ( n23154 , n23150 , n23153 );
and ( n23155 , n23065 , n23153 );
or ( n23156 , n23151 , n23154 , n23155 );
and ( n23157 , n23029 , n23156 );
xor ( n23158 , n22855 , n22879 );
xor ( n23159 , n23158 , n22882 );
and ( n23160 , n23156 , n23159 );
and ( n23161 , n23029 , n23159 );
or ( n23162 , n23157 , n23160 , n23161 );
xor ( n23163 , n22804 , n22885 );
xor ( n23164 , n23163 , n22888 );
and ( n23165 , n23162 , n23164 );
xor ( n23166 , n22984 , n22986 );
xor ( n23167 , n23166 , n22989 );
and ( n23168 , n23164 , n23167 );
and ( n23169 , n23162 , n23167 );
or ( n23170 , n23165 , n23168 , n23169 );
xor ( n23171 , n22992 , n22994 );
xor ( n23172 , n23171 , n22997 );
and ( n23173 , n23170 , n23172 );
xor ( n23174 , n23162 , n23164 );
xor ( n23175 , n23174 , n23167 );
and ( n23176 , n21566 , n21663 );
and ( n23177 , n21712 , n21661 );
nor ( n23178 , n23176 , n23177 );
xnor ( n23179 , n23178 , n21673 );
and ( n23180 , n21226 , n21687 );
and ( n23181 , n21241 , n21685 );
nor ( n23182 , n23180 , n23181 );
xnor ( n23183 , n23182 , n21697 );
and ( n23184 , n23179 , n23183 );
and ( n23185 , n21252 , n21707 );
and ( n23186 , n21265 , n21705 );
nor ( n23187 , n23185 , n23186 );
xnor ( n23188 , n23187 , n21717 );
and ( n23189 , n23183 , n23188 );
and ( n23190 , n23179 , n23188 );
or ( n23191 , n23184 , n23189 , n23190 );
and ( n23192 , n21129 , n22114 );
and ( n23193 , n21216 , n22112 );
nor ( n23194 , n23192 , n23193 );
xnor ( n23195 , n23194 , n22124 );
xor ( n23196 , n23100 , n23104 );
xor ( n23197 , n23196 , n23109 );
and ( n23198 , n23195 , n23197 );
xor ( n23199 , n23066 , n23076 );
xor ( n23200 , n23199 , n23081 );
and ( n23201 , n23197 , n23200 );
and ( n23202 , n23195 , n23200 );
or ( n23203 , n23198 , n23201 , n23202 );
and ( n23204 , n23191 , n23203 );
and ( n23205 , n21406 , n22032 );
and ( n23206 , n21475 , n22029 );
nor ( n23207 , n23205 , n23206 );
xnor ( n23208 , n23207 , n22027 );
and ( n23209 , n23203 , n23208 );
and ( n23210 , n23191 , n23208 );
or ( n23211 , n23204 , n23209 , n23210 );
and ( n23212 , n21216 , n22114 );
and ( n23213 , n22077 , n22112 );
nor ( n23214 , n23212 , n23213 );
xnor ( n23215 , n23214 , n22124 );
xor ( n23216 , n23084 , n23088 );
xor ( n23217 , n23216 , n23093 );
and ( n23218 , n23215 , n23217 );
xor ( n23219 , n23112 , n23116 );
xor ( n23220 , n23219 , n23119 );
and ( n23221 , n23217 , n23220 );
and ( n23222 , n23215 , n23220 );
or ( n23223 , n23218 , n23221 , n23222 );
and ( n23224 , n23211 , n23223 );
xor ( n23225 , n23096 , n23122 );
xor ( n23226 , n23225 , n23127 );
and ( n23227 , n23223 , n23226 );
and ( n23228 , n23211 , n23226 );
or ( n23229 , n23224 , n23227 , n23228 );
and ( n23230 , n21534 , n21582 );
and ( n23231 , n21731 , n21580 );
nor ( n23232 , n23230 , n23231 );
xnor ( n23233 , n23232 , n21588 );
and ( n23234 , n21756 , n21783 );
and ( n23235 , n21519 , n21781 );
nor ( n23236 , n23234 , n23235 );
xnor ( n23237 , n23236 , n21793 );
and ( n23238 , n23233 , n23237 );
and ( n23239 , n21630 , n21739 );
and ( n23240 , n21645 , n21737 );
nor ( n23241 , n23239 , n23240 );
xnor ( n23242 , n23241 , n21749 );
and ( n23243 , n23237 , n23242 );
and ( n23244 , n23233 , n23242 );
or ( n23245 , n23238 , n23243 , n23244 );
and ( n23246 , n21655 , n21414 );
and ( n23247 , n21668 , n21412 );
nor ( n23248 , n23246 , n23247 );
xnor ( n23249 , n23248 , n21480 );
and ( n23250 , n23245 , n23249 );
and ( n23251 , n21679 , n21139 );
and ( n23252 , n21692 , n21137 );
nor ( n23253 , n23251 , n23252 );
xnor ( n23254 , n23253 , n21221 );
and ( n23255 , n23249 , n23254 );
and ( n23256 , n23245 , n23254 );
or ( n23257 , n23250 , n23255 , n23256 );
and ( n23258 , n21692 , n21139 );
and ( n23259 , n21655 , n21137 );
nor ( n23260 , n23258 , n23259 );
xnor ( n23261 , n23260 , n21221 );
and ( n23262 , n21241 , n21687 );
and ( n23263 , n21566 , n21685 );
nor ( n23264 , n23262 , n23263 );
xnor ( n23265 , n23264 , n21697 );
xor ( n23266 , n23261 , n23265 );
and ( n23267 , n21574 , n21236 );
and ( n23268 , n21252 , n21234 );
nor ( n23269 , n23267 , n23268 );
xnor ( n23270 , n23269 , n21246 );
xor ( n23271 , n23266 , n23270 );
and ( n23272 , n23257 , n23271 );
and ( n23273 , n21668 , n21414 );
and ( n23274 , n21129 , n21412 );
nor ( n23275 , n23273 , n23274 );
xnor ( n23276 , n23275 , n21480 );
and ( n23277 , n21265 , n21707 );
and ( n23278 , n21226 , n21705 );
nor ( n23279 , n23277 , n23278 );
xnor ( n23280 , n23279 , n21717 );
xor ( n23281 , n23276 , n23280 );
xor ( n23282 , n23033 , n23037 );
xor ( n23283 , n23282 , n23042 );
xor ( n23284 , n23281 , n23283 );
and ( n23285 , n23271 , n23284 );
and ( n23286 , n23257 , n23284 );
or ( n23287 , n23272 , n23285 , n23286 );
and ( n23288 , n23261 , n23265 );
and ( n23289 , n23265 , n23270 );
and ( n23290 , n23261 , n23270 );
or ( n23291 , n23288 , n23289 , n23290 );
and ( n23292 , n21475 , n22032 );
and ( n23293 , n21860 , n22029 );
nor ( n23294 , n23292 , n23293 );
xnor ( n23295 , n23294 , n22027 );
xor ( n23296 , n23291 , n23295 );
xor ( n23297 , n23134 , n23138 );
xor ( n23298 , n23297 , n23141 );
xor ( n23299 , n23296 , n23298 );
and ( n23300 , n23287 , n23299 );
xor ( n23301 , n23005 , n23007 );
xor ( n23302 , n23301 , n23010 );
and ( n23303 , n23299 , n23302 );
and ( n23304 , n23287 , n23302 );
or ( n23305 , n23300 , n23303 , n23304 );
and ( n23306 , n23229 , n23305 );
xor ( n23307 , n23130 , n23144 );
xor ( n23308 , n23307 , n23147 );
and ( n23309 , n23305 , n23308 );
and ( n23310 , n23229 , n23308 );
or ( n23311 , n23306 , n23309 , n23310 );
xor ( n23312 , n23070 , n23075 );
and ( n23313 , n23074 , n21551 );
and ( n23314 , n22813 , n21549 );
nor ( n23315 , n23313 , n23314 );
xnor ( n23316 , n23315 , n21557 );
xor ( n23317 , n20611 , n21090 );
buf ( n23318 , n23317 );
buf ( n23319 , n23318 );
buf ( n23320 , n23319 );
and ( n23321 , n23320 , n21513 );
and ( n23322 , n23316 , n23321 );
and ( n23323 , n23312 , n23322 );
and ( n23324 , n22813 , n21551 );
and ( n23325 , n21616 , n21549 );
nor ( n23326 , n23324 , n23325 );
xnor ( n23327 , n23326 , n21557 );
and ( n23328 , n23322 , n23327 );
and ( n23329 , n23312 , n23327 );
or ( n23330 , n23323 , n23328 , n23329 );
and ( n23331 , n21731 , n21582 );
and ( n23332 , n21744 , n21580 );
nor ( n23333 , n23331 , n23332 );
xnor ( n23334 , n23333 , n21588 );
and ( n23335 , n23330 , n23334 );
and ( n23336 , n21645 , n21739 );
and ( n23337 , n21756 , n21737 );
nor ( n23338 , n23336 , n23337 );
xnor ( n23339 , n23338 , n21749 );
and ( n23340 , n23334 , n23339 );
and ( n23341 , n23330 , n23339 );
or ( n23342 , n23335 , n23340 , n23341 );
xor ( n23343 , n23316 , n23321 );
and ( n23344 , n23320 , n21551 );
and ( n23345 , n23074 , n21549 );
nor ( n23346 , n23344 , n23345 );
xnor ( n23347 , n23346 , n21557 );
xor ( n23348 , n20613 , n21089 );
buf ( n23349 , n23348 );
buf ( n23350 , n23349 );
buf ( n23351 , n23350 );
and ( n23352 , n23351 , n21513 );
and ( n23353 , n23347 , n23352 );
and ( n23354 , n23343 , n23353 );
and ( n23355 , n21511 , n21625 );
and ( n23356 , n21599 , n21623 );
nor ( n23357 , n23355 , n23356 );
xnor ( n23358 , n23357 , n21635 );
and ( n23359 , n23353 , n23358 );
and ( n23360 , n23343 , n23358 );
or ( n23361 , n23354 , n23359 , n23360 );
and ( n23362 , n21486 , n21529 );
and ( n23363 , n21501 , n21527 );
nor ( n23364 , n23362 , n23363 );
xnor ( n23365 , n23364 , n21539 );
and ( n23366 , n23361 , n23365 );
and ( n23367 , n21599 , n21625 );
and ( n23368 , n21545 , n21623 );
nor ( n23369 , n23367 , n23368 );
xnor ( n23370 , n23369 , n21635 );
and ( n23371 , n23365 , n23370 );
and ( n23372 , n23361 , n23370 );
or ( n23373 , n23366 , n23371 , n23372 );
and ( n23374 , n21788 , n21236 );
and ( n23375 , n21574 , n21234 );
nor ( n23376 , n23374 , n23375 );
xnor ( n23377 , n23376 , n21246 );
and ( n23378 , n23373 , n23377 );
and ( n23379 , n22089 , n21260 );
and ( n23380 , n21777 , n21258 );
nor ( n23381 , n23379 , n23380 );
xnor ( n23382 , n23381 , n21270 );
and ( n23383 , n23377 , n23382 );
and ( n23384 , n23373 , n23382 );
or ( n23385 , n23378 , n23383 , n23384 );
and ( n23386 , n23342 , n23385 );
and ( n23387 , n21712 , n21663 );
and ( n23388 , n21679 , n21661 );
nor ( n23389 , n23387 , n23388 );
xnor ( n23390 , n23389 , n21673 );
and ( n23391 , n23385 , n23390 );
and ( n23392 , n23342 , n23390 );
or ( n23393 , n23386 , n23391 , n23392 );
and ( n23394 , n23276 , n23280 );
and ( n23395 , n23280 , n23283 );
and ( n23396 , n23276 , n23283 );
or ( n23397 , n23394 , n23395 , n23396 );
and ( n23398 , n23393 , n23397 );
xor ( n23399 , n23045 , n23049 );
xor ( n23400 , n23399 , n23054 );
and ( n23401 , n23397 , n23400 );
and ( n23402 , n23393 , n23400 );
or ( n23403 , n23398 , n23401 , n23402 );
and ( n23404 , n23291 , n23295 );
and ( n23405 , n23295 , n23298 );
and ( n23406 , n23291 , n23298 );
or ( n23407 , n23404 , n23405 , n23406 );
and ( n23408 , n23403 , n23407 );
xor ( n23409 , n23057 , n23059 );
xor ( n23410 , n23409 , n23062 );
and ( n23411 , n23407 , n23410 );
and ( n23412 , n23403 , n23410 );
or ( n23413 , n23408 , n23411 , n23412 );
and ( n23414 , n23311 , n23413 );
xor ( n23415 , n23065 , n23150 );
xor ( n23416 , n23415 , n23153 );
and ( n23417 , n23413 , n23416 );
and ( n23418 , n23311 , n23416 );
or ( n23419 , n23414 , n23417 , n23418 );
xor ( n23420 , n22976 , n22978 );
xor ( n23421 , n23420 , n22981 );
and ( n23422 , n23419 , n23421 );
xor ( n23423 , n23029 , n23156 );
xor ( n23424 , n23423 , n23159 );
and ( n23425 , n23421 , n23424 );
and ( n23426 , n23419 , n23424 );
or ( n23427 , n23422 , n23425 , n23426 );
and ( n23428 , n23175 , n23427 );
xor ( n23429 , n23419 , n23421 );
xor ( n23430 , n23429 , n23424 );
xor ( n23431 , n23013 , n23015 );
xor ( n23432 , n23431 , n23018 );
xor ( n23433 , n23229 , n23305 );
xor ( n23434 , n23433 , n23308 );
and ( n23435 , n23432 , n23434 );
xor ( n23436 , n23403 , n23407 );
xor ( n23437 , n23436 , n23410 );
and ( n23438 , n23434 , n23437 );
and ( n23439 , n23432 , n23437 );
or ( n23440 , n23435 , n23438 , n23439 );
xor ( n23441 , n23021 , n23023 );
xor ( n23442 , n23441 , n23026 );
and ( n23443 , n23440 , n23442 );
xor ( n23444 , n23311 , n23413 );
xor ( n23445 , n23444 , n23416 );
and ( n23446 , n23442 , n23445 );
and ( n23447 , n23440 , n23445 );
or ( n23448 , n23443 , n23446 , n23447 );
and ( n23449 , n23430 , n23448 );
xor ( n23450 , n23440 , n23442 );
xor ( n23451 , n23450 , n23445 );
xor ( n23452 , n23211 , n23223 );
xor ( n23453 , n23452 , n23226 );
xor ( n23454 , n23287 , n23299 );
xor ( n23455 , n23454 , n23302 );
and ( n23456 , n23453 , n23455 );
and ( n23457 , n21486 , n21739 );
and ( n23458 , n21501 , n21737 );
nor ( n23459 , n23457 , n23458 );
xnor ( n23460 , n23459 , n21749 );
and ( n23461 , n21599 , n21529 );
and ( n23462 , n21545 , n21527 );
nor ( n23463 , n23461 , n23462 );
xnor ( n23464 , n23463 , n21539 );
and ( n23465 , n23460 , n23464 );
and ( n23466 , n22813 , n21496 );
and ( n23467 , n21616 , n21494 );
nor ( n23468 , n23466 , n23467 );
xnor ( n23469 , n23468 , n21506 );
and ( n23470 , n23464 , n23469 );
and ( n23471 , n23460 , n23469 );
or ( n23472 , n23465 , n23470 , n23471 );
and ( n23473 , n21731 , n21260 );
and ( n23474 , n21744 , n21258 );
nor ( n23475 , n23473 , n23474 );
xnor ( n23476 , n23475 , n21270 );
and ( n23477 , n23472 , n23476 );
xor ( n23478 , n23343 , n23353 );
xor ( n23479 , n23478 , n23358 );
and ( n23480 , n23476 , n23479 );
and ( n23481 , n23472 , n23479 );
or ( n23482 , n23477 , n23480 , n23481 );
and ( n23483 , n21712 , n21139 );
and ( n23484 , n21679 , n21137 );
nor ( n23485 , n23483 , n23484 );
xnor ( n23486 , n23485 , n21221 );
and ( n23487 , n23482 , n23486 );
and ( n23488 , n21574 , n21707 );
and ( n23489 , n21252 , n21705 );
nor ( n23490 , n23488 , n23489 );
xnor ( n23491 , n23490 , n21717 );
and ( n23492 , n23486 , n23491 );
and ( n23493 , n23482 , n23491 );
or ( n23494 , n23487 , n23492 , n23493 );
xor ( n23495 , n23347 , n23352 );
and ( n23496 , n23074 , n21496 );
and ( n23497 , n22813 , n21494 );
nor ( n23498 , n23496 , n23497 );
xnor ( n23499 , n23498 , n21506 );
xor ( n23500 , n20615 , n21088 );
buf ( n23501 , n23500 );
buf ( n23502 , n23501 );
buf ( n23503 , n23502 );
and ( n23504 , n23503 , n21513 );
and ( n23505 , n23499 , n23504 );
and ( n23506 , n23495 , n23505 );
and ( n23507 , n21606 , n21625 );
and ( n23508 , n21511 , n21623 );
nor ( n23509 , n23507 , n23508 );
xnor ( n23510 , n23509 , n21635 );
and ( n23511 , n23505 , n23510 );
and ( n23512 , n23495 , n23510 );
or ( n23513 , n23506 , n23511 , n23512 );
and ( n23514 , n21519 , n21582 );
and ( n23515 , n21534 , n21580 );
nor ( n23516 , n23514 , n23515 );
xnor ( n23517 , n23516 , n21588 );
and ( n23518 , n23513 , n23517 );
and ( n23519 , n21645 , n21783 );
and ( n23520 , n21756 , n21781 );
nor ( n23521 , n23519 , n23520 );
xnor ( n23522 , n23521 , n21793 );
and ( n23523 , n23517 , n23522 );
and ( n23524 , n23513 , n23522 );
or ( n23525 , n23518 , n23523 , n23524 );
and ( n23526 , n21241 , n21663 );
and ( n23527 , n21566 , n21661 );
nor ( n23528 , n23526 , n23527 );
xnor ( n23529 , n23528 , n21673 );
and ( n23530 , n23525 , n23529 );
and ( n23531 , n21265 , n21687 );
and ( n23532 , n21226 , n21685 );
nor ( n23533 , n23531 , n23532 );
xnor ( n23534 , n23533 , n21697 );
and ( n23535 , n23529 , n23534 );
and ( n23536 , n23525 , n23534 );
or ( n23537 , n23530 , n23535 , n23536 );
and ( n23538 , n23494 , n23537 );
xor ( n23539 , n23179 , n23183 );
xor ( n23540 , n23539 , n23188 );
and ( n23541 , n23537 , n23540 );
and ( n23542 , n23494 , n23540 );
or ( n23543 , n23538 , n23541 , n23542 );
and ( n23544 , n21501 , n21739 );
and ( n23545 , n21630 , n21737 );
nor ( n23546 , n23544 , n23545 );
xnor ( n23547 , n23546 , n21749 );
and ( n23548 , n21545 , n21529 );
and ( n23549 , n21486 , n21527 );
nor ( n23550 , n23548 , n23549 );
xnor ( n23551 , n23550 , n21539 );
and ( n23552 , n23547 , n23551 );
and ( n23553 , n21616 , n21496 );
and ( n23554 , n21606 , n21494 );
nor ( n23555 , n23553 , n23554 );
xnor ( n23556 , n23555 , n21506 );
and ( n23557 , n23551 , n23556 );
and ( n23558 , n23547 , n23556 );
or ( n23559 , n23552 , n23557 , n23558 );
and ( n23560 , n21777 , n21236 );
and ( n23561 , n21788 , n21234 );
nor ( n23562 , n23560 , n23561 );
xnor ( n23563 , n23562 , n21246 );
and ( n23564 , n23559 , n23563 );
xor ( n23565 , n23312 , n23322 );
xor ( n23566 , n23565 , n23327 );
and ( n23567 , n23563 , n23566 );
and ( n23568 , n23559 , n23566 );
or ( n23569 , n23564 , n23567 , n23568 );
and ( n23570 , n21692 , n21414 );
and ( n23571 , n21655 , n21412 );
nor ( n23572 , n23570 , n23571 );
xnor ( n23573 , n23572 , n21480 );
and ( n23574 , n21744 , n21260 );
and ( n23575 , n22089 , n21258 );
nor ( n23576 , n23574 , n23575 );
xnor ( n23577 , n23576 , n21270 );
and ( n23578 , n23573 , n23577 );
xor ( n23579 , n23361 , n23365 );
xor ( n23580 , n23579 , n23370 );
and ( n23581 , n23577 , n23580 );
and ( n23582 , n23573 , n23580 );
or ( n23583 , n23578 , n23581 , n23582 );
and ( n23584 , n23569 , n23583 );
xor ( n23585 , n23330 , n23334 );
xor ( n23586 , n23585 , n23339 );
and ( n23587 , n23583 , n23586 );
and ( n23588 , n23569 , n23586 );
or ( n23589 , n23584 , n23587 , n23588 );
and ( n23590 , n23543 , n23589 );
xor ( n23591 , n23191 , n23203 );
xor ( n23592 , n23591 , n23208 );
and ( n23593 , n23589 , n23592 );
and ( n23594 , n23543 , n23592 );
or ( n23595 , n23590 , n23593 , n23594 );
and ( n23596 , n22077 , n22032 );
and ( n23597 , n21406 , n22029 );
nor ( n23598 , n23596 , n23597 );
xnor ( n23599 , n23598 , n22027 );
xor ( n23600 , n23373 , n23377 );
xor ( n23601 , n23600 , n23382 );
and ( n23602 , n23599 , n23601 );
xor ( n23603 , n23195 , n23197 );
xor ( n23604 , n23603 , n23200 );
and ( n23605 , n23601 , n23604 );
and ( n23606 , n23599 , n23604 );
or ( n23607 , n23602 , n23605 , n23606 );
xor ( n23608 , n23342 , n23385 );
xor ( n23609 , n23608 , n23390 );
and ( n23610 , n23607 , n23609 );
xor ( n23611 , n23215 , n23217 );
xor ( n23612 , n23611 , n23220 );
and ( n23613 , n23609 , n23612 );
and ( n23614 , n23607 , n23612 );
or ( n23615 , n23610 , n23613 , n23614 );
and ( n23616 , n23595 , n23615 );
xor ( n23617 , n23393 , n23397 );
xor ( n23618 , n23617 , n23400 );
and ( n23619 , n23615 , n23618 );
and ( n23620 , n23595 , n23618 );
or ( n23621 , n23616 , n23619 , n23620 );
and ( n23622 , n23456 , n23621 );
xor ( n23623 , n23432 , n23434 );
xor ( n23624 , n23623 , n23437 );
and ( n23625 , n23621 , n23624 );
and ( n23626 , n23456 , n23624 );
or ( n23627 , n23622 , n23625 , n23626 );
and ( n23628 , n23451 , n23627 );
xor ( n23629 , n23453 , n23455 );
xor ( n23630 , n23595 , n23615 );
xor ( n23631 , n23630 , n23618 );
and ( n23632 , n23629 , n23631 );
xor ( n23633 , n23543 , n23589 );
xor ( n23634 , n23633 , n23592 );
xor ( n23635 , n23607 , n23609 );
xor ( n23636 , n23635 , n23612 );
and ( n23637 , n23634 , n23636 );
and ( n23638 , n23631 , n23637 );
and ( n23639 , n23629 , n23637 );
or ( n23640 , n23632 , n23638 , n23639 );
xor ( n23641 , n23257 , n23271 );
xor ( n23642 , n23641 , n23284 );
xor ( n23643 , n23499 , n23504 );
and ( n23644 , n23320 , n21496 );
and ( n23645 , n23074 , n21494 );
nor ( n23646 , n23644 , n23645 );
xnor ( n23647 , n23646 , n21506 );
xor ( n23648 , n20734 , n21086 );
buf ( n23649 , n23648 );
buf ( n23650 , n23649 );
buf ( n23651 , n23650 );
and ( n23652 , n23651 , n21513 );
and ( n23653 , n23647 , n23652 );
and ( n23654 , n23643 , n23653 );
and ( n23655 , n23351 , n21551 );
and ( n23656 , n23320 , n21549 );
nor ( n23657 , n23655 , n23656 );
xnor ( n23658 , n23657 , n21557 );
and ( n23659 , n23653 , n23658 );
and ( n23660 , n23643 , n23658 );
or ( n23661 , n23654 , n23659 , n23660 );
and ( n23662 , n21756 , n21582 );
and ( n23663 , n21519 , n21580 );
nor ( n23664 , n23662 , n23663 );
xnor ( n23665 , n23664 , n21588 );
and ( n23666 , n23661 , n23665 );
and ( n23667 , n21630 , n21783 );
and ( n23668 , n21645 , n21781 );
nor ( n23669 , n23667 , n23668 );
xnor ( n23670 , n23669 , n21793 );
and ( n23671 , n23665 , n23670 );
and ( n23672 , n23661 , n23670 );
or ( n23673 , n23666 , n23671 , n23672 );
and ( n23674 , n21566 , n21139 );
and ( n23675 , n21712 , n21137 );
nor ( n23676 , n23674 , n23675 );
xnor ( n23677 , n23676 , n21221 );
and ( n23678 , n23673 , n23677 );
and ( n23679 , n21226 , n21663 );
and ( n23680 , n21241 , n21661 );
nor ( n23681 , n23679 , n23680 );
xnor ( n23682 , n23681 , n21673 );
and ( n23683 , n23677 , n23682 );
and ( n23684 , n23673 , n23682 );
or ( n23685 , n23678 , n23683 , n23684 );
and ( n23686 , n21216 , n22032 );
and ( n23687 , n22077 , n22029 );
nor ( n23688 , n23686 , n23687 );
xnor ( n23689 , n23688 , n22027 );
and ( n23690 , n23685 , n23689 );
xor ( n23691 , n23559 , n23563 );
xor ( n23692 , n23691 , n23566 );
and ( n23693 , n23689 , n23692 );
and ( n23694 , n23685 , n23692 );
or ( n23695 , n23690 , n23693 , n23694 );
and ( n23696 , n21129 , n22032 );
and ( n23697 , n21216 , n22029 );
nor ( n23698 , n23696 , n23697 );
xnor ( n23699 , n23698 , n22027 );
and ( n23700 , n21252 , n21687 );
and ( n23701 , n21265 , n21685 );
nor ( n23702 , n23700 , n23701 );
xnor ( n23703 , n23702 , n21697 );
and ( n23704 , n23699 , n23703 );
xor ( n23705 , n23513 , n23517 );
xor ( n23706 , n23705 , n23522 );
and ( n23707 , n23703 , n23706 );
and ( n23708 , n23699 , n23706 );
or ( n23709 , n23704 , n23707 , n23708 );
xor ( n23710 , n23525 , n23529 );
xor ( n23711 , n23710 , n23534 );
and ( n23712 , n23709 , n23711 );
xor ( n23713 , n23573 , n23577 );
xor ( n23714 , n23713 , n23580 );
and ( n23715 , n23711 , n23714 );
and ( n23716 , n23709 , n23714 );
or ( n23717 , n23712 , n23715 , n23716 );
and ( n23718 , n23695 , n23717 );
xor ( n23719 , n23599 , n23601 );
xor ( n23720 , n23719 , n23604 );
and ( n23721 , n23717 , n23720 );
and ( n23722 , n23695 , n23720 );
or ( n23723 , n23718 , n23721 , n23722 );
and ( n23724 , n23642 , n23723 );
xor ( n23725 , n23245 , n23249 );
xor ( n23726 , n23725 , n23254 );
and ( n23727 , n21668 , n22114 );
and ( n23728 , n21129 , n22112 );
nor ( n23729 , n23727 , n23728 );
xnor ( n23730 , n23729 , n22124 );
xor ( n23731 , n23233 , n23237 );
xor ( n23732 , n23731 , n23242 );
and ( n23733 , n23730 , n23732 );
and ( n23734 , n21788 , n21707 );
and ( n23735 , n21574 , n21705 );
nor ( n23736 , n23734 , n23735 );
xnor ( n23737 , n23736 , n21717 );
and ( n23738 , n22089 , n21236 );
and ( n23739 , n21777 , n21234 );
nor ( n23740 , n23738 , n23739 );
xnor ( n23741 , n23740 , n21246 );
and ( n23742 , n23737 , n23741 );
xor ( n23743 , n23547 , n23551 );
xor ( n23744 , n23743 , n23556 );
and ( n23745 , n23741 , n23744 );
and ( n23746 , n23737 , n23744 );
or ( n23747 , n23742 , n23745 , n23746 );
and ( n23748 , n23732 , n23747 );
and ( n23749 , n23730 , n23747 );
or ( n23750 , n23733 , n23748 , n23749 );
and ( n23751 , n23726 , n23750 );
xor ( n23752 , n23494 , n23537 );
xor ( n23753 , n23752 , n23540 );
and ( n23754 , n23750 , n23753 );
and ( n23755 , n23726 , n23753 );
or ( n23756 , n23751 , n23754 , n23755 );
and ( n23757 , n23723 , n23756 );
and ( n23758 , n23642 , n23756 );
or ( n23759 , n23724 , n23757 , n23758 );
xor ( n23760 , n23634 , n23636 );
xor ( n23761 , n23569 , n23583 );
xor ( n23762 , n23761 , n23586 );
xor ( n23763 , n23730 , n23732 );
xor ( n23764 , n23763 , n23747 );
xor ( n23765 , n23482 , n23486 );
xor ( n23766 , n23765 , n23491 );
and ( n23767 , n23764 , n23766 );
and ( n23768 , n21655 , n22114 );
and ( n23769 , n21668 , n22112 );
nor ( n23770 , n23768 , n23769 );
xnor ( n23771 , n23770 , n22124 );
and ( n23772 , n21679 , n21414 );
and ( n23773 , n21692 , n21412 );
nor ( n23774 , n23772 , n23773 );
xnor ( n23775 , n23774 , n21480 );
and ( n23776 , n23771 , n23775 );
and ( n23777 , n21545 , n21739 );
and ( n23778 , n21486 , n21737 );
nor ( n23779 , n23777 , n23778 );
xnor ( n23780 , n23779 , n21749 );
and ( n23781 , n21511 , n21529 );
and ( n23782 , n21599 , n21527 );
nor ( n23783 , n23781 , n23782 );
xnor ( n23784 , n23783 , n21539 );
and ( n23785 , n23780 , n23784 );
and ( n23786 , n21616 , n21625 );
and ( n23787 , n21606 , n21623 );
nor ( n23788 , n23786 , n23787 );
xnor ( n23789 , n23788 , n21635 );
and ( n23790 , n23784 , n23789 );
and ( n23791 , n23780 , n23789 );
or ( n23792 , n23785 , n23790 , n23791 );
and ( n23793 , n21534 , n21260 );
and ( n23794 , n21731 , n21258 );
nor ( n23795 , n23793 , n23794 );
xnor ( n23796 , n23795 , n21270 );
and ( n23797 , n23792 , n23796 );
xor ( n23798 , n23495 , n23505 );
xor ( n23799 , n23798 , n23510 );
and ( n23800 , n23796 , n23799 );
and ( n23801 , n23792 , n23799 );
or ( n23802 , n23797 , n23800 , n23801 );
and ( n23803 , n23775 , n23802 );
and ( n23804 , n23771 , n23802 );
or ( n23805 , n23776 , n23803 , n23804 );
and ( n23806 , n23766 , n23805 );
and ( n23807 , n23764 , n23805 );
or ( n23808 , n23767 , n23806 , n23807 );
and ( n23809 , n23762 , n23808 );
xor ( n23810 , n23695 , n23717 );
xor ( n23811 , n23810 , n23720 );
and ( n23812 , n23808 , n23811 );
and ( n23813 , n23762 , n23811 );
or ( n23814 , n23809 , n23812 , n23813 );
and ( n23815 , n23760 , n23814 );
xor ( n23816 , n23642 , n23723 );
xor ( n23817 , n23816 , n23756 );
and ( n23818 , n23814 , n23817 );
and ( n23819 , n23760 , n23817 );
or ( n23820 , n23815 , n23818 , n23819 );
and ( n23821 , n23759 , n23820 );
xor ( n23822 , n23629 , n23631 );
xor ( n23823 , n23822 , n23637 );
and ( n23824 , n23820 , n23823 );
and ( n23825 , n23759 , n23823 );
or ( n23826 , n23821 , n23824 , n23825 );
and ( n23827 , n23640 , n23826 );
xor ( n23828 , n23456 , n23621 );
xor ( n23829 , n23828 , n23624 );
and ( n23830 , n23826 , n23829 );
and ( n23831 , n23640 , n23829 );
or ( n23832 , n23827 , n23830 , n23831 );
and ( n23833 , n23627 , n23832 );
and ( n23834 , n23451 , n23832 );
or ( n23835 , n23628 , n23833 , n23834 );
and ( n23836 , n23448 , n23835 );
and ( n23837 , n23430 , n23835 );
or ( n23838 , n23449 , n23836 , n23837 );
and ( n23839 , n23427 , n23838 );
and ( n23840 , n23175 , n23838 );
or ( n23841 , n23428 , n23839 , n23840 );
and ( n23842 , n23172 , n23841 );
and ( n23843 , n23170 , n23841 );
or ( n23844 , n23173 , n23842 , n23843 );
and ( n23845 , n23000 , n23844 );
and ( n23846 , n22944 , n23844 );
or ( n23847 , n23001 , n23845 , n23846 );
xor ( n23848 , n22942 , n23847 );
xor ( n23849 , n22944 , n23000 );
xor ( n23850 , n23849 , n23844 );
xor ( n23851 , n23170 , n23172 );
xor ( n23852 , n23851 , n23841 );
xor ( n23853 , n23175 , n23427 );
xor ( n23854 , n23853 , n23838 );
xor ( n23855 , n23430 , n23448 );
xor ( n23856 , n23855 , n23835 );
xor ( n23857 , n23451 , n23627 );
xor ( n23858 , n23857 , n23832 );
xor ( n23859 , n23640 , n23826 );
xor ( n23860 , n23859 , n23829 );
xor ( n23861 , n23759 , n23820 );
xor ( n23862 , n23861 , n23823 );
xor ( n23863 , n23709 , n23711 );
xor ( n23864 , n23863 , n23714 );
xor ( n23865 , n23673 , n23677 );
xor ( n23866 , n23865 , n23682 );
xor ( n23867 , n23699 , n23703 );
xor ( n23868 , n23867 , n23706 );
and ( n23869 , n23866 , n23868 );
and ( n23870 , n23864 , n23869 );
xor ( n23871 , n23764 , n23766 );
xor ( n23872 , n23871 , n23805 );
and ( n23873 , n23869 , n23872 );
and ( n23874 , n23864 , n23872 );
or ( n23875 , n23870 , n23873 , n23874 );
xor ( n23876 , n23726 , n23750 );
xor ( n23877 , n23876 , n23753 );
and ( n23878 , n23875 , n23877 );
xor ( n23879 , n23647 , n23652 );
and ( n23880 , n23651 , n21551 );
and ( n23881 , n23503 , n21549 );
nor ( n23882 , n23880 , n23881 );
xnor ( n23883 , n23882 , n21557 );
xor ( n23884 , n20736 , n21085 );
buf ( n23885 , n23884 );
buf ( n23886 , n23885 );
buf ( n23887 , n23886 );
and ( n23888 , n23887 , n21513 );
and ( n23889 , n23883 , n23888 );
and ( n23890 , n23879 , n23889 );
and ( n23891 , n23503 , n21551 );
and ( n23892 , n23351 , n21549 );
nor ( n23893 , n23891 , n23892 );
xnor ( n23894 , n23893 , n21557 );
and ( n23895 , n23889 , n23894 );
and ( n23896 , n23879 , n23894 );
or ( n23897 , n23890 , n23895 , n23896 );
and ( n23898 , n21519 , n21260 );
and ( n23899 , n21534 , n21258 );
nor ( n23900 , n23898 , n23899 );
xnor ( n23901 , n23900 , n21270 );
and ( n23902 , n23897 , n23901 );
and ( n23903 , n21501 , n21783 );
and ( n23904 , n21630 , n21781 );
nor ( n23905 , n23903 , n23904 );
xnor ( n23906 , n23905 , n21793 );
and ( n23907 , n23901 , n23906 );
and ( n23908 , n23897 , n23906 );
or ( n23909 , n23902 , n23907 , n23908 );
and ( n23910 , n21777 , n21707 );
and ( n23911 , n21788 , n21705 );
nor ( n23912 , n23910 , n23911 );
xnor ( n23913 , n23912 , n21717 );
and ( n23914 , n23909 , n23913 );
and ( n23915 , n21744 , n21236 );
and ( n23916 , n22089 , n21234 );
nor ( n23917 , n23915 , n23916 );
xnor ( n23918 , n23917 , n21246 );
and ( n23919 , n23913 , n23918 );
and ( n23920 , n23909 , n23918 );
or ( n23921 , n23914 , n23919 , n23920 );
and ( n23922 , n21692 , n22114 );
and ( n23923 , n21655 , n22112 );
nor ( n23924 , n23922 , n23923 );
xnor ( n23925 , n23924 , n22124 );
and ( n23926 , n21574 , n21687 );
and ( n23927 , n21252 , n21685 );
nor ( n23928 , n23926 , n23927 );
xnor ( n23929 , n23928 , n21697 );
and ( n23930 , n23925 , n23929 );
xor ( n23931 , n23661 , n23665 );
xor ( n23932 , n23931 , n23670 );
and ( n23933 , n23929 , n23932 );
and ( n23934 , n23925 , n23932 );
or ( n23935 , n23930 , n23933 , n23934 );
and ( n23936 , n23921 , n23935 );
xor ( n23937 , n23472 , n23476 );
xor ( n23938 , n23937 , n23479 );
and ( n23939 , n23935 , n23938 );
and ( n23940 , n23921 , n23938 );
or ( n23941 , n23936 , n23939 , n23940 );
and ( n23942 , n23887 , n21551 );
and ( n23943 , n23651 , n21549 );
nor ( n23944 , n23942 , n23943 );
xnor ( n23945 , n23944 , n21557 );
xor ( n23946 , n20738 , n21084 );
buf ( n23947 , n23946 );
buf ( n23948 , n23947 );
buf ( n23949 , n23948 );
and ( n23950 , n23949 , n21513 );
and ( n23951 , n23945 , n23950 );
and ( n23952 , n23074 , n21625 );
and ( n23953 , n22813 , n21623 );
nor ( n23954 , n23952 , n23953 );
xnor ( n23955 , n23954 , n21635 );
and ( n23956 , n23951 , n23955 );
and ( n23957 , n23351 , n21496 );
and ( n23958 , n23320 , n21494 );
nor ( n23959 , n23957 , n23958 );
xnor ( n23960 , n23959 , n21506 );
and ( n23961 , n23955 , n23960 );
and ( n23962 , n23951 , n23960 );
or ( n23963 , n23956 , n23961 , n23962 );
and ( n23964 , n21606 , n21529 );
and ( n23965 , n21511 , n21527 );
nor ( n23966 , n23964 , n23965 );
xnor ( n23967 , n23966 , n21539 );
and ( n23968 , n23963 , n23967 );
and ( n23969 , n22813 , n21625 );
and ( n23970 , n21616 , n21623 );
nor ( n23971 , n23969 , n23970 );
xnor ( n23972 , n23971 , n21635 );
and ( n23973 , n23967 , n23972 );
and ( n23974 , n23963 , n23972 );
or ( n23975 , n23968 , n23973 , n23974 );
and ( n23976 , n21645 , n21582 );
and ( n23977 , n21756 , n21580 );
nor ( n23978 , n23976 , n23977 );
xnor ( n23979 , n23978 , n21588 );
and ( n23980 , n23975 , n23979 );
xor ( n23981 , n23643 , n23653 );
xor ( n23982 , n23981 , n23658 );
and ( n23983 , n23979 , n23982 );
and ( n23984 , n23975 , n23982 );
or ( n23985 , n23980 , n23983 , n23984 );
and ( n23986 , n21668 , n22032 );
and ( n23987 , n21129 , n22029 );
nor ( n23988 , n23986 , n23987 );
xnor ( n23989 , n23988 , n22027 );
and ( n23990 , n23985 , n23989 );
and ( n23991 , n21712 , n21414 );
and ( n23992 , n21679 , n21412 );
nor ( n23993 , n23991 , n23992 );
xnor ( n23994 , n23993 , n21480 );
and ( n23995 , n23989 , n23994 );
and ( n23996 , n23985 , n23994 );
or ( n23997 , n23990 , n23995 , n23996 );
and ( n23998 , n21241 , n21139 );
and ( n23999 , n21566 , n21137 );
nor ( n24000 , n23998 , n23999 );
xnor ( n24001 , n24000 , n21221 );
and ( n24002 , n21265 , n21663 );
and ( n24003 , n21226 , n21661 );
nor ( n24004 , n24002 , n24003 );
xnor ( n24005 , n24004 , n21673 );
and ( n24006 , n24001 , n24005 );
xor ( n24007 , n23460 , n23464 );
xor ( n24008 , n24007 , n23469 );
and ( n24009 , n24005 , n24008 );
and ( n24010 , n24001 , n24008 );
or ( n24011 , n24006 , n24009 , n24010 );
and ( n24012 , n23997 , n24011 );
xor ( n24013 , n23737 , n23741 );
xor ( n24014 , n24013 , n23744 );
and ( n24015 , n24011 , n24014 );
and ( n24016 , n23997 , n24014 );
or ( n24017 , n24012 , n24015 , n24016 );
and ( n24018 , n23941 , n24017 );
xor ( n24019 , n23685 , n23689 );
xor ( n24020 , n24019 , n23692 );
and ( n24021 , n24017 , n24020 );
and ( n24022 , n23941 , n24020 );
or ( n24023 , n24018 , n24021 , n24022 );
and ( n24024 , n23877 , n24023 );
and ( n24025 , n23875 , n24023 );
or ( n24026 , n23878 , n24024 , n24025 );
xor ( n24027 , n23760 , n23814 );
xor ( n24028 , n24027 , n23817 );
and ( n24029 , n24026 , n24028 );
xor ( n24030 , n23762 , n23808 );
xor ( n24031 , n24030 , n23811 );
and ( n24032 , n21756 , n21260 );
and ( n24033 , n21519 , n21258 );
nor ( n24034 , n24032 , n24033 );
xnor ( n24035 , n24034 , n21270 );
and ( n24036 , n21486 , n21783 );
and ( n24037 , n21501 , n21781 );
nor ( n24038 , n24036 , n24037 );
xnor ( n24039 , n24038 , n21793 );
and ( n24040 , n24035 , n24039 );
and ( n24041 , n21599 , n21739 );
and ( n24042 , n21545 , n21737 );
nor ( n24043 , n24041 , n24042 );
xnor ( n24044 , n24043 , n21749 );
and ( n24045 , n24039 , n24044 );
and ( n24046 , n24035 , n24044 );
or ( n24047 , n24040 , n24045 , n24046 );
and ( n24048 , n21226 , n21139 );
and ( n24049 , n21241 , n21137 );
nor ( n24050 , n24048 , n24049 );
xnor ( n24051 , n24050 , n21221 );
and ( n24052 , n24047 , n24051 );
and ( n24053 , n22089 , n21707 );
and ( n24054 , n21777 , n21705 );
nor ( n24055 , n24053 , n24054 );
xnor ( n24056 , n24055 , n21717 );
and ( n24057 , n24051 , n24056 );
and ( n24058 , n24047 , n24056 );
or ( n24059 , n24052 , n24057 , n24058 );
xor ( n24060 , n23909 , n23913 );
xor ( n24061 , n24060 , n23918 );
and ( n24062 , n24059 , n24061 );
xor ( n24063 , n23925 , n23929 );
xor ( n24064 , n24063 , n23932 );
and ( n24065 , n24061 , n24064 );
and ( n24066 , n24059 , n24064 );
or ( n24067 , n24062 , n24065 , n24066 );
and ( n24068 , n21788 , n21687 );
and ( n24069 , n21574 , n21685 );
nor ( n24070 , n24068 , n24069 );
xnor ( n24071 , n24070 , n21697 );
and ( n24072 , n21731 , n21236 );
and ( n24073 , n21744 , n21234 );
nor ( n24074 , n24072 , n24073 );
xnor ( n24075 , n24074 , n21246 );
and ( n24076 , n24071 , n24075 );
xor ( n24077 , n23780 , n23784 );
xor ( n24078 , n24077 , n23789 );
and ( n24079 , n24075 , n24078 );
and ( n24080 , n24071 , n24078 );
or ( n24081 , n24076 , n24079 , n24080 );
xor ( n24082 , n23883 , n23888 );
and ( n24083 , n21511 , n21739 );
and ( n24084 , n21599 , n21737 );
nor ( n24085 , n24083 , n24084 );
xnor ( n24086 , n24085 , n21749 );
and ( n24087 , n24082 , n24086 );
and ( n24088 , n21616 , n21529 );
and ( n24089 , n21606 , n21527 );
nor ( n24090 , n24088 , n24089 );
xnor ( n24091 , n24090 , n21539 );
and ( n24092 , n24086 , n24091 );
and ( n24093 , n24082 , n24091 );
or ( n24094 , n24087 , n24092 , n24093 );
and ( n24095 , n21630 , n21582 );
and ( n24096 , n21645 , n21580 );
nor ( n24097 , n24095 , n24096 );
xnor ( n24098 , n24097 , n21588 );
and ( n24099 , n24094 , n24098 );
xor ( n24100 , n23879 , n23889 );
xor ( n24101 , n24100 , n23894 );
and ( n24102 , n24098 , n24101 );
and ( n24103 , n24094 , n24101 );
or ( n24104 , n24099 , n24102 , n24103 );
and ( n24105 , n21252 , n21663 );
and ( n24106 , n21265 , n21661 );
nor ( n24107 , n24105 , n24106 );
xnor ( n24108 , n24107 , n21673 );
and ( n24109 , n24104 , n24108 );
xor ( n24110 , n23897 , n23901 );
xor ( n24111 , n24110 , n23906 );
and ( n24112 , n24108 , n24111 );
and ( n24113 , n24104 , n24111 );
or ( n24114 , n24109 , n24112 , n24113 );
and ( n24115 , n24081 , n24114 );
xor ( n24116 , n23792 , n23796 );
xor ( n24117 , n24116 , n23799 );
and ( n24118 , n24114 , n24117 );
and ( n24119 , n24081 , n24117 );
or ( n24120 , n24115 , n24118 , n24119 );
and ( n24121 , n24067 , n24120 );
xor ( n24122 , n23921 , n23935 );
xor ( n24123 , n24122 , n23938 );
and ( n24124 , n24120 , n24123 );
and ( n24125 , n24067 , n24123 );
or ( n24126 , n24121 , n24124 , n24125 );
xor ( n24127 , n23941 , n24017 );
xor ( n24128 , n24127 , n24020 );
and ( n24129 , n24126 , n24128 );
and ( n24130 , n24031 , n24129 );
xor ( n24131 , n23875 , n23877 );
xor ( n24132 , n24131 , n24023 );
and ( n24133 , n24129 , n24132 );
and ( n24134 , n24031 , n24132 );
or ( n24135 , n24130 , n24133 , n24134 );
and ( n24136 , n24028 , n24135 );
and ( n24137 , n24026 , n24135 );
or ( n24138 , n24029 , n24136 , n24137 );
and ( n24139 , n23862 , n24138 );
xor ( n24140 , n23862 , n24138 );
xor ( n24141 , n24026 , n24028 );
xor ( n24142 , n24141 , n24135 );
xor ( n24143 , n23864 , n23869 );
xor ( n24144 , n24143 , n23872 );
xor ( n24145 , n23771 , n23775 );
xor ( n24146 , n24145 , n23802 );
xor ( n24147 , n23866 , n23868 );
and ( n24148 , n24146 , n24147 );
xor ( n24149 , n23997 , n24011 );
xor ( n24150 , n24149 , n24014 );
and ( n24151 , n24147 , n24150 );
and ( n24152 , n24146 , n24150 );
or ( n24153 , n24148 , n24151 , n24152 );
and ( n24154 , n24144 , n24153 );
xor ( n24155 , n24126 , n24128 );
and ( n24156 , n24153 , n24155 );
and ( n24157 , n24144 , n24155 );
or ( n24158 , n24154 , n24156 , n24157 );
xor ( n24159 , n24031 , n24129 );
xor ( n24160 , n24159 , n24132 );
and ( n24161 , n24158 , n24160 );
and ( n24162 , n21265 , n21139 );
and ( n24163 , n21226 , n21137 );
nor ( n24164 , n24162 , n24163 );
xnor ( n24165 , n24164 , n21221 );
xor ( n24166 , n24035 , n24039 );
xor ( n24167 , n24166 , n24044 );
and ( n24168 , n24165 , n24167 );
xor ( n24169 , n24094 , n24098 );
xor ( n24170 , n24169 , n24101 );
and ( n24171 , n24167 , n24170 );
and ( n24172 , n24165 , n24170 );
or ( n24173 , n24168 , n24171 , n24172 );
xor ( n24174 , n24047 , n24051 );
xor ( n24175 , n24174 , n24056 );
and ( n24176 , n24173 , n24175 );
xor ( n24177 , n24071 , n24075 );
xor ( n24178 , n24177 , n24078 );
and ( n24179 , n24175 , n24178 );
and ( n24180 , n24173 , n24178 );
or ( n24181 , n24176 , n24179 , n24180 );
xor ( n24182 , n23985 , n23989 );
xor ( n24183 , n24182 , n23994 );
and ( n24184 , n24181 , n24183 );
xor ( n24185 , n24081 , n24114 );
xor ( n24186 , n24185 , n24117 );
and ( n24187 , n24183 , n24186 );
and ( n24188 , n24181 , n24186 );
or ( n24189 , n24184 , n24187 , n24188 );
and ( n24190 , n21692 , n22032 );
and ( n24191 , n21655 , n22029 );
nor ( n24192 , n24190 , n24191 );
xnor ( n24193 , n24192 , n22027 );
and ( n24194 , n21241 , n21414 );
and ( n24195 , n21566 , n21412 );
nor ( n24196 , n24194 , n24195 );
xnor ( n24197 , n24196 , n21480 );
and ( n24198 , n24193 , n24197 );
and ( n24199 , n21574 , n21663 );
and ( n24200 , n21252 , n21661 );
nor ( n24201 , n24199 , n24200 );
xnor ( n24202 , n24201 , n21673 );
and ( n24203 , n24197 , n24202 );
and ( n24204 , n24193 , n24202 );
or ( n24205 , n24198 , n24203 , n24204 );
and ( n24206 , n23949 , n21551 );
and ( n24207 , n23887 , n21549 );
nor ( n24208 , n24206 , n24207 );
xnor ( n24209 , n24208 , n21557 );
xor ( n24210 , n20811 , n21082 );
buf ( n24211 , n24210 );
buf ( n24212 , n24211 );
buf ( n24213 , n24212 );
and ( n24214 , n24213 , n21513 );
and ( n24215 , n24209 , n24214 );
and ( n24216 , n23320 , n21625 );
and ( n24217 , n23074 , n21623 );
nor ( n24218 , n24216 , n24217 );
xnor ( n24219 , n24218 , n21635 );
and ( n24220 , n24215 , n24219 );
and ( n24221 , n23503 , n21496 );
and ( n24222 , n23351 , n21494 );
nor ( n24223 , n24221 , n24222 );
xnor ( n24224 , n24223 , n21506 );
and ( n24225 , n24219 , n24224 );
and ( n24226 , n24215 , n24224 );
or ( n24227 , n24220 , n24225 , n24226 );
and ( n24228 , n21501 , n21582 );
and ( n24229 , n21630 , n21580 );
nor ( n24230 , n24228 , n24229 );
xnor ( n24231 , n24230 , n21588 );
and ( n24232 , n24227 , n24231 );
and ( n24233 , n21545 , n21783 );
and ( n24234 , n21486 , n21781 );
nor ( n24235 , n24233 , n24234 );
xnor ( n24236 , n24235 , n21793 );
and ( n24237 , n24231 , n24236 );
and ( n24238 , n24227 , n24236 );
or ( n24239 , n24232 , n24237 , n24238 );
and ( n24240 , n21534 , n21236 );
and ( n24241 , n21731 , n21234 );
nor ( n24242 , n24240 , n24241 );
xnor ( n24243 , n24242 , n21246 );
and ( n24244 , n24239 , n24243 );
xor ( n24245 , n23963 , n23967 );
xor ( n24246 , n24245 , n23972 );
and ( n24247 , n24243 , n24246 );
and ( n24248 , n24239 , n24246 );
or ( n24249 , n24244 , n24247 , n24248 );
and ( n24250 , n21679 , n22114 );
and ( n24251 , n21692 , n22112 );
nor ( n24252 , n24250 , n24251 );
xnor ( n24253 , n24252 , n22124 );
xor ( n24254 , n24249 , n24253 );
and ( n24255 , n21566 , n21414 );
and ( n24256 , n21712 , n21412 );
nor ( n24257 , n24255 , n24256 );
xnor ( n24258 , n24257 , n21480 );
xor ( n24259 , n24254 , n24258 );
and ( n24260 , n24205 , n24259 );
xor ( n24261 , n24104 , n24108 );
xor ( n24262 , n24261 , n24111 );
and ( n24263 , n24259 , n24262 );
and ( n24264 , n24205 , n24262 );
or ( n24265 , n24260 , n24263 , n24264 );
xor ( n24266 , n24059 , n24061 );
xor ( n24267 , n24266 , n24064 );
and ( n24268 , n24265 , n24267 );
and ( n24269 , n24249 , n24253 );
and ( n24270 , n24253 , n24258 );
and ( n24271 , n24249 , n24258 );
or ( n24272 , n24269 , n24270 , n24271 );
xor ( n24273 , n23945 , n23950 );
and ( n24274 , n21606 , n21739 );
and ( n24275 , n21511 , n21737 );
nor ( n24276 , n24274 , n24275 );
xnor ( n24277 , n24276 , n21749 );
and ( n24278 , n24273 , n24277 );
and ( n24279 , n22813 , n21529 );
and ( n24280 , n21616 , n21527 );
nor ( n24281 , n24279 , n24280 );
xnor ( n24282 , n24281 , n21539 );
and ( n24283 , n24277 , n24282 );
and ( n24284 , n24273 , n24282 );
or ( n24285 , n24278 , n24283 , n24284 );
and ( n24286 , n21519 , n21236 );
and ( n24287 , n21534 , n21234 );
nor ( n24288 , n24286 , n24287 );
xnor ( n24289 , n24288 , n21246 );
and ( n24290 , n24285 , n24289 );
xor ( n24291 , n23951 , n23955 );
xor ( n24292 , n24291 , n23960 );
and ( n24293 , n24289 , n24292 );
and ( n24294 , n24285 , n24292 );
or ( n24295 , n24290 , n24293 , n24294 );
and ( n24296 , n21777 , n21687 );
and ( n24297 , n21788 , n21685 );
nor ( n24298 , n24296 , n24297 );
xnor ( n24299 , n24298 , n21697 );
and ( n24300 , n24295 , n24299 );
and ( n24301 , n21744 , n21707 );
and ( n24302 , n22089 , n21705 );
nor ( n24303 , n24301 , n24302 );
xnor ( n24304 , n24303 , n21717 );
and ( n24305 , n24299 , n24304 );
and ( n24306 , n24295 , n24304 );
or ( n24307 , n24300 , n24305 , n24306 );
and ( n24308 , n21655 , n22032 );
and ( n24309 , n21668 , n22029 );
nor ( n24310 , n24308 , n24309 );
xnor ( n24311 , n24310 , n22027 );
and ( n24312 , n24307 , n24311 );
xor ( n24313 , n23975 , n23979 );
xor ( n24314 , n24313 , n23982 );
and ( n24315 , n24311 , n24314 );
and ( n24316 , n24307 , n24314 );
or ( n24317 , n24312 , n24315 , n24316 );
xor ( n24318 , n24272 , n24317 );
xor ( n24319 , n24001 , n24005 );
xor ( n24320 , n24319 , n24008 );
xor ( n24321 , n24318 , n24320 );
and ( n24322 , n24267 , n24321 );
and ( n24323 , n24265 , n24321 );
or ( n24324 , n24268 , n24322 , n24323 );
and ( n24325 , n24189 , n24324 );
xor ( n24326 , n24067 , n24120 );
xor ( n24327 , n24326 , n24123 );
and ( n24328 , n24324 , n24327 );
and ( n24329 , n24189 , n24327 );
or ( n24330 , n24325 , n24328 , n24329 );
and ( n24331 , n24272 , n24317 );
and ( n24332 , n24317 , n24320 );
and ( n24333 , n24272 , n24320 );
or ( n24334 , n24331 , n24332 , n24333 );
xor ( n24335 , n24146 , n24147 );
xor ( n24336 , n24335 , n24150 );
and ( n24337 , n24334 , n24336 );
xor ( n24338 , n24189 , n24324 );
xor ( n24339 , n24338 , n24327 );
and ( n24340 , n24336 , n24339 );
and ( n24341 , n24334 , n24339 );
or ( n24342 , n24337 , n24340 , n24341 );
and ( n24343 , n24330 , n24342 );
xor ( n24344 , n24144 , n24153 );
xor ( n24345 , n24344 , n24155 );
and ( n24346 , n24342 , n24345 );
and ( n24347 , n24330 , n24345 );
or ( n24348 , n24343 , n24346 , n24347 );
and ( n24349 , n24160 , n24348 );
and ( n24350 , n24158 , n24348 );
or ( n24351 , n24161 , n24349 , n24350 );
and ( n24352 , n24142 , n24351 );
xor ( n24353 , n24142 , n24351 );
xor ( n24354 , n24158 , n24160 );
xor ( n24355 , n24354 , n24348 );
xor ( n24356 , n24181 , n24183 );
xor ( n24357 , n24356 , n24186 );
and ( n24358 , n21731 , n21707 );
and ( n24359 , n21744 , n21705 );
nor ( n24360 , n24358 , n24359 );
xnor ( n24361 , n24360 , n21717 );
and ( n24362 , n21645 , n21260 );
and ( n24363 , n21756 , n21258 );
nor ( n24364 , n24362 , n24363 );
xnor ( n24365 , n24364 , n21270 );
and ( n24366 , n24361 , n24365 );
xor ( n24367 , n24082 , n24086 );
xor ( n24368 , n24367 , n24091 );
and ( n24369 , n24365 , n24368 );
and ( n24370 , n24361 , n24368 );
or ( n24371 , n24366 , n24369 , n24370 );
and ( n24372 , n21712 , n22114 );
and ( n24373 , n21679 , n22112 );
nor ( n24374 , n24372 , n24373 );
xnor ( n24375 , n24374 , n22124 );
and ( n24376 , n24371 , n24375 );
xor ( n24377 , n24239 , n24243 );
xor ( n24378 , n24377 , n24246 );
and ( n24379 , n24375 , n24378 );
and ( n24380 , n24371 , n24378 );
or ( n24381 , n24376 , n24379 , n24380 );
xor ( n24382 , n24307 , n24311 );
xor ( n24383 , n24382 , n24314 );
and ( n24384 , n24381 , n24383 );
and ( n24385 , n24357 , n24384 );
xor ( n24386 , n24265 , n24267 );
xor ( n24387 , n24386 , n24321 );
and ( n24388 , n24384 , n24387 );
and ( n24389 , n24357 , n24387 );
or ( n24390 , n24385 , n24388 , n24389 );
and ( n24391 , n21226 , n21414 );
and ( n24392 , n21241 , n21412 );
nor ( n24393 , n24391 , n24392 );
xnor ( n24394 , n24393 , n21480 );
and ( n24395 , n21252 , n21139 );
and ( n24396 , n21265 , n21137 );
nor ( n24397 , n24395 , n24396 );
xnor ( n24398 , n24397 , n21221 );
and ( n24399 , n24394 , n24398 );
xor ( n24400 , n24285 , n24289 );
xor ( n24401 , n24400 , n24292 );
and ( n24402 , n24398 , n24401 );
and ( n24403 , n24394 , n24401 );
or ( n24404 , n24399 , n24402 , n24403 );
xor ( n24405 , n24193 , n24197 );
xor ( n24406 , n24405 , n24202 );
and ( n24407 , n24404 , n24406 );
xor ( n24408 , n24165 , n24167 );
xor ( n24409 , n24408 , n24170 );
and ( n24410 , n24406 , n24409 );
and ( n24411 , n24404 , n24409 );
or ( n24412 , n24407 , n24410 , n24411 );
xor ( n24413 , n24173 , n24175 );
xor ( n24414 , n24413 , n24178 );
and ( n24415 , n24412 , n24414 );
xor ( n24416 , n24205 , n24259 );
xor ( n24417 , n24416 , n24262 );
and ( n24418 , n24414 , n24417 );
and ( n24419 , n24412 , n24417 );
or ( n24420 , n24415 , n24418 , n24419 );
and ( n24421 , n21566 , n22114 );
and ( n24422 , n21712 , n22112 );
nor ( n24423 , n24421 , n24422 );
xnor ( n24424 , n24423 , n22124 );
and ( n24425 , n21788 , n21663 );
and ( n24426 , n21574 , n21661 );
nor ( n24427 , n24425 , n24426 );
xnor ( n24428 , n24427 , n21673 );
and ( n24429 , n24424 , n24428 );
and ( n24430 , n21712 , n22032 );
and ( n24431 , n21679 , n22029 );
nor ( n24432 , n24430 , n24431 );
xnor ( n24433 , n24432 , n22027 );
and ( n24434 , n21241 , n22114 );
and ( n24435 , n21566 , n22112 );
nor ( n24436 , n24434 , n24435 );
xnor ( n24437 , n24436 , n22124 );
and ( n24438 , n24433 , n24437 );
and ( n24439 , n21777 , n21663 );
and ( n24440 , n21788 , n21661 );
nor ( n24441 , n24439 , n24440 );
xnor ( n24442 , n24441 , n21673 );
and ( n24443 , n24437 , n24442 );
and ( n24444 , n24433 , n24442 );
or ( n24445 , n24438 , n24443 , n24444 );
and ( n24446 , n24428 , n24445 );
and ( n24447 , n24424 , n24445 );
or ( n24448 , n24429 , n24446 , n24447 );
xor ( n24449 , n24295 , n24299 );
xor ( n24450 , n24449 , n24304 );
and ( n24451 , n24448 , n24450 );
xor ( n24452 , n24209 , n24214 );
and ( n24453 , n24213 , n21551 );
and ( n24454 , n23949 , n21549 );
nor ( n24455 , n24453 , n24454 );
xnor ( n24456 , n24455 , n21557 );
xor ( n24457 , n20813 , n21081 );
buf ( n24458 , n24457 );
buf ( n24459 , n24458 );
buf ( n24460 , n24459 );
and ( n24461 , n24460 , n21513 );
and ( n24462 , n24456 , n24461 );
and ( n24463 , n24452 , n24462 );
and ( n24464 , n23651 , n21496 );
and ( n24465 , n23503 , n21494 );
nor ( n24466 , n24464 , n24465 );
xnor ( n24467 , n24466 , n21506 );
and ( n24468 , n24462 , n24467 );
and ( n24469 , n24452 , n24467 );
or ( n24470 , n24463 , n24468 , n24469 );
and ( n24471 , n21486 , n21582 );
and ( n24472 , n21501 , n21580 );
nor ( n24473 , n24471 , n24472 );
xnor ( n24474 , n24473 , n21588 );
and ( n24475 , n24470 , n24474 );
and ( n24476 , n21599 , n21783 );
and ( n24477 , n21545 , n21781 );
nor ( n24478 , n24476 , n24477 );
xnor ( n24479 , n24478 , n21793 );
and ( n24480 , n24474 , n24479 );
and ( n24481 , n24470 , n24479 );
or ( n24482 , n24475 , n24480 , n24481 );
and ( n24483 , n21616 , n21739 );
and ( n24484 , n21606 , n21737 );
nor ( n24485 , n24483 , n24484 );
xnor ( n24486 , n24485 , n21749 );
and ( n24487 , n23074 , n21529 );
and ( n24488 , n22813 , n21527 );
nor ( n24489 , n24487 , n24488 );
xnor ( n24490 , n24489 , n21539 );
and ( n24491 , n24486 , n24490 );
and ( n24492 , n23351 , n21625 );
and ( n24493 , n23320 , n21623 );
nor ( n24494 , n24492 , n24493 );
xnor ( n24495 , n24494 , n21635 );
and ( n24496 , n24490 , n24495 );
and ( n24497 , n24486 , n24495 );
or ( n24498 , n24491 , n24496 , n24497 );
and ( n24499 , n21756 , n21236 );
and ( n24500 , n21519 , n21234 );
nor ( n24501 , n24499 , n24500 );
xnor ( n24502 , n24501 , n21246 );
and ( n24503 , n24498 , n24502 );
xor ( n24504 , n24215 , n24219 );
xor ( n24505 , n24504 , n24224 );
and ( n24506 , n24502 , n24505 );
and ( n24507 , n24498 , n24505 );
or ( n24508 , n24503 , n24506 , n24507 );
and ( n24509 , n24482 , n24508 );
and ( n24510 , n22089 , n21687 );
and ( n24511 , n21777 , n21685 );
nor ( n24512 , n24510 , n24511 );
xnor ( n24513 , n24512 , n21697 );
and ( n24514 , n24508 , n24513 );
and ( n24515 , n24482 , n24513 );
or ( n24516 , n24509 , n24514 , n24515 );
and ( n24517 , n24450 , n24516 );
and ( n24518 , n24448 , n24516 );
or ( n24519 , n24451 , n24517 , n24518 );
xor ( n24520 , n24381 , n24383 );
and ( n24521 , n24519 , n24520 );
and ( n24522 , n21534 , n21707 );
and ( n24523 , n21731 , n21705 );
nor ( n24524 , n24522 , n24523 );
xnor ( n24525 , n24524 , n21717 );
and ( n24526 , n21630 , n21260 );
and ( n24527 , n21645 , n21258 );
nor ( n24528 , n24526 , n24527 );
xnor ( n24529 , n24528 , n21270 );
and ( n24530 , n24525 , n24529 );
xor ( n24531 , n24273 , n24277 );
xor ( n24532 , n24531 , n24282 );
and ( n24533 , n24529 , n24532 );
and ( n24534 , n24525 , n24532 );
or ( n24535 , n24530 , n24533 , n24534 );
and ( n24536 , n21679 , n22032 );
and ( n24537 , n21692 , n22029 );
nor ( n24538 , n24536 , n24537 );
xnor ( n24539 , n24538 , n22027 );
and ( n24540 , n24535 , n24539 );
xor ( n24541 , n24361 , n24365 );
xor ( n24542 , n24541 , n24368 );
and ( n24543 , n24539 , n24542 );
and ( n24544 , n24535 , n24542 );
or ( n24545 , n24540 , n24543 , n24544 );
xor ( n24546 , n24371 , n24375 );
xor ( n24547 , n24546 , n24378 );
and ( n24548 , n24545 , n24547 );
and ( n24549 , n24520 , n24548 );
and ( n24550 , n24519 , n24548 );
or ( n24551 , n24521 , n24549 , n24550 );
and ( n24552 , n24420 , n24551 );
xor ( n24553 , n24424 , n24428 );
xor ( n24554 , n24553 , n24445 );
xor ( n24555 , n24227 , n24231 );
xor ( n24556 , n24555 , n24236 );
and ( n24557 , n24554 , n24556 );
and ( n24558 , n21519 , n21707 );
and ( n24559 , n21534 , n21705 );
nor ( n24560 , n24558 , n24559 );
xnor ( n24561 , n24560 , n21717 );
and ( n24562 , n21645 , n21236 );
and ( n24563 , n21756 , n21234 );
nor ( n24564 , n24562 , n24563 );
xnor ( n24565 , n24564 , n21246 );
and ( n24566 , n24561 , n24565 );
xor ( n24567 , n24486 , n24490 );
xor ( n24568 , n24567 , n24495 );
and ( n24569 , n24565 , n24568 );
and ( n24570 , n24561 , n24568 );
or ( n24571 , n24566 , n24569 , n24570 );
and ( n24572 , n21265 , n21414 );
and ( n24573 , n21226 , n21412 );
nor ( n24574 , n24572 , n24573 );
xnor ( n24575 , n24574 , n21480 );
and ( n24576 , n24571 , n24575 );
and ( n24577 , n21574 , n21139 );
and ( n24578 , n21252 , n21137 );
nor ( n24579 , n24577 , n24578 );
xnor ( n24580 , n24579 , n21221 );
and ( n24581 , n24575 , n24580 );
and ( n24582 , n24571 , n24580 );
or ( n24583 , n24576 , n24581 , n24582 );
and ( n24584 , n24556 , n24583 );
and ( n24585 , n24554 , n24583 );
or ( n24586 , n24557 , n24584 , n24585 );
xor ( n24587 , n24404 , n24406 );
xor ( n24588 , n24587 , n24409 );
and ( n24589 , n24586 , n24588 );
xor ( n24590 , n24482 , n24508 );
xor ( n24591 , n24590 , n24513 );
xor ( n24592 , n24394 , n24398 );
xor ( n24593 , n24592 , n24401 );
and ( n24594 , n24591 , n24593 );
xor ( n24595 , n24535 , n24539 );
xor ( n24596 , n24595 , n24542 );
and ( n24597 , n24593 , n24596 );
and ( n24598 , n24591 , n24596 );
or ( n24599 , n24594 , n24597 , n24598 );
and ( n24600 , n24588 , n24599 );
and ( n24601 , n24586 , n24599 );
or ( n24602 , n24589 , n24600 , n24601 );
xor ( n24603 , n24412 , n24414 );
xor ( n24604 , n24603 , n24417 );
and ( n24605 , n24602 , n24604 );
xor ( n24606 , n24448 , n24450 );
xor ( n24607 , n24606 , n24516 );
xor ( n24608 , n24545 , n24547 );
and ( n24609 , n24607 , n24608 );
xor ( n24610 , n24433 , n24437 );
xor ( n24611 , n24610 , n24442 );
xor ( n24612 , n24470 , n24474 );
xor ( n24613 , n24612 , n24479 );
and ( n24614 , n24611 , n24613 );
xor ( n24615 , n24571 , n24575 );
xor ( n24616 , n24615 , n24580 );
and ( n24617 , n24613 , n24616 );
and ( n24618 , n24611 , n24616 );
or ( n24619 , n24614 , n24617 , n24618 );
xor ( n24620 , n24554 , n24556 );
xor ( n24621 , n24620 , n24583 );
and ( n24622 , n24619 , n24621 );
xor ( n24623 , n24456 , n24461 );
and ( n24624 , n24460 , n21551 );
and ( n24625 , n24213 , n21549 );
nor ( n24626 , n24624 , n24625 );
xnor ( n24627 , n24626 , n21557 );
xor ( n24628 , n20855 , n21079 );
buf ( n24629 , n24628 );
buf ( n24630 , n24629 );
buf ( n24631 , n24630 );
and ( n24632 , n24631 , n21513 );
and ( n24633 , n24627 , n24632 );
and ( n24634 , n24623 , n24633 );
and ( n24635 , n23887 , n21496 );
and ( n24636 , n23651 , n21494 );
nor ( n24637 , n24635 , n24636 );
xnor ( n24638 , n24637 , n21506 );
and ( n24639 , n24633 , n24638 );
and ( n24640 , n24623 , n24638 );
or ( n24641 , n24634 , n24639 , n24640 );
and ( n24642 , n21501 , n21260 );
and ( n24643 , n21630 , n21258 );
nor ( n24644 , n24642 , n24643 );
xnor ( n24645 , n24644 , n21270 );
and ( n24646 , n24641 , n24645 );
and ( n24647 , n21511 , n21783 );
and ( n24648 , n21599 , n21781 );
nor ( n24649 , n24647 , n24648 );
xnor ( n24650 , n24649 , n21793 );
and ( n24651 , n24645 , n24650 );
and ( n24652 , n24641 , n24650 );
or ( n24653 , n24646 , n24651 , n24652 );
xor ( n24654 , n24627 , n24632 );
and ( n24655 , n24631 , n21551 );
and ( n24656 , n24460 , n21549 );
nor ( n24657 , n24655 , n24656 );
xnor ( n24658 , n24657 , n21557 );
xor ( n24659 , n20888 , n21077 );
buf ( n24660 , n24659 );
buf ( n24661 , n24660 );
buf ( n24662 , n24661 );
and ( n24663 , n24662 , n21513 );
and ( n24664 , n24658 , n24663 );
and ( n24665 , n24654 , n24664 );
and ( n24666 , n23949 , n21496 );
and ( n24667 , n23887 , n21494 );
nor ( n24668 , n24666 , n24667 );
xnor ( n24669 , n24668 , n21506 );
and ( n24670 , n24664 , n24669 );
and ( n24671 , n24654 , n24669 );
or ( n24672 , n24665 , n24670 , n24671 );
and ( n24673 , n23320 , n21529 );
and ( n24674 , n23074 , n21527 );
nor ( n24675 , n24673 , n24674 );
xnor ( n24676 , n24675 , n21539 );
and ( n24677 , n24672 , n24676 );
and ( n24678 , n23503 , n21625 );
and ( n24679 , n23351 , n21623 );
nor ( n24680 , n24678 , n24679 );
xnor ( n24681 , n24680 , n21635 );
and ( n24682 , n24676 , n24681 );
and ( n24683 , n24672 , n24681 );
or ( n24684 , n24677 , n24682 , n24683 );
and ( n24685 , n21545 , n21582 );
and ( n24686 , n21486 , n21580 );
nor ( n24687 , n24685 , n24686 );
xnor ( n24688 , n24687 , n21588 );
and ( n24689 , n24684 , n24688 );
xor ( n24690 , n24452 , n24462 );
xor ( n24691 , n24690 , n24467 );
and ( n24692 , n24688 , n24691 );
and ( n24693 , n24684 , n24691 );
or ( n24694 , n24689 , n24692 , n24693 );
and ( n24695 , n24653 , n24694 );
and ( n24696 , n21744 , n21687 );
and ( n24697 , n22089 , n21685 );
nor ( n24698 , n24696 , n24697 );
xnor ( n24699 , n24698 , n21697 );
and ( n24700 , n24694 , n24699 );
and ( n24701 , n24653 , n24699 );
or ( n24702 , n24695 , n24700 , n24701 );
and ( n24703 , n24621 , n24702 );
and ( n24704 , n24619 , n24702 );
or ( n24705 , n24622 , n24703 , n24704 );
and ( n24706 , n24608 , n24705 );
and ( n24707 , n24607 , n24705 );
or ( n24708 , n24609 , n24706 , n24707 );
and ( n24709 , n24604 , n24708 );
and ( n24710 , n24602 , n24708 );
or ( n24711 , n24605 , n24709 , n24710 );
and ( n24712 , n24551 , n24711 );
and ( n24713 , n24420 , n24711 );
or ( n24714 , n24552 , n24712 , n24713 );
and ( n24715 , n24390 , n24714 );
xor ( n24716 , n24334 , n24336 );
xor ( n24717 , n24716 , n24339 );
and ( n24718 , n24714 , n24717 );
and ( n24719 , n24390 , n24717 );
or ( n24720 , n24715 , n24718 , n24719 );
xor ( n24721 , n24330 , n24342 );
xor ( n24722 , n24721 , n24345 );
and ( n24723 , n24720 , n24722 );
xor ( n24724 , n24720 , n24722 );
xor ( n24725 , n24357 , n24384 );
xor ( n24726 , n24725 , n24387 );
xor ( n24727 , n24519 , n24520 );
xor ( n24728 , n24727 , n24548 );
xor ( n24729 , n24586 , n24588 );
xor ( n24730 , n24729 , n24599 );
xor ( n24731 , n24498 , n24502 );
xor ( n24732 , n24731 , n24505 );
and ( n24733 , n21566 , n22032 );
and ( n24734 , n21712 , n22029 );
nor ( n24735 , n24733 , n24734 );
xnor ( n24736 , n24735 , n22027 );
and ( n24737 , n21252 , n21414 );
and ( n24738 , n21265 , n21412 );
nor ( n24739 , n24737 , n24738 );
xnor ( n24740 , n24739 , n21480 );
and ( n24741 , n24736 , n24740 );
xor ( n24742 , n24561 , n24565 );
xor ( n24743 , n24742 , n24568 );
and ( n24744 , n24740 , n24743 );
and ( n24745 , n24736 , n24743 );
or ( n24746 , n24741 , n24744 , n24745 );
and ( n24747 , n24732 , n24746 );
and ( n24748 , n23074 , n21739 );
and ( n24749 , n22813 , n21737 );
nor ( n24750 , n24748 , n24749 );
xnor ( n24751 , n24750 , n21749 );
and ( n24752 , n23351 , n21529 );
and ( n24753 , n23320 , n21527 );
nor ( n24754 , n24752 , n24753 );
xnor ( n24755 , n24754 , n21539 );
and ( n24756 , n24751 , n24755 );
and ( n24757 , n23651 , n21625 );
and ( n24758 , n23503 , n21623 );
nor ( n24759 , n24757 , n24758 );
xnor ( n24760 , n24759 , n21635 );
and ( n24761 , n24755 , n24760 );
and ( n24762 , n24751 , n24760 );
or ( n24763 , n24756 , n24761 , n24762 );
and ( n24764 , n21606 , n21783 );
and ( n24765 , n21511 , n21781 );
nor ( n24766 , n24764 , n24765 );
xnor ( n24767 , n24766 , n21793 );
and ( n24768 , n24763 , n24767 );
and ( n24769 , n22813 , n21739 );
and ( n24770 , n21616 , n21737 );
nor ( n24771 , n24769 , n24770 );
xnor ( n24772 , n24771 , n21749 );
and ( n24773 , n24767 , n24772 );
and ( n24774 , n24763 , n24772 );
or ( n24775 , n24768 , n24773 , n24774 );
and ( n24776 , n21486 , n21260 );
and ( n24777 , n21501 , n21258 );
nor ( n24778 , n24776 , n24777 );
xnor ( n24779 , n24778 , n21270 );
and ( n24780 , n21599 , n21582 );
and ( n24781 , n21545 , n21580 );
nor ( n24782 , n24780 , n24781 );
xnor ( n24783 , n24782 , n21588 );
and ( n24784 , n24779 , n24783 );
xor ( n24785 , n24623 , n24633 );
xor ( n24786 , n24785 , n24638 );
and ( n24787 , n24783 , n24786 );
and ( n24788 , n24779 , n24786 );
or ( n24789 , n24784 , n24787 , n24788 );
and ( n24790 , n24775 , n24789 );
and ( n24791 , n21731 , n21687 );
and ( n24792 , n21744 , n21685 );
nor ( n24793 , n24791 , n24792 );
xnor ( n24794 , n24793 , n21697 );
and ( n24795 , n24789 , n24794 );
and ( n24796 , n24775 , n24794 );
or ( n24797 , n24790 , n24795 , n24796 );
and ( n24798 , n24746 , n24797 );
and ( n24799 , n24732 , n24797 );
or ( n24800 , n24747 , n24798 , n24799 );
xor ( n24801 , n24591 , n24593 );
xor ( n24802 , n24801 , n24596 );
and ( n24803 , n24800 , n24802 );
xor ( n24804 , n24658 , n24663 );
and ( n24805 , n24460 , n21496 );
and ( n24806 , n24213 , n21494 );
nor ( n24807 , n24805 , n24806 );
xnor ( n24808 , n24807 , n21506 );
xor ( n24809 , n20920 , n21075 );
buf ( n24810 , n24809 );
buf ( n24811 , n24810 );
buf ( n24812 , n24811 );
and ( n24813 , n24812 , n21513 );
and ( n24814 , n24808 , n24813 );
and ( n24815 , n24804 , n24814 );
and ( n24816 , n24213 , n21496 );
and ( n24817 , n23949 , n21494 );
nor ( n24818 , n24816 , n24817 );
xnor ( n24819 , n24818 , n21506 );
and ( n24820 , n24814 , n24819 );
and ( n24821 , n24804 , n24819 );
or ( n24822 , n24815 , n24820 , n24821 );
and ( n24823 , n21511 , n21582 );
and ( n24824 , n21599 , n21580 );
nor ( n24825 , n24823 , n24824 );
xnor ( n24826 , n24825 , n21588 );
and ( n24827 , n24822 , n24826 );
and ( n24828 , n21616 , n21783 );
and ( n24829 , n21606 , n21781 );
nor ( n24830 , n24828 , n24829 );
xnor ( n24831 , n24830 , n21793 );
and ( n24832 , n24826 , n24831 );
and ( n24833 , n24822 , n24831 );
or ( n24834 , n24827 , n24832 , n24833 );
and ( n24835 , n21756 , n21707 );
and ( n24836 , n21519 , n21705 );
nor ( n24837 , n24835 , n24836 );
xnor ( n24838 , n24837 , n21717 );
and ( n24839 , n24834 , n24838 );
xor ( n24840 , n24672 , n24676 );
xor ( n24841 , n24840 , n24681 );
and ( n24842 , n24838 , n24841 );
and ( n24843 , n24834 , n24841 );
or ( n24844 , n24839 , n24842 , n24843 );
and ( n24845 , n22089 , n21663 );
and ( n24846 , n21777 , n21661 );
nor ( n24847 , n24845 , n24846 );
xnor ( n24848 , n24847 , n21673 );
and ( n24849 , n24844 , n24848 );
xor ( n24850 , n24641 , n24645 );
xor ( n24851 , n24850 , n24650 );
and ( n24852 , n24848 , n24851 );
and ( n24853 , n24844 , n24851 );
or ( n24854 , n24849 , n24852 , n24853 );
xor ( n24855 , n24653 , n24694 );
xor ( n24856 , n24855 , n24699 );
and ( n24857 , n24854 , n24856 );
xor ( n24858 , n24525 , n24529 );
xor ( n24859 , n24858 , n24532 );
and ( n24860 , n24856 , n24859 );
and ( n24861 , n24854 , n24859 );
or ( n24862 , n24857 , n24860 , n24861 );
and ( n24863 , n24802 , n24862 );
and ( n24864 , n24800 , n24862 );
or ( n24865 , n24803 , n24863 , n24864 );
and ( n24866 , n24730 , n24865 );
xor ( n24867 , n24607 , n24608 );
xor ( n24868 , n24867 , n24705 );
and ( n24869 , n24865 , n24868 );
and ( n24870 , n24730 , n24868 );
or ( n24871 , n24866 , n24869 , n24870 );
and ( n24872 , n24728 , n24871 );
xor ( n24873 , n24602 , n24604 );
xor ( n24874 , n24873 , n24708 );
and ( n24875 , n24871 , n24874 );
and ( n24876 , n24728 , n24874 );
or ( n24877 , n24872 , n24875 , n24876 );
and ( n24878 , n24726 , n24877 );
xor ( n24879 , n24420 , n24551 );
xor ( n24880 , n24879 , n24711 );
and ( n24881 , n24877 , n24880 );
and ( n24882 , n24726 , n24880 );
or ( n24883 , n24878 , n24881 , n24882 );
xor ( n24884 , n24390 , n24714 );
xor ( n24885 , n24884 , n24717 );
and ( n24886 , n24883 , n24885 );
xor ( n24887 , n24883 , n24885 );
xor ( n24888 , n24726 , n24877 );
xor ( n24889 , n24888 , n24880 );
xor ( n24890 , n24728 , n24871 );
xor ( n24891 , n24890 , n24874 );
xor ( n24892 , n24611 , n24613 );
xor ( n24893 , n24892 , n24616 );
and ( n24894 , n21226 , n22114 );
and ( n24895 , n21241 , n22112 );
nor ( n24896 , n24894 , n24895 );
xnor ( n24897 , n24896 , n22124 );
and ( n24898 , n21788 , n21139 );
and ( n24899 , n21574 , n21137 );
nor ( n24900 , n24898 , n24899 );
xnor ( n24901 , n24900 , n21221 );
and ( n24902 , n24897 , n24901 );
xor ( n24903 , n24684 , n24688 );
xor ( n24904 , n24903 , n24691 );
and ( n24905 , n24901 , n24904 );
and ( n24906 , n24897 , n24904 );
or ( n24907 , n24902 , n24905 , n24906 );
and ( n24908 , n24893 , n24907 );
and ( n24909 , n21519 , n21687 );
and ( n24910 , n21534 , n21685 );
nor ( n24911 , n24909 , n24910 );
xnor ( n24912 , n24911 , n21697 );
and ( n24913 , n21545 , n21260 );
and ( n24914 , n21486 , n21258 );
nor ( n24915 , n24913 , n24914 );
xnor ( n24916 , n24915 , n21270 );
and ( n24917 , n24912 , n24916 );
xor ( n24918 , n24751 , n24755 );
xor ( n24919 , n24918 , n24760 );
and ( n24920 , n24916 , n24919 );
and ( n24921 , n24912 , n24919 );
or ( n24922 , n24917 , n24920 , n24921 );
and ( n24923 , n21744 , n21663 );
and ( n24924 , n22089 , n21661 );
nor ( n24925 , n24923 , n24924 );
xnor ( n24926 , n24925 , n21673 );
and ( n24927 , n24922 , n24926 );
and ( n24928 , n21534 , n21687 );
and ( n24929 , n21731 , n21685 );
nor ( n24930 , n24928 , n24929 );
xnor ( n24931 , n24930 , n21697 );
and ( n24932 , n24926 , n24931 );
and ( n24933 , n24922 , n24931 );
or ( n24934 , n24927 , n24932 , n24933 );
xor ( n24935 , n24736 , n24740 );
xor ( n24936 , n24935 , n24743 );
and ( n24937 , n24934 , n24936 );
xor ( n24938 , n24775 , n24789 );
xor ( n24939 , n24938 , n24794 );
and ( n24940 , n24936 , n24939 );
and ( n24941 , n24934 , n24939 );
or ( n24942 , n24937 , n24940 , n24941 );
and ( n24943 , n24907 , n24942 );
and ( n24944 , n24893 , n24942 );
or ( n24945 , n24908 , n24943 , n24944 );
xor ( n24946 , n24619 , n24621 );
xor ( n24947 , n24946 , n24702 );
and ( n24948 , n24945 , n24947 );
xor ( n24949 , n24732 , n24746 );
xor ( n24950 , n24949 , n24797 );
xor ( n24951 , n24854 , n24856 );
xor ( n24952 , n24951 , n24859 );
and ( n24953 , n24950 , n24952 );
and ( n24954 , n21265 , n22114 );
and ( n24955 , n21226 , n22112 );
nor ( n24956 , n24954 , n24955 );
xnor ( n24957 , n24956 , n22124 );
and ( n24958 , n21777 , n21139 );
and ( n24959 , n21788 , n21137 );
nor ( n24960 , n24958 , n24959 );
xnor ( n24961 , n24960 , n21221 );
and ( n24962 , n24957 , n24961 );
xor ( n24963 , n24779 , n24783 );
xor ( n24964 , n24963 , n24786 );
and ( n24965 , n24961 , n24964 );
and ( n24966 , n24957 , n24964 );
or ( n24967 , n24962 , n24965 , n24966 );
xor ( n24968 , n24844 , n24848 );
xor ( n24969 , n24968 , n24851 );
and ( n24970 , n24967 , n24969 );
xor ( n24971 , n24897 , n24901 );
xor ( n24972 , n24971 , n24904 );
and ( n24973 , n24969 , n24972 );
and ( n24974 , n24967 , n24972 );
or ( n24975 , n24970 , n24973 , n24974 );
and ( n24976 , n24952 , n24975 );
and ( n24977 , n24950 , n24975 );
or ( n24978 , n24953 , n24976 , n24977 );
and ( n24979 , n24947 , n24978 );
and ( n24980 , n24945 , n24978 );
or ( n24981 , n24948 , n24979 , n24980 );
xor ( n24982 , n24730 , n24865 );
xor ( n24983 , n24982 , n24868 );
and ( n24984 , n24981 , n24983 );
xor ( n24985 , n24800 , n24802 );
xor ( n24986 , n24985 , n24862 );
and ( n24987 , n23320 , n21739 );
and ( n24988 , n23074 , n21737 );
nor ( n24989 , n24987 , n24988 );
xnor ( n24990 , n24989 , n21749 );
and ( n24991 , n23503 , n21529 );
and ( n24992 , n23351 , n21527 );
nor ( n24993 , n24991 , n24992 );
xnor ( n24994 , n24993 , n21539 );
and ( n24995 , n24990 , n24994 );
and ( n24996 , n23887 , n21625 );
and ( n24997 , n23651 , n21623 );
nor ( n24998 , n24996 , n24997 );
xnor ( n24999 , n24998 , n21635 );
and ( n25000 , n24994 , n24999 );
and ( n25001 , n24990 , n24999 );
or ( n25002 , n24995 , n25000 , n25001 );
and ( n25003 , n21501 , n21236 );
and ( n25004 , n21630 , n21234 );
nor ( n25005 , n25003 , n25004 );
xnor ( n25006 , n25005 , n21246 );
and ( n25007 , n25002 , n25006 );
xor ( n25008 , n24654 , n24664 );
xor ( n25009 , n25008 , n24669 );
and ( n25010 , n25006 , n25009 );
and ( n25011 , n25002 , n25009 );
or ( n25012 , n25007 , n25010 , n25011 );
and ( n25013 , n21630 , n21236 );
and ( n25014 , n21645 , n21234 );
nor ( n25015 , n25013 , n25014 );
xnor ( n25016 , n25015 , n21246 );
and ( n25017 , n25012 , n25016 );
xor ( n25018 , n24763 , n24767 );
xor ( n25019 , n25018 , n24772 );
and ( n25020 , n25016 , n25019 );
and ( n25021 , n25012 , n25019 );
or ( n25022 , n25017 , n25020 , n25021 );
and ( n25023 , n21241 , n22032 );
and ( n25024 , n21566 , n22029 );
nor ( n25025 , n25023 , n25024 );
xnor ( n25026 , n25025 , n22027 );
and ( n25027 , n21574 , n21414 );
and ( n25028 , n21252 , n21412 );
nor ( n25029 , n25027 , n25028 );
xnor ( n25030 , n25029 , n21480 );
and ( n25031 , n25026 , n25030 );
xor ( n25032 , n24834 , n24838 );
xor ( n25033 , n25032 , n24841 );
and ( n25034 , n25030 , n25033 );
and ( n25035 , n25026 , n25033 );
or ( n25036 , n25031 , n25034 , n25035 );
and ( n25037 , n25022 , n25036 );
xor ( n25038 , n24934 , n24936 );
xor ( n25039 , n25038 , n24939 );
and ( n25040 , n25036 , n25039 );
and ( n25041 , n25022 , n25039 );
or ( n25042 , n25037 , n25040 , n25041 );
xor ( n25043 , n24893 , n24907 );
xor ( n25044 , n25043 , n24942 );
and ( n25045 , n25042 , n25044 );
xor ( n25046 , n24967 , n24969 );
xor ( n25047 , n25046 , n24972 );
and ( n25048 , n24631 , n21496 );
and ( n25049 , n24460 , n21494 );
nor ( n25050 , n25048 , n25049 );
xnor ( n25051 , n25050 , n21506 );
and ( n25052 , n24812 , n21551 );
and ( n25053 , n24662 , n21549 );
nor ( n25054 , n25052 , n25053 );
xnor ( n25055 , n25054 , n21557 );
and ( n25056 , n25051 , n25055 );
xor ( n25057 , n20948 , n21073 );
buf ( n25058 , n25057 );
buf ( n25059 , n25058 );
buf ( n25060 , n25059 );
and ( n25061 , n25060 , n21513 );
and ( n25062 , n25055 , n25061 );
and ( n25063 , n25051 , n25061 );
or ( n25064 , n25056 , n25062 , n25063 );
and ( n25065 , n23651 , n21529 );
and ( n25066 , n23503 , n21527 );
nor ( n25067 , n25065 , n25066 );
xnor ( n25068 , n25067 , n21539 );
and ( n25069 , n25064 , n25068 );
and ( n25070 , n23949 , n21625 );
and ( n25071 , n23887 , n21623 );
nor ( n25072 , n25070 , n25071 );
xnor ( n25073 , n25072 , n21635 );
and ( n25074 , n25068 , n25073 );
and ( n25075 , n25064 , n25073 );
or ( n25076 , n25069 , n25074 , n25075 );
and ( n25077 , n21486 , n21236 );
and ( n25078 , n21501 , n21234 );
nor ( n25079 , n25077 , n25078 );
xnor ( n25080 , n25079 , n21246 );
and ( n25081 , n25076 , n25080 );
xor ( n25082 , n24804 , n24814 );
xor ( n25083 , n25082 , n24819 );
and ( n25084 , n25080 , n25083 );
and ( n25085 , n25076 , n25083 );
or ( n25086 , n25081 , n25084 , n25085 );
and ( n25087 , n24662 , n21551 );
and ( n25088 , n24631 , n21549 );
nor ( n25089 , n25087 , n25088 );
xnor ( n25090 , n25089 , n21557 );
xor ( n25091 , n24808 , n24813 );
xor ( n25092 , n25090 , n25091 );
and ( n25093 , n23074 , n21783 );
and ( n25094 , n22813 , n21781 );
nor ( n25095 , n25093 , n25094 );
xnor ( n25096 , n25095 , n21793 );
and ( n25097 , n25092 , n25096 );
and ( n25098 , n23351 , n21739 );
and ( n25099 , n23320 , n21737 );
nor ( n25100 , n25098 , n25099 );
xnor ( n25101 , n25100 , n21749 );
and ( n25102 , n25096 , n25101 );
and ( n25103 , n25092 , n25101 );
or ( n25104 , n25097 , n25102 , n25103 );
and ( n25105 , n21599 , n21260 );
and ( n25106 , n21545 , n21258 );
nor ( n25107 , n25105 , n25106 );
xnor ( n25108 , n25107 , n21270 );
and ( n25109 , n25104 , n25108 );
xor ( n25110 , n24990 , n24994 );
xor ( n25111 , n25110 , n24999 );
and ( n25112 , n25108 , n25111 );
and ( n25113 , n25104 , n25111 );
or ( n25114 , n25109 , n25112 , n25113 );
and ( n25115 , n25086 , n25114 );
and ( n25116 , n21731 , n21663 );
and ( n25117 , n21744 , n21661 );
nor ( n25118 , n25116 , n25117 );
xnor ( n25119 , n25118 , n21673 );
and ( n25120 , n25114 , n25119 );
and ( n25121 , n25086 , n25119 );
or ( n25122 , n25115 , n25120 , n25121 );
and ( n25123 , n25090 , n25091 );
and ( n25124 , n21606 , n21582 );
and ( n25125 , n21511 , n21580 );
nor ( n25126 , n25124 , n25125 );
xnor ( n25127 , n25126 , n21588 );
and ( n25128 , n25123 , n25127 );
and ( n25129 , n22813 , n21783 );
and ( n25130 , n21616 , n21781 );
nor ( n25131 , n25129 , n25130 );
xnor ( n25132 , n25131 , n21793 );
and ( n25133 , n25127 , n25132 );
and ( n25134 , n25123 , n25132 );
or ( n25135 , n25128 , n25133 , n25134 );
and ( n25136 , n21645 , n21707 );
and ( n25137 , n21756 , n21705 );
nor ( n25138 , n25136 , n25137 );
xnor ( n25139 , n25138 , n21717 );
and ( n25140 , n25135 , n25139 );
xor ( n25141 , n24822 , n24826 );
xor ( n25142 , n25141 , n24831 );
and ( n25143 , n25139 , n25142 );
and ( n25144 , n25135 , n25142 );
or ( n25145 , n25140 , n25143 , n25144 );
and ( n25146 , n25122 , n25145 );
xor ( n25147 , n25012 , n25016 );
xor ( n25148 , n25147 , n25019 );
and ( n25149 , n25145 , n25148 );
and ( n25150 , n25122 , n25148 );
or ( n25151 , n25146 , n25149 , n25150 );
and ( n25152 , n25047 , n25151 );
and ( n25153 , n21788 , n21414 );
and ( n25154 , n21574 , n21412 );
nor ( n25155 , n25153 , n25154 );
xnor ( n25156 , n25155 , n21480 );
and ( n25157 , n22089 , n21139 );
and ( n25158 , n21777 , n21137 );
nor ( n25159 , n25157 , n25158 );
xnor ( n25160 , n25159 , n21221 );
and ( n25161 , n25156 , n25160 );
xor ( n25162 , n25002 , n25006 );
xor ( n25163 , n25162 , n25009 );
and ( n25164 , n25160 , n25163 );
and ( n25165 , n25156 , n25163 );
or ( n25166 , n25161 , n25164 , n25165 );
and ( n25167 , n24460 , n21625 );
and ( n25168 , n24213 , n21623 );
nor ( n25169 , n25167 , n25168 );
xnor ( n25170 , n25169 , n21635 );
and ( n25171 , n25060 , n21551 );
and ( n25172 , n24812 , n21549 );
nor ( n25173 , n25171 , n25172 );
xnor ( n25174 , n25173 , n21557 );
and ( n25175 , n25170 , n25174 );
xor ( n25176 , n20971 , n21071 );
buf ( n25177 , n25176 );
buf ( n25178 , n25177 );
buf ( n25179 , n25178 );
and ( n25180 , n25179 , n21513 );
and ( n25181 , n25174 , n25180 );
and ( n25182 , n25170 , n25180 );
or ( n25183 , n25175 , n25181 , n25182 );
and ( n25184 , n23887 , n21529 );
and ( n25185 , n23651 , n21527 );
nor ( n25186 , n25184 , n25185 );
xnor ( n25187 , n25186 , n21539 );
and ( n25188 , n25183 , n25187 );
and ( n25189 , n24213 , n21625 );
and ( n25190 , n23949 , n21623 );
nor ( n25191 , n25189 , n25190 );
xnor ( n25192 , n25191 , n21635 );
and ( n25193 , n25187 , n25192 );
and ( n25194 , n25183 , n25192 );
or ( n25195 , n25188 , n25193 , n25194 );
and ( n25196 , n21511 , n21260 );
and ( n25197 , n21599 , n21258 );
nor ( n25198 , n25196 , n25197 );
xnor ( n25199 , n25198 , n21270 );
and ( n25200 , n25195 , n25199 );
and ( n25201 , n21616 , n21582 );
and ( n25202 , n21606 , n21580 );
nor ( n25203 , n25201 , n25202 );
xnor ( n25204 , n25203 , n21588 );
and ( n25205 , n25199 , n25204 );
and ( n25206 , n25195 , n25204 );
or ( n25207 , n25200 , n25205 , n25206 );
and ( n25208 , n21756 , n21687 );
and ( n25209 , n21519 , n21685 );
nor ( n25210 , n25208 , n25209 );
xnor ( n25211 , n25210 , n21697 );
and ( n25212 , n25207 , n25211 );
and ( n25213 , n21630 , n21707 );
and ( n25214 , n21645 , n21705 );
nor ( n25215 , n25213 , n25214 );
xnor ( n25216 , n25215 , n21717 );
and ( n25217 , n25211 , n25216 );
and ( n25218 , n25207 , n25216 );
or ( n25219 , n25212 , n25217 , n25218 );
and ( n25220 , n21252 , n22114 );
and ( n25221 , n21265 , n22112 );
nor ( n25222 , n25220 , n25221 );
xnor ( n25223 , n25222 , n22124 );
and ( n25224 , n25219 , n25223 );
xor ( n25225 , n24912 , n24916 );
xor ( n25226 , n25225 , n24919 );
and ( n25227 , n25223 , n25226 );
and ( n25228 , n25219 , n25226 );
or ( n25229 , n25224 , n25227 , n25228 );
and ( n25230 , n25166 , n25229 );
xor ( n25231 , n24957 , n24961 );
xor ( n25232 , n25231 , n24964 );
and ( n25233 , n25229 , n25232 );
and ( n25234 , n25166 , n25232 );
or ( n25235 , n25230 , n25233 , n25234 );
and ( n25236 , n25151 , n25235 );
and ( n25237 , n25047 , n25235 );
or ( n25238 , n25152 , n25236 , n25237 );
and ( n25239 , n25044 , n25238 );
and ( n25240 , n25042 , n25238 );
or ( n25241 , n25045 , n25239 , n25240 );
and ( n25242 , n24986 , n25241 );
xor ( n25243 , n24945 , n24947 );
xor ( n25244 , n25243 , n24978 );
and ( n25245 , n25241 , n25244 );
and ( n25246 , n24986 , n25244 );
or ( n25247 , n25242 , n25245 , n25246 );
and ( n25248 , n24983 , n25247 );
and ( n25249 , n24981 , n25247 );
or ( n25250 , n24984 , n25248 , n25249 );
and ( n25251 , n24891 , n25250 );
xor ( n25252 , n24891 , n25250 );
xor ( n25253 , n24981 , n24983 );
xor ( n25254 , n25253 , n25247 );
xor ( n25255 , n24950 , n24952 );
xor ( n25256 , n25255 , n24975 );
and ( n25257 , n23320 , n21783 );
and ( n25258 , n23074 , n21781 );
nor ( n25259 , n25257 , n25258 );
xnor ( n25260 , n25259 , n21793 );
and ( n25261 , n23503 , n21739 );
and ( n25262 , n23351 , n21737 );
nor ( n25263 , n25261 , n25262 );
xnor ( n25264 , n25263 , n21749 );
and ( n25265 , n25260 , n25264 );
xor ( n25266 , n25051 , n25055 );
xor ( n25267 , n25266 , n25061 );
and ( n25268 , n25264 , n25267 );
and ( n25269 , n25260 , n25267 );
or ( n25270 , n25265 , n25268 , n25269 );
and ( n25271 , n21545 , n21236 );
and ( n25272 , n21486 , n21234 );
nor ( n25273 , n25271 , n25272 );
xnor ( n25274 , n25273 , n21246 );
and ( n25275 , n25270 , n25274 );
xor ( n25276 , n25064 , n25068 );
xor ( n25277 , n25276 , n25073 );
and ( n25278 , n25274 , n25277 );
and ( n25279 , n25270 , n25277 );
or ( n25280 , n25275 , n25278 , n25279 );
and ( n25281 , n21534 , n21663 );
and ( n25282 , n21731 , n21661 );
nor ( n25283 , n25281 , n25282 );
xnor ( n25284 , n25283 , n21673 );
and ( n25285 , n25280 , n25284 );
xor ( n25286 , n25123 , n25127 );
xor ( n25287 , n25286 , n25132 );
and ( n25288 , n25284 , n25287 );
and ( n25289 , n25280 , n25287 );
or ( n25290 , n25285 , n25288 , n25289 );
and ( n25291 , n21226 , n22032 );
and ( n25292 , n21241 , n22029 );
nor ( n25293 , n25291 , n25292 );
xnor ( n25294 , n25293 , n22027 );
and ( n25295 , n25290 , n25294 );
xor ( n25296 , n25135 , n25139 );
xor ( n25297 , n25296 , n25142 );
and ( n25298 , n25294 , n25297 );
and ( n25299 , n25290 , n25297 );
or ( n25300 , n25295 , n25298 , n25299 );
xor ( n25301 , n24922 , n24926 );
xor ( n25302 , n25301 , n24931 );
and ( n25303 , n25300 , n25302 );
xor ( n25304 , n25026 , n25030 );
xor ( n25305 , n25304 , n25033 );
and ( n25306 , n25302 , n25305 );
and ( n25307 , n25300 , n25305 );
or ( n25308 , n25303 , n25306 , n25307 );
xor ( n25309 , n25022 , n25036 );
xor ( n25310 , n25309 , n25039 );
and ( n25311 , n25308 , n25310 );
xor ( n25312 , n25166 , n25229 );
xor ( n25313 , n25312 , n25232 );
xor ( n25314 , n25300 , n25302 );
xor ( n25315 , n25314 , n25305 );
and ( n25316 , n25313 , n25315 );
and ( n25317 , n25310 , n25316 );
and ( n25318 , n25308 , n25316 );
or ( n25319 , n25311 , n25317 , n25318 );
and ( n25320 , n25256 , n25319 );
xor ( n25321 , n25042 , n25044 );
xor ( n25322 , n25321 , n25238 );
and ( n25323 , n25319 , n25322 );
and ( n25324 , n25256 , n25322 );
or ( n25325 , n25320 , n25323 , n25324 );
xor ( n25326 , n24986 , n25241 );
xor ( n25327 , n25326 , n25244 );
and ( n25328 , n25325 , n25327 );
xor ( n25329 , n25122 , n25145 );
xor ( n25330 , n25329 , n25148 );
and ( n25331 , n24631 , n21625 );
and ( n25332 , n24460 , n21623 );
nor ( n25333 , n25331 , n25332 );
xnor ( n25334 , n25333 , n21635 );
and ( n25335 , n25179 , n21551 );
and ( n25336 , n25060 , n21549 );
nor ( n25337 , n25335 , n25336 );
xnor ( n25338 , n25337 , n21557 );
and ( n25339 , n25334 , n25338 );
xor ( n25340 , n20993 , n21069 );
buf ( n25341 , n25340 );
buf ( n25342 , n25341 );
buf ( n25343 , n25342 );
and ( n25344 , n25343 , n21513 );
and ( n25345 , n25338 , n25344 );
and ( n25346 , n25334 , n25344 );
or ( n25347 , n25339 , n25345 , n25346 );
and ( n25348 , n23949 , n21529 );
and ( n25349 , n23887 , n21527 );
nor ( n25350 , n25348 , n25349 );
xnor ( n25351 , n25350 , n21539 );
and ( n25352 , n25347 , n25351 );
and ( n25353 , n24662 , n21496 );
and ( n25354 , n24631 , n21494 );
nor ( n25355 , n25353 , n25354 );
xnor ( n25356 , n25355 , n21506 );
and ( n25357 , n25351 , n25356 );
and ( n25358 , n25347 , n25356 );
or ( n25359 , n25352 , n25357 , n25358 );
and ( n25360 , n21606 , n21260 );
and ( n25361 , n21511 , n21258 );
nor ( n25362 , n25360 , n25361 );
xnor ( n25363 , n25362 , n21270 );
and ( n25364 , n25359 , n25363 );
and ( n25365 , n22813 , n21582 );
and ( n25366 , n21616 , n21580 );
nor ( n25367 , n25365 , n25366 );
xnor ( n25368 , n25367 , n21588 );
and ( n25369 , n25363 , n25368 );
and ( n25370 , n25359 , n25368 );
or ( n25371 , n25364 , n25369 , n25370 );
and ( n25372 , n21501 , n21707 );
and ( n25373 , n21630 , n21705 );
nor ( n25374 , n25372 , n25373 );
xnor ( n25375 , n25374 , n21717 );
and ( n25376 , n25371 , n25375 );
xor ( n25377 , n25092 , n25096 );
xor ( n25378 , n25377 , n25101 );
and ( n25379 , n25375 , n25378 );
and ( n25380 , n25371 , n25378 );
or ( n25381 , n25376 , n25379 , n25380 );
and ( n25382 , n21777 , n21414 );
and ( n25383 , n21788 , n21412 );
nor ( n25384 , n25382 , n25383 );
xnor ( n25385 , n25384 , n21480 );
and ( n25386 , n25381 , n25385 );
xor ( n25387 , n25076 , n25080 );
xor ( n25388 , n25387 , n25083 );
and ( n25389 , n25385 , n25388 );
and ( n25390 , n25381 , n25388 );
or ( n25391 , n25386 , n25389 , n25390 );
xor ( n25392 , n25086 , n25114 );
xor ( n25393 , n25392 , n25119 );
and ( n25394 , n25391 , n25393 );
xor ( n25395 , n25156 , n25160 );
xor ( n25396 , n25395 , n25163 );
and ( n25397 , n25393 , n25396 );
and ( n25398 , n25391 , n25396 );
or ( n25399 , n25394 , n25397 , n25398 );
and ( n25400 , n25330 , n25399 );
xor ( n25401 , n25219 , n25223 );
xor ( n25402 , n25401 , n25226 );
and ( n25403 , n21574 , n22114 );
and ( n25404 , n21252 , n22112 );
nor ( n25405 , n25403 , n25404 );
xnor ( n25406 , n25405 , n22124 );
and ( n25407 , n21744 , n21139 );
and ( n25408 , n22089 , n21137 );
nor ( n25409 , n25407 , n25408 );
xnor ( n25410 , n25409 , n21221 );
and ( n25411 , n25406 , n25410 );
xor ( n25412 , n25104 , n25108 );
xor ( n25413 , n25412 , n25111 );
and ( n25414 , n25410 , n25413 );
and ( n25415 , n25406 , n25413 );
or ( n25416 , n25411 , n25414 , n25415 );
and ( n25417 , n25402 , n25416 );
and ( n25418 , n21265 , n22032 );
and ( n25419 , n21226 , n22029 );
nor ( n25420 , n25418 , n25419 );
xnor ( n25421 , n25420 , n22027 );
xor ( n25422 , n25207 , n25211 );
xor ( n25423 , n25422 , n25216 );
and ( n25424 , n25421 , n25423 );
and ( n25425 , n21519 , n21663 );
and ( n25426 , n21534 , n21661 );
nor ( n25427 , n25425 , n25426 );
xnor ( n25428 , n25427 , n21673 );
and ( n25429 , n21645 , n21687 );
and ( n25430 , n21756 , n21685 );
nor ( n25431 , n25429 , n25430 );
xnor ( n25432 , n25431 , n21697 );
and ( n25433 , n25428 , n25432 );
xor ( n25434 , n25195 , n25199 );
xor ( n25435 , n25434 , n25204 );
and ( n25436 , n25432 , n25435 );
and ( n25437 , n25428 , n25435 );
or ( n25438 , n25433 , n25436 , n25437 );
and ( n25439 , n25423 , n25438 );
and ( n25440 , n25421 , n25438 );
or ( n25441 , n25424 , n25439 , n25440 );
and ( n25442 , n25416 , n25441 );
and ( n25443 , n25402 , n25441 );
or ( n25444 , n25417 , n25442 , n25443 );
and ( n25445 , n25399 , n25444 );
and ( n25446 , n25330 , n25444 );
or ( n25447 , n25400 , n25445 , n25446 );
xor ( n25448 , n25047 , n25151 );
xor ( n25449 , n25448 , n25235 );
and ( n25450 , n25447 , n25449 );
xor ( n25451 , n25313 , n25315 );
xor ( n25452 , n25391 , n25393 );
xor ( n25453 , n25452 , n25396 );
xor ( n25454 , n25381 , n25385 );
xor ( n25455 , n25454 , n25388 );
xor ( n25456 , n25406 , n25410 );
xor ( n25457 , n25456 , n25413 );
and ( n25458 , n25455 , n25457 );
and ( n25459 , n21534 , n21139 );
and ( n25460 , n21731 , n21137 );
nor ( n25461 , n25459 , n25460 );
xnor ( n25462 , n25461 , n21221 );
and ( n25463 , n21630 , n21687 );
and ( n25464 , n21645 , n21685 );
nor ( n25465 , n25463 , n25464 );
xnor ( n25466 , n25465 , n21697 );
and ( n25467 , n25462 , n25466 );
and ( n25468 , n23351 , n21783 );
and ( n25469 , n23320 , n21781 );
nor ( n25470 , n25468 , n25469 );
xnor ( n25471 , n25470 , n21793 );
and ( n25472 , n23651 , n21739 );
and ( n25473 , n23503 , n21737 );
nor ( n25474 , n25472 , n25473 );
xnor ( n25475 , n25474 , n21749 );
and ( n25476 , n25471 , n25475 );
xor ( n25477 , n25170 , n25174 );
xor ( n25478 , n25477 , n25180 );
and ( n25479 , n25475 , n25478 );
and ( n25480 , n25471 , n25478 );
or ( n25481 , n25476 , n25479 , n25480 );
and ( n25482 , n21599 , n21236 );
and ( n25483 , n21545 , n21234 );
nor ( n25484 , n25482 , n25483 );
xnor ( n25485 , n25484 , n21246 );
xor ( n25486 , n25481 , n25485 );
xor ( n25487 , n25183 , n25187 );
xor ( n25488 , n25487 , n25192 );
xor ( n25489 , n25486 , n25488 );
and ( n25490 , n25466 , n25489 );
and ( n25491 , n25462 , n25489 );
or ( n25492 , n25467 , n25490 , n25491 );
xor ( n25493 , n25428 , n25432 );
xor ( n25494 , n25493 , n25435 );
and ( n25495 , n25492 , n25494 );
and ( n25496 , n25481 , n25485 );
and ( n25497 , n25485 , n25488 );
and ( n25498 , n25481 , n25488 );
or ( n25499 , n25496 , n25497 , n25498 );
and ( n25500 , n21731 , n21139 );
and ( n25501 , n21744 , n21137 );
nor ( n25502 , n25500 , n25501 );
xnor ( n25503 , n25502 , n21221 );
xor ( n25504 , n25499 , n25503 );
xor ( n25505 , n25270 , n25274 );
xor ( n25506 , n25505 , n25277 );
xor ( n25507 , n25504 , n25506 );
and ( n25508 , n25494 , n25507 );
and ( n25509 , n25492 , n25507 );
or ( n25510 , n25495 , n25508 , n25509 );
and ( n25511 , n25457 , n25510 );
and ( n25512 , n25455 , n25510 );
or ( n25513 , n25458 , n25511 , n25512 );
and ( n25514 , n25453 , n25513 );
xor ( n25515 , n25402 , n25416 );
xor ( n25516 , n25515 , n25441 );
and ( n25517 , n25513 , n25516 );
and ( n25518 , n25453 , n25516 );
or ( n25519 , n25514 , n25517 , n25518 );
and ( n25520 , n25451 , n25519 );
xor ( n25521 , n25330 , n25399 );
xor ( n25522 , n25521 , n25444 );
and ( n25523 , n25519 , n25522 );
and ( n25524 , n25451 , n25522 );
or ( n25525 , n25520 , n25523 , n25524 );
and ( n25526 , n25449 , n25525 );
and ( n25527 , n25447 , n25525 );
or ( n25528 , n25450 , n25526 , n25527 );
xor ( n25529 , n25256 , n25319 );
xor ( n25530 , n25529 , n25322 );
and ( n25531 , n25528 , n25530 );
xor ( n25532 , n25308 , n25310 );
xor ( n25533 , n25532 , n25316 );
xor ( n25534 , n25447 , n25449 );
xor ( n25535 , n25534 , n25525 );
and ( n25536 , n25533 , n25535 );
and ( n25537 , n25179 , n21496 );
and ( n25538 , n25060 , n21494 );
nor ( n25539 , n25537 , n25538 );
xnor ( n25540 , n25539 , n21506 );
xor ( n25541 , n21010 , n21067 );
buf ( n25542 , n25541 );
buf ( n25543 , n25542 );
buf ( n25544 , n25543 );
and ( n25545 , n25544 , n21551 );
and ( n25546 , n25343 , n21549 );
nor ( n25547 , n25545 , n25546 );
xnor ( n25548 , n25547 , n21557 );
and ( n25549 , n25540 , n25548 );
xor ( n25550 , n21026 , n21065 );
buf ( n25551 , n25550 );
buf ( n25552 , n25551 );
buf ( n25553 , n25552 );
and ( n25554 , n25553 , n21513 );
and ( n25555 , n25548 , n25554 );
and ( n25556 , n25540 , n25554 );
or ( n25557 , n25549 , n25555 , n25556 );
and ( n25558 , n24460 , n21529 );
and ( n25559 , n24213 , n21527 );
nor ( n25560 , n25558 , n25559 );
xnor ( n25561 , n25560 , n21539 );
and ( n25562 , n25557 , n25561 );
and ( n25563 , n24662 , n21625 );
and ( n25564 , n24631 , n21623 );
nor ( n25565 , n25563 , n25564 );
xnor ( n25566 , n25565 , n21635 );
and ( n25567 , n25561 , n25566 );
and ( n25568 , n25557 , n25566 );
or ( n25569 , n25562 , n25567 , n25568 );
and ( n25570 , n23887 , n21739 );
and ( n25571 , n23651 , n21737 );
nor ( n25572 , n25570 , n25571 );
xnor ( n25573 , n25572 , n21749 );
and ( n25574 , n25569 , n25573 );
xor ( n25575 , n25334 , n25338 );
xor ( n25576 , n25575 , n25344 );
and ( n25577 , n25573 , n25576 );
and ( n25578 , n25569 , n25576 );
or ( n25579 , n25574 , n25577 , n25578 );
and ( n25580 , n21616 , n21260 );
and ( n25581 , n21606 , n21258 );
nor ( n25582 , n25580 , n25581 );
xnor ( n25583 , n25582 , n21270 );
and ( n25584 , n25579 , n25583 );
xor ( n25585 , n25347 , n25351 );
xor ( n25586 , n25585 , n25356 );
and ( n25587 , n25583 , n25586 );
and ( n25588 , n25579 , n25586 );
or ( n25589 , n25584 , n25587 , n25588 );
and ( n25590 , n21486 , n21707 );
and ( n25591 , n21501 , n21705 );
nor ( n25592 , n25590 , n25591 );
xnor ( n25593 , n25592 , n21717 );
and ( n25594 , n25589 , n25593 );
xor ( n25595 , n25260 , n25264 );
xor ( n25596 , n25595 , n25267 );
and ( n25597 , n25593 , n25596 );
and ( n25598 , n25589 , n25596 );
or ( n25599 , n25594 , n25597 , n25598 );
and ( n25600 , n21788 , n22114 );
and ( n25601 , n21574 , n22112 );
nor ( n25602 , n25600 , n25601 );
xnor ( n25603 , n25602 , n22124 );
and ( n25604 , n25599 , n25603 );
and ( n25605 , n22089 , n21414 );
and ( n25606 , n21777 , n21412 );
nor ( n25607 , n25605 , n25606 );
xnor ( n25608 , n25607 , n21480 );
and ( n25609 , n25603 , n25608 );
and ( n25610 , n25599 , n25608 );
or ( n25611 , n25604 , n25609 , n25610 );
and ( n25612 , n25499 , n25503 );
and ( n25613 , n25503 , n25506 );
and ( n25614 , n25499 , n25506 );
or ( n25615 , n25612 , n25613 , n25614 );
and ( n25616 , n25611 , n25615 );
xor ( n25617 , n25280 , n25284 );
xor ( n25618 , n25617 , n25287 );
and ( n25619 , n25615 , n25618 );
and ( n25620 , n25611 , n25618 );
or ( n25621 , n25616 , n25619 , n25620 );
xor ( n25622 , n25290 , n25294 );
xor ( n25623 , n25622 , n25297 );
and ( n25624 , n25621 , n25623 );
xor ( n25625 , n25451 , n25519 );
xor ( n25626 , n25625 , n25522 );
and ( n25627 , n25624 , n25626 );
and ( n25628 , n21252 , n22032 );
and ( n25629 , n21265 , n22029 );
nor ( n25630 , n25628 , n25629 );
xnor ( n25631 , n25630 , n22027 );
xor ( n25632 , n25371 , n25375 );
xor ( n25633 , n25632 , n25378 );
and ( n25634 , n25631 , n25633 );
and ( n25635 , n25060 , n21496 );
and ( n25636 , n24812 , n21494 );
nor ( n25637 , n25635 , n25636 );
xnor ( n25638 , n25637 , n21506 );
and ( n25639 , n25343 , n21551 );
and ( n25640 , n25179 , n21549 );
nor ( n25641 , n25639 , n25640 );
xnor ( n25642 , n25641 , n21557 );
and ( n25643 , n25638 , n25642 );
and ( n25644 , n25544 , n21513 );
and ( n25645 , n25642 , n25644 );
and ( n25646 , n25638 , n25644 );
or ( n25647 , n25643 , n25645 , n25646 );
and ( n25648 , n24213 , n21529 );
and ( n25649 , n23949 , n21527 );
nor ( n25650 , n25648 , n25649 );
xnor ( n25651 , n25650 , n21539 );
and ( n25652 , n25647 , n25651 );
and ( n25653 , n24812 , n21496 );
and ( n25654 , n24662 , n21494 );
nor ( n25655 , n25653 , n25654 );
xnor ( n25656 , n25655 , n21506 );
and ( n25657 , n25651 , n25656 );
and ( n25658 , n25647 , n25656 );
or ( n25659 , n25652 , n25657 , n25658 );
and ( n25660 , n21511 , n21236 );
and ( n25661 , n21599 , n21234 );
nor ( n25662 , n25660 , n25661 );
xnor ( n25663 , n25662 , n21246 );
and ( n25664 , n25659 , n25663 );
and ( n25665 , n23074 , n21582 );
and ( n25666 , n22813 , n21580 );
nor ( n25667 , n25665 , n25666 );
xnor ( n25668 , n25667 , n21588 );
and ( n25669 , n25663 , n25668 );
and ( n25670 , n25659 , n25668 );
or ( n25671 , n25664 , n25669 , n25670 );
and ( n25672 , n21756 , n21663 );
and ( n25673 , n21519 , n21661 );
nor ( n25674 , n25672 , n25673 );
xnor ( n25675 , n25674 , n21673 );
and ( n25676 , n25671 , n25675 );
xor ( n25677 , n25359 , n25363 );
xor ( n25678 , n25677 , n25368 );
and ( n25679 , n25675 , n25678 );
and ( n25680 , n25671 , n25678 );
or ( n25681 , n25676 , n25679 , n25680 );
and ( n25682 , n25633 , n25681 );
and ( n25683 , n25631 , n25681 );
or ( n25684 , n25634 , n25682 , n25683 );
xor ( n25685 , n25421 , n25423 );
xor ( n25686 , n25685 , n25438 );
and ( n25687 , n25684 , n25686 );
xor ( n25688 , n25455 , n25457 );
xor ( n25689 , n25688 , n25510 );
and ( n25690 , n25686 , n25689 );
and ( n25691 , n25684 , n25689 );
or ( n25692 , n25687 , n25690 , n25691 );
xor ( n25693 , n25453 , n25513 );
xor ( n25694 , n25693 , n25516 );
and ( n25695 , n25692 , n25694 );
xor ( n25696 , n25621 , n25623 );
and ( n25697 , n25694 , n25696 );
and ( n25698 , n25692 , n25696 );
or ( n25699 , n25695 , n25697 , n25698 );
and ( n25700 , n25626 , n25699 );
and ( n25701 , n25624 , n25699 );
or ( n25702 , n25627 , n25700 , n25701 );
and ( n25703 , n25535 , n25702 );
and ( n25704 , n25533 , n25702 );
or ( n25705 , n25536 , n25703 , n25704 );
and ( n25706 , n25530 , n25705 );
and ( n25707 , n25528 , n25705 );
or ( n25708 , n25531 , n25706 , n25707 );
and ( n25709 , n25327 , n25708 );
and ( n25710 , n25325 , n25708 );
or ( n25711 , n25328 , n25709 , n25710 );
and ( n25712 , n25254 , n25711 );
xor ( n25713 , n25254 , n25711 );
xor ( n25714 , n25325 , n25327 );
xor ( n25715 , n25714 , n25708 );
xor ( n25716 , n25528 , n25530 );
xor ( n25717 , n25716 , n25705 );
xor ( n25718 , n25533 , n25535 );
xor ( n25719 , n25718 , n25702 );
xor ( n25720 , n25624 , n25626 );
xor ( n25721 , n25720 , n25699 );
xor ( n25722 , n25611 , n25615 );
xor ( n25723 , n25722 , n25618 );
and ( n25724 , n23320 , n21582 );
and ( n25725 , n23074 , n21580 );
nor ( n25726 , n25724 , n25725 );
xnor ( n25727 , n25726 , n21588 );
and ( n25728 , n23503 , n21783 );
and ( n25729 , n23351 , n21781 );
nor ( n25730 , n25728 , n25729 );
xnor ( n25731 , n25730 , n21793 );
and ( n25732 , n25727 , n25731 );
xor ( n25733 , n25647 , n25651 );
xor ( n25734 , n25733 , n25656 );
and ( n25735 , n25731 , n25734 );
and ( n25736 , n25727 , n25734 );
or ( n25737 , n25732 , n25735 , n25736 );
and ( n25738 , n21501 , n21687 );
and ( n25739 , n21630 , n21685 );
nor ( n25740 , n25738 , n25739 );
xnor ( n25741 , n25740 , n21697 );
and ( n25742 , n25737 , n25741 );
xor ( n25743 , n25471 , n25475 );
xor ( n25744 , n25743 , n25478 );
and ( n25745 , n25741 , n25744 );
and ( n25746 , n25737 , n25744 );
or ( n25747 , n25742 , n25745 , n25746 );
and ( n25748 , n21777 , n22114 );
and ( n25749 , n21788 , n22112 );
nor ( n25750 , n25748 , n25749 );
xnor ( n25751 , n25750 , n22124 );
and ( n25752 , n25747 , n25751 );
and ( n25753 , n21744 , n21414 );
and ( n25754 , n22089 , n21412 );
nor ( n25755 , n25753 , n25754 );
xnor ( n25756 , n25755 , n21480 );
and ( n25757 , n25751 , n25756 );
and ( n25758 , n25747 , n25756 );
or ( n25759 , n25752 , n25757 , n25758 );
and ( n25760 , n25343 , n21496 );
and ( n25761 , n25179 , n21494 );
nor ( n25762 , n25760 , n25761 );
xnor ( n25763 , n25762 , n21506 );
and ( n25764 , n25553 , n21551 );
and ( n25765 , n25544 , n21549 );
nor ( n25766 , n25764 , n25765 );
xnor ( n25767 , n25766 , n21557 );
and ( n25768 , n25763 , n25767 );
xor ( n25769 , n21038 , n21063 );
buf ( n25770 , n25769 );
buf ( n25771 , n25770 );
buf ( n25772 , n25771 );
and ( n25773 , n25772 , n21513 );
and ( n25774 , n25767 , n25773 );
and ( n25775 , n25763 , n25773 );
or ( n25776 , n25768 , n25774 , n25775 );
and ( n25777 , n24631 , n21529 );
and ( n25778 , n24460 , n21527 );
nor ( n25779 , n25777 , n25778 );
xnor ( n25780 , n25779 , n21539 );
and ( n25781 , n25776 , n25780 );
xor ( n25782 , n25540 , n25548 );
xor ( n25783 , n25782 , n25554 );
and ( n25784 , n25780 , n25783 );
and ( n25785 , n25776 , n25783 );
or ( n25786 , n25781 , n25784 , n25785 );
and ( n25787 , n23949 , n21739 );
and ( n25788 , n23887 , n21737 );
nor ( n25789 , n25787 , n25788 );
xnor ( n25790 , n25789 , n21749 );
and ( n25791 , n25786 , n25790 );
xor ( n25792 , n25638 , n25642 );
xor ( n25793 , n25792 , n25644 );
and ( n25794 , n25790 , n25793 );
and ( n25795 , n25786 , n25793 );
or ( n25796 , n25791 , n25794 , n25795 );
and ( n25797 , n21606 , n21236 );
and ( n25798 , n21511 , n21234 );
nor ( n25799 , n25797 , n25798 );
xnor ( n25800 , n25799 , n21246 );
and ( n25801 , n25796 , n25800 );
and ( n25802 , n22813 , n21260 );
and ( n25803 , n21616 , n21258 );
nor ( n25804 , n25802 , n25803 );
xnor ( n25805 , n25804 , n21270 );
and ( n25806 , n25800 , n25805 );
and ( n25807 , n25796 , n25805 );
or ( n25808 , n25801 , n25806 , n25807 );
and ( n25809 , n21545 , n21707 );
and ( n25810 , n21486 , n21705 );
nor ( n25811 , n25809 , n25810 );
xnor ( n25812 , n25811 , n21717 );
and ( n25813 , n25808 , n25812 );
xor ( n25814 , n25659 , n25663 );
xor ( n25815 , n25814 , n25668 );
and ( n25816 , n25812 , n25815 );
and ( n25817 , n25808 , n25815 );
or ( n25818 , n25813 , n25816 , n25817 );
and ( n25819 , n21574 , n22032 );
and ( n25820 , n21252 , n22029 );
nor ( n25821 , n25819 , n25820 );
xnor ( n25822 , n25821 , n22027 );
and ( n25823 , n25818 , n25822 );
xor ( n25824 , n25589 , n25593 );
xor ( n25825 , n25824 , n25596 );
and ( n25826 , n25822 , n25825 );
and ( n25827 , n25818 , n25825 );
or ( n25828 , n25823 , n25826 , n25827 );
and ( n25829 , n25759 , n25828 );
xor ( n25830 , n25599 , n25603 );
xor ( n25831 , n25830 , n25608 );
and ( n25832 , n25828 , n25831 );
and ( n25833 , n25759 , n25831 );
or ( n25834 , n25829 , n25832 , n25833 );
and ( n25835 , n25723 , n25834 );
xor ( n25836 , n25492 , n25494 );
xor ( n25837 , n25836 , n25507 );
xor ( n25838 , n25631 , n25633 );
xor ( n25839 , n25838 , n25681 );
and ( n25840 , n25837 , n25839 );
and ( n25841 , n21519 , n21139 );
and ( n25842 , n21534 , n21137 );
nor ( n25843 , n25841 , n25842 );
xnor ( n25844 , n25843 , n21221 );
and ( n25845 , n21645 , n21663 );
and ( n25846 , n21756 , n21661 );
nor ( n25847 , n25845 , n25846 );
xnor ( n25848 , n25847 , n21673 );
and ( n25849 , n25844 , n25848 );
xor ( n25850 , n25579 , n25583 );
xor ( n25851 , n25850 , n25586 );
and ( n25852 , n25848 , n25851 );
and ( n25853 , n25844 , n25851 );
or ( n25854 , n25849 , n25852 , n25853 );
xor ( n25855 , n25671 , n25675 );
xor ( n25856 , n25855 , n25678 );
and ( n25857 , n25854 , n25856 );
xor ( n25858 , n25462 , n25466 );
xor ( n25859 , n25858 , n25489 );
and ( n25860 , n25856 , n25859 );
and ( n25861 , n25854 , n25859 );
or ( n25862 , n25857 , n25860 , n25861 );
and ( n25863 , n25839 , n25862 );
and ( n25864 , n25837 , n25862 );
or ( n25865 , n25840 , n25863 , n25864 );
and ( n25866 , n25834 , n25865 );
and ( n25867 , n25723 , n25865 );
or ( n25868 , n25835 , n25866 , n25867 );
xor ( n25869 , n25692 , n25694 );
xor ( n25870 , n25869 , n25696 );
and ( n25871 , n25868 , n25870 );
xor ( n25872 , n25684 , n25686 );
xor ( n25873 , n25872 , n25689 );
xor ( n25874 , n25723 , n25834 );
xor ( n25875 , n25874 , n25865 );
and ( n25876 , n25873 , n25875 );
and ( n25877 , n23320 , n21260 );
and ( n25878 , n23074 , n21258 );
nor ( n25879 , n25877 , n25878 );
xnor ( n25880 , n25879 , n21270 );
and ( n25881 , n23503 , n21582 );
and ( n25882 , n23351 , n21580 );
nor ( n25883 , n25881 , n25882 );
xnor ( n25884 , n25883 , n21588 );
and ( n25885 , n25880 , n25884 );
and ( n25886 , n25544 , n21496 );
and ( n25887 , n25343 , n21494 );
nor ( n25888 , n25886 , n25887 );
xnor ( n25889 , n25888 , n21506 );
and ( n25890 , n25772 , n21551 );
and ( n25891 , n25553 , n21549 );
nor ( n25892 , n25890 , n25891 );
xnor ( n25893 , n25892 , n21557 );
and ( n25894 , n25889 , n25893 );
xor ( n25895 , n21045 , n21061 );
buf ( n25896 , n25895 );
buf ( n25897 , n25896 );
buf ( n25898 , n25897 );
and ( n25899 , n25898 , n21513 );
and ( n25900 , n25893 , n25899 );
and ( n25901 , n25889 , n25899 );
or ( n25902 , n25894 , n25900 , n25901 );
and ( n25903 , n25060 , n21625 );
and ( n25904 , n24812 , n21623 );
nor ( n25905 , n25903 , n25904 );
xnor ( n25906 , n25905 , n21635 );
and ( n25907 , n25902 , n25906 );
xor ( n25908 , n25763 , n25767 );
xor ( n25909 , n25908 , n25773 );
and ( n25910 , n25906 , n25909 );
and ( n25911 , n25902 , n25909 );
or ( n25912 , n25907 , n25910 , n25911 );
and ( n25913 , n24213 , n21739 );
and ( n25914 , n23949 , n21737 );
nor ( n25915 , n25913 , n25914 );
xnor ( n25916 , n25915 , n21749 );
xor ( n25917 , n25912 , n25916 );
and ( n25918 , n24812 , n21625 );
and ( n25919 , n24662 , n21623 );
nor ( n25920 , n25918 , n25919 );
xnor ( n25921 , n25920 , n21635 );
xor ( n25922 , n25917 , n25921 );
and ( n25923 , n25884 , n25922 );
and ( n25924 , n25880 , n25922 );
or ( n25925 , n25885 , n25923 , n25924 );
and ( n25926 , n21501 , n21663 );
and ( n25927 , n21630 , n21661 );
nor ( n25928 , n25926 , n25927 );
xnor ( n25929 , n25928 , n21673 );
and ( n25930 , n25925 , n25929 );
and ( n25931 , n23074 , n21260 );
and ( n25932 , n22813 , n21258 );
nor ( n25933 , n25931 , n25932 );
xnor ( n25934 , n25933 , n21270 );
and ( n25935 , n23351 , n21582 );
and ( n25936 , n23320 , n21580 );
nor ( n25937 , n25935 , n25936 );
xnor ( n25938 , n25937 , n21588 );
xor ( n25939 , n25934 , n25938 );
and ( n25940 , n23651 , n21783 );
and ( n25941 , n23503 , n21781 );
nor ( n25942 , n25940 , n25941 );
xnor ( n25943 , n25942 , n21793 );
xor ( n25944 , n25939 , n25943 );
and ( n25945 , n25929 , n25944 );
and ( n25946 , n25925 , n25944 );
or ( n25947 , n25930 , n25945 , n25946 );
and ( n25948 , n21534 , n21414 );
and ( n25949 , n21731 , n21412 );
nor ( n25950 , n25948 , n25949 );
xnor ( n25951 , n25950 , n21480 );
and ( n25952 , n25947 , n25951 );
xor ( n25953 , n25796 , n25800 );
xor ( n25954 , n25953 , n25805 );
and ( n25955 , n25951 , n25954 );
and ( n25956 , n25947 , n25954 );
or ( n25957 , n25952 , n25955 , n25956 );
and ( n25958 , n21777 , n22032 );
and ( n25959 , n21788 , n22029 );
nor ( n25960 , n25958 , n25959 );
xnor ( n25961 , n25960 , n22027 );
and ( n25962 , n21744 , n22114 );
and ( n25963 , n22089 , n22112 );
nor ( n25964 , n25962 , n25963 );
xnor ( n25965 , n25964 , n22124 );
and ( n25966 , n25961 , n25965 );
and ( n25967 , n25934 , n25938 );
and ( n25968 , n25938 , n25943 );
and ( n25969 , n25934 , n25943 );
or ( n25970 , n25967 , n25968 , n25969 );
and ( n25971 , n21486 , n21687 );
and ( n25972 , n21501 , n21685 );
nor ( n25973 , n25971 , n25972 );
xnor ( n25974 , n25973 , n21697 );
xor ( n25975 , n25970 , n25974 );
xor ( n25976 , n25569 , n25573 );
xor ( n25977 , n25976 , n25576 );
xor ( n25978 , n25975 , n25977 );
and ( n25979 , n25965 , n25978 );
and ( n25980 , n25961 , n25978 );
or ( n25981 , n25966 , n25979 , n25980 );
and ( n25982 , n25957 , n25981 );
and ( n25983 , n25970 , n25974 );
and ( n25984 , n25974 , n25977 );
and ( n25985 , n25970 , n25977 );
or ( n25986 , n25983 , n25984 , n25985 );
and ( n25987 , n22089 , n22114 );
and ( n25988 , n21777 , n22112 );
nor ( n25989 , n25987 , n25988 );
xnor ( n25990 , n25989 , n22124 );
xor ( n25991 , n25986 , n25990 );
and ( n25992 , n21731 , n21414 );
and ( n25993 , n21744 , n21412 );
nor ( n25994 , n25992 , n25993 );
xnor ( n25995 , n25994 , n21480 );
xor ( n25996 , n25991 , n25995 );
and ( n25997 , n25981 , n25996 );
and ( n25998 , n25957 , n25996 );
or ( n25999 , n25982 , n25997 , n25998 );
buf ( n26000 , n21056 );
buf ( n26001 , n26000 );
buf ( n26002 , n26001 );
buf ( n26003 , n26002 );
and ( n26004 , n26003 , n21549 );
not ( n26005 , n26004 );
and ( n26006 , n26005 , n21557 );
and ( n26007 , n26003 , n21551 );
xor ( n26008 , n21055 , n21058 );
buf ( n26009 , n26008 );
buf ( n26010 , n26009 );
buf ( n26011 , n26010 );
and ( n26012 , n26011 , n21549 );
nor ( n26013 , n26007 , n26012 );
xnor ( n26014 , n26013 , n21557 );
and ( n26015 , n26006 , n26014 );
and ( n26016 , n26011 , n21551 );
xor ( n26017 , n21051 , n21059 );
buf ( n26018 , n26017 );
buf ( n26019 , n26018 );
buf ( n26020 , n26019 );
and ( n26021 , n26020 , n21549 );
nor ( n26022 , n26016 , n26021 );
xnor ( n26023 , n26022 , n21557 );
and ( n26024 , n26015 , n26023 );
and ( n26025 , n26003 , n21513 );
and ( n26026 , n26023 , n26025 );
and ( n26027 , n26015 , n26025 );
or ( n26028 , n26024 , n26026 , n26027 );
and ( n26029 , n26020 , n21551 );
and ( n26030 , n25898 , n21549 );
nor ( n26031 , n26029 , n26030 );
xnor ( n26032 , n26031 , n21557 );
and ( n26033 , n26028 , n26032 );
and ( n26034 , n26011 , n21513 );
and ( n26035 , n26032 , n26034 );
and ( n26036 , n26028 , n26034 );
or ( n26037 , n26033 , n26035 , n26036 );
and ( n26038 , n25898 , n21551 );
and ( n26039 , n25772 , n21549 );
nor ( n26040 , n26038 , n26039 );
xnor ( n26041 , n26040 , n21557 );
and ( n26042 , n26037 , n26041 );
and ( n26043 , n26020 , n21513 );
and ( n26044 , n26041 , n26043 );
and ( n26045 , n26037 , n26043 );
or ( n26046 , n26042 , n26044 , n26045 );
and ( n26047 , n25179 , n21625 );
and ( n26048 , n25060 , n21623 );
nor ( n26049 , n26047 , n26048 );
xnor ( n26050 , n26049 , n21635 );
and ( n26051 , n26046 , n26050 );
xor ( n26052 , n25889 , n25893 );
xor ( n26053 , n26052 , n25899 );
and ( n26054 , n26050 , n26053 );
and ( n26055 , n26046 , n26053 );
or ( n26056 , n26051 , n26054 , n26055 );
and ( n26057 , n24460 , n21739 );
and ( n26058 , n24213 , n21737 );
nor ( n26059 , n26057 , n26058 );
xnor ( n26060 , n26059 , n21749 );
and ( n26061 , n26056 , n26060 );
and ( n26062 , n24662 , n21529 );
and ( n26063 , n24631 , n21527 );
nor ( n26064 , n26062 , n26063 );
xnor ( n26065 , n26064 , n21539 );
and ( n26066 , n26060 , n26065 );
and ( n26067 , n26056 , n26065 );
or ( n26068 , n26061 , n26066 , n26067 );
and ( n26069 , n23887 , n21783 );
and ( n26070 , n23651 , n21781 );
nor ( n26071 , n26069 , n26070 );
xnor ( n26072 , n26071 , n21793 );
and ( n26073 , n26068 , n26072 );
xor ( n26074 , n25776 , n25780 );
xor ( n26075 , n26074 , n25783 );
and ( n26076 , n26072 , n26075 );
and ( n26077 , n26068 , n26075 );
or ( n26078 , n26073 , n26076 , n26077 );
and ( n26079 , n21511 , n21707 );
and ( n26080 , n21599 , n21705 );
nor ( n26081 , n26079 , n26080 );
xnor ( n26082 , n26081 , n21717 );
and ( n26083 , n26078 , n26082 );
xor ( n26084 , n25786 , n25790 );
xor ( n26085 , n26084 , n25793 );
and ( n26086 , n26082 , n26085 );
and ( n26087 , n26078 , n26085 );
or ( n26088 , n26083 , n26086 , n26087 );
and ( n26089 , n21756 , n21139 );
and ( n26090 , n21519 , n21137 );
nor ( n26091 , n26089 , n26090 );
xnor ( n26092 , n26091 , n21221 );
and ( n26093 , n26088 , n26092 );
and ( n26094 , n21630 , n21663 );
and ( n26095 , n21645 , n21661 );
nor ( n26096 , n26094 , n26095 );
xnor ( n26097 , n26096 , n21673 );
and ( n26098 , n26092 , n26097 );
and ( n26099 , n26088 , n26097 );
or ( n26100 , n26093 , n26098 , n26099 );
xor ( n26101 , n25808 , n25812 );
xor ( n26102 , n26101 , n25815 );
and ( n26103 , n26100 , n26102 );
xor ( n26104 , n25844 , n25848 );
xor ( n26105 , n26104 , n25851 );
and ( n26106 , n26102 , n26105 );
and ( n26107 , n26100 , n26105 );
or ( n26108 , n26103 , n26106 , n26107 );
and ( n26109 , n25999 , n26108 );
xor ( n26110 , n25747 , n25751 );
xor ( n26111 , n26110 , n25756 );
and ( n26112 , n26108 , n26111 );
and ( n26113 , n25999 , n26111 );
or ( n26114 , n26109 , n26112 , n26113 );
and ( n26115 , n25986 , n25990 );
and ( n26116 , n25990 , n25995 );
and ( n26117 , n25986 , n25995 );
or ( n26118 , n26115 , n26116 , n26117 );
and ( n26119 , n25912 , n25916 );
and ( n26120 , n25916 , n25921 );
and ( n26121 , n25912 , n25921 );
or ( n26122 , n26119 , n26120 , n26121 );
and ( n26123 , n21616 , n21236 );
and ( n26124 , n21606 , n21234 );
nor ( n26125 , n26123 , n26124 );
xnor ( n26126 , n26125 , n21246 );
and ( n26127 , n26122 , n26126 );
xor ( n26128 , n25557 , n25561 );
xor ( n26129 , n26128 , n25566 );
and ( n26130 , n26126 , n26129 );
and ( n26131 , n26122 , n26129 );
or ( n26132 , n26127 , n26130 , n26131 );
and ( n26133 , n21599 , n21707 );
and ( n26134 , n21545 , n21705 );
nor ( n26135 , n26133 , n26134 );
xnor ( n26136 , n26135 , n21717 );
and ( n26137 , n26132 , n26136 );
xor ( n26138 , n25727 , n25731 );
xor ( n26139 , n26138 , n25734 );
and ( n26140 , n26136 , n26139 );
and ( n26141 , n26132 , n26139 );
or ( n26142 , n26137 , n26140 , n26141 );
and ( n26143 , n21788 , n22032 );
and ( n26144 , n21574 , n22029 );
nor ( n26145 , n26143 , n26144 );
xnor ( n26146 , n26145 , n22027 );
and ( n26147 , n26142 , n26146 );
xor ( n26148 , n25737 , n25741 );
xor ( n26149 , n26148 , n25744 );
and ( n26150 , n26146 , n26149 );
and ( n26151 , n26142 , n26149 );
or ( n26152 , n26147 , n26150 , n26151 );
and ( n26153 , n26118 , n26152 );
xor ( n26154 , n25818 , n25822 );
xor ( n26155 , n26154 , n25825 );
and ( n26156 , n26152 , n26155 );
and ( n26157 , n26118 , n26155 );
or ( n26158 , n26153 , n26156 , n26157 );
and ( n26159 , n26114 , n26158 );
xor ( n26160 , n25759 , n25828 );
xor ( n26161 , n26160 , n25831 );
and ( n26162 , n26158 , n26161 );
and ( n26163 , n26114 , n26161 );
or ( n26164 , n26159 , n26162 , n26163 );
and ( n26165 , n25875 , n26164 );
and ( n26166 , n25873 , n26164 );
or ( n26167 , n25876 , n26165 , n26166 );
and ( n26168 , n25870 , n26167 );
and ( n26169 , n25868 , n26167 );
or ( n26170 , n25871 , n26168 , n26169 );
and ( n26171 , n25721 , n26170 );
xor ( n26172 , n25721 , n26170 );
xor ( n26173 , n25868 , n25870 );
xor ( n26174 , n26173 , n26167 );
xor ( n26175 , n25837 , n25839 );
xor ( n26176 , n26175 , n25862 );
xor ( n26177 , n26114 , n26158 );
xor ( n26178 , n26177 , n26161 );
and ( n26179 , n26176 , n26178 );
and ( n26180 , n23651 , n21582 );
and ( n26181 , n23503 , n21580 );
nor ( n26182 , n26180 , n26181 );
xnor ( n26183 , n26182 , n21588 );
and ( n26184 , n23949 , n21783 );
and ( n26185 , n23887 , n21781 );
nor ( n26186 , n26184 , n26185 );
xnor ( n26187 , n26186 , n21793 );
and ( n26188 , n26183 , n26187 );
xor ( n26189 , n25902 , n25906 );
xor ( n26190 , n26189 , n25909 );
and ( n26191 , n26187 , n26190 );
and ( n26192 , n26183 , n26190 );
or ( n26193 , n26188 , n26191 , n26192 );
and ( n26194 , n21606 , n21707 );
and ( n26195 , n21511 , n21705 );
nor ( n26196 , n26194 , n26195 );
xnor ( n26197 , n26196 , n21717 );
and ( n26198 , n26193 , n26197 );
and ( n26199 , n22813 , n21236 );
and ( n26200 , n21616 , n21234 );
nor ( n26201 , n26199 , n26200 );
xnor ( n26202 , n26201 , n21246 );
and ( n26203 , n26197 , n26202 );
and ( n26204 , n26193 , n26202 );
or ( n26205 , n26198 , n26203 , n26204 );
and ( n26206 , n21519 , n21414 );
and ( n26207 , n21534 , n21412 );
nor ( n26208 , n26206 , n26207 );
xnor ( n26209 , n26208 , n21480 );
and ( n26210 , n26205 , n26209 );
and ( n26211 , n21545 , n21687 );
and ( n26212 , n21486 , n21685 );
nor ( n26213 , n26211 , n26212 );
xnor ( n26214 , n26213 , n21697 );
and ( n26215 , n26209 , n26214 );
and ( n26216 , n26205 , n26214 );
or ( n26217 , n26210 , n26215 , n26216 );
xor ( n26218 , n26088 , n26092 );
xor ( n26219 , n26218 , n26097 );
and ( n26220 , n26217 , n26219 );
xor ( n26221 , n26132 , n26136 );
xor ( n26222 , n26221 , n26139 );
and ( n26223 , n26219 , n26222 );
and ( n26224 , n26217 , n26222 );
or ( n26225 , n26220 , n26223 , n26224 );
xor ( n26226 , n26142 , n26146 );
xor ( n26227 , n26226 , n26149 );
and ( n26228 , n26225 , n26227 );
xor ( n26229 , n26100 , n26102 );
xor ( n26230 , n26229 , n26105 );
and ( n26231 , n26227 , n26230 );
and ( n26232 , n26225 , n26230 );
or ( n26233 , n26228 , n26231 , n26232 );
xor ( n26234 , n25854 , n25856 );
xor ( n26235 , n26234 , n25859 );
and ( n26236 , n26233 , n26235 );
xor ( n26237 , n26118 , n26152 );
xor ( n26238 , n26237 , n26155 );
and ( n26239 , n26235 , n26238 );
and ( n26240 , n26233 , n26238 );
or ( n26241 , n26236 , n26239 , n26240 );
and ( n26242 , n26178 , n26241 );
and ( n26243 , n26176 , n26241 );
or ( n26244 , n26179 , n26242 , n26243 );
xor ( n26245 , n25873 , n25875 );
xor ( n26246 , n26245 , n26164 );
and ( n26247 , n26244 , n26246 );
xor ( n26248 , n25999 , n26108 );
xor ( n26249 , n26248 , n26111 );
xor ( n26250 , n25957 , n25981 );
xor ( n26251 , n26250 , n25996 );
and ( n26252 , n21731 , n22114 );
and ( n26253 , n21744 , n22112 );
nor ( n26254 , n26252 , n26253 );
xnor ( n26255 , n26254 , n22124 );
and ( n26256 , n21744 , n22032 );
and ( n26257 , n22089 , n22029 );
nor ( n26258 , n26256 , n26257 );
xnor ( n26259 , n26258 , n22027 );
and ( n26260 , n21534 , n22114 );
and ( n26261 , n21731 , n22112 );
nor ( n26262 , n26260 , n26261 );
xnor ( n26263 , n26262 , n22124 );
and ( n26264 , n26259 , n26263 );
and ( n26265 , n21731 , n22032 );
and ( n26266 , n21744 , n22029 );
nor ( n26267 , n26265 , n26266 );
xnor ( n26268 , n26267 , n22027 );
and ( n26269 , n21645 , n21414 );
and ( n26270 , n21756 , n21412 );
nor ( n26271 , n26269 , n26270 );
xnor ( n26272 , n26271 , n21480 );
and ( n26273 , n26268 , n26272 );
and ( n26274 , n21545 , n21663 );
and ( n26275 , n21486 , n21661 );
nor ( n26276 , n26274 , n26275 );
xnor ( n26277 , n26276 , n21673 );
and ( n26278 , n26272 , n26277 );
and ( n26279 , n26268 , n26277 );
or ( n26280 , n26273 , n26278 , n26279 );
and ( n26281 , n26263 , n26280 );
and ( n26282 , n26259 , n26280 );
or ( n26283 , n26264 , n26281 , n26282 );
and ( n26284 , n26255 , n26283 );
and ( n26285 , n23074 , n21236 );
and ( n26286 , n22813 , n21234 );
nor ( n26287 , n26285 , n26286 );
xnor ( n26288 , n26287 , n21246 );
and ( n26289 , n23351 , n21260 );
and ( n26290 , n23320 , n21258 );
nor ( n26291 , n26289 , n26290 );
xnor ( n26292 , n26291 , n21270 );
and ( n26293 , n26288 , n26292 );
and ( n26294 , n21534 , n22032 );
and ( n26295 , n21731 , n22029 );
nor ( n26296 , n26294 , n26295 );
xnor ( n26297 , n26296 , n22027 );
and ( n26298 , n21630 , n21414 );
and ( n26299 , n21645 , n21412 );
nor ( n26300 , n26298 , n26299 );
xnor ( n26301 , n26300 , n21480 );
and ( n26302 , n26297 , n26301 );
and ( n26303 , n26292 , n26302 );
and ( n26304 , n26288 , n26302 );
or ( n26305 , n26293 , n26303 , n26304 );
and ( n26306 , n21756 , n22114 );
and ( n26307 , n21519 , n22112 );
nor ( n26308 , n26306 , n26307 );
xnor ( n26309 , n26308 , n22124 );
and ( n26310 , n21486 , n21139 );
and ( n26311 , n21501 , n21137 );
nor ( n26312 , n26310 , n26311 );
xnor ( n26313 , n26312 , n21221 );
and ( n26314 , n26309 , n26313 );
and ( n26315 , n21599 , n21663 );
and ( n26316 , n21545 , n21661 );
nor ( n26317 , n26315 , n26316 );
xnor ( n26318 , n26317 , n21673 );
and ( n26319 , n26313 , n26318 );
and ( n26320 , n26309 , n26318 );
or ( n26321 , n26314 , n26319 , n26320 );
and ( n26322 , n23320 , n21236 );
and ( n26323 , n23074 , n21234 );
nor ( n26324 , n26322 , n26323 );
xnor ( n26325 , n26324 , n21246 );
and ( n26326 , n23503 , n21260 );
and ( n26327 , n23351 , n21258 );
nor ( n26328 , n26326 , n26327 );
xnor ( n26329 , n26328 , n21270 );
and ( n26330 , n26325 , n26329 );
and ( n26331 , n23887 , n21582 );
and ( n26332 , n23651 , n21580 );
nor ( n26333 , n26331 , n26332 );
xnor ( n26334 , n26333 , n21588 );
and ( n26335 , n26329 , n26334 );
and ( n26336 , n26325 , n26334 );
or ( n26337 , n26330 , n26335 , n26336 );
and ( n26338 , n26321 , n26337 );
xor ( n26339 , n26268 , n26272 );
xor ( n26340 , n26339 , n26277 );
and ( n26341 , n26337 , n26340 );
and ( n26342 , n26321 , n26340 );
or ( n26343 , n26338 , n26341 , n26342 );
and ( n26344 , n26305 , n26343 );
xor ( n26345 , n26259 , n26263 );
xor ( n26346 , n26345 , n26280 );
and ( n26347 , n26343 , n26346 );
and ( n26348 , n26305 , n26346 );
or ( n26349 , n26344 , n26347 , n26348 );
and ( n26350 , n26283 , n26349 );
and ( n26351 , n26255 , n26349 );
or ( n26352 , n26284 , n26350 , n26351 );
xor ( n26353 , n26255 , n26283 );
xor ( n26354 , n26353 , n26349 );
xor ( n26355 , n25925 , n25929 );
xor ( n26356 , n26355 , n25944 );
and ( n26357 , n26354 , n26356 );
xor ( n26358 , n26297 , n26301 );
and ( n26359 , n21511 , n21663 );
and ( n26360 , n21599 , n21661 );
nor ( n26361 , n26359 , n26360 );
xnor ( n26362 , n26361 , n21673 );
and ( n26363 , n21616 , n21687 );
and ( n26364 , n21606 , n21685 );
nor ( n26365 , n26363 , n26364 );
xnor ( n26366 , n26365 , n21697 );
and ( n26367 , n26362 , n26366 );
and ( n26368 , n26358 , n26367 );
and ( n26369 , n21519 , n22032 );
and ( n26370 , n21534 , n22029 );
nor ( n26371 , n26369 , n26370 );
xnor ( n26372 , n26371 , n22027 );
and ( n26373 , n21645 , n22114 );
and ( n26374 , n21756 , n22112 );
nor ( n26375 , n26373 , n26374 );
xnor ( n26376 , n26375 , n22124 );
and ( n26377 , n26372 , n26376 );
and ( n26378 , n21501 , n21414 );
and ( n26379 , n21630 , n21412 );
nor ( n26380 , n26378 , n26379 );
xnor ( n26381 , n26380 , n21480 );
and ( n26382 , n26376 , n26381 );
and ( n26383 , n26372 , n26381 );
or ( n26384 , n26377 , n26382 , n26383 );
and ( n26385 , n26367 , n26384 );
and ( n26386 , n26358 , n26384 );
or ( n26387 , n26368 , n26385 , n26386 );
and ( n26388 , n21545 , n21139 );
and ( n26389 , n21486 , n21137 );
nor ( n26390 , n26388 , n26389 );
xnor ( n26391 , n26390 , n21221 );
and ( n26392 , n23074 , n21707 );
and ( n26393 , n22813 , n21705 );
nor ( n26394 , n26392 , n26393 );
xnor ( n26395 , n26394 , n21717 );
and ( n26396 , n26391 , n26395 );
and ( n26397 , n23351 , n21236 );
and ( n26398 , n23320 , n21234 );
nor ( n26399 , n26397 , n26398 );
xnor ( n26400 , n26399 , n21246 );
and ( n26401 , n26395 , n26400 );
and ( n26402 , n26391 , n26400 );
or ( n26403 , n26396 , n26401 , n26402 );
xor ( n26404 , n26309 , n26313 );
xor ( n26405 , n26404 , n26318 );
and ( n26406 , n26403 , n26405 );
xor ( n26407 , n26325 , n26329 );
xor ( n26408 , n26407 , n26334 );
and ( n26409 , n26405 , n26408 );
and ( n26410 , n26403 , n26408 );
or ( n26411 , n26406 , n26409 , n26410 );
and ( n26412 , n26387 , n26411 );
xor ( n26413 , n26288 , n26292 );
xor ( n26414 , n26413 , n26302 );
and ( n26415 , n26411 , n26414 );
and ( n26416 , n26387 , n26414 );
or ( n26417 , n26412 , n26415 , n26416 );
xor ( n26418 , n26305 , n26343 );
xor ( n26419 , n26418 , n26346 );
and ( n26420 , n26417 , n26419 );
xor ( n26421 , n25880 , n25884 );
xor ( n26422 , n26421 , n25922 );
and ( n26423 , n26419 , n26422 );
and ( n26424 , n26417 , n26422 );
or ( n26425 , n26420 , n26423 , n26424 );
and ( n26426 , n26356 , n26425 );
and ( n26427 , n26354 , n26425 );
or ( n26428 , n26357 , n26426 , n26427 );
and ( n26429 , n26352 , n26428 );
and ( n26430 , n21616 , n21707 );
and ( n26431 , n21606 , n21705 );
nor ( n26432 , n26430 , n26431 );
xnor ( n26433 , n26432 , n21717 );
xor ( n26434 , n26183 , n26187 );
xor ( n26435 , n26434 , n26190 );
and ( n26436 , n26433 , n26435 );
xor ( n26437 , n26321 , n26337 );
xor ( n26438 , n26437 , n26340 );
and ( n26439 , n24460 , n21783 );
and ( n26440 , n24213 , n21781 );
nor ( n26441 , n26439 , n26440 );
xnor ( n26442 , n26441 , n21793 );
and ( n26443 , n24662 , n21739 );
and ( n26444 , n24631 , n21737 );
nor ( n26445 , n26443 , n26444 );
xnor ( n26446 , n26445 , n21749 );
and ( n26447 , n26442 , n26446 );
xor ( n26448 , n26362 , n26366 );
and ( n26449 , n26446 , n26448 );
and ( n26450 , n26442 , n26448 );
or ( n26451 , n26447 , n26449 , n26450 );
and ( n26452 , n21756 , n22032 );
and ( n26453 , n21519 , n22029 );
nor ( n26454 , n26452 , n26453 );
xnor ( n26455 , n26454 , n22027 );
and ( n26456 , n21630 , n22114 );
and ( n26457 , n21645 , n22112 );
nor ( n26458 , n26456 , n26457 );
xnor ( n26459 , n26458 , n22124 );
and ( n26460 , n26455 , n26459 );
and ( n26461 , n21486 , n21414 );
and ( n26462 , n21501 , n21412 );
nor ( n26463 , n26461 , n26462 );
xnor ( n26464 , n26463 , n21480 );
and ( n26465 , n21599 , n21139 );
and ( n26466 , n21545 , n21137 );
nor ( n26467 , n26465 , n26466 );
xnor ( n26468 , n26467 , n21221 );
and ( n26469 , n26464 , n26468 );
and ( n26470 , n21606 , n21663 );
and ( n26471 , n21511 , n21661 );
nor ( n26472 , n26470 , n26471 );
xnor ( n26473 , n26472 , n21673 );
and ( n26474 , n26468 , n26473 );
and ( n26475 , n26464 , n26473 );
or ( n26476 , n26469 , n26474 , n26475 );
and ( n26477 , n26460 , n26476 );
and ( n26478 , n22813 , n21687 );
and ( n26479 , n21616 , n21685 );
nor ( n26480 , n26478 , n26479 );
xnor ( n26481 , n26480 , n21697 );
and ( n26482 , n23320 , n21707 );
and ( n26483 , n23074 , n21705 );
nor ( n26484 , n26482 , n26483 );
xnor ( n26485 , n26484 , n21717 );
and ( n26486 , n26481 , n26485 );
and ( n26487 , n23503 , n21236 );
and ( n26488 , n23351 , n21234 );
nor ( n26489 , n26487 , n26488 );
xnor ( n26490 , n26489 , n21246 );
and ( n26491 , n26485 , n26490 );
and ( n26492 , n26481 , n26490 );
or ( n26493 , n26486 , n26491 , n26492 );
and ( n26494 , n26476 , n26493 );
and ( n26495 , n26460 , n26493 );
or ( n26496 , n26477 , n26494 , n26495 );
and ( n26497 , n26451 , n26496 );
and ( n26498 , n23887 , n21260 );
and ( n26499 , n23651 , n21258 );
nor ( n26500 , n26498 , n26499 );
xnor ( n26501 , n26500 , n21270 );
and ( n26502 , n24213 , n21582 );
and ( n26503 , n23949 , n21580 );
nor ( n26504 , n26502 , n26503 );
xnor ( n26505 , n26504 , n21588 );
and ( n26506 , n26501 , n26505 );
and ( n26507 , n24631 , n21783 );
and ( n26508 , n24460 , n21781 );
nor ( n26509 , n26507 , n26508 );
xnor ( n26510 , n26509 , n21793 );
and ( n26511 , n26505 , n26510 );
and ( n26512 , n26501 , n26510 );
or ( n26513 , n26506 , n26511 , n26512 );
xor ( n26514 , n26372 , n26376 );
xor ( n26515 , n26514 , n26381 );
and ( n26516 , n26513 , n26515 );
xor ( n26517 , n26391 , n26395 );
xor ( n26518 , n26517 , n26400 );
and ( n26519 , n26515 , n26518 );
and ( n26520 , n26513 , n26518 );
or ( n26521 , n26516 , n26519 , n26520 );
and ( n26522 , n26496 , n26521 );
and ( n26523 , n26451 , n26521 );
or ( n26524 , n26497 , n26522 , n26523 );
and ( n26525 , n26438 , n26524 );
xor ( n26526 , n26387 , n26411 );
xor ( n26527 , n26526 , n26414 );
and ( n26528 , n26524 , n26527 );
and ( n26529 , n26438 , n26527 );
or ( n26530 , n26525 , n26528 , n26529 );
and ( n26531 , n26436 , n26530 );
and ( n26532 , n21756 , n21414 );
and ( n26533 , n21519 , n21412 );
nor ( n26534 , n26532 , n26533 );
xnor ( n26535 , n26534 , n21480 );
and ( n26536 , n21630 , n21139 );
and ( n26537 , n21645 , n21137 );
nor ( n26538 , n26536 , n26537 );
xnor ( n26539 , n26538 , n21221 );
xor ( n26540 , n26535 , n26539 );
xor ( n26541 , n26193 , n26197 );
xor ( n26542 , n26541 , n26202 );
xor ( n26543 , n26540 , n26542 );
and ( n26544 , n26530 , n26543 );
and ( n26545 , n26436 , n26543 );
or ( n26546 , n26531 , n26544 , n26545 );
xor ( n26547 , n26354 , n26356 );
xor ( n26548 , n26547 , n26425 );
and ( n26549 , n26546 , n26548 );
xor ( n26550 , n26433 , n26435 );
xor ( n26551 , n26358 , n26367 );
xor ( n26552 , n26551 , n26384 );
xor ( n26553 , n26403 , n26405 );
xor ( n26554 , n26553 , n26408 );
and ( n26555 , n26552 , n26554 );
and ( n26556 , n24812 , n21739 );
and ( n26557 , n24662 , n21737 );
nor ( n26558 , n26556 , n26557 );
xnor ( n26559 , n26558 , n21749 );
and ( n26560 , n25179 , n21529 );
and ( n26561 , n25060 , n21527 );
nor ( n26562 , n26560 , n26561 );
xnor ( n26563 , n26562 , n21539 );
and ( n26564 , n26559 , n26563 );
xor ( n26565 , n26455 , n26459 );
and ( n26566 , n26563 , n26565 );
and ( n26567 , n26559 , n26565 );
or ( n26568 , n26564 , n26566 , n26567 );
and ( n26569 , n21645 , n22032 );
and ( n26570 , n21756 , n22029 );
nor ( n26571 , n26569 , n26570 );
xnor ( n26572 , n26571 , n22027 );
and ( n26573 , n21501 , n22114 );
and ( n26574 , n21630 , n22112 );
nor ( n26575 , n26573 , n26574 );
xnor ( n26576 , n26575 , n22124 );
and ( n26577 , n26572 , n26576 );
and ( n26578 , n21545 , n21414 );
and ( n26579 , n21486 , n21412 );
nor ( n26580 , n26578 , n26579 );
xnor ( n26581 , n26580 , n21480 );
and ( n26582 , n26576 , n26581 );
and ( n26583 , n26572 , n26581 );
or ( n26584 , n26577 , n26582 , n26583 );
and ( n26585 , n21511 , n21139 );
and ( n26586 , n21599 , n21137 );
nor ( n26587 , n26585 , n26586 );
xnor ( n26588 , n26587 , n21221 );
and ( n26589 , n21616 , n21663 );
and ( n26590 , n21606 , n21661 );
nor ( n26591 , n26589 , n26590 );
xnor ( n26592 , n26591 , n21673 );
and ( n26593 , n26588 , n26592 );
and ( n26594 , n23074 , n21687 );
and ( n26595 , n22813 , n21685 );
nor ( n26596 , n26594 , n26595 );
xnor ( n26597 , n26596 , n21697 );
and ( n26598 , n26592 , n26597 );
and ( n26599 , n26588 , n26597 );
or ( n26600 , n26593 , n26598 , n26599 );
and ( n26601 , n26584 , n26600 );
and ( n26602 , n23351 , n21707 );
and ( n26603 , n23320 , n21705 );
nor ( n26604 , n26602 , n26603 );
xnor ( n26605 , n26604 , n21717 );
and ( n26606 , n23651 , n21236 );
and ( n26607 , n23503 , n21234 );
nor ( n26608 , n26606 , n26607 );
xnor ( n26609 , n26608 , n21246 );
and ( n26610 , n26605 , n26609 );
and ( n26611 , n23949 , n21260 );
and ( n26612 , n23887 , n21258 );
nor ( n26613 , n26611 , n26612 );
xnor ( n26614 , n26613 , n21270 );
and ( n26615 , n26609 , n26614 );
and ( n26616 , n26605 , n26614 );
or ( n26617 , n26610 , n26615 , n26616 );
and ( n26618 , n26600 , n26617 );
and ( n26619 , n26584 , n26617 );
or ( n26620 , n26601 , n26618 , n26619 );
and ( n26621 , n26568 , n26620 );
and ( n26622 , n24460 , n21582 );
and ( n26623 , n24213 , n21580 );
nor ( n26624 , n26622 , n26623 );
xnor ( n26625 , n26624 , n21588 );
and ( n26626 , n24662 , n21783 );
and ( n26627 , n24631 , n21781 );
nor ( n26628 , n26626 , n26627 );
xnor ( n26629 , n26628 , n21793 );
and ( n26630 , n26625 , n26629 );
and ( n26631 , n25060 , n21739 );
and ( n26632 , n24812 , n21737 );
nor ( n26633 , n26631 , n26632 );
xnor ( n26634 , n26633 , n21749 );
and ( n26635 , n26629 , n26634 );
and ( n26636 , n26625 , n26634 );
or ( n26637 , n26630 , n26635 , n26636 );
xor ( n26638 , n26464 , n26468 );
xor ( n26639 , n26638 , n26473 );
and ( n26640 , n26637 , n26639 );
xor ( n26641 , n26481 , n26485 );
xor ( n26642 , n26641 , n26490 );
and ( n26643 , n26639 , n26642 );
and ( n26644 , n26637 , n26642 );
or ( n26645 , n26640 , n26643 , n26644 );
and ( n26646 , n26620 , n26645 );
and ( n26647 , n26568 , n26645 );
or ( n26648 , n26621 , n26646 , n26647 );
and ( n26649 , n26554 , n26648 );
and ( n26650 , n26552 , n26648 );
or ( n26651 , n26555 , n26649 , n26650 );
and ( n26652 , n26550 , n26651 );
xor ( n26653 , n26438 , n26524 );
xor ( n26654 , n26653 , n26527 );
and ( n26655 , n26651 , n26654 );
and ( n26656 , n26550 , n26654 );
or ( n26657 , n26652 , n26655 , n26656 );
xor ( n26658 , n26417 , n26419 );
xor ( n26659 , n26658 , n26422 );
and ( n26660 , n26657 , n26659 );
xor ( n26661 , n26436 , n26530 );
xor ( n26662 , n26661 , n26543 );
and ( n26663 , n26659 , n26662 );
and ( n26664 , n26657 , n26662 );
or ( n26665 , n26660 , n26663 , n26664 );
and ( n26666 , n26548 , n26665 );
and ( n26667 , n26546 , n26665 );
or ( n26668 , n26549 , n26666 , n26667 );
and ( n26669 , n26428 , n26668 );
and ( n26670 , n26352 , n26668 );
or ( n26671 , n26429 , n26669 , n26670 );
and ( n26672 , n26251 , n26671 );
and ( n26673 , n21645 , n21139 );
and ( n26674 , n21756 , n21137 );
nor ( n26675 , n26673 , n26674 );
xnor ( n26676 , n26675 , n21221 );
xor ( n26677 , n26122 , n26126 );
xor ( n26678 , n26677 , n26129 );
and ( n26679 , n26676 , n26678 );
xor ( n26680 , n26078 , n26082 );
xor ( n26681 , n26680 , n26085 );
and ( n26682 , n26678 , n26681 );
and ( n26683 , n26676 , n26681 );
or ( n26684 , n26679 , n26682 , n26683 );
xor ( n26685 , n25947 , n25951 );
xor ( n26686 , n26685 , n25954 );
and ( n26687 , n26684 , n26686 );
and ( n26688 , n26671 , n26687 );
and ( n26689 , n26251 , n26687 );
or ( n26690 , n26672 , n26688 , n26689 );
and ( n26691 , n26249 , n26690 );
xor ( n26692 , n26233 , n26235 );
xor ( n26693 , n26692 , n26238 );
and ( n26694 , n26690 , n26693 );
and ( n26695 , n26249 , n26693 );
or ( n26696 , n26691 , n26694 , n26695 );
xor ( n26697 , n26176 , n26178 );
xor ( n26698 , n26697 , n26241 );
and ( n26699 , n26696 , n26698 );
xor ( n26700 , n26225 , n26227 );
xor ( n26701 , n26700 , n26230 );
and ( n26702 , n25544 , n21625 );
and ( n26703 , n25343 , n21623 );
nor ( n26704 , n26702 , n26703 );
xnor ( n26705 , n26704 , n21635 );
and ( n26706 , n25772 , n21496 );
and ( n26707 , n25553 , n21494 );
nor ( n26708 , n26706 , n26707 );
xnor ( n26709 , n26708 , n21506 );
and ( n26710 , n26705 , n26709 );
xor ( n26711 , n26028 , n26032 );
xor ( n26712 , n26711 , n26034 );
and ( n26713 , n26709 , n26712 );
and ( n26714 , n26705 , n26712 );
or ( n26715 , n26710 , n26713 , n26714 );
and ( n26716 , n25060 , n21529 );
and ( n26717 , n24812 , n21527 );
nor ( n26718 , n26716 , n26717 );
xnor ( n26719 , n26718 , n21539 );
and ( n26720 , n26715 , n26719 );
and ( n26721 , n25343 , n21625 );
and ( n26722 , n25179 , n21623 );
nor ( n26723 , n26721 , n26722 );
xnor ( n26724 , n26723 , n21635 );
and ( n26725 , n25553 , n21496 );
and ( n26726 , n25544 , n21494 );
nor ( n26727 , n26725 , n26726 );
xnor ( n26728 , n26727 , n21506 );
xor ( n26729 , n26724 , n26728 );
xor ( n26730 , n26037 , n26041 );
xor ( n26731 , n26730 , n26043 );
xor ( n26732 , n26729 , n26731 );
and ( n26733 , n26719 , n26732 );
and ( n26734 , n26715 , n26732 );
or ( n26735 , n26720 , n26733 , n26734 );
and ( n26736 , n24213 , n21783 );
and ( n26737 , n23949 , n21781 );
nor ( n26738 , n26736 , n26737 );
xnor ( n26739 , n26738 , n21793 );
and ( n26740 , n26735 , n26739 );
xor ( n26741 , n26046 , n26050 );
xor ( n26742 , n26741 , n26053 );
and ( n26743 , n26739 , n26742 );
and ( n26744 , n26735 , n26742 );
or ( n26745 , n26740 , n26743 , n26744 );
and ( n26746 , n21511 , n21687 );
and ( n26747 , n21599 , n21685 );
nor ( n26748 , n26746 , n26747 );
xnor ( n26749 , n26748 , n21697 );
and ( n26750 , n26745 , n26749 );
xor ( n26751 , n26056 , n26060 );
xor ( n26752 , n26751 , n26065 );
and ( n26753 , n26749 , n26752 );
and ( n26754 , n26745 , n26752 );
or ( n26755 , n26750 , n26753 , n26754 );
and ( n26756 , n21486 , n21663 );
and ( n26757 , n21501 , n21661 );
nor ( n26758 , n26756 , n26757 );
xnor ( n26759 , n26758 , n21673 );
and ( n26760 , n26755 , n26759 );
and ( n26761 , n21599 , n21687 );
and ( n26762 , n21545 , n21685 );
nor ( n26763 , n26761 , n26762 );
xnor ( n26764 , n26763 , n21697 );
and ( n26765 , n26759 , n26764 );
and ( n26766 , n26755 , n26764 );
or ( n26767 , n26760 , n26765 , n26766 );
and ( n26768 , n22089 , n22032 );
and ( n26769 , n21777 , n22029 );
nor ( n26770 , n26768 , n26769 );
xnor ( n26771 , n26770 , n22027 );
and ( n26772 , n26767 , n26771 );
xor ( n26773 , n26205 , n26209 );
xor ( n26774 , n26773 , n26214 );
and ( n26775 , n26771 , n26774 );
and ( n26776 , n26767 , n26774 );
or ( n26777 , n26772 , n26775 , n26776 );
xor ( n26778 , n25961 , n25965 );
xor ( n26779 , n26778 , n25978 );
and ( n26780 , n26777 , n26779 );
xor ( n26781 , n26217 , n26219 );
xor ( n26782 , n26781 , n26222 );
and ( n26783 , n26779 , n26782 );
and ( n26784 , n26777 , n26782 );
or ( n26785 , n26780 , n26783 , n26784 );
and ( n26786 , n26701 , n26785 );
xor ( n26787 , n26352 , n26428 );
xor ( n26788 , n26787 , n26668 );
xor ( n26789 , n26684 , n26686 );
and ( n26790 , n26788 , n26789 );
and ( n26791 , n26535 , n26539 );
and ( n26792 , n26539 , n26542 );
and ( n26793 , n26535 , n26542 );
or ( n26794 , n26791 , n26792 , n26793 );
xor ( n26795 , n26676 , n26678 );
xor ( n26796 , n26795 , n26681 );
and ( n26797 , n26794 , n26796 );
and ( n26798 , n26789 , n26797 );
and ( n26799 , n26788 , n26797 );
or ( n26800 , n26790 , n26798 , n26799 );
and ( n26801 , n26785 , n26800 );
and ( n26802 , n26701 , n26800 );
or ( n26803 , n26786 , n26801 , n26802 );
xor ( n26804 , n26251 , n26671 );
xor ( n26805 , n26804 , n26687 );
xor ( n26806 , n26777 , n26779 );
xor ( n26807 , n26806 , n26782 );
xor ( n26808 , n26068 , n26072 );
xor ( n26809 , n26808 , n26075 );
xor ( n26810 , n26442 , n26446 );
xor ( n26811 , n26810 , n26448 );
xor ( n26812 , n26460 , n26476 );
xor ( n26813 , n26812 , n26493 );
and ( n26814 , n26811 , n26813 );
xor ( n26815 , n26513 , n26515 );
xor ( n26816 , n26815 , n26518 );
and ( n26817 , n26813 , n26816 );
and ( n26818 , n26811 , n26816 );
or ( n26819 , n26814 , n26817 , n26818 );
xor ( n26820 , n26451 , n26496 );
xor ( n26821 , n26820 , n26521 );
and ( n26822 , n26819 , n26821 );
xor ( n26823 , n26501 , n26505 );
xor ( n26824 , n26823 , n26510 );
and ( n26825 , n25343 , n21529 );
and ( n26826 , n25179 , n21527 );
nor ( n26827 , n26825 , n26826 );
xnor ( n26828 , n26827 , n21539 );
and ( n26829 , n25553 , n21625 );
and ( n26830 , n25544 , n21623 );
nor ( n26831 , n26829 , n26830 );
xnor ( n26832 , n26831 , n21635 );
and ( n26833 , n26828 , n26832 );
and ( n26834 , n21630 , n22032 );
and ( n26835 , n21645 , n22029 );
nor ( n26836 , n26834 , n26835 );
xnor ( n26837 , n26836 , n22027 );
and ( n26838 , n21486 , n22114 );
and ( n26839 , n21501 , n22112 );
nor ( n26840 , n26838 , n26839 );
xnor ( n26841 , n26840 , n22124 );
and ( n26842 , n26837 , n26841 );
and ( n26843 , n21599 , n21414 );
and ( n26844 , n21545 , n21412 );
nor ( n26845 , n26843 , n26844 );
xnor ( n26846 , n26845 , n21480 );
and ( n26847 , n26841 , n26846 );
and ( n26848 , n26837 , n26846 );
or ( n26849 , n26842 , n26847 , n26848 );
and ( n26850 , n26832 , n26849 );
and ( n26851 , n26828 , n26849 );
or ( n26852 , n26833 , n26850 , n26851 );
and ( n26853 , n26824 , n26852 );
and ( n26854 , n21606 , n21139 );
and ( n26855 , n21511 , n21137 );
nor ( n26856 , n26854 , n26855 );
xnor ( n26857 , n26856 , n21221 );
and ( n26858 , n22813 , n21663 );
and ( n26859 , n21616 , n21661 );
nor ( n26860 , n26858 , n26859 );
xnor ( n26861 , n26860 , n21673 );
and ( n26862 , n26857 , n26861 );
and ( n26863 , n23320 , n21687 );
and ( n26864 , n23074 , n21685 );
nor ( n26865 , n26863 , n26864 );
xnor ( n26866 , n26865 , n21697 );
and ( n26867 , n26861 , n26866 );
and ( n26868 , n26857 , n26866 );
or ( n26869 , n26862 , n26867 , n26868 );
and ( n26870 , n23503 , n21707 );
and ( n26871 , n23351 , n21705 );
nor ( n26872 , n26870 , n26871 );
xnor ( n26873 , n26872 , n21717 );
and ( n26874 , n23887 , n21236 );
and ( n26875 , n23651 , n21234 );
nor ( n26876 , n26874 , n26875 );
xnor ( n26877 , n26876 , n21246 );
and ( n26878 , n26873 , n26877 );
and ( n26879 , n24213 , n21260 );
and ( n26880 , n23949 , n21258 );
nor ( n26881 , n26879 , n26880 );
xnor ( n26882 , n26881 , n21270 );
and ( n26883 , n26877 , n26882 );
and ( n26884 , n26873 , n26882 );
or ( n26885 , n26878 , n26883 , n26884 );
and ( n26886 , n26869 , n26885 );
and ( n26887 , n24631 , n21582 );
and ( n26888 , n24460 , n21580 );
nor ( n26889 , n26887 , n26888 );
xnor ( n26890 , n26889 , n21588 );
and ( n26891 , n24812 , n21783 );
and ( n26892 , n24662 , n21781 );
nor ( n26893 , n26891 , n26892 );
xnor ( n26894 , n26893 , n21793 );
and ( n26895 , n26890 , n26894 );
and ( n26896 , n25179 , n21739 );
and ( n26897 , n25060 , n21737 );
nor ( n26898 , n26896 , n26897 );
xnor ( n26899 , n26898 , n21749 );
and ( n26900 , n26894 , n26899 );
and ( n26901 , n26890 , n26899 );
or ( n26902 , n26895 , n26900 , n26901 );
and ( n26903 , n26885 , n26902 );
and ( n26904 , n26869 , n26902 );
or ( n26905 , n26886 , n26903 , n26904 );
and ( n26906 , n26852 , n26905 );
and ( n26907 , n26824 , n26905 );
or ( n26908 , n26853 , n26906 , n26907 );
xor ( n26909 , n26572 , n26576 );
xor ( n26910 , n26909 , n26581 );
xor ( n26911 , n26588 , n26592 );
xor ( n26912 , n26911 , n26597 );
and ( n26913 , n26910 , n26912 );
xor ( n26914 , n26605 , n26609 );
xor ( n26915 , n26914 , n26614 );
and ( n26916 , n26912 , n26915 );
and ( n26917 , n26910 , n26915 );
or ( n26918 , n26913 , n26916 , n26917 );
xor ( n26919 , n26559 , n26563 );
xor ( n26920 , n26919 , n26565 );
and ( n26921 , n26918 , n26920 );
xor ( n26922 , n26584 , n26600 );
xor ( n26923 , n26922 , n26617 );
and ( n26924 , n26920 , n26923 );
and ( n26925 , n26918 , n26923 );
or ( n26926 , n26921 , n26924 , n26925 );
and ( n26927 , n26908 , n26926 );
xor ( n26928 , n26568 , n26620 );
xor ( n26929 , n26928 , n26645 );
and ( n26930 , n26926 , n26929 );
and ( n26931 , n26908 , n26929 );
or ( n26932 , n26927 , n26930 , n26931 );
and ( n26933 , n26821 , n26932 );
and ( n26934 , n26819 , n26932 );
or ( n26935 , n26822 , n26933 , n26934 );
xor ( n26936 , n26550 , n26651 );
xor ( n26937 , n26936 , n26654 );
and ( n26938 , n26935 , n26937 );
and ( n26939 , n26724 , n26728 );
and ( n26940 , n26728 , n26731 );
and ( n26941 , n26724 , n26731 );
or ( n26942 , n26939 , n26940 , n26941 );
and ( n26943 , n24631 , n21739 );
and ( n26944 , n24460 , n21737 );
nor ( n26945 , n26943 , n26944 );
xnor ( n26946 , n26945 , n21749 );
and ( n26947 , n26942 , n26946 );
and ( n26948 , n24812 , n21529 );
and ( n26949 , n24662 , n21527 );
nor ( n26950 , n26948 , n26949 );
xnor ( n26951 , n26950 , n21539 );
and ( n26952 , n26946 , n26951 );
and ( n26953 , n26942 , n26951 );
or ( n26954 , n26947 , n26952 , n26953 );
and ( n26955 , n26937 , n26954 );
and ( n26956 , n26935 , n26954 );
or ( n26957 , n26938 , n26955 , n26956 );
and ( n26958 , n26809 , n26957 );
xor ( n26959 , n26657 , n26659 );
xor ( n26960 , n26959 , n26662 );
and ( n26961 , n26957 , n26960 );
and ( n26962 , n26809 , n26960 );
or ( n26963 , n26958 , n26961 , n26962 );
xor ( n26964 , n26546 , n26548 );
xor ( n26965 , n26964 , n26665 );
and ( n26966 , n26963 , n26965 );
xor ( n26967 , n26767 , n26771 );
xor ( n26968 , n26967 , n26774 );
and ( n26969 , n26965 , n26968 );
and ( n26970 , n26963 , n26968 );
or ( n26971 , n26966 , n26969 , n26970 );
and ( n26972 , n26807 , n26971 );
xor ( n26973 , n26788 , n26789 );
xor ( n26974 , n26973 , n26797 );
and ( n26975 , n26971 , n26974 );
and ( n26976 , n26807 , n26974 );
or ( n26977 , n26972 , n26975 , n26976 );
and ( n26978 , n26805 , n26977 );
xor ( n26979 , n26701 , n26785 );
xor ( n26980 , n26979 , n26800 );
and ( n26981 , n26977 , n26980 );
and ( n26982 , n26805 , n26980 );
or ( n26983 , n26978 , n26981 , n26982 );
and ( n26984 , n26803 , n26983 );
xor ( n26985 , n26249 , n26690 );
xor ( n26986 , n26985 , n26693 );
and ( n26987 , n26983 , n26986 );
and ( n26988 , n26803 , n26986 );
or ( n26989 , n26984 , n26987 , n26988 );
and ( n26990 , n26698 , n26989 );
and ( n26991 , n26696 , n26989 );
or ( n26992 , n26699 , n26990 , n26991 );
and ( n26993 , n26246 , n26992 );
and ( n26994 , n26244 , n26992 );
or ( n26995 , n26247 , n26993 , n26994 );
and ( n26996 , n26174 , n26995 );
xor ( n26997 , n26174 , n26995 );
xor ( n26998 , n26244 , n26246 );
xor ( n26999 , n26998 , n26992 );
xor ( n27000 , n26696 , n26698 );
xor ( n27001 , n27000 , n26989 );
xor ( n27002 , n26803 , n26983 );
xor ( n27003 , n27002 , n26986 );
xor ( n27004 , n26805 , n26977 );
xor ( n27005 , n27004 , n26980 );
xor ( n27006 , n26794 , n26796 );
xor ( n27007 , n26552 , n26554 );
xor ( n27008 , n27007 , n26648 );
xor ( n27009 , n26811 , n26813 );
xor ( n27010 , n27009 , n26816 );
xor ( n27011 , n26637 , n26639 );
xor ( n27012 , n27011 , n26642 );
and ( n27013 , n25898 , n21496 );
and ( n27014 , n25772 , n21494 );
nor ( n27015 , n27013 , n27014 );
xnor ( n27016 , n27015 , n21506 );
xor ( n27017 , n26015 , n26023 );
xor ( n27018 , n27017 , n26025 );
and ( n27019 , n27016 , n27018 );
and ( n27020 , n27012 , n27019 );
xor ( n27021 , n26625 , n26629 );
xor ( n27022 , n27021 , n26634 );
and ( n27023 , n26020 , n21496 );
and ( n27024 , n25898 , n21494 );
nor ( n27025 , n27023 , n27024 );
xnor ( n27026 , n27025 , n21506 );
xor ( n27027 , n26006 , n26014 );
and ( n27028 , n27026 , n27027 );
and ( n27029 , n27022 , n27028 );
and ( n27030 , n25544 , n21529 );
and ( n27031 , n25343 , n21527 );
nor ( n27032 , n27030 , n27031 );
xnor ( n27033 , n27032 , n21539 );
and ( n27034 , n25772 , n21625 );
and ( n27035 , n25553 , n21623 );
nor ( n27036 , n27034 , n27035 );
xnor ( n27037 , n27036 , n21635 );
and ( n27038 , n27033 , n27037 );
and ( n27039 , n26011 , n21496 );
and ( n27040 , n26020 , n21494 );
nor ( n27041 , n27039 , n27040 );
xnor ( n27042 , n27041 , n21506 );
and ( n27043 , n27042 , n26004 );
and ( n27044 , n27037 , n27043 );
and ( n27045 , n27033 , n27043 );
or ( n27046 , n27038 , n27044 , n27045 );
and ( n27047 , n27028 , n27046 );
and ( n27048 , n27022 , n27046 );
or ( n27049 , n27029 , n27047 , n27048 );
and ( n27050 , n27019 , n27049 );
and ( n27051 , n27012 , n27049 );
or ( n27052 , n27020 , n27050 , n27051 );
and ( n27053 , n27010 , n27052 );
and ( n27054 , n21501 , n22032 );
and ( n27055 , n21630 , n22029 );
nor ( n27056 , n27054 , n27055 );
xnor ( n27057 , n27056 , n22027 );
and ( n27058 , n23651 , n21707 );
and ( n27059 , n23503 , n21705 );
nor ( n27060 , n27058 , n27059 );
xnor ( n27061 , n27060 , n21717 );
and ( n27062 , n27057 , n27061 );
and ( n27063 , n23949 , n21236 );
and ( n27064 , n23887 , n21234 );
nor ( n27065 , n27063 , n27064 );
xnor ( n27066 , n27065 , n21246 );
and ( n27067 , n27061 , n27066 );
and ( n27068 , n27057 , n27066 );
or ( n27069 , n27062 , n27067 , n27068 );
and ( n27070 , n25060 , n21783 );
and ( n27071 , n24812 , n21781 );
nor ( n27072 , n27070 , n27071 );
xnor ( n27073 , n27072 , n21793 );
and ( n27074 , n25343 , n21739 );
and ( n27075 , n25179 , n21737 );
nor ( n27076 , n27074 , n27075 );
xnor ( n27077 , n27076 , n21749 );
and ( n27078 , n27073 , n27077 );
and ( n27079 , n25553 , n21529 );
and ( n27080 , n25544 , n21527 );
nor ( n27081 , n27079 , n27080 );
xnor ( n27082 , n27081 , n21539 );
and ( n27083 , n27077 , n27082 );
and ( n27084 , n27073 , n27082 );
or ( n27085 , n27078 , n27083 , n27084 );
and ( n27086 , n27069 , n27085 );
xor ( n27087 , n26837 , n26841 );
xor ( n27088 , n27087 , n26846 );
and ( n27089 , n27085 , n27088 );
and ( n27090 , n27069 , n27088 );
or ( n27091 , n27086 , n27089 , n27090 );
xor ( n27092 , n26857 , n26861 );
xor ( n27093 , n27092 , n26866 );
xor ( n27094 , n26873 , n26877 );
xor ( n27095 , n27094 , n26882 );
and ( n27096 , n27093 , n27095 );
xor ( n27097 , n26890 , n26894 );
xor ( n27098 , n27097 , n26899 );
and ( n27099 , n27095 , n27098 );
and ( n27100 , n27093 , n27098 );
or ( n27101 , n27096 , n27099 , n27100 );
and ( n27102 , n27091 , n27101 );
xor ( n27103 , n26828 , n26832 );
xor ( n27104 , n27103 , n26849 );
and ( n27105 , n27101 , n27104 );
and ( n27106 , n27091 , n27104 );
or ( n27107 , n27102 , n27105 , n27106 );
xor ( n27108 , n26824 , n26852 );
xor ( n27109 , n27108 , n26905 );
and ( n27110 , n27107 , n27109 );
xor ( n27111 , n26918 , n26920 );
xor ( n27112 , n27111 , n26923 );
and ( n27113 , n27109 , n27112 );
and ( n27114 , n27107 , n27112 );
or ( n27115 , n27110 , n27113 , n27114 );
and ( n27116 , n27052 , n27115 );
and ( n27117 , n27010 , n27115 );
or ( n27118 , n27053 , n27116 , n27117 );
and ( n27119 , n27008 , n27118 );
xor ( n27120 , n26819 , n26821 );
xor ( n27121 , n27120 , n26932 );
and ( n27122 , n27118 , n27121 );
and ( n27123 , n27008 , n27121 );
or ( n27124 , n27119 , n27122 , n27123 );
xor ( n27125 , n26942 , n26946 );
xor ( n27126 , n27125 , n26951 );
xor ( n27127 , n26908 , n26926 );
xor ( n27128 , n27127 , n26929 );
xor ( n27129 , n26705 , n26709 );
xor ( n27130 , n27129 , n26712 );
xor ( n27131 , n26869 , n26885 );
xor ( n27132 , n27131 , n26902 );
xor ( n27133 , n26910 , n26912 );
xor ( n27134 , n27133 , n26915 );
and ( n27135 , n27132 , n27134 );
xor ( n27136 , n27016 , n27018 );
and ( n27137 , n27134 , n27136 );
and ( n27138 , n27132 , n27136 );
or ( n27139 , n27135 , n27137 , n27138 );
and ( n27140 , n27130 , n27139 );
xor ( n27141 , n27026 , n27027 );
and ( n27142 , n25898 , n21625 );
and ( n27143 , n25772 , n21623 );
nor ( n27144 , n27142 , n27143 );
xnor ( n27145 , n27144 , n21635 );
xor ( n27146 , n27042 , n26004 );
and ( n27147 , n27145 , n27146 );
and ( n27148 , n26003 , n21494 );
not ( n27149 , n27148 );
and ( n27150 , n27149 , n21506 );
and ( n27151 , n26003 , n21496 );
and ( n27152 , n26011 , n21494 );
nor ( n27153 , n27151 , n27152 );
xnor ( n27154 , n27153 , n21506 );
and ( n27155 , n27150 , n27154 );
and ( n27156 , n27146 , n27155 );
and ( n27157 , n27145 , n27155 );
or ( n27158 , n27147 , n27156 , n27157 );
and ( n27159 , n27141 , n27158 );
xor ( n27160 , n27033 , n27037 );
xor ( n27161 , n27160 , n27043 );
and ( n27162 , n27158 , n27161 );
and ( n27163 , n27141 , n27161 );
or ( n27164 , n27159 , n27162 , n27163 );
xor ( n27165 , n27022 , n27028 );
xor ( n27166 , n27165 , n27046 );
and ( n27167 , n27164 , n27166 );
xor ( n27168 , n27091 , n27101 );
xor ( n27169 , n27168 , n27104 );
and ( n27170 , n27166 , n27169 );
and ( n27171 , n27164 , n27169 );
or ( n27172 , n27167 , n27170 , n27171 );
and ( n27173 , n27139 , n27172 );
and ( n27174 , n27130 , n27172 );
or ( n27175 , n27140 , n27173 , n27174 );
and ( n27176 , n27128 , n27175 );
xor ( n27177 , n27010 , n27052 );
xor ( n27178 , n27177 , n27115 );
and ( n27179 , n27175 , n27178 );
and ( n27180 , n27128 , n27178 );
or ( n27181 , n27176 , n27179 , n27180 );
and ( n27182 , n27126 , n27181 );
xor ( n27183 , n27008 , n27118 );
xor ( n27184 , n27183 , n27121 );
and ( n27185 , n27181 , n27184 );
and ( n27186 , n27126 , n27184 );
or ( n27187 , n27182 , n27185 , n27186 );
and ( n27188 , n27124 , n27187 );
xor ( n27189 , n26935 , n26937 );
xor ( n27190 , n27189 , n26954 );
and ( n27191 , n27187 , n27190 );
and ( n27192 , n27124 , n27190 );
or ( n27193 , n27188 , n27191 , n27192 );
xor ( n27194 , n26809 , n26957 );
xor ( n27195 , n27194 , n26960 );
and ( n27196 , n27193 , n27195 );
xor ( n27197 , n26755 , n26759 );
xor ( n27198 , n27197 , n26764 );
and ( n27199 , n27195 , n27198 );
and ( n27200 , n27193 , n27198 );
or ( n27201 , n27196 , n27199 , n27200 );
and ( n27202 , n27006 , n27201 );
and ( n27203 , n23651 , n21260 );
and ( n27204 , n23503 , n21258 );
nor ( n27205 , n27203 , n27204 );
xnor ( n27206 , n27205 , n21270 );
and ( n27207 , n23949 , n21582 );
and ( n27208 , n23887 , n21580 );
nor ( n27209 , n27207 , n27208 );
xnor ( n27210 , n27209 , n21588 );
and ( n27211 , n27206 , n27210 );
xor ( n27212 , n26715 , n26719 );
xor ( n27213 , n27212 , n26732 );
and ( n27214 , n27210 , n27213 );
and ( n27215 , n27206 , n27213 );
or ( n27216 , n27211 , n27214 , n27215 );
and ( n27217 , n21606 , n21687 );
and ( n27218 , n21511 , n21685 );
nor ( n27219 , n27217 , n27218 );
xnor ( n27220 , n27219 , n21697 );
and ( n27221 , n27216 , n27220 );
and ( n27222 , n22813 , n21707 );
and ( n27223 , n21616 , n21705 );
nor ( n27224 , n27222 , n27223 );
xnor ( n27225 , n27224 , n21717 );
and ( n27226 , n27220 , n27225 );
and ( n27227 , n27216 , n27225 );
or ( n27228 , n27221 , n27226 , n27227 );
and ( n27229 , n21519 , n22114 );
and ( n27230 , n21534 , n22112 );
nor ( n27231 , n27229 , n27230 );
xnor ( n27232 , n27231 , n22124 );
and ( n27233 , n27228 , n27232 );
and ( n27234 , n21501 , n21139 );
and ( n27235 , n21630 , n21137 );
nor ( n27236 , n27234 , n27235 );
xnor ( n27237 , n27236 , n21221 );
and ( n27238 , n27232 , n27237 );
and ( n27239 , n27228 , n27237 );
or ( n27240 , n27233 , n27238 , n27239 );
xor ( n27241 , n26745 , n26749 );
xor ( n27242 , n27241 , n26752 );
xor ( n27243 , n27124 , n27187 );
xor ( n27244 , n27243 , n27190 );
and ( n27245 , n27242 , n27244 );
xor ( n27246 , n27228 , n27232 );
xor ( n27247 , n27246 , n27237 );
and ( n27248 , n27244 , n27247 );
and ( n27249 , n27242 , n27247 );
or ( n27250 , n27245 , n27248 , n27249 );
and ( n27251 , n27240 , n27250 );
xor ( n27252 , n27193 , n27195 );
xor ( n27253 , n27252 , n27198 );
and ( n27254 , n27250 , n27253 );
and ( n27255 , n27240 , n27253 );
or ( n27256 , n27251 , n27254 , n27255 );
and ( n27257 , n27201 , n27256 );
and ( n27258 , n27006 , n27256 );
or ( n27259 , n27202 , n27257 , n27258 );
xor ( n27260 , n26807 , n26971 );
xor ( n27261 , n27260 , n26974 );
and ( n27262 , n27259 , n27261 );
xor ( n27263 , n27259 , n27261 );
xor ( n27264 , n26963 , n26965 );
xor ( n27265 , n27264 , n26968 );
xor ( n27266 , n27006 , n27201 );
xor ( n27267 , n27266 , n27256 );
and ( n27268 , n27265 , n27267 );
xor ( n27269 , n27265 , n27267 );
xor ( n27270 , n27240 , n27250 );
xor ( n27271 , n27270 , n27253 );
xor ( n27272 , n26735 , n26739 );
xor ( n27273 , n27272 , n26742 );
xor ( n27274 , n27126 , n27181 );
xor ( n27275 , n27274 , n27184 );
and ( n27276 , n27273 , n27275 );
xor ( n27277 , n27216 , n27220 );
xor ( n27278 , n27277 , n27225 );
and ( n27279 , n27275 , n27278 );
and ( n27280 , n27273 , n27278 );
or ( n27281 , n27276 , n27279 , n27280 );
xor ( n27282 , n27242 , n27244 );
xor ( n27283 , n27282 , n27247 );
and ( n27284 , n27281 , n27283 );
xor ( n27285 , n27281 , n27283 );
xor ( n27286 , n27012 , n27019 );
xor ( n27287 , n27286 , n27049 );
xor ( n27288 , n27107 , n27109 );
xor ( n27289 , n27288 , n27112 );
and ( n27290 , n27287 , n27289 );
xor ( n27291 , n27069 , n27085 );
xor ( n27292 , n27291 , n27088 );
xor ( n27293 , n27093 , n27095 );
xor ( n27294 , n27293 , n27098 );
and ( n27295 , n27292 , n27294 );
xor ( n27296 , n27057 , n27061 );
xor ( n27297 , n27296 , n27066 );
xor ( n27298 , n27073 , n27077 );
xor ( n27299 , n27298 , n27082 );
and ( n27300 , n27297 , n27299 );
xor ( n27301 , n27145 , n27146 );
xor ( n27302 , n27301 , n27155 );
and ( n27303 , n27299 , n27302 );
and ( n27304 , n27297 , n27302 );
or ( n27305 , n27300 , n27303 , n27304 );
and ( n27306 , n27294 , n27305 );
and ( n27307 , n27292 , n27305 );
or ( n27308 , n27295 , n27306 , n27307 );
xor ( n27309 , n27132 , n27134 );
xor ( n27310 , n27309 , n27136 );
and ( n27311 , n27308 , n27310 );
xor ( n27312 , n27164 , n27166 );
xor ( n27313 , n27312 , n27169 );
and ( n27314 , n27310 , n27313 );
and ( n27315 , n27308 , n27313 );
or ( n27316 , n27311 , n27314 , n27315 );
and ( n27317 , n27289 , n27316 );
and ( n27318 , n27287 , n27316 );
or ( n27319 , n27290 , n27317 , n27318 );
xor ( n27320 , n27128 , n27175 );
xor ( n27321 , n27320 , n27178 );
and ( n27322 , n27319 , n27321 );
xor ( n27323 , n27206 , n27210 );
xor ( n27324 , n27323 , n27213 );
and ( n27325 , n27321 , n27324 );
and ( n27326 , n27319 , n27324 );
or ( n27327 , n27322 , n27325 , n27326 );
xor ( n27328 , n27273 , n27275 );
xor ( n27329 , n27328 , n27278 );
and ( n27330 , n27327 , n27329 );
xor ( n27331 , n27327 , n27329 );
xor ( n27332 , n27319 , n27321 );
xor ( n27333 , n27332 , n27324 );
xor ( n27334 , n27130 , n27139 );
xor ( n27335 , n27334 , n27172 );
xor ( n27336 , n27287 , n27289 );
xor ( n27337 , n27336 , n27316 );
and ( n27338 , n27335 , n27337 );
xor ( n27339 , n27308 , n27310 );
xor ( n27340 , n27339 , n27313 );
xor ( n27341 , n27141 , n27158 );
xor ( n27342 , n27341 , n27161 );
xor ( n27343 , n27292 , n27294 );
xor ( n27344 , n27343 , n27305 );
and ( n27345 , n27342 , n27344 );
xor ( n27346 , n27150 , n27154 );
and ( n27347 , n26003 , n21623 );
not ( n27348 , n27347 );
and ( n27349 , n27348 , n21635 );
and ( n27350 , n26003 , n21625 );
and ( n27351 , n26011 , n21623 );
nor ( n27352 , n27350 , n27351 );
xnor ( n27353 , n27352 , n21635 );
and ( n27354 , n27349 , n27353 );
and ( n27355 , n26011 , n21625 );
and ( n27356 , n26020 , n21623 );
nor ( n27357 , n27355 , n27356 );
xnor ( n27358 , n27357 , n21635 );
and ( n27359 , n27354 , n27358 );
and ( n27360 , n27358 , n27148 );
and ( n27361 , n27354 , n27148 );
or ( n27362 , n27359 , n27360 , n27361 );
and ( n27363 , n27346 , n27362 );
and ( n27364 , n26020 , n21625 );
and ( n27365 , n25898 , n21623 );
nor ( n27366 , n27364 , n27365 );
xnor ( n27367 , n27366 , n21635 );
and ( n27368 , n27362 , n27367 );
and ( n27369 , n27346 , n27367 );
or ( n27370 , n27363 , n27368 , n27369 );
xor ( n27371 , n27297 , n27299 );
xor ( n27372 , n27371 , n27302 );
and ( n27373 , n27370 , n27372 );
and ( n27374 , n25544 , n21739 );
and ( n27375 , n25343 , n21737 );
nor ( n27376 , n27374 , n27375 );
xnor ( n27377 , n27376 , n21749 );
and ( n27378 , n25772 , n21529 );
and ( n27379 , n25553 , n21527 );
nor ( n27380 , n27378 , n27379 );
xnor ( n27381 , n27380 , n21539 );
and ( n27382 , n27377 , n27381 );
xor ( n27383 , n27346 , n27362 );
xor ( n27384 , n27383 , n27367 );
and ( n27385 , n27381 , n27384 );
and ( n27386 , n27377 , n27384 );
or ( n27387 , n27382 , n27385 , n27386 );
and ( n27388 , n27372 , n27387 );
and ( n27389 , n27370 , n27387 );
or ( n27390 , n27373 , n27388 , n27389 );
and ( n27391 , n27344 , n27390 );
and ( n27392 , n27342 , n27390 );
or ( n27393 , n27345 , n27391 , n27392 );
and ( n27394 , n27340 , n27393 );
xor ( n27395 , n27349 , n27353 );
and ( n27396 , n26003 , n21527 );
not ( n27397 , n27396 );
and ( n27398 , n27397 , n21539 );
and ( n27399 , n26003 , n21529 );
and ( n27400 , n26011 , n21527 );
nor ( n27401 , n27399 , n27400 );
xnor ( n27402 , n27401 , n21539 );
and ( n27403 , n27398 , n27402 );
and ( n27404 , n26011 , n21529 );
and ( n27405 , n26020 , n21527 );
nor ( n27406 , n27404 , n27405 );
xnor ( n27407 , n27406 , n21539 );
and ( n27408 , n27403 , n27407 );
and ( n27409 , n27407 , n27347 );
and ( n27410 , n27403 , n27347 );
or ( n27411 , n27408 , n27409 , n27410 );
and ( n27412 , n27395 , n27411 );
and ( n27413 , n26020 , n21529 );
and ( n27414 , n25898 , n21527 );
nor ( n27415 , n27413 , n27414 );
xnor ( n27416 , n27415 , n21539 );
and ( n27417 , n27411 , n27416 );
and ( n27418 , n27395 , n27416 );
or ( n27419 , n27412 , n27417 , n27418 );
and ( n27420 , n25898 , n21529 );
and ( n27421 , n25772 , n21527 );
nor ( n27422 , n27420 , n27421 );
xnor ( n27423 , n27422 , n21539 );
and ( n27424 , n27419 , n27423 );
xor ( n27425 , n27354 , n27358 );
xor ( n27426 , n27425 , n27148 );
and ( n27427 , n27423 , n27426 );
and ( n27428 , n27419 , n27426 );
or ( n27429 , n27424 , n27427 , n27428 );
and ( n27430 , n25179 , n21783 );
and ( n27431 , n25060 , n21781 );
nor ( n27432 , n27430 , n27431 );
xnor ( n27433 , n27432 , n21793 );
and ( n27434 , n27429 , n27433 );
xor ( n27435 , n27377 , n27381 );
xor ( n27436 , n27435 , n27384 );
and ( n27437 , n27433 , n27436 );
and ( n27438 , n27429 , n27436 );
or ( n27439 , n27434 , n27437 , n27438 );
and ( n27440 , n24460 , n21260 );
and ( n27441 , n24213 , n21258 );
nor ( n27442 , n27440 , n27441 );
xnor ( n27443 , n27442 , n21270 );
and ( n27444 , n27439 , n27443 );
and ( n27445 , n24662 , n21582 );
and ( n27446 , n24631 , n21580 );
nor ( n27447 , n27445 , n27446 );
xnor ( n27448 , n27447 , n21588 );
and ( n27449 , n27443 , n27448 );
and ( n27450 , n27439 , n27448 );
or ( n27451 , n27444 , n27449 , n27450 );
xor ( n27452 , n27342 , n27344 );
xor ( n27453 , n27452 , n27390 );
and ( n27454 , n27451 , n27453 );
and ( n27455 , n25343 , n21783 );
and ( n27456 , n25179 , n21781 );
nor ( n27457 , n27455 , n27456 );
xnor ( n27458 , n27457 , n21793 );
and ( n27459 , n25553 , n21739 );
and ( n27460 , n25544 , n21737 );
nor ( n27461 , n27459 , n27460 );
xnor ( n27462 , n27461 , n21749 );
and ( n27463 , n27458 , n27462 );
xor ( n27464 , n27419 , n27423 );
xor ( n27465 , n27464 , n27426 );
and ( n27466 , n27462 , n27465 );
and ( n27467 , n27458 , n27465 );
or ( n27468 , n27463 , n27466 , n27467 );
and ( n27469 , n24631 , n21260 );
and ( n27470 , n24460 , n21258 );
nor ( n27471 , n27469 , n27470 );
xnor ( n27472 , n27471 , n21270 );
and ( n27473 , n27468 , n27472 );
and ( n27474 , n24812 , n21582 );
and ( n27475 , n24662 , n21580 );
nor ( n27476 , n27474 , n27475 );
xnor ( n27477 , n27476 , n21588 );
and ( n27478 , n27472 , n27477 );
and ( n27479 , n27468 , n27477 );
or ( n27480 , n27473 , n27478 , n27479 );
and ( n27481 , n23074 , n21663 );
and ( n27482 , n22813 , n21661 );
nor ( n27483 , n27481 , n27482 );
xnor ( n27484 , n27483 , n21673 );
and ( n27485 , n27480 , n27484 );
xor ( n27486 , n27439 , n27443 );
xor ( n27487 , n27486 , n27448 );
and ( n27488 , n27484 , n27487 );
and ( n27489 , n27480 , n27487 );
or ( n27490 , n27485 , n27488 , n27489 );
and ( n27491 , n27453 , n27490 );
and ( n27492 , n27451 , n27490 );
or ( n27493 , n27454 , n27491 , n27492 );
and ( n27494 , n27393 , n27493 );
and ( n27495 , n27340 , n27493 );
or ( n27496 , n27394 , n27494 , n27495 );
and ( n27497 , n27337 , n27496 );
and ( n27498 , n27335 , n27496 );
or ( n27499 , n27338 , n27497 , n27498 );
and ( n27500 , n27333 , n27499 );
xor ( n27501 , n27333 , n27499 );
xor ( n27502 , n27335 , n27337 );
xor ( n27503 , n27502 , n27496 );
xor ( n27504 , n27398 , n27402 );
and ( n27505 , n26003 , n21737 );
not ( n27506 , n27505 );
and ( n27507 , n27506 , n21749 );
and ( n27508 , n26003 , n21739 );
and ( n27509 , n26011 , n21737 );
nor ( n27510 , n27508 , n27509 );
xnor ( n27511 , n27510 , n21749 );
and ( n27512 , n27507 , n27511 );
and ( n27513 , n26011 , n21739 );
and ( n27514 , n26020 , n21737 );
nor ( n27515 , n27513 , n27514 );
xnor ( n27516 , n27515 , n21749 );
and ( n27517 , n27512 , n27516 );
and ( n27518 , n27516 , n27396 );
and ( n27519 , n27512 , n27396 );
or ( n27520 , n27517 , n27518 , n27519 );
and ( n27521 , n27504 , n27520 );
and ( n27522 , n26020 , n21739 );
and ( n27523 , n25898 , n21737 );
nor ( n27524 , n27522 , n27523 );
xnor ( n27525 , n27524 , n21749 );
and ( n27526 , n27520 , n27525 );
and ( n27527 , n27504 , n27525 );
or ( n27528 , n27521 , n27526 , n27527 );
and ( n27529 , n25898 , n21739 );
and ( n27530 , n25772 , n21737 );
nor ( n27531 , n27529 , n27530 );
xnor ( n27532 , n27531 , n21749 );
and ( n27533 , n27528 , n27532 );
xor ( n27534 , n27403 , n27407 );
xor ( n27535 , n27534 , n27347 );
and ( n27536 , n27532 , n27535 );
and ( n27537 , n27528 , n27535 );
or ( n27538 , n27533 , n27536 , n27537 );
and ( n27539 , n25179 , n21582 );
and ( n27540 , n25060 , n21580 );
nor ( n27541 , n27539 , n27540 );
xnor ( n27542 , n27541 , n21588 );
and ( n27543 , n27538 , n27542 );
and ( n27544 , n25544 , n21783 );
and ( n27545 , n25343 , n21781 );
nor ( n27546 , n27544 , n27545 );
xnor ( n27547 , n27546 , n21793 );
and ( n27548 , n25772 , n21739 );
and ( n27549 , n25553 , n21737 );
nor ( n27550 , n27548 , n27549 );
xnor ( n27551 , n27550 , n21749 );
xor ( n27552 , n27547 , n27551 );
xor ( n27553 , n27395 , n27411 );
xor ( n27554 , n27553 , n27416 );
xor ( n27555 , n27552 , n27554 );
and ( n27556 , n27542 , n27555 );
and ( n27557 , n27538 , n27555 );
or ( n27558 , n27543 , n27556 , n27557 );
and ( n27559 , n24460 , n21236 );
and ( n27560 , n24213 , n21234 );
nor ( n27561 , n27559 , n27560 );
xnor ( n27562 , n27561 , n21246 );
and ( n27563 , n27558 , n27562 );
and ( n27564 , n24662 , n21260 );
and ( n27565 , n24631 , n21258 );
nor ( n27566 , n27564 , n27565 );
xnor ( n27567 , n27566 , n21270 );
and ( n27568 , n27562 , n27567 );
and ( n27569 , n27558 , n27567 );
or ( n27570 , n27563 , n27568 , n27569 );
and ( n27571 , n23887 , n21707 );
and ( n27572 , n23651 , n21705 );
nor ( n27573 , n27571 , n27572 );
xnor ( n27574 , n27573 , n21717 );
and ( n27575 , n27570 , n27574 );
xor ( n27576 , n27468 , n27472 );
xor ( n27577 , n27576 , n27477 );
and ( n27578 , n27574 , n27577 );
and ( n27579 , n27570 , n27577 );
or ( n27580 , n27575 , n27578 , n27579 );
and ( n27581 , n21511 , n21414 );
and ( n27582 , n21599 , n21412 );
nor ( n27583 , n27581 , n27582 );
xnor ( n27584 , n27583 , n21480 );
and ( n27585 , n27580 , n27584 );
and ( n27586 , n21616 , n21139 );
and ( n27587 , n21606 , n21137 );
nor ( n27588 , n27586 , n27587 );
xnor ( n27589 , n27588 , n21221 );
and ( n27590 , n27584 , n27589 );
and ( n27591 , n27580 , n27589 );
or ( n27592 , n27585 , n27590 , n27591 );
and ( n27593 , n27547 , n27551 );
and ( n27594 , n27551 , n27554 );
and ( n27595 , n27547 , n27554 );
or ( n27596 , n27593 , n27594 , n27595 );
and ( n27597 , n25060 , n21582 );
and ( n27598 , n24812 , n21580 );
nor ( n27599 , n27597 , n27598 );
xnor ( n27600 , n27599 , n21588 );
and ( n27601 , n27596 , n27600 );
xor ( n27602 , n27458 , n27462 );
xor ( n27603 , n27602 , n27465 );
and ( n27604 , n27600 , n27603 );
and ( n27605 , n27596 , n27603 );
or ( n27606 , n27601 , n27604 , n27605 );
and ( n27607 , n24213 , n21236 );
and ( n27608 , n23949 , n21234 );
nor ( n27609 , n27607 , n27608 );
xnor ( n27610 , n27609 , n21246 );
and ( n27611 , n27606 , n27610 );
xor ( n27612 , n27429 , n27433 );
xor ( n27613 , n27612 , n27436 );
and ( n27614 , n27610 , n27613 );
and ( n27615 , n27606 , n27613 );
or ( n27616 , n27611 , n27614 , n27615 );
and ( n27617 , n23351 , n21687 );
and ( n27618 , n23320 , n21685 );
nor ( n27619 , n27617 , n27618 );
xnor ( n27620 , n27619 , n21697 );
and ( n27621 , n27616 , n27620 );
and ( n27622 , n27592 , n27621 );
xor ( n27623 , n27451 , n27453 );
xor ( n27624 , n27623 , n27490 );
and ( n27625 , n27621 , n27624 );
and ( n27626 , n27592 , n27624 );
or ( n27627 , n27622 , n27625 , n27626 );
xor ( n27628 , n27340 , n27393 );
xor ( n27629 , n27628 , n27493 );
and ( n27630 , n27627 , n27629 );
and ( n27631 , n23320 , n21663 );
and ( n27632 , n23074 , n21661 );
nor ( n27633 , n27631 , n27632 );
xnor ( n27634 , n27633 , n21673 );
and ( n27635 , n23503 , n21687 );
and ( n27636 , n23351 , n21685 );
nor ( n27637 , n27635 , n27636 );
xnor ( n27638 , n27637 , n21697 );
and ( n27639 , n27634 , n27638 );
xor ( n27640 , n27606 , n27610 );
xor ( n27641 , n27640 , n27613 );
and ( n27642 , n27638 , n27641 );
and ( n27643 , n27634 , n27641 );
or ( n27644 , n27639 , n27642 , n27643 );
and ( n27645 , n21545 , n22114 );
and ( n27646 , n21486 , n22112 );
nor ( n27647 , n27645 , n27646 );
xnor ( n27648 , n27647 , n22124 );
and ( n27649 , n27644 , n27648 );
xor ( n27650 , n27480 , n27484 );
xor ( n27651 , n27650 , n27487 );
and ( n27652 , n27648 , n27651 );
and ( n27653 , n27644 , n27651 );
or ( n27654 , n27649 , n27652 , n27653 );
xor ( n27655 , n27370 , n27372 );
xor ( n27656 , n27655 , n27387 );
xor ( n27657 , n27616 , n27620 );
and ( n27658 , n27656 , n27657 );
and ( n27659 , n25343 , n21582 );
and ( n27660 , n25179 , n21580 );
nor ( n27661 , n27659 , n27660 );
xnor ( n27662 , n27661 , n21588 );
and ( n27663 , n25553 , n21783 );
and ( n27664 , n25544 , n21781 );
nor ( n27665 , n27663 , n27664 );
xnor ( n27666 , n27665 , n21793 );
and ( n27667 , n27662 , n27666 );
xor ( n27668 , n27528 , n27532 );
xor ( n27669 , n27668 , n27535 );
and ( n27670 , n27666 , n27669 );
and ( n27671 , n27662 , n27669 );
or ( n27672 , n27667 , n27670 , n27671 );
and ( n27673 , n24631 , n21236 );
and ( n27674 , n24460 , n21234 );
nor ( n27675 , n27673 , n27674 );
xnor ( n27676 , n27675 , n21246 );
and ( n27677 , n27672 , n27676 );
and ( n27678 , n24812 , n21260 );
and ( n27679 , n24662 , n21258 );
nor ( n27680 , n27678 , n27679 );
xnor ( n27681 , n27680 , n21270 );
and ( n27682 , n27676 , n27681 );
and ( n27683 , n27672 , n27681 );
or ( n27684 , n27677 , n27682 , n27683 );
and ( n27685 , n23949 , n21707 );
and ( n27686 , n23887 , n21705 );
nor ( n27687 , n27685 , n27686 );
xnor ( n27688 , n27687 , n21717 );
and ( n27689 , n27684 , n27688 );
xor ( n27690 , n27596 , n27600 );
xor ( n27691 , n27690 , n27603 );
and ( n27692 , n27688 , n27691 );
and ( n27693 , n27684 , n27691 );
or ( n27694 , n27689 , n27692 , n27693 );
and ( n27695 , n21606 , n21414 );
and ( n27696 , n21511 , n21412 );
nor ( n27697 , n27695 , n27696 );
xnor ( n27698 , n27697 , n21480 );
and ( n27699 , n27694 , n27698 );
and ( n27700 , n22813 , n21139 );
and ( n27701 , n21616 , n21137 );
nor ( n27702 , n27700 , n27701 );
xnor ( n27703 , n27702 , n21221 );
and ( n27704 , n27698 , n27703 );
and ( n27705 , n27694 , n27703 );
or ( n27706 , n27699 , n27704 , n27705 );
and ( n27707 , n27657 , n27706 );
and ( n27708 , n27656 , n27706 );
or ( n27709 , n27658 , n27707 , n27708 );
and ( n27710 , n27654 , n27709 );
xor ( n27711 , n27592 , n27621 );
xor ( n27712 , n27711 , n27624 );
and ( n27713 , n27709 , n27712 );
and ( n27714 , n27654 , n27712 );
or ( n27715 , n27710 , n27713 , n27714 );
and ( n27716 , n27629 , n27715 );
and ( n27717 , n27627 , n27715 );
or ( n27718 , n27630 , n27716 , n27717 );
and ( n27719 , n27503 , n27718 );
xor ( n27720 , n27503 , n27718 );
xor ( n27721 , n27627 , n27629 );
xor ( n27722 , n27721 , n27715 );
and ( n27723 , n23351 , n21663 );
and ( n27724 , n23320 , n21661 );
nor ( n27725 , n27723 , n27724 );
xnor ( n27726 , n27725 , n21673 );
and ( n27727 , n23651 , n21687 );
and ( n27728 , n23503 , n21685 );
nor ( n27729 , n27727 , n27728 );
xnor ( n27730 , n27729 , n21697 );
and ( n27731 , n27726 , n27730 );
xor ( n27732 , n27558 , n27562 );
xor ( n27733 , n27732 , n27567 );
and ( n27734 , n27730 , n27733 );
and ( n27735 , n27726 , n27733 );
or ( n27736 , n27731 , n27734 , n27735 );
and ( n27737 , n21486 , n22032 );
and ( n27738 , n21501 , n22029 );
nor ( n27739 , n27737 , n27738 );
xnor ( n27740 , n27739 , n22027 );
and ( n27741 , n27736 , n27740 );
xor ( n27742 , n27570 , n27574 );
xor ( n27743 , n27742 , n27577 );
and ( n27744 , n27740 , n27743 );
and ( n27745 , n27736 , n27743 );
or ( n27746 , n27741 , n27744 , n27745 );
and ( n27747 , n25544 , n21582 );
and ( n27748 , n25343 , n21580 );
nor ( n27749 , n27747 , n27748 );
xnor ( n27750 , n27749 , n21588 );
and ( n27751 , n25772 , n21783 );
and ( n27752 , n25553 , n21781 );
nor ( n27753 , n27751 , n27752 );
xnor ( n27754 , n27753 , n21793 );
and ( n27755 , n27750 , n27754 );
xor ( n27756 , n27504 , n27520 );
xor ( n27757 , n27756 , n27525 );
and ( n27758 , n27754 , n27757 );
and ( n27759 , n27750 , n27757 );
or ( n27760 , n27755 , n27758 , n27759 );
and ( n27761 , n25060 , n21260 );
and ( n27762 , n24812 , n21258 );
nor ( n27763 , n27761 , n27762 );
xnor ( n27764 , n27763 , n21270 );
and ( n27765 , n27760 , n27764 );
xor ( n27766 , n27662 , n27666 );
xor ( n27767 , n27766 , n27669 );
and ( n27768 , n27764 , n27767 );
and ( n27769 , n27760 , n27767 );
or ( n27770 , n27765 , n27768 , n27769 );
and ( n27771 , n24213 , n21707 );
and ( n27772 , n23949 , n21705 );
nor ( n27773 , n27771 , n27772 );
xnor ( n27774 , n27773 , n21717 );
and ( n27775 , n27770 , n27774 );
xor ( n27776 , n27538 , n27542 );
xor ( n27777 , n27776 , n27555 );
and ( n27778 , n27774 , n27777 );
and ( n27779 , n27770 , n27777 );
or ( n27780 , n27775 , n27778 , n27779 );
and ( n27781 , n23074 , n21139 );
and ( n27782 , n22813 , n21137 );
nor ( n27783 , n27781 , n27782 );
xnor ( n27784 , n27783 , n21221 );
and ( n27785 , n27780 , n27784 );
xor ( n27786 , n27684 , n27688 );
xor ( n27787 , n27786 , n27691 );
and ( n27788 , n27784 , n27787 );
and ( n27789 , n27780 , n27787 );
or ( n27790 , n27785 , n27788 , n27789 );
and ( n27791 , n21599 , n22114 );
and ( n27792 , n21545 , n22112 );
nor ( n27793 , n27791 , n27792 );
xnor ( n27794 , n27793 , n22124 );
and ( n27795 , n27790 , n27794 );
xor ( n27796 , n27634 , n27638 );
xor ( n27797 , n27796 , n27641 );
and ( n27798 , n27794 , n27797 );
and ( n27799 , n27790 , n27797 );
or ( n27800 , n27795 , n27798 , n27799 );
and ( n27801 , n27746 , n27800 );
xor ( n27802 , n27580 , n27584 );
xor ( n27803 , n27802 , n27589 );
and ( n27804 , n27800 , n27803 );
and ( n27805 , n27746 , n27803 );
or ( n27806 , n27801 , n27804 , n27805 );
xor ( n27807 , n27654 , n27709 );
xor ( n27808 , n27807 , n27712 );
and ( n27809 , n27806 , n27808 );
xor ( n27810 , n27644 , n27648 );
xor ( n27811 , n27810 , n27651 );
xor ( n27812 , n27656 , n27657 );
xor ( n27813 , n27812 , n27706 );
and ( n27814 , n27811 , n27813 );
xor ( n27815 , n27746 , n27800 );
xor ( n27816 , n27815 , n27803 );
and ( n27817 , n27813 , n27816 );
and ( n27818 , n27811 , n27816 );
or ( n27819 , n27814 , n27817 , n27818 );
and ( n27820 , n27808 , n27819 );
and ( n27821 , n27806 , n27819 );
or ( n27822 , n27809 , n27820 , n27821 );
and ( n27823 , n27722 , n27822 );
xor ( n27824 , n27722 , n27822 );
xor ( n27825 , n27507 , n27511 );
and ( n27826 , n26003 , n21781 );
not ( n27827 , n27826 );
and ( n27828 , n27827 , n21793 );
and ( n27829 , n26003 , n21783 );
and ( n27830 , n26011 , n21781 );
nor ( n27831 , n27829 , n27830 );
xnor ( n27832 , n27831 , n21793 );
and ( n27833 , n27828 , n27832 );
and ( n27834 , n26011 , n21783 );
and ( n27835 , n26020 , n21781 );
nor ( n27836 , n27834 , n27835 );
xnor ( n27837 , n27836 , n21793 );
and ( n27838 , n27833 , n27837 );
and ( n27839 , n27837 , n27505 );
and ( n27840 , n27833 , n27505 );
or ( n27841 , n27838 , n27839 , n27840 );
and ( n27842 , n27825 , n27841 );
and ( n27843 , n26020 , n21783 );
and ( n27844 , n25898 , n21781 );
nor ( n27845 , n27843 , n27844 );
xnor ( n27846 , n27845 , n21793 );
and ( n27847 , n27841 , n27846 );
and ( n27848 , n27825 , n27846 );
or ( n27849 , n27842 , n27847 , n27848 );
and ( n27850 , n25898 , n21783 );
and ( n27851 , n25772 , n21781 );
nor ( n27852 , n27850 , n27851 );
xnor ( n27853 , n27852 , n21793 );
and ( n27854 , n27849 , n27853 );
xor ( n27855 , n27512 , n27516 );
xor ( n27856 , n27855 , n27396 );
and ( n27857 , n27853 , n27856 );
and ( n27858 , n27849 , n27856 );
or ( n27859 , n27854 , n27857 , n27858 );
and ( n27860 , n25179 , n21260 );
and ( n27861 , n25060 , n21258 );
nor ( n27862 , n27860 , n27861 );
xnor ( n27863 , n27862 , n21270 );
and ( n27864 , n27859 , n27863 );
xor ( n27865 , n27750 , n27754 );
xor ( n27866 , n27865 , n27757 );
and ( n27867 , n27863 , n27866 );
and ( n27868 , n27859 , n27866 );
or ( n27869 , n27864 , n27867 , n27868 );
and ( n27870 , n24460 , n21707 );
and ( n27871 , n24213 , n21705 );
nor ( n27872 , n27870 , n27871 );
xnor ( n27873 , n27872 , n21717 );
and ( n27874 , n27869 , n27873 );
and ( n27875 , n24662 , n21236 );
and ( n27876 , n24631 , n21234 );
nor ( n27877 , n27875 , n27876 );
xnor ( n27878 , n27877 , n21246 );
and ( n27879 , n27873 , n27878 );
and ( n27880 , n27869 , n27878 );
or ( n27881 , n27874 , n27879 , n27880 );
and ( n27882 , n23887 , n21687 );
and ( n27883 , n23651 , n21685 );
nor ( n27884 , n27882 , n27883 );
xnor ( n27885 , n27884 , n21697 );
and ( n27886 , n27881 , n27885 );
xor ( n27887 , n27672 , n27676 );
xor ( n27888 , n27887 , n27681 );
and ( n27889 , n27885 , n27888 );
and ( n27890 , n27881 , n27888 );
or ( n27891 , n27886 , n27889 , n27890 );
and ( n27892 , n21511 , n22114 );
and ( n27893 , n21599 , n22112 );
nor ( n27894 , n27892 , n27893 );
xnor ( n27895 , n27894 , n22124 );
and ( n27896 , n27891 , n27895 );
and ( n27897 , n21616 , n21414 );
and ( n27898 , n21606 , n21412 );
nor ( n27899 , n27897 , n27898 );
xnor ( n27900 , n27899 , n21480 );
and ( n27901 , n27895 , n27900 );
and ( n27902 , n27891 , n27900 );
or ( n27903 , n27896 , n27901 , n27902 );
and ( n27904 , n23320 , n21139 );
and ( n27905 , n23074 , n21137 );
nor ( n27906 , n27904 , n27905 );
xnor ( n27907 , n27906 , n21221 );
and ( n27908 , n23503 , n21663 );
and ( n27909 , n23351 , n21661 );
nor ( n27910 , n27908 , n27909 );
xnor ( n27911 , n27910 , n21673 );
and ( n27912 , n27907 , n27911 );
xor ( n27913 , n27770 , n27774 );
xor ( n27914 , n27913 , n27777 );
and ( n27915 , n27911 , n27914 );
and ( n27916 , n27907 , n27914 );
or ( n27917 , n27912 , n27915 , n27916 );
and ( n27918 , n21545 , n22032 );
and ( n27919 , n21486 , n22029 );
nor ( n27920 , n27918 , n27919 );
xnor ( n27921 , n27920 , n22027 );
and ( n27922 , n27917 , n27921 );
xor ( n27923 , n27726 , n27730 );
xor ( n27924 , n27923 , n27733 );
and ( n27925 , n27921 , n27924 );
and ( n27926 , n27917 , n27924 );
or ( n27927 , n27922 , n27925 , n27926 );
and ( n27928 , n27903 , n27927 );
xor ( n27929 , n27694 , n27698 );
xor ( n27930 , n27929 , n27703 );
and ( n27931 , n27927 , n27930 );
and ( n27932 , n27903 , n27930 );
or ( n27933 , n27928 , n27931 , n27932 );
and ( n27934 , n25343 , n21260 );
and ( n27935 , n25179 , n21258 );
nor ( n27936 , n27934 , n27935 );
xnor ( n27937 , n27936 , n21270 );
and ( n27938 , n25553 , n21582 );
and ( n27939 , n25544 , n21580 );
nor ( n27940 , n27938 , n27939 );
xnor ( n27941 , n27940 , n21588 );
and ( n27942 , n27937 , n27941 );
xor ( n27943 , n27849 , n27853 );
xor ( n27944 , n27943 , n27856 );
and ( n27945 , n27941 , n27944 );
and ( n27946 , n27937 , n27944 );
or ( n27947 , n27942 , n27945 , n27946 );
and ( n27948 , n24812 , n21236 );
and ( n27949 , n24662 , n21234 );
nor ( n27950 , n27948 , n27949 );
xnor ( n27951 , n27950 , n21246 );
and ( n27952 , n27947 , n27951 );
xor ( n27953 , n27859 , n27863 );
xor ( n27954 , n27953 , n27866 );
and ( n27955 , n27951 , n27954 );
and ( n27956 , n27947 , n27954 );
or ( n27957 , n27952 , n27955 , n27956 );
and ( n27958 , n23949 , n21687 );
and ( n27959 , n23887 , n21685 );
nor ( n27960 , n27958 , n27959 );
xnor ( n27961 , n27960 , n21697 );
and ( n27962 , n27957 , n27961 );
xor ( n27963 , n27760 , n27764 );
xor ( n27964 , n27963 , n27767 );
and ( n27965 , n27961 , n27964 );
and ( n27966 , n27957 , n27964 );
or ( n27967 , n27962 , n27965 , n27966 );
and ( n27968 , n21606 , n22114 );
and ( n27969 , n21511 , n22112 );
nor ( n27970 , n27968 , n27969 );
xnor ( n27971 , n27970 , n22124 );
and ( n27972 , n27967 , n27971 );
and ( n27973 , n22813 , n21414 );
and ( n27974 , n21616 , n21412 );
nor ( n27975 , n27973 , n27974 );
xnor ( n27976 , n27975 , n21480 );
and ( n27977 , n27971 , n27976 );
and ( n27978 , n27967 , n27976 );
or ( n27979 , n27972 , n27977 , n27978 );
xor ( n27980 , n27891 , n27895 );
xor ( n27981 , n27980 , n27900 );
and ( n27982 , n27979 , n27981 );
xor ( n27983 , n27780 , n27784 );
xor ( n27984 , n27983 , n27787 );
and ( n27985 , n27981 , n27984 );
and ( n27986 , n27979 , n27984 );
or ( n27987 , n27982 , n27985 , n27986 );
xor ( n27988 , n27736 , n27740 );
xor ( n27989 , n27988 , n27743 );
and ( n27990 , n27987 , n27989 );
xor ( n27991 , n27790 , n27794 );
xor ( n27992 , n27991 , n27797 );
and ( n27993 , n27989 , n27992 );
and ( n27994 , n27987 , n27992 );
or ( n27995 , n27990 , n27993 , n27994 );
and ( n27996 , n27933 , n27995 );
and ( n27997 , n23074 , n21414 );
and ( n27998 , n22813 , n21412 );
nor ( n27999 , n27997 , n27998 );
xnor ( n28000 , n27999 , n21480 );
and ( n28001 , n23651 , n21663 );
and ( n28002 , n23503 , n21661 );
nor ( n28003 , n28001 , n28002 );
xnor ( n28004 , n28003 , n21673 );
and ( n28005 , n28000 , n28004 );
xor ( n28006 , n27869 , n27873 );
xor ( n28007 , n28006 , n27878 );
and ( n28008 , n28004 , n28007 );
and ( n28009 , n28000 , n28007 );
or ( n28010 , n28005 , n28008 , n28009 );
and ( n28011 , n21599 , n22032 );
and ( n28012 , n21545 , n22029 );
nor ( n28013 , n28011 , n28012 );
xnor ( n28014 , n28013 , n22027 );
and ( n28015 , n28010 , n28014 );
xor ( n28016 , n27881 , n27885 );
xor ( n28017 , n28016 , n27888 );
and ( n28018 , n28014 , n28017 );
and ( n28019 , n28010 , n28017 );
or ( n28020 , n28015 , n28018 , n28019 );
and ( n28021 , n25544 , n21260 );
and ( n28022 , n25343 , n21258 );
nor ( n28023 , n28021 , n28022 );
xnor ( n28024 , n28023 , n21270 );
and ( n28025 , n25772 , n21582 );
and ( n28026 , n25553 , n21580 );
nor ( n28027 , n28025 , n28026 );
xnor ( n28028 , n28027 , n21588 );
and ( n28029 , n28024 , n28028 );
xor ( n28030 , n27825 , n27841 );
xor ( n28031 , n28030 , n27846 );
and ( n28032 , n28028 , n28031 );
and ( n28033 , n28024 , n28031 );
or ( n28034 , n28029 , n28032 , n28033 );
and ( n28035 , n25060 , n21236 );
and ( n28036 , n24812 , n21234 );
nor ( n28037 , n28035 , n28036 );
xnor ( n28038 , n28037 , n21246 );
and ( n28039 , n28034 , n28038 );
xor ( n28040 , n27937 , n27941 );
xor ( n28041 , n28040 , n27944 );
and ( n28042 , n28038 , n28041 );
and ( n28043 , n28034 , n28041 );
or ( n28044 , n28039 , n28042 , n28043 );
and ( n28045 , n24213 , n21687 );
and ( n28046 , n23949 , n21685 );
nor ( n28047 , n28045 , n28046 );
xnor ( n28048 , n28047 , n21697 );
and ( n28049 , n28044 , n28048 );
and ( n28050 , n24631 , n21707 );
and ( n28051 , n24460 , n21705 );
nor ( n28052 , n28050 , n28051 );
xnor ( n28053 , n28052 , n21717 );
and ( n28054 , n28048 , n28053 );
and ( n28055 , n28044 , n28053 );
or ( n28056 , n28049 , n28054 , n28055 );
and ( n28057 , n21616 , n22114 );
and ( n28058 , n21606 , n22112 );
nor ( n28059 , n28057 , n28058 );
xnor ( n28060 , n28059 , n22124 );
and ( n28061 , n28056 , n28060 );
and ( n28062 , n23351 , n21139 );
and ( n28063 , n23320 , n21137 );
nor ( n28064 , n28062 , n28063 );
xnor ( n28065 , n28064 , n21221 );
and ( n28066 , n28060 , n28065 );
and ( n28067 , n28056 , n28065 );
or ( n28068 , n28061 , n28066 , n28067 );
xor ( n28069 , n27828 , n27832 );
and ( n28070 , n26003 , n21580 );
not ( n28071 , n28070 );
and ( n28072 , n28071 , n21588 );
and ( n28073 , n26003 , n21582 );
and ( n28074 , n26011 , n21580 );
nor ( n28075 , n28073 , n28074 );
xnor ( n28076 , n28075 , n21588 );
and ( n28077 , n28072 , n28076 );
and ( n28078 , n26011 , n21582 );
and ( n28079 , n26020 , n21580 );
nor ( n28080 , n28078 , n28079 );
xnor ( n28081 , n28080 , n21588 );
and ( n28082 , n28077 , n28081 );
and ( n28083 , n28081 , n27826 );
and ( n28084 , n28077 , n27826 );
or ( n28085 , n28082 , n28083 , n28084 );
and ( n28086 , n28069 , n28085 );
and ( n28087 , n26020 , n21582 );
and ( n28088 , n25898 , n21580 );
nor ( n28089 , n28087 , n28088 );
xnor ( n28090 , n28089 , n21588 );
and ( n28091 , n28085 , n28090 );
and ( n28092 , n28069 , n28090 );
or ( n28093 , n28086 , n28091 , n28092 );
and ( n28094 , n25898 , n21582 );
and ( n28095 , n25772 , n21580 );
nor ( n28096 , n28094 , n28095 );
xnor ( n28097 , n28096 , n21588 );
and ( n28098 , n28093 , n28097 );
xor ( n28099 , n27833 , n27837 );
xor ( n28100 , n28099 , n27505 );
and ( n28101 , n28097 , n28100 );
and ( n28102 , n28093 , n28100 );
or ( n28103 , n28098 , n28101 , n28102 );
and ( n28104 , n25179 , n21236 );
and ( n28105 , n25060 , n21234 );
nor ( n28106 , n28104 , n28105 );
xnor ( n28107 , n28106 , n21246 );
and ( n28108 , n28103 , n28107 );
xor ( n28109 , n28024 , n28028 );
xor ( n28110 , n28109 , n28031 );
and ( n28111 , n28107 , n28110 );
and ( n28112 , n28103 , n28110 );
or ( n28113 , n28108 , n28111 , n28112 );
and ( n28114 , n24460 , n21687 );
and ( n28115 , n24213 , n21685 );
nor ( n28116 , n28114 , n28115 );
xnor ( n28117 , n28116 , n21697 );
and ( n28118 , n28113 , n28117 );
and ( n28119 , n24662 , n21707 );
and ( n28120 , n24631 , n21705 );
nor ( n28121 , n28119 , n28120 );
xnor ( n28122 , n28121 , n21717 );
and ( n28123 , n28117 , n28122 );
and ( n28124 , n28113 , n28122 );
or ( n28125 , n28118 , n28123 , n28124 );
and ( n28126 , n23887 , n21663 );
and ( n28127 , n23651 , n21661 );
nor ( n28128 , n28126 , n28127 );
xnor ( n28129 , n28128 , n21673 );
and ( n28130 , n28125 , n28129 );
xor ( n28131 , n27947 , n27951 );
xor ( n28132 , n28131 , n27954 );
and ( n28133 , n28129 , n28132 );
and ( n28134 , n28125 , n28132 );
or ( n28135 , n28130 , n28133 , n28134 );
and ( n28136 , n21511 , n22032 );
and ( n28137 , n21599 , n22029 );
nor ( n28138 , n28136 , n28137 );
xnor ( n28139 , n28138 , n22027 );
and ( n28140 , n28135 , n28139 );
xor ( n28141 , n27957 , n27961 );
xor ( n28142 , n28141 , n27964 );
and ( n28143 , n28139 , n28142 );
and ( n28144 , n28135 , n28142 );
or ( n28145 , n28140 , n28143 , n28144 );
and ( n28146 , n28068 , n28145 );
xor ( n28147 , n27907 , n27911 );
xor ( n28148 , n28147 , n27914 );
and ( n28149 , n28145 , n28148 );
and ( n28150 , n28068 , n28148 );
or ( n28151 , n28146 , n28149 , n28150 );
and ( n28152 , n28020 , n28151 );
xor ( n28153 , n27917 , n27921 );
xor ( n28154 , n28153 , n27924 );
and ( n28155 , n28151 , n28154 );
and ( n28156 , n28020 , n28154 );
or ( n28157 , n28152 , n28155 , n28156 );
xor ( n28158 , n27903 , n27927 );
xor ( n28159 , n28158 , n27930 );
and ( n28160 , n28157 , n28159 );
xor ( n28161 , n27987 , n27989 );
xor ( n28162 , n28161 , n27992 );
and ( n28163 , n28159 , n28162 );
and ( n28164 , n28157 , n28162 );
or ( n28165 , n28160 , n28163 , n28164 );
and ( n28166 , n27995 , n28165 );
and ( n28167 , n27933 , n28165 );
or ( n28168 , n27996 , n28166 , n28167 );
xor ( n28169 , n27806 , n27808 );
xor ( n28170 , n28169 , n27819 );
and ( n28171 , n28168 , n28170 );
xor ( n28172 , n28168 , n28170 );
xor ( n28173 , n27811 , n27813 );
xor ( n28174 , n28173 , n27816 );
xor ( n28175 , n27933 , n27995 );
xor ( n28176 , n28175 , n28165 );
and ( n28177 , n28174 , n28176 );
xor ( n28178 , n28174 , n28176 );
xor ( n28179 , n28157 , n28159 );
xor ( n28180 , n28179 , n28162 );
and ( n28181 , n23651 , n21139 );
and ( n28182 , n23503 , n21137 );
nor ( n28183 , n28181 , n28182 );
xnor ( n28184 , n28183 , n21221 );
and ( n28185 , n23949 , n21663 );
and ( n28186 , n23887 , n21661 );
nor ( n28187 , n28185 , n28186 );
xnor ( n28188 , n28187 , n21673 );
and ( n28189 , n28184 , n28188 );
xor ( n28190 , n28034 , n28038 );
xor ( n28191 , n28190 , n28041 );
and ( n28192 , n28188 , n28191 );
and ( n28193 , n28184 , n28191 );
or ( n28194 , n28189 , n28192 , n28193 );
and ( n28195 , n21606 , n22032 );
and ( n28196 , n21511 , n22029 );
nor ( n28197 , n28195 , n28196 );
xnor ( n28198 , n28197 , n22027 );
and ( n28199 , n28194 , n28198 );
and ( n28200 , n22813 , n22114 );
and ( n28201 , n21616 , n22112 );
nor ( n28202 , n28200 , n28201 );
xnor ( n28203 , n28202 , n22124 );
and ( n28204 , n28198 , n28203 );
and ( n28205 , n28194 , n28203 );
or ( n28206 , n28199 , n28204 , n28205 );
and ( n28207 , n23320 , n21414 );
and ( n28208 , n23074 , n21412 );
nor ( n28209 , n28207 , n28208 );
xnor ( n28210 , n28209 , n21480 );
and ( n28211 , n23503 , n21139 );
and ( n28212 , n23351 , n21137 );
nor ( n28213 , n28211 , n28212 );
xnor ( n28214 , n28213 , n21221 );
and ( n28215 , n28210 , n28214 );
xor ( n28216 , n28044 , n28048 );
xor ( n28217 , n28216 , n28053 );
and ( n28218 , n28214 , n28217 );
and ( n28219 , n28210 , n28217 );
or ( n28220 , n28215 , n28218 , n28219 );
and ( n28221 , n28206 , n28220 );
xor ( n28222 , n28000 , n28004 );
xor ( n28223 , n28222 , n28007 );
and ( n28224 , n28220 , n28223 );
and ( n28225 , n28206 , n28223 );
or ( n28226 , n28221 , n28224 , n28225 );
xor ( n28227 , n27967 , n27971 );
xor ( n28228 , n28227 , n27976 );
and ( n28229 , n28226 , n28228 );
xor ( n28230 , n28010 , n28014 );
xor ( n28231 , n28230 , n28017 );
and ( n28232 , n28228 , n28231 );
and ( n28233 , n28226 , n28231 );
or ( n28234 , n28229 , n28232 , n28233 );
xor ( n28235 , n28020 , n28151 );
xor ( n28236 , n28235 , n28154 );
and ( n28237 , n28234 , n28236 );
xor ( n28238 , n27979 , n27981 );
xor ( n28239 , n28238 , n27984 );
and ( n28240 , n28236 , n28239 );
and ( n28241 , n28234 , n28239 );
or ( n28242 , n28237 , n28240 , n28241 );
and ( n28243 , n28180 , n28242 );
xor ( n28244 , n28180 , n28242 );
xor ( n28245 , n28234 , n28236 );
xor ( n28246 , n28245 , n28239 );
and ( n28247 , n25343 , n21236 );
and ( n28248 , n25179 , n21234 );
nor ( n28249 , n28247 , n28248 );
xnor ( n28250 , n28249 , n21246 );
and ( n28251 , n25553 , n21260 );
and ( n28252 , n25544 , n21258 );
nor ( n28253 , n28251 , n28252 );
xnor ( n28254 , n28253 , n21270 );
and ( n28255 , n28250 , n28254 );
xor ( n28256 , n28093 , n28097 );
xor ( n28257 , n28256 , n28100 );
and ( n28258 , n28254 , n28257 );
and ( n28259 , n28250 , n28257 );
or ( n28260 , n28255 , n28258 , n28259 );
and ( n28261 , n24631 , n21687 );
and ( n28262 , n24460 , n21685 );
nor ( n28263 , n28261 , n28262 );
xnor ( n28264 , n28263 , n21697 );
and ( n28265 , n28260 , n28264 );
xor ( n28266 , n28103 , n28107 );
xor ( n28267 , n28266 , n28110 );
and ( n28268 , n28264 , n28267 );
and ( n28269 , n28260 , n28267 );
or ( n28270 , n28265 , n28268 , n28269 );
and ( n28271 , n23074 , n22114 );
and ( n28272 , n22813 , n22112 );
nor ( n28273 , n28271 , n28272 );
xnor ( n28274 , n28273 , n22124 );
and ( n28275 , n28270 , n28274 );
and ( n28276 , n23351 , n21414 );
and ( n28277 , n23320 , n21412 );
nor ( n28278 , n28276 , n28277 );
xnor ( n28279 , n28278 , n21480 );
and ( n28280 , n28274 , n28279 );
and ( n28281 , n28270 , n28279 );
or ( n28282 , n28275 , n28280 , n28281 );
xor ( n28283 , n28210 , n28214 );
xor ( n28284 , n28283 , n28217 );
and ( n28285 , n28282 , n28284 );
xor ( n28286 , n28125 , n28129 );
xor ( n28287 , n28286 , n28132 );
and ( n28288 , n28284 , n28287 );
and ( n28289 , n28282 , n28287 );
or ( n28290 , n28285 , n28288 , n28289 );
xor ( n28291 , n28056 , n28060 );
xor ( n28292 , n28291 , n28065 );
and ( n28293 , n28290 , n28292 );
xor ( n28294 , n28135 , n28139 );
xor ( n28295 , n28294 , n28142 );
and ( n28296 , n28292 , n28295 );
and ( n28297 , n28290 , n28295 );
or ( n28298 , n28293 , n28296 , n28297 );
xor ( n28299 , n28226 , n28228 );
xor ( n28300 , n28299 , n28231 );
and ( n28301 , n28298 , n28300 );
xor ( n28302 , n28068 , n28145 );
xor ( n28303 , n28302 , n28148 );
and ( n28304 , n28300 , n28303 );
and ( n28305 , n28298 , n28303 );
or ( n28306 , n28301 , n28304 , n28305 );
and ( n28307 , n28246 , n28306 );
xor ( n28308 , n28246 , n28306 );
xor ( n28309 , n28298 , n28300 );
xor ( n28310 , n28309 , n28303 );
and ( n28311 , n25544 , n21236 );
and ( n28312 , n25343 , n21234 );
nor ( n28313 , n28311 , n28312 );
xnor ( n28314 , n28313 , n21246 );
and ( n28315 , n25772 , n21260 );
and ( n28316 , n25553 , n21258 );
nor ( n28317 , n28315 , n28316 );
xnor ( n28318 , n28317 , n21270 );
and ( n28319 , n28314 , n28318 );
xor ( n28320 , n28069 , n28085 );
xor ( n28321 , n28320 , n28090 );
and ( n28322 , n28318 , n28321 );
and ( n28323 , n28314 , n28321 );
or ( n28324 , n28319 , n28322 , n28323 );
and ( n28325 , n25060 , n21707 );
and ( n28326 , n24812 , n21705 );
nor ( n28327 , n28325 , n28326 );
xnor ( n28328 , n28327 , n21717 );
and ( n28329 , n28324 , n28328 );
xor ( n28330 , n28250 , n28254 );
xor ( n28331 , n28330 , n28257 );
and ( n28332 , n28328 , n28331 );
and ( n28333 , n28324 , n28331 );
or ( n28334 , n28329 , n28332 , n28333 );
and ( n28335 , n24213 , n21663 );
and ( n28336 , n23949 , n21661 );
nor ( n28337 , n28335 , n28336 );
xnor ( n28338 , n28337 , n21673 );
and ( n28339 , n28334 , n28338 );
and ( n28340 , n24812 , n21707 );
and ( n28341 , n24662 , n21705 );
nor ( n28342 , n28340 , n28341 );
xnor ( n28343 , n28342 , n21717 );
and ( n28344 , n28338 , n28343 );
and ( n28345 , n28334 , n28343 );
or ( n28346 , n28339 , n28344 , n28345 );
and ( n28347 , n21616 , n22032 );
and ( n28348 , n21606 , n22029 );
nor ( n28349 , n28347 , n28348 );
xnor ( n28350 , n28349 , n22027 );
and ( n28351 , n28346 , n28350 );
xor ( n28352 , n28113 , n28117 );
xor ( n28353 , n28352 , n28122 );
and ( n28354 , n28350 , n28353 );
and ( n28355 , n28346 , n28353 );
or ( n28356 , n28351 , n28354 , n28355 );
xor ( n28357 , n28072 , n28076 );
and ( n28358 , n26003 , n21258 );
not ( n28359 , n28358 );
and ( n28360 , n28359 , n21270 );
and ( n28361 , n26003 , n21260 );
and ( n28362 , n26011 , n21258 );
nor ( n28363 , n28361 , n28362 );
xnor ( n28364 , n28363 , n21270 );
and ( n28365 , n28360 , n28364 );
and ( n28366 , n26011 , n21260 );
and ( n28367 , n26020 , n21258 );
nor ( n28368 , n28366 , n28367 );
xnor ( n28369 , n28368 , n21270 );
and ( n28370 , n28365 , n28369 );
and ( n28371 , n28369 , n28070 );
and ( n28372 , n28365 , n28070 );
or ( n28373 , n28370 , n28371 , n28372 );
and ( n28374 , n28357 , n28373 );
and ( n28375 , n26020 , n21260 );
and ( n28376 , n25898 , n21258 );
nor ( n28377 , n28375 , n28376 );
xnor ( n28378 , n28377 , n21270 );
and ( n28379 , n28373 , n28378 );
and ( n28380 , n28357 , n28378 );
or ( n28381 , n28374 , n28379 , n28380 );
and ( n28382 , n25898 , n21260 );
and ( n28383 , n25772 , n21258 );
nor ( n28384 , n28382 , n28383 );
xnor ( n28385 , n28384 , n21270 );
and ( n28386 , n28381 , n28385 );
xor ( n28387 , n28077 , n28081 );
xor ( n28388 , n28387 , n27826 );
and ( n28389 , n28385 , n28388 );
and ( n28390 , n28381 , n28388 );
or ( n28391 , n28386 , n28389 , n28390 );
and ( n28392 , n25179 , n21707 );
and ( n28393 , n25060 , n21705 );
nor ( n28394 , n28392 , n28393 );
xnor ( n28395 , n28394 , n21717 );
and ( n28396 , n28391 , n28395 );
xor ( n28397 , n28314 , n28318 );
xor ( n28398 , n28397 , n28321 );
and ( n28399 , n28395 , n28398 );
and ( n28400 , n28391 , n28398 );
or ( n28401 , n28396 , n28399 , n28400 );
and ( n28402 , n24460 , n21663 );
and ( n28403 , n24213 , n21661 );
nor ( n28404 , n28402 , n28403 );
xnor ( n28405 , n28404 , n21673 );
and ( n28406 , n28401 , n28405 );
and ( n28407 , n24662 , n21687 );
and ( n28408 , n24631 , n21685 );
nor ( n28409 , n28407 , n28408 );
xnor ( n28410 , n28409 , n21697 );
and ( n28411 , n28405 , n28410 );
and ( n28412 , n28401 , n28410 );
or ( n28413 , n28406 , n28411 , n28412 );
and ( n28414 , n23320 , n22114 );
and ( n28415 , n23074 , n22112 );
nor ( n28416 , n28414 , n28415 );
xnor ( n28417 , n28416 , n22124 );
and ( n28418 , n28413 , n28417 );
and ( n28419 , n23887 , n21139 );
and ( n28420 , n23651 , n21137 );
nor ( n28421 , n28419 , n28420 );
xnor ( n28422 , n28421 , n21221 );
and ( n28423 , n28417 , n28422 );
and ( n28424 , n28413 , n28422 );
or ( n28425 , n28418 , n28423 , n28424 );
xor ( n28426 , n28270 , n28274 );
xor ( n28427 , n28426 , n28279 );
and ( n28428 , n28425 , n28427 );
xor ( n28429 , n28184 , n28188 );
xor ( n28430 , n28429 , n28191 );
and ( n28431 , n28427 , n28430 );
and ( n28432 , n28425 , n28430 );
or ( n28433 , n28428 , n28431 , n28432 );
and ( n28434 , n28356 , n28433 );
xor ( n28435 , n28194 , n28198 );
xor ( n28436 , n28435 , n28203 );
and ( n28437 , n28433 , n28436 );
and ( n28438 , n28356 , n28436 );
or ( n28439 , n28434 , n28437 , n28438 );
xor ( n28440 , n28206 , n28220 );
xor ( n28441 , n28440 , n28223 );
and ( n28442 , n28439 , n28441 );
xor ( n28443 , n28290 , n28292 );
xor ( n28444 , n28443 , n28295 );
and ( n28445 , n28441 , n28444 );
and ( n28446 , n28439 , n28444 );
or ( n28447 , n28442 , n28445 , n28446 );
and ( n28448 , n28310 , n28447 );
xor ( n28449 , n28310 , n28447 );
and ( n28450 , n23074 , n22032 );
and ( n28451 , n22813 , n22029 );
nor ( n28452 , n28450 , n28451 );
xnor ( n28453 , n28452 , n22027 );
and ( n28454 , n23651 , n21414 );
and ( n28455 , n23503 , n21412 );
nor ( n28456 , n28454 , n28455 );
xnor ( n28457 , n28456 , n21480 );
and ( n28458 , n28453 , n28457 );
xor ( n28459 , n28401 , n28405 );
xor ( n28460 , n28459 , n28410 );
and ( n28461 , n28457 , n28460 );
and ( n28462 , n28453 , n28460 );
or ( n28463 , n28458 , n28461 , n28462 );
and ( n28464 , n25343 , n21707 );
and ( n28465 , n25179 , n21705 );
nor ( n28466 , n28464 , n28465 );
xnor ( n28467 , n28466 , n21717 );
and ( n28468 , n25553 , n21236 );
and ( n28469 , n25544 , n21234 );
nor ( n28470 , n28468 , n28469 );
xnor ( n28471 , n28470 , n21246 );
and ( n28472 , n28467 , n28471 );
xor ( n28473 , n28381 , n28385 );
xor ( n28474 , n28473 , n28388 );
and ( n28475 , n28471 , n28474 );
and ( n28476 , n28467 , n28474 );
or ( n28477 , n28472 , n28475 , n28476 );
and ( n28478 , n24631 , n21663 );
and ( n28479 , n24460 , n21661 );
nor ( n28480 , n28478 , n28479 );
xnor ( n28481 , n28480 , n21673 );
and ( n28482 , n28477 , n28481 );
xor ( n28483 , n28391 , n28395 );
xor ( n28484 , n28483 , n28398 );
and ( n28485 , n28481 , n28484 );
and ( n28486 , n28477 , n28484 );
or ( n28487 , n28482 , n28485 , n28486 );
and ( n28488 , n23949 , n21139 );
and ( n28489 , n23887 , n21137 );
nor ( n28490 , n28488 , n28489 );
xnor ( n28491 , n28490 , n21221 );
and ( n28492 , n28487 , n28491 );
xor ( n28493 , n28324 , n28328 );
xor ( n28494 , n28493 , n28331 );
and ( n28495 , n28491 , n28494 );
and ( n28496 , n28487 , n28494 );
or ( n28497 , n28492 , n28495 , n28496 );
and ( n28498 , n28463 , n28497 );
and ( n28499 , n22813 , n22032 );
and ( n28500 , n21616 , n22029 );
nor ( n28501 , n28499 , n28500 );
xnor ( n28502 , n28501 , n22027 );
and ( n28503 , n28497 , n28502 );
and ( n28504 , n28463 , n28502 );
or ( n28505 , n28498 , n28503 , n28504 );
and ( n28506 , n23503 , n21414 );
and ( n28507 , n23351 , n21412 );
nor ( n28508 , n28506 , n28507 );
xnor ( n28509 , n28508 , n21480 );
xor ( n28510 , n28334 , n28338 );
xor ( n28511 , n28510 , n28343 );
and ( n28512 , n28509 , n28511 );
xor ( n28513 , n28260 , n28264 );
xor ( n28514 , n28513 , n28267 );
and ( n28515 , n28511 , n28514 );
and ( n28516 , n28509 , n28514 );
or ( n28517 , n28512 , n28515 , n28516 );
and ( n28518 , n28505 , n28517 );
xor ( n28519 , n28346 , n28350 );
xor ( n28520 , n28519 , n28353 );
and ( n28521 , n28517 , n28520 );
and ( n28522 , n28505 , n28520 );
or ( n28523 , n28518 , n28521 , n28522 );
xor ( n28524 , n28356 , n28433 );
xor ( n28525 , n28524 , n28436 );
and ( n28526 , n28523 , n28525 );
xor ( n28527 , n28282 , n28284 );
xor ( n28528 , n28527 , n28287 );
and ( n28529 , n28525 , n28528 );
and ( n28530 , n28523 , n28528 );
or ( n28531 , n28526 , n28529 , n28530 );
xor ( n28532 , n28439 , n28441 );
xor ( n28533 , n28532 , n28444 );
and ( n28534 , n28531 , n28533 );
xor ( n28535 , n28531 , n28533 );
xor ( n28536 , n28523 , n28525 );
xor ( n28537 , n28536 , n28528 );
and ( n28538 , n25544 , n21707 );
and ( n28539 , n25343 , n21705 );
nor ( n28540 , n28538 , n28539 );
xnor ( n28541 , n28540 , n21717 );
and ( n28542 , n25772 , n21236 );
and ( n28543 , n25553 , n21234 );
nor ( n28544 , n28542 , n28543 );
xnor ( n28545 , n28544 , n21246 );
and ( n28546 , n28541 , n28545 );
xor ( n28547 , n28357 , n28373 );
xor ( n28548 , n28547 , n28378 );
and ( n28549 , n28545 , n28548 );
and ( n28550 , n28541 , n28548 );
or ( n28551 , n28546 , n28549 , n28550 );
and ( n28552 , n25060 , n21687 );
and ( n28553 , n24812 , n21685 );
nor ( n28554 , n28552 , n28553 );
xnor ( n28555 , n28554 , n21697 );
and ( n28556 , n28551 , n28555 );
xor ( n28557 , n28467 , n28471 );
xor ( n28558 , n28557 , n28474 );
and ( n28559 , n28555 , n28558 );
and ( n28560 , n28551 , n28558 );
or ( n28561 , n28556 , n28559 , n28560 );
and ( n28562 , n24213 , n21139 );
and ( n28563 , n23949 , n21137 );
nor ( n28564 , n28562 , n28563 );
xnor ( n28565 , n28564 , n21221 );
and ( n28566 , n28561 , n28565 );
and ( n28567 , n24812 , n21687 );
and ( n28568 , n24662 , n21685 );
nor ( n28569 , n28567 , n28568 );
xnor ( n28570 , n28569 , n21697 );
and ( n28571 , n28565 , n28570 );
and ( n28572 , n28561 , n28570 );
or ( n28573 , n28566 , n28571 , n28572 );
and ( n28574 , n23351 , n22114 );
and ( n28575 , n23320 , n22112 );
nor ( n28576 , n28574 , n28575 );
xnor ( n28577 , n28576 , n22124 );
and ( n28578 , n28573 , n28577 );
xor ( n28579 , n28487 , n28491 );
xor ( n28580 , n28579 , n28494 );
and ( n28581 , n28577 , n28580 );
and ( n28582 , n28573 , n28580 );
or ( n28583 , n28578 , n28581 , n28582 );
xor ( n28584 , n28413 , n28417 );
xor ( n28585 , n28584 , n28422 );
and ( n28586 , n28583 , n28585 );
xor ( n28587 , n28509 , n28511 );
xor ( n28588 , n28587 , n28514 );
and ( n28589 , n28585 , n28588 );
and ( n28590 , n28583 , n28588 );
or ( n28591 , n28586 , n28589 , n28590 );
xor ( n28592 , n28505 , n28517 );
xor ( n28593 , n28592 , n28520 );
and ( n28594 , n28591 , n28593 );
xor ( n28595 , n28425 , n28427 );
xor ( n28596 , n28595 , n28430 );
and ( n28597 , n28593 , n28596 );
and ( n28598 , n28591 , n28596 );
or ( n28599 , n28594 , n28597 , n28598 );
and ( n28600 , n28537 , n28599 );
xor ( n28601 , n28537 , n28599 );
xor ( n28602 , n28591 , n28593 );
xor ( n28603 , n28602 , n28596 );
and ( n28604 , n23320 , n22032 );
and ( n28605 , n23074 , n22029 );
nor ( n28606 , n28604 , n28605 );
xnor ( n28607 , n28606 , n22027 );
and ( n28608 , n23503 , n22114 );
and ( n28609 , n23351 , n22112 );
nor ( n28610 , n28608 , n28609 );
xnor ( n28611 , n28610 , n22124 );
and ( n28612 , n28607 , n28611 );
xor ( n28613 , n28561 , n28565 );
xor ( n28614 , n28613 , n28570 );
and ( n28615 , n28611 , n28614 );
and ( n28616 , n28607 , n28614 );
or ( n28617 , n28612 , n28615 , n28616 );
xor ( n28618 , n28360 , n28364 );
and ( n28619 , n26003 , n21234 );
not ( n28620 , n28619 );
and ( n28621 , n28620 , n21246 );
and ( n28622 , n26003 , n21236 );
and ( n28623 , n26011 , n21234 );
nor ( n28624 , n28622 , n28623 );
xnor ( n28625 , n28624 , n21246 );
and ( n28626 , n28621 , n28625 );
and ( n28627 , n26011 , n21236 );
and ( n28628 , n26020 , n21234 );
nor ( n28629 , n28627 , n28628 );
xnor ( n28630 , n28629 , n21246 );
and ( n28631 , n28626 , n28630 );
and ( n28632 , n28630 , n28358 );
and ( n28633 , n28626 , n28358 );
or ( n28634 , n28631 , n28632 , n28633 );
and ( n28635 , n28618 , n28634 );
and ( n28636 , n26020 , n21236 );
and ( n28637 , n25898 , n21234 );
nor ( n28638 , n28636 , n28637 );
xnor ( n28639 , n28638 , n21246 );
and ( n28640 , n28634 , n28639 );
and ( n28641 , n28618 , n28639 );
or ( n28642 , n28635 , n28640 , n28641 );
and ( n28643 , n25898 , n21236 );
and ( n28644 , n25772 , n21234 );
nor ( n28645 , n28643 , n28644 );
xnor ( n28646 , n28645 , n21246 );
and ( n28647 , n28642 , n28646 );
xor ( n28648 , n28365 , n28369 );
xor ( n28649 , n28648 , n28070 );
and ( n28650 , n28646 , n28649 );
and ( n28651 , n28642 , n28649 );
or ( n28652 , n28647 , n28650 , n28651 );
and ( n28653 , n25179 , n21687 );
and ( n28654 , n25060 , n21685 );
nor ( n28655 , n28653 , n28654 );
xnor ( n28656 , n28655 , n21697 );
and ( n28657 , n28652 , n28656 );
xor ( n28658 , n28541 , n28545 );
xor ( n28659 , n28658 , n28548 );
and ( n28660 , n28656 , n28659 );
and ( n28661 , n28652 , n28659 );
or ( n28662 , n28657 , n28660 , n28661 );
and ( n28663 , n24460 , n21139 );
and ( n28664 , n24213 , n21137 );
nor ( n28665 , n28663 , n28664 );
xnor ( n28666 , n28665 , n21221 );
and ( n28667 , n28662 , n28666 );
and ( n28668 , n24662 , n21663 );
and ( n28669 , n24631 , n21661 );
nor ( n28670 , n28668 , n28669 );
xnor ( n28671 , n28670 , n21673 );
and ( n28672 , n28666 , n28671 );
and ( n28673 , n28662 , n28671 );
or ( n28674 , n28667 , n28672 , n28673 );
and ( n28675 , n23887 , n21414 );
and ( n28676 , n23651 , n21412 );
nor ( n28677 , n28675 , n28676 );
xnor ( n28678 , n28677 , n21480 );
and ( n28679 , n28674 , n28678 );
xor ( n28680 , n28477 , n28481 );
xor ( n28681 , n28680 , n28484 );
and ( n28682 , n28678 , n28681 );
and ( n28683 , n28674 , n28681 );
or ( n28684 , n28679 , n28682 , n28683 );
and ( n28685 , n28617 , n28684 );
xor ( n28686 , n28453 , n28457 );
xor ( n28687 , n28686 , n28460 );
and ( n28688 , n28684 , n28687 );
and ( n28689 , n28617 , n28687 );
or ( n28690 , n28685 , n28688 , n28689 );
xor ( n28691 , n28463 , n28497 );
xor ( n28692 , n28691 , n28502 );
and ( n28693 , n28690 , n28692 );
xor ( n28694 , n28583 , n28585 );
xor ( n28695 , n28694 , n28588 );
and ( n28696 , n28692 , n28695 );
and ( n28697 , n28690 , n28695 );
or ( n28698 , n28693 , n28696 , n28697 );
and ( n28699 , n28603 , n28698 );
xor ( n28700 , n28603 , n28698 );
xor ( n28701 , n28690 , n28692 );
xor ( n28702 , n28701 , n28695 );
and ( n28703 , n23351 , n22032 );
and ( n28704 , n23320 , n22029 );
nor ( n28705 , n28703 , n28704 );
xnor ( n28706 , n28705 , n22027 );
and ( n28707 , n23651 , n22114 );
and ( n28708 , n23503 , n22112 );
nor ( n28709 , n28707 , n28708 );
xnor ( n28710 , n28709 , n22124 );
and ( n28711 , n28706 , n28710 );
xor ( n28712 , n28662 , n28666 );
xor ( n28713 , n28712 , n28671 );
and ( n28714 , n28710 , n28713 );
and ( n28715 , n28706 , n28713 );
or ( n28716 , n28711 , n28714 , n28715 );
and ( n28717 , n25343 , n21687 );
and ( n28718 , n25179 , n21685 );
nor ( n28719 , n28717 , n28718 );
xnor ( n28720 , n28719 , n21697 );
and ( n28721 , n25553 , n21707 );
and ( n28722 , n25544 , n21705 );
nor ( n28723 , n28721 , n28722 );
xnor ( n28724 , n28723 , n21717 );
and ( n28725 , n28720 , n28724 );
xor ( n28726 , n28642 , n28646 );
xor ( n28727 , n28726 , n28649 );
and ( n28728 , n28724 , n28727 );
and ( n28729 , n28720 , n28727 );
or ( n28730 , n28725 , n28728 , n28729 );
and ( n28731 , n24631 , n21139 );
and ( n28732 , n24460 , n21137 );
nor ( n28733 , n28731 , n28732 );
xnor ( n28734 , n28733 , n21221 );
and ( n28735 , n28730 , n28734 );
and ( n28736 , n24812 , n21663 );
and ( n28737 , n24662 , n21661 );
nor ( n28738 , n28736 , n28737 );
xnor ( n28739 , n28738 , n21673 );
and ( n28740 , n28734 , n28739 );
and ( n28741 , n28730 , n28739 );
or ( n28742 , n28735 , n28740 , n28741 );
and ( n28743 , n23949 , n21414 );
and ( n28744 , n23887 , n21412 );
nor ( n28745 , n28743 , n28744 );
xnor ( n28746 , n28745 , n21480 );
and ( n28747 , n28742 , n28746 );
xor ( n28748 , n28551 , n28555 );
xor ( n28749 , n28748 , n28558 );
and ( n28750 , n28746 , n28749 );
and ( n28751 , n28742 , n28749 );
or ( n28752 , n28747 , n28750 , n28751 );
and ( n28753 , n28716 , n28752 );
xor ( n28754 , n28674 , n28678 );
xor ( n28755 , n28754 , n28681 );
and ( n28756 , n28752 , n28755 );
and ( n28757 , n28716 , n28755 );
or ( n28758 , n28753 , n28756 , n28757 );
xor ( n28759 , n28617 , n28684 );
xor ( n28760 , n28759 , n28687 );
and ( n28761 , n28758 , n28760 );
xor ( n28762 , n28573 , n28577 );
xor ( n28763 , n28762 , n28580 );
and ( n28764 , n28760 , n28763 );
and ( n28765 , n28758 , n28763 );
or ( n28766 , n28761 , n28764 , n28765 );
and ( n28767 , n28702 , n28766 );
xor ( n28768 , n28702 , n28766 );
xor ( n28769 , n28621 , n28625 );
and ( n28770 , n26003 , n21705 );
not ( n28771 , n28770 );
and ( n28772 , n28771 , n21717 );
and ( n28773 , n26003 , n21707 );
and ( n28774 , n26011 , n21705 );
nor ( n28775 , n28773 , n28774 );
xnor ( n28776 , n28775 , n21717 );
and ( n28777 , n28772 , n28776 );
and ( n28778 , n26011 , n21707 );
and ( n28779 , n26020 , n21705 );
nor ( n28780 , n28778 , n28779 );
xnor ( n28781 , n28780 , n21717 );
and ( n28782 , n28777 , n28781 );
and ( n28783 , n28781 , n28619 );
and ( n28784 , n28777 , n28619 );
or ( n28785 , n28782 , n28783 , n28784 );
and ( n28786 , n28769 , n28785 );
and ( n28787 , n26020 , n21707 );
and ( n28788 , n25898 , n21705 );
nor ( n28789 , n28787 , n28788 );
xnor ( n28790 , n28789 , n21717 );
and ( n28791 , n28785 , n28790 );
and ( n28792 , n28769 , n28790 );
or ( n28793 , n28786 , n28791 , n28792 );
and ( n28794 , n25898 , n21707 );
and ( n28795 , n25772 , n21705 );
nor ( n28796 , n28794 , n28795 );
xnor ( n28797 , n28796 , n21717 );
and ( n28798 , n28793 , n28797 );
xor ( n28799 , n28626 , n28630 );
xor ( n28800 , n28799 , n28358 );
and ( n28801 , n28797 , n28800 );
and ( n28802 , n28793 , n28800 );
or ( n28803 , n28798 , n28801 , n28802 );
and ( n28804 , n25179 , n21663 );
and ( n28805 , n25060 , n21661 );
nor ( n28806 , n28804 , n28805 );
xnor ( n28807 , n28806 , n21673 );
and ( n28808 , n28803 , n28807 );
and ( n28809 , n25544 , n21687 );
and ( n28810 , n25343 , n21685 );
nor ( n28811 , n28809 , n28810 );
xnor ( n28812 , n28811 , n21697 );
and ( n28813 , n25772 , n21707 );
and ( n28814 , n25553 , n21705 );
nor ( n28815 , n28813 , n28814 );
xnor ( n28816 , n28815 , n21717 );
xor ( n28817 , n28812 , n28816 );
xor ( n28818 , n28618 , n28634 );
xor ( n28819 , n28818 , n28639 );
xor ( n28820 , n28817 , n28819 );
and ( n28821 , n28807 , n28820 );
and ( n28822 , n28803 , n28820 );
or ( n28823 , n28808 , n28821 , n28822 );
and ( n28824 , n24460 , n21414 );
and ( n28825 , n24213 , n21412 );
nor ( n28826 , n28824 , n28825 );
xnor ( n28827 , n28826 , n21480 );
and ( n28828 , n28823 , n28827 );
and ( n28829 , n24662 , n21139 );
and ( n28830 , n24631 , n21137 );
nor ( n28831 , n28829 , n28830 );
xnor ( n28832 , n28831 , n21221 );
and ( n28833 , n28827 , n28832 );
and ( n28834 , n28823 , n28832 );
or ( n28835 , n28828 , n28833 , n28834 );
and ( n28836 , n23503 , n22032 );
and ( n28837 , n23351 , n22029 );
nor ( n28838 , n28836 , n28837 );
xnor ( n28839 , n28838 , n22027 );
and ( n28840 , n28835 , n28839 );
and ( n28841 , n23887 , n22114 );
and ( n28842 , n23651 , n22112 );
nor ( n28843 , n28841 , n28842 );
xnor ( n28844 , n28843 , n22124 );
and ( n28845 , n28839 , n28844 );
and ( n28846 , n28835 , n28844 );
or ( n28847 , n28840 , n28845 , n28846 );
and ( n28848 , n28812 , n28816 );
and ( n28849 , n28816 , n28819 );
and ( n28850 , n28812 , n28819 );
or ( n28851 , n28848 , n28849 , n28850 );
and ( n28852 , n25060 , n21663 );
and ( n28853 , n24812 , n21661 );
nor ( n28854 , n28852 , n28853 );
xnor ( n28855 , n28854 , n21673 );
and ( n28856 , n28851 , n28855 );
xor ( n28857 , n28720 , n28724 );
xor ( n28858 , n28857 , n28727 );
and ( n28859 , n28855 , n28858 );
and ( n28860 , n28851 , n28858 );
or ( n28861 , n28856 , n28859 , n28860 );
and ( n28862 , n24213 , n21414 );
and ( n28863 , n23949 , n21412 );
nor ( n28864 , n28862 , n28863 );
xnor ( n28865 , n28864 , n21480 );
and ( n28866 , n28861 , n28865 );
xor ( n28867 , n28652 , n28656 );
xor ( n28868 , n28867 , n28659 );
and ( n28869 , n28865 , n28868 );
and ( n28870 , n28861 , n28868 );
or ( n28871 , n28866 , n28869 , n28870 );
and ( n28872 , n28847 , n28871 );
xor ( n28873 , n28742 , n28746 );
xor ( n28874 , n28873 , n28749 );
and ( n28875 , n28871 , n28874 );
and ( n28876 , n28847 , n28874 );
or ( n28877 , n28872 , n28875 , n28876 );
xor ( n28878 , n28607 , n28611 );
xor ( n28879 , n28878 , n28614 );
and ( n28880 , n28877 , n28879 );
xor ( n28881 , n28716 , n28752 );
xor ( n28882 , n28881 , n28755 );
and ( n28883 , n28879 , n28882 );
and ( n28884 , n28877 , n28882 );
or ( n28885 , n28880 , n28883 , n28884 );
xor ( n28886 , n28758 , n28760 );
xor ( n28887 , n28886 , n28763 );
and ( n28888 , n28885 , n28887 );
xor ( n28889 , n28885 , n28887 );
xor ( n28890 , n28877 , n28879 );
xor ( n28891 , n28890 , n28882 );
and ( n28892 , n23651 , n22032 );
and ( n28893 , n23503 , n22029 );
nor ( n28894 , n28892 , n28893 );
xnor ( n28895 , n28894 , n22027 );
and ( n28896 , n23949 , n22114 );
and ( n28897 , n23887 , n22112 );
nor ( n28898 , n28896 , n28897 );
xnor ( n28899 , n28898 , n22124 );
and ( n28900 , n28895 , n28899 );
xor ( n28901 , n28851 , n28855 );
xor ( n28902 , n28901 , n28858 );
and ( n28903 , n28899 , n28902 );
and ( n28904 , n28895 , n28902 );
or ( n28905 , n28900 , n28903 , n28904 );
xor ( n28906 , n28730 , n28734 );
xor ( n28907 , n28906 , n28739 );
and ( n28908 , n28905 , n28907 );
xor ( n28909 , n28861 , n28865 );
xor ( n28910 , n28909 , n28868 );
and ( n28911 , n28907 , n28910 );
and ( n28912 , n28905 , n28910 );
or ( n28913 , n28908 , n28911 , n28912 );
xor ( n28914 , n28706 , n28710 );
xor ( n28915 , n28914 , n28713 );
and ( n28916 , n28913 , n28915 );
xor ( n28917 , n28847 , n28871 );
xor ( n28918 , n28917 , n28874 );
and ( n28919 , n28915 , n28918 );
and ( n28920 , n28913 , n28918 );
or ( n28921 , n28916 , n28919 , n28920 );
and ( n28922 , n28891 , n28921 );
xor ( n28923 , n28891 , n28921 );
xor ( n28924 , n28913 , n28915 );
xor ( n28925 , n28924 , n28918 );
and ( n28926 , n25544 , n21663 );
and ( n28927 , n25343 , n21661 );
nor ( n28928 , n28926 , n28927 );
xnor ( n28929 , n28928 , n21673 );
and ( n28930 , n25772 , n21687 );
and ( n28931 , n25553 , n21685 );
nor ( n28932 , n28930 , n28931 );
xnor ( n28933 , n28932 , n21697 );
and ( n28934 , n28929 , n28933 );
xor ( n28935 , n28769 , n28785 );
xor ( n28936 , n28935 , n28790 );
and ( n28937 , n28933 , n28936 );
and ( n28938 , n28929 , n28936 );
or ( n28939 , n28934 , n28937 , n28938 );
and ( n28940 , n25060 , n21139 );
and ( n28941 , n24812 , n21137 );
nor ( n28942 , n28940 , n28941 );
xnor ( n28943 , n28942 , n21221 );
and ( n28944 , n28939 , n28943 );
and ( n28945 , n25343 , n21663 );
and ( n28946 , n25179 , n21661 );
nor ( n28947 , n28945 , n28946 );
xnor ( n28948 , n28947 , n21673 );
and ( n28949 , n25553 , n21687 );
and ( n28950 , n25544 , n21685 );
nor ( n28951 , n28949 , n28950 );
xnor ( n28952 , n28951 , n21697 );
xor ( n28953 , n28948 , n28952 );
xor ( n28954 , n28793 , n28797 );
xor ( n28955 , n28954 , n28800 );
xor ( n28956 , n28953 , n28955 );
and ( n28957 , n28943 , n28956 );
and ( n28958 , n28939 , n28956 );
or ( n28959 , n28944 , n28957 , n28958 );
and ( n28960 , n24213 , n22114 );
and ( n28961 , n23949 , n22112 );
nor ( n28962 , n28960 , n28961 );
xnor ( n28963 , n28962 , n22124 );
and ( n28964 , n28959 , n28963 );
and ( n28965 , n24812 , n21139 );
and ( n28966 , n24662 , n21137 );
nor ( n28967 , n28965 , n28966 );
xnor ( n28968 , n28967 , n21221 );
and ( n28969 , n28963 , n28968 );
and ( n28970 , n28959 , n28968 );
or ( n28971 , n28964 , n28969 , n28970 );
and ( n28972 , n28948 , n28952 );
and ( n28973 , n28952 , n28955 );
and ( n28974 , n28948 , n28955 );
or ( n28975 , n28972 , n28973 , n28974 );
and ( n28976 , n24631 , n21414 );
and ( n28977 , n24460 , n21412 );
nor ( n28978 , n28976 , n28977 );
xnor ( n28979 , n28978 , n21480 );
and ( n28980 , n28975 , n28979 );
xor ( n28981 , n28803 , n28807 );
xor ( n28982 , n28981 , n28820 );
and ( n28983 , n28979 , n28982 );
and ( n28984 , n28975 , n28982 );
or ( n28985 , n28980 , n28983 , n28984 );
and ( n28986 , n28971 , n28985 );
xor ( n28987 , n28823 , n28827 );
xor ( n28988 , n28987 , n28832 );
and ( n28989 , n28985 , n28988 );
and ( n28990 , n28971 , n28988 );
or ( n28991 , n28986 , n28989 , n28990 );
xor ( n28992 , n28835 , n28839 );
xor ( n28993 , n28992 , n28844 );
and ( n28994 , n28991 , n28993 );
xor ( n28995 , n28905 , n28907 );
xor ( n28996 , n28995 , n28910 );
and ( n28997 , n28993 , n28996 );
and ( n28998 , n28991 , n28996 );
or ( n28999 , n28994 , n28997 , n28998 );
and ( n29000 , n28925 , n28999 );
xor ( n29001 , n28925 , n28999 );
xor ( n29002 , n28991 , n28993 );
xor ( n29003 , n29002 , n28996 );
xor ( n29004 , n28772 , n28776 );
and ( n29005 , n26003 , n21685 );
not ( n29006 , n29005 );
and ( n29007 , n29006 , n21697 );
and ( n29008 , n26003 , n21687 );
and ( n29009 , n26011 , n21685 );
nor ( n29010 , n29008 , n29009 );
xnor ( n29011 , n29010 , n21697 );
and ( n29012 , n29007 , n29011 );
and ( n29013 , n26011 , n21687 );
and ( n29014 , n26020 , n21685 );
nor ( n29015 , n29013 , n29014 );
xnor ( n29016 , n29015 , n21697 );
and ( n29017 , n29012 , n29016 );
and ( n29018 , n29016 , n28770 );
and ( n29019 , n29012 , n28770 );
or ( n29020 , n29017 , n29018 , n29019 );
and ( n29021 , n29004 , n29020 );
and ( n29022 , n26020 , n21687 );
and ( n29023 , n25898 , n21685 );
nor ( n29024 , n29022 , n29023 );
xnor ( n29025 , n29024 , n21697 );
and ( n29026 , n29020 , n29025 );
and ( n29027 , n29004 , n29025 );
or ( n29028 , n29021 , n29026 , n29027 );
and ( n29029 , n25898 , n21687 );
and ( n29030 , n25772 , n21685 );
nor ( n29031 , n29029 , n29030 );
xnor ( n29032 , n29031 , n21697 );
and ( n29033 , n29028 , n29032 );
xor ( n29034 , n28777 , n28781 );
xor ( n29035 , n29034 , n28619 );
and ( n29036 , n29032 , n29035 );
and ( n29037 , n29028 , n29035 );
or ( n29038 , n29033 , n29036 , n29037 );
and ( n29039 , n25179 , n21139 );
and ( n29040 , n25060 , n21137 );
nor ( n29041 , n29039 , n29040 );
xnor ( n29042 , n29041 , n21221 );
and ( n29043 , n29038 , n29042 );
xor ( n29044 , n28929 , n28933 );
xor ( n29045 , n29044 , n28936 );
and ( n29046 , n29042 , n29045 );
and ( n29047 , n29038 , n29045 );
or ( n29048 , n29043 , n29046 , n29047 );
and ( n29049 , n24460 , n22114 );
and ( n29050 , n24213 , n22112 );
nor ( n29051 , n29049 , n29050 );
xnor ( n29052 , n29051 , n22124 );
and ( n29053 , n29048 , n29052 );
and ( n29054 , n24662 , n21414 );
and ( n29055 , n24631 , n21412 );
nor ( n29056 , n29054 , n29055 );
xnor ( n29057 , n29056 , n21480 );
and ( n29058 , n29052 , n29057 );
and ( n29059 , n29048 , n29057 );
or ( n29060 , n29053 , n29058 , n29059 );
and ( n29061 , n23887 , n22032 );
and ( n29062 , n23651 , n22029 );
nor ( n29063 , n29061 , n29062 );
xnor ( n29064 , n29063 , n22027 );
and ( n29065 , n29060 , n29064 );
xor ( n29066 , n28975 , n28979 );
xor ( n29067 , n29066 , n28982 );
and ( n29068 , n29064 , n29067 );
and ( n29069 , n29060 , n29067 );
or ( n29070 , n29065 , n29068 , n29069 );
xor ( n29071 , n28971 , n28985 );
xor ( n29072 , n29071 , n28988 );
and ( n29073 , n29070 , n29072 );
xor ( n29074 , n28895 , n28899 );
xor ( n29075 , n29074 , n28902 );
and ( n29076 , n29072 , n29075 );
and ( n29077 , n29070 , n29075 );
or ( n29078 , n29073 , n29076 , n29077 );
and ( n29079 , n29003 , n29078 );
xor ( n29080 , n29003 , n29078 );
and ( n29081 , n25343 , n21139 );
and ( n29082 , n25179 , n21137 );
nor ( n29083 , n29081 , n29082 );
xnor ( n29084 , n29083 , n21221 );
and ( n29085 , n25553 , n21663 );
and ( n29086 , n25544 , n21661 );
nor ( n29087 , n29085 , n29086 );
xnor ( n29088 , n29087 , n21673 );
and ( n29089 , n29084 , n29088 );
xor ( n29090 , n29028 , n29032 );
xor ( n29091 , n29090 , n29035 );
and ( n29092 , n29088 , n29091 );
and ( n29093 , n29084 , n29091 );
or ( n29094 , n29089 , n29092 , n29093 );
and ( n29095 , n24631 , n22114 );
and ( n29096 , n24460 , n22112 );
nor ( n29097 , n29095 , n29096 );
xnor ( n29098 , n29097 , n22124 );
and ( n29099 , n29094 , n29098 );
xor ( n29100 , n29038 , n29042 );
xor ( n29101 , n29100 , n29045 );
and ( n29102 , n29098 , n29101 );
and ( n29103 , n29094 , n29101 );
or ( n29104 , n29099 , n29102 , n29103 );
and ( n29105 , n23949 , n22032 );
and ( n29106 , n23887 , n22029 );
nor ( n29107 , n29105 , n29106 );
xnor ( n29108 , n29107 , n22027 );
and ( n29109 , n29104 , n29108 );
xor ( n29110 , n28939 , n28943 );
xor ( n29111 , n29110 , n28956 );
and ( n29112 , n29108 , n29111 );
and ( n29113 , n29104 , n29111 );
or ( n29114 , n29109 , n29112 , n29113 );
xor ( n29115 , n28959 , n28963 );
xor ( n29116 , n29115 , n28968 );
and ( n29117 , n29114 , n29116 );
xor ( n29118 , n29060 , n29064 );
xor ( n29119 , n29118 , n29067 );
and ( n29120 , n29116 , n29119 );
and ( n29121 , n29114 , n29119 );
or ( n29122 , n29117 , n29120 , n29121 );
xor ( n29123 , n29070 , n29072 );
xor ( n29124 , n29123 , n29075 );
and ( n29125 , n29122 , n29124 );
xor ( n29126 , n29122 , n29124 );
xor ( n29127 , n29114 , n29116 );
xor ( n29128 , n29127 , n29119 );
and ( n29129 , n25544 , n21139 );
and ( n29130 , n25343 , n21137 );
nor ( n29131 , n29129 , n29130 );
xnor ( n29132 , n29131 , n21221 );
and ( n29133 , n25772 , n21663 );
and ( n29134 , n25553 , n21661 );
nor ( n29135 , n29133 , n29134 );
xnor ( n29136 , n29135 , n21673 );
and ( n29137 , n29132 , n29136 );
xor ( n29138 , n29004 , n29020 );
xor ( n29139 , n29138 , n29025 );
and ( n29140 , n29136 , n29139 );
and ( n29141 , n29132 , n29139 );
or ( n29142 , n29137 , n29140 , n29141 );
and ( n29143 , n25060 , n21414 );
and ( n29144 , n24812 , n21412 );
nor ( n29145 , n29143 , n29144 );
xnor ( n29146 , n29145 , n21480 );
and ( n29147 , n29142 , n29146 );
xor ( n29148 , n29084 , n29088 );
xor ( n29149 , n29148 , n29091 );
and ( n29150 , n29146 , n29149 );
and ( n29151 , n29142 , n29149 );
or ( n29152 , n29147 , n29150 , n29151 );
and ( n29153 , n24213 , n22032 );
and ( n29154 , n23949 , n22029 );
nor ( n29155 , n29153 , n29154 );
xnor ( n29156 , n29155 , n22027 );
and ( n29157 , n29152 , n29156 );
and ( n29158 , n24812 , n21414 );
and ( n29159 , n24662 , n21412 );
nor ( n29160 , n29158 , n29159 );
xnor ( n29161 , n29160 , n21480 );
and ( n29162 , n29156 , n29161 );
and ( n29163 , n29152 , n29161 );
or ( n29164 , n29157 , n29162 , n29163 );
xor ( n29165 , n29048 , n29052 );
xor ( n29166 , n29165 , n29057 );
and ( n29167 , n29164 , n29166 );
xor ( n29168 , n29104 , n29108 );
xor ( n29169 , n29168 , n29111 );
and ( n29170 , n29166 , n29169 );
and ( n29171 , n29164 , n29169 );
or ( n29172 , n29167 , n29170 , n29171 );
and ( n29173 , n29128 , n29172 );
xor ( n29174 , n29128 , n29172 );
xor ( n29175 , n29164 , n29166 );
xor ( n29176 , n29175 , n29169 );
xor ( n29177 , n29007 , n29011 );
and ( n29178 , n26003 , n21661 );
not ( n29179 , n29178 );
and ( n29180 , n29179 , n21673 );
and ( n29181 , n26003 , n21663 );
and ( n29182 , n26011 , n21661 );
nor ( n29183 , n29181 , n29182 );
xnor ( n29184 , n29183 , n21673 );
and ( n29185 , n29180 , n29184 );
and ( n29186 , n26011 , n21663 );
and ( n29187 , n26020 , n21661 );
nor ( n29188 , n29186 , n29187 );
xnor ( n29189 , n29188 , n21673 );
and ( n29190 , n29185 , n29189 );
and ( n29191 , n29189 , n29005 );
and ( n29192 , n29185 , n29005 );
or ( n29193 , n29190 , n29191 , n29192 );
and ( n29194 , n29177 , n29193 );
and ( n29195 , n26020 , n21663 );
and ( n29196 , n25898 , n21661 );
nor ( n29197 , n29195 , n29196 );
xnor ( n29198 , n29197 , n21673 );
and ( n29199 , n29193 , n29198 );
and ( n29200 , n29177 , n29198 );
or ( n29201 , n29194 , n29199 , n29200 );
and ( n29202 , n25898 , n21663 );
and ( n29203 , n25772 , n21661 );
nor ( n29204 , n29202 , n29203 );
xnor ( n29205 , n29204 , n21673 );
and ( n29206 , n29201 , n29205 );
xor ( n29207 , n29012 , n29016 );
xor ( n29208 , n29207 , n28770 );
and ( n29209 , n29205 , n29208 );
and ( n29210 , n29201 , n29208 );
or ( n29211 , n29206 , n29209 , n29210 );
and ( n29212 , n25179 , n21414 );
and ( n29213 , n25060 , n21412 );
nor ( n29214 , n29212 , n29213 );
xnor ( n29215 , n29214 , n21480 );
and ( n29216 , n29211 , n29215 );
xor ( n29217 , n29132 , n29136 );
xor ( n29218 , n29217 , n29139 );
and ( n29219 , n29215 , n29218 );
and ( n29220 , n29211 , n29218 );
or ( n29221 , n29216 , n29219 , n29220 );
and ( n29222 , n24460 , n22032 );
and ( n29223 , n24213 , n22029 );
nor ( n29224 , n29222 , n29223 );
xnor ( n29225 , n29224 , n22027 );
and ( n29226 , n29221 , n29225 );
and ( n29227 , n24662 , n22114 );
and ( n29228 , n24631 , n22112 );
nor ( n29229 , n29227 , n29228 );
xnor ( n29230 , n29229 , n22124 );
and ( n29231 , n29225 , n29230 );
and ( n29232 , n29221 , n29230 );
or ( n29233 , n29226 , n29231 , n29232 );
xor ( n29234 , n29152 , n29156 );
xor ( n29235 , n29234 , n29161 );
and ( n29236 , n29233 , n29235 );
xor ( n29237 , n29094 , n29098 );
xor ( n29238 , n29237 , n29101 );
and ( n29239 , n29235 , n29238 );
and ( n29240 , n29233 , n29238 );
or ( n29241 , n29236 , n29239 , n29240 );
and ( n29242 , n29176 , n29241 );
xor ( n29243 , n29176 , n29241 );
and ( n29244 , n25343 , n21414 );
and ( n29245 , n25179 , n21412 );
nor ( n29246 , n29244 , n29245 );
xnor ( n29247 , n29246 , n21480 );
and ( n29248 , n25553 , n21139 );
and ( n29249 , n25544 , n21137 );
nor ( n29250 , n29248 , n29249 );
xnor ( n29251 , n29250 , n21221 );
and ( n29252 , n29247 , n29251 );
xor ( n29253 , n29201 , n29205 );
xor ( n29254 , n29253 , n29208 );
and ( n29255 , n29251 , n29254 );
and ( n29256 , n29247 , n29254 );
or ( n29257 , n29252 , n29255 , n29256 );
and ( n29258 , n24812 , n22114 );
and ( n29259 , n24662 , n22112 );
nor ( n29260 , n29258 , n29259 );
xnor ( n29261 , n29260 , n22124 );
and ( n29262 , n29257 , n29261 );
xor ( n29263 , n29211 , n29215 );
xor ( n29264 , n29263 , n29218 );
and ( n29265 , n29261 , n29264 );
and ( n29266 , n29257 , n29264 );
or ( n29267 , n29262 , n29265 , n29266 );
xor ( n29268 , n29221 , n29225 );
xor ( n29269 , n29268 , n29230 );
and ( n29270 , n29267 , n29269 );
xor ( n29271 , n29142 , n29146 );
xor ( n29272 , n29271 , n29149 );
and ( n29273 , n29269 , n29272 );
and ( n29274 , n29267 , n29272 );
or ( n29275 , n29270 , n29273 , n29274 );
xor ( n29276 , n29233 , n29235 );
xor ( n29277 , n29276 , n29238 );
and ( n29278 , n29275 , n29277 );
xor ( n29279 , n29275 , n29277 );
xor ( n29280 , n29267 , n29269 );
xor ( n29281 , n29280 , n29272 );
and ( n29282 , n25544 , n21414 );
and ( n29283 , n25343 , n21412 );
nor ( n29284 , n29282 , n29283 );
xnor ( n29285 , n29284 , n21480 );
and ( n29286 , n25772 , n21139 );
and ( n29287 , n25553 , n21137 );
nor ( n29288 , n29286 , n29287 );
xnor ( n29289 , n29288 , n21221 );
and ( n29290 , n29285 , n29289 );
xor ( n29291 , n29177 , n29193 );
xor ( n29292 , n29291 , n29198 );
and ( n29293 , n29289 , n29292 );
and ( n29294 , n29285 , n29292 );
or ( n29295 , n29290 , n29293 , n29294 );
and ( n29296 , n25060 , n22114 );
and ( n29297 , n24812 , n22112 );
nor ( n29298 , n29296 , n29297 );
xnor ( n29299 , n29298 , n22124 );
and ( n29300 , n29295 , n29299 );
xor ( n29301 , n29247 , n29251 );
xor ( n29302 , n29301 , n29254 );
and ( n29303 , n29299 , n29302 );
and ( n29304 , n29295 , n29302 );
or ( n29305 , n29300 , n29303 , n29304 );
and ( n29306 , n24631 , n22032 );
and ( n29307 , n24460 , n22029 );
nor ( n29308 , n29306 , n29307 );
xnor ( n29309 , n29308 , n22027 );
and ( n29310 , n29305 , n29309 );
xor ( n29311 , n29257 , n29261 );
xor ( n29312 , n29311 , n29264 );
and ( n29313 , n29309 , n29312 );
and ( n29314 , n29305 , n29312 );
or ( n29315 , n29310 , n29313 , n29314 );
and ( n29316 , n29281 , n29315 );
xor ( n29317 , n29281 , n29315 );
xor ( n29318 , n29305 , n29309 );
xor ( n29319 , n29318 , n29312 );
xor ( n29320 , n29180 , n29184 );
and ( n29321 , n26003 , n21137 );
not ( n29322 , n29321 );
and ( n29323 , n29322 , n21221 );
and ( n29324 , n26003 , n21139 );
and ( n29325 , n26011 , n21137 );
nor ( n29326 , n29324 , n29325 );
xnor ( n29327 , n29326 , n21221 );
and ( n29328 , n29323 , n29327 );
and ( n29329 , n26011 , n21139 );
and ( n29330 , n26020 , n21137 );
nor ( n29331 , n29329 , n29330 );
xnor ( n29332 , n29331 , n21221 );
and ( n29333 , n29328 , n29332 );
and ( n29334 , n29332 , n29178 );
and ( n29335 , n29328 , n29178 );
or ( n29336 , n29333 , n29334 , n29335 );
and ( n29337 , n29320 , n29336 );
and ( n29338 , n26020 , n21139 );
and ( n29339 , n25898 , n21137 );
nor ( n29340 , n29338 , n29339 );
xnor ( n29341 , n29340 , n21221 );
and ( n29342 , n29336 , n29341 );
and ( n29343 , n29320 , n29341 );
or ( n29344 , n29337 , n29342 , n29343 );
and ( n29345 , n25898 , n21139 );
and ( n29346 , n25772 , n21137 );
nor ( n29347 , n29345 , n29346 );
xnor ( n29348 , n29347 , n21221 );
and ( n29349 , n29344 , n29348 );
xor ( n29350 , n29185 , n29189 );
xor ( n29351 , n29350 , n29005 );
and ( n29352 , n29348 , n29351 );
and ( n29353 , n29344 , n29351 );
or ( n29354 , n29349 , n29352 , n29353 );
and ( n29355 , n25179 , n22114 );
and ( n29356 , n25060 , n22112 );
nor ( n29357 , n29355 , n29356 );
xnor ( n29358 , n29357 , n22124 );
and ( n29359 , n29354 , n29358 );
xor ( n29360 , n29285 , n29289 );
xor ( n29361 , n29360 , n29292 );
and ( n29362 , n29358 , n29361 );
and ( n29363 , n29354 , n29361 );
or ( n29364 , n29359 , n29362 , n29363 );
and ( n29365 , n24662 , n22032 );
and ( n29366 , n24631 , n22029 );
nor ( n29367 , n29365 , n29366 );
xnor ( n29368 , n29367 , n22027 );
and ( n29369 , n29364 , n29368 );
xor ( n29370 , n29295 , n29299 );
xor ( n29371 , n29370 , n29302 );
and ( n29372 , n29368 , n29371 );
and ( n29373 , n29364 , n29371 );
or ( n29374 , n29369 , n29372 , n29373 );
and ( n29375 , n29319 , n29374 );
xor ( n29376 , n29319 , n29374 );
and ( n29377 , n25343 , n22114 );
and ( n29378 , n25179 , n22112 );
nor ( n29379 , n29377 , n29378 );
xnor ( n29380 , n29379 , n22124 );
and ( n29381 , n25553 , n21414 );
and ( n29382 , n25544 , n21412 );
nor ( n29383 , n29381 , n29382 );
xnor ( n29384 , n29383 , n21480 );
and ( n29385 , n29380 , n29384 );
xor ( n29386 , n29344 , n29348 );
xor ( n29387 , n29386 , n29351 );
and ( n29388 , n29384 , n29387 );
and ( n29389 , n29380 , n29387 );
or ( n29390 , n29385 , n29388 , n29389 );
and ( n29391 , n24812 , n22032 );
and ( n29392 , n24662 , n22029 );
nor ( n29393 , n29391 , n29392 );
xnor ( n29394 , n29393 , n22027 );
and ( n29395 , n29390 , n29394 );
xor ( n29396 , n29354 , n29358 );
xor ( n29397 , n29396 , n29361 );
and ( n29398 , n29394 , n29397 );
and ( n29399 , n29390 , n29397 );
or ( n29400 , n29395 , n29398 , n29399 );
xor ( n29401 , n29364 , n29368 );
xor ( n29402 , n29401 , n29371 );
and ( n29403 , n29400 , n29402 );
xor ( n29404 , n29400 , n29402 );
xor ( n29405 , n29390 , n29394 );
xor ( n29406 , n29405 , n29397 );
and ( n29407 , n25544 , n22114 );
and ( n29408 , n25343 , n22112 );
nor ( n29409 , n29407 , n29408 );
xnor ( n29410 , n29409 , n22124 );
and ( n29411 , n25772 , n21414 );
and ( n29412 , n25553 , n21412 );
nor ( n29413 , n29411 , n29412 );
xnor ( n29414 , n29413 , n21480 );
and ( n29415 , n29410 , n29414 );
xor ( n29416 , n29320 , n29336 );
xor ( n29417 , n29416 , n29341 );
and ( n29418 , n29414 , n29417 );
and ( n29419 , n29410 , n29417 );
or ( n29420 , n29415 , n29418 , n29419 );
and ( n29421 , n25060 , n22032 );
and ( n29422 , n24812 , n22029 );
nor ( n29423 , n29421 , n29422 );
xnor ( n29424 , n29423 , n22027 );
and ( n29425 , n29420 , n29424 );
xor ( n29426 , n29380 , n29384 );
xor ( n29427 , n29426 , n29387 );
and ( n29428 , n29424 , n29427 );
and ( n29429 , n29420 , n29427 );
or ( n29430 , n29425 , n29428 , n29429 );
and ( n29431 , n29406 , n29430 );
xor ( n29432 , n29406 , n29430 );
xor ( n29433 , n29323 , n29327 );
and ( n29434 , n26003 , n21412 );
not ( n29435 , n29434 );
and ( n29436 , n29435 , n21480 );
and ( n29437 , n26003 , n21414 );
and ( n29438 , n26011 , n21412 );
nor ( n29439 , n29437 , n29438 );
xnor ( n29440 , n29439 , n21480 );
and ( n29441 , n29436 , n29440 );
and ( n29442 , n26011 , n21414 );
and ( n29443 , n26020 , n21412 );
nor ( n29444 , n29442 , n29443 );
xnor ( n29445 , n29444 , n21480 );
and ( n29446 , n29441 , n29445 );
and ( n29447 , n29445 , n29321 );
and ( n29448 , n29441 , n29321 );
or ( n29449 , n29446 , n29447 , n29448 );
and ( n29450 , n29433 , n29449 );
and ( n29451 , n26020 , n21414 );
and ( n29452 , n25898 , n21412 );
nor ( n29453 , n29451 , n29452 );
xnor ( n29454 , n29453 , n21480 );
and ( n29455 , n29449 , n29454 );
and ( n29456 , n29433 , n29454 );
or ( n29457 , n29450 , n29455 , n29456 );
and ( n29458 , n25898 , n21414 );
and ( n29459 , n25772 , n21412 );
nor ( n29460 , n29458 , n29459 );
xnor ( n29461 , n29460 , n21480 );
and ( n29462 , n29457 , n29461 );
xor ( n29463 , n29328 , n29332 );
xor ( n29464 , n29463 , n29178 );
and ( n29465 , n29461 , n29464 );
and ( n29466 , n29457 , n29464 );
or ( n29467 , n29462 , n29465 , n29466 );
and ( n29468 , n25179 , n22032 );
and ( n29469 , n25060 , n22029 );
nor ( n29470 , n29468 , n29469 );
xnor ( n29471 , n29470 , n22027 );
and ( n29472 , n29467 , n29471 );
xor ( n29473 , n29410 , n29414 );
xor ( n29474 , n29473 , n29417 );
and ( n29475 , n29471 , n29474 );
and ( n29476 , n29467 , n29474 );
or ( n29477 , n29472 , n29475 , n29476 );
xor ( n29478 , n29420 , n29424 );
xor ( n29479 , n29478 , n29427 );
and ( n29480 , n29477 , n29479 );
xor ( n29481 , n29477 , n29479 );
xor ( n29482 , n29467 , n29471 );
xor ( n29483 , n29482 , n29474 );
and ( n29484 , n25343 , n22032 );
and ( n29485 , n25179 , n22029 );
nor ( n29486 , n29484 , n29485 );
xnor ( n29487 , n29486 , n22027 );
and ( n29488 , n25553 , n22114 );
and ( n29489 , n25544 , n22112 );
nor ( n29490 , n29488 , n29489 );
xnor ( n29491 , n29490 , n22124 );
and ( n29492 , n29487 , n29491 );
xor ( n29493 , n29457 , n29461 );
xor ( n29494 , n29493 , n29464 );
and ( n29495 , n29491 , n29494 );
and ( n29496 , n29487 , n29494 );
or ( n29497 , n29492 , n29495 , n29496 );
and ( n29498 , n29483 , n29497 );
xor ( n29499 , n29483 , n29497 );
and ( n29500 , n25544 , n22032 );
and ( n29501 , n25343 , n22029 );
nor ( n29502 , n29500 , n29501 );
xnor ( n29503 , n29502 , n22027 );
and ( n29504 , n25772 , n22114 );
and ( n29505 , n25553 , n22112 );
nor ( n29506 , n29504 , n29505 );
xnor ( n29507 , n29506 , n22124 );
and ( n29508 , n29503 , n29507 );
xor ( n29509 , n29433 , n29449 );
xor ( n29510 , n29509 , n29454 );
and ( n29511 , n29507 , n29510 );
and ( n29512 , n29503 , n29510 );
or ( n29513 , n29508 , n29511 , n29512 );
xor ( n29514 , n29487 , n29491 );
xor ( n29515 , n29514 , n29494 );
and ( n29516 , n29513 , n29515 );
xor ( n29517 , n29513 , n29515 );
xor ( n29518 , n29503 , n29507 );
xor ( n29519 , n29518 , n29510 );
xor ( n29520 , n29436 , n29440 );
and ( n29521 , n26003 , n22112 );
not ( n29522 , n29521 );
and ( n29523 , n29522 , n22124 );
and ( n29524 , n26003 , n22114 );
and ( n29525 , n26011 , n22112 );
nor ( n29526 , n29524 , n29525 );
xnor ( n29527 , n29526 , n22124 );
and ( n29528 , n29523 , n29527 );
and ( n29529 , n26011 , n22114 );
and ( n29530 , n26020 , n22112 );
nor ( n29531 , n29529 , n29530 );
xnor ( n29532 , n29531 , n22124 );
and ( n29533 , n29528 , n29532 );
and ( n29534 , n29532 , n29434 );
and ( n29535 , n29528 , n29434 );
or ( n29536 , n29533 , n29534 , n29535 );
and ( n29537 , n29520 , n29536 );
and ( n29538 , n26020 , n22114 );
and ( n29539 , n25898 , n22112 );
nor ( n29540 , n29538 , n29539 );
xnor ( n29541 , n29540 , n22124 );
and ( n29542 , n29536 , n29541 );
and ( n29543 , n29520 , n29541 );
or ( n29544 , n29537 , n29542 , n29543 );
and ( n29545 , n25898 , n22114 );
and ( n29546 , n25772 , n22112 );
nor ( n29547 , n29545 , n29546 );
xnor ( n29548 , n29547 , n22124 );
and ( n29549 , n29544 , n29548 );
xor ( n29550 , n29441 , n29445 );
xor ( n29551 , n29550 , n29321 );
and ( n29552 , n29548 , n29551 );
and ( n29553 , n29544 , n29551 );
or ( n29554 , n29549 , n29552 , n29553 );
and ( n29555 , n29519 , n29554 );
xor ( n29556 , n29519 , n29554 );
and ( n29557 , n25553 , n22032 );
and ( n29558 , n25544 , n22029 );
nor ( n29559 , n29557 , n29558 );
xnor ( n29560 , n29559 , n22027 );
xor ( n29561 , n29544 , n29548 );
xor ( n29562 , n29561 , n29551 );
and ( n29563 , n29560 , n29562 );
xor ( n29564 , n29560 , n29562 );
and ( n29565 , n25772 , n22032 );
and ( n29566 , n25553 , n22029 );
nor ( n29567 , n29565 , n29566 );
xnor ( n29568 , n29567 , n22027 );
xor ( n29569 , n29520 , n29536 );
xor ( n29570 , n29569 , n29541 );
and ( n29571 , n29568 , n29570 );
xor ( n29572 , n29568 , n29570 );
and ( n29573 , n25898 , n22032 );
and ( n29574 , n25772 , n22029 );
nor ( n29575 , n29573 , n29574 );
xnor ( n29576 , n29575 , n22027 );
xor ( n29577 , n29528 , n29532 );
xor ( n29578 , n29577 , n29434 );
and ( n29579 , n29576 , n29578 );
xor ( n29580 , n29576 , n29578 );
and ( n29581 , n26020 , n22032 );
and ( n29582 , n25898 , n22029 );
nor ( n29583 , n29581 , n29582 );
xnor ( n29584 , n29583 , n22027 );
xor ( n29585 , n29523 , n29527 );
and ( n29586 , n29584 , n29585 );
xor ( n29587 , n29584 , n29585 );
and ( n29588 , n26011 , n22032 );
and ( n29589 , n26020 , n22029 );
nor ( n29590 , n29588 , n29589 );
xnor ( n29591 , n29590 , n22027 );
and ( n29592 , n29591 , n29521 );
xor ( n29593 , n29591 , n29521 );
and ( n29594 , n26003 , n22032 );
and ( n29595 , n26011 , n22029 );
nor ( n29596 , n29594 , n29595 );
xnor ( n29597 , n29596 , n22027 );
and ( n29598 , n26003 , n22029 );
not ( n29599 , n29598 );
and ( n29600 , n29599 , n22027 );
and ( n29601 , n29597 , n29600 );
and ( n29602 , n29593 , n29601 );
or ( n29603 , n29592 , n29602 );
and ( n29604 , n29587 , n29603 );
or ( n29605 , n29586 , n29604 );
and ( n29606 , n29580 , n29605 );
or ( n29607 , n29579 , n29606 );
and ( n29608 , n29572 , n29607 );
or ( n29609 , n29571 , n29608 );
and ( n29610 , n29564 , n29609 );
or ( n29611 , n29563 , n29610 );
and ( n29612 , n29556 , n29611 );
or ( n29613 , n29555 , n29612 );
and ( n29614 , n29517 , n29613 );
or ( n29615 , n29516 , n29614 );
and ( n29616 , n29499 , n29615 );
or ( n29617 , n29498 , n29616 );
and ( n29618 , n29481 , n29617 );
or ( n29619 , n29480 , n29618 );
and ( n29620 , n29432 , n29619 );
or ( n29621 , n29431 , n29620 );
and ( n29622 , n29404 , n29621 );
or ( n29623 , n29403 , n29622 );
and ( n29624 , n29376 , n29623 );
or ( n29625 , n29375 , n29624 );
and ( n29626 , n29317 , n29625 );
or ( n29627 , n29316 , n29626 );
and ( n29628 , n29279 , n29627 );
or ( n29629 , n29278 , n29628 );
and ( n29630 , n29243 , n29629 );
or ( n29631 , n29242 , n29630 );
and ( n29632 , n29174 , n29631 );
or ( n29633 , n29173 , n29632 );
and ( n29634 , n29126 , n29633 );
or ( n29635 , n29125 , n29634 );
and ( n29636 , n29080 , n29635 );
or ( n29637 , n29079 , n29636 );
and ( n29638 , n29001 , n29637 );
or ( n29639 , n29000 , n29638 );
and ( n29640 , n28923 , n29639 );
or ( n29641 , n28922 , n29640 );
and ( n29642 , n28889 , n29641 );
or ( n29643 , n28888 , n29642 );
and ( n29644 , n28768 , n29643 );
or ( n29645 , n28767 , n29644 );
and ( n29646 , n28700 , n29645 );
or ( n29647 , n28699 , n29646 );
and ( n29648 , n28601 , n29647 );
or ( n29649 , n28600 , n29648 );
and ( n29650 , n28535 , n29649 );
or ( n29651 , n28534 , n29650 );
and ( n29652 , n28449 , n29651 );
or ( n29653 , n28448 , n29652 );
and ( n29654 , n28308 , n29653 );
or ( n29655 , n28307 , n29654 );
and ( n29656 , n28244 , n29655 );
or ( n29657 , n28243 , n29656 );
and ( n29658 , n28178 , n29657 );
or ( n29659 , n28177 , n29658 );
and ( n29660 , n28172 , n29659 );
or ( n29661 , n28171 , n29660 );
and ( n29662 , n27824 , n29661 );
or ( n29663 , n27823 , n29662 );
and ( n29664 , n27720 , n29663 );
or ( n29665 , n27719 , n29664 );
and ( n29666 , n27501 , n29665 );
or ( n29667 , n27500 , n29666 );
and ( n29668 , n27331 , n29667 );
or ( n29669 , n27330 , n29668 );
and ( n29670 , n27285 , n29669 );
or ( n29671 , n27284 , n29670 );
and ( n29672 , n27271 , n29671 );
and ( n29673 , n27269 , n29672 );
or ( n29674 , n27268 , n29673 );
and ( n29675 , n27263 , n29674 );
or ( n29676 , n27262 , n29675 );
and ( n29677 , n27005 , n29676 );
and ( n29678 , n27003 , n29677 );
and ( n29679 , n27001 , n29678 );
and ( n29680 , n26999 , n29679 );
and ( n29681 , n26997 , n29680 );
or ( n29682 , n26996 , n29681 );
and ( n29683 , n26172 , n29682 );
or ( n29684 , n26171 , n29683 );
and ( n29685 , n25719 , n29684 );
and ( n29686 , n25717 , n29685 );
and ( n29687 , n25715 , n29686 );
and ( n29688 , n25713 , n29687 );
or ( n29689 , n25712 , n29688 );
and ( n29690 , n25252 , n29689 );
or ( n29691 , n25251 , n29690 );
and ( n29692 , n24889 , n29691 );
and ( n29693 , n24887 , n29692 );
or ( n29694 , n24886 , n29693 );
and ( n29695 , n24724 , n29694 );
or ( n29696 , n24723 , n29695 );
and ( n29697 , n24355 , n29696 );
and ( n29698 , n24353 , n29697 );
or ( n29699 , n24352 , n29698 );
and ( n29700 , n24140 , n29699 );
or ( n29701 , n24139 , n29700 );
and ( n29702 , n23860 , n29701 );
and ( n29703 , n23858 , n29702 );
and ( n29704 , n23856 , n29703 );
and ( n29705 , n23854 , n29704 );
and ( n29706 , n23852 , n29705 );
and ( n29707 , n23850 , n29706 );
xor ( n29708 , n23848 , n29707 );
buf ( n29709 , n29708 );
buf ( n29710 , n29709 );
xor ( n29711 , n23850 , n29706 );
buf ( n29712 , n29711 );
buf ( n29713 , n29712 );
xor ( n29714 , n23852 , n29705 );
buf ( n29715 , n29714 );
buf ( n29716 , n29715 );
xor ( n29717 , n23854 , n29704 );
buf ( n29718 , n29717 );
buf ( n29719 , n29718 );
xor ( n29720 , n23856 , n29703 );
buf ( n29721 , n29720 );
buf ( n29722 , n29721 );
xor ( n29723 , n23858 , n29702 );
buf ( n29724 , n29723 );
buf ( n29725 , n29724 );
xor ( n29726 , n23860 , n29701 );
buf ( n29727 , n29726 );
buf ( n29728 , n29727 );
xor ( n29729 , n24140 , n29699 );
buf ( n29730 , n29729 );
buf ( n29731 , n29730 );
xor ( n29732 , n24353 , n29697 );
buf ( n29733 , n29732 );
buf ( n29734 , n29733 );
xor ( n29735 , n24355 , n29696 );
buf ( n29736 , n29735 );
buf ( n29737 , n29736 );
xor ( n29738 , n24724 , n29694 );
buf ( n29739 , n29738 );
buf ( n29740 , n29739 );
xor ( n29741 , n24887 , n29692 );
buf ( n29742 , n29741 );
buf ( n29743 , n29742 );
xor ( n29744 , n24889 , n29691 );
buf ( n29745 , n29744 );
buf ( n29746 , n29745 );
xor ( n29747 , n25252 , n29689 );
buf ( n29748 , n29747 );
buf ( n29749 , n29748 );
xor ( n29750 , n25713 , n29687 );
buf ( n29751 , n29750 );
buf ( n29752 , n29751 );
xor ( n29753 , n25715 , n29686 );
buf ( n29754 , n29753 );
buf ( n29755 , n29754 );
xor ( n29756 , n25717 , n29685 );
buf ( n29757 , n29756 );
buf ( n29758 , n29757 );
xor ( n29759 , n25719 , n29684 );
buf ( n29760 , n29759 );
buf ( n29761 , n29760 );
xor ( n29762 , n26172 , n29682 );
buf ( n29763 , n29762 );
buf ( n29764 , n29763 );
xor ( n29765 , n26997 , n29680 );
buf ( n29766 , n29765 );
buf ( n29767 , n29766 );
xor ( n29768 , n26999 , n29679 );
buf ( n29769 , n29768 );
buf ( n29770 , n29769 );
xor ( n29771 , n27001 , n29678 );
buf ( n29772 , n29771 );
buf ( n29773 , n29772 );
xor ( n29774 , n27003 , n29677 );
buf ( n29775 , n29774 );
buf ( n29776 , n29775 );
xor ( n29777 , n27005 , n29676 );
buf ( n29778 , n29777 );
buf ( n29779 , n29778 );
xor ( n29780 , n27263 , n29674 );
buf ( n29781 , n29780 );
buf ( n29782 , n29781 );
xor ( n29783 , n27269 , n29672 );
buf ( n29784 , n29783 );
buf ( n29785 , n29784 );
xor ( n29786 , n27271 , n29671 );
buf ( n29787 , n29786 );
buf ( n29788 , n29787 );
xor ( n29789 , n27285 , n29669 );
buf ( n29790 , n29789 );
buf ( n29791 , n29790 );
xor ( n29792 , n27331 , n29667 );
buf ( n29793 , n29792 );
buf ( n29794 , n29793 );
xor ( n29795 , n27501 , n29665 );
buf ( n29796 , n29795 );
buf ( n29797 , n29796 );
xor ( n29798 , n27720 , n29663 );
buf ( n29799 , n29798 );
buf ( n29800 , n29799 );
xor ( n29801 , n27824 , n29661 );
buf ( n29802 , n29801 );
buf ( n29803 , n29802 );
xor ( n29804 , n28172 , n29659 );
buf ( n29805 , n29804 );
buf ( n29806 , n29805 );
xor ( n29807 , n28178 , n29657 );
buf ( n29808 , n29807 );
buf ( n29809 , n29808 );
xor ( n29810 , n28244 , n29655 );
buf ( n29811 , n29810 );
buf ( n29812 , n29811 );
xor ( n29813 , n28308 , n29653 );
buf ( n29814 , n29813 );
buf ( n29815 , n29814 );
xor ( n29816 , n28449 , n29651 );
buf ( n29817 , n29816 );
buf ( n29818 , n29817 );
xor ( n29819 , n28535 , n29649 );
buf ( n29820 , n29819 );
buf ( n29821 , n29820 );
xor ( n29822 , n28601 , n29647 );
buf ( n29823 , n29822 );
buf ( n29824 , n29823 );
xor ( n29825 , n28700 , n29645 );
buf ( n29826 , n29825 );
buf ( n29827 , n29826 );
xor ( n29828 , n28768 , n29643 );
buf ( n29829 , n29828 );
buf ( n29830 , n29829 );
xor ( n29831 , n28889 , n29641 );
buf ( n29832 , n29831 );
buf ( n29833 , n29832 );
xor ( n29834 , n28923 , n29639 );
buf ( n29835 , n29834 );
buf ( n29836 , n29835 );
xor ( n29837 , n29001 , n29637 );
buf ( n29838 , n29837 );
buf ( n29839 , n29838 );
xor ( n29840 , n29080 , n29635 );
buf ( n29841 , n29840 );
buf ( n29842 , n29841 );
xor ( n29843 , n29126 , n29633 );
buf ( n29844 , n29843 );
buf ( n29845 , n29844 );
xor ( n29846 , n29174 , n29631 );
buf ( n29847 , n29846 );
buf ( n29848 , n29847 );
xor ( n29849 , n29243 , n29629 );
buf ( n29850 , n29849 );
buf ( n29851 , n29850 );
xor ( n29852 , n29279 , n29627 );
buf ( n29853 , n29852 );
buf ( n29854 , n29853 );
xor ( n29855 , n29317 , n29625 );
buf ( n29856 , n29855 );
buf ( n29857 , n29856 );
xor ( n29858 , n29376 , n29623 );
buf ( n29859 , n29858 );
buf ( n29860 , n29859 );
xor ( n29861 , n29404 , n29621 );
buf ( n29862 , n29861 );
buf ( n29863 , n29862 );
xor ( n29864 , n29432 , n29619 );
buf ( n29865 , n29864 );
buf ( n29866 , n29865 );
xor ( n29867 , n29481 , n29617 );
buf ( n29868 , n29867 );
buf ( n29869 , n29868 );
xor ( n29870 , n29499 , n29615 );
buf ( n29871 , n29870 );
buf ( n29872 , n29871 );
xor ( n29873 , n29517 , n29613 );
buf ( n29874 , n29873 );
buf ( n29875 , n29874 );
xor ( n29876 , n29556 , n29611 );
buf ( n29877 , n29876 );
buf ( n29878 , n29877 );
xor ( n29879 , n29564 , n29609 );
buf ( n29880 , n29879 );
buf ( n29881 , n29880 );
xor ( n29882 , n29572 , n29607 );
buf ( n29883 , n29882 );
buf ( n29884 , n29883 );
xor ( n29885 , n29580 , n29605 );
buf ( n29886 , n29885 );
buf ( n29887 , n29886 );
xor ( n29888 , n29587 , n29603 );
buf ( n29889 , n29888 );
buf ( n29890 , n29889 );
xor ( n29891 , n29593 , n29601 );
buf ( n29892 , n29891 );
buf ( n29893 , n29892 );
xor ( n29894 , n29597 , n29600 );
buf ( n29895 , n29894 );
buf ( n29896 , n29895 );
buf ( n29897 , n29598 );
buf ( n29898 , n29897 );
buf ( n29899 , n29898 );
and ( n29900 , n15770 , n29710 );
and ( n29901 , n15773 , n29713 );
and ( n29902 , n15776 , n29716 );
and ( n29903 , n15779 , n29719 );
and ( n29904 , n15782 , n29722 );
and ( n29905 , n15785 , n29725 );
and ( n29906 , n15788 , n29728 );
and ( n29907 , n15791 , n29731 );
and ( n29908 , n15794 , n29734 );
and ( n29909 , n15797 , n29737 );
and ( n29910 , n15800 , n29740 );
and ( n29911 , n15803 , n29743 );
and ( n29912 , n15806 , n29746 );
and ( n29913 , n15809 , n29749 );
and ( n29914 , n15812 , n29752 );
and ( n29915 , n15815 , n29755 );
and ( n29916 , n15818 , n29758 );
and ( n29917 , n15821 , n29761 );
and ( n29918 , n15824 , n29764 );
and ( n29919 , n15827 , n29767 );
and ( n29920 , n15830 , n29770 );
and ( n29921 , n15833 , n29773 );
and ( n29922 , n15836 , n29776 );
and ( n29923 , n15839 , n29779 );
and ( n29924 , n15842 , n29782 );
and ( n29925 , n15845 , n29785 );
and ( n29926 , n15848 , n29788 );
and ( n29927 , n15851 , n29791 );
and ( n29928 , n15854 , n29794 );
and ( n29929 , n15857 , n29797 );
and ( n29930 , n15860 , n29800 );
and ( n29931 , n15863 , n29803 );
and ( n29932 , n15866 , n29806 );
and ( n29933 , n15869 , n29809 );
and ( n29934 , n15872 , n29812 );
and ( n29935 , n15875 , n29815 );
and ( n29936 , n15878 , n29818 );
and ( n29937 , n15881 , n29821 );
and ( n29938 , n15884 , n29824 );
and ( n29939 , n15887 , n29827 );
and ( n29940 , n15890 , n29830 );
and ( n29941 , n15893 , n29833 );
and ( n29942 , n15896 , n29836 );
and ( n29943 , n15899 , n29839 );
and ( n29944 , n15902 , n29842 );
and ( n29945 , n15905 , n29845 );
and ( n29946 , n15908 , n29848 );
and ( n29947 , n15911 , n29851 );
and ( n29948 , n15914 , n29854 );
and ( n29949 , n15917 , n29857 );
and ( n29950 , n15920 , n29860 );
and ( n29951 , n15923 , n29863 );
and ( n29952 , n15926 , n29866 );
and ( n29953 , n15929 , n29869 );
and ( n29954 , n15932 , n29872 );
and ( n29955 , n15935 , n29875 );
and ( n29956 , n15938 , n29878 );
and ( n29957 , n15941 , n29881 );
and ( n29958 , n15944 , n29884 );
and ( n29959 , n15947 , n29887 );
and ( n29960 , n15950 , n29890 );
and ( n29961 , n15953 , n29893 );
and ( n29962 , n15956 , n29896 );
and ( n29963 , n15959 , n29899 );
and ( n29964 , n29896 , n29963 );
and ( n29965 , n15956 , n29963 );
or ( n29966 , n29962 , n29964 , n29965 );
and ( n29967 , n29893 , n29966 );
and ( n29968 , n15953 , n29966 );
or ( n29969 , n29961 , n29967 , n29968 );
and ( n29970 , n29890 , n29969 );
and ( n29971 , n15950 , n29969 );
or ( n29972 , n29960 , n29970 , n29971 );
and ( n29973 , n29887 , n29972 );
and ( n29974 , n15947 , n29972 );
or ( n29975 , n29959 , n29973 , n29974 );
and ( n29976 , n29884 , n29975 );
and ( n29977 , n15944 , n29975 );
or ( n29978 , n29958 , n29976 , n29977 );
and ( n29979 , n29881 , n29978 );
and ( n29980 , n15941 , n29978 );
or ( n29981 , n29957 , n29979 , n29980 );
and ( n29982 , n29878 , n29981 );
and ( n29983 , n15938 , n29981 );
or ( n29984 , n29956 , n29982 , n29983 );
and ( n29985 , n29875 , n29984 );
and ( n29986 , n15935 , n29984 );
or ( n29987 , n29955 , n29985 , n29986 );
and ( n29988 , n29872 , n29987 );
and ( n29989 , n15932 , n29987 );
or ( n29990 , n29954 , n29988 , n29989 );
and ( n29991 , n29869 , n29990 );
and ( n29992 , n15929 , n29990 );
or ( n29993 , n29953 , n29991 , n29992 );
and ( n29994 , n29866 , n29993 );
and ( n29995 , n15926 , n29993 );
or ( n29996 , n29952 , n29994 , n29995 );
and ( n29997 , n29863 , n29996 );
and ( n29998 , n15923 , n29996 );
or ( n29999 , n29951 , n29997 , n29998 );
and ( n30000 , n29860 , n29999 );
and ( n30001 , n15920 , n29999 );
or ( n30002 , n29950 , n30000 , n30001 );
and ( n30003 , n29857 , n30002 );
and ( n30004 , n15917 , n30002 );
or ( n30005 , n29949 , n30003 , n30004 );
and ( n30006 , n29854 , n30005 );
and ( n30007 , n15914 , n30005 );
or ( n30008 , n29948 , n30006 , n30007 );
and ( n30009 , n29851 , n30008 );
and ( n30010 , n15911 , n30008 );
or ( n30011 , n29947 , n30009 , n30010 );
and ( n30012 , n29848 , n30011 );
and ( n30013 , n15908 , n30011 );
or ( n30014 , n29946 , n30012 , n30013 );
and ( n30015 , n29845 , n30014 );
and ( n30016 , n15905 , n30014 );
or ( n30017 , n29945 , n30015 , n30016 );
and ( n30018 , n29842 , n30017 );
and ( n30019 , n15902 , n30017 );
or ( n30020 , n29944 , n30018 , n30019 );
and ( n30021 , n29839 , n30020 );
and ( n30022 , n15899 , n30020 );
or ( n30023 , n29943 , n30021 , n30022 );
and ( n30024 , n29836 , n30023 );
and ( n30025 , n15896 , n30023 );
or ( n30026 , n29942 , n30024 , n30025 );
and ( n30027 , n29833 , n30026 );
and ( n30028 , n15893 , n30026 );
or ( n30029 , n29941 , n30027 , n30028 );
and ( n30030 , n29830 , n30029 );
and ( n30031 , n15890 , n30029 );
or ( n30032 , n29940 , n30030 , n30031 );
and ( n30033 , n29827 , n30032 );
and ( n30034 , n15887 , n30032 );
or ( n30035 , n29939 , n30033 , n30034 );
and ( n30036 , n29824 , n30035 );
and ( n30037 , n15884 , n30035 );
or ( n30038 , n29938 , n30036 , n30037 );
and ( n30039 , n29821 , n30038 );
and ( n30040 , n15881 , n30038 );
or ( n30041 , n29937 , n30039 , n30040 );
and ( n30042 , n29818 , n30041 );
and ( n30043 , n15878 , n30041 );
or ( n30044 , n29936 , n30042 , n30043 );
and ( n30045 , n29815 , n30044 );
and ( n30046 , n15875 , n30044 );
or ( n30047 , n29935 , n30045 , n30046 );
and ( n30048 , n29812 , n30047 );
and ( n30049 , n15872 , n30047 );
or ( n30050 , n29934 , n30048 , n30049 );
and ( n30051 , n29809 , n30050 );
and ( n30052 , n15869 , n30050 );
or ( n30053 , n29933 , n30051 , n30052 );
and ( n30054 , n29806 , n30053 );
and ( n30055 , n15866 , n30053 );
or ( n30056 , n29932 , n30054 , n30055 );
and ( n30057 , n29803 , n30056 );
and ( n30058 , n15863 , n30056 );
or ( n30059 , n29931 , n30057 , n30058 );
and ( n30060 , n29800 , n30059 );
and ( n30061 , n15860 , n30059 );
or ( n30062 , n29930 , n30060 , n30061 );
and ( n30063 , n29797 , n30062 );
and ( n30064 , n15857 , n30062 );
or ( n30065 , n29929 , n30063 , n30064 );
and ( n30066 , n29794 , n30065 );
and ( n30067 , n15854 , n30065 );
or ( n30068 , n29928 , n30066 , n30067 );
and ( n30069 , n29791 , n30068 );
and ( n30070 , n15851 , n30068 );
or ( n30071 , n29927 , n30069 , n30070 );
and ( n30072 , n29788 , n30071 );
and ( n30073 , n15848 , n30071 );
or ( n30074 , n29926 , n30072 , n30073 );
and ( n30075 , n29785 , n30074 );
and ( n30076 , n15845 , n30074 );
or ( n30077 , n29925 , n30075 , n30076 );
and ( n30078 , n29782 , n30077 );
and ( n30079 , n15842 , n30077 );
or ( n30080 , n29924 , n30078 , n30079 );
and ( n30081 , n29779 , n30080 );
and ( n30082 , n15839 , n30080 );
or ( n30083 , n29923 , n30081 , n30082 );
and ( n30084 , n29776 , n30083 );
and ( n30085 , n15836 , n30083 );
or ( n30086 , n29922 , n30084 , n30085 );
and ( n30087 , n29773 , n30086 );
and ( n30088 , n15833 , n30086 );
or ( n30089 , n29921 , n30087 , n30088 );
and ( n30090 , n29770 , n30089 );
and ( n30091 , n15830 , n30089 );
or ( n30092 , n29920 , n30090 , n30091 );
and ( n30093 , n29767 , n30092 );
and ( n30094 , n15827 , n30092 );
or ( n30095 , n29919 , n30093 , n30094 );
and ( n30096 , n29764 , n30095 );
and ( n30097 , n15824 , n30095 );
or ( n30098 , n29918 , n30096 , n30097 );
and ( n30099 , n29761 , n30098 );
and ( n30100 , n15821 , n30098 );
or ( n30101 , n29917 , n30099 , n30100 );
and ( n30102 , n29758 , n30101 );
and ( n30103 , n15818 , n30101 );
or ( n30104 , n29916 , n30102 , n30103 );
and ( n30105 , n29755 , n30104 );
and ( n30106 , n15815 , n30104 );
or ( n30107 , n29915 , n30105 , n30106 );
and ( n30108 , n29752 , n30107 );
and ( n30109 , n15812 , n30107 );
or ( n30110 , n29914 , n30108 , n30109 );
and ( n30111 , n29749 , n30110 );
and ( n30112 , n15809 , n30110 );
or ( n30113 , n29913 , n30111 , n30112 );
and ( n30114 , n29746 , n30113 );
and ( n30115 , n15806 , n30113 );
or ( n30116 , n29912 , n30114 , n30115 );
and ( n30117 , n29743 , n30116 );
and ( n30118 , n15803 , n30116 );
or ( n30119 , n29911 , n30117 , n30118 );
and ( n30120 , n29740 , n30119 );
and ( n30121 , n15800 , n30119 );
or ( n30122 , n29910 , n30120 , n30121 );
and ( n30123 , n29737 , n30122 );
and ( n30124 , n15797 , n30122 );
or ( n30125 , n29909 , n30123 , n30124 );
and ( n30126 , n29734 , n30125 );
and ( n30127 , n15794 , n30125 );
or ( n30128 , n29908 , n30126 , n30127 );
and ( n30129 , n29731 , n30128 );
and ( n30130 , n15791 , n30128 );
or ( n30131 , n29907 , n30129 , n30130 );
and ( n30132 , n29728 , n30131 );
and ( n30133 , n15788 , n30131 );
or ( n30134 , n29906 , n30132 , n30133 );
and ( n30135 , n29725 , n30134 );
and ( n30136 , n15785 , n30134 );
or ( n30137 , n29905 , n30135 , n30136 );
and ( n30138 , n29722 , n30137 );
and ( n30139 , n15782 , n30137 );
or ( n30140 , n29904 , n30138 , n30139 );
and ( n30141 , n29719 , n30140 );
and ( n30142 , n15779 , n30140 );
or ( n30143 , n29903 , n30141 , n30142 );
and ( n30144 , n29716 , n30143 );
and ( n30145 , n15776 , n30143 );
or ( n30146 , n29902 , n30144 , n30145 );
and ( n30147 , n29713 , n30146 );
and ( n30148 , n15773 , n30146 );
or ( n30149 , n29901 , n30147 , n30148 );
and ( n30150 , n29710 , n30149 );
and ( n30151 , n15770 , n30149 );
or ( n30152 , n29900 , n30150 , n30151 );
buf ( n30153 , n30152 );
xor ( n30154 , n15770 , n29710 );
xor ( n30155 , n30154 , n30149 );
buf ( n30156 , n30155 );
xor ( n30157 , n15773 , n29713 );
xor ( n30158 , n30157 , n30146 );
buf ( n30159 , n30158 );
xor ( n30160 , n15776 , n29716 );
xor ( n30161 , n30160 , n30143 );
buf ( n30162 , n30161 );
xor ( n30163 , n15779 , n29719 );
xor ( n30164 , n30163 , n30140 );
buf ( n30165 , n30164 );
xor ( n30166 , n15782 , n29722 );
xor ( n30167 , n30166 , n30137 );
buf ( n30168 , n30167 );
xor ( n30169 , n15785 , n29725 );
xor ( n30170 , n30169 , n30134 );
buf ( n30171 , n30170 );
xor ( n30172 , n15788 , n29728 );
xor ( n30173 , n30172 , n30131 );
buf ( n30174 , n30173 );
xor ( n30175 , n15791 , n29731 );
xor ( n30176 , n30175 , n30128 );
buf ( n30177 , n30176 );
xor ( n30178 , n15794 , n29734 );
xor ( n30179 , n30178 , n30125 );
buf ( n30180 , n30179 );
xor ( n30181 , n15797 , n29737 );
xor ( n30182 , n30181 , n30122 );
buf ( n30183 , n30182 );
xor ( n30184 , n15800 , n29740 );
xor ( n30185 , n30184 , n30119 );
buf ( n30186 , n30185 );
xor ( n30187 , n15803 , n29743 );
xor ( n30188 , n30187 , n30116 );
buf ( n30189 , n30188 );
xor ( n30190 , n15806 , n29746 );
xor ( n30191 , n30190 , n30113 );
buf ( n30192 , n30191 );
xor ( n30193 , n15809 , n29749 );
xor ( n30194 , n30193 , n30110 );
buf ( n30195 , n30194 );
xor ( n30196 , n15812 , n29752 );
xor ( n30197 , n30196 , n30107 );
buf ( n30198 , n30197 );
xor ( n30199 , n15815 , n29755 );
xor ( n30200 , n30199 , n30104 );
buf ( n30201 , n30200 );
xor ( n30202 , n15818 , n29758 );
xor ( n30203 , n30202 , n30101 );
buf ( n30204 , n30203 );
xor ( n30205 , n15821 , n29761 );
xor ( n30206 , n30205 , n30098 );
buf ( n30207 , n30206 );
xor ( n30208 , n15824 , n29764 );
xor ( n30209 , n30208 , n30095 );
buf ( n30210 , n30209 );
xor ( n30211 , n15827 , n29767 );
xor ( n30212 , n30211 , n30092 );
buf ( n30213 , n30212 );
xor ( n30214 , n15830 , n29770 );
xor ( n30215 , n30214 , n30089 );
buf ( n30216 , n30215 );
xor ( n30217 , n15833 , n29773 );
xor ( n30218 , n30217 , n30086 );
buf ( n30219 , n30218 );
xor ( n30220 , n15836 , n29776 );
xor ( n30221 , n30220 , n30083 );
buf ( n30222 , n30221 );
xor ( n30223 , n15839 , n29779 );
xor ( n30224 , n30223 , n30080 );
buf ( n30225 , n30224 );
xor ( n30226 , n15842 , n29782 );
xor ( n30227 , n30226 , n30077 );
buf ( n30228 , n30227 );
xor ( n30229 , n15845 , n29785 );
xor ( n30230 , n30229 , n30074 );
buf ( n30231 , n30230 );
xor ( n30232 , n15848 , n29788 );
xor ( n30233 , n30232 , n30071 );
buf ( n30234 , n30233 );
xor ( n30235 , n15851 , n29791 );
xor ( n30236 , n30235 , n30068 );
buf ( n30237 , n30236 );
xor ( n30238 , n15854 , n29794 );
xor ( n30239 , n30238 , n30065 );
buf ( n30240 , n30239 );
xor ( n30241 , n15857 , n29797 );
xor ( n30242 , n30241 , n30062 );
buf ( n30243 , n30242 );
xor ( n30244 , n15860 , n29800 );
xor ( n30245 , n30244 , n30059 );
buf ( n30246 , n30245 );
xor ( n30247 , n15863 , n29803 );
xor ( n30248 , n30247 , n30056 );
buf ( n30249 , n30248 );
xor ( n30250 , n15866 , n29806 );
xor ( n30251 , n30250 , n30053 );
buf ( n30252 , n30251 );
xor ( n30253 , n15869 , n29809 );
xor ( n30254 , n30253 , n30050 );
buf ( n30255 , n30254 );
xor ( n30256 , n15872 , n29812 );
xor ( n30257 , n30256 , n30047 );
buf ( n30258 , n30257 );
xor ( n30259 , n15875 , n29815 );
xor ( n30260 , n30259 , n30044 );
buf ( n30261 , n30260 );
xor ( n30262 , n15878 , n29818 );
xor ( n30263 , n30262 , n30041 );
buf ( n30264 , n30263 );
xor ( n30265 , n15881 , n29821 );
xor ( n30266 , n30265 , n30038 );
buf ( n30267 , n30266 );
xor ( n30268 , n15884 , n29824 );
xor ( n30269 , n30268 , n30035 );
buf ( n30270 , n30269 );
xor ( n30271 , n15887 , n29827 );
xor ( n30272 , n30271 , n30032 );
buf ( n30273 , n30272 );
xor ( n30274 , n15890 , n29830 );
xor ( n30275 , n30274 , n30029 );
buf ( n30276 , n30275 );
xor ( n30277 , n15893 , n29833 );
xor ( n30278 , n30277 , n30026 );
buf ( n30279 , n30278 );
xor ( n30280 , n15896 , n29836 );
xor ( n30281 , n30280 , n30023 );
buf ( n30282 , n30281 );
xor ( n30283 , n15899 , n29839 );
xor ( n30284 , n30283 , n30020 );
buf ( n30285 , n30284 );
xor ( n30286 , n15902 , n29842 );
xor ( n30287 , n30286 , n30017 );
buf ( n30288 , n30287 );
xor ( n30289 , n15905 , n29845 );
xor ( n30290 , n30289 , n30014 );
buf ( n30291 , n30290 );
xor ( n30292 , n15908 , n29848 );
xor ( n30293 , n30292 , n30011 );
buf ( n30294 , n30293 );
xor ( n30295 , n15911 , n29851 );
xor ( n30296 , n30295 , n30008 );
buf ( n30297 , n30296 );
xor ( n30298 , n15914 , n29854 );
xor ( n30299 , n30298 , n30005 );
buf ( n30300 , n30299 );
xor ( n30301 , n15917 , n29857 );
xor ( n30302 , n30301 , n30002 );
buf ( n30303 , n30302 );
xor ( n30304 , n15920 , n29860 );
xor ( n30305 , n30304 , n29999 );
buf ( n30306 , n30305 );
xor ( n30307 , n15923 , n29863 );
xor ( n30308 , n30307 , n29996 );
buf ( n30309 , n30308 );
xor ( n30310 , n15926 , n29866 );
xor ( n30311 , n30310 , n29993 );
buf ( n30312 , n30311 );
xor ( n30313 , n15929 , n29869 );
xor ( n30314 , n30313 , n29990 );
buf ( n30315 , n30314 );
xor ( n30316 , n15932 , n29872 );
xor ( n30317 , n30316 , n29987 );
buf ( n30318 , n30317 );
xor ( n30319 , n15935 , n29875 );
xor ( n30320 , n30319 , n29984 );
buf ( n30321 , n30320 );
xor ( n30322 , n15938 , n29878 );
xor ( n30323 , n30322 , n29981 );
buf ( n30324 , n30323 );
xor ( n30325 , n15941 , n29881 );
xor ( n30326 , n30325 , n29978 );
buf ( n30327 , n30326 );
xor ( n30328 , n15944 , n29884 );
xor ( n30329 , n30328 , n29975 );
buf ( n30330 , n30329 );
xor ( n30331 , n15947 , n29887 );
xor ( n30332 , n30331 , n29972 );
buf ( n30333 , n30332 );
xor ( n30334 , n15950 , n29890 );
xor ( n30335 , n30334 , n29969 );
buf ( n30336 , n30335 );
xor ( n30337 , n15953 , n29893 );
xor ( n30338 , n30337 , n29966 );
buf ( n30339 , n30338 );
xor ( n30340 , n15956 , n29896 );
xor ( n30341 , n30340 , n29963 );
buf ( n30342 , n30341 );
xor ( n30343 , n15959 , n29899 );
buf ( n30344 , n30343 );
buf ( n30345 , n30153 );
buf ( n30346 , n30156 );
buf ( n30347 , n30159 );
buf ( n30348 , n30162 );
buf ( n30349 , n30165 );
buf ( n30350 , n30168 );
buf ( n30351 , n30171 );
buf ( n30352 , n30174 );
buf ( n30353 , n30177 );
buf ( n30354 , n30180 );
buf ( n30355 , n30183 );
buf ( n30356 , n30186 );
buf ( n30357 , n30189 );
buf ( n30358 , n30192 );
buf ( n30359 , n30195 );
buf ( n30360 , n30198 );
buf ( n30361 , n30201 );
buf ( n30362 , n30204 );
buf ( n30363 , n30207 );
buf ( n30364 , n30210 );
buf ( n30365 , n30213 );
buf ( n30366 , n30216 );
buf ( n30367 , n30219 );
buf ( n30368 , n30222 );
buf ( n30369 , n30225 );
buf ( n30370 , n30228 );
buf ( n30371 , n30231 );
buf ( n30372 , n30234 );
buf ( n30373 , n30237 );
buf ( n30374 , n30240 );
buf ( n30375 , n30243 );
buf ( n30376 , n30246 );
buf ( n30377 , n30249 );
buf ( n30378 , n30252 );
buf ( n30379 , n30255 );
buf ( n30380 , n30258 );
buf ( n30381 , n30261 );
buf ( n30382 , n30264 );
buf ( n30383 , n30267 );
buf ( n30384 , n30270 );
buf ( n30385 , n30273 );
buf ( n30386 , n30276 );
buf ( n30387 , n30279 );
buf ( n30388 , n30282 );
buf ( n30389 , n30285 );
buf ( n30390 , n30288 );
buf ( n30391 , n30291 );
buf ( n30392 , n30294 );
buf ( n30393 , n30297 );
buf ( n30394 , n30300 );
buf ( n30395 , n30303 );
buf ( n30396 , n30306 );
buf ( n30397 , n30309 );
buf ( n30398 , n30312 );
buf ( n30399 , n30315 );
buf ( n30400 , n30318 );
buf ( n30401 , n30321 );
buf ( n30402 , n30324 );
buf ( n30403 , n30327 );
buf ( n30404 , n30330 );
buf ( n30405 , n30333 );
buf ( n30406 , n30336 );
buf ( n30407 , n30339 );
buf ( n30408 , n30342 );
buf ( n30409 , n30344 );
buf ( n30410 , n15769 );
buf ( n30411 , n30410 );
buf ( n30412 , n1218 );
buf ( n30413 , n30412 );
buf ( n30414 , n30413 );
buf ( n30415 , n15772 );
buf ( n30416 , n30415 );
and ( n30417 , n30414 , n30416 );
buf ( n30418 , n1219 );
buf ( n30419 , n30418 );
buf ( n30420 , n1218 );
buf ( n30421 , n30420 );
and ( n30422 , n30419 , n30421 );
buf ( n30423 , n1219 );
buf ( n30424 , n30423 );
and ( n30425 , n30413 , n30424 );
and ( n30426 , n30422 , n30425 );
buf ( n30427 , n15775 );
buf ( n30428 , n30427 );
and ( n30429 , n30425 , n30428 );
and ( n30430 , n30422 , n30428 );
or ( n30431 , n30426 , n30429 , n30430 );
and ( n30432 , n30416 , n30431 );
and ( n30433 , n30414 , n30431 );
or ( n30434 , n30417 , n30432 , n30433 );
and ( n30435 , n30411 , n30434 );
xor ( n30436 , n30414 , n30416 );
xor ( n30437 , n30436 , n30431 );
buf ( n30438 , n1220 );
buf ( n30439 , n30438 );
and ( n30440 , n30413 , n30439 );
buf ( n30441 , n1220 );
buf ( n30442 , n30441 );
and ( n30443 , n30442 , n30421 );
and ( n30444 , n30440 , n30443 );
xor ( n30445 , n30422 , n30425 );
xor ( n30446 , n30445 , n30428 );
and ( n30447 , n30444 , n30446 );
buf ( n30448 , n30419 );
buf ( n30449 , n15778 );
buf ( n30450 , n30449 );
and ( n30451 , n30448 , n30450 );
xor ( n30452 , n30440 , n30443 );
and ( n30453 , n30450 , n30452 );
and ( n30454 , n30448 , n30452 );
or ( n30455 , n30451 , n30453 , n30454 );
and ( n30456 , n30446 , n30455 );
and ( n30457 , n30444 , n30455 );
or ( n30458 , n30447 , n30456 , n30457 );
and ( n30459 , n30437 , n30458 );
buf ( n30460 , n1221 );
buf ( n30461 , n30460 );
and ( n30462 , n30413 , n30461 );
buf ( n30463 , n1221 );
buf ( n30464 , n30463 );
and ( n30465 , n30464 , n30421 );
and ( n30466 , n30462 , n30465 );
buf ( n30467 , n1222 );
buf ( n30468 , n30467 );
and ( n30469 , n30468 , n30421 );
and ( n30470 , n30464 , n30424 );
or ( n30471 , n30469 , n30470 );
buf ( n30472 , n1222 );
buf ( n30473 , n30472 );
and ( n30474 , n30413 , n30473 );
and ( n30475 , n30419 , n30461 );
or ( n30476 , n30474 , n30475 );
and ( n30477 , n30471 , n30476 );
and ( n30478 , n30466 , n30477 );
and ( n30479 , n30442 , n30424 );
and ( n30480 , n30419 , n30439 );
and ( n30481 , n30479 , n30480 );
xor ( n30482 , n30462 , n30465 );
and ( n30483 , n30480 , n30482 );
and ( n30484 , n30479 , n30482 );
or ( n30485 , n30481 , n30483 , n30484 );
and ( n30486 , n30477 , n30485 );
and ( n30487 , n30466 , n30485 );
or ( n30488 , n30478 , n30486 , n30487 );
xor ( n30489 , n30444 , n30446 );
xor ( n30490 , n30489 , n30455 );
and ( n30491 , n30488 , n30490 );
xor ( n30492 , n30448 , n30450 );
xor ( n30493 , n30492 , n30452 );
xnor ( n30494 , n30469 , n30470 );
xnor ( n30495 , n30474 , n30475 );
and ( n30496 , n30494 , n30495 );
buf ( n30497 , n15781 );
buf ( n30498 , n30497 );
or ( n30499 , n30496 , n30498 );
and ( n30500 , n30493 , n30499 );
xor ( n30501 , n30471 , n30476 );
buf ( n30502 , n1223 );
buf ( n30503 , n30502 );
and ( n30504 , n30503 , n30421 );
and ( n30505 , n30468 , n30424 );
or ( n30506 , n30504 , n30505 );
buf ( n30507 , n1223 );
buf ( n30508 , n30507 );
and ( n30509 , n30413 , n30508 );
and ( n30510 , n30419 , n30473 );
or ( n30511 , n30509 , n30510 );
and ( n30512 , n30506 , n30511 );
and ( n30513 , n30501 , n30512 );
buf ( n30514 , n30442 );
buf ( n30515 , n15784 );
buf ( n30516 , n30515 );
and ( n30517 , n30514 , n30516 );
and ( n30518 , n30464 , n30439 );
and ( n30519 , n30442 , n30461 );
and ( n30520 , n30518 , n30519 );
buf ( n30521 , n15787 );
buf ( n30522 , n30521 );
and ( n30523 , n30519 , n30522 );
and ( n30524 , n30518 , n30522 );
or ( n30525 , n30520 , n30523 , n30524 );
and ( n30526 , n30516 , n30525 );
and ( n30527 , n30514 , n30525 );
or ( n30528 , n30517 , n30526 , n30527 );
and ( n30529 , n30512 , n30528 );
and ( n30530 , n30501 , n30528 );
or ( n30531 , n30513 , n30529 , n30530 );
and ( n30532 , n30499 , n30531 );
and ( n30533 , n30493 , n30531 );
or ( n30534 , n30500 , n30532 , n30533 );
and ( n30535 , n30490 , n30534 );
and ( n30536 , n30488 , n30534 );
or ( n30537 , n30491 , n30535 , n30536 );
and ( n30538 , n30458 , n30537 );
and ( n30539 , n30437 , n30537 );
or ( n30540 , n30459 , n30538 , n30539 );
and ( n30541 , n30434 , n30540 );
and ( n30542 , n30411 , n30540 );
or ( n30543 , n30435 , n30541 , n30542 );
xor ( n30544 , n30411 , n30434 );
xor ( n30545 , n30544 , n30540 );
xor ( n30546 , n30437 , n30458 );
xor ( n30547 , n30546 , n30537 );
xor ( n30548 , n30466 , n30477 );
xor ( n30549 , n30548 , n30485 );
xor ( n30550 , n30479 , n30480 );
xor ( n30551 , n30550 , n30482 );
xnor ( n30552 , n30496 , n30498 );
and ( n30553 , n30551 , n30552 );
xor ( n30554 , n30506 , n30511 );
xor ( n30555 , n30494 , n30495 );
and ( n30556 , n30554 , n30555 );
buf ( n30557 , n1224 );
buf ( n30558 , n30557 );
and ( n30559 , n30558 , n30421 );
and ( n30560 , n30468 , n30439 );
or ( n30561 , n30559 , n30560 );
buf ( n30562 , n1224 );
buf ( n30563 , n30562 );
and ( n30564 , n30413 , n30563 );
and ( n30565 , n30442 , n30473 );
or ( n30566 , n30564 , n30565 );
and ( n30567 , n30561 , n30566 );
and ( n30568 , n30555 , n30567 );
and ( n30569 , n30554 , n30567 );
or ( n30570 , n30556 , n30568 , n30569 );
and ( n30571 , n30552 , n30570 );
and ( n30572 , n30551 , n30570 );
or ( n30573 , n30553 , n30571 , n30572 );
and ( n30574 , n30549 , n30573 );
xor ( n30575 , n30493 , n30499 );
xor ( n30576 , n30575 , n30531 );
and ( n30577 , n30573 , n30576 );
and ( n30578 , n30549 , n30576 );
or ( n30579 , n30574 , n30577 , n30578 );
xor ( n30580 , n30488 , n30490 );
xor ( n30581 , n30580 , n30534 );
and ( n30582 , n30579 , n30581 );
xor ( n30583 , n30501 , n30512 );
xor ( n30584 , n30583 , n30528 );
xnor ( n30585 , n30504 , n30505 );
xnor ( n30586 , n30509 , n30510 );
and ( n30587 , n30585 , n30586 );
xor ( n30588 , n30514 , n30516 );
xor ( n30589 , n30588 , n30525 );
and ( n30590 , n30587 , n30589 );
buf ( n30591 , n1225 );
buf ( n30592 , n30591 );
and ( n30593 , n30413 , n30592 );
and ( n30594 , n30419 , n30563 );
and ( n30595 , n30593 , n30594 );
and ( n30596 , n30442 , n30508 );
and ( n30597 , n30594 , n30596 );
and ( n30598 , n30593 , n30596 );
or ( n30599 , n30595 , n30597 , n30598 );
and ( n30600 , n30503 , n30424 );
and ( n30601 , n30599 , n30600 );
buf ( n30602 , n1225 );
buf ( n30603 , n30602 );
and ( n30604 , n30603 , n30421 );
and ( n30605 , n30558 , n30424 );
and ( n30606 , n30604 , n30605 );
and ( n30607 , n30503 , n30439 );
and ( n30608 , n30605 , n30607 );
and ( n30609 , n30604 , n30607 );
or ( n30610 , n30606 , n30608 , n30609 );
and ( n30611 , n30419 , n30508 );
and ( n30612 , n30610 , n30611 );
and ( n30613 , n30601 , n30612 );
and ( n30614 , n30589 , n30613 );
and ( n30615 , n30587 , n30613 );
or ( n30616 , n30590 , n30614 , n30615 );
and ( n30617 , n30584 , n30616 );
xor ( n30618 , n30551 , n30552 );
xor ( n30619 , n30618 , n30570 );
and ( n30620 , n30616 , n30619 );
and ( n30621 , n30584 , n30619 );
or ( n30622 , n30617 , n30620 , n30621 );
xor ( n30623 , n30549 , n30573 );
xor ( n30624 , n30623 , n30576 );
and ( n30625 , n30622 , n30624 );
xor ( n30626 , n30518 , n30519 );
xor ( n30627 , n30626 , n30522 );
xor ( n30628 , n30561 , n30566 );
and ( n30629 , n30627 , n30628 );
xor ( n30630 , n30585 , n30586 );
and ( n30631 , n30628 , n30630 );
and ( n30632 , n30627 , n30630 );
or ( n30633 , n30629 , n30631 , n30632 );
xor ( n30634 , n30554 , n30555 );
xor ( n30635 , n30634 , n30567 );
and ( n30636 , n30633 , n30635 );
xnor ( n30637 , n30559 , n30560 );
xnor ( n30638 , n30564 , n30565 );
and ( n30639 , n30637 , n30638 );
buf ( n30640 , n30464 );
buf ( n30641 , n15790 );
buf ( n30642 , n30641 );
and ( n30643 , n30640 , n30642 );
and ( n30644 , n30468 , n30461 );
and ( n30645 , n30464 , n30473 );
and ( n30646 , n30644 , n30645 );
buf ( n30647 , n15793 );
buf ( n30648 , n30647 );
and ( n30649 , n30645 , n30648 );
and ( n30650 , n30644 , n30648 );
or ( n30651 , n30646 , n30649 , n30650 );
and ( n30652 , n30642 , n30651 );
and ( n30653 , n30640 , n30651 );
or ( n30654 , n30643 , n30652 , n30653 );
and ( n30655 , n30639 , n30654 );
xor ( n30656 , n30601 , n30612 );
and ( n30657 , n30654 , n30656 );
and ( n30658 , n30639 , n30656 );
or ( n30659 , n30655 , n30657 , n30658 );
and ( n30660 , n30635 , n30659 );
and ( n30661 , n30633 , n30659 );
or ( n30662 , n30636 , n30660 , n30661 );
xor ( n30663 , n30584 , n30616 );
xor ( n30664 , n30663 , n30619 );
and ( n30665 , n30662 , n30664 );
xor ( n30666 , n30599 , n30600 );
xor ( n30667 , n30610 , n30611 );
and ( n30668 , n30666 , n30667 );
xor ( n30669 , n30637 , n30638 );
and ( n30670 , n30603 , n30424 );
and ( n30671 , n30503 , n30461 );
or ( n30672 , n30670 , n30671 );
and ( n30673 , n30419 , n30592 );
and ( n30674 , n30464 , n30508 );
or ( n30675 , n30673 , n30674 );
and ( n30676 , n30672 , n30675 );
and ( n30677 , n30669 , n30676 );
xor ( n30678 , n30604 , n30605 );
xor ( n30679 , n30678 , n30607 );
xor ( n30680 , n30593 , n30594 );
xor ( n30681 , n30680 , n30596 );
and ( n30682 , n30679 , n30681 );
and ( n30683 , n30676 , n30682 );
and ( n30684 , n30669 , n30682 );
or ( n30685 , n30677 , n30683 , n30684 );
and ( n30686 , n30668 , n30685 );
xor ( n30687 , n30627 , n30628 );
xor ( n30688 , n30687 , n30630 );
and ( n30689 , n30685 , n30688 );
and ( n30690 , n30668 , n30688 );
or ( n30691 , n30686 , n30689 , n30690 );
xor ( n30692 , n30587 , n30589 );
xor ( n30693 , n30692 , n30613 );
and ( n30694 , n30691 , n30693 );
xor ( n30695 , n30640 , n30642 );
xor ( n30696 , n30695 , n30651 );
xor ( n30697 , n30666 , n30667 );
and ( n30698 , n30696 , n30697 );
buf ( n30699 , n1226 );
buf ( n30700 , n30699 );
and ( n30701 , n30419 , n30700 );
and ( n30702 , n30442 , n30592 );
and ( n30703 , n30701 , n30702 );
and ( n30704 , n30464 , n30563 );
and ( n30705 , n30702 , n30704 );
and ( n30706 , n30701 , n30704 );
or ( n30707 , n30703 , n30705 , n30706 );
buf ( n30708 , n1226 );
buf ( n30709 , n30708 );
and ( n30710 , n30709 , n30421 );
and ( n30711 , n30707 , n30710 );
and ( n30712 , n30558 , n30439 );
and ( n30713 , n30710 , n30712 );
and ( n30714 , n30707 , n30712 );
or ( n30715 , n30711 , n30713 , n30714 );
and ( n30716 , n30709 , n30424 );
and ( n30717 , n30603 , n30439 );
and ( n30718 , n30716 , n30717 );
and ( n30719 , n30558 , n30461 );
and ( n30720 , n30717 , n30719 );
and ( n30721 , n30716 , n30719 );
or ( n30722 , n30718 , n30720 , n30721 );
and ( n30723 , n30413 , n30700 );
and ( n30724 , n30722 , n30723 );
and ( n30725 , n30442 , n30563 );
and ( n30726 , n30723 , n30725 );
and ( n30727 , n30722 , n30725 );
or ( n30728 , n30724 , n30726 , n30727 );
and ( n30729 , n30715 , n30728 );
and ( n30730 , n30697 , n30729 );
and ( n30731 , n30696 , n30729 );
or ( n30732 , n30698 , n30730 , n30731 );
xor ( n30733 , n30639 , n30654 );
xor ( n30734 , n30733 , n30656 );
and ( n30735 , n30732 , n30734 );
xor ( n30736 , n30668 , n30685 );
xor ( n30737 , n30736 , n30688 );
and ( n30738 , n30734 , n30737 );
and ( n30739 , n30732 , n30737 );
or ( n30740 , n30735 , n30738 , n30739 );
and ( n30741 , n30693 , n30740 );
and ( n30742 , n30691 , n30740 );
or ( n30743 , n30694 , n30741 , n30742 );
and ( n30744 , n30664 , n30743 );
and ( n30745 , n30662 , n30743 );
or ( n30746 , n30665 , n30744 , n30745 );
and ( n30747 , n30624 , n30746 );
and ( n30748 , n30622 , n30746 );
or ( n30749 , n30625 , n30747 , n30748 );
and ( n30750 , n30581 , n30749 );
and ( n30751 , n30579 , n30749 );
or ( n30752 , n30582 , n30750 , n30751 );
or ( n30753 , n30547 , n30752 );
or ( n30754 , n30545 , n30753 );
xor ( n30755 , n30543 , n30754 );
not ( n30756 , n30755 );
xnor ( n30757 , n30545 , n30753 );
xnor ( n30758 , n30547 , n30752 );
xor ( n30759 , n30579 , n30581 );
xor ( n30760 , n30759 , n30749 );
not ( n30761 , n30760 );
xor ( n30762 , n30622 , n30624 );
xor ( n30763 , n30762 , n30746 );
xor ( n30764 , n30662 , n30664 );
xor ( n30765 , n30764 , n30743 );
xor ( n30766 , n30633 , n30635 );
xor ( n30767 , n30766 , n30659 );
xor ( n30768 , n30691 , n30693 );
xor ( n30769 , n30768 , n30740 );
and ( n30770 , n30767 , n30769 );
xor ( n30771 , n30644 , n30645 );
xor ( n30772 , n30771 , n30648 );
xor ( n30773 , n30672 , n30675 );
and ( n30774 , n30772 , n30773 );
xor ( n30775 , n30679 , n30681 );
and ( n30776 , n30773 , n30775 );
and ( n30777 , n30772 , n30775 );
or ( n30778 , n30774 , n30776 , n30777 );
xor ( n30779 , n30669 , n30676 );
xor ( n30780 , n30779 , n30682 );
and ( n30781 , n30778 , n30780 );
xnor ( n30782 , n30670 , n30671 );
xnor ( n30783 , n30673 , n30674 );
and ( n30784 , n30782 , n30783 );
xor ( n30785 , n30715 , n30728 );
and ( n30786 , n30784 , n30785 );
buf ( n30787 , n1228 );
buf ( n30788 , n30787 );
and ( n30789 , n30413 , n30788 );
buf ( n30790 , n1227 );
buf ( n30791 , n30790 );
and ( n30792 , n30419 , n30791 );
and ( n30793 , n30789 , n30792 );
and ( n30794 , n30464 , n30592 );
and ( n30795 , n30792 , n30794 );
and ( n30796 , n30789 , n30794 );
or ( n30797 , n30793 , n30795 , n30796 );
buf ( n30798 , n1227 );
buf ( n30799 , n30798 );
and ( n30800 , n30799 , n30421 );
or ( n30801 , n30797 , n30800 );
buf ( n30802 , n1228 );
buf ( n30803 , n30802 );
and ( n30804 , n30803 , n30421 );
and ( n30805 , n30799 , n30424 );
and ( n30806 , n30804 , n30805 );
and ( n30807 , n30603 , n30461 );
and ( n30808 , n30805 , n30807 );
and ( n30809 , n30804 , n30807 );
or ( n30810 , n30806 , n30808 , n30809 );
and ( n30811 , n30413 , n30791 );
or ( n30812 , n30810 , n30811 );
and ( n30813 , n30801 , n30812 );
and ( n30814 , n30785 , n30813 );
and ( n30815 , n30784 , n30813 );
or ( n30816 , n30786 , n30814 , n30815 );
and ( n30817 , n30780 , n30816 );
and ( n30818 , n30778 , n30816 );
or ( n30819 , n30781 , n30817 , n30818 );
xor ( n30820 , n30732 , n30734 );
xor ( n30821 , n30820 , n30737 );
and ( n30822 , n30819 , n30821 );
xor ( n30823 , n30707 , n30710 );
xor ( n30824 , n30823 , n30712 );
xor ( n30825 , n30722 , n30723 );
xor ( n30826 , n30825 , n30725 );
and ( n30827 , n30824 , n30826 );
buf ( n30828 , n30468 );
buf ( n30829 , n15796 );
buf ( n30830 , n30829 );
and ( n30831 , n30828 , n30830 );
xor ( n30832 , n30782 , n30783 );
and ( n30833 , n30830 , n30832 );
and ( n30834 , n30828 , n30832 );
or ( n30835 , n30831 , n30833 , n30834 );
and ( n30836 , n30827 , n30835 );
xor ( n30837 , n30772 , n30773 );
xor ( n30838 , n30837 , n30775 );
and ( n30839 , n30835 , n30838 );
and ( n30840 , n30827 , n30838 );
or ( n30841 , n30836 , n30839 , n30840 );
xor ( n30842 , n30696 , n30697 );
xor ( n30843 , n30842 , n30729 );
and ( n30844 , n30841 , n30843 );
and ( n30845 , n30709 , n30439 );
and ( n30846 , n30558 , n30473 );
or ( n30847 , n30845 , n30846 );
and ( n30848 , n30442 , n30700 );
and ( n30849 , n30468 , n30563 );
or ( n30850 , n30848 , n30849 );
and ( n30851 , n30847 , n30850 );
xor ( n30852 , n30716 , n30717 );
xor ( n30853 , n30852 , n30719 );
xor ( n30854 , n30701 , n30702 );
xor ( n30855 , n30854 , n30704 );
and ( n30856 , n30853 , n30855 );
and ( n30857 , n30851 , n30856 );
xor ( n30858 , n30801 , n30812 );
and ( n30859 , n30856 , n30858 );
and ( n30860 , n30851 , n30858 );
or ( n30861 , n30857 , n30859 , n30860 );
xor ( n30862 , n30824 , n30826 );
xnor ( n30863 , n30845 , n30846 );
xnor ( n30864 , n30848 , n30849 );
and ( n30865 , n30863 , n30864 );
not ( n30866 , n30865 );
buf ( n30867 , n15799 );
buf ( n30868 , n30867 );
and ( n30869 , n30866 , n30868 );
and ( n30870 , n30862 , n30869 );
buf ( n30871 , n30865 );
and ( n30872 , n30869 , n30871 );
and ( n30873 , n30862 , n30871 );
or ( n30874 , n30870 , n30872 , n30873 );
and ( n30875 , n30861 , n30874 );
xnor ( n30876 , n30797 , n30800 );
xnor ( n30877 , n30810 , n30811 );
and ( n30878 , n30876 , n30877 );
and ( n30879 , n30503 , n30473 );
and ( n30880 , n30468 , n30508 );
and ( n30881 , n30879 , n30880 );
xor ( n30882 , n30847 , n30850 );
and ( n30883 , n30880 , n30882 );
and ( n30884 , n30879 , n30882 );
or ( n30885 , n30881 , n30883 , n30884 );
and ( n30886 , n30878 , n30885 );
xor ( n30887 , n30853 , n30855 );
buf ( n30888 , n1229 );
buf ( n30889 , n30888 );
and ( n30890 , n30889 , n30421 );
and ( n30891 , n30709 , n30461 );
and ( n30892 , n30890 , n30891 );
and ( n30893 , n30603 , n30473 );
and ( n30894 , n30891 , n30893 );
and ( n30895 , n30890 , n30893 );
or ( n30896 , n30892 , n30894 , n30895 );
buf ( n30897 , n1229 );
buf ( n30898 , n30897 );
and ( n30899 , n30413 , n30898 );
and ( n30900 , n30464 , n30700 );
and ( n30901 , n30899 , n30900 );
and ( n30902 , n30468 , n30592 );
and ( n30903 , n30900 , n30902 );
and ( n30904 , n30899 , n30902 );
or ( n30905 , n30901 , n30903 , n30904 );
and ( n30906 , n30896 , n30905 );
and ( n30907 , n30887 , n30906 );
and ( n30908 , n30803 , n30424 );
and ( n30909 , n30799 , n30439 );
or ( n30910 , n30908 , n30909 );
and ( n30911 , n30419 , n30788 );
and ( n30912 , n30442 , n30791 );
or ( n30913 , n30911 , n30912 );
and ( n30914 , n30910 , n30913 );
and ( n30915 , n30906 , n30914 );
and ( n30916 , n30887 , n30914 );
or ( n30917 , n30907 , n30915 , n30916 );
and ( n30918 , n30885 , n30917 );
and ( n30919 , n30878 , n30917 );
or ( n30920 , n30886 , n30918 , n30919 );
and ( n30921 , n30874 , n30920 );
and ( n30922 , n30861 , n30920 );
or ( n30923 , n30875 , n30921 , n30922 );
and ( n30924 , n30843 , n30923 );
and ( n30925 , n30841 , n30923 );
or ( n30926 , n30844 , n30924 , n30925 );
and ( n30927 , n30821 , n30926 );
and ( n30928 , n30819 , n30926 );
or ( n30929 , n30822 , n30927 , n30928 );
and ( n30930 , n30769 , n30929 );
and ( n30931 , n30767 , n30929 );
or ( n30932 , n30770 , n30930 , n30931 );
or ( n30933 , n30765 , n30932 );
and ( n30934 , n30763 , n30933 );
xor ( n30935 , n30763 , n30933 );
xnor ( n30936 , n30765 , n30932 );
xor ( n30937 , n30767 , n30769 );
xor ( n30938 , n30937 , n30929 );
xor ( n30939 , n30778 , n30780 );
xor ( n30940 , n30939 , n30816 );
xor ( n30941 , n30784 , n30785 );
xor ( n30942 , n30941 , n30813 );
xor ( n30943 , n30827 , n30835 );
xor ( n30944 , n30943 , n30838 );
and ( n30945 , n30942 , n30944 );
xor ( n30946 , n30828 , n30830 );
xor ( n30947 , n30946 , n30832 );
xor ( n30948 , n30804 , n30805 );
xor ( n30949 , n30948 , n30807 );
xor ( n30950 , n30789 , n30792 );
xor ( n30951 , n30950 , n30794 );
and ( n30952 , n30949 , n30951 );
xor ( n30953 , n30866 , n30868 );
and ( n30954 , n30952 , n30953 );
xor ( n30955 , n30876 , n30877 );
and ( n30956 , n30953 , n30955 );
and ( n30957 , n30952 , n30955 );
or ( n30958 , n30954 , n30956 , n30957 );
and ( n30959 , n30947 , n30958 );
and ( n30960 , n30419 , n30898 );
and ( n30961 , n30442 , n30788 );
and ( n30962 , n30960 , n30961 );
and ( n30963 , n30468 , n30700 );
and ( n30964 , n30961 , n30963 );
and ( n30965 , n30960 , n30963 );
or ( n30966 , n30962 , n30964 , n30965 );
xor ( n30967 , n30899 , n30900 );
xor ( n30968 , n30967 , n30902 );
or ( n30969 , n30966 , n30968 );
and ( n30970 , n30889 , n30424 );
and ( n30971 , n30803 , n30439 );
and ( n30972 , n30970 , n30971 );
and ( n30973 , n30709 , n30473 );
and ( n30974 , n30971 , n30973 );
and ( n30975 , n30970 , n30973 );
or ( n30976 , n30972 , n30974 , n30975 );
xor ( n30977 , n30890 , n30891 );
xor ( n30978 , n30977 , n30893 );
or ( n30979 , n30976 , n30978 );
and ( n30980 , n30969 , n30979 );
buf ( n30981 , n30503 );
buf ( n30982 , n15802 );
buf ( n30983 , n30982 );
and ( n30984 , n30981 , n30983 );
xor ( n30985 , n30896 , n30905 );
and ( n30986 , n30983 , n30985 );
and ( n30987 , n30981 , n30985 );
or ( n30988 , n30984 , n30986 , n30987 );
and ( n30989 , n30980 , n30988 );
xor ( n30990 , n30910 , n30913 );
xor ( n30991 , n30949 , n30951 );
and ( n30992 , n30990 , n30991 );
xor ( n30993 , n30863 , n30864 );
and ( n30994 , n30991 , n30993 );
and ( n30995 , n30990 , n30993 );
or ( n30996 , n30992 , n30994 , n30995 );
and ( n30997 , n30988 , n30996 );
and ( n30998 , n30980 , n30996 );
or ( n30999 , n30989 , n30997 , n30998 );
and ( n31000 , n30958 , n30999 );
and ( n31001 , n30947 , n30999 );
or ( n31002 , n30959 , n31000 , n31001 );
and ( n31003 , n30944 , n31002 );
and ( n31004 , n30942 , n31002 );
or ( n31005 , n30945 , n31003 , n31004 );
and ( n31006 , n30940 , n31005 );
xor ( n31007 , n30841 , n30843 );
xor ( n31008 , n31007 , n30923 );
and ( n31009 , n31005 , n31008 );
and ( n31010 , n30940 , n31008 );
or ( n31011 , n31006 , n31009 , n31010 );
xor ( n31012 , n30819 , n30821 );
xor ( n31013 , n31012 , n30926 );
and ( n31014 , n31011 , n31013 );
xor ( n31015 , n30851 , n30856 );
xor ( n31016 , n31015 , n30858 );
xor ( n31017 , n30862 , n30869 );
xor ( n31018 , n31017 , n30871 );
and ( n31019 , n31016 , n31018 );
xor ( n31020 , n30878 , n30885 );
xor ( n31021 , n31020 , n30917 );
and ( n31022 , n31018 , n31021 );
and ( n31023 , n31016 , n31021 );
or ( n31024 , n31019 , n31022 , n31023 );
xor ( n31025 , n30861 , n30874 );
xor ( n31026 , n31025 , n30920 );
and ( n31027 , n31024 , n31026 );
xor ( n31028 , n30879 , n30880 );
xor ( n31029 , n31028 , n30882 );
xor ( n31030 , n30887 , n30906 );
xor ( n31031 , n31030 , n30914 );
and ( n31032 , n31029 , n31031 );
and ( n31033 , n30799 , n30461 );
and ( n31034 , n30603 , n30508 );
or ( n31035 , n31033 , n31034 );
and ( n31036 , n30464 , n30791 );
and ( n31037 , n30503 , n30592 );
or ( n31038 , n31036 , n31037 );
and ( n31039 , n31035 , n31038 );
xnor ( n31040 , n30908 , n30909 );
xnor ( n31041 , n30911 , n30912 );
and ( n31042 , n31040 , n31041 );
and ( n31043 , n31039 , n31042 );
xor ( n31044 , n30969 , n30979 );
and ( n31045 , n31042 , n31044 );
and ( n31046 , n31039 , n31044 );
or ( n31047 , n31043 , n31045 , n31046 );
and ( n31048 , n31031 , n31047 );
and ( n31049 , n31029 , n31047 );
or ( n31050 , n31032 , n31048 , n31049 );
and ( n31051 , n30442 , n30898 );
and ( n31052 , n30464 , n30788 );
and ( n31053 , n31051 , n31052 );
and ( n31054 , n30468 , n30791 );
and ( n31055 , n31052 , n31054 );
and ( n31056 , n31051 , n31054 );
or ( n31057 , n31053 , n31055 , n31056 );
xor ( n31058 , n30960 , n30961 );
xor ( n31059 , n31058 , n30963 );
or ( n31060 , n31057 , n31059 );
and ( n31061 , n30889 , n30439 );
and ( n31062 , n30803 , n30461 );
and ( n31063 , n31061 , n31062 );
and ( n31064 , n30799 , n30473 );
and ( n31065 , n31062 , n31064 );
and ( n31066 , n31061 , n31064 );
or ( n31067 , n31063 , n31065 , n31066 );
xor ( n31068 , n30970 , n30971 );
xor ( n31069 , n31068 , n30973 );
or ( n31070 , n31067 , n31069 );
and ( n31071 , n31060 , n31070 );
buf ( n31072 , n1231 );
buf ( n31073 , n31072 );
and ( n31074 , n30413 , n31073 );
buf ( n31075 , n1230 );
buf ( n31076 , n31075 );
and ( n31077 , n30419 , n31076 );
and ( n31078 , n31074 , n31077 );
and ( n31079 , n30503 , n30700 );
and ( n31080 , n31077 , n31079 );
and ( n31081 , n31074 , n31079 );
or ( n31082 , n31078 , n31080 , n31081 );
buf ( n31083 , n1230 );
buf ( n31084 , n31083 );
and ( n31085 , n31084 , n30421 );
or ( n31086 , n31082 , n31085 );
buf ( n31087 , n1231 );
buf ( n31088 , n31087 );
and ( n31089 , n31088 , n30421 );
and ( n31090 , n31084 , n30424 );
and ( n31091 , n31089 , n31090 );
and ( n31092 , n30709 , n30508 );
and ( n31093 , n31090 , n31092 );
and ( n31094 , n31089 , n31092 );
or ( n31095 , n31091 , n31093 , n31094 );
and ( n31096 , n30413 , n31076 );
or ( n31097 , n31095 , n31096 );
and ( n31098 , n31086 , n31097 );
and ( n31099 , n31071 , n31098 );
xnor ( n31100 , n30966 , n30968 );
xnor ( n31101 , n30976 , n30978 );
and ( n31102 , n31100 , n31101 );
and ( n31103 , n31098 , n31102 );
and ( n31104 , n31071 , n31102 );
or ( n31105 , n31099 , n31103 , n31104 );
and ( n31106 , n30558 , n30508 );
and ( n31107 , n30503 , n30563 );
and ( n31108 , n31106 , n31107 );
xor ( n31109 , n31035 , n31038 );
and ( n31110 , n31107 , n31109 );
and ( n31111 , n31106 , n31109 );
or ( n31112 , n31108 , n31110 , n31111 );
xor ( n31113 , n30981 , n30983 );
xor ( n31114 , n31113 , n30985 );
and ( n31115 , n31112 , n31114 );
xor ( n31116 , n30990 , n30991 );
xor ( n31117 , n31116 , n30993 );
and ( n31118 , n31114 , n31117 );
and ( n31119 , n31112 , n31117 );
or ( n31120 , n31115 , n31118 , n31119 );
and ( n31121 , n31105 , n31120 );
xor ( n31122 , n30952 , n30953 );
xor ( n31123 , n31122 , n30955 );
and ( n31124 , n31120 , n31123 );
and ( n31125 , n31105 , n31123 );
or ( n31126 , n31121 , n31124 , n31125 );
and ( n31127 , n31050 , n31126 );
xor ( n31128 , n30947 , n30958 );
xor ( n31129 , n31128 , n30999 );
and ( n31130 , n31126 , n31129 );
and ( n31131 , n31050 , n31129 );
or ( n31132 , n31127 , n31130 , n31131 );
and ( n31133 , n31026 , n31132 );
and ( n31134 , n31024 , n31132 );
or ( n31135 , n31027 , n31133 , n31134 );
xor ( n31136 , n30940 , n31005 );
xor ( n31137 , n31136 , n31008 );
and ( n31138 , n31135 , n31137 );
xor ( n31139 , n30942 , n30944 );
xor ( n31140 , n31139 , n31002 );
xor ( n31141 , n31016 , n31018 );
xor ( n31142 , n31141 , n31021 );
xor ( n31143 , n30980 , n30988 );
xor ( n31144 , n31143 , n30996 );
xnor ( n31145 , n31036 , n31037 );
xnor ( n31146 , n31067 , n31069 );
or ( n31147 , n31145 , n31146 );
xnor ( n31148 , n31033 , n31034 );
xnor ( n31149 , n31057 , n31059 );
or ( n31150 , n31148 , n31149 );
and ( n31151 , n31147 , n31150 );
xor ( n31152 , n31040 , n31041 );
buf ( n31153 , n30558 );
buf ( n31154 , n15808 );
buf ( n31155 , n31154 );
and ( n31156 , n31153 , n31155 );
and ( n31157 , n30603 , n30563 );
and ( n31158 , n30558 , n30592 );
and ( n31159 , n31157 , n31158 );
buf ( n31160 , n15811 );
buf ( n31161 , n31160 );
and ( n31162 , n31158 , n31161 );
and ( n31163 , n31157 , n31161 );
or ( n31164 , n31159 , n31162 , n31163 );
and ( n31165 , n31155 , n31164 );
and ( n31166 , n31153 , n31164 );
or ( n31167 , n31156 , n31165 , n31166 );
and ( n31168 , n31152 , n31167 );
xor ( n31169 , n31060 , n31070 );
and ( n31170 , n31167 , n31169 );
and ( n31171 , n31152 , n31169 );
or ( n31172 , n31168 , n31170 , n31171 );
and ( n31173 , n31151 , n31172 );
xor ( n31174 , n31086 , n31097 );
xor ( n31175 , n31100 , n31101 );
and ( n31176 , n31174 , n31175 );
xnor ( n31177 , n31082 , n31085 );
xnor ( n31178 , n31095 , n31096 );
and ( n31179 , n31177 , n31178 );
and ( n31180 , n31175 , n31179 );
and ( n31181 , n31174 , n31179 );
or ( n31182 , n31176 , n31180 , n31181 );
and ( n31183 , n31172 , n31182 );
and ( n31184 , n31151 , n31182 );
or ( n31185 , n31173 , n31183 , n31184 );
and ( n31186 , n31144 , n31185 );
xor ( n31187 , n31039 , n31042 );
xor ( n31188 , n31187 , n31044 );
xor ( n31189 , n31071 , n31098 );
xor ( n31190 , n31189 , n31102 );
and ( n31191 , n31188 , n31190 );
xor ( n31192 , n31112 , n31114 );
xor ( n31193 , n31192 , n31117 );
and ( n31194 , n31190 , n31193 );
and ( n31195 , n31188 , n31193 );
or ( n31196 , n31191 , n31194 , n31195 );
and ( n31197 , n31185 , n31196 );
and ( n31198 , n31144 , n31196 );
or ( n31199 , n31186 , n31197 , n31198 );
and ( n31200 , n31142 , n31199 );
xor ( n31201 , n31050 , n31126 );
xor ( n31202 , n31201 , n31129 );
and ( n31203 , n31199 , n31202 );
and ( n31204 , n31142 , n31202 );
or ( n31205 , n31200 , n31203 , n31204 );
and ( n31206 , n31140 , n31205 );
xor ( n31207 , n31024 , n31026 );
xor ( n31208 , n31207 , n31132 );
and ( n31209 , n31205 , n31208 );
and ( n31210 , n31140 , n31208 );
or ( n31211 , n31206 , n31209 , n31210 );
and ( n31212 , n31137 , n31211 );
and ( n31213 , n31135 , n31211 );
or ( n31214 , n31138 , n31212 , n31213 );
and ( n31215 , n31013 , n31214 );
and ( n31216 , n31011 , n31214 );
or ( n31217 , n31014 , n31215 , n31216 );
and ( n31218 , n30938 , n31217 );
xor ( n31219 , n30938 , n31217 );
xor ( n31220 , n31011 , n31013 );
xor ( n31221 , n31220 , n31214 );
xor ( n31222 , n31135 , n31137 );
xor ( n31223 , n31222 , n31211 );
xor ( n31224 , n31140 , n31205 );
xor ( n31225 , n31224 , n31208 );
xor ( n31226 , n31029 , n31031 );
xor ( n31227 , n31226 , n31047 );
xor ( n31228 , n31105 , n31120 );
xor ( n31229 , n31228 , n31123 );
and ( n31230 , n31227 , n31229 );
xnor ( n31231 , n31145 , n31146 );
xnor ( n31232 , n31148 , n31149 );
and ( n31233 , n31231 , n31232 );
buf ( n31234 , n15805 );
buf ( n31235 , n31234 );
or ( n31236 , n31233 , n31235 );
buf ( n31237 , n1232 );
buf ( n31238 , n31237 );
and ( n31239 , n31238 , n30421 );
and ( n31240 , n30889 , n30461 );
and ( n31241 , n31239 , n31240 );
and ( n31242 , n30799 , n30508 );
and ( n31243 , n31240 , n31242 );
and ( n31244 , n31239 , n31242 );
or ( n31245 , n31241 , n31243 , n31244 );
buf ( n31246 , n1232 );
buf ( n31247 , n31246 );
and ( n31248 , n30413 , n31247 );
and ( n31249 , n30464 , n30898 );
and ( n31250 , n31248 , n31249 );
and ( n31251 , n30503 , n30791 );
and ( n31252 , n31249 , n31251 );
and ( n31253 , n31248 , n31251 );
or ( n31254 , n31250 , n31252 , n31253 );
and ( n31255 , n31245 , n31254 );
and ( n31256 , n30803 , n30473 );
and ( n31257 , n30709 , n30563 );
or ( n31258 , n31256 , n31257 );
and ( n31259 , n30468 , n30788 );
and ( n31260 , n30558 , n30700 );
or ( n31261 , n31259 , n31260 );
and ( n31262 , n31258 , n31261 );
and ( n31263 , n31255 , n31262 );
xor ( n31264 , n31153 , n31155 );
xor ( n31265 , n31264 , n31164 );
and ( n31266 , n31262 , n31265 );
and ( n31267 , n31255 , n31265 );
or ( n31268 , n31263 , n31266 , n31267 );
xor ( n31269 , n31106 , n31107 );
xor ( n31270 , n31269 , n31109 );
and ( n31271 , n31268 , n31270 );
xor ( n31272 , n31147 , n31150 );
and ( n31273 , n31270 , n31272 );
and ( n31274 , n31268 , n31272 );
or ( n31275 , n31271 , n31273 , n31274 );
and ( n31276 , n31236 , n31275 );
buf ( n31277 , n1233 );
buf ( n31278 , n31277 );
and ( n31279 , n31278 , n30421 );
and ( n31280 , n30889 , n30473 );
and ( n31281 , n31279 , n31280 );
and ( n31282 , n30803 , n30508 );
and ( n31283 , n31280 , n31282 );
and ( n31284 , n31279 , n31282 );
or ( n31285 , n31281 , n31283 , n31284 );
and ( n31286 , n30419 , n31073 );
and ( n31287 , n31285 , n31286 );
and ( n31288 , n30442 , n31076 );
and ( n31289 , n31286 , n31288 );
and ( n31290 , n31285 , n31288 );
or ( n31291 , n31287 , n31289 , n31290 );
xor ( n31292 , n31089 , n31090 );
xor ( n31293 , n31292 , n31092 );
and ( n31294 , n31291 , n31293 );
xor ( n31295 , n31061 , n31062 );
xor ( n31296 , n31295 , n31064 );
and ( n31297 , n31293 , n31296 );
and ( n31298 , n31291 , n31296 );
or ( n31299 , n31294 , n31297 , n31298 );
buf ( n31300 , n1233 );
buf ( n31301 , n31300 );
and ( n31302 , n30413 , n31301 );
and ( n31303 , n30468 , n30898 );
and ( n31304 , n31302 , n31303 );
and ( n31305 , n30503 , n30788 );
and ( n31306 , n31303 , n31305 );
and ( n31307 , n31302 , n31305 );
or ( n31308 , n31304 , n31306 , n31307 );
and ( n31309 , n31088 , n30424 );
and ( n31310 , n31308 , n31309 );
and ( n31311 , n31084 , n30439 );
and ( n31312 , n31309 , n31311 );
and ( n31313 , n31308 , n31311 );
or ( n31314 , n31310 , n31312 , n31313 );
xor ( n31315 , n31074 , n31077 );
xor ( n31316 , n31315 , n31079 );
and ( n31317 , n31314 , n31316 );
xor ( n31318 , n31051 , n31052 );
xor ( n31319 , n31318 , n31054 );
and ( n31320 , n31316 , n31319 );
and ( n31321 , n31314 , n31319 );
or ( n31322 , n31317 , n31320 , n31321 );
and ( n31323 , n31299 , n31322 );
xor ( n31324 , n31177 , n31178 );
xor ( n31325 , n31157 , n31158 );
xor ( n31326 , n31325 , n31161 );
xor ( n31327 , n31245 , n31254 );
and ( n31328 , n31326 , n31327 );
xor ( n31329 , n31258 , n31261 );
and ( n31330 , n31327 , n31329 );
and ( n31331 , n31326 , n31329 );
or ( n31332 , n31328 , n31330 , n31331 );
and ( n31333 , n31324 , n31332 );
and ( n31334 , n31238 , n30424 );
and ( n31335 , n31088 , n30439 );
and ( n31336 , n31334 , n31335 );
and ( n31337 , n30799 , n30563 );
and ( n31338 , n31335 , n31337 );
and ( n31339 , n31334 , n31337 );
or ( n31340 , n31336 , n31338 , n31339 );
and ( n31341 , n30419 , n31247 );
and ( n31342 , n30442 , n31073 );
and ( n31343 , n31341 , n31342 );
and ( n31344 , n30558 , n30791 );
and ( n31345 , n31342 , n31344 );
and ( n31346 , n31341 , n31344 );
or ( n31347 , n31343 , n31345 , n31346 );
and ( n31348 , n31340 , n31347 );
xnor ( n31349 , n31256 , n31257 );
xnor ( n31350 , n31259 , n31260 );
and ( n31351 , n31349 , n31350 );
and ( n31352 , n31348 , n31351 );
buf ( n31353 , n30603 );
buf ( n31354 , n15814 );
buf ( n31355 , n31354 );
and ( n31356 , n31353 , n31355 );
and ( n31357 , n30464 , n31076 );
and ( n31358 , n31084 , n30461 );
and ( n31359 , n31357 , n31358 );
and ( n31360 , n31355 , n31359 );
and ( n31361 , n31353 , n31359 );
or ( n31362 , n31356 , n31360 , n31361 );
and ( n31363 , n31351 , n31362 );
and ( n31364 , n31348 , n31362 );
or ( n31365 , n31352 , n31363 , n31364 );
and ( n31366 , n31332 , n31365 );
and ( n31367 , n31324 , n31365 );
or ( n31368 , n31333 , n31366 , n31367 );
and ( n31369 , n31323 , n31368 );
xor ( n31370 , n31152 , n31167 );
xor ( n31371 , n31370 , n31169 );
and ( n31372 , n31368 , n31371 );
and ( n31373 , n31323 , n31371 );
or ( n31374 , n31369 , n31372 , n31373 );
and ( n31375 , n31275 , n31374 );
and ( n31376 , n31236 , n31374 );
or ( n31377 , n31276 , n31375 , n31376 );
and ( n31378 , n31229 , n31377 );
and ( n31379 , n31227 , n31377 );
or ( n31380 , n31230 , n31378 , n31379 );
xor ( n31381 , n31142 , n31199 );
xor ( n31382 , n31381 , n31202 );
and ( n31383 , n31380 , n31382 );
xor ( n31384 , n31144 , n31185 );
xor ( n31385 , n31384 , n31196 );
xor ( n31386 , n31151 , n31172 );
xor ( n31387 , n31386 , n31182 );
xor ( n31388 , n31188 , n31190 );
xor ( n31389 , n31388 , n31193 );
and ( n31390 , n31387 , n31389 );
xor ( n31391 , n31174 , n31175 );
xor ( n31392 , n31391 , n31179 );
xnor ( n31393 , n31233 , n31235 );
and ( n31394 , n31392 , n31393 );
xor ( n31395 , n31255 , n31262 );
xor ( n31396 , n31395 , n31265 );
xor ( n31397 , n31299 , n31322 );
and ( n31398 , n31396 , n31397 );
xor ( n31399 , n31231 , n31232 );
and ( n31400 , n31397 , n31399 );
and ( n31401 , n31396 , n31399 );
or ( n31402 , n31398 , n31400 , n31401 );
and ( n31403 , n31393 , n31402 );
and ( n31404 , n31392 , n31402 );
or ( n31405 , n31394 , n31403 , n31404 );
and ( n31406 , n31389 , n31405 );
and ( n31407 , n31387 , n31405 );
or ( n31408 , n31390 , n31406 , n31407 );
and ( n31409 , n31385 , n31408 );
xor ( n31410 , n31227 , n31229 );
xor ( n31411 , n31410 , n31377 );
and ( n31412 , n31408 , n31411 );
and ( n31413 , n31385 , n31411 );
or ( n31414 , n31409 , n31412 , n31413 );
and ( n31415 , n31382 , n31414 );
and ( n31416 , n31380 , n31414 );
or ( n31417 , n31383 , n31415 , n31416 );
or ( n31418 , n31225 , n31417 );
and ( n31419 , n31223 , n31418 );
xor ( n31420 , n31223 , n31418 );
xnor ( n31421 , n31225 , n31417 );
xor ( n31422 , n31380 , n31382 );
xor ( n31423 , n31422 , n31414 );
xor ( n31424 , n31248 , n31249 );
xor ( n31425 , n31424 , n31251 );
xor ( n31426 , n31285 , n31286 );
xor ( n31427 , n31426 , n31288 );
or ( n31428 , n31425 , n31427 );
xor ( n31429 , n31239 , n31240 );
xor ( n31430 , n31429 , n31242 );
xor ( n31431 , n31308 , n31309 );
xor ( n31432 , n31431 , n31311 );
or ( n31433 , n31430 , n31432 );
and ( n31434 , n31428 , n31433 );
xor ( n31435 , n31291 , n31293 );
xor ( n31436 , n31435 , n31296 );
xor ( n31437 , n31314 , n31316 );
xor ( n31438 , n31437 , n31319 );
and ( n31439 , n31436 , n31438 );
and ( n31440 , n31434 , n31439 );
buf ( n31441 , n1234 );
buf ( n31442 , n31441 );
and ( n31443 , n30413 , n31442 );
and ( n31444 , n30419 , n31301 );
and ( n31445 , n31443 , n31444 );
and ( n31446 , n30468 , n31076 );
and ( n31447 , n31444 , n31446 );
and ( n31448 , n31443 , n31446 );
or ( n31449 , n31445 , n31447 , n31448 );
and ( n31450 , n30442 , n31247 );
and ( n31451 , n30464 , n31073 );
and ( n31452 , n31450 , n31451 );
and ( n31453 , n30558 , n30788 );
and ( n31454 , n31451 , n31453 );
and ( n31455 , n31450 , n31453 );
or ( n31456 , n31452 , n31454 , n31455 );
and ( n31457 , n31449 , n31456 );
xor ( n31458 , n31334 , n31335 );
xor ( n31459 , n31458 , n31337 );
and ( n31460 , n31456 , n31459 );
and ( n31461 , n31449 , n31459 );
or ( n31462 , n31457 , n31460 , n31461 );
buf ( n31463 , n1234 );
buf ( n31464 , n31463 );
and ( n31465 , n31464 , n30421 );
and ( n31466 , n31278 , n30424 );
and ( n31467 , n31465 , n31466 );
and ( n31468 , n31084 , n30473 );
and ( n31469 , n31466 , n31468 );
and ( n31470 , n31465 , n31468 );
or ( n31471 , n31467 , n31469 , n31470 );
and ( n31472 , n31238 , n30439 );
and ( n31473 , n31088 , n30461 );
and ( n31474 , n31472 , n31473 );
and ( n31475 , n30803 , n30563 );
and ( n31476 , n31473 , n31475 );
and ( n31477 , n31472 , n31475 );
or ( n31478 , n31474 , n31476 , n31477 );
and ( n31479 , n31471 , n31478 );
xor ( n31480 , n31341 , n31342 );
xor ( n31481 , n31480 , n31344 );
and ( n31482 , n31478 , n31481 );
and ( n31483 , n31471 , n31481 );
or ( n31484 , n31479 , n31482 , n31483 );
and ( n31485 , n31462 , n31484 );
xor ( n31486 , n31340 , n31347 );
xor ( n31487 , n31349 , n31350 );
and ( n31488 , n31486 , n31487 );
and ( n31489 , n30889 , n30508 );
and ( n31490 , n30799 , n30592 );
or ( n31491 , n31489 , n31490 );
and ( n31492 , n30503 , n30898 );
and ( n31493 , n30603 , n30791 );
or ( n31494 , n31492 , n31493 );
and ( n31495 , n31491 , n31494 );
and ( n31496 , n31487 , n31495 );
and ( n31497 , n31486 , n31495 );
or ( n31498 , n31488 , n31496 , n31497 );
and ( n31499 , n31485 , n31498 );
xor ( n31500 , n31279 , n31280 );
xor ( n31501 , n31500 , n31282 );
xor ( n31502 , n31302 , n31303 );
xor ( n31503 , n31502 , n31305 );
and ( n31504 , n31501 , n31503 );
and ( n31505 , n30709 , n30592 );
and ( n31506 , n30603 , n30700 );
and ( n31507 , n31505 , n31506 );
xor ( n31508 , n31357 , n31358 );
and ( n31509 , n31506 , n31508 );
and ( n31510 , n31505 , n31508 );
or ( n31511 , n31507 , n31509 , n31510 );
and ( n31512 , n31504 , n31511 );
xor ( n31513 , n31353 , n31355 );
xor ( n31514 , n31513 , n31359 );
and ( n31515 , n31511 , n31514 );
and ( n31516 , n31504 , n31514 );
or ( n31517 , n31512 , n31515 , n31516 );
and ( n31518 , n31498 , n31517 );
and ( n31519 , n31485 , n31517 );
or ( n31520 , n31499 , n31518 , n31519 );
and ( n31521 , n31439 , n31520 );
and ( n31522 , n31434 , n31520 );
or ( n31523 , n31440 , n31521 , n31522 );
xor ( n31524 , n31268 , n31270 );
xor ( n31525 , n31524 , n31272 );
and ( n31526 , n31523 , n31525 );
xor ( n31527 , n31323 , n31368 );
xor ( n31528 , n31527 , n31371 );
and ( n31529 , n31525 , n31528 );
and ( n31530 , n31523 , n31528 );
or ( n31531 , n31526 , n31529 , n31530 );
xor ( n31532 , n31236 , n31275 );
xor ( n31533 , n31532 , n31374 );
and ( n31534 , n31531 , n31533 );
xor ( n31535 , n31324 , n31332 );
xor ( n31536 , n31535 , n31365 );
xor ( n31537 , n31326 , n31327 );
xor ( n31538 , n31537 , n31329 );
xor ( n31539 , n31348 , n31351 );
xor ( n31540 , n31539 , n31362 );
and ( n31541 , n31538 , n31540 );
xor ( n31542 , n31428 , n31433 );
and ( n31543 , n31540 , n31542 );
and ( n31544 , n31538 , n31542 );
or ( n31545 , n31541 , n31543 , n31544 );
and ( n31546 , n31536 , n31545 );
xor ( n31547 , n31436 , n31438 );
xnor ( n31548 , n31425 , n31427 );
xnor ( n31549 , n31430 , n31432 );
and ( n31550 , n31548 , n31549 );
and ( n31551 , n31547 , n31550 );
xor ( n31552 , n31462 , n31484 );
xnor ( n31553 , n31489 , n31490 );
xnor ( n31554 , n31492 , n31493 );
and ( n31555 , n31553 , n31554 );
not ( n31556 , n31555 );
buf ( n31557 , n15817 );
buf ( n31558 , n31557 );
and ( n31559 , n31556 , n31558 );
and ( n31560 , n31552 , n31559 );
buf ( n31561 , n31555 );
and ( n31562 , n31559 , n31561 );
and ( n31563 , n31552 , n31561 );
or ( n31564 , n31560 , n31562 , n31563 );
and ( n31565 , n31550 , n31564 );
and ( n31566 , n31547 , n31564 );
or ( n31567 , n31551 , n31565 , n31566 );
and ( n31568 , n31545 , n31567 );
and ( n31569 , n31536 , n31567 );
or ( n31570 , n31546 , n31568 , n31569 );
xor ( n31571 , n31443 , n31444 );
xor ( n31572 , n31571 , n31446 );
xor ( n31573 , n31450 , n31451 );
xor ( n31574 , n31573 , n31453 );
or ( n31575 , n31572 , n31574 );
xor ( n31576 , n31465 , n31466 );
xor ( n31577 , n31576 , n31468 );
xor ( n31578 , n31472 , n31473 );
xor ( n31579 , n31578 , n31475 );
or ( n31580 , n31577 , n31579 );
and ( n31581 , n31575 , n31580 );
and ( n31582 , n30442 , n31301 );
and ( n31583 , n30464 , n31247 );
and ( n31584 , n31582 , n31583 );
and ( n31585 , n30603 , n30788 );
and ( n31586 , n31583 , n31585 );
and ( n31587 , n31582 , n31585 );
or ( n31588 , n31584 , n31586 , n31587 );
buf ( n31589 , n1235 );
buf ( n31590 , n31589 );
and ( n31591 , n30413 , n31590 );
and ( n31592 , n30419 , n31442 );
and ( n31593 , n31591 , n31592 );
and ( n31594 , n30558 , n30898 );
and ( n31595 , n31592 , n31594 );
and ( n31596 , n31591 , n31594 );
or ( n31597 , n31593 , n31595 , n31596 );
and ( n31598 , n31588 , n31597 );
and ( n31599 , n31278 , n30439 );
and ( n31600 , n31238 , n30461 );
and ( n31601 , n31599 , n31600 );
and ( n31602 , n30803 , n30592 );
and ( n31603 , n31600 , n31602 );
and ( n31604 , n31599 , n31602 );
or ( n31605 , n31601 , n31603 , n31604 );
buf ( n31606 , n1235 );
buf ( n31607 , n31606 );
and ( n31608 , n31607 , n30421 );
and ( n31609 , n31464 , n30424 );
and ( n31610 , n31608 , n31609 );
and ( n31611 , n30889 , n30563 );
and ( n31612 , n31609 , n31611 );
and ( n31613 , n31608 , n31611 );
or ( n31614 , n31610 , n31612 , n31613 );
and ( n31615 , n31605 , n31614 );
and ( n31616 , n31598 , n31615 );
and ( n31617 , n31581 , n31616 );
xor ( n31618 , n31449 , n31456 );
xor ( n31619 , n31618 , n31459 );
xor ( n31620 , n31471 , n31478 );
xor ( n31621 , n31620 , n31481 );
and ( n31622 , n31619 , n31621 );
and ( n31623 , n31616 , n31622 );
and ( n31624 , n31581 , n31622 );
or ( n31625 , n31617 , n31623 , n31624 );
xor ( n31626 , n31491 , n31494 );
xor ( n31627 , n31501 , n31503 );
and ( n31628 , n31626 , n31627 );
and ( n31629 , n31088 , n30473 );
and ( n31630 , n31084 , n30508 );
or ( n31631 , n31629 , n31630 );
and ( n31632 , n30468 , n31073 );
and ( n31633 , n30503 , n31076 );
or ( n31634 , n31632 , n31633 );
and ( n31635 , n31631 , n31634 );
and ( n31636 , n31627 , n31635 );
and ( n31637 , n31626 , n31635 );
or ( n31638 , n31628 , n31636 , n31637 );
xor ( n31639 , n31486 , n31487 );
xor ( n31640 , n31639 , n31495 );
and ( n31641 , n31638 , n31640 );
xor ( n31642 , n31504 , n31511 );
xor ( n31643 , n31642 , n31514 );
and ( n31644 , n31640 , n31643 );
and ( n31645 , n31638 , n31643 );
or ( n31646 , n31641 , n31644 , n31645 );
and ( n31647 , n31625 , n31646 );
xor ( n31648 , n31485 , n31498 );
xor ( n31649 , n31648 , n31517 );
and ( n31650 , n31646 , n31649 );
and ( n31651 , n31625 , n31649 );
or ( n31652 , n31647 , n31650 , n31651 );
xor ( n31653 , n31396 , n31397 );
xor ( n31654 , n31653 , n31399 );
and ( n31655 , n31652 , n31654 );
xor ( n31656 , n31434 , n31439 );
xor ( n31657 , n31656 , n31520 );
and ( n31658 , n31654 , n31657 );
and ( n31659 , n31652 , n31657 );
or ( n31660 , n31655 , n31658 , n31659 );
and ( n31661 , n31570 , n31660 );
xor ( n31662 , n31392 , n31393 );
xor ( n31663 , n31662 , n31402 );
and ( n31664 , n31660 , n31663 );
and ( n31665 , n31570 , n31663 );
or ( n31666 , n31661 , n31664 , n31665 );
and ( n31667 , n31533 , n31666 );
and ( n31668 , n31531 , n31666 );
or ( n31669 , n31534 , n31667 , n31668 );
xor ( n31670 , n31385 , n31408 );
xor ( n31671 , n31670 , n31411 );
and ( n31672 , n31669 , n31671 );
xor ( n31673 , n31387 , n31389 );
xor ( n31674 , n31673 , n31405 );
xor ( n31675 , n31523 , n31525 );
xor ( n31676 , n31675 , n31528 );
xor ( n31677 , n31548 , n31549 );
buf ( n31678 , n30709 );
buf ( n31679 , n15820 );
buf ( n31680 , n31679 );
and ( n31681 , n31678 , n31680 );
and ( n31682 , n30799 , n30700 );
and ( n31683 , n30709 , n30791 );
and ( n31684 , n31682 , n31683 );
buf ( n31685 , n15823 );
buf ( n31686 , n31685 );
and ( n31687 , n31683 , n31686 );
and ( n31688 , n31682 , n31686 );
or ( n31689 , n31684 , n31687 , n31688 );
and ( n31690 , n31680 , n31689 );
and ( n31691 , n31678 , n31689 );
or ( n31692 , n31681 , n31690 , n31691 );
xor ( n31693 , n31505 , n31506 );
xor ( n31694 , n31693 , n31508 );
and ( n31695 , n31692 , n31694 );
xor ( n31696 , n31556 , n31558 );
and ( n31697 , n31694 , n31696 );
and ( n31698 , n31692 , n31696 );
or ( n31699 , n31695 , n31697 , n31698 );
and ( n31700 , n31677 , n31699 );
xor ( n31701 , n31575 , n31580 );
xor ( n31702 , n31598 , n31615 );
and ( n31703 , n31701 , n31702 );
xor ( n31704 , n31619 , n31621 );
and ( n31705 , n31702 , n31704 );
and ( n31706 , n31701 , n31704 );
or ( n31707 , n31703 , n31705 , n31706 );
and ( n31708 , n31699 , n31707 );
and ( n31709 , n31677 , n31707 );
or ( n31710 , n31700 , n31708 , n31709 );
xor ( n31711 , n31582 , n31583 );
xor ( n31712 , n31711 , n31585 );
xor ( n31713 , n31591 , n31592 );
xor ( n31714 , n31713 , n31594 );
or ( n31715 , n31712 , n31714 );
xor ( n31716 , n31599 , n31600 );
xor ( n31717 , n31716 , n31602 );
xor ( n31718 , n31608 , n31609 );
xor ( n31719 , n31718 , n31611 );
or ( n31720 , n31717 , n31719 );
and ( n31721 , n31715 , n31720 );
xnor ( n31722 , n31572 , n31574 );
xnor ( n31723 , n31577 , n31579 );
and ( n31724 , n31722 , n31723 );
and ( n31725 , n31721 , n31724 );
xor ( n31726 , n31588 , n31597 );
xor ( n31727 , n31605 , n31614 );
and ( n31728 , n31726 , n31727 );
and ( n31729 , n31724 , n31728 );
and ( n31730 , n31721 , n31728 );
or ( n31731 , n31725 , n31729 , n31730 );
xor ( n31732 , n31631 , n31634 );
xor ( n31733 , n31553 , n31554 );
and ( n31734 , n31732 , n31733 );
buf ( n31735 , n1236 );
buf ( n31736 , n31735 );
and ( n31737 , n31736 , n30421 );
and ( n31738 , n31238 , n30473 );
and ( n31739 , n31737 , n31738 );
and ( n31740 , n30889 , n30592 );
and ( n31741 , n31738 , n31740 );
and ( n31742 , n31737 , n31740 );
or ( n31743 , n31739 , n31741 , n31742 );
buf ( n31744 , n1236 );
buf ( n31745 , n31744 );
and ( n31746 , n30413 , n31745 );
and ( n31747 , n30468 , n31247 );
and ( n31748 , n31746 , n31747 );
and ( n31749 , n30603 , n30898 );
and ( n31750 , n31747 , n31749 );
and ( n31751 , n31746 , n31749 );
or ( n31752 , n31748 , n31750 , n31751 );
and ( n31753 , n31743 , n31752 );
and ( n31754 , n31733 , n31753 );
and ( n31755 , n31732 , n31753 );
or ( n31756 , n31734 , n31754 , n31755 );
and ( n31757 , n31607 , n30424 );
and ( n31758 , n31464 , n30439 );
and ( n31759 , n31757 , n31758 );
and ( n31760 , n31088 , n30508 );
and ( n31761 , n31758 , n31760 );
and ( n31762 , n31757 , n31760 );
or ( n31763 , n31759 , n31761 , n31762 );
and ( n31764 , n30419 , n31590 );
and ( n31765 , n30442 , n31442 );
and ( n31766 , n31764 , n31765 );
and ( n31767 , n30503 , n31073 );
and ( n31768 , n31765 , n31767 );
and ( n31769 , n31764 , n31767 );
or ( n31770 , n31766 , n31768 , n31769 );
and ( n31771 , n31763 , n31770 );
and ( n31772 , n31084 , n30563 );
and ( n31773 , n30803 , n30700 );
or ( n31774 , n31772 , n31773 );
and ( n31775 , n30558 , n31076 );
and ( n31776 , n30709 , n30788 );
or ( n31777 , n31775 , n31776 );
and ( n31778 , n31774 , n31777 );
and ( n31779 , n31771 , n31778 );
xnor ( n31780 , n31629 , n31630 );
xnor ( n31781 , n31632 , n31633 );
and ( n31782 , n31780 , n31781 );
and ( n31783 , n31778 , n31782 );
and ( n31784 , n31771 , n31782 );
or ( n31785 , n31779 , n31783 , n31784 );
and ( n31786 , n31756 , n31785 );
xor ( n31787 , n31626 , n31627 );
xor ( n31788 , n31787 , n31635 );
and ( n31789 , n31785 , n31788 );
and ( n31790 , n31756 , n31788 );
or ( n31791 , n31786 , n31789 , n31790 );
and ( n31792 , n31731 , n31791 );
xor ( n31793 , n31552 , n31559 );
xor ( n31794 , n31793 , n31561 );
and ( n31795 , n31791 , n31794 );
and ( n31796 , n31731 , n31794 );
or ( n31797 , n31792 , n31795 , n31796 );
and ( n31798 , n31710 , n31797 );
xor ( n31799 , n31538 , n31540 );
xor ( n31800 , n31799 , n31542 );
and ( n31801 , n31797 , n31800 );
and ( n31802 , n31710 , n31800 );
or ( n31803 , n31798 , n31801 , n31802 );
xor ( n31804 , n31536 , n31545 );
xor ( n31805 , n31804 , n31567 );
and ( n31806 , n31803 , n31805 );
xor ( n31807 , n31652 , n31654 );
xor ( n31808 , n31807 , n31657 );
and ( n31809 , n31805 , n31808 );
and ( n31810 , n31803 , n31808 );
or ( n31811 , n31806 , n31809 , n31810 );
and ( n31812 , n31676 , n31811 );
xor ( n31813 , n31570 , n31660 );
xor ( n31814 , n31813 , n31663 );
and ( n31815 , n31811 , n31814 );
and ( n31816 , n31676 , n31814 );
or ( n31817 , n31812 , n31815 , n31816 );
or ( n31818 , n31674 , n31817 );
and ( n31819 , n31671 , n31818 );
and ( n31820 , n31669 , n31818 );
or ( n31821 , n31672 , n31819 , n31820 );
and ( n31822 , n31423 , n31821 );
xor ( n31823 , n31423 , n31821 );
xor ( n31824 , n31669 , n31671 );
xor ( n31825 , n31824 , n31818 );
not ( n31826 , n31825 );
xor ( n31827 , n31531 , n31533 );
xor ( n31828 , n31827 , n31666 );
xnor ( n31829 , n31674 , n31817 );
and ( n31830 , n31828 , n31829 );
xor ( n31831 , n31828 , n31829 );
xor ( n31832 , n31676 , n31811 );
xor ( n31833 , n31832 , n31814 );
xor ( n31834 , n31547 , n31550 );
xor ( n31835 , n31834 , n31564 );
xor ( n31836 , n31625 , n31646 );
xor ( n31837 , n31836 , n31649 );
and ( n31838 , n31835 , n31837 );
xor ( n31839 , n31581 , n31616 );
xor ( n31840 , n31839 , n31622 );
xor ( n31841 , n31638 , n31640 );
xor ( n31842 , n31841 , n31643 );
and ( n31843 , n31840 , n31842 );
xor ( n31844 , n31678 , n31680 );
xor ( n31845 , n31844 , n31689 );
xor ( n31846 , n31715 , n31720 );
and ( n31847 , n31845 , n31846 );
xor ( n31848 , n31722 , n31723 );
and ( n31849 , n31846 , n31848 );
and ( n31850 , n31845 , n31848 );
or ( n31851 , n31847 , n31849 , n31850 );
xor ( n31852 , n31726 , n31727 );
and ( n31853 , n30419 , n31745 );
and ( n31854 , n30442 , n31590 );
and ( n31855 , n31853 , n31854 );
and ( n31856 , n30603 , n31076 );
and ( n31857 , n31854 , n31856 );
and ( n31858 , n31853 , n31856 );
or ( n31859 , n31855 , n31857 , n31858 );
buf ( n31860 , n1237 );
buf ( n31861 , n31860 );
and ( n31862 , n30413 , n31861 );
and ( n31863 , n30503 , n31247 );
and ( n31864 , n31862 , n31863 );
and ( n31865 , n30558 , n31073 );
and ( n31866 , n31863 , n31865 );
and ( n31867 , n31862 , n31865 );
or ( n31868 , n31864 , n31866 , n31867 );
and ( n31869 , n31859 , n31868 );
xor ( n31870 , n31737 , n31738 );
xor ( n31871 , n31870 , n31740 );
and ( n31872 , n31868 , n31871 );
and ( n31873 , n31859 , n31871 );
or ( n31874 , n31869 , n31872 , n31873 );
and ( n31875 , n31736 , n30424 );
and ( n31876 , n31607 , n30439 );
and ( n31877 , n31875 , n31876 );
and ( n31878 , n31084 , n30592 );
and ( n31879 , n31876 , n31878 );
and ( n31880 , n31875 , n31878 );
or ( n31881 , n31877 , n31879 , n31880 );
buf ( n31882 , n1237 );
buf ( n31883 , n31882 );
and ( n31884 , n31883 , n30421 );
and ( n31885 , n31238 , n30508 );
and ( n31886 , n31884 , n31885 );
and ( n31887 , n31088 , n30563 );
and ( n31888 , n31885 , n31887 );
and ( n31889 , n31884 , n31887 );
or ( n31890 , n31886 , n31888 , n31889 );
and ( n31891 , n31881 , n31890 );
xor ( n31892 , n31746 , n31747 );
xor ( n31893 , n31892 , n31749 );
and ( n31894 , n31890 , n31893 );
and ( n31895 , n31881 , n31893 );
or ( n31896 , n31891 , n31894 , n31895 );
and ( n31897 , n31874 , n31896 );
and ( n31898 , n31852 , n31897 );
xnor ( n31899 , n31712 , n31714 );
xnor ( n31900 , n31717 , n31719 );
and ( n31901 , n31899 , n31900 );
and ( n31902 , n31897 , n31901 );
and ( n31903 , n31852 , n31901 );
or ( n31904 , n31898 , n31902 , n31903 );
and ( n31905 , n31851 , n31904 );
and ( n31906 , n30464 , n31301 );
and ( n31907 , n31278 , n30461 );
and ( n31908 , n31906 , n31907 );
xor ( n31909 , n31682 , n31683 );
xor ( n31910 , n31909 , n31686 );
and ( n31911 , n31908 , n31910 );
xor ( n31912 , n31743 , n31752 );
and ( n31913 , n31910 , n31912 );
and ( n31914 , n31908 , n31912 );
or ( n31915 , n31911 , n31913 , n31914 );
xor ( n31916 , n31763 , n31770 );
xor ( n31917 , n31774 , n31777 );
and ( n31918 , n31916 , n31917 );
xor ( n31919 , n31780 , n31781 );
and ( n31920 , n31917 , n31919 );
and ( n31921 , n31916 , n31919 );
or ( n31922 , n31918 , n31920 , n31921 );
and ( n31923 , n31915 , n31922 );
and ( n31924 , n31464 , n30461 );
and ( n31925 , n31278 , n30473 );
and ( n31926 , n31924 , n31925 );
and ( n31927 , n30889 , n30700 );
and ( n31928 , n31925 , n31927 );
and ( n31929 , n31924 , n31927 );
or ( n31930 , n31926 , n31928 , n31929 );
and ( n31931 , n30464 , n31442 );
and ( n31932 , n30468 , n31301 );
and ( n31933 , n31931 , n31932 );
and ( n31934 , n30709 , n30898 );
and ( n31935 , n31932 , n31934 );
and ( n31936 , n31931 , n31934 );
or ( n31937 , n31933 , n31935 , n31936 );
and ( n31938 , n31930 , n31937 );
xor ( n31939 , n31757 , n31758 );
xor ( n31940 , n31939 , n31760 );
xor ( n31941 , n31764 , n31765 );
xor ( n31942 , n31941 , n31767 );
and ( n31943 , n31940 , n31942 );
and ( n31944 , n31938 , n31943 );
xnor ( n31945 , n31772 , n31773 );
xnor ( n31946 , n31775 , n31776 );
and ( n31947 , n31945 , n31946 );
and ( n31948 , n31943 , n31947 );
and ( n31949 , n31938 , n31947 );
or ( n31950 , n31944 , n31948 , n31949 );
and ( n31951 , n31922 , n31950 );
and ( n31952 , n31915 , n31950 );
or ( n31953 , n31923 , n31951 , n31952 );
and ( n31954 , n31904 , n31953 );
and ( n31955 , n31851 , n31953 );
or ( n31956 , n31905 , n31954 , n31955 );
and ( n31957 , n31842 , n31956 );
and ( n31958 , n31840 , n31956 );
or ( n31959 , n31843 , n31957 , n31958 );
and ( n31960 , n31837 , n31959 );
and ( n31961 , n31835 , n31959 );
or ( n31962 , n31838 , n31960 , n31961 );
xor ( n31963 , n31803 , n31805 );
xor ( n31964 , n31963 , n31808 );
and ( n31965 , n31962 , n31964 );
xor ( n31966 , n31692 , n31694 );
xor ( n31967 , n31966 , n31696 );
xor ( n31968 , n31701 , n31702 );
xor ( n31969 , n31968 , n31704 );
and ( n31970 , n31967 , n31969 );
xor ( n31971 , n31721 , n31724 );
xor ( n31972 , n31971 , n31728 );
and ( n31973 , n31969 , n31972 );
and ( n31974 , n31967 , n31972 );
or ( n31975 , n31970 , n31973 , n31974 );
xor ( n31976 , n31677 , n31699 );
xor ( n31977 , n31976 , n31707 );
and ( n31978 , n31975 , n31977 );
xor ( n31979 , n31731 , n31791 );
xor ( n31980 , n31979 , n31794 );
and ( n31981 , n31977 , n31980 );
and ( n31982 , n31975 , n31980 );
or ( n31983 , n31978 , n31981 , n31982 );
xor ( n31984 , n31710 , n31797 );
xor ( n31985 , n31984 , n31800 );
and ( n31986 , n31983 , n31985 );
xor ( n31987 , n31756 , n31785 );
xor ( n31988 , n31987 , n31788 );
xor ( n31989 , n31732 , n31733 );
xor ( n31990 , n31989 , n31753 );
xor ( n31991 , n31771 , n31778 );
xor ( n31992 , n31991 , n31782 );
and ( n31993 , n31990 , n31992 );
and ( n31994 , n31736 , n30439 );
and ( n31995 , n31607 , n30461 );
and ( n31996 , n31994 , n31995 );
and ( n31997 , n31238 , n30563 );
and ( n31998 , n31995 , n31997 );
and ( n31999 , n31994 , n31997 );
or ( n32000 , n31996 , n31998 , n31999 );
xor ( n32001 , n31853 , n31854 );
xor ( n32002 , n32001 , n31856 );
and ( n32003 , n32000 , n32002 );
xor ( n32004 , n31931 , n31932 );
xor ( n32005 , n32004 , n31934 );
and ( n32006 , n32002 , n32005 );
and ( n32007 , n32000 , n32005 );
or ( n32008 , n32003 , n32006 , n32007 );
xor ( n32009 , n31881 , n31890 );
xor ( n32010 , n32009 , n31893 );
and ( n32011 , n32008 , n32010 );
and ( n32012 , n30442 , n31745 );
and ( n32013 , n30464 , n31590 );
and ( n32014 , n32012 , n32013 );
and ( n32015 , n30558 , n31247 );
and ( n32016 , n32013 , n32015 );
and ( n32017 , n32012 , n32015 );
or ( n32018 , n32014 , n32016 , n32017 );
xor ( n32019 , n31875 , n31876 );
xor ( n32020 , n32019 , n31878 );
and ( n32021 , n32018 , n32020 );
xor ( n32022 , n31924 , n31925 );
xor ( n32023 , n32022 , n31927 );
and ( n32024 , n32020 , n32023 );
and ( n32025 , n32018 , n32023 );
or ( n32026 , n32021 , n32024 , n32025 );
xor ( n32027 , n31859 , n31868 );
xor ( n32028 , n32027 , n31871 );
and ( n32029 , n32026 , n32028 );
and ( n32030 , n32011 , n32029 );
and ( n32031 , n31992 , n32030 );
and ( n32032 , n31990 , n32030 );
or ( n32033 , n31993 , n32031 , n32032 );
and ( n32034 , n31988 , n32033 );
buf ( n32035 , n30799 );
buf ( n32036 , n15826 );
buf ( n32037 , n32036 );
and ( n32038 , n32035 , n32037 );
xor ( n32039 , n31906 , n31907 );
and ( n32040 , n32037 , n32039 );
and ( n32041 , n32035 , n32039 );
or ( n32042 , n32038 , n32040 , n32041 );
xor ( n32043 , n31874 , n31896 );
and ( n32044 , n32042 , n32043 );
xor ( n32045 , n31899 , n31900 );
and ( n32046 , n32043 , n32045 );
and ( n32047 , n32042 , n32045 );
or ( n32048 , n32044 , n32046 , n32047 );
xor ( n32049 , n31930 , n31937 );
xor ( n32050 , n31940 , n31942 );
and ( n32051 , n32049 , n32050 );
xor ( n32052 , n31945 , n31946 );
and ( n32053 , n32050 , n32052 );
and ( n32054 , n32049 , n32052 );
or ( n32055 , n32051 , n32053 , n32054 );
buf ( n32056 , n1238 );
buf ( n32057 , n32056 );
and ( n32058 , n32057 , n30421 );
and ( n32059 , n31883 , n30424 );
and ( n32060 , n32058 , n32059 );
and ( n32061 , n31084 , n30700 );
and ( n32062 , n32059 , n32061 );
and ( n32063 , n32058 , n32061 );
or ( n32064 , n32060 , n32062 , n32063 );
buf ( n32065 , n1238 );
buf ( n32066 , n32065 );
and ( n32067 , n30413 , n32066 );
and ( n32068 , n30419 , n31861 );
and ( n32069 , n32067 , n32068 );
and ( n32070 , n30709 , n31076 );
and ( n32071 , n32068 , n32070 );
and ( n32072 , n32067 , n32070 );
or ( n32073 , n32069 , n32071 , n32072 );
and ( n32074 , n32064 , n32073 );
and ( n32075 , n31088 , n30592 );
and ( n32076 , n30889 , n30791 );
or ( n32077 , n32075 , n32076 );
and ( n32078 , n30603 , n31073 );
and ( n32079 , n30799 , n30898 );
or ( n32080 , n32078 , n32079 );
and ( n32081 , n32077 , n32080 );
and ( n32082 , n32074 , n32081 );
xor ( n32083 , n32035 , n32037 );
xor ( n32084 , n32083 , n32039 );
and ( n32085 , n32081 , n32084 );
and ( n32086 , n32074 , n32084 );
or ( n32087 , n32082 , n32085 , n32086 );
and ( n32088 , n32055 , n32087 );
xor ( n32089 , n31908 , n31910 );
xor ( n32090 , n32089 , n31912 );
and ( n32091 , n32087 , n32090 );
and ( n32092 , n32055 , n32090 );
or ( n32093 , n32088 , n32091 , n32092 );
and ( n32094 , n32048 , n32093 );
xor ( n32095 , n31845 , n31846 );
xor ( n32096 , n32095 , n31848 );
and ( n32097 , n32093 , n32096 );
and ( n32098 , n32048 , n32096 );
or ( n32099 , n32094 , n32097 , n32098 );
and ( n32100 , n32033 , n32099 );
and ( n32101 , n31988 , n32099 );
or ( n32102 , n32034 , n32100 , n32101 );
xor ( n32103 , n31840 , n31842 );
xor ( n32104 , n32103 , n31956 );
and ( n32105 , n32102 , n32104 );
xor ( n32106 , n31975 , n31977 );
xor ( n32107 , n32106 , n31980 );
and ( n32108 , n32104 , n32107 );
and ( n32109 , n32102 , n32107 );
or ( n32110 , n32105 , n32108 , n32109 );
and ( n32111 , n31985 , n32110 );
and ( n32112 , n31983 , n32110 );
or ( n32113 , n31986 , n32111 , n32112 );
and ( n32114 , n31964 , n32113 );
and ( n32115 , n31962 , n32113 );
or ( n32116 , n31965 , n32114 , n32115 );
and ( n32117 , n31833 , n32116 );
xor ( n32118 , n31833 , n32116 );
xor ( n32119 , n31962 , n31964 );
xor ( n32120 , n32119 , n32113 );
xor ( n32121 , n31835 , n31837 );
xor ( n32122 , n32121 , n31959 );
xor ( n32123 , n31983 , n31985 );
xor ( n32124 , n32123 , n32110 );
and ( n32125 , n32122 , n32124 );
xor ( n32126 , n31851 , n31904 );
xor ( n32127 , n32126 , n31953 );
xor ( n32128 , n31967 , n31969 );
xor ( n32129 , n32128 , n31972 );
and ( n32130 , n32127 , n32129 );
xor ( n32131 , n31852 , n31897 );
xor ( n32132 , n32131 , n31901 );
xor ( n32133 , n31915 , n31922 );
xor ( n32134 , n32133 , n31950 );
and ( n32135 , n32132 , n32134 );
xor ( n32136 , n31916 , n31917 );
xor ( n32137 , n32136 , n31919 );
xor ( n32138 , n31938 , n31943 );
xor ( n32139 , n32138 , n31947 );
and ( n32140 , n32137 , n32139 );
xor ( n32141 , n32011 , n32029 );
and ( n32142 , n32139 , n32141 );
and ( n32143 , n32137 , n32141 );
or ( n32144 , n32140 , n32142 , n32143 );
and ( n32145 , n32134 , n32144 );
and ( n32146 , n32132 , n32144 );
or ( n32147 , n32135 , n32145 , n32146 );
and ( n32148 , n32129 , n32147 );
and ( n32149 , n32127 , n32147 );
or ( n32150 , n32130 , n32148 , n32149 );
xor ( n32151 , n32102 , n32104 );
xor ( n32152 , n32151 , n32107 );
and ( n32153 , n32150 , n32152 );
buf ( n32154 , n1239 );
buf ( n32155 , n32154 );
and ( n32156 , n32155 , n30421 );
and ( n32157 , n32057 , n30424 );
and ( n32158 , n32156 , n32157 );
and ( n32159 , n31238 , n30592 );
and ( n32160 , n32157 , n32159 );
and ( n32161 , n32156 , n32159 );
or ( n32162 , n32158 , n32160 , n32161 );
and ( n32163 , n30468 , n31442 );
and ( n32164 , n32162 , n32163 );
and ( n32165 , n30503 , n31301 );
and ( n32166 , n32163 , n32165 );
and ( n32167 , n32162 , n32165 );
or ( n32168 , n32164 , n32166 , n32167 );
xor ( n32169 , n31862 , n31863 );
xor ( n32170 , n32169 , n31865 );
or ( n32171 , n32168 , n32170 );
buf ( n32172 , n1239 );
buf ( n32173 , n32172 );
and ( n32174 , n30413 , n32173 );
and ( n32175 , n30419 , n32066 );
and ( n32176 , n32174 , n32175 );
and ( n32177 , n30603 , n31247 );
and ( n32178 , n32175 , n32177 );
and ( n32179 , n32174 , n32177 );
or ( n32180 , n32176 , n32178 , n32179 );
and ( n32181 , n31464 , n30473 );
and ( n32182 , n32180 , n32181 );
and ( n32183 , n31278 , n30508 );
and ( n32184 , n32181 , n32183 );
and ( n32185 , n32180 , n32183 );
or ( n32186 , n32182 , n32184 , n32185 );
xor ( n32187 , n31884 , n31885 );
xor ( n32188 , n32187 , n31887 );
or ( n32189 , n32186 , n32188 );
and ( n32190 , n32171 , n32189 );
xor ( n32191 , n32008 , n32010 );
xor ( n32192 , n32026 , n32028 );
and ( n32193 , n32191 , n32192 );
and ( n32194 , n32190 , n32193 );
xnor ( n32195 , n32075 , n32076 );
xnor ( n32196 , n32078 , n32079 );
and ( n32197 , n32195 , n32196 );
buf ( n32198 , n15829 );
buf ( n32199 , n32198 );
or ( n32200 , n32197 , n32199 );
xor ( n32201 , n32067 , n32068 );
xor ( n32202 , n32201 , n32070 );
xor ( n32203 , n32012 , n32013 );
xor ( n32204 , n32203 , n32015 );
or ( n32205 , n32202 , n32204 );
xor ( n32206 , n32058 , n32059 );
xor ( n32207 , n32206 , n32061 );
xor ( n32208 , n31994 , n31995 );
xor ( n32209 , n32208 , n31997 );
or ( n32210 , n32207 , n32209 );
and ( n32211 , n32205 , n32210 );
and ( n32212 , n32200 , n32211 );
xor ( n32213 , n32018 , n32020 );
xor ( n32214 , n32213 , n32023 );
xor ( n32215 , n32000 , n32002 );
xor ( n32216 , n32215 , n32005 );
and ( n32217 , n32214 , n32216 );
and ( n32218 , n32211 , n32217 );
and ( n32219 , n32200 , n32217 );
or ( n32220 , n32212 , n32218 , n32219 );
and ( n32221 , n32193 , n32220 );
and ( n32222 , n32190 , n32220 );
or ( n32223 , n32194 , n32221 , n32222 );
and ( n32224 , n30803 , n30791 );
and ( n32225 , n30799 , n30788 );
and ( n32226 , n32224 , n32225 );
xor ( n32227 , n32064 , n32073 );
and ( n32228 , n32225 , n32227 );
and ( n32229 , n32224 , n32227 );
or ( n32230 , n32226 , n32228 , n32229 );
xor ( n32231 , n32077 , n32080 );
and ( n32232 , n31883 , n30439 );
and ( n32233 , n31736 , n30461 );
and ( n32234 , n32232 , n32233 );
and ( n32235 , n31088 , n30700 );
and ( n32236 , n32233 , n32235 );
and ( n32237 , n32232 , n32235 );
or ( n32238 , n32234 , n32236 , n32237 );
and ( n32239 , n30442 , n31861 );
and ( n32240 , n30464 , n31745 );
and ( n32241 , n32239 , n32240 );
and ( n32242 , n30709 , n31073 );
and ( n32243 , n32240 , n32242 );
and ( n32244 , n32239 , n32242 );
or ( n32245 , n32241 , n32243 , n32244 );
and ( n32246 , n32238 , n32245 );
and ( n32247 , n32231 , n32246 );
and ( n32248 , n31607 , n30473 );
and ( n32249 , n31464 , n30508 );
and ( n32250 , n32248 , n32249 );
and ( n32251 , n31084 , n30791 );
and ( n32252 , n32249 , n32251 );
and ( n32253 , n32248 , n32251 );
or ( n32254 , n32250 , n32252 , n32253 );
and ( n32255 , n30468 , n31590 );
and ( n32256 , n30503 , n31442 );
and ( n32257 , n32255 , n32256 );
and ( n32258 , n30799 , n31076 );
and ( n32259 , n32256 , n32258 );
and ( n32260 , n32255 , n32258 );
or ( n32261 , n32257 , n32259 , n32260 );
and ( n32262 , n32254 , n32261 );
and ( n32263 , n32246 , n32262 );
and ( n32264 , n32231 , n32262 );
or ( n32265 , n32247 , n32263 , n32264 );
and ( n32266 , n32230 , n32265 );
xor ( n32267 , n32049 , n32050 );
xor ( n32268 , n32267 , n32052 );
and ( n32269 , n32265 , n32268 );
and ( n32270 , n32230 , n32268 );
or ( n32271 , n32266 , n32269 , n32270 );
xor ( n32272 , n32042 , n32043 );
xor ( n32273 , n32272 , n32045 );
and ( n32274 , n32271 , n32273 );
xor ( n32275 , n32055 , n32087 );
xor ( n32276 , n32275 , n32090 );
and ( n32277 , n32273 , n32276 );
and ( n32278 , n32271 , n32276 );
or ( n32279 , n32274 , n32277 , n32278 );
and ( n32280 , n32223 , n32279 );
xor ( n32281 , n31990 , n31992 );
xor ( n32282 , n32281 , n32030 );
and ( n32283 , n32279 , n32282 );
and ( n32284 , n32223 , n32282 );
or ( n32285 , n32280 , n32283 , n32284 );
xor ( n32286 , n31988 , n32033 );
xor ( n32287 , n32286 , n32099 );
and ( n32288 , n32285 , n32287 );
xor ( n32289 , n32048 , n32093 );
xor ( n32290 , n32289 , n32096 );
xor ( n32291 , n32074 , n32081 );
xor ( n32292 , n32291 , n32084 );
xor ( n32293 , n32171 , n32189 );
and ( n32294 , n32292 , n32293 );
xor ( n32295 , n32191 , n32192 );
and ( n32296 , n32293 , n32295 );
and ( n32297 , n32292 , n32295 );
or ( n32298 , n32294 , n32296 , n32297 );
xnor ( n32299 , n32168 , n32170 );
xnor ( n32300 , n32186 , n32188 );
and ( n32301 , n32299 , n32300 );
buf ( n32302 , n30803 );
buf ( n32303 , n15832 );
buf ( n32304 , n32303 );
and ( n32305 , n32302 , n32304 );
and ( n32306 , n30889 , n30788 );
and ( n32307 , n30803 , n30898 );
and ( n32308 , n32306 , n32307 );
buf ( n32309 , n15835 );
buf ( n32310 , n32309 );
and ( n32311 , n32307 , n32310 );
and ( n32312 , n32306 , n32310 );
or ( n32313 , n32308 , n32311 , n32312 );
and ( n32314 , n32304 , n32313 );
and ( n32315 , n32302 , n32313 );
or ( n32316 , n32305 , n32314 , n32315 );
xnor ( n32317 , n32197 , n32199 );
and ( n32318 , n32316 , n32317 );
xor ( n32319 , n32205 , n32210 );
and ( n32320 , n32317 , n32319 );
and ( n32321 , n32316 , n32319 );
or ( n32322 , n32318 , n32320 , n32321 );
and ( n32323 , n32301 , n32322 );
xor ( n32324 , n32214 , n32216 );
xor ( n32325 , n32232 , n32233 );
xor ( n32326 , n32325 , n32235 );
xor ( n32327 , n32248 , n32249 );
xor ( n32328 , n32327 , n32251 );
and ( n32329 , n32326 , n32328 );
xor ( n32330 , n32156 , n32157 );
xor ( n32331 , n32330 , n32159 );
and ( n32332 , n32328 , n32331 );
and ( n32333 , n32326 , n32331 );
or ( n32334 , n32329 , n32332 , n32333 );
xor ( n32335 , n32239 , n32240 );
xor ( n32336 , n32335 , n32242 );
xor ( n32337 , n32255 , n32256 );
xor ( n32338 , n32337 , n32258 );
and ( n32339 , n32336 , n32338 );
xor ( n32340 , n32174 , n32175 );
xor ( n32341 , n32340 , n32177 );
and ( n32342 , n32338 , n32341 );
and ( n32343 , n32336 , n32341 );
or ( n32344 , n32339 , n32342 , n32343 );
and ( n32345 , n32334 , n32344 );
and ( n32346 , n32324 , n32345 );
buf ( n32347 , n1240 );
buf ( n32348 , n32347 );
and ( n32349 , n30413 , n32348 );
and ( n32350 , n30503 , n31590 );
and ( n32351 , n32349 , n32350 );
and ( n32352 , n30558 , n31442 );
and ( n32353 , n32350 , n32352 );
and ( n32354 , n32349 , n32352 );
or ( n32355 , n32351 , n32353 , n32354 );
and ( n32356 , n30464 , n31861 );
and ( n32357 , n30468 , n31745 );
and ( n32358 , n32356 , n32357 );
and ( n32359 , n30603 , n31301 );
and ( n32360 , n32357 , n32359 );
and ( n32361 , n32356 , n32359 );
or ( n32362 , n32358 , n32360 , n32361 );
or ( n32363 , n32355 , n32362 );
buf ( n32364 , n1240 );
buf ( n32365 , n32364 );
and ( n32366 , n32365 , n30421 );
and ( n32367 , n31607 , n30508 );
and ( n32368 , n32366 , n32367 );
and ( n32369 , n31464 , n30563 );
and ( n32370 , n32367 , n32369 );
and ( n32371 , n32366 , n32369 );
or ( n32372 , n32368 , n32370 , n32371 );
and ( n32373 , n31883 , n30461 );
and ( n32374 , n31736 , n30473 );
and ( n32375 , n32373 , n32374 );
and ( n32376 , n31278 , n30592 );
and ( n32377 , n32374 , n32376 );
and ( n32378 , n32373 , n32376 );
or ( n32379 , n32375 , n32377 , n32378 );
or ( n32380 , n32372 , n32379 );
and ( n32381 , n32363 , n32380 );
and ( n32382 , n32345 , n32381 );
and ( n32383 , n32324 , n32381 );
or ( n32384 , n32346 , n32382 , n32383 );
and ( n32385 , n32322 , n32384 );
and ( n32386 , n32301 , n32384 );
or ( n32387 , n32323 , n32385 , n32386 );
and ( n32388 , n32298 , n32387 );
and ( n32389 , n30419 , n32173 );
and ( n32390 , n30442 , n32066 );
and ( n32391 , n32389 , n32390 );
and ( n32392 , n30799 , n31073 );
and ( n32393 , n32390 , n32392 );
and ( n32394 , n32389 , n32392 );
or ( n32395 , n32391 , n32393 , n32394 );
not ( n32396 , n32395 );
and ( n32397 , n31278 , n30563 );
and ( n32398 , n32396 , n32397 );
and ( n32399 , n32155 , n30424 );
and ( n32400 , n32057 , n30439 );
and ( n32401 , n32399 , n32400 );
and ( n32402 , n31088 , n30791 );
and ( n32403 , n32400 , n32402 );
and ( n32404 , n32399 , n32402 );
or ( n32405 , n32401 , n32403 , n32404 );
not ( n32406 , n32405 );
and ( n32407 , n30558 , n31301 );
and ( n32408 , n32406 , n32407 );
and ( n32409 , n32398 , n32408 );
buf ( n32410 , n32395 );
buf ( n32411 , n32405 );
and ( n32412 , n32410 , n32411 );
and ( n32413 , n32409 , n32412 );
xor ( n32414 , n32180 , n32181 );
xor ( n32415 , n32414 , n32183 );
xor ( n32416 , n32162 , n32163 );
xor ( n32417 , n32416 , n32165 );
and ( n32418 , n32415 , n32417 );
and ( n32419 , n32412 , n32418 );
and ( n32420 , n32409 , n32418 );
or ( n32421 , n32413 , n32419 , n32420 );
xnor ( n32422 , n32202 , n32204 );
xnor ( n32423 , n32207 , n32209 );
and ( n32424 , n32422 , n32423 );
xor ( n32425 , n32238 , n32245 );
xor ( n32426 , n32254 , n32261 );
and ( n32427 , n32425 , n32426 );
xor ( n32428 , n32195 , n32196 );
and ( n32429 , n32426 , n32428 );
and ( n32430 , n32425 , n32428 );
or ( n32431 , n32427 , n32429 , n32430 );
and ( n32432 , n32424 , n32431 );
xor ( n32433 , n32224 , n32225 );
xor ( n32434 , n32433 , n32227 );
and ( n32435 , n32431 , n32434 );
and ( n32436 , n32424 , n32434 );
or ( n32437 , n32432 , n32435 , n32436 );
and ( n32438 , n32421 , n32437 );
xor ( n32439 , n32200 , n32211 );
xor ( n32440 , n32439 , n32217 );
and ( n32441 , n32437 , n32440 );
and ( n32442 , n32421 , n32440 );
or ( n32443 , n32438 , n32441 , n32442 );
and ( n32444 , n32387 , n32443 );
and ( n32445 , n32298 , n32443 );
or ( n32446 , n32388 , n32444 , n32445 );
and ( n32447 , n32290 , n32446 );
xor ( n32448 , n32137 , n32139 );
xor ( n32449 , n32448 , n32141 );
xor ( n32450 , n32190 , n32193 );
xor ( n32451 , n32450 , n32220 );
and ( n32452 , n32449 , n32451 );
xor ( n32453 , n32271 , n32273 );
xor ( n32454 , n32453 , n32276 );
and ( n32455 , n32451 , n32454 );
and ( n32456 , n32449 , n32454 );
or ( n32457 , n32452 , n32455 , n32456 );
and ( n32458 , n32446 , n32457 );
and ( n32459 , n32290 , n32457 );
or ( n32460 , n32447 , n32458 , n32459 );
and ( n32461 , n32287 , n32460 );
and ( n32462 , n32285 , n32460 );
or ( n32463 , n32288 , n32461 , n32462 );
and ( n32464 , n32152 , n32463 );
and ( n32465 , n32150 , n32463 );
or ( n32466 , n32153 , n32464 , n32465 );
and ( n32467 , n32124 , n32466 );
and ( n32468 , n32122 , n32466 );
or ( n32469 , n32125 , n32467 , n32468 );
and ( n32470 , n32120 , n32469 );
xor ( n32471 , n32120 , n32469 );
xor ( n32472 , n32122 , n32124 );
xor ( n32473 , n32472 , n32466 );
xor ( n32474 , n32127 , n32129 );
xor ( n32475 , n32474 , n32147 );
xor ( n32476 , n32132 , n32134 );
xor ( n32477 , n32476 , n32144 );
xor ( n32478 , n32223 , n32279 );
xor ( n32479 , n32478 , n32282 );
and ( n32480 , n32477 , n32479 );
xor ( n32481 , n32230 , n32265 );
xor ( n32482 , n32481 , n32268 );
xor ( n32483 , n32231 , n32246 );
xor ( n32484 , n32483 , n32262 );
xor ( n32485 , n32299 , n32300 );
and ( n32486 , n32484 , n32485 );
and ( n32487 , n31238 , n30700 );
and ( n32488 , n31084 , n30788 );
or ( n32489 , n32487 , n32488 );
and ( n32490 , n30709 , n31247 );
and ( n32491 , n30803 , n31076 );
or ( n32492 , n32490 , n32491 );
and ( n32493 , n32489 , n32492 );
xor ( n32494 , n32302 , n32304 );
xor ( n32495 , n32494 , n32313 );
and ( n32496 , n32493 , n32495 );
xor ( n32497 , n32334 , n32344 );
and ( n32498 , n32495 , n32497 );
and ( n32499 , n32493 , n32497 );
or ( n32500 , n32496 , n32498 , n32499 );
and ( n32501 , n32485 , n32500 );
and ( n32502 , n32484 , n32500 );
or ( n32503 , n32486 , n32501 , n32502 );
and ( n32504 , n32482 , n32503 );
xor ( n32505 , n32363 , n32380 );
xor ( n32506 , n32398 , n32408 );
and ( n32507 , n32505 , n32506 );
xor ( n32508 , n32410 , n32411 );
and ( n32509 , n32506 , n32508 );
and ( n32510 , n32505 , n32508 );
or ( n32511 , n32507 , n32509 , n32510 );
xor ( n32512 , n32415 , n32417 );
xor ( n32513 , n32422 , n32423 );
and ( n32514 , n32512 , n32513 );
and ( n32515 , n30464 , n32066 );
and ( n32516 , n30468 , n31861 );
and ( n32517 , n32515 , n32516 );
and ( n32518 , n30799 , n31247 );
and ( n32519 , n32516 , n32518 );
and ( n32520 , n32515 , n32518 );
or ( n32521 , n32517 , n32519 , n32520 );
xor ( n32522 , n32366 , n32367 );
xor ( n32523 , n32522 , n32369 );
and ( n32524 , n32521 , n32523 );
xor ( n32525 , n32399 , n32400 );
xor ( n32526 , n32525 , n32402 );
and ( n32527 , n32523 , n32526 );
and ( n32528 , n32521 , n32526 );
or ( n32529 , n32524 , n32527 , n32528 );
and ( n32530 , n32057 , n30461 );
and ( n32531 , n31883 , n30473 );
and ( n32532 , n32530 , n32531 );
and ( n32533 , n31238 , n30791 );
and ( n32534 , n32531 , n32533 );
and ( n32535 , n32530 , n32533 );
or ( n32536 , n32532 , n32534 , n32535 );
xor ( n32537 , n32349 , n32350 );
xor ( n32538 , n32537 , n32352 );
and ( n32539 , n32536 , n32538 );
xor ( n32540 , n32389 , n32390 );
xor ( n32541 , n32540 , n32392 );
and ( n32542 , n32538 , n32541 );
and ( n32543 , n32536 , n32541 );
or ( n32544 , n32539 , n32542 , n32543 );
and ( n32545 , n32529 , n32544 );
and ( n32546 , n32513 , n32545 );
and ( n32547 , n32512 , n32545 );
or ( n32548 , n32514 , n32546 , n32547 );
and ( n32549 , n32511 , n32548 );
and ( n32550 , n30503 , n31745 );
and ( n32551 , n30558 , n31590 );
and ( n32552 , n32550 , n32551 );
and ( n32553 , n30803 , n31073 );
and ( n32554 , n32551 , n32553 );
and ( n32555 , n32550 , n32553 );
or ( n32556 , n32552 , n32554 , n32555 );
and ( n32557 , n30419 , n32348 );
and ( n32558 , n30442 , n32173 );
and ( n32559 , n32557 , n32558 );
and ( n32560 , n30709 , n31301 );
and ( n32561 , n32558 , n32560 );
and ( n32562 , n32557 , n32560 );
or ( n32563 , n32559 , n32561 , n32562 );
or ( n32564 , n32556 , n32563 );
and ( n32565 , n31736 , n30508 );
and ( n32566 , n31607 , n30563 );
and ( n32567 , n32565 , n32566 );
and ( n32568 , n31088 , n30788 );
and ( n32569 , n32566 , n32568 );
and ( n32570 , n32565 , n32568 );
or ( n32571 , n32567 , n32569 , n32570 );
and ( n32572 , n32365 , n30424 );
and ( n32573 , n32155 , n30439 );
and ( n32574 , n32572 , n32573 );
and ( n32575 , n31278 , n30700 );
and ( n32576 , n32573 , n32575 );
and ( n32577 , n32572 , n32575 );
or ( n32578 , n32574 , n32576 , n32577 );
or ( n32579 , n32571 , n32578 );
and ( n32580 , n32564 , n32579 );
xor ( n32581 , n32326 , n32328 );
xor ( n32582 , n32581 , n32331 );
xor ( n32583 , n32336 , n32338 );
xor ( n32584 , n32583 , n32341 );
and ( n32585 , n32582 , n32584 );
and ( n32586 , n32580 , n32585 );
xnor ( n32587 , n32355 , n32362 );
xnor ( n32588 , n32372 , n32379 );
and ( n32589 , n32587 , n32588 );
and ( n32590 , n32585 , n32589 );
and ( n32591 , n32580 , n32589 );
or ( n32592 , n32586 , n32590 , n32591 );
and ( n32593 , n32548 , n32592 );
and ( n32594 , n32511 , n32592 );
or ( n32595 , n32549 , n32593 , n32594 );
and ( n32596 , n32503 , n32595 );
and ( n32597 , n32482 , n32595 );
or ( n32598 , n32504 , n32596 , n32597 );
xor ( n32599 , n32396 , n32397 );
xor ( n32600 , n32406 , n32407 );
and ( n32601 , n32599 , n32600 );
xor ( n32602 , n32306 , n32307 );
xor ( n32603 , n32602 , n32310 );
xor ( n32604 , n32489 , n32492 );
and ( n32605 , n32603 , n32604 );
xnor ( n32606 , n32487 , n32488 );
xnor ( n32607 , n32490 , n32491 );
and ( n32608 , n32606 , n32607 );
and ( n32609 , n32604 , n32608 );
and ( n32610 , n32603 , n32608 );
or ( n32611 , n32605 , n32609 , n32610 );
and ( n32612 , n32601 , n32611 );
xor ( n32613 , n32425 , n32426 );
xor ( n32614 , n32613 , n32428 );
and ( n32615 , n32611 , n32614 );
and ( n32616 , n32601 , n32614 );
or ( n32617 , n32612 , n32615 , n32616 );
xor ( n32618 , n32316 , n32317 );
xor ( n32619 , n32618 , n32319 );
and ( n32620 , n32617 , n32619 );
xor ( n32621 , n32324 , n32345 );
xor ( n32622 , n32621 , n32381 );
and ( n32623 , n32619 , n32622 );
and ( n32624 , n32617 , n32622 );
or ( n32625 , n32620 , n32623 , n32624 );
xor ( n32626 , n32292 , n32293 );
xor ( n32627 , n32626 , n32295 );
and ( n32628 , n32625 , n32627 );
xor ( n32629 , n32301 , n32322 );
xor ( n32630 , n32629 , n32384 );
and ( n32631 , n32627 , n32630 );
and ( n32632 , n32625 , n32630 );
or ( n32633 , n32628 , n32631 , n32632 );
and ( n32634 , n32598 , n32633 );
xor ( n32635 , n32298 , n32387 );
xor ( n32636 , n32635 , n32443 );
and ( n32637 , n32633 , n32636 );
and ( n32638 , n32598 , n32636 );
or ( n32639 , n32634 , n32637 , n32638 );
and ( n32640 , n32479 , n32639 );
and ( n32641 , n32477 , n32639 );
or ( n32642 , n32480 , n32640 , n32641 );
and ( n32643 , n32475 , n32642 );
xor ( n32644 , n32285 , n32287 );
xor ( n32645 , n32644 , n32460 );
and ( n32646 , n32642 , n32645 );
and ( n32647 , n32475 , n32645 );
or ( n32648 , n32643 , n32646 , n32647 );
xor ( n32649 , n32150 , n32152 );
xor ( n32650 , n32649 , n32463 );
and ( n32651 , n32648 , n32650 );
xor ( n32652 , n32290 , n32446 );
xor ( n32653 , n32652 , n32457 );
xor ( n32654 , n32449 , n32451 );
xor ( n32655 , n32654 , n32454 );
xor ( n32656 , n32421 , n32437 );
xor ( n32657 , n32656 , n32440 );
xor ( n32658 , n32409 , n32412 );
xor ( n32659 , n32658 , n32418 );
xor ( n32660 , n32424 , n32431 );
xor ( n32661 , n32660 , n32434 );
and ( n32662 , n32659 , n32661 );
and ( n32663 , n32057 , n30473 );
and ( n32664 , n31883 , n30508 );
and ( n32665 , n32663 , n32664 );
and ( n32666 , n31464 , n30700 );
and ( n32667 , n32664 , n32666 );
and ( n32668 , n32663 , n32666 );
or ( n32669 , n32665 , n32667 , n32668 );
buf ( n32670 , n1241 );
buf ( n32671 , n32670 );
and ( n32672 , n30413 , n32671 );
and ( n32673 , n32669 , n32672 );
and ( n32674 , n30603 , n31442 );
and ( n32675 , n32672 , n32674 );
and ( n32676 , n32669 , n32674 );
or ( n32677 , n32673 , n32675 , n32676 );
xor ( n32678 , n32356 , n32357 );
xor ( n32679 , n32678 , n32359 );
or ( n32680 , n32677 , n32679 );
and ( n32681 , n30468 , n32066 );
and ( n32682 , n30503 , n31861 );
and ( n32683 , n32681 , n32682 );
and ( n32684 , n30709 , n31442 );
and ( n32685 , n32682 , n32684 );
and ( n32686 , n32681 , n32684 );
or ( n32687 , n32683 , n32685 , n32686 );
buf ( n32688 , n1241 );
buf ( n32689 , n32688 );
and ( n32690 , n32689 , n30421 );
and ( n32691 , n32687 , n32690 );
and ( n32692 , n31464 , n30592 );
and ( n32693 , n32690 , n32692 );
and ( n32694 , n32687 , n32692 );
or ( n32695 , n32691 , n32693 , n32694 );
xor ( n32696 , n32373 , n32374 );
xor ( n32697 , n32696 , n32376 );
or ( n32698 , n32695 , n32697 );
and ( n32699 , n32680 , n32698 );
xor ( n32700 , n32529 , n32544 );
xor ( n32701 , n32564 , n32579 );
and ( n32702 , n32700 , n32701 );
xor ( n32703 , n32582 , n32584 );
and ( n32704 , n32701 , n32703 );
and ( n32705 , n32700 , n32703 );
or ( n32706 , n32702 , n32704 , n32705 );
and ( n32707 , n32699 , n32706 );
xor ( n32708 , n32587 , n32588 );
xor ( n32709 , n32599 , n32600 );
and ( n32710 , n32708 , n32709 );
and ( n32711 , n30442 , n32348 );
and ( n32712 , n30464 , n32173 );
and ( n32713 , n32711 , n32712 );
and ( n32714 , n30803 , n31247 );
and ( n32715 , n32712 , n32714 );
and ( n32716 , n32711 , n32714 );
or ( n32717 , n32713 , n32715 , n32716 );
buf ( n32718 , n1242 );
buf ( n32719 , n32718 );
and ( n32720 , n30413 , n32719 );
and ( n32721 , n30419 , n32671 );
and ( n32722 , n32720 , n32721 );
and ( n32723 , n30603 , n31590 );
and ( n32724 , n32721 , n32723 );
and ( n32725 , n32720 , n32723 );
or ( n32726 , n32722 , n32724 , n32725 );
or ( n32727 , n32717 , n32726 );
and ( n32728 , n32365 , n30439 );
and ( n32729 , n32155 , n30461 );
and ( n32730 , n32728 , n32729 );
and ( n32731 , n31238 , n30788 );
and ( n32732 , n32729 , n32731 );
and ( n32733 , n32728 , n32731 );
or ( n32734 , n32730 , n32732 , n32733 );
buf ( n32735 , n1242 );
buf ( n32736 , n32735 );
and ( n32737 , n32736 , n30421 );
and ( n32738 , n32689 , n30424 );
and ( n32739 , n32737 , n32738 );
and ( n32740 , n31607 , n30592 );
and ( n32741 , n32738 , n32740 );
and ( n32742 , n32737 , n32740 );
or ( n32743 , n32739 , n32741 , n32742 );
or ( n32744 , n32734 , n32743 );
and ( n32745 , n32727 , n32744 );
and ( n32746 , n32709 , n32745 );
and ( n32747 , n32708 , n32745 );
or ( n32748 , n32710 , n32746 , n32747 );
and ( n32749 , n32706 , n32748 );
and ( n32750 , n32699 , n32748 );
or ( n32751 , n32707 , n32749 , n32750 );
and ( n32752 , n32661 , n32751 );
and ( n32753 , n32659 , n32751 );
or ( n32754 , n32662 , n32752 , n32753 );
and ( n32755 , n32657 , n32754 );
xor ( n32756 , n32550 , n32551 );
xor ( n32757 , n32756 , n32553 );
xor ( n32758 , n32515 , n32516 );
xor ( n32759 , n32758 , n32518 );
or ( n32760 , n32757 , n32759 );
xor ( n32761 , n32565 , n32566 );
xor ( n32762 , n32761 , n32568 );
xor ( n32763 , n32530 , n32531 );
xor ( n32764 , n32763 , n32533 );
or ( n32765 , n32762 , n32764 );
and ( n32766 , n32760 , n32765 );
xor ( n32767 , n32521 , n32523 );
xor ( n32768 , n32767 , n32526 );
xor ( n32769 , n32536 , n32538 );
xor ( n32770 , n32769 , n32541 );
and ( n32771 , n32768 , n32770 );
and ( n32772 , n32766 , n32771 );
xnor ( n32773 , n32556 , n32563 );
xnor ( n32774 , n32571 , n32578 );
and ( n32775 , n32773 , n32774 );
and ( n32776 , n32771 , n32775 );
and ( n32777 , n32766 , n32775 );
or ( n32778 , n32772 , n32776 , n32777 );
xor ( n32779 , n32493 , n32495 );
xor ( n32780 , n32779 , n32497 );
and ( n32781 , n32778 , n32780 );
xor ( n32782 , n32505 , n32506 );
xor ( n32783 , n32782 , n32508 );
and ( n32784 , n32780 , n32783 );
and ( n32785 , n32778 , n32783 );
or ( n32786 , n32781 , n32784 , n32785 );
xor ( n32787 , n32512 , n32513 );
xor ( n32788 , n32787 , n32545 );
xor ( n32789 , n32580 , n32585 );
xor ( n32790 , n32789 , n32589 );
and ( n32791 , n32788 , n32790 );
xor ( n32792 , n32601 , n32611 );
xor ( n32793 , n32792 , n32614 );
and ( n32794 , n32790 , n32793 );
and ( n32795 , n32788 , n32793 );
or ( n32796 , n32791 , n32794 , n32795 );
and ( n32797 , n32786 , n32796 );
xor ( n32798 , n32484 , n32485 );
xor ( n32799 , n32798 , n32500 );
and ( n32800 , n32796 , n32799 );
and ( n32801 , n32786 , n32799 );
or ( n32802 , n32797 , n32800 , n32801 );
and ( n32803 , n32754 , n32802 );
and ( n32804 , n32657 , n32802 );
or ( n32805 , n32755 , n32803 , n32804 );
and ( n32806 , n32655 , n32805 );
xor ( n32807 , n32598 , n32633 );
xor ( n32808 , n32807 , n32636 );
and ( n32809 , n32805 , n32808 );
and ( n32810 , n32655 , n32808 );
or ( n32811 , n32806 , n32809 , n32810 );
and ( n32812 , n32653 , n32811 );
xor ( n32813 , n32477 , n32479 );
xor ( n32814 , n32813 , n32639 );
and ( n32815 , n32811 , n32814 );
and ( n32816 , n32653 , n32814 );
or ( n32817 , n32812 , n32815 , n32816 );
xor ( n32818 , n32475 , n32642 );
xor ( n32819 , n32818 , n32645 );
and ( n32820 , n32817 , n32819 );
xor ( n32821 , n32653 , n32811 );
xor ( n32822 , n32821 , n32814 );
xor ( n32823 , n32482 , n32503 );
xor ( n32824 , n32823 , n32595 );
xor ( n32825 , n32625 , n32627 );
xor ( n32826 , n32825 , n32630 );
and ( n32827 , n32824 , n32826 );
xor ( n32828 , n32511 , n32548 );
xor ( n32829 , n32828 , n32592 );
xor ( n32830 , n32617 , n32619 );
xor ( n32831 , n32830 , n32622 );
and ( n32832 , n32829 , n32831 );
buf ( n32833 , n30889 );
buf ( n32834 , n15838 );
buf ( n32835 , n32834 );
and ( n32836 , n32833 , n32835 );
xor ( n32837 , n32606 , n32607 );
and ( n32838 , n32835 , n32837 );
and ( n32839 , n32833 , n32837 );
or ( n32840 , n32836 , n32838 , n32839 );
xor ( n32841 , n32603 , n32604 );
xor ( n32842 , n32841 , n32608 );
and ( n32843 , n32840 , n32842 );
xor ( n32844 , n32680 , n32698 );
and ( n32845 , n32842 , n32844 );
and ( n32846 , n32840 , n32844 );
or ( n32847 , n32843 , n32845 , n32846 );
xor ( n32848 , n32557 , n32558 );
xor ( n32849 , n32848 , n32560 );
xor ( n32850 , n32669 , n32672 );
xor ( n32851 , n32850 , n32674 );
or ( n32852 , n32849 , n32851 );
xor ( n32853 , n32572 , n32573 );
xor ( n32854 , n32853 , n32575 );
xor ( n32855 , n32687 , n32690 );
xor ( n32856 , n32855 , n32692 );
or ( n32857 , n32854 , n32856 );
and ( n32858 , n32852 , n32857 );
xnor ( n32859 , n32677 , n32679 );
xnor ( n32860 , n32695 , n32697 );
and ( n32861 , n32859 , n32860 );
and ( n32862 , n32858 , n32861 );
and ( n32863 , n31278 , n30791 );
and ( n32864 , n31088 , n30898 );
or ( n32865 , n32863 , n32864 );
and ( n32866 , n30799 , n31301 );
and ( n32867 , n30889 , n31073 );
or ( n32868 , n32866 , n32867 );
and ( n32869 , n32865 , n32868 );
xor ( n32870 , n32727 , n32744 );
and ( n32871 , n32869 , n32870 );
xor ( n32872 , n32760 , n32765 );
and ( n32873 , n32870 , n32872 );
and ( n32874 , n32869 , n32872 );
or ( n32875 , n32871 , n32873 , n32874 );
and ( n32876 , n32861 , n32875 );
and ( n32877 , n32858 , n32875 );
or ( n32878 , n32862 , n32876 , n32877 );
and ( n32879 , n32847 , n32878 );
xor ( n32880 , n32768 , n32770 );
xor ( n32881 , n32773 , n32774 );
and ( n32882 , n32880 , n32881 );
xnor ( n32883 , n32863 , n32864 );
xnor ( n32884 , n32866 , n32867 );
and ( n32885 , n32883 , n32884 );
buf ( n32886 , n15841 );
buf ( n32887 , n32886 );
or ( n32888 , n32885 , n32887 );
and ( n32889 , n32881 , n32888 );
and ( n32890 , n32880 , n32888 );
or ( n32891 , n32882 , n32889 , n32890 );
and ( n32892 , n30468 , n32173 );
and ( n32893 , n30503 , n32066 );
and ( n32894 , n32892 , n32893 );
and ( n32895 , n30803 , n31301 );
and ( n32896 , n32893 , n32895 );
and ( n32897 , n32892 , n32895 );
or ( n32898 , n32894 , n32896 , n32897 );
and ( n32899 , n30442 , n32671 );
and ( n32900 , n30464 , n32348 );
and ( n32901 , n32899 , n32900 );
and ( n32902 , n30799 , n31442 );
and ( n32903 , n32900 , n32902 );
and ( n32904 , n32899 , n32902 );
or ( n32905 , n32901 , n32903 , n32904 );
and ( n32906 , n32898 , n32905 );
and ( n32907 , n31736 , n30563 );
and ( n32908 , n32905 , n32907 );
and ( n32909 , n32898 , n32907 );
or ( n32910 , n32906 , n32908 , n32909 );
and ( n32911 , n32155 , n30473 );
and ( n32912 , n32057 , n30508 );
and ( n32913 , n32911 , n32912 );
and ( n32914 , n31278 , n30788 );
and ( n32915 , n32912 , n32914 );
and ( n32916 , n32911 , n32914 );
or ( n32917 , n32913 , n32915 , n32916 );
and ( n32918 , n32689 , n30439 );
and ( n32919 , n32365 , n30461 );
and ( n32920 , n32918 , n32919 );
and ( n32921 , n31464 , n30791 );
and ( n32922 , n32919 , n32921 );
and ( n32923 , n32918 , n32921 );
or ( n32924 , n32920 , n32922 , n32923 );
and ( n32925 , n32917 , n32924 );
and ( n32926 , n30558 , n31745 );
and ( n32927 , n32924 , n32926 );
and ( n32928 , n32917 , n32926 );
or ( n32929 , n32925 , n32927 , n32928 );
and ( n32930 , n32910 , n32929 );
buf ( n32931 , n1243 );
buf ( n32932 , n32931 );
and ( n32933 , n30413 , n32932 );
and ( n32934 , n30419 , n32719 );
and ( n32935 , n32933 , n32934 );
and ( n32936 , n30709 , n31590 );
and ( n32937 , n32934 , n32936 );
and ( n32938 , n32933 , n32936 );
or ( n32939 , n32935 , n32937 , n32938 );
and ( n32940 , n30558 , n31861 );
and ( n32941 , n30603 , n31745 );
and ( n32942 , n32940 , n32941 );
and ( n32943 , n30889 , n31247 );
and ( n32944 , n32941 , n32943 );
and ( n32945 , n32940 , n32943 );
or ( n32946 , n32942 , n32944 , n32945 );
or ( n32947 , n32939 , n32946 );
buf ( n32948 , n1243 );
buf ( n32949 , n32948 );
and ( n32950 , n32949 , n30421 );
and ( n32951 , n32736 , n30424 );
and ( n32952 , n32950 , n32951 );
and ( n32953 , n31607 , n30700 );
and ( n32954 , n32951 , n32953 );
and ( n32955 , n32950 , n32953 );
or ( n32956 , n32952 , n32954 , n32955 );
and ( n32957 , n31883 , n30563 );
and ( n32958 , n31736 , n30592 );
and ( n32959 , n32957 , n32958 );
and ( n32960 , n31238 , n30898 );
and ( n32961 , n32958 , n32960 );
and ( n32962 , n32957 , n32960 );
or ( n32963 , n32959 , n32961 , n32962 );
or ( n32964 , n32956 , n32963 );
and ( n32965 , n32947 , n32964 );
and ( n32966 , n32930 , n32965 );
xor ( n32967 , n32711 , n32712 );
xor ( n32968 , n32967 , n32714 );
xor ( n32969 , n32720 , n32721 );
xor ( n32970 , n32969 , n32723 );
and ( n32971 , n32968 , n32970 );
xor ( n32972 , n32728 , n32729 );
xor ( n32973 , n32972 , n32731 );
xor ( n32974 , n32737 , n32738 );
xor ( n32975 , n32974 , n32740 );
and ( n32976 , n32973 , n32975 );
and ( n32977 , n32971 , n32976 );
and ( n32978 , n32965 , n32977 );
and ( n32979 , n32930 , n32977 );
or ( n32980 , n32966 , n32978 , n32979 );
and ( n32981 , n32891 , n32980 );
xnor ( n32982 , n32717 , n32726 );
xnor ( n32983 , n32734 , n32743 );
and ( n32984 , n32982 , n32983 );
xnor ( n32985 , n32757 , n32759 );
xnor ( n32986 , n32762 , n32764 );
and ( n32987 , n32985 , n32986 );
and ( n32988 , n32984 , n32987 );
and ( n32989 , n31084 , n30898 );
and ( n32990 , n30889 , n31076 );
and ( n32991 , n32989 , n32990 );
xor ( n32992 , n32865 , n32868 );
and ( n32993 , n32990 , n32992 );
and ( n32994 , n32989 , n32992 );
or ( n32995 , n32991 , n32993 , n32994 );
and ( n32996 , n32987 , n32995 );
and ( n32997 , n32984 , n32995 );
or ( n32998 , n32988 , n32996 , n32997 );
and ( n32999 , n32980 , n32998 );
and ( n33000 , n32891 , n32998 );
or ( n33001 , n32981 , n32999 , n33000 );
and ( n33002 , n32878 , n33001 );
and ( n33003 , n32847 , n33001 );
or ( n33004 , n32879 , n33002 , n33003 );
and ( n33005 , n32831 , n33004 );
and ( n33006 , n32829 , n33004 );
or ( n33007 , n32832 , n33005 , n33006 );
and ( n33008 , n32826 , n33007 );
and ( n33009 , n32824 , n33007 );
or ( n33010 , n32827 , n33008 , n33009 );
xor ( n33011 , n32655 , n32805 );
xor ( n33012 , n33011 , n32808 );
and ( n33013 , n33010 , n33012 );
xor ( n33014 , n32700 , n32701 );
xor ( n33015 , n33014 , n32703 );
xor ( n33016 , n32708 , n32709 );
xor ( n33017 , n33016 , n32745 );
and ( n33018 , n33015 , n33017 );
xor ( n33019 , n32766 , n32771 );
xor ( n33020 , n33019 , n32775 );
and ( n33021 , n33017 , n33020 );
and ( n33022 , n33015 , n33020 );
or ( n33023 , n33018 , n33021 , n33022 );
xor ( n33024 , n32699 , n32706 );
xor ( n33025 , n33024 , n32748 );
and ( n33026 , n33023 , n33025 );
xor ( n33027 , n32778 , n32780 );
xor ( n33028 , n33027 , n32783 );
and ( n33029 , n33025 , n33028 );
and ( n33030 , n33023 , n33028 );
or ( n33031 , n33026 , n33029 , n33030 );
xor ( n33032 , n32659 , n32661 );
xor ( n33033 , n33032 , n32751 );
and ( n33034 , n33031 , n33033 );
xor ( n33035 , n32786 , n32796 );
xor ( n33036 , n33035 , n32799 );
and ( n33037 , n33033 , n33036 );
and ( n33038 , n33031 , n33036 );
or ( n33039 , n33034 , n33037 , n33038 );
xor ( n33040 , n32657 , n32754 );
xor ( n33041 , n33040 , n32802 );
and ( n33042 , n33039 , n33041 );
xor ( n33043 , n32788 , n32790 );
xor ( n33044 , n33043 , n32793 );
xor ( n33045 , n32833 , n32835 );
xor ( n33046 , n33045 , n32837 );
xor ( n33047 , n32852 , n32857 );
and ( n33048 , n33046 , n33047 );
xor ( n33049 , n32859 , n32860 );
and ( n33050 , n33047 , n33049 );
and ( n33051 , n33046 , n33049 );
or ( n33052 , n33048 , n33050 , n33051 );
xor ( n33053 , n32968 , n32970 );
xor ( n33054 , n32973 , n32975 );
and ( n33055 , n33053 , n33054 );
xnor ( n33056 , n32885 , n32887 );
and ( n33057 , n33055 , n33056 );
xor ( n33058 , n32892 , n32893 );
xor ( n33059 , n33058 , n32895 );
xor ( n33060 , n32940 , n32941 );
xor ( n33061 , n33060 , n32943 );
and ( n33062 , n33059 , n33061 );
xor ( n33063 , n32899 , n32900 );
xor ( n33064 , n33063 , n32902 );
and ( n33065 , n33061 , n33064 );
and ( n33066 , n33059 , n33064 );
or ( n33067 , n33062 , n33065 , n33066 );
xor ( n33068 , n32681 , n32682 );
xor ( n33069 , n33068 , n32684 );
or ( n33070 , n33067 , n33069 );
xor ( n33071 , n32911 , n32912 );
xor ( n33072 , n33071 , n32914 );
xor ( n33073 , n32957 , n32958 );
xor ( n33074 , n33073 , n32960 );
and ( n33075 , n33072 , n33074 );
xor ( n33076 , n32918 , n32919 );
xor ( n33077 , n33076 , n32921 );
and ( n33078 , n33074 , n33077 );
and ( n33079 , n33072 , n33077 );
or ( n33080 , n33075 , n33078 , n33079 );
xor ( n33081 , n32663 , n32664 );
xor ( n33082 , n33081 , n32666 );
or ( n33083 , n33080 , n33082 );
and ( n33084 , n33070 , n33083 );
and ( n33085 , n33057 , n33084 );
and ( n33086 , n32949 , n30424 );
and ( n33087 , n32736 , n30439 );
and ( n33088 , n33086 , n33087 );
and ( n33089 , n31736 , n30700 );
and ( n33090 , n33087 , n33089 );
and ( n33091 , n33086 , n33089 );
or ( n33092 , n33088 , n33090 , n33091 );
and ( n33093 , n32689 , n30461 );
and ( n33094 , n32365 , n30473 );
and ( n33095 , n33093 , n33094 );
and ( n33096 , n31278 , n30898 );
and ( n33097 , n33094 , n33096 );
and ( n33098 , n33093 , n33096 );
or ( n33099 , n33095 , n33097 , n33098 );
and ( n33100 , n33092 , n33099 );
xor ( n33101 , n32933 , n32934 );
xor ( n33102 , n33101 , n32936 );
and ( n33103 , n33099 , n33102 );
and ( n33104 , n33092 , n33102 );
or ( n33105 , n33100 , n33103 , n33104 );
xor ( n33106 , n32917 , n32924 );
xor ( n33107 , n33106 , n32926 );
and ( n33108 , n33105 , n33107 );
and ( n33109 , n30419 , n32932 );
and ( n33110 , n30442 , n32719 );
and ( n33111 , n33109 , n33110 );
and ( n33112 , n30709 , n31745 );
and ( n33113 , n33110 , n33112 );
and ( n33114 , n33109 , n33112 );
or ( n33115 , n33111 , n33113 , n33114 );
and ( n33116 , n30464 , n32671 );
and ( n33117 , n30468 , n32348 );
and ( n33118 , n33116 , n33117 );
and ( n33119 , n30889 , n31301 );
and ( n33120 , n33117 , n33119 );
and ( n33121 , n33116 , n33119 );
or ( n33122 , n33118 , n33120 , n33121 );
and ( n33123 , n33115 , n33122 );
xor ( n33124 , n32950 , n32951 );
xor ( n33125 , n33124 , n32953 );
and ( n33126 , n33122 , n33125 );
and ( n33127 , n33115 , n33125 );
or ( n33128 , n33123 , n33126 , n33127 );
xor ( n33129 , n32898 , n32905 );
xor ( n33130 , n33129 , n32907 );
and ( n33131 , n33128 , n33130 );
and ( n33132 , n33108 , n33131 );
and ( n33133 , n33084 , n33132 );
and ( n33134 , n33057 , n33132 );
or ( n33135 , n33085 , n33133 , n33134 );
and ( n33136 , n33052 , n33135 );
xnor ( n33137 , n32849 , n32851 );
xnor ( n33138 , n32854 , n32856 );
and ( n33139 , n33137 , n33138 );
buf ( n33140 , n31084 );
buf ( n33141 , n15844 );
buf ( n33142 , n33141 );
and ( n33143 , n33140 , n33142 );
and ( n33144 , n31088 , n31076 );
and ( n33145 , n31084 , n31073 );
and ( n33146 , n33144 , n33145 );
buf ( n33147 , n15847 );
buf ( n33148 , n33147 );
and ( n33149 , n33145 , n33148 );
and ( n33150 , n33144 , n33148 );
or ( n33151 , n33146 , n33149 , n33150 );
and ( n33152 , n33142 , n33151 );
and ( n33153 , n33140 , n33151 );
or ( n33154 , n33143 , n33152 , n33153 );
xor ( n33155 , n32910 , n32929 );
and ( n33156 , n33154 , n33155 );
xor ( n33157 , n32947 , n32964 );
and ( n33158 , n33155 , n33157 );
and ( n33159 , n33154 , n33157 );
or ( n33160 , n33156 , n33158 , n33159 );
and ( n33161 , n33139 , n33160 );
xor ( n33162 , n32971 , n32976 );
xor ( n33163 , n32982 , n32983 );
and ( n33164 , n33162 , n33163 );
xor ( n33165 , n32985 , n32986 );
and ( n33166 , n33163 , n33165 );
and ( n33167 , n33162 , n33165 );
or ( n33168 , n33164 , n33166 , n33167 );
and ( n33169 , n33160 , n33168 );
and ( n33170 , n33139 , n33168 );
or ( n33171 , n33161 , n33169 , n33170 );
and ( n33172 , n33135 , n33171 );
and ( n33173 , n33052 , n33171 );
or ( n33174 , n33136 , n33172 , n33173 );
and ( n33175 , n33044 , n33174 );
xnor ( n33176 , n32939 , n32946 );
xnor ( n33177 , n32956 , n32963 );
and ( n33178 , n33176 , n33177 );
xor ( n33179 , n32883 , n32884 );
and ( n33180 , n32155 , n30508 );
and ( n33181 , n32057 , n30563 );
and ( n33182 , n33180 , n33181 );
and ( n33183 , n31607 , n30791 );
and ( n33184 , n33181 , n33183 );
and ( n33185 , n33180 , n33183 );
or ( n33186 , n33182 , n33184 , n33185 );
and ( n33187 , n30503 , n32173 );
and ( n33188 , n30558 , n32066 );
and ( n33189 , n33187 , n33188 );
and ( n33190 , n30799 , n31590 );
and ( n33191 , n33188 , n33190 );
and ( n33192 , n33187 , n33190 );
or ( n33193 , n33189 , n33191 , n33192 );
and ( n33194 , n33186 , n33193 );
and ( n33195 , n33179 , n33194 );
and ( n33196 , n31464 , n30788 );
and ( n33197 , n31238 , n31076 );
or ( n33198 , n33196 , n33197 );
and ( n33199 , n30803 , n31442 );
and ( n33200 , n31084 , n31247 );
or ( n33201 , n33199 , n33200 );
and ( n33202 , n33198 , n33201 );
and ( n33203 , n33194 , n33202 );
and ( n33204 , n33179 , n33202 );
or ( n33205 , n33195 , n33203 , n33204 );
and ( n33206 , n33178 , n33205 );
xor ( n33207 , n32989 , n32990 );
xor ( n33208 , n33207 , n32992 );
and ( n33209 , n33205 , n33208 );
and ( n33210 , n33178 , n33208 );
or ( n33211 , n33206 , n33209 , n33210 );
xor ( n33212 , n32869 , n32870 );
xor ( n33213 , n33212 , n32872 );
and ( n33214 , n33211 , n33213 );
xor ( n33215 , n32880 , n32881 );
xor ( n33216 , n33215 , n32888 );
and ( n33217 , n33213 , n33216 );
and ( n33218 , n33211 , n33216 );
or ( n33219 , n33214 , n33217 , n33218 );
xor ( n33220 , n32840 , n32842 );
xor ( n33221 , n33220 , n32844 );
and ( n33222 , n33219 , n33221 );
xor ( n33223 , n32858 , n32861 );
xor ( n33224 , n33223 , n32875 );
and ( n33225 , n33221 , n33224 );
and ( n33226 , n33219 , n33224 );
or ( n33227 , n33222 , n33225 , n33226 );
and ( n33228 , n33174 , n33227 );
and ( n33229 , n33044 , n33227 );
or ( n33230 , n33175 , n33228 , n33229 );
xor ( n33231 , n32829 , n32831 );
xor ( n33232 , n33231 , n33004 );
and ( n33233 , n33230 , n33232 );
xor ( n33234 , n33031 , n33033 );
xor ( n33235 , n33234 , n33036 );
and ( n33236 , n33232 , n33235 );
and ( n33237 , n33230 , n33235 );
or ( n33238 , n33233 , n33236 , n33237 );
and ( n33239 , n33041 , n33238 );
and ( n33240 , n33039 , n33238 );
or ( n33241 , n33042 , n33239 , n33240 );
and ( n33242 , n33012 , n33241 );
and ( n33243 , n33010 , n33241 );
or ( n33244 , n33013 , n33242 , n33243 );
and ( n33245 , n32822 , n33244 );
xor ( n33246 , n33010 , n33012 );
xor ( n33247 , n33246 , n33241 );
xor ( n33248 , n32824 , n32826 );
xor ( n33249 , n33248 , n33007 );
xor ( n33250 , n33039 , n33041 );
xor ( n33251 , n33250 , n33238 );
and ( n33252 , n33249 , n33251 );
xor ( n33253 , n32847 , n32878 );
xor ( n33254 , n33253 , n33001 );
xor ( n33255 , n33023 , n33025 );
xor ( n33256 , n33255 , n33028 );
and ( n33257 , n33254 , n33256 );
xor ( n33258 , n32891 , n32980 );
xor ( n33259 , n33258 , n32998 );
xor ( n33260 , n33015 , n33017 );
xor ( n33261 , n33260 , n33020 );
and ( n33262 , n33259 , n33261 );
xor ( n33263 , n32930 , n32965 );
xor ( n33264 , n33263 , n32977 );
xor ( n33265 , n32984 , n32987 );
xor ( n33266 , n33265 , n32995 );
and ( n33267 , n33264 , n33266 );
xor ( n33268 , n33055 , n33056 );
xor ( n33269 , n33070 , n33083 );
and ( n33270 , n33268 , n33269 );
xor ( n33271 , n33108 , n33131 );
and ( n33272 , n33269 , n33271 );
and ( n33273 , n33268 , n33271 );
or ( n33274 , n33270 , n33272 , n33273 );
and ( n33275 , n33266 , n33274 );
and ( n33276 , n33264 , n33274 );
or ( n33277 , n33267 , n33275 , n33276 );
and ( n33278 , n33261 , n33277 );
and ( n33279 , n33259 , n33277 );
or ( n33280 , n33262 , n33278 , n33279 );
and ( n33281 , n33256 , n33280 );
and ( n33282 , n33254 , n33280 );
or ( n33283 , n33257 , n33281 , n33282 );
xor ( n33284 , n33230 , n33232 );
xor ( n33285 , n33284 , n33235 );
and ( n33286 , n33283 , n33285 );
xor ( n33287 , n33137 , n33138 );
and ( n33288 , n32949 , n30439 );
and ( n33289 , n32736 , n30461 );
and ( n33290 , n33288 , n33289 );
and ( n33291 , n31736 , n30791 );
and ( n33292 , n33289 , n33291 );
and ( n33293 , n33288 , n33291 );
or ( n33294 , n33290 , n33292 , n33293 );
buf ( n33295 , n1244 );
buf ( n33296 , n33295 );
and ( n33297 , n30413 , n33296 );
and ( n33298 , n33294 , n33297 );
and ( n33299 , n30603 , n31861 );
and ( n33300 , n33297 , n33299 );
and ( n33301 , n33294 , n33299 );
or ( n33302 , n33298 , n33300 , n33301 );
buf ( n33303 , n1245 );
buf ( n33304 , n33303 );
and ( n33305 , n33304 , n30421 );
and ( n33306 , n31883 , n30700 );
and ( n33307 , n33305 , n33306 );
and ( n33308 , n31278 , n31076 );
and ( n33309 , n33306 , n33308 );
and ( n33310 , n33305 , n33308 );
or ( n33311 , n33307 , n33309 , n33310 );
and ( n33312 , n32689 , n30473 );
and ( n33313 , n32365 , n30508 );
and ( n33314 , n33312 , n33313 );
and ( n33315 , n31607 , n30788 );
and ( n33316 , n33313 , n33315 );
and ( n33317 , n33312 , n33315 );
or ( n33318 , n33314 , n33316 , n33317 );
and ( n33319 , n33311 , n33318 );
and ( n33320 , n32155 , n30563 );
and ( n33321 , n32057 , n30592 );
and ( n33322 , n33320 , n33321 );
and ( n33323 , n31464 , n30898 );
and ( n33324 , n33321 , n33323 );
and ( n33325 , n33320 , n33323 );
or ( n33326 , n33322 , n33324 , n33325 );
and ( n33327 , n33318 , n33326 );
and ( n33328 , n33311 , n33326 );
or ( n33329 , n33319 , n33327 , n33328 );
or ( n33330 , n33302 , n33329 );
and ( n33331 , n30442 , n32932 );
and ( n33332 , n30464 , n32719 );
and ( n33333 , n33331 , n33332 );
and ( n33334 , n30799 , n31745 );
and ( n33335 , n33332 , n33334 );
and ( n33336 , n33331 , n33334 );
or ( n33337 , n33333 , n33335 , n33336 );
buf ( n33338 , n1244 );
buf ( n33339 , n33338 );
and ( n33340 , n33339 , n30421 );
and ( n33341 , n33337 , n33340 );
and ( n33342 , n31883 , n30592 );
and ( n33343 , n33340 , n33342 );
and ( n33344 , n33337 , n33342 );
or ( n33345 , n33341 , n33343 , n33344 );
buf ( n33346 , n1245 );
buf ( n33347 , n33346 );
and ( n33348 , n30413 , n33347 );
and ( n33349 , n30709 , n31861 );
and ( n33350 , n33348 , n33349 );
and ( n33351 , n31084 , n31301 );
and ( n33352 , n33349 , n33351 );
and ( n33353 , n33348 , n33351 );
or ( n33354 , n33350 , n33352 , n33353 );
and ( n33355 , n30468 , n32671 );
and ( n33356 , n30503 , n32348 );
and ( n33357 , n33355 , n33356 );
and ( n33358 , n30803 , n31590 );
and ( n33359 , n33356 , n33358 );
and ( n33360 , n33355 , n33358 );
or ( n33361 , n33357 , n33359 , n33360 );
and ( n33362 , n33354 , n33361 );
and ( n33363 , n30558 , n32173 );
and ( n33364 , n30603 , n32066 );
and ( n33365 , n33363 , n33364 );
and ( n33366 , n30889 , n31442 );
and ( n33367 , n33364 , n33366 );
and ( n33368 , n33363 , n33366 );
or ( n33369 , n33365 , n33367 , n33368 );
and ( n33370 , n33361 , n33369 );
and ( n33371 , n33354 , n33369 );
or ( n33372 , n33362 , n33370 , n33371 );
or ( n33373 , n33345 , n33372 );
and ( n33374 , n33330 , n33373 );
and ( n33375 , n33287 , n33374 );
xor ( n33376 , n33092 , n33099 );
xor ( n33377 , n33376 , n33102 );
xor ( n33378 , n33059 , n33061 );
xor ( n33379 , n33378 , n33064 );
or ( n33380 , n33377 , n33379 );
xor ( n33381 , n33115 , n33122 );
xor ( n33382 , n33381 , n33125 );
xor ( n33383 , n33072 , n33074 );
xor ( n33384 , n33383 , n33077 );
or ( n33385 , n33382 , n33384 );
and ( n33386 , n33380 , n33385 );
and ( n33387 , n33374 , n33386 );
and ( n33388 , n33287 , n33386 );
or ( n33389 , n33375 , n33387 , n33388 );
xnor ( n33390 , n33067 , n33069 );
xnor ( n33391 , n33080 , n33082 );
and ( n33392 , n33390 , n33391 );
xor ( n33393 , n33105 , n33107 );
xor ( n33394 , n33128 , n33130 );
and ( n33395 , n33393 , n33394 );
and ( n33396 , n33392 , n33395 );
xor ( n33397 , n33140 , n33142 );
xor ( n33398 , n33397 , n33151 );
xor ( n33399 , n33176 , n33177 );
and ( n33400 , n33398 , n33399 );
xor ( n33401 , n33053 , n33054 );
and ( n33402 , n33399 , n33401 );
and ( n33403 , n33398 , n33401 );
or ( n33404 , n33400 , n33402 , n33403 );
and ( n33405 , n33395 , n33404 );
and ( n33406 , n33392 , n33404 );
or ( n33407 , n33396 , n33405 , n33406 );
and ( n33408 , n33389 , n33407 );
xor ( n33409 , n33144 , n33145 );
xor ( n33410 , n33409 , n33148 );
xor ( n33411 , n33186 , n33193 );
and ( n33412 , n33410 , n33411 );
xor ( n33413 , n33198 , n33201 );
and ( n33414 , n33411 , n33413 );
and ( n33415 , n33410 , n33413 );
or ( n33416 , n33412 , n33414 , n33415 );
xor ( n33417 , n33180 , n33181 );
xor ( n33418 , n33417 , n33183 );
xor ( n33419 , n33187 , n33188 );
xor ( n33420 , n33419 , n33190 );
and ( n33421 , n33418 , n33420 );
xnor ( n33422 , n33196 , n33197 );
xnor ( n33423 , n33199 , n33200 );
and ( n33424 , n33422 , n33423 );
and ( n33425 , n33421 , n33424 );
buf ( n33426 , n31088 );
buf ( n33427 , n15850 );
buf ( n33428 , n33427 );
and ( n33429 , n33426 , n33428 );
and ( n33430 , n30419 , n33296 );
and ( n33431 , n33339 , n30424 );
and ( n33432 , n33430 , n33431 );
and ( n33433 , n33428 , n33432 );
and ( n33434 , n33426 , n33432 );
or ( n33435 , n33429 , n33433 , n33434 );
and ( n33436 , n33424 , n33435 );
and ( n33437 , n33421 , n33435 );
or ( n33438 , n33425 , n33436 , n33437 );
and ( n33439 , n33416 , n33438 );
xor ( n33440 , n33179 , n33194 );
xor ( n33441 , n33440 , n33202 );
and ( n33442 , n33438 , n33441 );
and ( n33443 , n33416 , n33441 );
or ( n33444 , n33439 , n33442 , n33443 );
xor ( n33445 , n33154 , n33155 );
xor ( n33446 , n33445 , n33157 );
and ( n33447 , n33444 , n33446 );
xor ( n33448 , n33162 , n33163 );
xor ( n33449 , n33448 , n33165 );
and ( n33450 , n33446 , n33449 );
and ( n33451 , n33444 , n33449 );
or ( n33452 , n33447 , n33450 , n33451 );
and ( n33453 , n33407 , n33452 );
and ( n33454 , n33389 , n33452 );
or ( n33455 , n33408 , n33453 , n33454 );
xor ( n33456 , n33046 , n33047 );
xor ( n33457 , n33456 , n33049 );
xor ( n33458 , n33057 , n33084 );
xor ( n33459 , n33458 , n33132 );
and ( n33460 , n33457 , n33459 );
xor ( n33461 , n33139 , n33160 );
xor ( n33462 , n33461 , n33168 );
and ( n33463 , n33459 , n33462 );
and ( n33464 , n33457 , n33462 );
or ( n33465 , n33460 , n33463 , n33464 );
and ( n33466 , n33455 , n33465 );
xor ( n33467 , n33052 , n33135 );
xor ( n33468 , n33467 , n33171 );
and ( n33469 , n33465 , n33468 );
and ( n33470 , n33455 , n33468 );
or ( n33471 , n33466 , n33469 , n33470 );
xor ( n33472 , n33044 , n33174 );
xor ( n33473 , n33472 , n33227 );
and ( n33474 , n33471 , n33473 );
xor ( n33475 , n33219 , n33221 );
xor ( n33476 , n33475 , n33224 );
xor ( n33477 , n33211 , n33213 );
xor ( n33478 , n33477 , n33216 );
xor ( n33479 , n33178 , n33205 );
xor ( n33480 , n33479 , n33208 );
xor ( n33481 , n33330 , n33373 );
xor ( n33482 , n33380 , n33385 );
and ( n33483 , n33481 , n33482 );
xor ( n33484 , n33390 , n33391 );
and ( n33485 , n33482 , n33484 );
and ( n33486 , n33481 , n33484 );
or ( n33487 , n33483 , n33485 , n33486 );
and ( n33488 , n33480 , n33487 );
xor ( n33489 , n33393 , n33394 );
xor ( n33490 , n33086 , n33087 );
xor ( n33491 , n33490 , n33089 );
xor ( n33492 , n33093 , n33094 );
xor ( n33493 , n33492 , n33096 );
and ( n33494 , n33491 , n33493 );
xor ( n33495 , n33337 , n33340 );
xor ( n33496 , n33495 , n33342 );
and ( n33497 , n33493 , n33496 );
and ( n33498 , n33491 , n33496 );
or ( n33499 , n33494 , n33497 , n33498 );
xor ( n33500 , n33109 , n33110 );
xor ( n33501 , n33500 , n33112 );
xor ( n33502 , n33116 , n33117 );
xor ( n33503 , n33502 , n33119 );
and ( n33504 , n33501 , n33503 );
xor ( n33505 , n33294 , n33297 );
xor ( n33506 , n33505 , n33299 );
and ( n33507 , n33503 , n33506 );
and ( n33508 , n33501 , n33506 );
or ( n33509 , n33504 , n33507 , n33508 );
and ( n33510 , n33499 , n33509 );
and ( n33511 , n33489 , n33510 );
and ( n33512 , n33339 , n30439 );
and ( n33513 , n32949 , n30461 );
and ( n33514 , n33512 , n33513 );
and ( n33515 , n31883 , n30791 );
and ( n33516 , n33513 , n33515 );
and ( n33517 , n33512 , n33515 );
or ( n33518 , n33514 , n33516 , n33517 );
and ( n33519 , n32736 , n30473 );
and ( n33520 , n32689 , n30508 );
and ( n33521 , n33519 , n33520 );
and ( n33522 , n31464 , n31076 );
and ( n33523 , n33520 , n33522 );
and ( n33524 , n33519 , n33522 );
or ( n33525 , n33521 , n33523 , n33524 );
and ( n33526 , n33518 , n33525 );
and ( n33527 , n32365 , n30563 );
and ( n33528 , n32155 , n30592 );
and ( n33529 , n33527 , n33528 );
and ( n33530 , n31736 , n30788 );
and ( n33531 , n33528 , n33530 );
and ( n33532 , n33527 , n33530 );
or ( n33533 , n33529 , n33531 , n33532 );
and ( n33534 , n33525 , n33533 );
and ( n33535 , n33518 , n33533 );
or ( n33536 , n33526 , n33534 , n33535 );
xor ( n33537 , n33311 , n33318 );
xor ( n33538 , n33537 , n33326 );
or ( n33539 , n33536 , n33538 );
and ( n33540 , n30442 , n33296 );
and ( n33541 , n30464 , n32932 );
and ( n33542 , n33540 , n33541 );
and ( n33543 , n30799 , n31861 );
and ( n33544 , n33541 , n33543 );
and ( n33545 , n33540 , n33543 );
or ( n33546 , n33542 , n33544 , n33545 );
and ( n33547 , n30468 , n32719 );
and ( n33548 , n30503 , n32671 );
and ( n33549 , n33547 , n33548 );
and ( n33550 , n31084 , n31442 );
and ( n33551 , n33548 , n33550 );
and ( n33552 , n33547 , n33550 );
or ( n33553 , n33549 , n33551 , n33552 );
and ( n33554 , n33546 , n33553 );
and ( n33555 , n30558 , n32348 );
and ( n33556 , n30603 , n32173 );
and ( n33557 , n33555 , n33556 );
and ( n33558 , n30803 , n31745 );
and ( n33559 , n33556 , n33558 );
and ( n33560 , n33555 , n33558 );
or ( n33561 , n33557 , n33559 , n33560 );
and ( n33562 , n33553 , n33561 );
and ( n33563 , n33546 , n33561 );
or ( n33564 , n33554 , n33562 , n33563 );
xor ( n33565 , n33354 , n33361 );
xor ( n33566 , n33565 , n33369 );
or ( n33567 , n33564 , n33566 );
and ( n33568 , n33539 , n33567 );
and ( n33569 , n33510 , n33568 );
and ( n33570 , n33489 , n33568 );
or ( n33571 , n33511 , n33569 , n33570 );
and ( n33572 , n33487 , n33571 );
and ( n33573 , n33480 , n33571 );
or ( n33574 , n33488 , n33572 , n33573 );
and ( n33575 , n33478 , n33574 );
xnor ( n33576 , n33302 , n33329 );
xnor ( n33577 , n33345 , n33372 );
and ( n33578 , n33576 , n33577 );
xnor ( n33579 , n33377 , n33379 );
xnor ( n33580 , n33382 , n33384 );
and ( n33581 , n33579 , n33580 );
and ( n33582 , n33578 , n33581 );
xor ( n33583 , n33355 , n33356 );
xor ( n33584 , n33583 , n33358 );
xor ( n33585 , n33363 , n33364 );
xor ( n33586 , n33585 , n33366 );
or ( n33587 , n33584 , n33586 );
xor ( n33588 , n33312 , n33313 );
xor ( n33589 , n33588 , n33315 );
xor ( n33590 , n33320 , n33321 );
xor ( n33591 , n33590 , n33323 );
or ( n33592 , n33589 , n33591 );
and ( n33593 , n33587 , n33592 );
and ( n33594 , n31238 , n31073 );
and ( n33595 , n31088 , n31247 );
and ( n33596 , n33594 , n33595 );
buf ( n33597 , n15853 );
buf ( n33598 , n33597 );
and ( n33599 , n33595 , n33598 );
and ( n33600 , n33594 , n33598 );
or ( n33601 , n33596 , n33599 , n33600 );
xor ( n33602 , n33418 , n33420 );
and ( n33603 , n33601 , n33602 );
xor ( n33604 , n33422 , n33423 );
and ( n33605 , n33602 , n33604 );
and ( n33606 , n33601 , n33604 );
or ( n33607 , n33603 , n33605 , n33606 );
and ( n33608 , n33593 , n33607 );
xor ( n33609 , n33410 , n33411 );
xor ( n33610 , n33609 , n33413 );
and ( n33611 , n33607 , n33610 );
and ( n33612 , n33593 , n33610 );
or ( n33613 , n33608 , n33611 , n33612 );
and ( n33614 , n33581 , n33613 );
and ( n33615 , n33578 , n33613 );
or ( n33616 , n33582 , n33614 , n33615 );
xor ( n33617 , n33268 , n33269 );
xor ( n33618 , n33617 , n33271 );
and ( n33619 , n33616 , n33618 );
xor ( n33620 , n33287 , n33374 );
xor ( n33621 , n33620 , n33386 );
and ( n33622 , n33618 , n33621 );
and ( n33623 , n33616 , n33621 );
or ( n33624 , n33619 , n33622 , n33623 );
and ( n33625 , n33574 , n33624 );
and ( n33626 , n33478 , n33624 );
or ( n33627 , n33575 , n33625 , n33626 );
and ( n33628 , n33476 , n33627 );
xor ( n33629 , n33264 , n33266 );
xor ( n33630 , n33629 , n33274 );
xor ( n33631 , n33389 , n33407 );
xor ( n33632 , n33631 , n33452 );
and ( n33633 , n33630 , n33632 );
xor ( n33634 , n33457 , n33459 );
xor ( n33635 , n33634 , n33462 );
and ( n33636 , n33632 , n33635 );
and ( n33637 , n33630 , n33635 );
or ( n33638 , n33633 , n33636 , n33637 );
and ( n33639 , n33627 , n33638 );
and ( n33640 , n33476 , n33638 );
or ( n33641 , n33628 , n33639 , n33640 );
and ( n33642 , n33473 , n33641 );
and ( n33643 , n33471 , n33641 );
or ( n33644 , n33474 , n33642 , n33643 );
and ( n33645 , n33285 , n33644 );
and ( n33646 , n33283 , n33644 );
or ( n33647 , n33286 , n33645 , n33646 );
and ( n33648 , n33251 , n33647 );
and ( n33649 , n33249 , n33647 );
or ( n33650 , n33252 , n33648 , n33649 );
or ( n33651 , n33247 , n33650 );
and ( n33652 , n33244 , n33651 );
and ( n33653 , n32822 , n33651 );
or ( n33654 , n33245 , n33652 , n33653 );
and ( n33655 , n32819 , n33654 );
and ( n33656 , n32817 , n33654 );
or ( n33657 , n32820 , n33655 , n33656 );
and ( n33658 , n32650 , n33657 );
and ( n33659 , n32648 , n33657 );
or ( n33660 , n32651 , n33658 , n33659 );
and ( n33661 , n32473 , n33660 );
xor ( n33662 , n32473 , n33660 );
xor ( n33663 , n32648 , n32650 );
xor ( n33664 , n33663 , n33657 );
not ( n33665 , n33664 );
xor ( n33666 , n32817 , n32819 );
xor ( n33667 , n33666 , n33654 );
not ( n33668 , n33667 );
xor ( n33669 , n32822 , n33244 );
xor ( n33670 , n33669 , n33651 );
xnor ( n33671 , n33247 , n33650 );
xor ( n33672 , n33249 , n33251 );
xor ( n33673 , n33672 , n33647 );
xor ( n33674 , n33254 , n33256 );
xor ( n33675 , n33674 , n33280 );
xor ( n33676 , n33259 , n33261 );
xor ( n33677 , n33676 , n33277 );
xor ( n33678 , n33455 , n33465 );
xor ( n33679 , n33678 , n33468 );
and ( n33680 , n33677 , n33679 );
xor ( n33681 , n33392 , n33395 );
xor ( n33682 , n33681 , n33404 );
xor ( n33683 , n33444 , n33446 );
xor ( n33684 , n33683 , n33449 );
and ( n33685 , n33682 , n33684 );
xor ( n33686 , n33398 , n33399 );
xor ( n33687 , n33686 , n33401 );
xor ( n33688 , n33416 , n33438 );
xor ( n33689 , n33688 , n33441 );
and ( n33690 , n33687 , n33689 );
buf ( n33691 , n1246 );
buf ( n33692 , n33691 );
and ( n33693 , n33692 , n30421 );
and ( n33694 , n33304 , n30424 );
and ( n33695 , n33693 , n33694 );
and ( n33696 , n32057 , n30700 );
and ( n33697 , n33694 , n33696 );
and ( n33698 , n33693 , n33696 );
or ( n33699 , n33695 , n33697 , n33698 );
xor ( n33700 , n33348 , n33349 );
xor ( n33701 , n33700 , n33351 );
and ( n33702 , n33699 , n33701 );
xor ( n33703 , n33331 , n33332 );
xor ( n33704 , n33703 , n33334 );
and ( n33705 , n33701 , n33704 );
and ( n33706 , n33699 , n33704 );
or ( n33707 , n33702 , n33705 , n33706 );
xor ( n33708 , n33501 , n33503 );
xor ( n33709 , n33708 , n33506 );
or ( n33710 , n33707 , n33709 );
buf ( n33711 , n1246 );
buf ( n33712 , n33711 );
and ( n33713 , n30413 , n33712 );
and ( n33714 , n30419 , n33347 );
and ( n33715 , n33713 , n33714 );
and ( n33716 , n30709 , n32066 );
and ( n33717 , n33714 , n33716 );
and ( n33718 , n33713 , n33716 );
or ( n33719 , n33715 , n33717 , n33718 );
xor ( n33720 , n33305 , n33306 );
xor ( n33721 , n33720 , n33308 );
and ( n33722 , n33719 , n33721 );
xor ( n33723 , n33288 , n33289 );
xor ( n33724 , n33723 , n33291 );
and ( n33725 , n33721 , n33724 );
and ( n33726 , n33719 , n33724 );
or ( n33727 , n33722 , n33725 , n33726 );
xor ( n33728 , n33491 , n33493 );
xor ( n33729 , n33728 , n33496 );
or ( n33730 , n33727 , n33729 );
and ( n33731 , n33710 , n33730 );
and ( n33732 , n33689 , n33731 );
and ( n33733 , n33687 , n33731 );
or ( n33734 , n33690 , n33732 , n33733 );
and ( n33735 , n33684 , n33734 );
and ( n33736 , n33682 , n33734 );
or ( n33737 , n33685 , n33735 , n33736 );
xor ( n33738 , n33421 , n33424 );
xor ( n33739 , n33738 , n33435 );
xor ( n33740 , n33499 , n33509 );
and ( n33741 , n33739 , n33740 );
xor ( n33742 , n33539 , n33567 );
and ( n33743 , n33740 , n33742 );
and ( n33744 , n33739 , n33742 );
or ( n33745 , n33741 , n33743 , n33744 );
xor ( n33746 , n33576 , n33577 );
xor ( n33747 , n33579 , n33580 );
and ( n33748 , n33746 , n33747 );
and ( n33749 , n32949 , n30473 );
and ( n33750 , n32736 , n30508 );
and ( n33751 , n33749 , n33750 );
and ( n33752 , n31883 , n30788 );
and ( n33753 , n33750 , n33752 );
and ( n33754 , n33749 , n33752 );
or ( n33755 , n33751 , n33753 , n33754 );
and ( n33756 , n32689 , n30563 );
and ( n33757 , n32365 , n30592 );
and ( n33758 , n33756 , n33757 );
and ( n33759 , n31736 , n30898 );
and ( n33760 , n33757 , n33759 );
and ( n33761 , n33756 , n33759 );
or ( n33762 , n33758 , n33760 , n33761 );
and ( n33763 , n33755 , n33762 );
xor ( n33764 , n33555 , n33556 );
xor ( n33765 , n33764 , n33558 );
and ( n33766 , n33762 , n33765 );
and ( n33767 , n33755 , n33765 );
or ( n33768 , n33763 , n33766 , n33767 );
xor ( n33769 , n33699 , n33701 );
xor ( n33770 , n33769 , n33704 );
or ( n33771 , n33768 , n33770 );
and ( n33772 , n30468 , n32932 );
and ( n33773 , n30503 , n32719 );
and ( n33774 , n33772 , n33773 );
and ( n33775 , n30803 , n31861 );
and ( n33776 , n33773 , n33775 );
and ( n33777 , n33772 , n33775 );
or ( n33778 , n33774 , n33776 , n33777 );
and ( n33779 , n30558 , n32671 );
and ( n33780 , n30603 , n32348 );
and ( n33781 , n33779 , n33780 );
and ( n33782 , n30889 , n31745 );
and ( n33783 , n33780 , n33782 );
and ( n33784 , n33779 , n33782 );
or ( n33785 , n33781 , n33783 , n33784 );
and ( n33786 , n33778 , n33785 );
xor ( n33787 , n33527 , n33528 );
xor ( n33788 , n33787 , n33530 );
and ( n33789 , n33785 , n33788 );
and ( n33790 , n33778 , n33788 );
or ( n33791 , n33786 , n33789 , n33790 );
xor ( n33792 , n33719 , n33721 );
xor ( n33793 , n33792 , n33724 );
or ( n33794 , n33791 , n33793 );
and ( n33795 , n33771 , n33794 );
and ( n33796 , n33747 , n33795 );
and ( n33797 , n33746 , n33795 );
or ( n33798 , n33748 , n33796 , n33797 );
and ( n33799 , n33745 , n33798 );
xnor ( n33800 , n33536 , n33538 );
xnor ( n33801 , n33564 , n33566 );
and ( n33802 , n33800 , n33801 );
and ( n33803 , n31607 , n30898 );
and ( n33804 , n31278 , n31073 );
or ( n33805 , n33803 , n33804 );
and ( n33806 , n30889 , n31590 );
and ( n33807 , n31088 , n31301 );
or ( n33808 , n33806 , n33807 );
and ( n33809 , n33805 , n33808 );
xor ( n33810 , n33426 , n33428 );
xor ( n33811 , n33810 , n33432 );
and ( n33812 , n33809 , n33811 );
xor ( n33813 , n33587 , n33592 );
and ( n33814 , n33811 , n33813 );
and ( n33815 , n33809 , n33813 );
or ( n33816 , n33812 , n33814 , n33815 );
and ( n33817 , n33802 , n33816 );
xor ( n33818 , n33713 , n33714 );
xor ( n33819 , n33818 , n33716 );
xor ( n33820 , n33540 , n33541 );
xor ( n33821 , n33820 , n33543 );
or ( n33822 , n33819 , n33821 );
xor ( n33823 , n33693 , n33694 );
xor ( n33824 , n33823 , n33696 );
xor ( n33825 , n33512 , n33513 );
xor ( n33826 , n33825 , n33515 );
or ( n33827 , n33824 , n33826 );
and ( n33828 , n33822 , n33827 );
xor ( n33829 , n33546 , n33553 );
xor ( n33830 , n33829 , n33561 );
xor ( n33831 , n33518 , n33525 );
xor ( n33832 , n33831 , n33533 );
and ( n33833 , n33830 , n33832 );
and ( n33834 , n33828 , n33833 );
xnor ( n33835 , n33584 , n33586 );
xnor ( n33836 , n33589 , n33591 );
and ( n33837 , n33835 , n33836 );
and ( n33838 , n33833 , n33837 );
and ( n33839 , n33828 , n33837 );
or ( n33840 , n33834 , n33838 , n33839 );
and ( n33841 , n33816 , n33840 );
and ( n33842 , n33802 , n33840 );
or ( n33843 , n33817 , n33841 , n33842 );
and ( n33844 , n33798 , n33843 );
and ( n33845 , n33745 , n33843 );
or ( n33846 , n33799 , n33844 , n33845 );
xor ( n33847 , n33481 , n33482 );
xor ( n33848 , n33847 , n33484 );
xor ( n33849 , n33489 , n33510 );
xor ( n33850 , n33849 , n33568 );
and ( n33851 , n33848 , n33850 );
xor ( n33852 , n33578 , n33581 );
xor ( n33853 , n33852 , n33613 );
and ( n33854 , n33850 , n33853 );
and ( n33855 , n33848 , n33853 );
or ( n33856 , n33851 , n33854 , n33855 );
and ( n33857 , n33846 , n33856 );
xor ( n33858 , n33480 , n33487 );
xor ( n33859 , n33858 , n33571 );
and ( n33860 , n33856 , n33859 );
and ( n33861 , n33846 , n33859 );
or ( n33862 , n33857 , n33860 , n33861 );
and ( n33863 , n33737 , n33862 );
xor ( n33864 , n33478 , n33574 );
xor ( n33865 , n33864 , n33624 );
and ( n33866 , n33862 , n33865 );
and ( n33867 , n33737 , n33865 );
or ( n33868 , n33863 , n33866 , n33867 );
and ( n33869 , n33679 , n33868 );
and ( n33870 , n33677 , n33868 );
or ( n33871 , n33680 , n33869 , n33870 );
and ( n33872 , n33675 , n33871 );
xor ( n33873 , n33471 , n33473 );
xor ( n33874 , n33873 , n33641 );
and ( n33875 , n33871 , n33874 );
and ( n33876 , n33675 , n33874 );
or ( n33877 , n33872 , n33875 , n33876 );
xor ( n33878 , n33283 , n33285 );
xor ( n33879 , n33878 , n33644 );
and ( n33880 , n33877 , n33879 );
xor ( n33881 , n33476 , n33627 );
xor ( n33882 , n33881 , n33638 );
xor ( n33883 , n33630 , n33632 );
xor ( n33884 , n33883 , n33635 );
xor ( n33885 , n33616 , n33618 );
xor ( n33886 , n33885 , n33621 );
xor ( n33887 , n33430 , n33431 );
xor ( n33888 , n33594 , n33595 );
xor ( n33889 , n33888 , n33598 );
and ( n33890 , n33887 , n33889 );
xor ( n33891 , n33805 , n33808 );
and ( n33892 , n33889 , n33891 );
and ( n33893 , n33887 , n33891 );
or ( n33894 , n33890 , n33892 , n33893 );
buf ( n33895 , n1247 );
buf ( n33896 , n33895 );
and ( n33897 , n33896 , n30421 );
and ( n33898 , n32155 , n30700 );
and ( n33899 , n33897 , n33898 );
and ( n33900 , n31607 , n31076 );
and ( n33901 , n33898 , n33900 );
and ( n33902 , n33897 , n33900 );
or ( n33903 , n33899 , n33901 , n33902 );
buf ( n33904 , n1247 );
buf ( n33905 , n33904 );
and ( n33906 , n30413 , n33905 );
and ( n33907 , n30709 , n32173 );
and ( n33908 , n33906 , n33907 );
and ( n33909 , n31084 , n31590 );
and ( n33910 , n33907 , n33909 );
and ( n33911 , n33906 , n33909 );
or ( n33912 , n33908 , n33910 , n33911 );
and ( n33913 , n33903 , n33912 );
and ( n33914 , n33692 , n30424 );
and ( n33915 , n32057 , n30791 );
and ( n33916 , n33914 , n33915 );
and ( n33917 , n31464 , n31073 );
and ( n33918 , n33915 , n33917 );
and ( n33919 , n33914 , n33917 );
or ( n33920 , n33916 , n33918 , n33919 );
and ( n33921 , n30419 , n33712 );
and ( n33922 , n30799 , n32066 );
and ( n33923 , n33921 , n33922 );
and ( n33924 , n31088 , n31442 );
and ( n33925 , n33922 , n33924 );
and ( n33926 , n33921 , n33924 );
or ( n33927 , n33923 , n33925 , n33926 );
and ( n33928 , n33920 , n33927 );
and ( n33929 , n33913 , n33928 );
and ( n33930 , n33304 , n30439 );
and ( n33931 , n33339 , n30461 );
or ( n33932 , n33930 , n33931 );
and ( n33933 , n30442 , n33347 );
and ( n33934 , n30464 , n33296 );
or ( n33935 , n33933 , n33934 );
and ( n33936 , n33932 , n33935 );
and ( n33937 , n33928 , n33936 );
and ( n33938 , n33913 , n33936 );
or ( n33939 , n33929 , n33937 , n33938 );
and ( n33940 , n33894 , n33939 );
xor ( n33941 , n33519 , n33520 );
xor ( n33942 , n33941 , n33522 );
xor ( n33943 , n33547 , n33548 );
xor ( n33944 , n33943 , n33550 );
and ( n33945 , n33942 , n33944 );
xnor ( n33946 , n33803 , n33804 );
xnor ( n33947 , n33806 , n33807 );
and ( n33948 , n33946 , n33947 );
and ( n33949 , n33945 , n33948 );
buf ( n33950 , n31238 );
buf ( n33951 , n15856 );
buf ( n33952 , n33951 );
and ( n33953 , n33950 , n33952 );
and ( n33954 , n31278 , n31247 );
and ( n33955 , n31238 , n31301 );
and ( n33956 , n33954 , n33955 );
buf ( n33957 , n15859 );
buf ( n33958 , n33957 );
and ( n33959 , n33955 , n33958 );
and ( n33960 , n33954 , n33958 );
or ( n33961 , n33956 , n33959 , n33960 );
and ( n33962 , n33952 , n33961 );
and ( n33963 , n33950 , n33961 );
or ( n33964 , n33953 , n33962 , n33963 );
and ( n33965 , n33948 , n33964 );
and ( n33966 , n33945 , n33964 );
or ( n33967 , n33949 , n33965 , n33966 );
and ( n33968 , n33939 , n33967 );
and ( n33969 , n33894 , n33967 );
or ( n33970 , n33940 , n33968 , n33969 );
xor ( n33971 , n33593 , n33607 );
xor ( n33972 , n33971 , n33610 );
and ( n33973 , n33970 , n33972 );
xor ( n33974 , n33710 , n33730 );
and ( n33975 , n33972 , n33974 );
and ( n33976 , n33970 , n33974 );
or ( n33977 , n33973 , n33975 , n33976 );
xnor ( n33978 , n33707 , n33709 );
xnor ( n33979 , n33727 , n33729 );
and ( n33980 , n33978 , n33979 );
xor ( n33981 , n33601 , n33602 );
xor ( n33982 , n33981 , n33604 );
xor ( n33983 , n33771 , n33794 );
and ( n33984 , n33982 , n33983 );
xor ( n33985 , n33800 , n33801 );
and ( n33986 , n33983 , n33985 );
and ( n33987 , n33982 , n33985 );
or ( n33988 , n33984 , n33986 , n33987 );
and ( n33989 , n33980 , n33988 );
and ( n33990 , n33339 , n30473 );
and ( n33991 , n32057 , n30788 );
and ( n33992 , n33990 , n33991 );
and ( n33993 , n31607 , n31073 );
and ( n33994 , n33991 , n33993 );
and ( n33995 , n33990 , n33993 );
or ( n33996 , n33992 , n33994 , n33995 );
and ( n33997 , n33692 , n30439 );
and ( n33998 , n33304 , n30461 );
and ( n33999 , n33997 , n33998 );
and ( n34000 , n32155 , n30791 );
and ( n34001 , n33998 , n34000 );
and ( n34002 , n33997 , n34000 );
or ( n34003 , n33999 , n34001 , n34002 );
and ( n34004 , n33996 , n34003 );
xor ( n34005 , n33921 , n33922 );
xor ( n34006 , n34005 , n33924 );
and ( n34007 , n34003 , n34006 );
and ( n34008 , n33996 , n34006 );
or ( n34009 , n34004 , n34007 , n34008 );
not ( n34010 , n34009 );
xor ( n34011 , n33755 , n33762 );
xor ( n34012 , n34011 , n33765 );
and ( n34013 , n34010 , n34012 );
and ( n34014 , n30468 , n33296 );
and ( n34015 , n30803 , n32066 );
and ( n34016 , n34014 , n34015 );
and ( n34017 , n31088 , n31590 );
and ( n34018 , n34015 , n34017 );
and ( n34019 , n34014 , n34017 );
or ( n34020 , n34016 , n34018 , n34019 );
and ( n34021 , n30442 , n33712 );
and ( n34022 , n30464 , n33347 );
and ( n34023 , n34021 , n34022 );
and ( n34024 , n30799 , n32173 );
and ( n34025 , n34022 , n34024 );
and ( n34026 , n34021 , n34024 );
or ( n34027 , n34023 , n34025 , n34026 );
and ( n34028 , n34020 , n34027 );
xor ( n34029 , n33914 , n33915 );
xor ( n34030 , n34029 , n33917 );
and ( n34031 , n34027 , n34030 );
and ( n34032 , n34020 , n34030 );
or ( n34033 , n34028 , n34031 , n34032 );
not ( n34034 , n34033 );
xor ( n34035 , n33778 , n33785 );
xor ( n34036 , n34035 , n33788 );
and ( n34037 , n34034 , n34036 );
and ( n34038 , n34013 , n34037 );
buf ( n34039 , n34009 );
buf ( n34040 , n34033 );
and ( n34041 , n34039 , n34040 );
and ( n34042 , n34038 , n34041 );
xnor ( n34043 , n33768 , n33770 );
xnor ( n34044 , n33791 , n33793 );
and ( n34045 , n34043 , n34044 );
and ( n34046 , n34041 , n34045 );
and ( n34047 , n34038 , n34045 );
or ( n34048 , n34042 , n34046 , n34047 );
and ( n34049 , n33988 , n34048 );
and ( n34050 , n33980 , n34048 );
or ( n34051 , n33989 , n34049 , n34050 );
and ( n34052 , n33977 , n34051 );
xor ( n34053 , n33822 , n33827 );
xor ( n34054 , n33830 , n33832 );
and ( n34055 , n34053 , n34054 );
xor ( n34056 , n33835 , n33836 );
and ( n34057 , n34054 , n34056 );
and ( n34058 , n34053 , n34056 );
or ( n34059 , n34055 , n34057 , n34058 );
xor ( n34060 , n33749 , n33750 );
xor ( n34061 , n34060 , n33752 );
xor ( n34062 , n33756 , n33757 );
xor ( n34063 , n34062 , n33759 );
and ( n34064 , n34061 , n34063 );
xor ( n34065 , n33897 , n33898 );
xor ( n34066 , n34065 , n33900 );
and ( n34067 , n34063 , n34066 );
and ( n34068 , n34061 , n34066 );
or ( n34069 , n34064 , n34067 , n34068 );
xor ( n34070 , n33772 , n33773 );
xor ( n34071 , n34070 , n33775 );
xor ( n34072 , n33779 , n33780 );
xor ( n34073 , n34072 , n33782 );
and ( n34074 , n34071 , n34073 );
xor ( n34075 , n33906 , n33907 );
xor ( n34076 , n34075 , n33909 );
and ( n34077 , n34073 , n34076 );
and ( n34078 , n34071 , n34076 );
or ( n34079 , n34074 , n34077 , n34078 );
and ( n34080 , n34069 , n34079 );
buf ( n34081 , n1248 );
buf ( n34082 , n34081 );
and ( n34083 , n30413 , n34082 );
and ( n34084 , n30603 , n32671 );
and ( n34085 , n34083 , n34084 );
and ( n34086 , n30709 , n32348 );
and ( n34087 , n34084 , n34086 );
and ( n34088 , n34083 , n34086 );
or ( n34089 , n34085 , n34087 , n34088 );
and ( n34090 , n30503 , n32932 );
and ( n34091 , n30558 , n32719 );
and ( n34092 , n34090 , n34091 );
and ( n34093 , n30889 , n31861 );
and ( n34094 , n34091 , n34093 );
and ( n34095 , n34090 , n34093 );
or ( n34096 , n34092 , n34094 , n34095 );
or ( n34097 , n34089 , n34096 );
buf ( n34098 , n1248 );
buf ( n34099 , n34098 );
and ( n34100 , n34099 , n30421 );
and ( n34101 , n32689 , n30592 );
and ( n34102 , n34100 , n34101 );
and ( n34103 , n32365 , n30700 );
and ( n34104 , n34101 , n34103 );
and ( n34105 , n34100 , n34103 );
or ( n34106 , n34102 , n34104 , n34105 );
and ( n34107 , n32949 , n30508 );
and ( n34108 , n32736 , n30563 );
and ( n34109 , n34107 , n34108 );
and ( n34110 , n31883 , n30898 );
and ( n34111 , n34108 , n34110 );
and ( n34112 , n34107 , n34110 );
or ( n34113 , n34109 , n34111 , n34112 );
or ( n34114 , n34106 , n34113 );
and ( n34115 , n34097 , n34114 );
and ( n34116 , n34080 , n34115 );
xnor ( n34117 , n33819 , n33821 );
xnor ( n34118 , n33824 , n33826 );
and ( n34119 , n34117 , n34118 );
and ( n34120 , n34115 , n34119 );
and ( n34121 , n34080 , n34119 );
or ( n34122 , n34116 , n34120 , n34121 );
and ( n34123 , n34059 , n34122 );
xor ( n34124 , n33903 , n33912 );
xor ( n34125 , n33920 , n33927 );
and ( n34126 , n34124 , n34125 );
xor ( n34127 , n33932 , n33935 );
and ( n34128 , n34125 , n34127 );
and ( n34129 , n34124 , n34127 );
or ( n34130 , n34126 , n34128 , n34129 );
xor ( n34131 , n33942 , n33944 );
xor ( n34132 , n33946 , n33947 );
and ( n34133 , n34131 , n34132 );
and ( n34134 , n31736 , n31076 );
and ( n34135 , n31464 , n31247 );
or ( n34136 , n34134 , n34135 );
and ( n34137 , n31084 , n31745 );
and ( n34138 , n31238 , n31442 );
or ( n34139 , n34137 , n34138 );
and ( n34140 , n34136 , n34139 );
and ( n34141 , n34132 , n34140 );
and ( n34142 , n34131 , n34140 );
or ( n34143 , n34133 , n34141 , n34142 );
and ( n34144 , n34130 , n34143 );
xor ( n34145 , n33887 , n33889 );
xor ( n34146 , n34145 , n33891 );
and ( n34147 , n34143 , n34146 );
and ( n34148 , n34130 , n34146 );
or ( n34149 , n34144 , n34147 , n34148 );
and ( n34150 , n34122 , n34149 );
and ( n34151 , n34059 , n34149 );
or ( n34152 , n34123 , n34150 , n34151 );
xor ( n34153 , n33809 , n33811 );
xor ( n34154 , n34153 , n33813 );
xor ( n34155 , n33828 , n33833 );
xor ( n34156 , n34155 , n33837 );
and ( n34157 , n34154 , n34156 );
xor ( n34158 , n33894 , n33939 );
xor ( n34159 , n34158 , n33967 );
and ( n34160 , n34156 , n34159 );
and ( n34161 , n34154 , n34159 );
or ( n34162 , n34157 , n34160 , n34161 );
and ( n34163 , n34152 , n34162 );
xor ( n34164 , n33739 , n33740 );
xor ( n34165 , n34164 , n33742 );
and ( n34166 , n34162 , n34165 );
and ( n34167 , n34152 , n34165 );
or ( n34168 , n34163 , n34166 , n34167 );
and ( n34169 , n34051 , n34168 );
and ( n34170 , n33977 , n34168 );
or ( n34171 , n34052 , n34169 , n34170 );
and ( n34172 , n33886 , n34171 );
xor ( n34173 , n33687 , n33689 );
xor ( n34174 , n34173 , n33731 );
xor ( n34175 , n33745 , n33798 );
xor ( n34176 , n34175 , n33843 );
and ( n34177 , n34174 , n34176 );
xor ( n34178 , n33848 , n33850 );
xor ( n34179 , n34178 , n33853 );
and ( n34180 , n34176 , n34179 );
and ( n34181 , n34174 , n34179 );
or ( n34182 , n34177 , n34180 , n34181 );
and ( n34183 , n34171 , n34182 );
and ( n34184 , n33886 , n34182 );
or ( n34185 , n34172 , n34183 , n34184 );
and ( n34186 , n33884 , n34185 );
xor ( n34187 , n33737 , n33862 );
xor ( n34188 , n34187 , n33865 );
and ( n34189 , n34185 , n34188 );
and ( n34190 , n33884 , n34188 );
or ( n34191 , n34186 , n34189 , n34190 );
and ( n34192 , n33882 , n34191 );
xor ( n34193 , n33677 , n33679 );
xor ( n34194 , n34193 , n33868 );
and ( n34195 , n34191 , n34194 );
and ( n34196 , n33882 , n34194 );
or ( n34197 , n34192 , n34195 , n34196 );
xor ( n34198 , n33675 , n33871 );
xor ( n34199 , n34198 , n33874 );
and ( n34200 , n34197 , n34199 );
xor ( n34201 , n33882 , n34191 );
xor ( n34202 , n34201 , n34194 );
xor ( n34203 , n33682 , n33684 );
xor ( n34204 , n34203 , n33734 );
xor ( n34205 , n33846 , n33856 );
xor ( n34206 , n34205 , n33859 );
and ( n34207 , n34204 , n34206 );
xor ( n34208 , n33746 , n33747 );
xor ( n34209 , n34208 , n33795 );
xor ( n34210 , n33802 , n33816 );
xor ( n34211 , n34210 , n33840 );
and ( n34212 , n34209 , n34211 );
xor ( n34213 , n33978 , n33979 );
xor ( n34214 , n33913 , n33928 );
xor ( n34215 , n34214 , n33936 );
xor ( n34216 , n33945 , n33948 );
xor ( n34217 , n34216 , n33964 );
and ( n34218 , n34215 , n34217 );
xor ( n34219 , n34013 , n34037 );
and ( n34220 , n34217 , n34219 );
and ( n34221 , n34215 , n34219 );
or ( n34222 , n34218 , n34220 , n34221 );
and ( n34223 , n34213 , n34222 );
xor ( n34224 , n34039 , n34040 );
xor ( n34225 , n34043 , n34044 );
and ( n34226 , n34224 , n34225 );
xor ( n34227 , n34010 , n34012 );
xor ( n34228 , n34034 , n34036 );
and ( n34229 , n34227 , n34228 );
and ( n34230 , n34225 , n34229 );
and ( n34231 , n34224 , n34229 );
or ( n34232 , n34226 , n34230 , n34231 );
and ( n34233 , n34222 , n34232 );
and ( n34234 , n34213 , n34232 );
or ( n34235 , n34223 , n34233 , n34234 );
and ( n34236 , n34211 , n34235 );
and ( n34237 , n34209 , n34235 );
or ( n34238 , n34212 , n34236 , n34237 );
xnor ( n34239 , n33930 , n33931 );
xnor ( n34240 , n33933 , n33934 );
and ( n34241 , n34239 , n34240 );
xor ( n34242 , n33950 , n33952 );
xor ( n34243 , n34242 , n33961 );
and ( n34244 , n34241 , n34243 );
xor ( n34245 , n34069 , n34079 );
and ( n34246 , n34243 , n34245 );
and ( n34247 , n34241 , n34245 );
or ( n34248 , n34244 , n34246 , n34247 );
xor ( n34249 , n34097 , n34114 );
xor ( n34250 , n34117 , n34118 );
and ( n34251 , n34249 , n34250 );
buf ( n34252 , n1249 );
buf ( n34253 , n34252 );
and ( n34254 , n30413 , n34253 );
and ( n34255 , n30709 , n32671 );
and ( n34256 , n34254 , n34255 );
and ( n34257 , n31088 , n31745 );
and ( n34258 , n34255 , n34257 );
and ( n34259 , n34254 , n34257 );
or ( n34260 , n34256 , n34258 , n34259 );
and ( n34261 , n30558 , n32932 );
and ( n34262 , n30603 , n32719 );
and ( n34263 , n34261 , n34262 );
and ( n34264 , n31084 , n31861 );
and ( n34265 , n34262 , n34264 );
and ( n34266 , n34261 , n34264 );
or ( n34267 , n34263 , n34265 , n34266 );
and ( n34268 , n34260 , n34267 );
and ( n34269 , n30419 , n34082 );
and ( n34270 , n30442 , n33905 );
and ( n34271 , n34269 , n34270 );
and ( n34272 , n30799 , n32348 );
and ( n34273 , n34270 , n34272 );
and ( n34274 , n34269 , n34272 );
or ( n34275 , n34271 , n34273 , n34274 );
and ( n34276 , n34267 , n34275 );
and ( n34277 , n34260 , n34275 );
or ( n34278 , n34268 , n34276 , n34277 );
buf ( n34279 , n1249 );
buf ( n34280 , n34279 );
and ( n34281 , n34280 , n30421 );
and ( n34282 , n32689 , n30700 );
and ( n34283 , n34281 , n34282 );
and ( n34284 , n31736 , n31073 );
and ( n34285 , n34282 , n34284 );
and ( n34286 , n34281 , n34284 );
or ( n34287 , n34283 , n34285 , n34286 );
and ( n34288 , n32949 , n30563 );
and ( n34289 , n32736 , n30592 );
and ( n34290 , n34288 , n34289 );
and ( n34291 , n31883 , n31076 );
and ( n34292 , n34289 , n34291 );
and ( n34293 , n34288 , n34291 );
or ( n34294 , n34290 , n34292 , n34293 );
and ( n34295 , n34287 , n34294 );
and ( n34296 , n34099 , n30424 );
and ( n34297 , n33896 , n30439 );
and ( n34298 , n34296 , n34297 );
and ( n34299 , n32365 , n30791 );
and ( n34300 , n34297 , n34299 );
and ( n34301 , n34296 , n34299 );
or ( n34302 , n34298 , n34300 , n34301 );
and ( n34303 , n34294 , n34302 );
and ( n34304 , n34287 , n34302 );
or ( n34305 , n34295 , n34303 , n34304 );
and ( n34306 , n34278 , n34305 );
and ( n34307 , n34250 , n34306 );
and ( n34308 , n34249 , n34306 );
or ( n34309 , n34251 , n34307 , n34308 );
and ( n34310 , n34248 , n34309 );
xor ( n34311 , n33990 , n33991 );
xor ( n34312 , n34311 , n33993 );
xor ( n34313 , n34107 , n34108 );
xor ( n34314 , n34313 , n34110 );
and ( n34315 , n34312 , n34314 );
xor ( n34316 , n33997 , n33998 );
xor ( n34317 , n34316 , n34000 );
and ( n34318 , n34314 , n34317 );
and ( n34319 , n34312 , n34317 );
or ( n34320 , n34315 , n34318 , n34319 );
xor ( n34321 , n34014 , n34015 );
xor ( n34322 , n34321 , n34017 );
xor ( n34323 , n34090 , n34091 );
xor ( n34324 , n34323 , n34093 );
and ( n34325 , n34322 , n34324 );
xor ( n34326 , n34021 , n34022 );
xor ( n34327 , n34326 , n34024 );
and ( n34328 , n34324 , n34327 );
and ( n34329 , n34322 , n34327 );
or ( n34330 , n34325 , n34328 , n34329 );
and ( n34331 , n34320 , n34330 );
and ( n34332 , n30803 , n32173 );
and ( n34333 , n31238 , n31590 );
and ( n34334 , n34332 , n34333 );
and ( n34335 , n31278 , n31442 );
and ( n34336 , n34333 , n34335 );
and ( n34337 , n34332 , n34335 );
or ( n34338 , n34334 , n34336 , n34337 );
and ( n34339 , n33896 , n30424 );
or ( n34340 , n34338 , n34339 );
and ( n34341 , n32155 , n30788 );
and ( n34342 , n31607 , n31247 );
and ( n34343 , n34341 , n34342 );
and ( n34344 , n31464 , n31301 );
and ( n34345 , n34342 , n34344 );
and ( n34346 , n34341 , n34344 );
or ( n34347 , n34343 , n34345 , n34346 );
and ( n34348 , n30419 , n33905 );
or ( n34349 , n34347 , n34348 );
and ( n34350 , n34340 , n34349 );
and ( n34351 , n34331 , n34350 );
and ( n34352 , n30468 , n33347 );
and ( n34353 , n30503 , n33296 );
and ( n34354 , n34352 , n34353 );
and ( n34355 , n30889 , n32066 );
and ( n34356 , n34353 , n34355 );
and ( n34357 , n34352 , n34355 );
or ( n34358 , n34354 , n34356 , n34357 );
xor ( n34359 , n34083 , n34084 );
xor ( n34360 , n34359 , n34086 );
or ( n34361 , n34358 , n34360 );
and ( n34362 , n33304 , n30473 );
and ( n34363 , n33339 , n30508 );
and ( n34364 , n34362 , n34363 );
and ( n34365 , n32057 , n30898 );
and ( n34366 , n34363 , n34365 );
and ( n34367 , n34362 , n34365 );
or ( n34368 , n34364 , n34366 , n34367 );
xor ( n34369 , n34100 , n34101 );
xor ( n34370 , n34369 , n34103 );
or ( n34371 , n34368 , n34370 );
and ( n34372 , n34361 , n34371 );
and ( n34373 , n34350 , n34372 );
and ( n34374 , n34331 , n34372 );
or ( n34375 , n34351 , n34373 , n34374 );
and ( n34376 , n34309 , n34375 );
and ( n34377 , n34248 , n34375 );
or ( n34378 , n34310 , n34376 , n34377 );
xor ( n34379 , n34061 , n34063 );
xor ( n34380 , n34379 , n34066 );
xor ( n34381 , n34071 , n34073 );
xor ( n34382 , n34381 , n34076 );
and ( n34383 , n34380 , n34382 );
xor ( n34384 , n34020 , n34027 );
xor ( n34385 , n34384 , n34030 );
xor ( n34386 , n33996 , n34003 );
xor ( n34387 , n34386 , n34006 );
and ( n34388 , n34385 , n34387 );
and ( n34389 , n34383 , n34388 );
xnor ( n34390 , n34089 , n34096 );
xnor ( n34391 , n34106 , n34113 );
and ( n34392 , n34390 , n34391 );
and ( n34393 , n34388 , n34392 );
and ( n34394 , n34383 , n34392 );
or ( n34395 , n34389 , n34393 , n34394 );
xor ( n34396 , n33954 , n33955 );
xor ( n34397 , n34396 , n33958 );
xor ( n34398 , n34136 , n34139 );
and ( n34399 , n34397 , n34398 );
xor ( n34400 , n34239 , n34240 );
and ( n34401 , n34398 , n34400 );
and ( n34402 , n34397 , n34400 );
or ( n34403 , n34399 , n34401 , n34402 );
xor ( n34404 , n34124 , n34125 );
xor ( n34405 , n34404 , n34127 );
and ( n34406 , n34403 , n34405 );
xor ( n34407 , n34131 , n34132 );
xor ( n34408 , n34407 , n34140 );
and ( n34409 , n34405 , n34408 );
and ( n34410 , n34403 , n34408 );
or ( n34411 , n34406 , n34409 , n34410 );
and ( n34412 , n34395 , n34411 );
xor ( n34413 , n34053 , n34054 );
xor ( n34414 , n34413 , n34056 );
and ( n34415 , n34411 , n34414 );
and ( n34416 , n34395 , n34414 );
or ( n34417 , n34412 , n34415 , n34416 );
and ( n34418 , n34378 , n34417 );
xor ( n34419 , n33982 , n33983 );
xor ( n34420 , n34419 , n33985 );
and ( n34421 , n34417 , n34420 );
and ( n34422 , n34378 , n34420 );
or ( n34423 , n34418 , n34421 , n34422 );
xor ( n34424 , n34038 , n34041 );
xor ( n34425 , n34424 , n34045 );
xor ( n34426 , n34059 , n34122 );
xor ( n34427 , n34426 , n34149 );
and ( n34428 , n34425 , n34427 );
xor ( n34429 , n34154 , n34156 );
xor ( n34430 , n34429 , n34159 );
and ( n34431 , n34427 , n34430 );
and ( n34432 , n34425 , n34430 );
or ( n34433 , n34428 , n34431 , n34432 );
and ( n34434 , n34423 , n34433 );
xor ( n34435 , n33970 , n33972 );
xor ( n34436 , n34435 , n33974 );
and ( n34437 , n34433 , n34436 );
and ( n34438 , n34423 , n34436 );
or ( n34439 , n34434 , n34437 , n34438 );
and ( n34440 , n34238 , n34439 );
xor ( n34441 , n33977 , n34051 );
xor ( n34442 , n34441 , n34168 );
and ( n34443 , n34439 , n34442 );
and ( n34444 , n34238 , n34442 );
or ( n34445 , n34440 , n34443 , n34444 );
and ( n34446 , n34206 , n34445 );
and ( n34447 , n34204 , n34445 );
or ( n34448 , n34207 , n34446 , n34447 );
xor ( n34449 , n33884 , n34185 );
xor ( n34450 , n34449 , n34188 );
and ( n34451 , n34448 , n34450 );
xor ( n34452 , n33886 , n34171 );
xor ( n34453 , n34452 , n34182 );
xor ( n34454 , n34174 , n34176 );
xor ( n34455 , n34454 , n34179 );
xor ( n34456 , n33980 , n33988 );
xor ( n34457 , n34456 , n34048 );
xor ( n34458 , n34152 , n34162 );
xor ( n34459 , n34458 , n34165 );
and ( n34460 , n34457 , n34459 );
xor ( n34461 , n34080 , n34115 );
xor ( n34462 , n34461 , n34119 );
xor ( n34463 , n34130 , n34143 );
xor ( n34464 , n34463 , n34146 );
and ( n34465 , n34462 , n34464 );
xor ( n34466 , n34227 , n34228 );
buf ( n34467 , n31278 );
buf ( n34468 , n15862 );
buf ( n34469 , n34468 );
and ( n34470 , n34467 , n34469 );
not ( n34471 , n34470 );
xnor ( n34472 , n34338 , n34339 );
xnor ( n34473 , n34347 , n34348 );
and ( n34474 , n34472 , n34473 );
and ( n34475 , n34471 , n34474 );
and ( n34476 , n34466 , n34475 );
buf ( n34477 , n34470 );
and ( n34478 , n34475 , n34477 );
and ( n34479 , n34466 , n34477 );
or ( n34480 , n34476 , n34478 , n34479 );
and ( n34481 , n34464 , n34480 );
and ( n34482 , n34462 , n34480 );
or ( n34483 , n34465 , n34481 , n34482 );
and ( n34484 , n33692 , n30473 );
and ( n34485 , n33304 , n30508 );
and ( n34486 , n34484 , n34485 );
and ( n34487 , n32365 , n30788 );
and ( n34488 , n34485 , n34487 );
and ( n34489 , n34484 , n34487 );
or ( n34490 , n34486 , n34488 , n34489 );
xor ( n34491 , n34352 , n34353 );
xor ( n34492 , n34491 , n34355 );
and ( n34493 , n34490 , n34492 );
xor ( n34494 , n34332 , n34333 );
xor ( n34495 , n34494 , n34335 );
and ( n34496 , n34492 , n34495 );
and ( n34497 , n34490 , n34495 );
or ( n34498 , n34493 , n34496 , n34497 );
xor ( n34499 , n34287 , n34294 );
xor ( n34500 , n34499 , n34302 );
or ( n34501 , n34498 , n34500 );
and ( n34502 , n30468 , n33712 );
and ( n34503 , n30503 , n33347 );
and ( n34504 , n34502 , n34503 );
and ( n34505 , n30803 , n32348 );
and ( n34506 , n34503 , n34505 );
and ( n34507 , n34502 , n34505 );
or ( n34508 , n34504 , n34506 , n34507 );
xor ( n34509 , n34362 , n34363 );
xor ( n34510 , n34509 , n34365 );
and ( n34511 , n34508 , n34510 );
xor ( n34512 , n34341 , n34342 );
xor ( n34513 , n34512 , n34344 );
and ( n34514 , n34510 , n34513 );
and ( n34515 , n34508 , n34513 );
or ( n34516 , n34511 , n34514 , n34515 );
xor ( n34517 , n34260 , n34267 );
xor ( n34518 , n34517 , n34275 );
or ( n34519 , n34516 , n34518 );
and ( n34520 , n34501 , n34519 );
xor ( n34521 , n34322 , n34324 );
xor ( n34522 , n34521 , n34327 );
xnor ( n34523 , n34368 , n34370 );
or ( n34524 , n34522 , n34523 );
xor ( n34525 , n34312 , n34314 );
xor ( n34526 , n34525 , n34317 );
xnor ( n34527 , n34358 , n34360 );
or ( n34528 , n34526 , n34527 );
and ( n34529 , n34524 , n34528 );
and ( n34530 , n34520 , n34529 );
and ( n34531 , n30464 , n33712 );
and ( n34532 , n33692 , n30461 );
and ( n34533 , n34531 , n34532 );
xor ( n34534 , n34467 , n34469 );
and ( n34535 , n34533 , n34534 );
xnor ( n34536 , n34134 , n34135 );
xnor ( n34537 , n34137 , n34138 );
and ( n34538 , n34536 , n34537 );
and ( n34539 , n34535 , n34538 );
xor ( n34540 , n34278 , n34305 );
and ( n34541 , n34538 , n34540 );
and ( n34542 , n34535 , n34540 );
or ( n34543 , n34539 , n34541 , n34542 );
and ( n34544 , n34529 , n34543 );
and ( n34545 , n34520 , n34543 );
or ( n34546 , n34530 , n34544 , n34545 );
xor ( n34547 , n34320 , n34330 );
xor ( n34548 , n34340 , n34349 );
and ( n34549 , n34547 , n34548 );
xor ( n34550 , n34361 , n34371 );
and ( n34551 , n34548 , n34550 );
and ( n34552 , n34547 , n34550 );
or ( n34553 , n34549 , n34551 , n34552 );
xor ( n34554 , n34380 , n34382 );
xor ( n34555 , n34385 , n34387 );
and ( n34556 , n34554 , n34555 );
xor ( n34557 , n34390 , n34391 );
and ( n34558 , n34555 , n34557 );
and ( n34559 , n34554 , n34557 );
or ( n34560 , n34556 , n34558 , n34559 );
and ( n34561 , n34553 , n34560 );
xor ( n34562 , n34254 , n34255 );
xor ( n34563 , n34562 , n34257 );
xor ( n34564 , n34261 , n34262 );
xor ( n34565 , n34564 , n34264 );
and ( n34566 , n34563 , n34565 );
xor ( n34567 , n34281 , n34282 );
xor ( n34568 , n34567 , n34284 );
xor ( n34569 , n34288 , n34289 );
xor ( n34570 , n34569 , n34291 );
and ( n34571 , n34568 , n34570 );
and ( n34572 , n34566 , n34571 );
xor ( n34573 , n34533 , n34534 );
xor ( n34574 , n34536 , n34537 );
and ( n34575 , n34573 , n34574 );
and ( n34576 , n34099 , n30439 );
and ( n34577 , n33896 , n30461 );
and ( n34578 , n34576 , n34577 );
and ( n34579 , n30442 , n34082 );
and ( n34580 , n30464 , n33905 );
and ( n34581 , n34579 , n34580 );
and ( n34582 , n34578 , n34581 );
and ( n34583 , n34574 , n34582 );
and ( n34584 , n34573 , n34582 );
or ( n34585 , n34575 , n34583 , n34584 );
and ( n34586 , n34572 , n34585 );
xor ( n34587 , n34397 , n34398 );
xor ( n34588 , n34587 , n34400 );
and ( n34589 , n34585 , n34588 );
and ( n34590 , n34572 , n34588 );
or ( n34591 , n34586 , n34589 , n34590 );
and ( n34592 , n34560 , n34591 );
and ( n34593 , n34553 , n34591 );
or ( n34594 , n34561 , n34592 , n34593 );
and ( n34595 , n34546 , n34594 );
xor ( n34596 , n34241 , n34243 );
xor ( n34597 , n34596 , n34245 );
xor ( n34598 , n34249 , n34250 );
xor ( n34599 , n34598 , n34306 );
and ( n34600 , n34597 , n34599 );
xor ( n34601 , n34331 , n34350 );
xor ( n34602 , n34601 , n34372 );
and ( n34603 , n34599 , n34602 );
and ( n34604 , n34597 , n34602 );
or ( n34605 , n34600 , n34603 , n34604 );
and ( n34606 , n34594 , n34605 );
and ( n34607 , n34546 , n34605 );
or ( n34608 , n34595 , n34606 , n34607 );
and ( n34609 , n34483 , n34608 );
xor ( n34610 , n34215 , n34217 );
xor ( n34611 , n34610 , n34219 );
xor ( n34612 , n34224 , n34225 );
xor ( n34613 , n34612 , n34229 );
and ( n34614 , n34611 , n34613 );
xor ( n34615 , n34248 , n34309 );
xor ( n34616 , n34615 , n34375 );
and ( n34617 , n34613 , n34616 );
and ( n34618 , n34611 , n34616 );
or ( n34619 , n34614 , n34617 , n34618 );
and ( n34620 , n34608 , n34619 );
and ( n34621 , n34483 , n34619 );
or ( n34622 , n34609 , n34620 , n34621 );
and ( n34623 , n34459 , n34622 );
and ( n34624 , n34457 , n34622 );
or ( n34625 , n34460 , n34623 , n34624 );
and ( n34626 , n34455 , n34625 );
xor ( n34627 , n34213 , n34222 );
xor ( n34628 , n34627 , n34232 );
xor ( n34629 , n34378 , n34417 );
xor ( n34630 , n34629 , n34420 );
and ( n34631 , n34628 , n34630 );
xor ( n34632 , n34425 , n34427 );
xor ( n34633 , n34632 , n34430 );
and ( n34634 , n34630 , n34633 );
and ( n34635 , n34628 , n34633 );
or ( n34636 , n34631 , n34634 , n34635 );
xor ( n34637 , n34209 , n34211 );
xor ( n34638 , n34637 , n34235 );
and ( n34639 , n34636 , n34638 );
xor ( n34640 , n34423 , n34433 );
xor ( n34641 , n34640 , n34436 );
and ( n34642 , n34638 , n34641 );
and ( n34643 , n34636 , n34641 );
or ( n34644 , n34639 , n34642 , n34643 );
and ( n34645 , n34625 , n34644 );
and ( n34646 , n34455 , n34644 );
or ( n34647 , n34626 , n34645 , n34646 );
and ( n34648 , n34453 , n34647 );
xor ( n34649 , n34204 , n34206 );
xor ( n34650 , n34649 , n34445 );
and ( n34651 , n34647 , n34650 );
and ( n34652 , n34453 , n34650 );
or ( n34653 , n34648 , n34651 , n34652 );
and ( n34654 , n34450 , n34653 );
and ( n34655 , n34448 , n34653 );
or ( n34656 , n34451 , n34654 , n34655 );
and ( n34657 , n34202 , n34656 );
xor ( n34658 , n34448 , n34450 );
xor ( n34659 , n34658 , n34653 );
xor ( n34660 , n34238 , n34439 );
xor ( n34661 , n34660 , n34442 );
xor ( n34662 , n34395 , n34411 );
xor ( n34663 , n34662 , n34414 );
xor ( n34664 , n34383 , n34388 );
xor ( n34665 , n34664 , n34392 );
xor ( n34666 , n34403 , n34405 );
xor ( n34667 , n34666 , n34408 );
and ( n34668 , n34665 , n34667 );
and ( n34669 , n30603 , n32932 );
and ( n34670 , n30709 , n32719 );
and ( n34671 , n34669 , n34670 );
and ( n34672 , n31084 , n32066 );
and ( n34673 , n34670 , n34672 );
and ( n34674 , n34669 , n34672 );
or ( n34675 , n34671 , n34673 , n34674 );
and ( n34676 , n30558 , n33296 );
and ( n34677 , n30889 , n32173 );
and ( n34678 , n34676 , n34677 );
and ( n34679 , n31238 , n31745 );
and ( n34680 , n34677 , n34679 );
and ( n34681 , n34676 , n34679 );
or ( n34682 , n34678 , n34680 , n34681 );
and ( n34683 , n34675 , n34682 );
and ( n34684 , n30419 , n34253 );
and ( n34685 , n30799 , n32671 );
and ( n34686 , n34684 , n34685 );
and ( n34687 , n31088 , n31861 );
and ( n34688 , n34685 , n34687 );
and ( n34689 , n34684 , n34687 );
or ( n34690 , n34686 , n34688 , n34689 );
and ( n34691 , n34682 , n34690 );
and ( n34692 , n34675 , n34690 );
or ( n34693 , n34683 , n34691 , n34692 );
and ( n34694 , n32949 , n30592 );
and ( n34695 , n32736 , n30700 );
and ( n34696 , n34694 , n34695 );
and ( n34697 , n32057 , n31076 );
and ( n34698 , n34695 , n34697 );
and ( n34699 , n34694 , n34697 );
or ( n34700 , n34696 , n34698 , n34699 );
and ( n34701 , n33339 , n30563 );
and ( n34702 , n32155 , n30898 );
and ( n34703 , n34701 , n34702 );
and ( n34704 , n31736 , n31247 );
and ( n34705 , n34702 , n34704 );
and ( n34706 , n34701 , n34704 );
or ( n34707 , n34703 , n34705 , n34706 );
and ( n34708 , n34700 , n34707 );
and ( n34709 , n34280 , n30424 );
and ( n34710 , n32689 , n30791 );
and ( n34711 , n34709 , n34710 );
and ( n34712 , n31883 , n31073 );
and ( n34713 , n34710 , n34712 );
and ( n34714 , n34709 , n34712 );
or ( n34715 , n34711 , n34713 , n34714 );
and ( n34716 , n34707 , n34715 );
and ( n34717 , n34700 , n34715 );
or ( n34718 , n34708 , n34716 , n34717 );
and ( n34719 , n34693 , n34718 );
xor ( n34720 , n34471 , n34474 );
or ( n34721 , n34719 , n34720 );
and ( n34722 , n34667 , n34721 );
and ( n34723 , n34665 , n34721 );
or ( n34724 , n34668 , n34722 , n34723 );
and ( n34725 , n34663 , n34724 );
xor ( n34726 , n34501 , n34519 );
xor ( n34727 , n34524 , n34528 );
and ( n34728 , n34726 , n34727 );
and ( n34729 , n33896 , n30473 );
and ( n34730 , n33692 , n30508 );
and ( n34731 , n34729 , n34730 );
and ( n34732 , n32155 , n31076 );
and ( n34733 , n34730 , n34732 );
and ( n34734 , n34729 , n34732 );
or ( n34735 , n34731 , n34733 , n34734 );
and ( n34736 , n32949 , n30700 );
and ( n34737 , n32736 , n30791 );
and ( n34738 , n34736 , n34737 );
and ( n34739 , n31883 , n31247 );
and ( n34740 , n34737 , n34739 );
and ( n34741 , n34736 , n34739 );
or ( n34742 , n34738 , n34740 , n34741 );
and ( n34743 , n34735 , n34742 );
and ( n34744 , n33304 , n30563 );
and ( n34745 , n33339 , n30592 );
and ( n34746 , n34744 , n34745 );
and ( n34747 , n32057 , n31073 );
and ( n34748 , n34745 , n34747 );
and ( n34749 , n34744 , n34747 );
or ( n34750 , n34746 , n34748 , n34749 );
and ( n34751 , n34742 , n34750 );
and ( n34752 , n34735 , n34750 );
or ( n34753 , n34743 , n34751 , n34752 );
xor ( n34754 , n34269 , n34270 );
xor ( n34755 , n34754 , n34272 );
or ( n34756 , n34753 , n34755 );
and ( n34757 , n30468 , n33905 );
and ( n34758 , n30503 , n33712 );
and ( n34759 , n34757 , n34758 );
and ( n34760 , n31084 , n32173 );
and ( n34761 , n34758 , n34760 );
and ( n34762 , n34757 , n34760 );
or ( n34763 , n34759 , n34761 , n34762 );
and ( n34764 , n30709 , n32932 );
and ( n34765 , n30799 , n32719 );
and ( n34766 , n34764 , n34765 );
and ( n34767 , n31238 , n31861 );
and ( n34768 , n34765 , n34767 );
and ( n34769 , n34764 , n34767 );
or ( n34770 , n34766 , n34768 , n34769 );
and ( n34771 , n34763 , n34770 );
and ( n34772 , n30558 , n33347 );
and ( n34773 , n30603 , n33296 );
and ( n34774 , n34772 , n34773 );
and ( n34775 , n31088 , n32066 );
and ( n34776 , n34773 , n34775 );
and ( n34777 , n34772 , n34775 );
or ( n34778 , n34774 , n34776 , n34777 );
and ( n34779 , n34770 , n34778 );
and ( n34780 , n34763 , n34778 );
or ( n34781 , n34771 , n34779 , n34780 );
xor ( n34782 , n34296 , n34297 );
xor ( n34783 , n34782 , n34299 );
or ( n34784 , n34781 , n34783 );
and ( n34785 , n34756 , n34784 );
and ( n34786 , n34727 , n34785 );
and ( n34787 , n34726 , n34785 );
or ( n34788 , n34728 , n34786 , n34787 );
xnor ( n34789 , n34498 , n34500 );
xnor ( n34790 , n34516 , n34518 );
and ( n34791 , n34789 , n34790 );
xnor ( n34792 , n34522 , n34523 );
xnor ( n34793 , n34526 , n34527 );
and ( n34794 , n34792 , n34793 );
and ( n34795 , n34791 , n34794 );
xor ( n34796 , n34693 , n34718 );
xor ( n34797 , n34566 , n34571 );
and ( n34798 , n34796 , n34797 );
xor ( n34799 , n34472 , n34473 );
and ( n34800 , n34797 , n34799 );
and ( n34801 , n34796 , n34799 );
or ( n34802 , n34798 , n34800 , n34801 );
and ( n34803 , n34794 , n34802 );
and ( n34804 , n34791 , n34802 );
or ( n34805 , n34795 , n34803 , n34804 );
and ( n34806 , n34788 , n34805 );
xor ( n34807 , n34502 , n34503 );
xor ( n34808 , n34807 , n34505 );
xor ( n34809 , n34669 , n34670 );
xor ( n34810 , n34809 , n34672 );
or ( n34811 , n34808 , n34810 );
xor ( n34812 , n34484 , n34485 );
xor ( n34813 , n34812 , n34487 );
xor ( n34814 , n34694 , n34695 );
xor ( n34815 , n34814 , n34697 );
or ( n34816 , n34813 , n34815 );
and ( n34817 , n34811 , n34816 );
and ( n34818 , n30442 , n34253 );
and ( n34819 , n30464 , n34082 );
and ( n34820 , n34818 , n34819 );
and ( n34821 , n30803 , n32671 );
and ( n34822 , n34819 , n34821 );
and ( n34823 , n34818 , n34821 );
or ( n34824 , n34820 , n34822 , n34823 );
and ( n34825 , n30889 , n32348 );
and ( n34826 , n31278 , n31745 );
and ( n34827 , n34825 , n34826 );
and ( n34828 , n31464 , n31590 );
and ( n34829 , n34826 , n34828 );
and ( n34830 , n34825 , n34828 );
or ( n34831 , n34827 , n34829 , n34830 );
or ( n34832 , n34824 , n34831 );
and ( n34833 , n34280 , n30439 );
and ( n34834 , n34099 , n30461 );
and ( n34835 , n34833 , n34834 );
and ( n34836 , n32689 , n30788 );
and ( n34837 , n34834 , n34836 );
and ( n34838 , n34833 , n34836 );
or ( n34839 , n34835 , n34837 , n34838 );
and ( n34840 , n32365 , n30898 );
and ( n34841 , n31736 , n31301 );
and ( n34842 , n34840 , n34841 );
and ( n34843 , n31607 , n31442 );
and ( n34844 , n34841 , n34843 );
and ( n34845 , n34840 , n34843 );
or ( n34846 , n34842 , n34844 , n34845 );
or ( n34847 , n34839 , n34846 );
and ( n34848 , n34832 , n34847 );
and ( n34849 , n34817 , n34848 );
xor ( n34850 , n34676 , n34677 );
xor ( n34851 , n34850 , n34679 );
xor ( n34852 , n34684 , n34685 );
xor ( n34853 , n34852 , n34687 );
or ( n34854 , n34851 , n34853 );
xor ( n34855 , n34701 , n34702 );
xor ( n34856 , n34855 , n34704 );
xor ( n34857 , n34709 , n34710 );
xor ( n34858 , n34857 , n34712 );
or ( n34859 , n34856 , n34858 );
and ( n34860 , n34854 , n34859 );
and ( n34861 , n34848 , n34860 );
and ( n34862 , n34817 , n34860 );
or ( n34863 , n34849 , n34861 , n34862 );
xor ( n34864 , n34675 , n34682 );
xor ( n34865 , n34864 , n34690 );
xor ( n34866 , n34700 , n34707 );
xor ( n34867 , n34866 , n34715 );
and ( n34868 , n34865 , n34867 );
xor ( n34869 , n34508 , n34510 );
xor ( n34870 , n34869 , n34513 );
xor ( n34871 , n34490 , n34492 );
xor ( n34872 , n34871 , n34495 );
and ( n34873 , n34870 , n34872 );
and ( n34874 , n34868 , n34873 );
xor ( n34875 , n34563 , n34565 );
xor ( n34876 , n34568 , n34570 );
and ( n34877 , n34875 , n34876 );
and ( n34878 , n34873 , n34877 );
and ( n34879 , n34868 , n34877 );
or ( n34880 , n34874 , n34878 , n34879 );
and ( n34881 , n34863 , n34880 );
xor ( n34882 , n34535 , n34538 );
xor ( n34883 , n34882 , n34540 );
and ( n34884 , n34880 , n34883 );
and ( n34885 , n34863 , n34883 );
or ( n34886 , n34881 , n34884 , n34885 );
and ( n34887 , n34805 , n34886 );
and ( n34888 , n34788 , n34886 );
or ( n34889 , n34806 , n34887 , n34888 );
and ( n34890 , n34724 , n34889 );
and ( n34891 , n34663 , n34889 );
or ( n34892 , n34725 , n34890 , n34891 );
xor ( n34893 , n34547 , n34548 );
xor ( n34894 , n34893 , n34550 );
xor ( n34895 , n34554 , n34555 );
xor ( n34896 , n34895 , n34557 );
and ( n34897 , n34894 , n34896 );
xor ( n34898 , n34572 , n34585 );
xor ( n34899 , n34898 , n34588 );
and ( n34900 , n34896 , n34899 );
and ( n34901 , n34894 , n34899 );
or ( n34902 , n34897 , n34900 , n34901 );
xor ( n34903 , n34466 , n34475 );
xor ( n34904 , n34903 , n34477 );
and ( n34905 , n34902 , n34904 );
xor ( n34906 , n34520 , n34529 );
xor ( n34907 , n34906 , n34543 );
and ( n34908 , n34904 , n34907 );
and ( n34909 , n34902 , n34907 );
or ( n34910 , n34905 , n34908 , n34909 );
xor ( n34911 , n34462 , n34464 );
xor ( n34912 , n34911 , n34480 );
and ( n34913 , n34910 , n34912 );
xor ( n34914 , n34546 , n34594 );
xor ( n34915 , n34914 , n34605 );
and ( n34916 , n34912 , n34915 );
and ( n34917 , n34910 , n34915 );
or ( n34918 , n34913 , n34916 , n34917 );
and ( n34919 , n34892 , n34918 );
xor ( n34920 , n34483 , n34608 );
xor ( n34921 , n34920 , n34619 );
and ( n34922 , n34918 , n34921 );
and ( n34923 , n34892 , n34921 );
or ( n34924 , n34919 , n34922 , n34923 );
xor ( n34925 , n34457 , n34459 );
xor ( n34926 , n34925 , n34622 );
and ( n34927 , n34924 , n34926 );
xor ( n34928 , n34636 , n34638 );
xor ( n34929 , n34928 , n34641 );
and ( n34930 , n34926 , n34929 );
and ( n34931 , n34924 , n34929 );
or ( n34932 , n34927 , n34930 , n34931 );
and ( n34933 , n34661 , n34932 );
xor ( n34934 , n34455 , n34625 );
xor ( n34935 , n34934 , n34644 );
and ( n34936 , n34932 , n34935 );
and ( n34937 , n34661 , n34935 );
or ( n34938 , n34933 , n34936 , n34937 );
xor ( n34939 , n34453 , n34647 );
xor ( n34940 , n34939 , n34650 );
and ( n34941 , n34938 , n34940 );
xor ( n34942 , n34661 , n34932 );
xor ( n34943 , n34942 , n34935 );
xor ( n34944 , n34628 , n34630 );
xor ( n34945 , n34944 , n34633 );
xor ( n34946 , n34611 , n34613 );
xor ( n34947 , n34946 , n34616 );
xor ( n34948 , n34553 , n34560 );
xor ( n34949 , n34948 , n34591 );
xor ( n34950 , n34597 , n34599 );
xor ( n34951 , n34950 , n34602 );
and ( n34952 , n34949 , n34951 );
xnor ( n34953 , n34719 , n34720 );
xor ( n34954 , n34531 , n34532 );
buf ( n34955 , n31464 );
buf ( n34956 , n15868 );
buf ( n34957 , n34956 );
and ( n34958 , n34955 , n34957 );
and ( n34959 , n34954 , n34958 );
xor ( n34960 , n34578 , n34581 );
and ( n34961 , n34958 , n34960 );
and ( n34962 , n34954 , n34960 );
or ( n34963 , n34959 , n34961 , n34962 );
xor ( n34964 , n34573 , n34574 );
xor ( n34965 , n34964 , n34582 );
and ( n34966 , n34963 , n34965 );
xor ( n34967 , n34756 , n34784 );
and ( n34968 , n34965 , n34967 );
and ( n34969 , n34963 , n34967 );
or ( n34970 , n34966 , n34968 , n34969 );
and ( n34971 , n34953 , n34970 );
xor ( n34972 , n34789 , n34790 );
xor ( n34973 , n34792 , n34793 );
and ( n34974 , n34972 , n34973 );
xor ( n34975 , n34955 , n34957 );
and ( n34976 , n31464 , n31745 );
and ( n34977 , n31736 , n31442 );
and ( n34978 , n34976 , n34977 );
buf ( n34979 , n15871 );
buf ( n34980 , n34979 );
and ( n34981 , n34978 , n34980 );
and ( n34982 , n34975 , n34981 );
and ( n34983 , n32949 , n30791 );
and ( n34984 , n32736 , n30788 );
and ( n34985 , n34983 , n34984 );
and ( n34986 , n32057 , n31247 );
and ( n34987 , n34984 , n34986 );
and ( n34988 , n34983 , n34986 );
or ( n34989 , n34985 , n34987 , n34988 );
and ( n34990 , n30799 , n32932 );
and ( n34991 , n30803 , n32719 );
and ( n34992 , n34990 , n34991 );
and ( n34993 , n31238 , n32066 );
and ( n34994 , n34991 , n34993 );
and ( n34995 , n34990 , n34993 );
or ( n34996 , n34992 , n34994 , n34995 );
and ( n34997 , n34989 , n34996 );
and ( n34998 , n34981 , n34997 );
and ( n34999 , n34975 , n34997 );
or ( n35000 , n34982 , n34998 , n34999 );
not ( n35001 , n35000 );
xnor ( n35002 , n34851 , n34853 );
xnor ( n35003 , n34856 , n34858 );
and ( n35004 , n35002 , n35003 );
and ( n35005 , n35001 , n35004 );
and ( n35006 , n34973 , n35005 );
and ( n35007 , n34972 , n35005 );
or ( n35008 , n34974 , n35006 , n35007 );
and ( n35009 , n34970 , n35008 );
and ( n35010 , n34953 , n35008 );
or ( n35011 , n34971 , n35009 , n35010 );
and ( n35012 , n34951 , n35011 );
and ( n35013 , n34949 , n35011 );
or ( n35014 , n34952 , n35012 , n35013 );
and ( n35015 , n34947 , n35014 );
buf ( n35016 , n35000 );
and ( n35017 , n31607 , n31301 );
xnor ( n35018 , n34839 , n34846 );
or ( n35019 , n35017 , n35018 );
and ( n35020 , n31278 , n31590 );
xnor ( n35021 , n34824 , n34831 );
or ( n35022 , n35020 , n35021 );
and ( n35023 , n35019 , n35022 );
and ( n35024 , n35016 , n35023 );
and ( n35025 , n34099 , n30473 );
and ( n35026 , n33896 , n30508 );
and ( n35027 , n35025 , n35026 );
and ( n35028 , n32689 , n30898 );
and ( n35029 , n35026 , n35028 );
and ( n35030 , n35025 , n35028 );
or ( n35031 , n35027 , n35029 , n35030 );
and ( n35032 , n33692 , n30563 );
and ( n35033 , n32365 , n31076 );
and ( n35034 , n35032 , n35033 );
and ( n35035 , n31883 , n31301 );
and ( n35036 , n35033 , n35035 );
and ( n35037 , n35032 , n35035 );
or ( n35038 , n35034 , n35036 , n35037 );
and ( n35039 , n35031 , n35038 );
and ( n35040 , n33304 , n30592 );
and ( n35041 , n33339 , n30700 );
and ( n35042 , n35040 , n35041 );
and ( n35043 , n32155 , n31073 );
and ( n35044 , n35041 , n35043 );
and ( n35045 , n35040 , n35043 );
or ( n35046 , n35042 , n35044 , n35045 );
and ( n35047 , n35038 , n35046 );
and ( n35048 , n35031 , n35046 );
or ( n35049 , n35039 , n35047 , n35048 );
xor ( n35050 , n34735 , n34742 );
xor ( n35051 , n35050 , n34750 );
or ( n35052 , n35049 , n35051 );
and ( n35053 , n30468 , n34082 );
and ( n35054 , n30503 , n33905 );
and ( n35055 , n35053 , n35054 );
and ( n35056 , n30889 , n32671 );
and ( n35057 , n35054 , n35056 );
and ( n35058 , n35053 , n35056 );
or ( n35059 , n35055 , n35057 , n35058 );
and ( n35060 , n30558 , n33712 );
and ( n35061 , n31084 , n32348 );
and ( n35062 , n35060 , n35061 );
and ( n35063 , n31278 , n31861 );
and ( n35064 , n35061 , n35063 );
and ( n35065 , n35060 , n35063 );
or ( n35066 , n35062 , n35064 , n35065 );
and ( n35067 , n35059 , n35066 );
and ( n35068 , n30603 , n33347 );
and ( n35069 , n30709 , n33296 );
and ( n35070 , n35068 , n35069 );
and ( n35071 , n31088 , n32173 );
and ( n35072 , n35069 , n35071 );
and ( n35073 , n35068 , n35071 );
or ( n35074 , n35070 , n35072 , n35073 );
and ( n35075 , n35066 , n35074 );
and ( n35076 , n35059 , n35074 );
or ( n35077 , n35067 , n35075 , n35076 );
xor ( n35078 , n34763 , n34770 );
xor ( n35079 , n35078 , n34778 );
or ( n35080 , n35077 , n35079 );
and ( n35081 , n35052 , n35080 );
and ( n35082 , n35023 , n35081 );
and ( n35083 , n35016 , n35081 );
or ( n35084 , n35024 , n35082 , n35083 );
xnor ( n35085 , n34753 , n34755 );
xnor ( n35086 , n34781 , n34783 );
and ( n35087 , n35085 , n35086 );
xor ( n35088 , n34576 , n34577 );
xor ( n35089 , n34579 , n34580 );
and ( n35090 , n35088 , n35089 );
xor ( n35091 , n34811 , n34816 );
and ( n35092 , n35090 , n35091 );
xor ( n35093 , n34832 , n34847 );
and ( n35094 , n35091 , n35093 );
and ( n35095 , n35090 , n35093 );
or ( n35096 , n35092 , n35094 , n35095 );
and ( n35097 , n35087 , n35096 );
xor ( n35098 , n34854 , n34859 );
xor ( n35099 , n34865 , n34867 );
and ( n35100 , n35098 , n35099 );
xor ( n35101 , n34870 , n34872 );
and ( n35102 , n35099 , n35101 );
and ( n35103 , n35098 , n35101 );
or ( n35104 , n35100 , n35102 , n35103 );
and ( n35105 , n35096 , n35104 );
and ( n35106 , n35087 , n35104 );
or ( n35107 , n35097 , n35105 , n35106 );
and ( n35108 , n35084 , n35107 );
xor ( n35109 , n34875 , n34876 );
xor ( n35110 , n34833 , n34834 );
xor ( n35111 , n35110 , n34836 );
xor ( n35112 , n34840 , n34841 );
xor ( n35113 , n35112 , n34843 );
and ( n35114 , n35111 , n35113 );
xor ( n35115 , n34729 , n34730 );
xor ( n35116 , n35115 , n34732 );
and ( n35117 , n35113 , n35116 );
and ( n35118 , n35111 , n35116 );
or ( n35119 , n35114 , n35117 , n35118 );
xor ( n35120 , n34818 , n34819 );
xor ( n35121 , n35120 , n34821 );
xor ( n35122 , n34825 , n34826 );
xor ( n35123 , n35122 , n34828 );
and ( n35124 , n35121 , n35123 );
xor ( n35125 , n34757 , n34758 );
xor ( n35126 , n35125 , n34760 );
and ( n35127 , n35123 , n35126 );
and ( n35128 , n35121 , n35126 );
or ( n35129 , n35124 , n35127 , n35128 );
and ( n35130 , n35119 , n35129 );
and ( n35131 , n35109 , n35130 );
xor ( n35132 , n34764 , n34765 );
xor ( n35133 , n35132 , n34767 );
xor ( n35134 , n34772 , n34773 );
xor ( n35135 , n35134 , n34775 );
or ( n35136 , n35133 , n35135 );
xor ( n35137 , n34736 , n34737 );
xor ( n35138 , n35137 , n34739 );
xor ( n35139 , n34744 , n34745 );
xor ( n35140 , n35139 , n34747 );
or ( n35141 , n35138 , n35140 );
and ( n35142 , n35136 , n35141 );
and ( n35143 , n35130 , n35142 );
and ( n35144 , n35109 , n35142 );
or ( n35145 , n35131 , n35143 , n35144 );
xor ( n35146 , n34796 , n34797 );
xor ( n35147 , n35146 , n34799 );
and ( n35148 , n35145 , n35147 );
xor ( n35149 , n34817 , n34848 );
xor ( n35150 , n35149 , n34860 );
and ( n35151 , n35147 , n35150 );
and ( n35152 , n35145 , n35150 );
or ( n35153 , n35148 , n35151 , n35152 );
and ( n35154 , n35107 , n35153 );
and ( n35155 , n35084 , n35153 );
or ( n35156 , n35108 , n35154 , n35155 );
xor ( n35157 , n34726 , n34727 );
xor ( n35158 , n35157 , n34785 );
xor ( n35159 , n34791 , n34794 );
xor ( n35160 , n35159 , n34802 );
and ( n35161 , n35158 , n35160 );
xor ( n35162 , n34863 , n34880 );
xor ( n35163 , n35162 , n34883 );
and ( n35164 , n35160 , n35163 );
and ( n35165 , n35158 , n35163 );
or ( n35166 , n35161 , n35164 , n35165 );
and ( n35167 , n35156 , n35166 );
xor ( n35168 , n34665 , n34667 );
xor ( n35169 , n35168 , n34721 );
and ( n35170 , n35166 , n35169 );
and ( n35171 , n35156 , n35169 );
or ( n35172 , n35167 , n35170 , n35171 );
and ( n35173 , n35014 , n35172 );
and ( n35174 , n34947 , n35172 );
or ( n35175 , n35015 , n35173 , n35174 );
and ( n35176 , n34945 , n35175 );
xor ( n35177 , n34892 , n34918 );
xor ( n35178 , n35177 , n34921 );
and ( n35179 , n35175 , n35178 );
and ( n35180 , n34945 , n35178 );
or ( n35181 , n35176 , n35179 , n35180 );
xor ( n35182 , n34924 , n34926 );
xor ( n35183 , n35182 , n34929 );
and ( n35184 , n35181 , n35183 );
xor ( n35185 , n34663 , n34724 );
xor ( n35186 , n35185 , n34889 );
xor ( n35187 , n34910 , n34912 );
xor ( n35188 , n35187 , n34915 );
and ( n35189 , n35186 , n35188 );
xor ( n35190 , n34788 , n34805 );
xor ( n35191 , n35190 , n34886 );
xor ( n35192 , n34902 , n34904 );
xor ( n35193 , n35192 , n34907 );
and ( n35194 , n35191 , n35193 );
xor ( n35195 , n34894 , n34896 );
xor ( n35196 , n35195 , n34899 );
xor ( n35197 , n34868 , n34873 );
xor ( n35198 , n35197 , n34877 );
xnor ( n35199 , n35017 , n35018 );
xnor ( n35200 , n35020 , n35021 );
and ( n35201 , n35199 , n35200 );
not ( n35202 , n35201 );
buf ( n35203 , n15865 );
buf ( n35204 , n35203 );
and ( n35205 , n35202 , n35204 );
and ( n35206 , n35198 , n35205 );
buf ( n35207 , n35201 );
and ( n35208 , n35205 , n35207 );
and ( n35209 , n35198 , n35207 );
or ( n35210 , n35206 , n35208 , n35209 );
and ( n35211 , n35196 , n35210 );
xnor ( n35212 , n34808 , n34810 );
xnor ( n35213 , n34813 , n34815 );
and ( n35214 , n35212 , n35213 );
xor ( n35215 , n34954 , n34958 );
xor ( n35216 , n35215 , n34960 );
and ( n35217 , n35214 , n35216 );
xor ( n35218 , n35001 , n35004 );
and ( n35219 , n35216 , n35218 );
and ( n35220 , n35214 , n35218 );
or ( n35221 , n35217 , n35219 , n35220 );
xor ( n35222 , n35019 , n35022 );
xor ( n35223 , n35052 , n35080 );
and ( n35224 , n35222 , n35223 );
xor ( n35225 , n35085 , n35086 );
and ( n35226 , n35223 , n35225 );
and ( n35227 , n35222 , n35225 );
or ( n35228 , n35224 , n35226 , n35227 );
and ( n35229 , n35221 , n35228 );
xor ( n35230 , n34978 , n34980 );
buf ( n35231 , n31607 );
buf ( n35232 , n15874 );
buf ( n35233 , n35232 );
and ( n35234 , n35231 , n35233 );
and ( n35235 , n35230 , n35234 );
and ( n35236 , n30464 , n34253 );
and ( n35237 , n34280 , n30461 );
and ( n35238 , n35236 , n35237 );
and ( n35239 , n35234 , n35238 );
and ( n35240 , n35230 , n35238 );
or ( n35241 , n35235 , n35239 , n35240 );
xnor ( n35242 , n35133 , n35135 );
xnor ( n35243 , n35138 , n35140 );
and ( n35244 , n35242 , n35243 );
or ( n35245 , n35241 , n35244 );
and ( n35246 , n34280 , n30473 );
and ( n35247 , n32736 , n30898 );
and ( n35248 , n35246 , n35247 );
and ( n35249 , n32057 , n31301 );
and ( n35250 , n35247 , n35249 );
and ( n35251 , n35246 , n35249 );
or ( n35252 , n35248 , n35250 , n35251 );
and ( n35253 , n33339 , n30791 );
and ( n35254 , n32949 , n30788 );
and ( n35255 , n35253 , n35254 );
and ( n35256 , n32155 , n31247 );
and ( n35257 , n35254 , n35256 );
and ( n35258 , n35253 , n35256 );
or ( n35259 , n35255 , n35257 , n35258 );
and ( n35260 , n35252 , n35259 );
and ( n35261 , n32689 , n31076 );
and ( n35262 , n31883 , n31442 );
and ( n35263 , n35261 , n35262 );
and ( n35264 , n31736 , n31590 );
and ( n35265 , n35262 , n35264 );
and ( n35266 , n35261 , n35264 );
or ( n35267 , n35263 , n35265 , n35266 );
and ( n35268 , n35259 , n35267 );
and ( n35269 , n35252 , n35267 );
or ( n35270 , n35260 , n35268 , n35269 );
xor ( n35271 , n35031 , n35038 );
xor ( n35272 , n35271 , n35046 );
or ( n35273 , n35270 , n35272 );
and ( n35274 , n30468 , n34253 );
and ( n35275 , n30889 , n32719 );
and ( n35276 , n35274 , n35275 );
and ( n35277 , n31278 , n32066 );
and ( n35278 , n35275 , n35277 );
and ( n35279 , n35274 , n35277 );
or ( n35280 , n35276 , n35278 , n35279 );
and ( n35281 , n30799 , n33296 );
and ( n35282 , n30803 , n32932 );
and ( n35283 , n35281 , n35282 );
and ( n35284 , n31238 , n32173 );
and ( n35285 , n35282 , n35284 );
and ( n35286 , n35281 , n35284 );
or ( n35287 , n35283 , n35285 , n35286 );
and ( n35288 , n35280 , n35287 );
and ( n35289 , n31084 , n32671 );
and ( n35290 , n31464 , n31861 );
and ( n35291 , n35289 , n35290 );
and ( n35292 , n31607 , n31745 );
and ( n35293 , n35290 , n35292 );
and ( n35294 , n35289 , n35292 );
or ( n35295 , n35291 , n35293 , n35294 );
and ( n35296 , n35287 , n35295 );
and ( n35297 , n35280 , n35295 );
or ( n35298 , n35288 , n35296 , n35297 );
xor ( n35299 , n35059 , n35066 );
xor ( n35300 , n35299 , n35074 );
or ( n35301 , n35298 , n35300 );
and ( n35302 , n35273 , n35301 );
and ( n35303 , n35245 , n35302 );
xnor ( n35304 , n35049 , n35051 );
xnor ( n35305 , n35077 , n35079 );
and ( n35306 , n35304 , n35305 );
and ( n35307 , n35302 , n35306 );
and ( n35308 , n35245 , n35306 );
or ( n35309 , n35303 , n35307 , n35308 );
and ( n35310 , n35228 , n35309 );
and ( n35311 , n35221 , n35309 );
or ( n35312 , n35229 , n35310 , n35311 );
and ( n35313 , n35210 , n35312 );
and ( n35314 , n35196 , n35312 );
or ( n35315 , n35211 , n35313 , n35314 );
and ( n35316 , n35193 , n35315 );
and ( n35317 , n35191 , n35315 );
or ( n35318 , n35194 , n35316 , n35317 );
and ( n35319 , n35188 , n35318 );
and ( n35320 , n35186 , n35318 );
or ( n35321 , n35189 , n35319 , n35320 );
xor ( n35322 , n34945 , n35175 );
xor ( n35323 , n35322 , n35178 );
and ( n35324 , n35321 , n35323 );
xor ( n35325 , n35088 , n35089 );
xor ( n35326 , n34975 , n34981 );
xor ( n35327 , n35326 , n34997 );
and ( n35328 , n35325 , n35327 );
xor ( n35329 , n35119 , n35129 );
and ( n35330 , n35327 , n35329 );
and ( n35331 , n35325 , n35329 );
or ( n35332 , n35328 , n35330 , n35331 );
xor ( n35333 , n35136 , n35141 );
xor ( n35334 , n35212 , n35213 );
and ( n35335 , n35333 , n35334 );
xor ( n35336 , n35002 , n35003 );
and ( n35337 , n35334 , n35336 );
and ( n35338 , n35333 , n35336 );
or ( n35339 , n35335 , n35337 , n35338 );
and ( n35340 , n35332 , n35339 );
and ( n35341 , n30603 , n33712 );
and ( n35342 , n30709 , n33347 );
and ( n35343 , n35341 , n35342 );
and ( n35344 , n31088 , n32348 );
and ( n35345 , n35342 , n35344 );
and ( n35346 , n35341 , n35344 );
or ( n35347 , n35343 , n35345 , n35346 );
xor ( n35348 , n35025 , n35026 );
xor ( n35349 , n35348 , n35028 );
and ( n35350 , n35347 , n35349 );
xor ( n35351 , n34983 , n34984 );
xor ( n35352 , n35351 , n34986 );
and ( n35353 , n35349 , n35352 );
and ( n35354 , n35347 , n35352 );
or ( n35355 , n35350 , n35353 , n35354 );
and ( n35356 , n33692 , n30592 );
and ( n35357 , n33304 , n30700 );
and ( n35358 , n35356 , n35357 );
and ( n35359 , n32365 , n31073 );
and ( n35360 , n35357 , n35359 );
and ( n35361 , n35356 , n35359 );
or ( n35362 , n35358 , n35360 , n35361 );
xor ( n35363 , n35053 , n35054 );
xor ( n35364 , n35363 , n35056 );
and ( n35365 , n35362 , n35364 );
xor ( n35366 , n34990 , n34991 );
xor ( n35367 , n35366 , n34993 );
and ( n35368 , n35364 , n35367 );
and ( n35369 , n35362 , n35367 );
or ( n35370 , n35365 , n35368 , n35369 );
and ( n35371 , n35355 , n35370 );
xor ( n35372 , n35060 , n35061 );
xor ( n35373 , n35372 , n35063 );
xor ( n35374 , n35068 , n35069 );
xor ( n35375 , n35374 , n35071 );
or ( n35376 , n35373 , n35375 );
xor ( n35377 , n35032 , n35033 );
xor ( n35378 , n35377 , n35035 );
xor ( n35379 , n35040 , n35041 );
xor ( n35380 , n35379 , n35043 );
or ( n35381 , n35378 , n35380 );
and ( n35382 , n35376 , n35381 );
and ( n35383 , n35371 , n35382 );
xor ( n35384 , n35111 , n35113 );
xor ( n35385 , n35384 , n35116 );
xor ( n35386 , n35121 , n35123 );
xor ( n35387 , n35386 , n35126 );
and ( n35388 , n35385 , n35387 );
and ( n35389 , n35382 , n35388 );
and ( n35390 , n35371 , n35388 );
or ( n35391 , n35383 , n35389 , n35390 );
and ( n35392 , n35339 , n35391 );
and ( n35393 , n35332 , n35391 );
or ( n35394 , n35340 , n35392 , n35393 );
xor ( n35395 , n35090 , n35091 );
xor ( n35396 , n35395 , n35093 );
xor ( n35397 , n35098 , n35099 );
xor ( n35398 , n35397 , n35101 );
and ( n35399 , n35396 , n35398 );
xor ( n35400 , n35109 , n35130 );
xor ( n35401 , n35400 , n35142 );
and ( n35402 , n35398 , n35401 );
and ( n35403 , n35396 , n35401 );
or ( n35404 , n35399 , n35402 , n35403 );
and ( n35405 , n35394 , n35404 );
xor ( n35406 , n34963 , n34965 );
xor ( n35407 , n35406 , n34967 );
and ( n35408 , n35404 , n35407 );
and ( n35409 , n35394 , n35407 );
or ( n35410 , n35405 , n35408 , n35409 );
xor ( n35411 , n34972 , n34973 );
xor ( n35412 , n35411 , n35005 );
xor ( n35413 , n35016 , n35023 );
xor ( n35414 , n35413 , n35081 );
and ( n35415 , n35412 , n35414 );
xor ( n35416 , n35087 , n35096 );
xor ( n35417 , n35416 , n35104 );
and ( n35418 , n35414 , n35417 );
and ( n35419 , n35412 , n35417 );
or ( n35420 , n35415 , n35418 , n35419 );
and ( n35421 , n35410 , n35420 );
xor ( n35422 , n34953 , n34970 );
xor ( n35423 , n35422 , n35008 );
and ( n35424 , n35420 , n35423 );
and ( n35425 , n35410 , n35423 );
or ( n35426 , n35421 , n35424 , n35425 );
xor ( n35427 , n34949 , n34951 );
xor ( n35428 , n35427 , n35011 );
and ( n35429 , n35426 , n35428 );
xor ( n35430 , n35156 , n35166 );
xor ( n35431 , n35430 , n35169 );
and ( n35432 , n35428 , n35431 );
and ( n35433 , n35426 , n35431 );
or ( n35434 , n35429 , n35432 , n35433 );
xor ( n35435 , n34947 , n35014 );
xor ( n35436 , n35435 , n35172 );
and ( n35437 , n35434 , n35436 );
xor ( n35438 , n35084 , n35107 );
xor ( n35439 , n35438 , n35153 );
xor ( n35440 , n35158 , n35160 );
xor ( n35441 , n35440 , n35163 );
and ( n35442 , n35439 , n35441 );
xor ( n35443 , n35145 , n35147 );
xor ( n35444 , n35443 , n35150 );
xor ( n35445 , n35202 , n35204 );
xor ( n35446 , n34989 , n34996 );
and ( n35447 , n34099 , n30508 );
and ( n35448 , n33896 , n30563 );
or ( n35449 , n35447 , n35448 );
and ( n35450 , n30503 , n34082 );
and ( n35451 , n30558 , n33905 );
or ( n35452 , n35450 , n35451 );
and ( n35453 , n35449 , n35452 );
and ( n35454 , n35446 , n35453 );
xor ( n35455 , n35231 , n35233 );
xor ( n35456 , n35236 , n35237 );
and ( n35457 , n35455 , n35456 );
xor ( n35458 , n34976 , n34977 );
and ( n35459 , n35456 , n35458 );
and ( n35460 , n35455 , n35458 );
or ( n35461 , n35457 , n35459 , n35460 );
and ( n35462 , n35453 , n35461 );
and ( n35463 , n35446 , n35461 );
or ( n35464 , n35454 , n35462 , n35463 );
xnor ( n35465 , n35241 , n35244 );
and ( n35466 , n35464 , n35465 );
xor ( n35467 , n35273 , n35301 );
and ( n35468 , n35465 , n35467 );
and ( n35469 , n35464 , n35467 );
or ( n35470 , n35466 , n35468 , n35469 );
and ( n35471 , n35445 , n35470 );
xor ( n35472 , n35199 , n35200 );
xor ( n35473 , n35304 , n35305 );
and ( n35474 , n35472 , n35473 );
xnor ( n35475 , n35270 , n35272 );
xnor ( n35476 , n35298 , n35300 );
and ( n35477 , n35475 , n35476 );
and ( n35478 , n35473 , n35477 );
and ( n35479 , n35472 , n35477 );
or ( n35480 , n35474 , n35478 , n35479 );
and ( n35481 , n35470 , n35480 );
and ( n35482 , n35445 , n35480 );
or ( n35483 , n35471 , n35481 , n35482 );
and ( n35484 , n35444 , n35483 );
xor ( n35485 , n35230 , n35234 );
xor ( n35486 , n35485 , n35238 );
xor ( n35487 , n35355 , n35370 );
and ( n35488 , n35486 , n35487 );
xor ( n35489 , n35376 , n35381 );
and ( n35490 , n35487 , n35489 );
and ( n35491 , n35486 , n35489 );
or ( n35492 , n35488 , n35490 , n35491 );
xor ( n35493 , n35385 , n35387 );
xor ( n35494 , n35242 , n35243 );
and ( n35495 , n35493 , n35494 );
xor ( n35496 , n35246 , n35247 );
xor ( n35497 , n35496 , n35249 );
xor ( n35498 , n35356 , n35357 );
xor ( n35499 , n35498 , n35359 );
and ( n35500 , n35497 , n35499 );
xor ( n35501 , n35253 , n35254 );
xor ( n35502 , n35501 , n35256 );
and ( n35503 , n35499 , n35502 );
and ( n35504 , n35497 , n35502 );
or ( n35505 , n35500 , n35503 , n35504 );
xor ( n35506 , n35274 , n35275 );
xor ( n35507 , n35506 , n35277 );
xor ( n35508 , n35341 , n35342 );
xor ( n35509 , n35508 , n35344 );
and ( n35510 , n35507 , n35509 );
xor ( n35511 , n35281 , n35282 );
xor ( n35512 , n35511 , n35284 );
and ( n35513 , n35509 , n35512 );
and ( n35514 , n35507 , n35512 );
or ( n35515 , n35510 , n35513 , n35514 );
and ( n35516 , n35505 , n35515 );
and ( n35517 , n35494 , n35516 );
and ( n35518 , n35493 , n35516 );
or ( n35519 , n35495 , n35517 , n35518 );
and ( n35520 , n35492 , n35519 );
and ( n35521 , n30803 , n33296 );
and ( n35522 , n30889 , n32932 );
and ( n35523 , n35521 , n35522 );
and ( n35524 , n31278 , n32173 );
and ( n35525 , n35522 , n35524 );
and ( n35526 , n35521 , n35524 );
or ( n35527 , n35523 , n35525 , n35526 );
and ( n35528 , n30709 , n33712 );
and ( n35529 , n30799 , n33347 );
and ( n35530 , n35528 , n35529 );
and ( n35531 , n31238 , n32348 );
and ( n35532 , n35529 , n35531 );
and ( n35533 , n35528 , n35531 );
or ( n35534 , n35530 , n35532 , n35533 );
or ( n35535 , n35527 , n35534 );
and ( n35536 , n33339 , n30788 );
and ( n35537 , n32949 , n30898 );
and ( n35538 , n35536 , n35537 );
and ( n35539 , n32155 , n31301 );
and ( n35540 , n35537 , n35539 );
and ( n35541 , n35536 , n35539 );
or ( n35542 , n35538 , n35540 , n35541 );
and ( n35543 , n33692 , n30700 );
and ( n35544 , n33304 , n30791 );
and ( n35545 , n35543 , n35544 );
and ( n35546 , n32365 , n31247 );
and ( n35547 , n35544 , n35546 );
and ( n35548 , n35543 , n35546 );
or ( n35549 , n35545 , n35547 , n35548 );
or ( n35550 , n35542 , n35549 );
and ( n35551 , n35535 , n35550 );
and ( n35552 , n30603 , n33905 );
and ( n35553 , n31088 , n32671 );
and ( n35554 , n35552 , n35553 );
and ( n35555 , n31464 , n32066 );
and ( n35556 , n35553 , n35555 );
and ( n35557 , n35552 , n35555 );
or ( n35558 , n35554 , n35556 , n35557 );
and ( n35559 , n30503 , n34253 );
and ( n35560 , n30558 , n34082 );
and ( n35561 , n35559 , n35560 );
and ( n35562 , n31084 , n32719 );
and ( n35563 , n35560 , n35562 );
and ( n35564 , n35559 , n35562 );
or ( n35565 , n35561 , n35563 , n35564 );
or ( n35566 , n35558 , n35565 );
and ( n35567 , n33896 , n30592 );
and ( n35568 , n32689 , n31073 );
and ( n35569 , n35567 , n35568 );
and ( n35570 , n32057 , n31442 );
and ( n35571 , n35568 , n35570 );
and ( n35572 , n35567 , n35570 );
or ( n35573 , n35569 , n35571 , n35572 );
and ( n35574 , n34280 , n30508 );
and ( n35575 , n34099 , n30563 );
and ( n35576 , n35574 , n35575 );
and ( n35577 , n32736 , n31076 );
and ( n35578 , n35575 , n35577 );
and ( n35579 , n35574 , n35577 );
or ( n35580 , n35576 , n35578 , n35579 );
or ( n35581 , n35573 , n35580 );
and ( n35582 , n35566 , n35581 );
and ( n35583 , n35551 , n35582 );
xor ( n35584 , n35280 , n35287 );
xor ( n35585 , n35584 , n35295 );
xor ( n35586 , n35252 , n35259 );
xor ( n35587 , n35586 , n35267 );
and ( n35588 , n35585 , n35587 );
and ( n35589 , n35582 , n35588 );
and ( n35590 , n35551 , n35588 );
or ( n35591 , n35583 , n35589 , n35590 );
and ( n35592 , n35519 , n35591 );
and ( n35593 , n35492 , n35591 );
or ( n35594 , n35520 , n35592 , n35593 );
xor ( n35595 , n35347 , n35349 );
xor ( n35596 , n35595 , n35352 );
xor ( n35597 , n35362 , n35364 );
xor ( n35598 , n35597 , n35367 );
and ( n35599 , n35596 , n35598 );
xnor ( n35600 , n35373 , n35375 );
xnor ( n35601 , n35378 , n35380 );
and ( n35602 , n35600 , n35601 );
and ( n35603 , n35599 , n35602 );
xor ( n35604 , n35449 , n35452 );
xnor ( n35605 , n35447 , n35448 );
xnor ( n35606 , n35450 , n35451 );
and ( n35607 , n35605 , n35606 );
and ( n35608 , n35604 , n35607 );
xor ( n35609 , n35455 , n35456 );
xor ( n35610 , n35609 , n35458 );
and ( n35611 , n35607 , n35610 );
and ( n35612 , n35604 , n35610 );
or ( n35613 , n35608 , n35611 , n35612 );
and ( n35614 , n35602 , n35613 );
and ( n35615 , n35599 , n35613 );
or ( n35616 , n35603 , n35614 , n35615 );
xor ( n35617 , n35325 , n35327 );
xor ( n35618 , n35617 , n35329 );
and ( n35619 , n35616 , n35618 );
xor ( n35620 , n35333 , n35334 );
xor ( n35621 , n35620 , n35336 );
and ( n35622 , n35618 , n35621 );
and ( n35623 , n35616 , n35621 );
or ( n35624 , n35619 , n35622 , n35623 );
and ( n35625 , n35594 , n35624 );
xor ( n35626 , n35214 , n35216 );
xor ( n35627 , n35626 , n35218 );
and ( n35628 , n35624 , n35627 );
and ( n35629 , n35594 , n35627 );
or ( n35630 , n35625 , n35628 , n35629 );
and ( n35631 , n35483 , n35630 );
and ( n35632 , n35444 , n35630 );
or ( n35633 , n35484 , n35631 , n35632 );
and ( n35634 , n35441 , n35633 );
and ( n35635 , n35439 , n35633 );
or ( n35636 , n35442 , n35634 , n35635 );
xor ( n35637 , n35222 , n35223 );
xor ( n35638 , n35637 , n35225 );
xor ( n35639 , n35245 , n35302 );
xor ( n35640 , n35639 , n35306 );
and ( n35641 , n35638 , n35640 );
xor ( n35642 , n35332 , n35339 );
xor ( n35643 , n35642 , n35391 );
and ( n35644 , n35640 , n35643 );
and ( n35645 , n35638 , n35643 );
or ( n35646 , n35641 , n35644 , n35645 );
xor ( n35647 , n35198 , n35205 );
xor ( n35648 , n35647 , n35207 );
and ( n35649 , n35646 , n35648 );
xor ( n35650 , n35221 , n35228 );
xor ( n35651 , n35650 , n35309 );
and ( n35652 , n35648 , n35651 );
and ( n35653 , n35646 , n35651 );
or ( n35654 , n35649 , n35652 , n35653 );
xor ( n35655 , n35196 , n35210 );
xor ( n35656 , n35655 , n35312 );
and ( n35657 , n35654 , n35656 );
xor ( n35658 , n35410 , n35420 );
xor ( n35659 , n35658 , n35423 );
and ( n35660 , n35656 , n35659 );
and ( n35661 , n35654 , n35659 );
or ( n35662 , n35657 , n35660 , n35661 );
and ( n35663 , n35636 , n35662 );
xor ( n35664 , n35191 , n35193 );
xor ( n35665 , n35664 , n35315 );
and ( n35666 , n35662 , n35665 );
and ( n35667 , n35636 , n35665 );
or ( n35668 , n35663 , n35666 , n35667 );
and ( n35669 , n35436 , n35668 );
and ( n35670 , n35434 , n35668 );
or ( n35671 , n35437 , n35669 , n35670 );
and ( n35672 , n35323 , n35671 );
and ( n35673 , n35321 , n35671 );
or ( n35674 , n35324 , n35672 , n35673 );
and ( n35675 , n35183 , n35674 );
and ( n35676 , n35181 , n35674 );
or ( n35677 , n35184 , n35675 , n35676 );
or ( n35678 , n34943 , n35677 );
and ( n35679 , n34940 , n35678 );
and ( n35680 , n34938 , n35678 );
or ( n35681 , n34941 , n35679 , n35680 );
or ( n35682 , n34659 , n35681 );
and ( n35683 , n34656 , n35682 );
and ( n35684 , n34202 , n35682 );
or ( n35685 , n34657 , n35683 , n35684 );
and ( n35686 , n34199 , n35685 );
and ( n35687 , n34197 , n35685 );
or ( n35688 , n34200 , n35686 , n35687 );
and ( n35689 , n33879 , n35688 );
and ( n35690 , n33877 , n35688 );
or ( n35691 , n33880 , n35689 , n35690 );
and ( n35692 , n33673 , n35691 );
xor ( n35693 , n33673 , n35691 );
xor ( n35694 , n33877 , n33879 );
xor ( n35695 , n35694 , n35688 );
xor ( n35696 , n34197 , n34199 );
xor ( n35697 , n35696 , n35685 );
xor ( n35698 , n34202 , n34656 );
xor ( n35699 , n35698 , n35682 );
not ( n35700 , n35699 );
xnor ( n35701 , n34659 , n35681 );
xor ( n35702 , n34938 , n34940 );
xor ( n35703 , n35702 , n35678 );
not ( n35704 , n35703 );
xnor ( n35705 , n34943 , n35677 );
xor ( n35706 , n35181 , n35183 );
xor ( n35707 , n35706 , n35674 );
xor ( n35708 , n35186 , n35188 );
xor ( n35709 , n35708 , n35318 );
xor ( n35710 , n35426 , n35428 );
xor ( n35711 , n35710 , n35431 );
xor ( n35712 , n35394 , n35404 );
xor ( n35713 , n35712 , n35407 );
xor ( n35714 , n35412 , n35414 );
xor ( n35715 , n35714 , n35417 );
and ( n35716 , n35713 , n35715 );
xor ( n35717 , n35396 , n35398 );
xor ( n35718 , n35717 , n35401 );
xor ( n35719 , n35371 , n35382 );
xor ( n35720 , n35719 , n35388 );
xor ( n35721 , n35446 , n35453 );
xor ( n35722 , n35721 , n35461 );
xor ( n35723 , n35475 , n35476 );
and ( n35724 , n35722 , n35723 );
and ( n35725 , n34099 , n30592 );
and ( n35726 , n33896 , n30700 );
and ( n35727 , n35725 , n35726 );
and ( n35728 , n32689 , n31247 );
and ( n35729 , n35726 , n35728 );
and ( n35730 , n35725 , n35728 );
or ( n35731 , n35727 , n35729 , n35730 );
and ( n35732 , n33692 , n30791 );
and ( n35733 , n33304 , n30788 );
and ( n35734 , n35732 , n35733 );
and ( n35735 , n32365 , n31301 );
and ( n35736 , n35733 , n35735 );
and ( n35737 , n35732 , n35735 );
or ( n35738 , n35734 , n35736 , n35737 );
and ( n35739 , n35731 , n35738 );
and ( n35740 , n33339 , n30898 );
and ( n35741 , n32949 , n31076 );
and ( n35742 , n35740 , n35741 );
and ( n35743 , n32155 , n31442 );
and ( n35744 , n35741 , n35743 );
and ( n35745 , n35740 , n35743 );
or ( n35746 , n35742 , n35744 , n35745 );
and ( n35747 , n35738 , n35746 );
and ( n35748 , n35731 , n35746 );
or ( n35749 , n35739 , n35747 , n35748 );
xor ( n35750 , n35289 , n35290 );
xor ( n35751 , n35750 , n35292 );
or ( n35752 , n35749 , n35751 );
and ( n35753 , n30603 , n34082 );
and ( n35754 , n30709 , n33905 );
and ( n35755 , n35753 , n35754 );
and ( n35756 , n31238 , n32671 );
and ( n35757 , n35754 , n35756 );
and ( n35758 , n35753 , n35756 );
or ( n35759 , n35755 , n35757 , n35758 );
and ( n35760 , n30799 , n33712 );
and ( n35761 , n30803 , n33347 );
and ( n35762 , n35760 , n35761 );
and ( n35763 , n31278 , n32348 );
and ( n35764 , n35761 , n35763 );
and ( n35765 , n35760 , n35763 );
or ( n35766 , n35762 , n35764 , n35765 );
and ( n35767 , n35759 , n35766 );
and ( n35768 , n30889 , n33296 );
and ( n35769 , n31084 , n32932 );
and ( n35770 , n35768 , n35769 );
and ( n35771 , n31464 , n32173 );
and ( n35772 , n35769 , n35771 );
and ( n35773 , n35768 , n35771 );
or ( n35774 , n35770 , n35772 , n35773 );
and ( n35775 , n35766 , n35774 );
and ( n35776 , n35759 , n35774 );
or ( n35777 , n35767 , n35775 , n35776 );
xor ( n35778 , n35261 , n35262 );
xor ( n35779 , n35778 , n35264 );
or ( n35780 , n35777 , n35779 );
and ( n35781 , n35752 , n35780 );
and ( n35782 , n35723 , n35781 );
and ( n35783 , n35722 , n35781 );
or ( n35784 , n35724 , n35782 , n35783 );
and ( n35785 , n35720 , n35784 );
xor ( n35786 , n35552 , n35553 );
xor ( n35787 , n35786 , n35555 );
xor ( n35788 , n35559 , n35560 );
xor ( n35789 , n35788 , n35562 );
and ( n35790 , n35787 , n35789 );
xor ( n35791 , n35521 , n35522 );
xor ( n35792 , n35791 , n35524 );
and ( n35793 , n35789 , n35792 );
and ( n35794 , n35787 , n35792 );
or ( n35795 , n35790 , n35793 , n35794 );
not ( n35796 , n35795 );
xnor ( n35797 , n35542 , n35549 );
and ( n35798 , n35796 , n35797 );
xor ( n35799 , n35567 , n35568 );
xor ( n35800 , n35799 , n35570 );
xor ( n35801 , n35574 , n35575 );
xor ( n35802 , n35801 , n35577 );
and ( n35803 , n35800 , n35802 );
xor ( n35804 , n35536 , n35537 );
xor ( n35805 , n35804 , n35539 );
and ( n35806 , n35802 , n35805 );
and ( n35807 , n35800 , n35805 );
or ( n35808 , n35803 , n35806 , n35807 );
not ( n35809 , n35808 );
xnor ( n35810 , n35527 , n35534 );
and ( n35811 , n35809 , n35810 );
and ( n35812 , n35798 , n35811 );
buf ( n35813 , n35795 );
buf ( n35814 , n35808 );
and ( n35815 , n35813 , n35814 );
and ( n35816 , n35812 , n35815 );
xor ( n35817 , n35505 , n35515 );
xor ( n35818 , n35535 , n35550 );
and ( n35819 , n35817 , n35818 );
xor ( n35820 , n35566 , n35581 );
and ( n35821 , n35818 , n35820 );
and ( n35822 , n35817 , n35820 );
or ( n35823 , n35819 , n35821 , n35822 );
and ( n35824 , n35815 , n35823 );
and ( n35825 , n35812 , n35823 );
or ( n35826 , n35816 , n35824 , n35825 );
and ( n35827 , n35784 , n35826 );
and ( n35828 , n35720 , n35826 );
or ( n35829 , n35785 , n35827 , n35828 );
and ( n35830 , n35718 , n35829 );
xor ( n35831 , n35585 , n35587 );
xor ( n35832 , n35596 , n35598 );
and ( n35833 , n35831 , n35832 );
xor ( n35834 , n35600 , n35601 );
and ( n35835 , n35832 , n35834 );
and ( n35836 , n35831 , n35834 );
or ( n35837 , n35833 , n35835 , n35836 );
xor ( n35838 , n35497 , n35499 );
xor ( n35839 , n35838 , n35502 );
xor ( n35840 , n35507 , n35509 );
xor ( n35841 , n35840 , n35512 );
and ( n35842 , n35839 , n35841 );
xnor ( n35843 , n35558 , n35565 );
xnor ( n35844 , n35573 , n35580 );
and ( n35845 , n35843 , n35844 );
and ( n35846 , n35842 , n35845 );
buf ( n35847 , n15877 );
buf ( n35848 , n35847 );
and ( n35849 , n31607 , n31861 );
and ( n35850 , n31883 , n31590 );
and ( n35851 , n35849 , n35850 );
and ( n35852 , n35848 , n35851 );
xor ( n35853 , n35605 , n35606 );
and ( n35854 , n35851 , n35853 );
and ( n35855 , n35848 , n35853 );
or ( n35856 , n35852 , n35854 , n35855 );
and ( n35857 , n35845 , n35856 );
and ( n35858 , n35842 , n35856 );
or ( n35859 , n35846 , n35857 , n35858 );
and ( n35860 , n35837 , n35859 );
xor ( n35861 , n35486 , n35487 );
xor ( n35862 , n35861 , n35489 );
and ( n35863 , n35859 , n35862 );
and ( n35864 , n35837 , n35862 );
or ( n35865 , n35860 , n35863 , n35864 );
xor ( n35866 , n35493 , n35494 );
xor ( n35867 , n35866 , n35516 );
xor ( n35868 , n35551 , n35582 );
xor ( n35869 , n35868 , n35588 );
and ( n35870 , n35867 , n35869 );
xor ( n35871 , n35599 , n35602 );
xor ( n35872 , n35871 , n35613 );
and ( n35873 , n35869 , n35872 );
and ( n35874 , n35867 , n35872 );
or ( n35875 , n35870 , n35873 , n35874 );
and ( n35876 , n35865 , n35875 );
xor ( n35877 , n35464 , n35465 );
xor ( n35878 , n35877 , n35467 );
and ( n35879 , n35875 , n35878 );
and ( n35880 , n35865 , n35878 );
or ( n35881 , n35876 , n35879 , n35880 );
and ( n35882 , n35829 , n35881 );
and ( n35883 , n35718 , n35881 );
or ( n35884 , n35830 , n35882 , n35883 );
and ( n35885 , n35715 , n35884 );
and ( n35886 , n35713 , n35884 );
or ( n35887 , n35716 , n35885 , n35886 );
xor ( n35888 , n35472 , n35473 );
xor ( n35889 , n35888 , n35477 );
xor ( n35890 , n35492 , n35519 );
xor ( n35891 , n35890 , n35591 );
and ( n35892 , n35889 , n35891 );
xor ( n35893 , n35616 , n35618 );
xor ( n35894 , n35893 , n35621 );
and ( n35895 , n35891 , n35894 );
and ( n35896 , n35889 , n35894 );
or ( n35897 , n35892 , n35895 , n35896 );
xor ( n35898 , n35445 , n35470 );
xor ( n35899 , n35898 , n35480 );
and ( n35900 , n35897 , n35899 );
xor ( n35901 , n35594 , n35624 );
xor ( n35902 , n35901 , n35627 );
and ( n35903 , n35899 , n35902 );
and ( n35904 , n35897 , n35902 );
or ( n35905 , n35900 , n35903 , n35904 );
xor ( n35906 , n35444 , n35483 );
xor ( n35907 , n35906 , n35630 );
and ( n35908 , n35905 , n35907 );
xor ( n35909 , n35646 , n35648 );
xor ( n35910 , n35909 , n35651 );
and ( n35911 , n35907 , n35910 );
and ( n35912 , n35905 , n35910 );
or ( n35913 , n35908 , n35911 , n35912 );
and ( n35914 , n35887 , n35913 );
xor ( n35915 , n35439 , n35441 );
xor ( n35916 , n35915 , n35633 );
and ( n35917 , n35913 , n35916 );
and ( n35918 , n35887 , n35916 );
or ( n35919 , n35914 , n35917 , n35918 );
and ( n35920 , n35711 , n35919 );
xor ( n35921 , n35636 , n35662 );
xor ( n35922 , n35921 , n35665 );
and ( n35923 , n35919 , n35922 );
and ( n35924 , n35711 , n35922 );
or ( n35925 , n35920 , n35923 , n35924 );
and ( n35926 , n35709 , n35925 );
xor ( n35927 , n35434 , n35436 );
xor ( n35928 , n35927 , n35668 );
and ( n35929 , n35925 , n35928 );
and ( n35930 , n35709 , n35928 );
or ( n35931 , n35926 , n35929 , n35930 );
xor ( n35932 , n35321 , n35323 );
xor ( n35933 , n35932 , n35671 );
and ( n35934 , n35931 , n35933 );
xor ( n35935 , n35654 , n35656 );
xor ( n35936 , n35935 , n35659 );
xor ( n35937 , n35638 , n35640 );
xor ( n35938 , n35937 , n35643 );
and ( n35939 , n32736 , n31073 );
and ( n35940 , n32057 , n31590 );
and ( n35941 , n35939 , n35940 );
and ( n35942 , n31883 , n31745 );
and ( n35943 , n35940 , n35942 );
and ( n35944 , n35939 , n35942 );
or ( n35945 , n35941 , n35943 , n35944 );
and ( n35946 , n31088 , n32719 );
and ( n35947 , n31607 , n32066 );
and ( n35948 , n35946 , n35947 );
and ( n35949 , n31736 , n31861 );
and ( n35950 , n35947 , n35949 );
and ( n35951 , n35946 , n35949 );
or ( n35952 , n35948 , n35950 , n35951 );
and ( n35953 , n35945 , n35952 );
xor ( n35954 , n35543 , n35544 );
xor ( n35955 , n35954 , n35546 );
xor ( n35956 , n35528 , n35529 );
xor ( n35957 , n35956 , n35531 );
and ( n35958 , n35955 , n35957 );
and ( n35959 , n35953 , n35958 );
buf ( n35960 , n31736 );
buf ( n35961 , n15880 );
buf ( n35962 , n35961 );
and ( n35963 , n35960 , n35962 );
xor ( n35964 , n35849 , n35850 );
and ( n35965 , n35962 , n35964 );
and ( n35966 , n35960 , n35964 );
or ( n35967 , n35963 , n35965 , n35966 );
and ( n35968 , n35958 , n35967 );
and ( n35969 , n35953 , n35967 );
or ( n35970 , n35959 , n35968 , n35969 );
xor ( n35971 , n35604 , n35607 );
xor ( n35972 , n35971 , n35610 );
and ( n35973 , n35970 , n35972 );
xor ( n35974 , n35752 , n35780 );
and ( n35975 , n35972 , n35974 );
and ( n35976 , n35970 , n35974 );
or ( n35977 , n35973 , n35975 , n35976 );
xor ( n35978 , n35798 , n35811 );
xor ( n35979 , n35813 , n35814 );
and ( n35980 , n35978 , n35979 );
and ( n35981 , n34099 , n30700 );
and ( n35982 , n32736 , n31247 );
and ( n35983 , n35981 , n35982 );
and ( n35984 , n32155 , n31590 );
and ( n35985 , n35982 , n35984 );
and ( n35986 , n35981 , n35984 );
or ( n35987 , n35983 , n35985 , n35986 );
and ( n35988 , n33304 , n30898 );
and ( n35989 , n33339 , n31076 );
and ( n35990 , n35988 , n35989 );
and ( n35991 , n32365 , n31442 );
and ( n35992 , n35989 , n35991 );
and ( n35993 , n35988 , n35991 );
or ( n35994 , n35990 , n35992 , n35993 );
and ( n35995 , n35987 , n35994 );
and ( n35996 , n33896 , n30791 );
and ( n35997 , n33692 , n30788 );
and ( n35998 , n35996 , n35997 );
and ( n35999 , n32689 , n31301 );
and ( n36000 , n35997 , n35999 );
and ( n36001 , n35996 , n35999 );
or ( n36002 , n35998 , n36000 , n36001 );
and ( n36003 , n35994 , n36002 );
and ( n36004 , n35987 , n36002 );
or ( n36005 , n35995 , n36003 , n36004 );
xor ( n36006 , n35731 , n35738 );
xor ( n36007 , n36006 , n35746 );
and ( n36008 , n36005 , n36007 );
and ( n36009 , n30709 , n34082 );
and ( n36010 , n31238 , n32719 );
and ( n36011 , n36009 , n36010 );
and ( n36012 , n31607 , n32173 );
and ( n36013 , n36010 , n36012 );
and ( n36014 , n36009 , n36012 );
or ( n36015 , n36011 , n36013 , n36014 );
and ( n36016 , n30889 , n33347 );
and ( n36017 , n31084 , n33296 );
and ( n36018 , n36016 , n36017 );
and ( n36019 , n31464 , n32348 );
and ( n36020 , n36017 , n36019 );
and ( n36021 , n36016 , n36019 );
or ( n36022 , n36018 , n36020 , n36021 );
and ( n36023 , n36015 , n36022 );
and ( n36024 , n30799 , n33905 );
and ( n36025 , n30803 , n33712 );
and ( n36026 , n36024 , n36025 );
and ( n36027 , n31278 , n32671 );
and ( n36028 , n36025 , n36027 );
and ( n36029 , n36024 , n36027 );
or ( n36030 , n36026 , n36028 , n36029 );
and ( n36031 , n36022 , n36030 );
and ( n36032 , n36015 , n36030 );
or ( n36033 , n36023 , n36031 , n36032 );
xor ( n36034 , n35759 , n35766 );
xor ( n36035 , n36034 , n35774 );
and ( n36036 , n36033 , n36035 );
and ( n36037 , n36008 , n36036 );
and ( n36038 , n35979 , n36037 );
and ( n36039 , n35978 , n36037 );
or ( n36040 , n35980 , n36038 , n36039 );
and ( n36041 , n35977 , n36040 );
xnor ( n36042 , n35749 , n35751 );
xnor ( n36043 , n35777 , n35779 );
and ( n36044 , n36042 , n36043 );
xor ( n36045 , n35796 , n35797 );
xor ( n36046 , n35809 , n35810 );
and ( n36047 , n36045 , n36046 );
and ( n36048 , n36044 , n36047 );
xor ( n36049 , n35839 , n35841 );
xor ( n36050 , n35843 , n35844 );
and ( n36051 , n36049 , n36050 );
xor ( n36052 , n35753 , n35754 );
xor ( n36053 , n36052 , n35756 );
xor ( n36054 , n35760 , n35761 );
xor ( n36055 , n36054 , n35763 );
and ( n36056 , n36053 , n36055 );
xor ( n36057 , n35725 , n35726 );
xor ( n36058 , n36057 , n35728 );
xor ( n36059 , n35732 , n35733 );
xor ( n36060 , n36059 , n35735 );
and ( n36061 , n36058 , n36060 );
and ( n36062 , n36056 , n36061 );
and ( n36063 , n36050 , n36062 );
and ( n36064 , n36049 , n36062 );
or ( n36065 , n36051 , n36063 , n36064 );
and ( n36066 , n36047 , n36065 );
and ( n36067 , n36044 , n36065 );
or ( n36068 , n36048 , n36066 , n36067 );
and ( n36069 , n36040 , n36068 );
and ( n36070 , n35977 , n36068 );
or ( n36071 , n36041 , n36069 , n36070 );
xor ( n36072 , n35946 , n35947 );
xor ( n36073 , n36072 , n35949 );
xor ( n36074 , n35768 , n35769 );
xor ( n36075 , n36074 , n35771 );
and ( n36076 , n36073 , n36075 );
xor ( n36077 , n35939 , n35940 );
xor ( n36078 , n36077 , n35942 );
xor ( n36079 , n35740 , n35741 );
xor ( n36080 , n36079 , n35743 );
and ( n36081 , n36078 , n36080 );
and ( n36082 , n36076 , n36081 );
xor ( n36083 , n35800 , n35802 );
xor ( n36084 , n36083 , n35805 );
xor ( n36085 , n35787 , n35789 );
xor ( n36086 , n36085 , n35792 );
and ( n36087 , n36084 , n36086 );
and ( n36088 , n36082 , n36087 );
and ( n36089 , n30558 , n34253 );
and ( n36090 , n34280 , n30563 );
and ( n36091 , n36089 , n36090 );
xor ( n36092 , n35945 , n35952 );
and ( n36093 , n36091 , n36092 );
xor ( n36094 , n35955 , n35957 );
and ( n36095 , n36092 , n36094 );
and ( n36096 , n36091 , n36094 );
or ( n36097 , n36093 , n36095 , n36096 );
and ( n36098 , n36087 , n36097 );
and ( n36099 , n36082 , n36097 );
or ( n36100 , n36088 , n36098 , n36099 );
and ( n36101 , n31736 , n32066 );
and ( n36102 , n32057 , n31745 );
and ( n36103 , n36101 , n36102 );
buf ( n36104 , n15883 );
buf ( n36105 , n36104 );
and ( n36106 , n36103 , n36105 );
and ( n36107 , n34280 , n30592 );
and ( n36108 , n32949 , n31073 );
or ( n36109 , n36107 , n36108 );
and ( n36110 , n30603 , n34253 );
and ( n36111 , n31088 , n32932 );
or ( n36112 , n36110 , n36111 );
and ( n36113 , n36109 , n36112 );
and ( n36114 , n36106 , n36113 );
xor ( n36115 , n35960 , n35962 );
xor ( n36116 , n36115 , n35964 );
and ( n36117 , n36113 , n36116 );
and ( n36118 , n36106 , n36116 );
or ( n36119 , n36114 , n36117 , n36118 );
xor ( n36120 , n35848 , n35851 );
xor ( n36121 , n36120 , n35853 );
and ( n36122 , n36119 , n36121 );
xor ( n36123 , n35953 , n35958 );
xor ( n36124 , n36123 , n35967 );
and ( n36125 , n36121 , n36124 );
and ( n36126 , n36119 , n36124 );
or ( n36127 , n36122 , n36125 , n36126 );
and ( n36128 , n36100 , n36127 );
xor ( n36129 , n35817 , n35818 );
xor ( n36130 , n36129 , n35820 );
and ( n36131 , n36127 , n36130 );
and ( n36132 , n36100 , n36130 );
or ( n36133 , n36128 , n36131 , n36132 );
xor ( n36134 , n35722 , n35723 );
xor ( n36135 , n36134 , n35781 );
and ( n36136 , n36133 , n36135 );
xor ( n36137 , n35812 , n35815 );
xor ( n36138 , n36137 , n35823 );
and ( n36139 , n36135 , n36138 );
and ( n36140 , n36133 , n36138 );
or ( n36141 , n36136 , n36139 , n36140 );
and ( n36142 , n36071 , n36141 );
xor ( n36143 , n35720 , n35784 );
xor ( n36144 , n36143 , n35826 );
and ( n36145 , n36141 , n36144 );
and ( n36146 , n36071 , n36144 );
or ( n36147 , n36142 , n36145 , n36146 );
and ( n36148 , n35938 , n36147 );
xor ( n36149 , n35718 , n35829 );
xor ( n36150 , n36149 , n35881 );
and ( n36151 , n36147 , n36150 );
and ( n36152 , n35938 , n36150 );
or ( n36153 , n36148 , n36151 , n36152 );
xor ( n36154 , n35713 , n35715 );
xor ( n36155 , n36154 , n35884 );
and ( n36156 , n36153 , n36155 );
xor ( n36157 , n35905 , n35907 );
xor ( n36158 , n36157 , n35910 );
and ( n36159 , n36155 , n36158 );
and ( n36160 , n36153 , n36158 );
or ( n36161 , n36156 , n36159 , n36160 );
and ( n36162 , n35936 , n36161 );
xor ( n36163 , n35887 , n35913 );
xor ( n36164 , n36163 , n35916 );
and ( n36165 , n36161 , n36164 );
and ( n36166 , n35936 , n36164 );
or ( n36167 , n36162 , n36165 , n36166 );
xor ( n36168 , n35711 , n35919 );
xor ( n36169 , n36168 , n35922 );
or ( n36170 , n36167 , n36169 );
xor ( n36171 , n35709 , n35925 );
xor ( n36172 , n36171 , n35928 );
or ( n36173 , n36170 , n36172 );
and ( n36174 , n35933 , n36173 );
and ( n36175 , n35931 , n36173 );
or ( n36176 , n35934 , n36174 , n36175 );
and ( n36177 , n35707 , n36176 );
xor ( n36178 , n35707 , n36176 );
xor ( n36179 , n35931 , n35933 );
xor ( n36180 , n36179 , n36173 );
xnor ( n36181 , n36170 , n36172 );
xnor ( n36182 , n36167 , n36169 );
xor ( n36183 , n35936 , n36161 );
xor ( n36184 , n36183 , n36164 );
xor ( n36185 , n35897 , n35899 );
xor ( n36186 , n36185 , n35902 );
xor ( n36187 , n35865 , n35875 );
xor ( n36188 , n36187 , n35878 );
xor ( n36189 , n35889 , n35891 );
xor ( n36190 , n36189 , n35894 );
and ( n36191 , n36188 , n36190 );
xor ( n36192 , n35837 , n35859 );
xor ( n36193 , n36192 , n35862 );
xor ( n36194 , n35867 , n35869 );
xor ( n36195 , n36194 , n35872 );
and ( n36196 , n36193 , n36195 );
xor ( n36197 , n35831 , n35832 );
xor ( n36198 , n36197 , n35834 );
xor ( n36199 , n35842 , n35845 );
xor ( n36200 , n36199 , n35856 );
and ( n36201 , n36198 , n36200 );
xor ( n36202 , n36008 , n36036 );
xor ( n36203 , n36042 , n36043 );
and ( n36204 , n36202 , n36203 );
xor ( n36205 , n36045 , n36046 );
and ( n36206 , n36203 , n36205 );
and ( n36207 , n36202 , n36205 );
or ( n36208 , n36204 , n36206 , n36207 );
and ( n36209 , n36200 , n36208 );
and ( n36210 , n36198 , n36208 );
or ( n36211 , n36201 , n36209 , n36210 );
and ( n36212 , n36195 , n36211 );
and ( n36213 , n36193 , n36211 );
or ( n36214 , n36196 , n36212 , n36213 );
and ( n36215 , n36190 , n36214 );
and ( n36216 , n36188 , n36214 );
or ( n36217 , n36191 , n36215 , n36216 );
and ( n36218 , n36186 , n36217 );
xor ( n36219 , n35938 , n36147 );
xor ( n36220 , n36219 , n36150 );
and ( n36221 , n36217 , n36220 );
and ( n36222 , n36186 , n36220 );
or ( n36223 , n36218 , n36221 , n36222 );
xor ( n36224 , n36153 , n36155 );
xor ( n36225 , n36224 , n36158 );
and ( n36226 , n36223 , n36225 );
xor ( n36227 , n36005 , n36007 );
xor ( n36228 , n36033 , n36035 );
and ( n36229 , n36227 , n36228 );
xor ( n36230 , n36056 , n36061 );
xor ( n36231 , n36076 , n36081 );
and ( n36232 , n36230 , n36231 );
xor ( n36233 , n36084 , n36086 );
and ( n36234 , n36231 , n36233 );
and ( n36235 , n36230 , n36233 );
or ( n36236 , n36232 , n36234 , n36235 );
and ( n36237 , n36229 , n36236 );
xor ( n36238 , n35981 , n35982 );
xor ( n36239 , n36238 , n35984 );
xor ( n36240 , n35988 , n35989 );
xor ( n36241 , n36240 , n35991 );
and ( n36242 , n36239 , n36241 );
xor ( n36243 , n35996 , n35997 );
xor ( n36244 , n36243 , n35999 );
and ( n36245 , n36241 , n36244 );
and ( n36246 , n36239 , n36244 );
or ( n36247 , n36242 , n36245 , n36246 );
xor ( n36248 , n36009 , n36010 );
xor ( n36249 , n36248 , n36012 );
xor ( n36250 , n36016 , n36017 );
xor ( n36251 , n36250 , n36019 );
and ( n36252 , n36249 , n36251 );
xor ( n36253 , n36024 , n36025 );
xor ( n36254 , n36253 , n36027 );
and ( n36255 , n36251 , n36254 );
and ( n36256 , n36249 , n36254 );
or ( n36257 , n36252 , n36255 , n36256 );
and ( n36258 , n36247 , n36257 );
and ( n36259 , n31238 , n32932 );
and ( n36260 , n31736 , n32173 );
and ( n36261 , n36259 , n36260 );
and ( n36262 , n31883 , n32066 );
and ( n36263 , n36260 , n36262 );
and ( n36264 , n36259 , n36262 );
or ( n36265 , n36261 , n36263 , n36264 );
and ( n36266 , n30709 , n34253 );
and ( n36267 , n30799 , n34082 );
and ( n36268 , n36266 , n36267 );
and ( n36269 , n31278 , n32719 );
and ( n36270 , n36267 , n36269 );
and ( n36271 , n36266 , n36269 );
or ( n36272 , n36268 , n36270 , n36271 );
or ( n36273 , n36265 , n36272 );
and ( n36274 , n32949 , n31247 );
and ( n36275 , n32155 , n31745 );
and ( n36276 , n36274 , n36275 );
and ( n36277 , n32057 , n31861 );
and ( n36278 , n36275 , n36277 );
and ( n36279 , n36274 , n36277 );
or ( n36280 , n36276 , n36278 , n36279 );
and ( n36281 , n34280 , n30700 );
and ( n36282 , n34099 , n30791 );
and ( n36283 , n36281 , n36282 );
and ( n36284 , n32736 , n31301 );
and ( n36285 , n36282 , n36284 );
and ( n36286 , n36281 , n36284 );
or ( n36287 , n36283 , n36285 , n36286 );
or ( n36288 , n36280 , n36287 );
and ( n36289 , n36273 , n36288 );
and ( n36290 , n36258 , n36289 );
and ( n36291 , n31084 , n33347 );
and ( n36292 , n31088 , n33296 );
and ( n36293 , n36291 , n36292 );
and ( n36294 , n31607 , n32348 );
and ( n36295 , n36292 , n36294 );
and ( n36296 , n36291 , n36294 );
or ( n36297 , n36293 , n36295 , n36296 );
and ( n36298 , n30803 , n33905 );
and ( n36299 , n30889 , n33712 );
and ( n36300 , n36298 , n36299 );
and ( n36301 , n31464 , n32671 );
and ( n36302 , n36299 , n36301 );
and ( n36303 , n36298 , n36301 );
or ( n36304 , n36300 , n36302 , n36303 );
and ( n36305 , n36297 , n36304 );
and ( n36306 , n33304 , n31076 );
and ( n36307 , n33339 , n31073 );
and ( n36308 , n36306 , n36307 );
and ( n36309 , n32365 , n31590 );
and ( n36310 , n36307 , n36309 );
and ( n36311 , n36306 , n36309 );
or ( n36312 , n36308 , n36310 , n36311 );
and ( n36313 , n33896 , n30788 );
and ( n36314 , n33692 , n30898 );
and ( n36315 , n36313 , n36314 );
and ( n36316 , n32689 , n31442 );
and ( n36317 , n36314 , n36316 );
and ( n36318 , n36313 , n36316 );
or ( n36319 , n36315 , n36317 , n36318 );
and ( n36320 , n36312 , n36319 );
and ( n36321 , n36305 , n36320 );
and ( n36322 , n36289 , n36321 );
and ( n36323 , n36258 , n36321 );
or ( n36324 , n36290 , n36322 , n36323 );
and ( n36325 , n36236 , n36324 );
and ( n36326 , n36229 , n36324 );
or ( n36327 , n36237 , n36325 , n36326 );
xor ( n36328 , n36015 , n36022 );
xor ( n36329 , n36328 , n36030 );
xor ( n36330 , n35987 , n35994 );
xor ( n36331 , n36330 , n36002 );
and ( n36332 , n36329 , n36331 );
xor ( n36333 , n36053 , n36055 );
xor ( n36334 , n36058 , n36060 );
and ( n36335 , n36333 , n36334 );
and ( n36336 , n36332 , n36335 );
xor ( n36337 , n36073 , n36075 );
xor ( n36338 , n36078 , n36080 );
and ( n36339 , n36337 , n36338 );
and ( n36340 , n36335 , n36339 );
and ( n36341 , n36332 , n36339 );
or ( n36342 , n36336 , n36340 , n36341 );
xor ( n36343 , n36089 , n36090 );
buf ( n36344 , n31883 );
buf ( n36345 , n15886 );
buf ( n36346 , n36345 );
and ( n36347 , n36344 , n36346 );
and ( n36348 , n36343 , n36347 );
xor ( n36349 , n36109 , n36112 );
and ( n36350 , n36347 , n36349 );
and ( n36351 , n36343 , n36349 );
or ( n36352 , n36348 , n36350 , n36351 );
xor ( n36353 , n36091 , n36092 );
xor ( n36354 , n36353 , n36094 );
and ( n36355 , n36352 , n36354 );
xor ( n36356 , n36106 , n36113 );
xor ( n36357 , n36356 , n36116 );
and ( n36358 , n36354 , n36357 );
and ( n36359 , n36352 , n36357 );
or ( n36360 , n36355 , n36358 , n36359 );
and ( n36361 , n36342 , n36360 );
xor ( n36362 , n36049 , n36050 );
xor ( n36363 , n36362 , n36062 );
and ( n36364 , n36360 , n36363 );
and ( n36365 , n36342 , n36363 );
or ( n36366 , n36361 , n36364 , n36365 );
and ( n36367 , n36327 , n36366 );
xor ( n36368 , n35970 , n35972 );
xor ( n36369 , n36368 , n35974 );
and ( n36370 , n36366 , n36369 );
and ( n36371 , n36327 , n36369 );
or ( n36372 , n36367 , n36370 , n36371 );
xor ( n36373 , n35978 , n35979 );
xor ( n36374 , n36373 , n36037 );
xor ( n36375 , n36044 , n36047 );
xor ( n36376 , n36375 , n36065 );
and ( n36377 , n36374 , n36376 );
xor ( n36378 , n36100 , n36127 );
xor ( n36379 , n36378 , n36130 );
and ( n36380 , n36376 , n36379 );
and ( n36381 , n36374 , n36379 );
or ( n36382 , n36377 , n36380 , n36381 );
and ( n36383 , n36372 , n36382 );
xor ( n36384 , n35977 , n36040 );
xor ( n36385 , n36384 , n36068 );
and ( n36386 , n36382 , n36385 );
and ( n36387 , n36372 , n36385 );
or ( n36388 , n36383 , n36386 , n36387 );
xor ( n36389 , n36071 , n36141 );
xor ( n36390 , n36389 , n36144 );
and ( n36391 , n36388 , n36390 );
xor ( n36392 , n36133 , n36135 );
xor ( n36393 , n36392 , n36138 );
xor ( n36394 , n36082 , n36087 );
xor ( n36395 , n36394 , n36097 );
xor ( n36396 , n36119 , n36121 );
xor ( n36397 , n36396 , n36124 );
and ( n36398 , n36395 , n36397 );
xor ( n36399 , n36227 , n36228 );
xor ( n36400 , n36344 , n36346 );
and ( n36401 , n31883 , n32173 );
and ( n36402 , n32155 , n31861 );
and ( n36403 , n36401 , n36402 );
buf ( n36404 , n15889 );
buf ( n36405 , n36404 );
and ( n36406 , n36403 , n36405 );
and ( n36407 , n36400 , n36406 );
and ( n36408 , n33692 , n31076 );
and ( n36409 , n33304 , n31073 );
and ( n36410 , n36408 , n36409 );
and ( n36411 , n32689 , n31590 );
and ( n36412 , n36409 , n36411 );
and ( n36413 , n36408 , n36411 );
or ( n36414 , n36410 , n36412 , n36413 );
and ( n36415 , n31084 , n33712 );
and ( n36416 , n31088 , n33347 );
and ( n36417 , n36415 , n36416 );
and ( n36418 , n31607 , n32671 );
and ( n36419 , n36416 , n36418 );
and ( n36420 , n36415 , n36418 );
or ( n36421 , n36417 , n36419 , n36420 );
and ( n36422 , n36414 , n36421 );
and ( n36423 , n36406 , n36422 );
and ( n36424 , n36400 , n36422 );
or ( n36425 , n36407 , n36423 , n36424 );
xor ( n36426 , n36306 , n36307 );
xor ( n36427 , n36426 , n36309 );
xor ( n36428 , n36313 , n36314 );
xor ( n36429 , n36428 , n36316 );
and ( n36430 , n36427 , n36429 );
xor ( n36431 , n36274 , n36275 );
xor ( n36432 , n36431 , n36277 );
and ( n36433 , n36429 , n36432 );
and ( n36434 , n36427 , n36432 );
or ( n36435 , n36430 , n36433 , n36434 );
xor ( n36436 , n36291 , n36292 );
xor ( n36437 , n36436 , n36294 );
xor ( n36438 , n36298 , n36299 );
xor ( n36439 , n36438 , n36301 );
and ( n36440 , n36437 , n36439 );
xor ( n36441 , n36259 , n36260 );
xor ( n36442 , n36441 , n36262 );
and ( n36443 , n36439 , n36442 );
and ( n36444 , n36437 , n36442 );
or ( n36445 , n36440 , n36443 , n36444 );
and ( n36446 , n36435 , n36445 );
and ( n36447 , n36425 , n36446 );
and ( n36448 , n36399 , n36447 );
xor ( n36449 , n36297 , n36304 );
xor ( n36450 , n36312 , n36319 );
and ( n36451 , n36449 , n36450 );
xor ( n36452 , n36103 , n36105 );
and ( n36453 , n36451 , n36452 );
and ( n36454 , n36447 , n36453 );
and ( n36455 , n36399 , n36453 );
or ( n36456 , n36448 , n36454 , n36455 );
and ( n36457 , n36397 , n36456 );
and ( n36458 , n36395 , n36456 );
or ( n36459 , n36398 , n36457 , n36458 );
xnor ( n36460 , n36110 , n36111 );
xnor ( n36461 , n36280 , n36287 );
or ( n36462 , n36460 , n36461 );
xnor ( n36463 , n36107 , n36108 );
xnor ( n36464 , n36265 , n36272 );
or ( n36465 , n36463 , n36464 );
and ( n36466 , n36462 , n36465 );
and ( n36467 , n34280 , n30791 );
and ( n36468 , n32949 , n31301 );
and ( n36469 , n36467 , n36468 );
and ( n36470 , n32365 , n31745 );
and ( n36471 , n36468 , n36470 );
and ( n36472 , n36467 , n36470 );
or ( n36473 , n36469 , n36471 , n36472 );
and ( n36474 , n34099 , n30788 );
and ( n36475 , n33896 , n30898 );
and ( n36476 , n36474 , n36475 );
and ( n36477 , n32736 , n31442 );
and ( n36478 , n36475 , n36477 );
and ( n36479 , n36474 , n36477 );
or ( n36480 , n36476 , n36478 , n36479 );
and ( n36481 , n36473 , n36480 );
xor ( n36482 , n36266 , n36267 );
xor ( n36483 , n36482 , n36269 );
and ( n36484 , n36480 , n36483 );
and ( n36485 , n36473 , n36483 );
or ( n36486 , n36481 , n36484 , n36485 );
xor ( n36487 , n36249 , n36251 );
xor ( n36488 , n36487 , n36254 );
and ( n36489 , n36486 , n36488 );
and ( n36490 , n30799 , n34253 );
and ( n36491 , n31278 , n32932 );
and ( n36492 , n36490 , n36491 );
and ( n36493 , n31736 , n32348 );
and ( n36494 , n36491 , n36493 );
and ( n36495 , n36490 , n36493 );
or ( n36496 , n36492 , n36494 , n36495 );
and ( n36497 , n30803 , n34082 );
and ( n36498 , n30889 , n33905 );
and ( n36499 , n36497 , n36498 );
and ( n36500 , n31464 , n32719 );
and ( n36501 , n36498 , n36500 );
and ( n36502 , n36497 , n36500 );
or ( n36503 , n36499 , n36501 , n36502 );
and ( n36504 , n36496 , n36503 );
xor ( n36505 , n36281 , n36282 );
xor ( n36506 , n36505 , n36284 );
and ( n36507 , n36503 , n36506 );
and ( n36508 , n36496 , n36506 );
or ( n36509 , n36504 , n36507 , n36508 );
xor ( n36510 , n36239 , n36241 );
xor ( n36511 , n36510 , n36244 );
and ( n36512 , n36509 , n36511 );
and ( n36513 , n36489 , n36512 );
and ( n36514 , n36466 , n36513 );
xor ( n36515 , n36247 , n36257 );
xor ( n36516 , n36273 , n36288 );
and ( n36517 , n36515 , n36516 );
xor ( n36518 , n36305 , n36320 );
and ( n36519 , n36516 , n36518 );
and ( n36520 , n36515 , n36518 );
or ( n36521 , n36517 , n36519 , n36520 );
and ( n36522 , n36513 , n36521 );
and ( n36523 , n36466 , n36521 );
or ( n36524 , n36514 , n36522 , n36523 );
xor ( n36525 , n36329 , n36331 );
xor ( n36526 , n36333 , n36334 );
and ( n36527 , n36525 , n36526 );
xor ( n36528 , n36337 , n36338 );
and ( n36529 , n36526 , n36528 );
and ( n36530 , n36525 , n36528 );
or ( n36531 , n36527 , n36529 , n36530 );
xor ( n36532 , n36230 , n36231 );
xor ( n36533 , n36532 , n36233 );
and ( n36534 , n36531 , n36533 );
xor ( n36535 , n36258 , n36289 );
xor ( n36536 , n36535 , n36321 );
and ( n36537 , n36533 , n36536 );
and ( n36538 , n36531 , n36536 );
or ( n36539 , n36534 , n36537 , n36538 );
and ( n36540 , n36524 , n36539 );
xor ( n36541 , n36202 , n36203 );
xor ( n36542 , n36541 , n36205 );
and ( n36543 , n36539 , n36542 );
and ( n36544 , n36524 , n36542 );
or ( n36545 , n36540 , n36543 , n36544 );
and ( n36546 , n36459 , n36545 );
xor ( n36547 , n36198 , n36200 );
xor ( n36548 , n36547 , n36208 );
and ( n36549 , n36545 , n36548 );
and ( n36550 , n36459 , n36548 );
or ( n36551 , n36546 , n36549 , n36550 );
and ( n36552 , n36393 , n36551 );
xor ( n36553 , n36193 , n36195 );
xor ( n36554 , n36553 , n36211 );
and ( n36555 , n36551 , n36554 );
and ( n36556 , n36393 , n36554 );
or ( n36557 , n36552 , n36555 , n36556 );
and ( n36558 , n36390 , n36557 );
and ( n36559 , n36388 , n36557 );
or ( n36560 , n36391 , n36558 , n36559 );
xor ( n36561 , n36186 , n36217 );
xor ( n36562 , n36561 , n36220 );
and ( n36563 , n36560 , n36562 );
xor ( n36564 , n36188 , n36190 );
xor ( n36565 , n36564 , n36214 );
xor ( n36566 , n36372 , n36382 );
xor ( n36567 , n36566 , n36385 );
xor ( n36568 , n36327 , n36366 );
xor ( n36569 , n36568 , n36369 );
xor ( n36570 , n36374 , n36376 );
xor ( n36571 , n36570 , n36379 );
and ( n36572 , n36569 , n36571 );
xor ( n36573 , n36229 , n36236 );
xor ( n36574 , n36573 , n36324 );
xor ( n36575 , n36342 , n36360 );
xor ( n36576 , n36575 , n36363 );
and ( n36577 , n36574 , n36576 );
xor ( n36578 , n36332 , n36335 );
xor ( n36579 , n36578 , n36339 );
xor ( n36580 , n36352 , n36354 );
xor ( n36581 , n36580 , n36357 );
and ( n36582 , n36579 , n36581 );
xor ( n36583 , n36486 , n36488 );
xor ( n36584 , n36509 , n36511 );
and ( n36585 , n36583 , n36584 );
xor ( n36586 , n36451 , n36452 );
and ( n36587 , n36585 , n36586 );
and ( n36588 , n36581 , n36587 );
and ( n36589 , n36579 , n36587 );
or ( n36590 , n36582 , n36588 , n36589 );
and ( n36591 , n36576 , n36590 );
and ( n36592 , n36574 , n36590 );
or ( n36593 , n36577 , n36591 , n36592 );
and ( n36594 , n36571 , n36593 );
and ( n36595 , n36569 , n36593 );
or ( n36596 , n36572 , n36594 , n36595 );
and ( n36597 , n36567 , n36596 );
xor ( n36598 , n36393 , n36551 );
xor ( n36599 , n36598 , n36554 );
and ( n36600 , n36596 , n36599 );
and ( n36601 , n36567 , n36599 );
or ( n36602 , n36597 , n36600 , n36601 );
and ( n36603 , n36565 , n36602 );
xor ( n36604 , n36388 , n36390 );
xor ( n36605 , n36604 , n36557 );
and ( n36606 , n36602 , n36605 );
and ( n36607 , n36565 , n36605 );
or ( n36608 , n36603 , n36606 , n36607 );
and ( n36609 , n36562 , n36608 );
and ( n36610 , n36560 , n36608 );
or ( n36611 , n36563 , n36609 , n36610 );
and ( n36612 , n36225 , n36611 );
and ( n36613 , n36223 , n36611 );
or ( n36614 , n36226 , n36612 , n36613 );
and ( n36615 , n36184 , n36614 );
xor ( n36616 , n36184 , n36614 );
xor ( n36617 , n36223 , n36225 );
xor ( n36618 , n36617 , n36611 );
xor ( n36619 , n36560 , n36562 );
xor ( n36620 , n36619 , n36608 );
xor ( n36621 , n36565 , n36602 );
xor ( n36622 , n36621 , n36605 );
xor ( n36623 , n36343 , n36347 );
xor ( n36624 , n36623 , n36349 );
xor ( n36625 , n36425 , n36446 );
and ( n36626 , n36624 , n36625 );
xor ( n36627 , n36462 , n36465 );
and ( n36628 , n36625 , n36627 );
and ( n36629 , n36624 , n36627 );
or ( n36630 , n36626 , n36628 , n36629 );
xor ( n36631 , n36489 , n36512 );
xor ( n36632 , n36403 , n36405 );
buf ( n36633 , n32057 );
buf ( n36634 , n15892 );
buf ( n36635 , n36634 );
and ( n36636 , n36633 , n36635 );
and ( n36637 , n36632 , n36636 );
and ( n36638 , n31238 , n33296 );
and ( n36639 , n33339 , n31247 );
and ( n36640 , n36638 , n36639 );
and ( n36641 , n36636 , n36640 );
and ( n36642 , n36632 , n36640 );
or ( n36643 , n36637 , n36641 , n36642 );
and ( n36644 , n30889 , n34082 );
and ( n36645 , n31084 , n33905 );
and ( n36646 , n36644 , n36645 );
and ( n36647 , n31607 , n32719 );
and ( n36648 , n36645 , n36647 );
and ( n36649 , n36644 , n36647 );
or ( n36650 , n36646 , n36648 , n36649 );
and ( n36651 , n31088 , n33712 );
and ( n36652 , n31238 , n33347 );
and ( n36653 , n36651 , n36652 );
and ( n36654 , n31736 , n32671 );
and ( n36655 , n36652 , n36654 );
and ( n36656 , n36651 , n36654 );
or ( n36657 , n36653 , n36655 , n36656 );
and ( n36658 , n36650 , n36657 );
and ( n36659 , n31278 , n33296 );
and ( n36660 , n31883 , n32348 );
and ( n36661 , n36659 , n36660 );
and ( n36662 , n32057 , n32173 );
and ( n36663 , n36660 , n36662 );
and ( n36664 , n36659 , n36662 );
or ( n36665 , n36661 , n36663 , n36664 );
and ( n36666 , n36657 , n36665 );
and ( n36667 , n36650 , n36665 );
or ( n36668 , n36658 , n36666 , n36667 );
and ( n36669 , n34099 , n30898 );
and ( n36670 , n33896 , n31076 );
and ( n36671 , n36669 , n36670 );
and ( n36672 , n32736 , n31590 );
and ( n36673 , n36670 , n36672 );
and ( n36674 , n36669 , n36672 );
or ( n36675 , n36671 , n36673 , n36674 );
and ( n36676 , n33692 , n31073 );
and ( n36677 , n33304 , n31247 );
and ( n36678 , n36676 , n36677 );
and ( n36679 , n32689 , n31745 );
and ( n36680 , n36677 , n36679 );
and ( n36681 , n36676 , n36679 );
or ( n36682 , n36678 , n36680 , n36681 );
and ( n36683 , n36675 , n36682 );
and ( n36684 , n33339 , n31301 );
and ( n36685 , n32365 , n31861 );
and ( n36686 , n36684 , n36685 );
and ( n36687 , n32155 , n32066 );
and ( n36688 , n36685 , n36687 );
and ( n36689 , n36684 , n36687 );
or ( n36690 , n36686 , n36688 , n36689 );
and ( n36691 , n36682 , n36690 );
and ( n36692 , n36675 , n36690 );
or ( n36693 , n36683 , n36691 , n36692 );
and ( n36694 , n36668 , n36693 );
and ( n36695 , n36643 , n36694 );
xor ( n36696 , n36400 , n36406 );
xor ( n36697 , n36696 , n36422 );
and ( n36698 , n36694 , n36697 );
and ( n36699 , n36643 , n36697 );
or ( n36700 , n36695 , n36698 , n36699 );
and ( n36701 , n36631 , n36700 );
xor ( n36702 , n36473 , n36480 );
xor ( n36703 , n36702 , n36483 );
xor ( n36704 , n36437 , n36439 );
xor ( n36705 , n36704 , n36442 );
and ( n36706 , n36703 , n36705 );
xor ( n36707 , n36496 , n36503 );
xor ( n36708 , n36707 , n36506 );
xor ( n36709 , n36427 , n36429 );
xor ( n36710 , n36709 , n36432 );
and ( n36711 , n36708 , n36710 );
and ( n36712 , n36706 , n36711 );
and ( n36713 , n36700 , n36712 );
and ( n36714 , n36631 , n36712 );
or ( n36715 , n36701 , n36713 , n36714 );
and ( n36716 , n36630 , n36715 );
xnor ( n36717 , n36460 , n36461 );
xnor ( n36718 , n36463 , n36464 );
and ( n36719 , n36717 , n36718 );
xor ( n36720 , n36101 , n36102 );
xor ( n36721 , n36435 , n36445 );
and ( n36722 , n36720 , n36721 );
xor ( n36723 , n36449 , n36450 );
and ( n36724 , n36721 , n36723 );
and ( n36725 , n36720 , n36723 );
or ( n36726 , n36722 , n36724 , n36725 );
and ( n36727 , n36719 , n36726 );
xor ( n36728 , n36515 , n36516 );
xor ( n36729 , n36728 , n36518 );
and ( n36730 , n36726 , n36729 );
and ( n36731 , n36719 , n36729 );
or ( n36732 , n36727 , n36730 , n36731 );
and ( n36733 , n36715 , n36732 );
and ( n36734 , n36630 , n36732 );
or ( n36735 , n36716 , n36733 , n36734 );
xor ( n36736 , n36399 , n36447 );
xor ( n36737 , n36736 , n36453 );
xor ( n36738 , n36466 , n36513 );
xor ( n36739 , n36738 , n36521 );
and ( n36740 , n36737 , n36739 );
xor ( n36741 , n36531 , n36533 );
xor ( n36742 , n36741 , n36536 );
and ( n36743 , n36739 , n36742 );
and ( n36744 , n36737 , n36742 );
or ( n36745 , n36740 , n36743 , n36744 );
and ( n36746 , n36735 , n36745 );
xor ( n36747 , n36395 , n36397 );
xor ( n36748 , n36747 , n36456 );
and ( n36749 , n36745 , n36748 );
and ( n36750 , n36735 , n36748 );
or ( n36751 , n36746 , n36749 , n36750 );
xor ( n36752 , n36459 , n36545 );
xor ( n36753 , n36752 , n36548 );
and ( n36754 , n36751 , n36753 );
xor ( n36755 , n36524 , n36539 );
xor ( n36756 , n36755 , n36542 );
xor ( n36757 , n36525 , n36526 );
xor ( n36758 , n36757 , n36528 );
xor ( n36759 , n36585 , n36586 );
and ( n36760 , n36758 , n36759 );
xor ( n36761 , n36490 , n36491 );
xor ( n36762 , n36761 , n36493 );
xor ( n36763 , n36497 , n36498 );
xor ( n36764 , n36763 , n36500 );
and ( n36765 , n36762 , n36764 );
xor ( n36766 , n36467 , n36468 );
xor ( n36767 , n36766 , n36470 );
xor ( n36768 , n36474 , n36475 );
xor ( n36769 , n36768 , n36477 );
and ( n36770 , n36767 , n36769 );
and ( n36771 , n36765 , n36770 );
xor ( n36772 , n36414 , n36421 );
and ( n36773 , n34280 , n30788 );
and ( n36774 , n32949 , n31442 );
or ( n36775 , n36773 , n36774 );
and ( n36776 , n30803 , n34253 );
and ( n36777 , n31464 , n32932 );
or ( n36778 , n36776 , n36777 );
and ( n36779 , n36775 , n36778 );
and ( n36780 , n36772 , n36779 );
xor ( n36781 , n36408 , n36409 );
xor ( n36782 , n36781 , n36411 );
xor ( n36783 , n36415 , n36416 );
xor ( n36784 , n36783 , n36418 );
and ( n36785 , n36782 , n36784 );
and ( n36786 , n36779 , n36785 );
and ( n36787 , n36772 , n36785 );
or ( n36788 , n36780 , n36786 , n36787 );
and ( n36789 , n36771 , n36788 );
xor ( n36790 , n36643 , n36694 );
xor ( n36791 , n36790 , n36697 );
and ( n36792 , n36788 , n36791 );
and ( n36793 , n36771 , n36791 );
or ( n36794 , n36789 , n36792 , n36793 );
and ( n36795 , n36759 , n36794 );
and ( n36796 , n36758 , n36794 );
or ( n36797 , n36760 , n36795 , n36796 );
xor ( n36798 , n36706 , n36711 );
xor ( n36799 , n36717 , n36718 );
and ( n36800 , n36798 , n36799 );
xor ( n36801 , n36583 , n36584 );
and ( n36802 , n36799 , n36801 );
and ( n36803 , n36798 , n36801 );
or ( n36804 , n36800 , n36802 , n36803 );
and ( n36805 , n33896 , n31073 );
and ( n36806 , n33692 , n31247 );
and ( n36807 , n36805 , n36806 );
and ( n36808 , n32736 , n31745 );
and ( n36809 , n36806 , n36808 );
and ( n36810 , n36805 , n36808 );
or ( n36811 , n36807 , n36809 , n36810 );
xor ( n36812 , n36644 , n36645 );
xor ( n36813 , n36812 , n36647 );
and ( n36814 , n36811 , n36813 );
xor ( n36815 , n36651 , n36652 );
xor ( n36816 , n36815 , n36654 );
and ( n36817 , n36813 , n36816 );
and ( n36818 , n36811 , n36816 );
or ( n36819 , n36814 , n36817 , n36818 );
xor ( n36820 , n36675 , n36682 );
xor ( n36821 , n36820 , n36690 );
or ( n36822 , n36819 , n36821 );
and ( n36823 , n31088 , n33905 );
and ( n36824 , n31238 , n33712 );
and ( n36825 , n36823 , n36824 );
and ( n36826 , n31736 , n32719 );
and ( n36827 , n36824 , n36826 );
and ( n36828 , n36823 , n36826 );
or ( n36829 , n36825 , n36827 , n36828 );
xor ( n36830 , n36669 , n36670 );
xor ( n36831 , n36830 , n36672 );
and ( n36832 , n36829 , n36831 );
xor ( n36833 , n36676 , n36677 );
xor ( n36834 , n36833 , n36679 );
and ( n36835 , n36831 , n36834 );
and ( n36836 , n36829 , n36834 );
or ( n36837 , n36832 , n36835 , n36836 );
xor ( n36838 , n36650 , n36657 );
xor ( n36839 , n36838 , n36665 );
or ( n36840 , n36837 , n36839 );
and ( n36841 , n36822 , n36840 );
xor ( n36842 , n36703 , n36705 );
xor ( n36843 , n36708 , n36710 );
and ( n36844 , n36842 , n36843 );
and ( n36845 , n36841 , n36844 );
xor ( n36846 , n36633 , n36635 );
xor ( n36847 , n36638 , n36639 );
and ( n36848 , n36846 , n36847 );
xor ( n36849 , n36401 , n36402 );
and ( n36850 , n36847 , n36849 );
and ( n36851 , n36846 , n36849 );
or ( n36852 , n36848 , n36850 , n36851 );
xor ( n36853 , n36632 , n36636 );
xor ( n36854 , n36853 , n36640 );
and ( n36855 , n36852 , n36854 );
xor ( n36856 , n36668 , n36693 );
and ( n36857 , n36854 , n36856 );
and ( n36858 , n36852 , n36856 );
or ( n36859 , n36855 , n36857 , n36858 );
and ( n36860 , n36844 , n36859 );
and ( n36861 , n36841 , n36859 );
or ( n36862 , n36845 , n36860 , n36861 );
and ( n36863 , n36804 , n36862 );
xor ( n36864 , n36765 , n36770 );
and ( n36865 , n30889 , n34253 );
and ( n36866 , n31084 , n34082 );
and ( n36867 , n36865 , n36866 );
and ( n36868 , n31607 , n32932 );
and ( n36869 , n36866 , n36868 );
and ( n36870 , n36865 , n36868 );
or ( n36871 , n36867 , n36869 , n36870 );
and ( n36872 , n31278 , n33347 );
and ( n36873 , n31464 , n33296 );
and ( n36874 , n36872 , n36873 );
and ( n36875 , n31883 , n32671 );
and ( n36876 , n36873 , n36875 );
and ( n36877 , n36872 , n36875 );
or ( n36878 , n36874 , n36876 , n36877 );
or ( n36879 , n36871 , n36878 );
and ( n36880 , n34280 , n30898 );
and ( n36881 , n34099 , n31076 );
and ( n36882 , n36880 , n36881 );
and ( n36883 , n32949 , n31590 );
and ( n36884 , n36881 , n36883 );
and ( n36885 , n36880 , n36883 );
or ( n36886 , n36882 , n36884 , n36885 );
and ( n36887 , n33304 , n31301 );
and ( n36888 , n33339 , n31442 );
and ( n36889 , n36887 , n36888 );
and ( n36890 , n32689 , n31861 );
and ( n36891 , n36888 , n36890 );
and ( n36892 , n36887 , n36890 );
or ( n36893 , n36889 , n36891 , n36892 );
or ( n36894 , n36886 , n36893 );
and ( n36895 , n36879 , n36894 );
and ( n36896 , n36864 , n36895 );
xor ( n36897 , n36762 , n36764 );
xor ( n36898 , n36767 , n36769 );
and ( n36899 , n36897 , n36898 );
and ( n36900 , n36895 , n36899 );
and ( n36901 , n36864 , n36899 );
or ( n36902 , n36896 , n36900 , n36901 );
xor ( n36903 , n36775 , n36778 );
xor ( n36904 , n36782 , n36784 );
and ( n36905 , n36903 , n36904 );
and ( n36906 , n32057 , n32348 );
and ( n36907 , n32365 , n32066 );
and ( n36908 , n36906 , n36907 );
buf ( n36909 , n15895 );
buf ( n36910 , n36909 );
and ( n36911 , n36908 , n36910 );
and ( n36912 , n36904 , n36911 );
and ( n36913 , n36903 , n36911 );
or ( n36914 , n36905 , n36912 , n36913 );
xor ( n36915 , n36684 , n36685 );
xor ( n36916 , n36915 , n36687 );
xor ( n36917 , n36659 , n36660 );
xor ( n36918 , n36917 , n36662 );
and ( n36919 , n36916 , n36918 );
xnor ( n36920 , n36773 , n36774 );
xnor ( n36921 , n36776 , n36777 );
and ( n36922 , n36920 , n36921 );
and ( n36923 , n36919 , n36922 );
xor ( n36924 , n36846 , n36847 );
xor ( n36925 , n36924 , n36849 );
and ( n36926 , n36922 , n36925 );
and ( n36927 , n36919 , n36925 );
or ( n36928 , n36923 , n36926 , n36927 );
and ( n36929 , n36914 , n36928 );
xor ( n36930 , n36772 , n36779 );
xor ( n36931 , n36930 , n36785 );
and ( n36932 , n36928 , n36931 );
and ( n36933 , n36914 , n36931 );
or ( n36934 , n36929 , n36932 , n36933 );
and ( n36935 , n36902 , n36934 );
xor ( n36936 , n36720 , n36721 );
xor ( n36937 , n36936 , n36723 );
and ( n36938 , n36934 , n36937 );
and ( n36939 , n36902 , n36937 );
or ( n36940 , n36935 , n36938 , n36939 );
and ( n36941 , n36862 , n36940 );
and ( n36942 , n36804 , n36940 );
or ( n36943 , n36863 , n36941 , n36942 );
and ( n36944 , n36797 , n36943 );
xor ( n36945 , n36624 , n36625 );
xor ( n36946 , n36945 , n36627 );
xor ( n36947 , n36631 , n36700 );
xor ( n36948 , n36947 , n36712 );
and ( n36949 , n36946 , n36948 );
xor ( n36950 , n36719 , n36726 );
xor ( n36951 , n36950 , n36729 );
and ( n36952 , n36948 , n36951 );
and ( n36953 , n36946 , n36951 );
or ( n36954 , n36949 , n36952 , n36953 );
and ( n36955 , n36943 , n36954 );
and ( n36956 , n36797 , n36954 );
or ( n36957 , n36944 , n36955 , n36956 );
and ( n36958 , n36756 , n36957 );
xor ( n36959 , n36579 , n36581 );
xor ( n36960 , n36959 , n36587 );
xor ( n36961 , n36630 , n36715 );
xor ( n36962 , n36961 , n36732 );
and ( n36963 , n36960 , n36962 );
xor ( n36964 , n36737 , n36739 );
xor ( n36965 , n36964 , n36742 );
and ( n36966 , n36962 , n36965 );
and ( n36967 , n36960 , n36965 );
or ( n36968 , n36963 , n36966 , n36967 );
and ( n36969 , n36957 , n36968 );
and ( n36970 , n36756 , n36968 );
or ( n36971 , n36958 , n36969 , n36970 );
and ( n36972 , n36753 , n36971 );
and ( n36973 , n36751 , n36971 );
or ( n36974 , n36754 , n36972 , n36973 );
xor ( n36975 , n36567 , n36596 );
xor ( n36976 , n36975 , n36599 );
and ( n36977 , n36974 , n36976 );
xor ( n36978 , n36569 , n36571 );
xor ( n36979 , n36978 , n36593 );
xor ( n36980 , n36574 , n36576 );
xor ( n36981 , n36980 , n36590 );
xor ( n36982 , n36735 , n36745 );
xor ( n36983 , n36982 , n36748 );
and ( n36984 , n36981 , n36983 );
xor ( n36985 , n36822 , n36840 );
xor ( n36986 , n36842 , n36843 );
and ( n36987 , n36985 , n36986 );
xnor ( n36988 , n36819 , n36821 );
xnor ( n36989 , n36837 , n36839 );
and ( n36990 , n36988 , n36989 );
and ( n36991 , n36986 , n36990 );
and ( n36992 , n36985 , n36990 );
or ( n36993 , n36987 , n36991 , n36992 );
xor ( n36994 , n36879 , n36894 );
xor ( n36995 , n36897 , n36898 );
and ( n36996 , n36994 , n36995 );
and ( n36997 , n31238 , n33905 );
and ( n36998 , n31278 , n33712 );
and ( n36999 , n36997 , n36998 );
and ( n37000 , n31883 , n32719 );
and ( n37001 , n36998 , n37000 );
and ( n37002 , n36997 , n37000 );
or ( n37003 , n36999 , n37001 , n37002 );
and ( n37004 , n31464 , n33347 );
and ( n37005 , n32057 , n32671 );
and ( n37006 , n37004 , n37005 );
and ( n37007 , n32155 , n32348 );
and ( n37008 , n37005 , n37007 );
and ( n37009 , n37004 , n37007 );
or ( n37010 , n37006 , n37008 , n37009 );
and ( n37011 , n37003 , n37010 );
xor ( n37012 , n36887 , n36888 );
xor ( n37013 , n37012 , n36890 );
and ( n37014 , n37010 , n37013 );
and ( n37015 , n37003 , n37013 );
or ( n37016 , n37011 , n37014 , n37015 );
and ( n37017 , n33896 , n31247 );
and ( n37018 , n33692 , n31301 );
and ( n37019 , n37017 , n37018 );
and ( n37020 , n32736 , n31861 );
and ( n37021 , n37018 , n37020 );
and ( n37022 , n37017 , n37020 );
or ( n37023 , n37019 , n37021 , n37022 );
and ( n37024 , n33304 , n31442 );
and ( n37025 , n32689 , n32066 );
and ( n37026 , n37024 , n37025 );
and ( n37027 , n32365 , n32173 );
and ( n37028 , n37025 , n37027 );
and ( n37029 , n37024 , n37027 );
or ( n37030 , n37026 , n37028 , n37029 );
and ( n37031 , n37023 , n37030 );
xor ( n37032 , n36872 , n36873 );
xor ( n37033 , n37032 , n36875 );
and ( n37034 , n37030 , n37033 );
and ( n37035 , n37023 , n37033 );
or ( n37036 , n37031 , n37034 , n37035 );
and ( n37037 , n37016 , n37036 );
and ( n37038 , n36995 , n37037 );
and ( n37039 , n36994 , n37037 );
or ( n37040 , n36996 , n37038 , n37039 );
xor ( n37041 , n36823 , n36824 );
xor ( n37042 , n37041 , n36826 );
xor ( n37043 , n36865 , n36866 );
xor ( n37044 , n37043 , n36868 );
or ( n37045 , n37042 , n37044 );
xor ( n37046 , n36805 , n36806 );
xor ( n37047 , n37046 , n36808 );
xor ( n37048 , n36880 , n36881 );
xor ( n37049 , n37048 , n36883 );
or ( n37050 , n37047 , n37049 );
and ( n37051 , n37045 , n37050 );
xor ( n37052 , n36829 , n36831 );
xor ( n37053 , n37052 , n36834 );
xor ( n37054 , n36811 , n36813 );
xor ( n37055 , n37054 , n36816 );
and ( n37056 , n37053 , n37055 );
and ( n37057 , n37051 , n37056 );
xnor ( n37058 , n36871 , n36878 );
xnor ( n37059 , n36886 , n36893 );
and ( n37060 , n37058 , n37059 );
and ( n37061 , n37056 , n37060 );
and ( n37062 , n37051 , n37060 );
or ( n37063 , n37057 , n37061 , n37062 );
and ( n37064 , n37040 , n37063 );
buf ( n37065 , n32155 );
buf ( n37066 , n15898 );
buf ( n37067 , n37066 );
or ( n37068 , n37065 , n37067 );
xor ( n37069 , n36908 , n36910 );
and ( n37070 , n37068 , n37069 );
xor ( n37071 , n36916 , n36918 );
and ( n37072 , n37069 , n37071 );
and ( n37073 , n37068 , n37071 );
or ( n37074 , n37070 , n37072 , n37073 );
xor ( n37075 , n36920 , n36921 );
and ( n37076 , n34280 , n31076 );
and ( n37077 , n34099 , n31073 );
and ( n37078 , n37076 , n37077 );
and ( n37079 , n32949 , n31745 );
and ( n37080 , n37077 , n37079 );
and ( n37081 , n37076 , n37079 );
or ( n37082 , n37078 , n37080 , n37081 );
and ( n37083 , n31084 , n34253 );
and ( n37084 , n31088 , n34082 );
and ( n37085 , n37083 , n37084 );
and ( n37086 , n31736 , n32932 );
and ( n37087 , n37084 , n37086 );
and ( n37088 , n37083 , n37086 );
or ( n37089 , n37085 , n37087 , n37088 );
and ( n37090 , n37082 , n37089 );
and ( n37091 , n37075 , n37090 );
xnor ( n37092 , n37065 , n37067 );
xor ( n37093 , n36906 , n36907 );
and ( n37094 , n37092 , n37093 );
and ( n37095 , n31607 , n33296 );
and ( n37096 , n33339 , n31590 );
and ( n37097 , n37095 , n37096 );
and ( n37098 , n37093 , n37097 );
and ( n37099 , n37092 , n37097 );
or ( n37100 , n37094 , n37098 , n37099 );
and ( n37101 , n37090 , n37100 );
and ( n37102 , n37075 , n37100 );
or ( n37103 , n37091 , n37101 , n37102 );
and ( n37104 , n37074 , n37103 );
xor ( n37105 , n36903 , n36904 );
xor ( n37106 , n37105 , n36911 );
and ( n37107 , n37103 , n37106 );
and ( n37108 , n37074 , n37106 );
or ( n37109 , n37104 , n37107 , n37108 );
and ( n37110 , n37063 , n37109 );
and ( n37111 , n37040 , n37109 );
or ( n37112 , n37064 , n37110 , n37111 );
and ( n37113 , n36993 , n37112 );
xor ( n37114 , n36852 , n36854 );
xor ( n37115 , n37114 , n36856 );
xor ( n37116 , n36864 , n36895 );
xor ( n37117 , n37116 , n36899 );
and ( n37118 , n37115 , n37117 );
xor ( n37119 , n36914 , n36928 );
xor ( n37120 , n37119 , n36931 );
and ( n37121 , n37117 , n37120 );
and ( n37122 , n37115 , n37120 );
or ( n37123 , n37118 , n37121 , n37122 );
and ( n37124 , n37112 , n37123 );
and ( n37125 , n36993 , n37123 );
or ( n37126 , n37113 , n37124 , n37125 );
xor ( n37127 , n36771 , n36788 );
xor ( n37128 , n37127 , n36791 );
xor ( n37129 , n36798 , n36799 );
xor ( n37130 , n37129 , n36801 );
and ( n37131 , n37128 , n37130 );
xor ( n37132 , n36841 , n36844 );
xor ( n37133 , n37132 , n36859 );
and ( n37134 , n37130 , n37133 );
and ( n37135 , n37128 , n37133 );
or ( n37136 , n37131 , n37134 , n37135 );
and ( n37137 , n37126 , n37136 );
xor ( n37138 , n36758 , n36759 );
xor ( n37139 , n37138 , n36794 );
and ( n37140 , n37136 , n37139 );
and ( n37141 , n37126 , n37139 );
or ( n37142 , n37137 , n37140 , n37141 );
xor ( n37143 , n36797 , n36943 );
xor ( n37144 , n37143 , n36954 );
and ( n37145 , n37142 , n37144 );
xor ( n37146 , n36960 , n36962 );
xor ( n37147 , n37146 , n36965 );
and ( n37148 , n37144 , n37147 );
and ( n37149 , n37142 , n37147 );
or ( n37150 , n37145 , n37148 , n37149 );
and ( n37151 , n36983 , n37150 );
and ( n37152 , n36981 , n37150 );
or ( n37153 , n36984 , n37151 , n37152 );
and ( n37154 , n36979 , n37153 );
xor ( n37155 , n36751 , n36753 );
xor ( n37156 , n37155 , n36971 );
and ( n37157 , n37153 , n37156 );
and ( n37158 , n36979 , n37156 );
or ( n37159 , n37154 , n37157 , n37158 );
and ( n37160 , n36976 , n37159 );
and ( n37161 , n36974 , n37159 );
or ( n37162 , n36977 , n37160 , n37161 );
or ( n37163 , n36622 , n37162 );
and ( n37164 , n36620 , n37163 );
xor ( n37165 , n36620 , n37163 );
xnor ( n37166 , n36622 , n37162 );
xor ( n37167 , n36974 , n36976 );
xor ( n37168 , n37167 , n37159 );
xor ( n37169 , n36979 , n37153 );
xor ( n37170 , n37169 , n37156 );
xor ( n37171 , n36756 , n36957 );
xor ( n37172 , n37171 , n36968 );
xor ( n37173 , n36981 , n36983 );
xor ( n37174 , n37173 , n37150 );
and ( n37175 , n37172 , n37174 );
xor ( n37176 , n36804 , n36862 );
xor ( n37177 , n37176 , n36940 );
xor ( n37178 , n36946 , n36948 );
xor ( n37179 , n37178 , n36951 );
and ( n37180 , n37177 , n37179 );
xor ( n37181 , n36902 , n36934 );
xor ( n37182 , n37181 , n36937 );
xor ( n37183 , n36919 , n36922 );
xor ( n37184 , n37183 , n36925 );
xor ( n37185 , n36988 , n36989 );
and ( n37186 , n37184 , n37185 );
and ( n37187 , n34099 , n31247 );
and ( n37188 , n33896 , n31301 );
and ( n37189 , n37187 , n37188 );
and ( n37190 , n32949 , n31861 );
and ( n37191 , n37188 , n37190 );
and ( n37192 , n37187 , n37190 );
or ( n37193 , n37189 , n37191 , n37192 );
and ( n37194 , n34280 , n31073 );
and ( n37195 , n33339 , n31745 );
and ( n37196 , n37194 , n37195 );
and ( n37197 , n32736 , n32066 );
and ( n37198 , n37195 , n37197 );
and ( n37199 , n37194 , n37197 );
or ( n37200 , n37196 , n37198 , n37199 );
and ( n37201 , n37193 , n37200 );
xor ( n37202 , n37083 , n37084 );
xor ( n37203 , n37202 , n37086 );
and ( n37204 , n37200 , n37203 );
and ( n37205 , n37193 , n37203 );
or ( n37206 , n37201 , n37204 , n37205 );
xor ( n37207 , n37023 , n37030 );
xor ( n37208 , n37207 , n37033 );
or ( n37209 , n37206 , n37208 );
and ( n37210 , n31238 , n34082 );
and ( n37211 , n31278 , n33905 );
and ( n37212 , n37210 , n37211 );
and ( n37213 , n31883 , n32932 );
and ( n37214 , n37211 , n37213 );
and ( n37215 , n37210 , n37213 );
or ( n37216 , n37212 , n37214 , n37215 );
and ( n37217 , n31088 , n34253 );
and ( n37218 , n31736 , n33296 );
and ( n37219 , n37217 , n37218 );
and ( n37220 , n32057 , n32719 );
and ( n37221 , n37218 , n37220 );
and ( n37222 , n37217 , n37220 );
or ( n37223 , n37219 , n37221 , n37222 );
and ( n37224 , n37216 , n37223 );
xor ( n37225 , n37076 , n37077 );
xor ( n37226 , n37225 , n37079 );
and ( n37227 , n37223 , n37226 );
and ( n37228 , n37216 , n37226 );
or ( n37229 , n37224 , n37227 , n37228 );
xor ( n37230 , n37003 , n37010 );
xor ( n37231 , n37230 , n37013 );
or ( n37232 , n37229 , n37231 );
and ( n37233 , n37209 , n37232 );
and ( n37234 , n37185 , n37233 );
and ( n37235 , n37184 , n37233 );
or ( n37236 , n37186 , n37234 , n37235 );
xor ( n37237 , n37016 , n37036 );
xor ( n37238 , n37045 , n37050 );
and ( n37239 , n37237 , n37238 );
xor ( n37240 , n37053 , n37055 );
and ( n37241 , n37238 , n37240 );
and ( n37242 , n37237 , n37240 );
or ( n37243 , n37239 , n37241 , n37242 );
xor ( n37244 , n37058 , n37059 );
xor ( n37245 , n36997 , n36998 );
xor ( n37246 , n37245 , n37000 );
xor ( n37247 , n37004 , n37005 );
xor ( n37248 , n37247 , n37007 );
or ( n37249 , n37246 , n37248 );
xor ( n37250 , n37017 , n37018 );
xor ( n37251 , n37250 , n37020 );
xor ( n37252 , n37024 , n37025 );
xor ( n37253 , n37252 , n37027 );
or ( n37254 , n37251 , n37253 );
and ( n37255 , n37249 , n37254 );
and ( n37256 , n37244 , n37255 );
xnor ( n37257 , n37042 , n37044 );
xnor ( n37258 , n37047 , n37049 );
and ( n37259 , n37257 , n37258 );
and ( n37260 , n37255 , n37259 );
and ( n37261 , n37244 , n37259 );
or ( n37262 , n37256 , n37260 , n37261 );
and ( n37263 , n37243 , n37262 );
xor ( n37264 , n37082 , n37089 );
and ( n37265 , n32155 , n32671 );
and ( n37266 , n32689 , n32173 );
and ( n37267 , n37265 , n37266 );
buf ( n37268 , n15901 );
buf ( n37269 , n37268 );
or ( n37270 , n37267 , n37269 );
and ( n37271 , n37264 , n37270 );
and ( n37272 , n33692 , n31442 );
and ( n37273 , n33304 , n31590 );
or ( n37274 , n37272 , n37273 );
and ( n37275 , n31464 , n33712 );
and ( n37276 , n31607 , n33347 );
or ( n37277 , n37275 , n37276 );
and ( n37278 , n37274 , n37277 );
and ( n37279 , n37270 , n37278 );
and ( n37280 , n37264 , n37278 );
or ( n37281 , n37271 , n37279 , n37280 );
xor ( n37282 , n37068 , n37069 );
xor ( n37283 , n37282 , n37071 );
and ( n37284 , n37281 , n37283 );
xor ( n37285 , n37075 , n37090 );
xor ( n37286 , n37285 , n37100 );
and ( n37287 , n37283 , n37286 );
and ( n37288 , n37281 , n37286 );
or ( n37289 , n37284 , n37287 , n37288 );
and ( n37290 , n37262 , n37289 );
and ( n37291 , n37243 , n37289 );
or ( n37292 , n37263 , n37290 , n37291 );
and ( n37293 , n37236 , n37292 );
xor ( n37294 , n36994 , n36995 );
xor ( n37295 , n37294 , n37037 );
xor ( n37296 , n37051 , n37056 );
xor ( n37297 , n37296 , n37060 );
and ( n37298 , n37295 , n37297 );
xor ( n37299 , n37074 , n37103 );
xor ( n37300 , n37299 , n37106 );
and ( n37301 , n37297 , n37300 );
and ( n37302 , n37295 , n37300 );
or ( n37303 , n37298 , n37301 , n37302 );
and ( n37304 , n37292 , n37303 );
and ( n37305 , n37236 , n37303 );
or ( n37306 , n37293 , n37304 , n37305 );
and ( n37307 , n37182 , n37306 );
xor ( n37308 , n36985 , n36986 );
xor ( n37309 , n37308 , n36990 );
xor ( n37310 , n37040 , n37063 );
xor ( n37311 , n37310 , n37109 );
and ( n37312 , n37309 , n37311 );
xor ( n37313 , n37115 , n37117 );
xor ( n37314 , n37313 , n37120 );
and ( n37315 , n37311 , n37314 );
and ( n37316 , n37309 , n37314 );
or ( n37317 , n37312 , n37315 , n37316 );
and ( n37318 , n37306 , n37317 );
and ( n37319 , n37182 , n37317 );
or ( n37320 , n37307 , n37318 , n37319 );
and ( n37321 , n37179 , n37320 );
and ( n37322 , n37177 , n37320 );
or ( n37323 , n37180 , n37321 , n37322 );
xor ( n37324 , n37142 , n37144 );
xor ( n37325 , n37324 , n37147 );
and ( n37326 , n37323 , n37325 );
xor ( n37327 , n37126 , n37136 );
xor ( n37328 , n37327 , n37139 );
xor ( n37329 , n36993 , n37112 );
xor ( n37330 , n37329 , n37123 );
xor ( n37331 , n37128 , n37130 );
xor ( n37332 , n37331 , n37133 );
and ( n37333 , n37330 , n37332 );
xor ( n37334 , n37209 , n37232 );
xnor ( n37335 , n37206 , n37208 );
xnor ( n37336 , n37229 , n37231 );
and ( n37337 , n37335 , n37336 );
and ( n37338 , n37334 , n37337 );
xor ( n37339 , n37092 , n37093 );
xor ( n37340 , n37339 , n37097 );
xor ( n37341 , n37249 , n37254 );
and ( n37342 , n37340 , n37341 );
xor ( n37343 , n37257 , n37258 );
and ( n37344 , n37341 , n37343 );
and ( n37345 , n37340 , n37343 );
or ( n37346 , n37342 , n37344 , n37345 );
and ( n37347 , n37337 , n37346 );
and ( n37348 , n37334 , n37346 );
or ( n37349 , n37338 , n37347 , n37348 );
buf ( n37350 , n32365 );
buf ( n37351 , n15904 );
buf ( n37352 , n37351 );
and ( n37353 , n37350 , n37352 );
xnor ( n37354 , n37272 , n37273 );
xnor ( n37355 , n37275 , n37276 );
and ( n37356 , n37354 , n37355 );
or ( n37357 , n37353 , n37356 );
and ( n37358 , n31238 , n34253 );
and ( n37359 , n31736 , n33347 );
and ( n37360 , n37358 , n37359 );
and ( n37361 , n31883 , n33296 );
and ( n37362 , n37359 , n37361 );
and ( n37363 , n37358 , n37361 );
or ( n37364 , n37360 , n37362 , n37363 );
xor ( n37365 , n37187 , n37188 );
xor ( n37366 , n37365 , n37190 );
and ( n37367 , n37364 , n37366 );
xor ( n37368 , n37194 , n37195 );
xor ( n37369 , n37368 , n37197 );
and ( n37370 , n37366 , n37369 );
and ( n37371 , n37364 , n37369 );
or ( n37372 , n37367 , n37370 , n37371 );
and ( n37373 , n34280 , n31247 );
and ( n37374 , n33304 , n31745 );
and ( n37375 , n37373 , n37374 );
and ( n37376 , n33339 , n31861 );
and ( n37377 , n37374 , n37376 );
and ( n37378 , n37373 , n37376 );
or ( n37379 , n37375 , n37377 , n37378 );
xor ( n37380 , n37210 , n37211 );
xor ( n37381 , n37380 , n37213 );
and ( n37382 , n37379 , n37381 );
xor ( n37383 , n37217 , n37218 );
xor ( n37384 , n37383 , n37220 );
and ( n37385 , n37381 , n37384 );
and ( n37386 , n37379 , n37384 );
or ( n37387 , n37382 , n37385 , n37386 );
and ( n37388 , n37372 , n37387 );
and ( n37389 , n37357 , n37388 );
and ( n37390 , n31607 , n33712 );
and ( n37391 , n32155 , n32719 );
and ( n37392 , n37390 , n37391 );
and ( n37393 , n32365 , n32671 );
and ( n37394 , n37391 , n37393 );
and ( n37395 , n37390 , n37393 );
or ( n37396 , n37392 , n37394 , n37395 );
not ( n37397 , n37396 );
and ( n37398 , n31278 , n34082 );
and ( n37399 , n31464 , n33905 );
and ( n37400 , n37398 , n37399 );
and ( n37401 , n32057 , n32932 );
and ( n37402 , n37399 , n37401 );
and ( n37403 , n37398 , n37401 );
or ( n37404 , n37400 , n37402 , n37403 );
and ( n37405 , n37397 , n37404 );
and ( n37406 , n33692 , n31590 );
and ( n37407 , n32736 , n32173 );
and ( n37408 , n37406 , n37407 );
and ( n37409 , n32689 , n32348 );
and ( n37410 , n37407 , n37409 );
and ( n37411 , n37406 , n37409 );
or ( n37412 , n37408 , n37410 , n37411 );
not ( n37413 , n37412 );
and ( n37414 , n34099 , n31301 );
and ( n37415 , n33896 , n31442 );
and ( n37416 , n37414 , n37415 );
and ( n37417 , n32949 , n32066 );
and ( n37418 , n37415 , n37417 );
and ( n37419 , n37414 , n37417 );
or ( n37420 , n37416 , n37418 , n37419 );
and ( n37421 , n37413 , n37420 );
and ( n37422 , n37405 , n37421 );
and ( n37423 , n37388 , n37422 );
and ( n37424 , n37357 , n37422 );
or ( n37425 , n37389 , n37423 , n37424 );
buf ( n37426 , n37396 );
buf ( n37427 , n37412 );
and ( n37428 , n37426 , n37427 );
xor ( n37429 , n37216 , n37223 );
xor ( n37430 , n37429 , n37226 );
xor ( n37431 , n37193 , n37200 );
xor ( n37432 , n37431 , n37203 );
and ( n37433 , n37430 , n37432 );
and ( n37434 , n37428 , n37433 );
xnor ( n37435 , n37246 , n37248 );
xnor ( n37436 , n37251 , n37253 );
and ( n37437 , n37435 , n37436 );
and ( n37438 , n37433 , n37437 );
and ( n37439 , n37428 , n37437 );
or ( n37440 , n37434 , n37438 , n37439 );
and ( n37441 , n37425 , n37440 );
xor ( n37442 , n37237 , n37238 );
xor ( n37443 , n37442 , n37240 );
and ( n37444 , n37440 , n37443 );
and ( n37445 , n37425 , n37443 );
or ( n37446 , n37441 , n37444 , n37445 );
and ( n37447 , n37349 , n37446 );
xor ( n37448 , n37184 , n37185 );
xor ( n37449 , n37448 , n37233 );
and ( n37450 , n37446 , n37449 );
and ( n37451 , n37349 , n37449 );
or ( n37452 , n37447 , n37450 , n37451 );
xor ( n37453 , n37236 , n37292 );
xor ( n37454 , n37453 , n37303 );
and ( n37455 , n37452 , n37454 );
xor ( n37456 , n37309 , n37311 );
xor ( n37457 , n37456 , n37314 );
and ( n37458 , n37454 , n37457 );
and ( n37459 , n37452 , n37457 );
or ( n37460 , n37455 , n37458 , n37459 );
and ( n37461 , n37332 , n37460 );
and ( n37462 , n37330 , n37460 );
or ( n37463 , n37333 , n37461 , n37462 );
and ( n37464 , n37328 , n37463 );
xor ( n37465 , n37177 , n37179 );
xor ( n37466 , n37465 , n37320 );
and ( n37467 , n37463 , n37466 );
and ( n37468 , n37328 , n37466 );
or ( n37469 , n37464 , n37467 , n37468 );
and ( n37470 , n37325 , n37469 );
and ( n37471 , n37323 , n37469 );
or ( n37472 , n37326 , n37470 , n37471 );
and ( n37473 , n37174 , n37472 );
and ( n37474 , n37172 , n37472 );
or ( n37475 , n37175 , n37473 , n37474 );
and ( n37476 , n37170 , n37475 );
xor ( n37477 , n37170 , n37475 );
xor ( n37478 , n37172 , n37174 );
xor ( n37479 , n37478 , n37472 );
not ( n37480 , n37479 );
xor ( n37481 , n37323 , n37325 );
xor ( n37482 , n37481 , n37469 );
xor ( n37483 , n37328 , n37463 );
xor ( n37484 , n37483 , n37466 );
xor ( n37485 , n37182 , n37306 );
xor ( n37486 , n37485 , n37317 );
xor ( n37487 , n37330 , n37332 );
xor ( n37488 , n37487 , n37460 );
and ( n37489 , n37486 , n37488 );
xor ( n37490 , n37243 , n37262 );
xor ( n37491 , n37490 , n37289 );
xor ( n37492 , n37295 , n37297 );
xor ( n37493 , n37492 , n37300 );
and ( n37494 , n37491 , n37493 );
xor ( n37495 , n37244 , n37255 );
xor ( n37496 , n37495 , n37259 );
xor ( n37497 , n37281 , n37283 );
xor ( n37498 , n37497 , n37286 );
and ( n37499 , n37496 , n37498 );
xor ( n37500 , n37264 , n37270 );
xor ( n37501 , n37500 , n37278 );
xor ( n37502 , n37335 , n37336 );
and ( n37503 , n37501 , n37502 );
xor ( n37504 , n37397 , n37404 );
xor ( n37505 , n37413 , n37420 );
and ( n37506 , n37504 , n37505 );
xnor ( n37507 , n37267 , n37269 );
and ( n37508 , n37506 , n37507 );
and ( n37509 , n37502 , n37508 );
and ( n37510 , n37501 , n37508 );
or ( n37511 , n37503 , n37509 , n37510 );
and ( n37512 , n37498 , n37511 );
and ( n37513 , n37496 , n37511 );
or ( n37514 , n37499 , n37512 , n37513 );
and ( n37515 , n37493 , n37514 );
and ( n37516 , n37491 , n37514 );
or ( n37517 , n37494 , n37515 , n37516 );
xor ( n37518 , n37452 , n37454 );
xor ( n37519 , n37518 , n37457 );
and ( n37520 , n37517 , n37519 );
and ( n37521 , n34280 , n31301 );
and ( n37522 , n34099 , n31442 );
and ( n37523 , n37521 , n37522 );
and ( n37524 , n33339 , n32066 );
and ( n37525 , n37522 , n37524 );
and ( n37526 , n37521 , n37524 );
or ( n37527 , n37523 , n37525 , n37526 );
xor ( n37528 , n37358 , n37359 );
xor ( n37529 , n37528 , n37361 );
and ( n37530 , n37527 , n37529 );
xor ( n37531 , n37390 , n37391 );
xor ( n37532 , n37531 , n37393 );
and ( n37533 , n37529 , n37532 );
and ( n37534 , n37527 , n37532 );
or ( n37535 , n37530 , n37533 , n37534 );
xor ( n37536 , n37379 , n37381 );
xor ( n37537 , n37536 , n37384 );
or ( n37538 , n37535 , n37537 );
and ( n37539 , n31278 , n34253 );
and ( n37540 , n31464 , n34082 );
and ( n37541 , n37539 , n37540 );
and ( n37542 , n32057 , n33296 );
and ( n37543 , n37540 , n37542 );
and ( n37544 , n37539 , n37542 );
or ( n37545 , n37541 , n37543 , n37544 );
xor ( n37546 , n37373 , n37374 );
xor ( n37547 , n37546 , n37376 );
and ( n37548 , n37545 , n37547 );
xor ( n37549 , n37406 , n37407 );
xor ( n37550 , n37549 , n37409 );
and ( n37551 , n37547 , n37550 );
and ( n37552 , n37545 , n37550 );
or ( n37553 , n37548 , n37551 , n37552 );
xor ( n37554 , n37364 , n37366 );
xor ( n37555 , n37554 , n37369 );
or ( n37556 , n37553 , n37555 );
and ( n37557 , n37538 , n37556 );
xor ( n37558 , n37095 , n37096 );
xor ( n37559 , n37274 , n37277 );
and ( n37560 , n37558 , n37559 );
xor ( n37561 , n37372 , n37387 );
and ( n37562 , n37559 , n37561 );
and ( n37563 , n37558 , n37561 );
or ( n37564 , n37560 , n37562 , n37563 );
and ( n37565 , n37557 , n37564 );
xor ( n37566 , n37405 , n37421 );
xor ( n37567 , n37426 , n37427 );
and ( n37568 , n37566 , n37567 );
xor ( n37569 , n37430 , n37432 );
and ( n37570 , n37567 , n37569 );
and ( n37571 , n37566 , n37569 );
or ( n37572 , n37568 , n37570 , n37571 );
and ( n37573 , n37564 , n37572 );
and ( n37574 , n37557 , n37572 );
or ( n37575 , n37565 , n37573 , n37574 );
xor ( n37576 , n37340 , n37341 );
xor ( n37577 , n37576 , n37343 );
xor ( n37578 , n37357 , n37388 );
xor ( n37579 , n37578 , n37422 );
and ( n37580 , n37577 , n37579 );
xor ( n37581 , n37428 , n37433 );
xor ( n37582 , n37581 , n37437 );
and ( n37583 , n37579 , n37582 );
and ( n37584 , n37577 , n37582 );
or ( n37585 , n37580 , n37583 , n37584 );
and ( n37586 , n37575 , n37585 );
xor ( n37587 , n37334 , n37337 );
xor ( n37588 , n37587 , n37346 );
and ( n37589 , n37585 , n37588 );
and ( n37590 , n37575 , n37588 );
or ( n37591 , n37586 , n37589 , n37590 );
xor ( n37592 , n37349 , n37446 );
xor ( n37593 , n37592 , n37449 );
and ( n37594 , n37591 , n37593 );
xor ( n37595 , n37425 , n37440 );
xor ( n37596 , n37595 , n37443 );
xor ( n37597 , n37506 , n37507 );
xor ( n37598 , n37350 , n37352 );
and ( n37599 , n32365 , n32719 );
and ( n37600 , n32736 , n32348 );
and ( n37601 , n37599 , n37600 );
buf ( n37602 , n15907 );
buf ( n37603 , n37602 );
and ( n37604 , n37601 , n37603 );
and ( n37605 , n37598 , n37604 );
and ( n37606 , n33692 , n31745 );
and ( n37607 , n33304 , n31861 );
and ( n37608 , n37606 , n37607 );
and ( n37609 , n32949 , n32173 );
and ( n37610 , n37607 , n37609 );
and ( n37611 , n37606 , n37609 );
or ( n37612 , n37608 , n37610 , n37611 );
and ( n37613 , n31736 , n33712 );
and ( n37614 , n31883 , n33347 );
and ( n37615 , n37613 , n37614 );
and ( n37616 , n32155 , n32932 );
and ( n37617 , n37614 , n37616 );
and ( n37618 , n37613 , n37616 );
or ( n37619 , n37615 , n37617 , n37618 );
and ( n37620 , n37612 , n37619 );
and ( n37621 , n37604 , n37620 );
and ( n37622 , n37598 , n37620 );
or ( n37623 , n37605 , n37621 , n37622 );
and ( n37624 , n37597 , n37623 );
xnor ( n37625 , n37353 , n37356 );
and ( n37626 , n37623 , n37625 );
and ( n37627 , n37597 , n37625 );
or ( n37628 , n37624 , n37626 , n37627 );
xor ( n37629 , n37601 , n37603 );
buf ( n37630 , n32689 );
buf ( n37631 , n15910 );
buf ( n37632 , n37631 );
and ( n37633 , n37630 , n37632 );
and ( n37634 , n37629 , n37633 );
and ( n37635 , n31607 , n33905 );
and ( n37636 , n33896 , n31590 );
and ( n37637 , n37635 , n37636 );
and ( n37638 , n37633 , n37637 );
and ( n37639 , n37629 , n37637 );
or ( n37640 , n37634 , n37638 , n37639 );
xor ( n37641 , n37414 , n37415 );
xor ( n37642 , n37641 , n37417 );
xor ( n37643 , n37398 , n37399 );
xor ( n37644 , n37643 , n37401 );
and ( n37645 , n37642 , n37644 );
and ( n37646 , n37640 , n37645 );
xor ( n37647 , n37598 , n37604 );
xor ( n37648 , n37647 , n37620 );
and ( n37649 , n37645 , n37648 );
and ( n37650 , n37640 , n37648 );
or ( n37651 , n37646 , n37649 , n37650 );
not ( n37652 , n37651 );
xnor ( n37653 , n37535 , n37537 );
xnor ( n37654 , n37553 , n37555 );
and ( n37655 , n37653 , n37654 );
and ( n37656 , n37652 , n37655 );
and ( n37657 , n37628 , n37656 );
buf ( n37658 , n37651 );
and ( n37659 , n37656 , n37658 );
and ( n37660 , n37628 , n37658 );
or ( n37661 , n37657 , n37659 , n37660 );
and ( n37662 , n37596 , n37661 );
xor ( n37663 , n37435 , n37436 );
xor ( n37664 , n37538 , n37556 );
and ( n37665 , n37663 , n37664 );
and ( n37666 , n34280 , n31442 );
and ( n37667 , n34099 , n31590 );
and ( n37668 , n37666 , n37667 );
and ( n37669 , n33339 , n32173 );
and ( n37670 , n37667 , n37669 );
and ( n37671 , n37666 , n37669 );
or ( n37672 , n37668 , n37670 , n37671 );
and ( n37673 , n33896 , n31745 );
and ( n37674 , n32949 , n32348 );
and ( n37675 , n37673 , n37674 );
and ( n37676 , n32736 , n32671 );
and ( n37677 , n37674 , n37676 );
and ( n37678 , n37673 , n37676 );
or ( n37679 , n37675 , n37677 , n37678 );
and ( n37680 , n37672 , n37679 );
xor ( n37681 , n37613 , n37614 );
xor ( n37682 , n37681 , n37616 );
and ( n37683 , n37679 , n37682 );
and ( n37684 , n37672 , n37682 );
or ( n37685 , n37680 , n37683 , n37684 );
xor ( n37686 , n37527 , n37529 );
xor ( n37687 , n37686 , n37532 );
or ( n37688 , n37685 , n37687 );
and ( n37689 , n31464 , n34253 );
and ( n37690 , n31607 , n34082 );
and ( n37691 , n37689 , n37690 );
and ( n37692 , n32155 , n33296 );
and ( n37693 , n37690 , n37692 );
and ( n37694 , n37689 , n37692 );
or ( n37695 , n37691 , n37693 , n37694 );
and ( n37696 , n31736 , n33905 );
and ( n37697 , n32365 , n32932 );
and ( n37698 , n37696 , n37697 );
and ( n37699 , n32689 , n32719 );
and ( n37700 , n37697 , n37699 );
and ( n37701 , n37696 , n37699 );
or ( n37702 , n37698 , n37700 , n37701 );
and ( n37703 , n37695 , n37702 );
xor ( n37704 , n37606 , n37607 );
xor ( n37705 , n37704 , n37609 );
and ( n37706 , n37702 , n37705 );
and ( n37707 , n37695 , n37705 );
or ( n37708 , n37703 , n37706 , n37707 );
xor ( n37709 , n37545 , n37547 );
xor ( n37710 , n37709 , n37550 );
or ( n37711 , n37708 , n37710 );
and ( n37712 , n37688 , n37711 );
and ( n37713 , n37664 , n37712 );
and ( n37714 , n37663 , n37712 );
or ( n37715 , n37665 , n37713 , n37714 );
xor ( n37716 , n37265 , n37266 );
xor ( n37717 , n37354 , n37355 );
and ( n37718 , n37716 , n37717 );
xor ( n37719 , n37504 , n37505 );
and ( n37720 , n37717 , n37719 );
and ( n37721 , n37716 , n37719 );
or ( n37722 , n37718 , n37720 , n37721 );
xor ( n37723 , n37558 , n37559 );
xor ( n37724 , n37723 , n37561 );
and ( n37725 , n37722 , n37724 );
xor ( n37726 , n37566 , n37567 );
xor ( n37727 , n37726 , n37569 );
and ( n37728 , n37724 , n37727 );
and ( n37729 , n37722 , n37727 );
or ( n37730 , n37725 , n37728 , n37729 );
and ( n37731 , n37715 , n37730 );
xor ( n37732 , n37501 , n37502 );
xor ( n37733 , n37732 , n37508 );
and ( n37734 , n37730 , n37733 );
and ( n37735 , n37715 , n37733 );
or ( n37736 , n37731 , n37734 , n37735 );
and ( n37737 , n37661 , n37736 );
and ( n37738 , n37596 , n37736 );
or ( n37739 , n37662 , n37737 , n37738 );
and ( n37740 , n37593 , n37739 );
and ( n37741 , n37591 , n37739 );
or ( n37742 , n37594 , n37740 , n37741 );
and ( n37743 , n37519 , n37742 );
and ( n37744 , n37517 , n37742 );
or ( n37745 , n37520 , n37743 , n37744 );
and ( n37746 , n37488 , n37745 );
and ( n37747 , n37486 , n37745 );
or ( n37748 , n37489 , n37746 , n37747 );
and ( n37749 , n37484 , n37748 );
xor ( n37750 , n37484 , n37748 );
xor ( n37751 , n37486 , n37488 );
xor ( n37752 , n37751 , n37745 );
xor ( n37753 , n37491 , n37493 );
xor ( n37754 , n37753 , n37514 );
xor ( n37755 , n37496 , n37498 );
xor ( n37756 , n37755 , n37511 );
xor ( n37757 , n37575 , n37585 );
xor ( n37758 , n37757 , n37588 );
and ( n37759 , n37756 , n37758 );
xor ( n37760 , n37557 , n37564 );
xor ( n37761 , n37760 , n37572 );
xor ( n37762 , n37577 , n37579 );
xor ( n37763 , n37762 , n37582 );
and ( n37764 , n37761 , n37763 );
xor ( n37765 , n37597 , n37623 );
xor ( n37766 , n37765 , n37625 );
xor ( n37767 , n37652 , n37655 );
and ( n37768 , n37766 , n37767 );
xor ( n37769 , n37612 , n37619 );
xor ( n37770 , n37642 , n37644 );
and ( n37771 , n37769 , n37770 );
and ( n37772 , n33692 , n31861 );
and ( n37773 , n33304 , n32066 );
or ( n37774 , n37772 , n37773 );
and ( n37775 , n31883 , n33712 );
and ( n37776 , n32057 , n33347 );
or ( n37777 , n37775 , n37776 );
and ( n37778 , n37774 , n37777 );
and ( n37779 , n37770 , n37778 );
and ( n37780 , n37769 , n37778 );
or ( n37781 , n37771 , n37779 , n37780 );
xor ( n37782 , n37640 , n37645 );
xor ( n37783 , n37782 , n37648 );
and ( n37784 , n37781 , n37783 );
xor ( n37785 , n37688 , n37711 );
and ( n37786 , n37783 , n37785 );
and ( n37787 , n37781 , n37785 );
or ( n37788 , n37784 , n37786 , n37787 );
and ( n37789 , n37767 , n37788 );
and ( n37790 , n37766 , n37788 );
or ( n37791 , n37768 , n37789 , n37790 );
and ( n37792 , n37763 , n37791 );
and ( n37793 , n37761 , n37791 );
or ( n37794 , n37764 , n37792 , n37793 );
and ( n37795 , n37758 , n37794 );
and ( n37796 , n37756 , n37794 );
or ( n37797 , n37759 , n37795 , n37796 );
and ( n37798 , n37754 , n37797 );
xor ( n37799 , n37591 , n37593 );
xor ( n37800 , n37799 , n37739 );
and ( n37801 , n37797 , n37800 );
and ( n37802 , n37754 , n37800 );
or ( n37803 , n37798 , n37801 , n37802 );
xor ( n37804 , n37517 , n37519 );
xor ( n37805 , n37804 , n37742 );
and ( n37806 , n37803 , n37805 );
xor ( n37807 , n37653 , n37654 );
xnor ( n37808 , n37685 , n37687 );
xnor ( n37809 , n37708 , n37710 );
and ( n37810 , n37808 , n37809 );
and ( n37811 , n37807 , n37810 );
xor ( n37812 , n37521 , n37522 );
xor ( n37813 , n37812 , n37524 );
xor ( n37814 , n37539 , n37540 );
xor ( n37815 , n37814 , n37542 );
and ( n37816 , n37813 , n37815 );
xor ( n37817 , n37629 , n37633 );
xor ( n37818 , n37817 , n37637 );
and ( n37819 , n37816 , n37818 );
xnor ( n37820 , n37772 , n37773 );
xnor ( n37821 , n37775 , n37776 );
and ( n37822 , n37820 , n37821 );
not ( n37823 , n37822 );
xor ( n37824 , n37630 , n37632 );
and ( n37825 , n37823 , n37824 );
and ( n37826 , n37818 , n37825 );
and ( n37827 , n37816 , n37825 );
or ( n37828 , n37819 , n37826 , n37827 );
and ( n37829 , n37810 , n37828 );
and ( n37830 , n37807 , n37828 );
or ( n37831 , n37811 , n37829 , n37830 );
buf ( n37832 , n37822 );
xor ( n37833 , n37689 , n37690 );
xor ( n37834 , n37833 , n37692 );
xor ( n37835 , n37696 , n37697 );
xor ( n37836 , n37835 , n37699 );
or ( n37837 , n37834 , n37836 );
xor ( n37838 , n37666 , n37667 );
xor ( n37839 , n37838 , n37669 );
xor ( n37840 , n37673 , n37674 );
xor ( n37841 , n37840 , n37676 );
or ( n37842 , n37839 , n37841 );
and ( n37843 , n37837 , n37842 );
and ( n37844 , n37832 , n37843 );
and ( n37845 , n31736 , n34082 );
and ( n37846 , n31883 , n33905 );
and ( n37847 , n37845 , n37846 );
and ( n37848 , n32365 , n33296 );
and ( n37849 , n37846 , n37848 );
and ( n37850 , n37845 , n37848 );
or ( n37851 , n37847 , n37849 , n37850 );
not ( n37852 , n37851 );
and ( n37853 , n31607 , n34253 );
and ( n37854 , n32057 , n33712 );
and ( n37855 , n37853 , n37854 );
and ( n37856 , n32155 , n33347 );
and ( n37857 , n37854 , n37856 );
and ( n37858 , n37853 , n37856 );
or ( n37859 , n37855 , n37857 , n37858 );
and ( n37860 , n37852 , n37859 );
and ( n37861 , n34099 , n31745 );
and ( n37862 , n33896 , n31861 );
and ( n37863 , n37861 , n37862 );
and ( n37864 , n33339 , n32348 );
and ( n37865 , n37862 , n37864 );
and ( n37866 , n37861 , n37864 );
or ( n37867 , n37863 , n37865 , n37866 );
not ( n37868 , n37867 );
and ( n37869 , n34280 , n31590 );
and ( n37870 , n33692 , n32066 );
and ( n37871 , n37869 , n37870 );
and ( n37872 , n33304 , n32173 );
and ( n37873 , n37870 , n37872 );
and ( n37874 , n37869 , n37872 );
or ( n37875 , n37871 , n37873 , n37874 );
and ( n37876 , n37868 , n37875 );
and ( n37877 , n37860 , n37876 );
and ( n37878 , n37843 , n37877 );
and ( n37879 , n37832 , n37877 );
or ( n37880 , n37844 , n37878 , n37879 );
buf ( n37881 , n37851 );
buf ( n37882 , n37867 );
and ( n37883 , n37881 , n37882 );
xor ( n37884 , n37695 , n37702 );
xor ( n37885 , n37884 , n37705 );
xor ( n37886 , n37672 , n37679 );
xor ( n37887 , n37886 , n37682 );
and ( n37888 , n37885 , n37887 );
and ( n37889 , n37883 , n37888 );
xor ( n37890 , n37635 , n37636 );
xor ( n37891 , n37599 , n37600 );
and ( n37892 , n37890 , n37891 );
xor ( n37893 , n37774 , n37777 );
and ( n37894 , n37891 , n37893 );
and ( n37895 , n37890 , n37893 );
or ( n37896 , n37892 , n37894 , n37895 );
and ( n37897 , n37888 , n37896 );
and ( n37898 , n37883 , n37896 );
or ( n37899 , n37889 , n37897 , n37898 );
and ( n37900 , n37880 , n37899 );
xor ( n37901 , n37716 , n37717 );
xor ( n37902 , n37901 , n37719 );
and ( n37903 , n37899 , n37902 );
and ( n37904 , n37880 , n37902 );
or ( n37905 , n37900 , n37903 , n37904 );
and ( n37906 , n37831 , n37905 );
xor ( n37907 , n37663 , n37664 );
xor ( n37908 , n37907 , n37712 );
and ( n37909 , n37905 , n37908 );
and ( n37910 , n37831 , n37908 );
or ( n37911 , n37906 , n37909 , n37910 );
xor ( n37912 , n37628 , n37656 );
xor ( n37913 , n37912 , n37658 );
and ( n37914 , n37911 , n37913 );
xor ( n37915 , n37715 , n37730 );
xor ( n37916 , n37915 , n37733 );
and ( n37917 , n37913 , n37916 );
and ( n37918 , n37911 , n37916 );
or ( n37919 , n37914 , n37917 , n37918 );
xor ( n37920 , n37596 , n37661 );
xor ( n37921 , n37920 , n37736 );
and ( n37922 , n37919 , n37921 );
xor ( n37923 , n37722 , n37724 );
xor ( n37924 , n37923 , n37727 );
xor ( n37925 , n37769 , n37770 );
xor ( n37926 , n37925 , n37778 );
xor ( n37927 , n37808 , n37809 );
and ( n37928 , n37926 , n37927 );
xor ( n37929 , n37813 , n37815 );
and ( n37930 , n32689 , n32932 );
and ( n37931 , n32949 , n32671 );
and ( n37932 , n37930 , n37931 );
buf ( n37933 , n15913 );
buf ( n37934 , n37933 );
and ( n37935 , n37932 , n37934 );
and ( n37936 , n37929 , n37935 );
xor ( n37937 , n37823 , n37824 );
and ( n37938 , n37935 , n37937 );
and ( n37939 , n37929 , n37937 );
or ( n37940 , n37936 , n37938 , n37939 );
and ( n37941 , n37927 , n37940 );
and ( n37942 , n37926 , n37940 );
or ( n37943 , n37928 , n37941 , n37942 );
xor ( n37944 , n37837 , n37842 );
xor ( n37945 , n37860 , n37876 );
and ( n37946 , n37944 , n37945 );
xor ( n37947 , n37881 , n37882 );
and ( n37948 , n37945 , n37947 );
and ( n37949 , n37944 , n37947 );
or ( n37950 , n37946 , n37948 , n37949 );
xor ( n37951 , n37885 , n37887 );
xor ( n37952 , n37932 , n37934 );
buf ( n37953 , n32736 );
buf ( n37954 , n15916 );
buf ( n37955 , n37954 );
and ( n37956 , n37953 , n37955 );
and ( n37957 , n37952 , n37956 );
and ( n37958 , n34099 , n31861 );
and ( n37959 , n33339 , n32671 );
and ( n37960 , n37958 , n37959 );
and ( n37961 , n32949 , n32719 );
and ( n37962 , n37959 , n37961 );
and ( n37963 , n37958 , n37961 );
or ( n37964 , n37960 , n37962 , n37963 );
and ( n37965 , n31883 , n34082 );
and ( n37966 , n32689 , n33296 );
and ( n37967 , n37965 , n37966 );
and ( n37968 , n32736 , n32932 );
and ( n37969 , n37966 , n37968 );
and ( n37970 , n37965 , n37968 );
or ( n37971 , n37967 , n37969 , n37970 );
and ( n37972 , n37964 , n37971 );
and ( n37973 , n37956 , n37972 );
and ( n37974 , n37952 , n37972 );
or ( n37975 , n37957 , n37973 , n37974 );
and ( n37976 , n37951 , n37975 );
and ( n37977 , n31736 , n34253 );
and ( n37978 , n32155 , n33712 );
and ( n37979 , n37977 , n37978 );
and ( n37980 , n32365 , n33347 );
and ( n37981 , n37978 , n37980 );
and ( n37982 , n37977 , n37980 );
or ( n37983 , n37979 , n37981 , n37982 );
xor ( n37984 , n37861 , n37862 );
xor ( n37985 , n37984 , n37864 );
and ( n37986 , n37983 , n37985 );
xor ( n37987 , n37869 , n37870 );
xor ( n37988 , n37987 , n37872 );
and ( n37989 , n37985 , n37988 );
and ( n37990 , n37983 , n37988 );
or ( n37991 , n37986 , n37989 , n37990 );
and ( n37992 , n34280 , n31745 );
and ( n37993 , n33692 , n32173 );
and ( n37994 , n37992 , n37993 );
and ( n37995 , n33304 , n32348 );
and ( n37996 , n37993 , n37995 );
and ( n37997 , n37992 , n37995 );
or ( n37998 , n37994 , n37996 , n37997 );
xor ( n37999 , n37845 , n37846 );
xor ( n38000 , n37999 , n37848 );
and ( n38001 , n37998 , n38000 );
xor ( n38002 , n37853 , n37854 );
xor ( n38003 , n38002 , n37856 );
and ( n38004 , n38000 , n38003 );
and ( n38005 , n37998 , n38003 );
or ( n38006 , n38001 , n38004 , n38005 );
and ( n38007 , n37991 , n38006 );
and ( n38008 , n37975 , n38007 );
and ( n38009 , n37951 , n38007 );
or ( n38010 , n37976 , n38008 , n38009 );
and ( n38011 , n37950 , n38010 );
xnor ( n38012 , n37834 , n37836 );
xnor ( n38013 , n37839 , n37841 );
and ( n38014 , n38012 , n38013 );
xor ( n38015 , n37852 , n37859 );
xor ( n38016 , n37868 , n37875 );
and ( n38017 , n38015 , n38016 );
and ( n38018 , n38014 , n38017 );
xor ( n38019 , n37890 , n37891 );
xor ( n38020 , n38019 , n37893 );
and ( n38021 , n38017 , n38020 );
and ( n38022 , n38014 , n38020 );
or ( n38023 , n38018 , n38021 , n38022 );
and ( n38024 , n38010 , n38023 );
and ( n38025 , n37950 , n38023 );
or ( n38026 , n38011 , n38024 , n38025 );
and ( n38027 , n37943 , n38026 );
xor ( n38028 , n37816 , n37818 );
xor ( n38029 , n38028 , n37825 );
xor ( n38030 , n37832 , n37843 );
xor ( n38031 , n38030 , n37877 );
and ( n38032 , n38029 , n38031 );
xor ( n38033 , n37883 , n37888 );
xor ( n38034 , n38033 , n37896 );
and ( n38035 , n38031 , n38034 );
and ( n38036 , n38029 , n38034 );
or ( n38037 , n38032 , n38035 , n38036 );
and ( n38038 , n38026 , n38037 );
and ( n38039 , n37943 , n38037 );
or ( n38040 , n38027 , n38038 , n38039 );
and ( n38041 , n37924 , n38040 );
xor ( n38042 , n37781 , n37783 );
xor ( n38043 , n38042 , n37785 );
xor ( n38044 , n37807 , n37810 );
xor ( n38045 , n38044 , n37828 );
and ( n38046 , n38043 , n38045 );
xor ( n38047 , n37880 , n37899 );
xor ( n38048 , n38047 , n37902 );
and ( n38049 , n38045 , n38048 );
and ( n38050 , n38043 , n38048 );
or ( n38051 , n38046 , n38049 , n38050 );
and ( n38052 , n38040 , n38051 );
and ( n38053 , n37924 , n38051 );
or ( n38054 , n38041 , n38052 , n38053 );
xor ( n38055 , n37761 , n37763 );
xor ( n38056 , n38055 , n37791 );
and ( n38057 , n38054 , n38056 );
xor ( n38058 , n37911 , n37913 );
xor ( n38059 , n38058 , n37916 );
and ( n38060 , n38056 , n38059 );
and ( n38061 , n38054 , n38059 );
or ( n38062 , n38057 , n38060 , n38061 );
and ( n38063 , n37921 , n38062 );
and ( n38064 , n37919 , n38062 );
or ( n38065 , n37922 , n38063 , n38064 );
xor ( n38066 , n37754 , n37797 );
xor ( n38067 , n38066 , n37800 );
and ( n38068 , n38065 , n38067 );
xor ( n38069 , n37756 , n37758 );
xor ( n38070 , n38069 , n37794 );
xor ( n38071 , n37919 , n37921 );
xor ( n38072 , n38071 , n38062 );
and ( n38073 , n38070 , n38072 );
xor ( n38074 , n37766 , n37767 );
xor ( n38075 , n38074 , n37788 );
xor ( n38076 , n37831 , n37905 );
xor ( n38077 , n38076 , n37908 );
and ( n38078 , n38075 , n38077 );
xor ( n38079 , n37953 , n37955 );
and ( n38080 , n32736 , n33296 );
and ( n38081 , n33339 , n32719 );
and ( n38082 , n38080 , n38081 );
buf ( n38083 , n15919 );
buf ( n38084 , n38083 );
and ( n38085 , n38082 , n38084 );
and ( n38086 , n38079 , n38085 );
and ( n38087 , n32057 , n33905 );
and ( n38088 , n33896 , n32066 );
and ( n38089 , n38087 , n38088 );
and ( n38090 , n38085 , n38089 );
and ( n38091 , n38079 , n38089 );
or ( n38092 , n38086 , n38090 , n38091 );
and ( n38093 , n32155 , n33905 );
and ( n38094 , n32365 , n33712 );
and ( n38095 , n38093 , n38094 );
and ( n38096 , n32689 , n33347 );
and ( n38097 , n38094 , n38096 );
and ( n38098 , n38093 , n38096 );
or ( n38099 , n38095 , n38097 , n38098 );
xor ( n38100 , n37992 , n37993 );
xor ( n38101 , n38100 , n37995 );
and ( n38102 , n38099 , n38101 );
xor ( n38103 , n37958 , n37959 );
xor ( n38104 , n38103 , n37961 );
and ( n38105 , n38101 , n38104 );
and ( n38106 , n38099 , n38104 );
or ( n38107 , n38102 , n38105 , n38106 );
and ( n38108 , n33896 , n32173 );
and ( n38109 , n33692 , n32348 );
and ( n38110 , n38108 , n38109 );
and ( n38111 , n33304 , n32671 );
and ( n38112 , n38109 , n38111 );
and ( n38113 , n38108 , n38111 );
or ( n38114 , n38110 , n38112 , n38113 );
xor ( n38115 , n37977 , n37978 );
xor ( n38116 , n38115 , n37980 );
and ( n38117 , n38114 , n38116 );
xor ( n38118 , n37965 , n37966 );
xor ( n38119 , n38118 , n37968 );
and ( n38120 , n38116 , n38119 );
and ( n38121 , n38114 , n38119 );
or ( n38122 , n38117 , n38120 , n38121 );
and ( n38123 , n38107 , n38122 );
and ( n38124 , n38092 , n38123 );
xor ( n38125 , n37952 , n37956 );
xor ( n38126 , n38125 , n37972 );
and ( n38127 , n38123 , n38126 );
and ( n38128 , n38092 , n38126 );
or ( n38129 , n38124 , n38127 , n38128 );
xor ( n38130 , n37820 , n37821 );
xor ( n38131 , n37991 , n38006 );
and ( n38132 , n38130 , n38131 );
xor ( n38133 , n38012 , n38013 );
and ( n38134 , n38131 , n38133 );
and ( n38135 , n38130 , n38133 );
or ( n38136 , n38132 , n38134 , n38135 );
and ( n38137 , n38129 , n38136 );
xor ( n38138 , n38015 , n38016 );
xor ( n38139 , n37983 , n37985 );
xor ( n38140 , n38139 , n37988 );
xor ( n38141 , n37998 , n38000 );
xor ( n38142 , n38141 , n38003 );
and ( n38143 , n38140 , n38142 );
and ( n38144 , n38138 , n38143 );
xor ( n38145 , n37930 , n37931 );
xor ( n38146 , n37964 , n37971 );
and ( n38147 , n38145 , n38146 );
and ( n38148 , n34280 , n31861 );
and ( n38149 , n34099 , n32066 );
or ( n38150 , n38148 , n38149 );
and ( n38151 , n31883 , n34253 );
and ( n38152 , n32057 , n34082 );
or ( n38153 , n38151 , n38152 );
and ( n38154 , n38150 , n38153 );
and ( n38155 , n38146 , n38154 );
and ( n38156 , n38145 , n38154 );
or ( n38157 , n38147 , n38155 , n38156 );
and ( n38158 , n38143 , n38157 );
and ( n38159 , n38138 , n38157 );
or ( n38160 , n38144 , n38158 , n38159 );
and ( n38161 , n38136 , n38160 );
and ( n38162 , n38129 , n38160 );
or ( n38163 , n38137 , n38161 , n38162 );
xor ( n38164 , n37929 , n37935 );
xor ( n38165 , n38164 , n37937 );
xor ( n38166 , n37944 , n37945 );
xor ( n38167 , n38166 , n37947 );
and ( n38168 , n38165 , n38167 );
xor ( n38169 , n37951 , n37975 );
xor ( n38170 , n38169 , n38007 );
and ( n38171 , n38167 , n38170 );
and ( n38172 , n38165 , n38170 );
or ( n38173 , n38168 , n38171 , n38172 );
and ( n38174 , n38163 , n38173 );
xor ( n38175 , n37926 , n37927 );
xor ( n38176 , n38175 , n37940 );
and ( n38177 , n38173 , n38176 );
and ( n38178 , n38163 , n38176 );
or ( n38179 , n38174 , n38177 , n38178 );
xor ( n38180 , n37943 , n38026 );
xor ( n38181 , n38180 , n38037 );
and ( n38182 , n38179 , n38181 );
xor ( n38183 , n38043 , n38045 );
xor ( n38184 , n38183 , n38048 );
and ( n38185 , n38181 , n38184 );
and ( n38186 , n38179 , n38184 );
or ( n38187 , n38182 , n38185 , n38186 );
and ( n38188 , n38077 , n38187 );
and ( n38189 , n38075 , n38187 );
or ( n38190 , n38078 , n38188 , n38189 );
xor ( n38191 , n38054 , n38056 );
xor ( n38192 , n38191 , n38059 );
and ( n38193 , n38190 , n38192 );
xor ( n38194 , n37924 , n38040 );
xor ( n38195 , n38194 , n38051 );
xor ( n38196 , n38075 , n38077 );
xor ( n38197 , n38196 , n38187 );
and ( n38198 , n38195 , n38197 );
xor ( n38199 , n37950 , n38010 );
xor ( n38200 , n38199 , n38023 );
xor ( n38201 , n38029 , n38031 );
xor ( n38202 , n38201 , n38034 );
and ( n38203 , n38200 , n38202 );
xor ( n38204 , n38014 , n38017 );
xor ( n38205 , n38204 , n38020 );
xor ( n38206 , n38092 , n38123 );
xor ( n38207 , n38206 , n38126 );
xor ( n38208 , n38079 , n38085 );
xor ( n38209 , n38208 , n38089 );
xor ( n38210 , n38107 , n38122 );
and ( n38211 , n38209 , n38210 );
xor ( n38212 , n38140 , n38142 );
and ( n38213 , n38210 , n38212 );
and ( n38214 , n38209 , n38212 );
or ( n38215 , n38211 , n38213 , n38214 );
and ( n38216 , n38207 , n38215 );
buf ( n38217 , n32949 );
buf ( n38218 , n15922 );
buf ( n38219 , n38218 );
and ( n38220 , n38217 , n38219 );
xnor ( n38221 , n38148 , n38149 );
xnor ( n38222 , n38151 , n38152 );
and ( n38223 , n38221 , n38222 );
or ( n38224 , n38220 , n38223 );
and ( n38225 , n32155 , n34082 );
and ( n38226 , n32365 , n33905 );
and ( n38227 , n38225 , n38226 );
and ( n38228 , n32689 , n33712 );
and ( n38229 , n38226 , n38228 );
and ( n38230 , n38225 , n38228 );
or ( n38231 , n38227 , n38229 , n38230 );
and ( n38232 , n32057 , n34253 );
and ( n38233 , n32736 , n33347 );
and ( n38234 , n38232 , n38233 );
and ( n38235 , n32949 , n33296 );
and ( n38236 , n38233 , n38235 );
and ( n38237 , n38232 , n38235 );
or ( n38238 , n38234 , n38236 , n38237 );
or ( n38239 , n38231 , n38238 );
and ( n38240 , n34099 , n32173 );
and ( n38241 , n33896 , n32348 );
and ( n38242 , n38240 , n38241 );
and ( n38243 , n33692 , n32671 );
and ( n38244 , n38241 , n38243 );
and ( n38245 , n38240 , n38243 );
or ( n38246 , n38242 , n38244 , n38245 );
and ( n38247 , n34280 , n32066 );
and ( n38248 , n33304 , n32719 );
and ( n38249 , n38247 , n38248 );
and ( n38250 , n33339 , n32932 );
and ( n38251 , n38248 , n38250 );
and ( n38252 , n38247 , n38250 );
or ( n38253 , n38249 , n38251 , n38252 );
or ( n38254 , n38246 , n38253 );
and ( n38255 , n38239 , n38254 );
and ( n38256 , n38224 , n38255 );
xor ( n38257 , n38087 , n38088 );
xor ( n38258 , n38082 , n38084 );
and ( n38259 , n38257 , n38258 );
xor ( n38260 , n38150 , n38153 );
and ( n38261 , n38258 , n38260 );
and ( n38262 , n38257 , n38260 );
or ( n38263 , n38259 , n38261 , n38262 );
and ( n38264 , n38255 , n38263 );
and ( n38265 , n38224 , n38263 );
or ( n38266 , n38256 , n38264 , n38265 );
and ( n38267 , n38215 , n38266 );
and ( n38268 , n38207 , n38266 );
or ( n38269 , n38216 , n38267 , n38268 );
and ( n38270 , n38205 , n38269 );
xor ( n38271 , n38129 , n38136 );
xor ( n38272 , n38271 , n38160 );
and ( n38273 , n38269 , n38272 );
and ( n38274 , n38205 , n38272 );
or ( n38275 , n38270 , n38273 , n38274 );
and ( n38276 , n38202 , n38275 );
and ( n38277 , n38200 , n38275 );
or ( n38278 , n38203 , n38276 , n38277 );
xor ( n38279 , n38179 , n38181 );
xor ( n38280 , n38279 , n38184 );
and ( n38281 , n38278 , n38280 );
xor ( n38282 , n38163 , n38173 );
xor ( n38283 , n38282 , n38176 );
xor ( n38284 , n38165 , n38167 );
xor ( n38285 , n38284 , n38170 );
xor ( n38286 , n38130 , n38131 );
xor ( n38287 , n38286 , n38133 );
xor ( n38288 , n38138 , n38143 );
xor ( n38289 , n38288 , n38157 );
and ( n38290 , n38287 , n38289 );
xnor ( n38291 , n38220 , n38223 );
xor ( n38292 , n38217 , n38219 );
and ( n38293 , n32949 , n33347 );
and ( n38294 , n33304 , n32932 );
and ( n38295 , n38293 , n38294 );
buf ( n38296 , n15925 );
buf ( n38297 , n38296 );
and ( n38298 , n38295 , n38297 );
and ( n38299 , n38292 , n38298 );
and ( n38300 , n34099 , n32348 );
and ( n38301 , n33896 , n32671 );
and ( n38302 , n38300 , n38301 );
and ( n38303 , n33692 , n32719 );
and ( n38304 , n38301 , n38303 );
and ( n38305 , n38300 , n38303 );
or ( n38306 , n38302 , n38304 , n38305 );
and ( n38307 , n32365 , n34082 );
and ( n38308 , n32689 , n33905 );
and ( n38309 , n38307 , n38308 );
and ( n38310 , n32736 , n33712 );
and ( n38311 , n38308 , n38310 );
and ( n38312 , n38307 , n38310 );
or ( n38313 , n38309 , n38311 , n38312 );
and ( n38314 , n38306 , n38313 );
and ( n38315 , n38298 , n38314 );
and ( n38316 , n38292 , n38314 );
or ( n38317 , n38299 , n38315 , n38316 );
and ( n38318 , n38291 , n38317 );
xor ( n38319 , n38108 , n38109 );
xor ( n38320 , n38319 , n38111 );
xor ( n38321 , n38093 , n38094 );
xor ( n38322 , n38321 , n38096 );
and ( n38323 , n38320 , n38322 );
and ( n38324 , n38317 , n38323 );
and ( n38325 , n38291 , n38323 );
or ( n38326 , n38318 , n38324 , n38325 );
xor ( n38327 , n38099 , n38101 );
xor ( n38328 , n38327 , n38104 );
xor ( n38329 , n38114 , n38116 );
xor ( n38330 , n38329 , n38119 );
and ( n38331 , n38328 , n38330 );
and ( n38332 , n38326 , n38331 );
and ( n38333 , n38289 , n38332 );
and ( n38334 , n38287 , n38332 );
or ( n38335 , n38290 , n38333 , n38334 );
and ( n38336 , n38285 , n38335 );
xor ( n38337 , n38205 , n38269 );
xor ( n38338 , n38337 , n38272 );
and ( n38339 , n38335 , n38338 );
and ( n38340 , n38285 , n38338 );
or ( n38341 , n38336 , n38339 , n38340 );
and ( n38342 , n38283 , n38341 );
xor ( n38343 , n38200 , n38202 );
xor ( n38344 , n38343 , n38275 );
and ( n38345 , n38341 , n38344 );
and ( n38346 , n38283 , n38344 );
or ( n38347 , n38342 , n38345 , n38346 );
and ( n38348 , n38280 , n38347 );
and ( n38349 , n38278 , n38347 );
or ( n38350 , n38281 , n38348 , n38349 );
and ( n38351 , n38197 , n38350 );
and ( n38352 , n38195 , n38350 );
or ( n38353 , n38198 , n38351 , n38352 );
and ( n38354 , n38192 , n38353 );
and ( n38355 , n38190 , n38353 );
or ( n38356 , n38193 , n38354 , n38355 );
and ( n38357 , n38072 , n38356 );
and ( n38358 , n38070 , n38356 );
or ( n38359 , n38073 , n38357 , n38358 );
and ( n38360 , n38067 , n38359 );
and ( n38361 , n38065 , n38359 );
or ( n38362 , n38068 , n38360 , n38361 );
and ( n38363 , n37805 , n38362 );
and ( n38364 , n37803 , n38362 );
or ( n38365 , n37806 , n38363 , n38364 );
and ( n38366 , n37752 , n38365 );
xor ( n38367 , n37752 , n38365 );
xor ( n38368 , n37803 , n37805 );
xor ( n38369 , n38368 , n38362 );
xor ( n38370 , n38065 , n38067 );
xor ( n38371 , n38370 , n38359 );
not ( n38372 , n38371 );
xor ( n38373 , n38070 , n38072 );
xor ( n38374 , n38373 , n38356 );
not ( n38375 , n38374 );
xor ( n38376 , n38190 , n38192 );
xor ( n38377 , n38376 , n38353 );
xor ( n38378 , n38195 , n38197 );
xor ( n38379 , n38378 , n38350 );
xor ( n38380 , n38278 , n38280 );
xor ( n38381 , n38380 , n38347 );
xor ( n38382 , n38283 , n38341 );
xor ( n38383 , n38382 , n38344 );
xor ( n38384 , n38145 , n38146 );
xor ( n38385 , n38384 , n38154 );
xor ( n38386 , n38239 , n38254 );
xor ( n38387 , n38328 , n38330 );
and ( n38388 , n38386 , n38387 );
xor ( n38389 , n38225 , n38226 );
xor ( n38390 , n38389 , n38228 );
xor ( n38391 , n38232 , n38233 );
xor ( n38392 , n38391 , n38235 );
or ( n38393 , n38390 , n38392 );
xor ( n38394 , n38240 , n38241 );
xor ( n38395 , n38394 , n38243 );
xor ( n38396 , n38247 , n38248 );
xor ( n38397 , n38396 , n38250 );
or ( n38398 , n38395 , n38397 );
and ( n38399 , n38393 , n38398 );
and ( n38400 , n38387 , n38399 );
and ( n38401 , n38386 , n38399 );
or ( n38402 , n38388 , n38400 , n38401 );
and ( n38403 , n38385 , n38402 );
xnor ( n38404 , n38231 , n38238 );
xnor ( n38405 , n38246 , n38253 );
and ( n38406 , n38404 , n38405 );
xor ( n38407 , n38080 , n38081 );
xor ( n38408 , n38320 , n38322 );
and ( n38409 , n38407 , n38408 );
xor ( n38410 , n38221 , n38222 );
and ( n38411 , n38408 , n38410 );
and ( n38412 , n38407 , n38410 );
or ( n38413 , n38409 , n38411 , n38412 );
and ( n38414 , n38406 , n38413 );
xor ( n38415 , n38257 , n38258 );
xor ( n38416 , n38415 , n38260 );
and ( n38417 , n38413 , n38416 );
and ( n38418 , n38406 , n38416 );
or ( n38419 , n38414 , n38417 , n38418 );
and ( n38420 , n38402 , n38419 );
and ( n38421 , n38385 , n38419 );
or ( n38422 , n38403 , n38420 , n38421 );
xor ( n38423 , n38207 , n38215 );
xor ( n38424 , n38423 , n38266 );
and ( n38425 , n38422 , n38424 );
xor ( n38426 , n38209 , n38210 );
xor ( n38427 , n38426 , n38212 );
xor ( n38428 , n38224 , n38255 );
xor ( n38429 , n38428 , n38263 );
and ( n38430 , n38427 , n38429 );
xor ( n38431 , n38326 , n38331 );
and ( n38432 , n38429 , n38431 );
and ( n38433 , n38427 , n38431 );
or ( n38434 , n38430 , n38432 , n38433 );
and ( n38435 , n38424 , n38434 );
and ( n38436 , n38422 , n38434 );
or ( n38437 , n38425 , n38435 , n38436 );
xor ( n38438 , n38285 , n38335 );
xor ( n38439 , n38438 , n38338 );
and ( n38440 , n38437 , n38439 );
xor ( n38441 , n38287 , n38289 );
xor ( n38442 , n38441 , n38332 );
xor ( n38443 , n38291 , n38317 );
xor ( n38444 , n38443 , n38323 );
xor ( n38445 , n38292 , n38298 );
xor ( n38446 , n38445 , n38314 );
xor ( n38447 , n38393 , n38398 );
and ( n38448 , n38446 , n38447 );
xor ( n38449 , n38404 , n38405 );
and ( n38450 , n38447 , n38449 );
and ( n38451 , n38446 , n38449 );
or ( n38452 , n38448 , n38450 , n38451 );
and ( n38453 , n38444 , n38452 );
xor ( n38454 , n38295 , n38297 );
buf ( n38455 , n33339 );
buf ( n38456 , n15928 );
buf ( n38457 , n38456 );
and ( n38458 , n38455 , n38457 );
and ( n38459 , n38454 , n38458 );
and ( n38460 , n32155 , n34253 );
and ( n38461 , n34280 , n32173 );
and ( n38462 , n38460 , n38461 );
and ( n38463 , n38458 , n38462 );
and ( n38464 , n38454 , n38462 );
or ( n38465 , n38459 , n38463 , n38464 );
and ( n38466 , n32736 , n33905 );
and ( n38467 , n32949 , n33712 );
and ( n38468 , n38466 , n38467 );
and ( n38469 , n33339 , n33347 );
and ( n38470 , n38467 , n38469 );
and ( n38471 , n38466 , n38469 );
or ( n38472 , n38468 , n38470 , n38471 );
xor ( n38473 , n38307 , n38308 );
xor ( n38474 , n38473 , n38310 );
or ( n38475 , n38472 , n38474 );
and ( n38476 , n33896 , n32719 );
and ( n38477 , n33692 , n32932 );
and ( n38478 , n38476 , n38477 );
and ( n38479 , n33304 , n33296 );
and ( n38480 , n38477 , n38479 );
and ( n38481 , n38476 , n38479 );
or ( n38482 , n38478 , n38480 , n38481 );
xor ( n38483 , n38300 , n38301 );
xor ( n38484 , n38483 , n38303 );
or ( n38485 , n38482 , n38484 );
and ( n38486 , n38475 , n38485 );
and ( n38487 , n38465 , n38486 );
xnor ( n38488 , n38390 , n38392 );
xnor ( n38489 , n38395 , n38397 );
and ( n38490 , n38488 , n38489 );
and ( n38491 , n38486 , n38490 );
and ( n38492 , n38465 , n38490 );
or ( n38493 , n38487 , n38491 , n38492 );
and ( n38494 , n38452 , n38493 );
and ( n38495 , n38444 , n38493 );
or ( n38496 , n38453 , n38494 , n38495 );
xor ( n38497 , n38385 , n38402 );
xor ( n38498 , n38497 , n38419 );
and ( n38499 , n38496 , n38498 );
xor ( n38500 , n38386 , n38387 );
xor ( n38501 , n38500 , n38399 );
xor ( n38502 , n38406 , n38413 );
xor ( n38503 , n38502 , n38416 );
and ( n38504 , n38501 , n38503 );
xor ( n38505 , n38407 , n38408 );
xor ( n38506 , n38505 , n38410 );
xor ( n38507 , n38306 , n38313 );
and ( n38508 , n34280 , n32348 );
and ( n38509 , n34099 , n32671 );
and ( n38510 , n38508 , n38509 );
and ( n38511 , n32365 , n34253 );
and ( n38512 , n32689 , n34082 );
and ( n38513 , n38511 , n38512 );
and ( n38514 , n38510 , n38513 );
and ( n38515 , n38507 , n38514 );
xor ( n38516 , n38454 , n38458 );
xor ( n38517 , n38516 , n38462 );
and ( n38518 , n38514 , n38517 );
and ( n38519 , n38507 , n38517 );
or ( n38520 , n38515 , n38518 , n38519 );
and ( n38521 , n38506 , n38520 );
xor ( n38522 , n38475 , n38485 );
xor ( n38523 , n38488 , n38489 );
and ( n38524 , n38522 , n38523 );
and ( n38525 , n33339 , n33712 );
and ( n38526 , n33692 , n33296 );
and ( n38527 , n38525 , n38526 );
buf ( n38528 , n15931 );
buf ( n38529 , n38528 );
and ( n38530 , n38527 , n38529 );
and ( n38531 , n34280 , n32671 );
and ( n38532 , n34099 , n32719 );
and ( n38533 , n38531 , n38532 );
and ( n38534 , n33896 , n32932 );
and ( n38535 , n38532 , n38534 );
and ( n38536 , n38531 , n38534 );
or ( n38537 , n38533 , n38535 , n38536 );
and ( n38538 , n32689 , n34253 );
and ( n38539 , n32736 , n34082 );
and ( n38540 , n38538 , n38539 );
and ( n38541 , n32949 , n33905 );
and ( n38542 , n38539 , n38541 );
and ( n38543 , n38538 , n38541 );
or ( n38544 , n38540 , n38542 , n38543 );
and ( n38545 , n38537 , n38544 );
or ( n38546 , n38530 , n38545 );
and ( n38547 , n38523 , n38546 );
and ( n38548 , n38522 , n38546 );
or ( n38549 , n38524 , n38547 , n38548 );
and ( n38550 , n38520 , n38549 );
and ( n38551 , n38506 , n38549 );
or ( n38552 , n38521 , n38550 , n38551 );
and ( n38553 , n38503 , n38552 );
and ( n38554 , n38501 , n38552 );
or ( n38555 , n38504 , n38553 , n38554 );
and ( n38556 , n38498 , n38555 );
and ( n38557 , n38496 , n38555 );
or ( n38558 , n38499 , n38556 , n38557 );
and ( n38559 , n38442 , n38558 );
xor ( n38560 , n38422 , n38424 );
xor ( n38561 , n38560 , n38434 );
and ( n38562 , n38558 , n38561 );
and ( n38563 , n38442 , n38561 );
or ( n38564 , n38559 , n38562 , n38563 );
and ( n38565 , n38439 , n38564 );
and ( n38566 , n38437 , n38564 );
or ( n38567 , n38440 , n38565 , n38566 );
and ( n38568 , n38383 , n38567 );
xor ( n38569 , n38437 , n38439 );
xor ( n38570 , n38569 , n38564 );
xor ( n38571 , n38427 , n38429 );
xor ( n38572 , n38571 , n38431 );
xor ( n38573 , n38508 , n38509 );
xor ( n38574 , n38511 , n38512 );
and ( n38575 , n38573 , n38574 );
xor ( n38576 , n38455 , n38457 );
and ( n38577 , n38575 , n38576 );
xnor ( n38578 , n38472 , n38474 );
xnor ( n38579 , n38482 , n38484 );
and ( n38580 , n38578 , n38579 );
and ( n38581 , n38577 , n38580 );
xor ( n38582 , n38460 , n38461 );
xor ( n38583 , n38293 , n38294 );
and ( n38584 , n38582 , n38583 );
xor ( n38585 , n38510 , n38513 );
and ( n38586 , n38583 , n38585 );
and ( n38587 , n38582 , n38585 );
or ( n38588 , n38584 , n38586 , n38587 );
and ( n38589 , n38580 , n38588 );
and ( n38590 , n38577 , n38588 );
or ( n38591 , n38581 , n38589 , n38590 );
xor ( n38592 , n38446 , n38447 );
xor ( n38593 , n38592 , n38449 );
and ( n38594 , n38591 , n38593 );
xor ( n38595 , n38465 , n38486 );
xor ( n38596 , n38595 , n38490 );
and ( n38597 , n38593 , n38596 );
and ( n38598 , n38591 , n38596 );
or ( n38599 , n38594 , n38597 , n38598 );
xor ( n38600 , n38444 , n38452 );
xor ( n38601 , n38600 , n38493 );
and ( n38602 , n38599 , n38601 );
xnor ( n38603 , n38530 , n38545 );
xor ( n38604 , n38575 , n38576 );
or ( n38605 , n38603 , n38604 );
xor ( n38606 , n38578 , n38579 );
xor ( n38607 , n38537 , n38544 );
xor ( n38608 , n38476 , n38477 );
xor ( n38609 , n38608 , n38479 );
xor ( n38610 , n38466 , n38467 );
xor ( n38611 , n38610 , n38469 );
xor ( n38612 , n38609 , n38611 );
and ( n38613 , n38607 , n38612 );
xor ( n38614 , n38573 , n38574 );
and ( n38615 , n38612 , n38614 );
and ( n38616 , n38607 , n38614 );
or ( n38617 , n38613 , n38615 , n38616 );
and ( n38618 , n38606 , n38617 );
xor ( n38619 , n38582 , n38583 );
xor ( n38620 , n38619 , n38585 );
and ( n38621 , n38617 , n38620 );
and ( n38622 , n38606 , n38620 );
or ( n38623 , n38618 , n38621 , n38622 );
and ( n38624 , n38605 , n38623 );
xor ( n38625 , n38507 , n38514 );
xor ( n38626 , n38625 , n38517 );
and ( n38627 , n38623 , n38626 );
and ( n38628 , n38605 , n38626 );
or ( n38629 , n38624 , n38627 , n38628 );
xor ( n38630 , n38506 , n38520 );
xor ( n38631 , n38630 , n38549 );
and ( n38632 , n38629 , n38631 );
xor ( n38633 , n38591 , n38593 );
xor ( n38634 , n38633 , n38596 );
and ( n38635 , n38631 , n38634 );
and ( n38636 , n38629 , n38634 );
or ( n38637 , n38632 , n38635 , n38636 );
and ( n38638 , n38601 , n38637 );
and ( n38639 , n38599 , n38637 );
or ( n38640 , n38602 , n38638 , n38639 );
and ( n38641 , n38572 , n38640 );
xor ( n38642 , n38496 , n38498 );
xor ( n38643 , n38642 , n38555 );
and ( n38644 , n38640 , n38643 );
and ( n38645 , n38572 , n38643 );
or ( n38646 , n38641 , n38644 , n38645 );
xor ( n38647 , n38442 , n38558 );
xor ( n38648 , n38647 , n38561 );
and ( n38649 , n38646 , n38648 );
xor ( n38650 , n38572 , n38640 );
xor ( n38651 , n38650 , n38643 );
xor ( n38652 , n38501 , n38503 );
xor ( n38653 , n38652 , n38552 );
xor ( n38654 , n38599 , n38601 );
xor ( n38655 , n38654 , n38637 );
and ( n38656 , n38653 , n38655 );
xor ( n38657 , n38522 , n38523 );
xor ( n38658 , n38657 , n38546 );
xor ( n38659 , n38577 , n38580 );
xor ( n38660 , n38659 , n38588 );
and ( n38661 , n38658 , n38660 );
xnor ( n38662 , n38603 , n38604 );
xor ( n38663 , n38527 , n38529 );
buf ( n38664 , n33304 );
buf ( n38665 , n15934 );
buf ( n38666 , n38665 );
and ( n38667 , n38664 , n38666 );
and ( n38668 , n38663 , n38667 );
and ( n38669 , n34099 , n32932 );
and ( n38670 , n33896 , n33296 );
and ( n38671 , n38669 , n38670 );
and ( n38672 , n33692 , n33347 );
and ( n38673 , n38670 , n38672 );
and ( n38674 , n38669 , n38672 );
or ( n38675 , n38671 , n38673 , n38674 );
and ( n38676 , n32949 , n34082 );
and ( n38677 , n33339 , n33905 );
and ( n38678 , n38676 , n38677 );
and ( n38679 , n33304 , n33712 );
and ( n38680 , n38677 , n38679 );
and ( n38681 , n38676 , n38679 );
or ( n38682 , n38678 , n38680 , n38681 );
and ( n38683 , n38675 , n38682 );
and ( n38684 , n38667 , n38683 );
and ( n38685 , n38663 , n38683 );
or ( n38686 , n38668 , n38684 , n38685 );
and ( n38687 , n38662 , n38686 );
and ( n38688 , n38609 , n38611 );
and ( n38689 , n38686 , n38688 );
and ( n38690 , n38662 , n38688 );
or ( n38691 , n38687 , n38689 , n38690 );
and ( n38692 , n38660 , n38691 );
and ( n38693 , n38658 , n38691 );
or ( n38694 , n38661 , n38692 , n38693 );
xor ( n38695 , n38629 , n38631 );
xor ( n38696 , n38695 , n38634 );
and ( n38697 , n38694 , n38696 );
xor ( n38698 , n38531 , n38532 );
xor ( n38699 , n38698 , n38534 );
xor ( n38700 , n38538 , n38539 );
xor ( n38701 , n38700 , n38541 );
and ( n38702 , n38699 , n38701 );
xor ( n38703 , n38664 , n38666 );
xor ( n38704 , n38525 , n38526 );
and ( n38705 , n38703 , n38704 );
and ( n38706 , n32736 , n34253 );
and ( n38707 , n34280 , n32719 );
and ( n38708 , n38706 , n38707 );
and ( n38709 , n38704 , n38708 );
and ( n38710 , n38703 , n38708 );
or ( n38711 , n38705 , n38709 , n38710 );
and ( n38712 , n38702 , n38711 );
xor ( n38713 , n38663 , n38667 );
xor ( n38714 , n38713 , n38683 );
and ( n38715 , n38711 , n38714 );
and ( n38716 , n38702 , n38714 );
or ( n38717 , n38712 , n38715 , n38716 );
xor ( n38718 , n38675 , n38682 );
xor ( n38719 , n38699 , n38701 );
and ( n38720 , n38718 , n38719 );
and ( n38721 , n33304 , n33905 );
and ( n38722 , n33896 , n33347 );
and ( n38723 , n38721 , n38722 );
buf ( n38724 , n15937 );
buf ( n38725 , n38724 );
or ( n38726 , n38723 , n38725 );
and ( n38727 , n38719 , n38726 );
and ( n38728 , n38718 , n38726 );
or ( n38729 , n38720 , n38727 , n38728 );
xnor ( n38730 , n38723 , n38725 );
buf ( n38731 , n38730 );
and ( n38732 , n34280 , n32932 );
and ( n38733 , n34099 , n33296 );
and ( n38734 , n38732 , n38733 );
and ( n38735 , n32949 , n34253 );
and ( n38736 , n33339 , n34082 );
and ( n38737 , n38735 , n38736 );
and ( n38738 , n38734 , n38737 );
and ( n38739 , n38731 , n38738 );
xor ( n38740 , n38669 , n38670 );
xor ( n38741 , n38740 , n38672 );
xor ( n38742 , n38676 , n38677 );
xor ( n38743 , n38742 , n38679 );
and ( n38744 , n38741 , n38743 );
and ( n38745 , n38738 , n38744 );
and ( n38746 , n38731 , n38744 );
or ( n38747 , n38739 , n38745 , n38746 );
and ( n38748 , n38729 , n38747 );
xor ( n38749 , n38607 , n38612 );
xor ( n38750 , n38749 , n38614 );
and ( n38751 , n38747 , n38750 );
and ( n38752 , n38729 , n38750 );
or ( n38753 , n38748 , n38751 , n38752 );
and ( n38754 , n38717 , n38753 );
xor ( n38755 , n38606 , n38617 );
xor ( n38756 , n38755 , n38620 );
and ( n38757 , n38753 , n38756 );
and ( n38758 , n38717 , n38756 );
or ( n38759 , n38754 , n38757 , n38758 );
xor ( n38760 , n38605 , n38623 );
xor ( n38761 , n38760 , n38626 );
and ( n38762 , n38759 , n38761 );
xor ( n38763 , n38662 , n38686 );
xor ( n38764 , n38763 , n38688 );
xor ( n38765 , n38703 , n38704 );
xor ( n38766 , n38765 , n38708 );
buf ( n38767 , n33692 );
buf ( n38768 , n15940 );
buf ( n38769 , n38768 );
and ( n38770 , n38767 , n38769 );
xor ( n38771 , n38732 , n38733 );
xor ( n38772 , n38735 , n38736 );
and ( n38773 , n38771 , n38772 );
and ( n38774 , n38770 , n38773 );
and ( n38775 , n38766 , n38774 );
xor ( n38776 , n38706 , n38707 );
xor ( n38777 , n38734 , n38737 );
and ( n38778 , n38776 , n38777 );
xor ( n38779 , n38741 , n38743 );
and ( n38780 , n38777 , n38779 );
and ( n38781 , n38776 , n38779 );
or ( n38782 , n38778 , n38780 , n38781 );
and ( n38783 , n38774 , n38782 );
and ( n38784 , n38766 , n38782 );
or ( n38785 , n38775 , n38783 , n38784 );
xor ( n38786 , n38702 , n38711 );
xor ( n38787 , n38786 , n38714 );
and ( n38788 , n38785 , n38787 );
xor ( n38789 , n38729 , n38747 );
xor ( n38790 , n38789 , n38750 );
and ( n38791 , n38787 , n38790 );
and ( n38792 , n38785 , n38790 );
or ( n38793 , n38788 , n38791 , n38792 );
and ( n38794 , n38764 , n38793 );
xor ( n38795 , n38717 , n38753 );
xor ( n38796 , n38795 , n38756 );
and ( n38797 , n38793 , n38796 );
and ( n38798 , n38764 , n38796 );
or ( n38799 , n38794 , n38797 , n38798 );
and ( n38800 , n38761 , n38799 );
and ( n38801 , n38759 , n38799 );
or ( n38802 , n38762 , n38800 , n38801 );
and ( n38803 , n38696 , n38802 );
and ( n38804 , n38694 , n38802 );
or ( n38805 , n38697 , n38803 , n38804 );
and ( n38806 , n38655 , n38805 );
and ( n38807 , n38653 , n38805 );
or ( n38808 , n38656 , n38806 , n38807 );
and ( n38809 , n38651 , n38808 );
xor ( n38810 , n38653 , n38655 );
xor ( n38811 , n38810 , n38805 );
xor ( n38812 , n38694 , n38696 );
xor ( n38813 , n38812 , n38802 );
xor ( n38814 , n38658 , n38660 );
xor ( n38815 , n38814 , n38691 );
xor ( n38816 , n38759 , n38761 );
xor ( n38817 , n38816 , n38799 );
and ( n38818 , n38815 , n38817 );
xor ( n38819 , n38764 , n38793 );
xor ( n38820 , n38819 , n38796 );
xor ( n38821 , n38718 , n38719 );
xor ( n38822 , n38821 , n38726 );
xor ( n38823 , n38731 , n38738 );
xor ( n38824 , n38823 , n38744 );
and ( n38825 , n38822 , n38824 );
xor ( n38826 , n38770 , n38773 );
not ( n38827 , n38730 );
and ( n38828 , n38826 , n38827 );
and ( n38829 , n34280 , n33296 );
and ( n38830 , n34099 , n33347 );
and ( n38831 , n38829 , n38830 );
and ( n38832 , n33896 , n33712 );
and ( n38833 , n38830 , n38832 );
and ( n38834 , n38829 , n38832 );
or ( n38835 , n38831 , n38833 , n38834 );
and ( n38836 , n33339 , n34253 );
and ( n38837 , n33304 , n34082 );
and ( n38838 , n38836 , n38837 );
and ( n38839 , n33692 , n33905 );
and ( n38840 , n38837 , n38839 );
and ( n38841 , n38836 , n38839 );
or ( n38842 , n38838 , n38840 , n38841 );
and ( n38843 , n38835 , n38842 );
and ( n38844 , n38827 , n38843 );
and ( n38845 , n38826 , n38843 );
or ( n38846 , n38828 , n38844 , n38845 );
and ( n38847 , n38824 , n38846 );
and ( n38848 , n38822 , n38846 );
or ( n38849 , n38825 , n38847 , n38848 );
xor ( n38850 , n38785 , n38787 );
xor ( n38851 , n38850 , n38790 );
and ( n38852 , n38849 , n38851 );
xor ( n38853 , n38767 , n38769 );
xor ( n38854 , n38721 , n38722 );
and ( n38855 , n38853 , n38854 );
xor ( n38856 , n38835 , n38842 );
and ( n38857 , n38854 , n38856 );
and ( n38858 , n38853 , n38856 );
or ( n38859 , n38855 , n38857 , n38858 );
xor ( n38860 , n38771 , n38772 );
buf ( n38861 , n33896 );
buf ( n38862 , n15946 );
buf ( n38863 , n38862 );
and ( n38864 , n38861 , n38863 );
and ( n38865 , n33304 , n34253 );
and ( n38866 , n34280 , n33347 );
and ( n38867 , n38865 , n38866 );
and ( n38868 , n38864 , n38867 );
and ( n38869 , n38860 , n38868 );
xor ( n38870 , n38829 , n38830 );
xor ( n38871 , n38870 , n38832 );
xor ( n38872 , n38836 , n38837 );
xor ( n38873 , n38872 , n38839 );
and ( n38874 , n38871 , n38873 );
and ( n38875 , n38868 , n38874 );
and ( n38876 , n38860 , n38874 );
or ( n38877 , n38869 , n38875 , n38876 );
and ( n38878 , n38859 , n38877 );
xor ( n38879 , n38776 , n38777 );
xor ( n38880 , n38879 , n38779 );
and ( n38881 , n38877 , n38880 );
and ( n38882 , n38859 , n38880 );
or ( n38883 , n38878 , n38881 , n38882 );
xor ( n38884 , n38766 , n38774 );
xor ( n38885 , n38884 , n38782 );
and ( n38886 , n38883 , n38885 );
xor ( n38887 , n38826 , n38827 );
xor ( n38888 , n38887 , n38843 );
buf ( n38889 , n15943 );
buf ( n38890 , n38889 );
and ( n38891 , n33692 , n34082 );
and ( n38892 , n34099 , n33712 );
and ( n38893 , n38891 , n38892 );
and ( n38894 , n38890 , n38893 );
xor ( n38895 , n38864 , n38867 );
and ( n38896 , n38893 , n38895 );
and ( n38897 , n38890 , n38895 );
or ( n38898 , n38894 , n38896 , n38897 );
xor ( n38899 , n38853 , n38854 );
xor ( n38900 , n38899 , n38856 );
and ( n38901 , n38898 , n38900 );
xor ( n38902 , n38860 , n38868 );
xor ( n38903 , n38902 , n38874 );
and ( n38904 , n38900 , n38903 );
and ( n38905 , n38898 , n38903 );
or ( n38906 , n38901 , n38904 , n38905 );
and ( n38907 , n38888 , n38906 );
xor ( n38908 , n38859 , n38877 );
xor ( n38909 , n38908 , n38880 );
and ( n38910 , n38906 , n38909 );
and ( n38911 , n38888 , n38909 );
or ( n38912 , n38907 , n38910 , n38911 );
and ( n38913 , n38885 , n38912 );
and ( n38914 , n38883 , n38912 );
or ( n38915 , n38886 , n38913 , n38914 );
and ( n38916 , n38851 , n38915 );
and ( n38917 , n38849 , n38915 );
or ( n38918 , n38852 , n38916 , n38917 );
and ( n38919 , n38820 , n38918 );
xor ( n38920 , n38849 , n38851 );
xor ( n38921 , n38920 , n38915 );
xor ( n38922 , n38822 , n38824 );
xor ( n38923 , n38922 , n38846 );
xor ( n38924 , n38883 , n38885 );
xor ( n38925 , n38924 , n38912 );
and ( n38926 , n38923 , n38925 );
xor ( n38927 , n38888 , n38906 );
xor ( n38928 , n38927 , n38909 );
xor ( n38929 , n38871 , n38873 );
and ( n38930 , n34280 , n33712 );
and ( n38931 , n34099 , n33905 );
or ( n38932 , n38930 , n38931 );
and ( n38933 , n33692 , n34253 );
and ( n38934 , n33896 , n34082 );
or ( n38935 , n38933 , n38934 );
and ( n38936 , n38932 , n38935 );
and ( n38937 , n38929 , n38936 );
xnor ( n38938 , n38930 , n38931 );
xnor ( n38939 , n38933 , n38934 );
and ( n38940 , n38938 , n38939 );
xor ( n38941 , n38861 , n38863 );
or ( n38942 , n38940 , n38941 );
and ( n38943 , n38936 , n38942 );
and ( n38944 , n38929 , n38942 );
or ( n38945 , n38937 , n38943 , n38944 );
xor ( n38946 , n38898 , n38900 );
xor ( n38947 , n38946 , n38903 );
and ( n38948 , n38945 , n38947 );
xor ( n38949 , n38865 , n38866 );
xor ( n38950 , n38891 , n38892 );
and ( n38951 , n38949 , n38950 );
xor ( n38952 , n38932 , n38935 );
and ( n38953 , n38950 , n38952 );
and ( n38954 , n38949 , n38952 );
or ( n38955 , n38951 , n38953 , n38954 );
xor ( n38956 , n38890 , n38893 );
xor ( n38957 , n38956 , n38895 );
and ( n38958 , n38955 , n38957 );
and ( n38959 , n33896 , n34253 );
and ( n38960 , n34280 , n33905 );
and ( n38961 , n38959 , n38960 );
buf ( n38962 , n15949 );
buf ( n38963 , n38962 );
and ( n38964 , n38961 , n38963 );
xnor ( n38965 , n38940 , n38941 );
or ( n38966 , n38964 , n38965 );
and ( n38967 , n38957 , n38966 );
and ( n38968 , n38955 , n38966 );
or ( n38969 , n38958 , n38967 , n38968 );
and ( n38970 , n38947 , n38969 );
and ( n38971 , n38945 , n38969 );
or ( n38972 , n38948 , n38970 , n38971 );
and ( n38973 , n38928 , n38972 );
xor ( n38974 , n38929 , n38936 );
xor ( n38975 , n38974 , n38942 );
buf ( n38976 , n34099 );
buf ( n38977 , n15952 );
buf ( n38978 , n38977 );
and ( n38979 , n38976 , n38978 );
xor ( n38980 , n38961 , n38963 );
or ( n38981 , n38979 , n38980 );
xor ( n38982 , n38949 , n38950 );
xor ( n38983 , n38982 , n38952 );
and ( n38984 , n38981 , n38983 );
xnor ( n38985 , n38964 , n38965 );
and ( n38986 , n38983 , n38985 );
and ( n38987 , n38981 , n38985 );
or ( n38988 , n38984 , n38986 , n38987 );
and ( n38989 , n38975 , n38988 );
xor ( n38990 , n38955 , n38957 );
xor ( n38991 , n38990 , n38966 );
and ( n38992 , n38988 , n38991 );
and ( n38993 , n38975 , n38991 );
or ( n38994 , n38989 , n38992 , n38993 );
xor ( n38995 , n38945 , n38947 );
xor ( n38996 , n38995 , n38969 );
or ( n38997 , n38994 , n38996 );
and ( n38998 , n38972 , n38997 );
and ( n38999 , n38928 , n38997 );
or ( n39000 , n38973 , n38998 , n38999 );
and ( n39001 , n38925 , n39000 );
and ( n39002 , n38923 , n39000 );
or ( n39003 , n38926 , n39001 , n39002 );
or ( n39004 , n38921 , n39003 );
and ( n39005 , n38918 , n39004 );
and ( n39006 , n38820 , n39004 );
or ( n39007 , n38919 , n39005 , n39006 );
and ( n39008 , n38817 , n39007 );
and ( n39009 , n38815 , n39007 );
or ( n39010 , n38818 , n39008 , n39009 );
or ( n39011 , n38813 , n39010 );
or ( n39012 , n38811 , n39011 );
and ( n39013 , n38808 , n39012 );
and ( n39014 , n38651 , n39012 );
or ( n39015 , n38809 , n39013 , n39014 );
and ( n39016 , n38648 , n39015 );
and ( n39017 , n38646 , n39015 );
or ( n39018 , n38649 , n39016 , n39017 );
or ( n39019 , n38570 , n39018 );
and ( n39020 , n38567 , n39019 );
and ( n39021 , n38383 , n39019 );
or ( n39022 , n38568 , n39020 , n39021 );
or ( n39023 , n38381 , n39022 );
and ( n39024 , n38379 , n39023 );
xor ( n39025 , n38379 , n39023 );
xnor ( n39026 , n38381 , n39022 );
xor ( n39027 , n38383 , n38567 );
xor ( n39028 , n39027 , n39019 );
not ( n39029 , n39028 );
xnor ( n39030 , n38570 , n39018 );
xor ( n39031 , n38646 , n38648 );
xor ( n39032 , n39031 , n39015 );
xor ( n39033 , n38651 , n38808 );
xor ( n39034 , n39033 , n39012 );
not ( n39035 , n39034 );
xnor ( n39036 , n38811 , n39011 );
xnor ( n39037 , n38813 , n39010 );
xor ( n39038 , n38815 , n38817 );
xor ( n39039 , n39038 , n39007 );
not ( n39040 , n39039 );
xor ( n39041 , n38820 , n38918 );
xor ( n39042 , n39041 , n39004 );
not ( n39043 , n39042 );
xnor ( n39044 , n38921 , n39003 );
xor ( n39045 , n38923 , n38925 );
xor ( n39046 , n39045 , n39000 );
xor ( n39047 , n38928 , n38972 );
xor ( n39048 , n39047 , n38997 );
not ( n39049 , n39048 );
xnor ( n39050 , n38994 , n38996 );
xor ( n39051 , n38975 , n38988 );
xor ( n39052 , n39051 , n38991 );
xor ( n39053 , n38938 , n38939 );
and ( n39054 , n34099 , n34253 );
and ( n39055 , n34280 , n34082 );
and ( n39056 , n39054 , n39055 );
xor ( n39057 , n38976 , n38978 );
or ( n39058 , n39056 , n39057 );
and ( n39059 , n39053 , n39058 );
xnor ( n39060 , n38979 , n38980 );
and ( n39061 , n39058 , n39060 );
and ( n39062 , n39053 , n39060 );
or ( n39063 , n39059 , n39061 , n39062 );
xor ( n39064 , n38981 , n38983 );
xor ( n39065 , n39064 , n38985 );
and ( n39066 , n39063 , n39065 );
xor ( n39067 , n39063 , n39065 );
xor ( n39068 , n38959 , n38960 );
xnor ( n39069 , n39056 , n39057 );
or ( n39070 , n39068 , n39069 );
xor ( n39071 , n39053 , n39058 );
xor ( n39072 , n39071 , n39060 );
and ( n39073 , n39070 , n39072 );
xor ( n39074 , n39070 , n39072 );
xnor ( n39075 , n39068 , n39069 );
buf ( n39076 , n15955 );
buf ( n39077 , n39076 );
xor ( n39078 , n39054 , n39055 );
and ( n39079 , n39077 , n39078 );
xor ( n39080 , n39077 , n39078 );
buf ( n39081 , n34280 );
buf ( n39082 , n15958 );
buf ( n39083 , n39082 );
and ( n39084 , n39081 , n39083 );
and ( n39085 , n39080 , n39084 );
or ( n39086 , n39079 , n39085 );
and ( n39087 , n39075 , n39086 );
and ( n39088 , n39074 , n39087 );
or ( n39089 , n39073 , n39088 );
and ( n39090 , n39067 , n39089 );
or ( n39091 , n39066 , n39090 );
and ( n39092 , n39052 , n39091 );
and ( n39093 , n39050 , n39092 );
and ( n39094 , n39049 , n39093 );
or ( n39095 , n39048 , n39094 );
and ( n39096 , n39046 , n39095 );
and ( n39097 , n39044 , n39096 );
and ( n39098 , n39043 , n39097 );
or ( n39099 , n39042 , n39098 );
and ( n39100 , n39040 , n39099 );
or ( n39101 , n39039 , n39100 );
and ( n39102 , n39037 , n39101 );
and ( n39103 , n39036 , n39102 );
and ( n39104 , n39035 , n39103 );
or ( n39105 , n39034 , n39104 );
and ( n39106 , n39032 , n39105 );
and ( n39107 , n39030 , n39106 );
and ( n39108 , n39029 , n39107 );
or ( n39109 , n39028 , n39108 );
and ( n39110 , n39026 , n39109 );
and ( n39111 , n39025 , n39110 );
or ( n39112 , n39024 , n39111 );
and ( n39113 , n38377 , n39112 );
and ( n39114 , n38375 , n39113 );
or ( n39115 , n38374 , n39114 );
and ( n39116 , n38372 , n39115 );
or ( n39117 , n38371 , n39116 );
and ( n39118 , n38369 , n39117 );
and ( n39119 , n38367 , n39118 );
or ( n39120 , n38366 , n39119 );
and ( n39121 , n37750 , n39120 );
or ( n39122 , n37749 , n39121 );
and ( n39123 , n37482 , n39122 );
and ( n39124 , n37480 , n39123 );
or ( n39125 , n37479 , n39124 );
and ( n39126 , n37477 , n39125 );
or ( n39127 , n37476 , n39126 );
and ( n39128 , n37168 , n39127 );
and ( n39129 , n37166 , n39128 );
and ( n39130 , n37165 , n39129 );
or ( n39131 , n37164 , n39130 );
and ( n39132 , n36618 , n39131 );
and ( n39133 , n36616 , n39132 );
or ( n39134 , n36615 , n39133 );
and ( n39135 , n36182 , n39134 );
and ( n39136 , n36181 , n39135 );
and ( n39137 , n36180 , n39136 );
and ( n39138 , n36178 , n39137 );
or ( n39139 , n36177 , n39138 );
and ( n39140 , n35705 , n39139 );
and ( n39141 , n35704 , n39140 );
or ( n39142 , n35703 , n39141 );
and ( n39143 , n35701 , n39142 );
and ( n39144 , n35700 , n39143 );
or ( n39145 , n35699 , n39144 );
and ( n39146 , n35697 , n39145 );
and ( n39147 , n35695 , n39146 );
and ( n39148 , n35693 , n39147 );
or ( n39149 , n35692 , n39148 );
and ( n39150 , n33671 , n39149 );
and ( n39151 , n33670 , n39150 );
and ( n39152 , n33668 , n39151 );
or ( n39153 , n33667 , n39152 );
and ( n39154 , n33665 , n39153 );
or ( n39155 , n33664 , n39154 );
and ( n39156 , n33662 , n39155 );
or ( n39157 , n33661 , n39156 );
and ( n39158 , n32471 , n39157 );
or ( n39159 , n32470 , n39158 );
and ( n39160 , n32118 , n39159 );
or ( n39161 , n32117 , n39160 );
and ( n39162 , n31831 , n39161 );
or ( n39163 , n31830 , n39162 );
and ( n39164 , n31826 , n39163 );
or ( n39165 , n31825 , n39164 );
and ( n39166 , n31823 , n39165 );
or ( n39167 , n31822 , n39166 );
and ( n39168 , n31421 , n39167 );
and ( n39169 , n31420 , n39168 );
or ( n39170 , n31419 , n39169 );
and ( n39171 , n31221 , n39170 );
and ( n39172 , n31219 , n39171 );
or ( n39173 , n31218 , n39172 );
and ( n39174 , n30936 , n39173 );
and ( n39175 , n30935 , n39174 );
or ( n39176 , n30934 , n39175 );
and ( n39177 , n30761 , n39176 );
or ( n39178 , n30760 , n39177 );
and ( n39179 , n30758 , n39178 );
and ( n39180 , n30757 , n39179 );
xor ( n39181 , n30756 , n39180 );
buf ( n39182 , n39181 );
buf ( n39183 , n39182 );
buf ( n39184 , n39183 );
buf ( n39185 , n1154 );
buf ( n39186 , n39185 );
buf ( n39187 , n1155 );
buf ( n39188 , n39187 );
xor ( n39189 , n39186 , n39188 );
buf ( n39190 , n1156 );
buf ( n39191 , n39190 );
xor ( n39192 , n39188 , n39191 );
not ( n39193 , n39192 );
and ( n39194 , n39189 , n39193 );
and ( n39195 , n39184 , n39194 );
not ( n39196 , n39195 );
and ( n39197 , n39188 , n39191 );
not ( n39198 , n39197 );
and ( n39199 , n39186 , n39198 );
xnor ( n39200 , n39196 , n39199 );
buf ( n39201 , n39200 );
not ( n39202 , n39199 );
and ( n39203 , n39201 , n39202 );
and ( n39204 , n39184 , n39186 );
and ( n39205 , n39202 , n39204 );
and ( n39206 , n39201 , n39204 );
or ( n39207 , n39203 , n39205 , n39206 );
buf ( n39208 , n39207 );
buf ( n39209 , n1157 );
buf ( n39210 , n39209 );
buf ( n39211 , n1158 );
buf ( n39212 , n39211 );
and ( n39213 , n39210 , n39212 );
not ( n39214 , n39213 );
and ( n39215 , n39191 , n39214 );
not ( n39216 , n39215 );
xor ( n39217 , n30757 , n39179 );
buf ( n39218 , n39217 );
buf ( n39219 , n39218 );
buf ( n39220 , n39219 );
and ( n39221 , n39220 , n39194 );
and ( n39222 , n39184 , n39192 );
nor ( n39223 , n39221 , n39222 );
xnor ( n39224 , n39223 , n39199 );
and ( n39225 , n39216 , n39224 );
xor ( n39226 , n30758 , n39178 );
buf ( n39227 , n39226 );
buf ( n39228 , n39227 );
buf ( n39229 , n39228 );
and ( n39230 , n39229 , n39186 );
and ( n39231 , n39224 , n39230 );
and ( n39232 , n39216 , n39230 );
or ( n39233 , n39225 , n39231 , n39232 );
not ( n39234 , n39200 );
and ( n39235 , n39233 , n39234 );
and ( n39236 , n39220 , n39186 );
and ( n39237 , n39234 , n39236 );
and ( n39238 , n39233 , n39236 );
or ( n39239 , n39235 , n39237 , n39238 );
buf ( n39240 , n39239 );
xor ( n39241 , n39201 , n39202 );
xor ( n39242 , n39241 , n39204 );
and ( n39243 , n39239 , n39242 );
buf ( n39244 , n39242 );
or ( n39245 , n39240 , n39243 , n39244 );
and ( n39246 , n39207 , n39245 );
buf ( n39247 , n39245 );
or ( n39248 , n39208 , n39246 , n39247 );
buf ( n39249 , n39248 );
not ( n39250 , n39207 );
xor ( n39251 , n39250 , n39245 );
xor ( n39252 , n39233 , n39234 );
xor ( n39253 , n39252 , n39236 );
buf ( n39254 , n39253 );
xor ( n39255 , n39191 , n39210 );
xor ( n39256 , n39210 , n39212 );
not ( n39257 , n39256 );
and ( n39258 , n39255 , n39257 );
and ( n39259 , n39184 , n39258 );
not ( n39260 , n39259 );
xnor ( n39261 , n39260 , n39215 );
not ( n39262 , n39261 );
and ( n39263 , n39229 , n39194 );
and ( n39264 , n39220 , n39192 );
nor ( n39265 , n39263 , n39264 );
xnor ( n39266 , n39265 , n39199 );
and ( n39267 , n39262 , n39266 );
xor ( n39268 , n30761 , n39176 );
buf ( n39269 , n39268 );
buf ( n39270 , n39269 );
buf ( n39271 , n39270 );
and ( n39272 , n39271 , n39186 );
and ( n39273 , n39266 , n39272 );
and ( n39274 , n39262 , n39272 );
or ( n39275 , n39267 , n39273 , n39274 );
buf ( n39276 , n39261 );
and ( n39277 , n39275 , n39276 );
xor ( n39278 , n39216 , n39224 );
xor ( n39279 , n39278 , n39230 );
and ( n39280 , n39276 , n39279 );
and ( n39281 , n39275 , n39279 );
or ( n39282 , n39277 , n39280 , n39281 );
and ( n39283 , n39253 , n39282 );
buf ( n39284 , n39282 );
or ( n39285 , n39254 , n39283 , n39284 );
not ( n39286 , n39239 );
xor ( n39287 , n39286 , n39242 );
and ( n39288 , n39285 , n39287 );
not ( n39289 , n39253 );
xor ( n39290 , n39289 , n39282 );
xor ( n39291 , n39275 , n39276 );
xor ( n39292 , n39291 , n39279 );
buf ( n39293 , n39292 );
buf ( n39294 , n1159 );
buf ( n39295 , n39294 );
buf ( n39296 , n1160 );
buf ( n39297 , n39296 );
and ( n39298 , n39295 , n39297 );
not ( n39299 , n39298 );
and ( n39300 , n39212 , n39299 );
not ( n39301 , n39300 );
and ( n39302 , n39220 , n39258 );
and ( n39303 , n39184 , n39256 );
nor ( n39304 , n39302 , n39303 );
xnor ( n39305 , n39304 , n39215 );
and ( n39306 , n39301 , n39305 );
xor ( n39307 , n30935 , n39174 );
buf ( n39308 , n39307 );
buf ( n39309 , n39308 );
buf ( n39310 , n39309 );
and ( n39311 , n39310 , n39186 );
and ( n39312 , n39305 , n39311 );
and ( n39313 , n39301 , n39311 );
or ( n39314 , n39306 , n39312 , n39313 );
and ( n39315 , n39229 , n39258 );
and ( n39316 , n39220 , n39256 );
nor ( n39317 , n39315 , n39316 );
xnor ( n39318 , n39317 , n39215 );
and ( n39319 , n39310 , n39194 );
and ( n39320 , n39271 , n39192 );
nor ( n39321 , n39319 , n39320 );
xnor ( n39322 , n39321 , n39199 );
and ( n39323 , n39318 , n39322 );
xor ( n39324 , n30936 , n39173 );
buf ( n39325 , n39324 );
buf ( n39326 , n39325 );
buf ( n39327 , n39326 );
and ( n39328 , n39327 , n39186 );
and ( n39329 , n39322 , n39328 );
and ( n39330 , n39318 , n39328 );
or ( n39331 , n39323 , n39329 , n39330 );
xor ( n39332 , n39212 , n39295 );
xor ( n39333 , n39295 , n39297 );
not ( n39334 , n39333 );
and ( n39335 , n39332 , n39334 );
and ( n39336 , n39184 , n39335 );
not ( n39337 , n39336 );
xnor ( n39338 , n39337 , n39300 );
buf ( n39339 , n39338 );
and ( n39340 , n39331 , n39339 );
and ( n39341 , n39271 , n39194 );
and ( n39342 , n39229 , n39192 );
nor ( n39343 , n39341 , n39342 );
xnor ( n39344 , n39343 , n39199 );
and ( n39345 , n39339 , n39344 );
and ( n39346 , n39331 , n39344 );
or ( n39347 , n39340 , n39345 , n39346 );
and ( n39348 , n39314 , n39347 );
xor ( n39349 , n39262 , n39266 );
xor ( n39350 , n39349 , n39272 );
and ( n39351 , n39347 , n39350 );
and ( n39352 , n39314 , n39350 );
or ( n39353 , n39348 , n39351 , n39352 );
and ( n39354 , n39292 , n39353 );
buf ( n39355 , n39353 );
or ( n39356 , n39293 , n39354 , n39355 );
and ( n39357 , n39290 , n39356 );
xor ( n39358 , n39314 , n39347 );
xor ( n39359 , n39358 , n39350 );
buf ( n39360 , n39359 );
buf ( n39361 , n1161 );
buf ( n39362 , n39361 );
buf ( n39363 , n1162 );
buf ( n39364 , n39363 );
and ( n39365 , n39362 , n39364 );
not ( n39366 , n39365 );
and ( n39367 , n39297 , n39366 );
not ( n39368 , n39367 );
and ( n39369 , n39220 , n39335 );
and ( n39370 , n39184 , n39333 );
nor ( n39371 , n39369 , n39370 );
xnor ( n39372 , n39371 , n39300 );
and ( n39373 , n39368 , n39372 );
and ( n39374 , n39327 , n39194 );
and ( n39375 , n39310 , n39192 );
nor ( n39376 , n39374 , n39375 );
xnor ( n39377 , n39376 , n39199 );
and ( n39378 , n39372 , n39377 );
and ( n39379 , n39368 , n39377 );
or ( n39380 , n39373 , n39378 , n39379 );
xor ( n39381 , n39297 , n39362 );
xor ( n39382 , n39362 , n39364 );
not ( n39383 , n39382 );
and ( n39384 , n39381 , n39383 );
and ( n39385 , n39184 , n39384 );
not ( n39386 , n39385 );
xnor ( n39387 , n39386 , n39367 );
buf ( n39388 , n39387 );
and ( n39389 , n39271 , n39258 );
and ( n39390 , n39229 , n39256 );
nor ( n39391 , n39389 , n39390 );
xnor ( n39392 , n39391 , n39215 );
and ( n39393 , n39388 , n39392 );
xor ( n39394 , n31219 , n39171 );
buf ( n39395 , n39394 );
buf ( n39396 , n39395 );
buf ( n39397 , n39396 );
and ( n39398 , n39397 , n39186 );
and ( n39399 , n39392 , n39398 );
and ( n39400 , n39388 , n39398 );
or ( n39401 , n39393 , n39399 , n39400 );
and ( n39402 , n39380 , n39401 );
not ( n39403 , n39338 );
and ( n39404 , n39401 , n39403 );
and ( n39405 , n39380 , n39403 );
or ( n39406 , n39402 , n39404 , n39405 );
xor ( n39407 , n39301 , n39305 );
xor ( n39408 , n39407 , n39311 );
and ( n39409 , n39406 , n39408 );
xor ( n39410 , n39331 , n39339 );
xor ( n39411 , n39410 , n39344 );
and ( n39412 , n39408 , n39411 );
and ( n39413 , n39406 , n39411 );
or ( n39414 , n39409 , n39412 , n39413 );
and ( n39415 , n39359 , n39414 );
buf ( n39416 , n39414 );
or ( n39417 , n39360 , n39415 , n39416 );
not ( n39418 , n39292 );
xor ( n39419 , n39418 , n39353 );
and ( n39420 , n39417 , n39419 );
and ( n39421 , n39229 , n39335 );
and ( n39422 , n39220 , n39333 );
nor ( n39423 , n39421 , n39422 );
xnor ( n39424 , n39423 , n39300 );
and ( n39425 , n39397 , n39194 );
and ( n39426 , n39327 , n39192 );
nor ( n39427 , n39425 , n39426 );
xnor ( n39428 , n39427 , n39199 );
and ( n39429 , n39424 , n39428 );
xor ( n39430 , n31221 , n39170 );
buf ( n39431 , n39430 );
buf ( n39432 , n39431 );
buf ( n39433 , n39432 );
and ( n39434 , n39433 , n39186 );
and ( n39435 , n39428 , n39434 );
and ( n39436 , n39424 , n39434 );
or ( n39437 , n39429 , n39435 , n39436 );
xor ( n39438 , n39368 , n39372 );
xor ( n39439 , n39438 , n39377 );
and ( n39440 , n39437 , n39439 );
xor ( n39441 , n39388 , n39392 );
xor ( n39442 , n39441 , n39398 );
and ( n39443 , n39439 , n39442 );
and ( n39444 , n39437 , n39442 );
or ( n39445 , n39440 , n39443 , n39444 );
xor ( n39446 , n39318 , n39322 );
xor ( n39447 , n39446 , n39328 );
and ( n39448 , n39445 , n39447 );
xor ( n39449 , n39380 , n39401 );
xor ( n39450 , n39449 , n39403 );
and ( n39451 , n39447 , n39450 );
and ( n39452 , n39445 , n39450 );
or ( n39453 , n39448 , n39451 , n39452 );
buf ( n39454 , n39453 );
xor ( n39455 , n39406 , n39408 );
xor ( n39456 , n39455 , n39411 );
and ( n39457 , n39453 , n39456 );
buf ( n39458 , n39456 );
or ( n39459 , n39454 , n39457 , n39458 );
not ( n39460 , n39359 );
xor ( n39461 , n39460 , n39414 );
and ( n39462 , n39459 , n39461 );
xor ( n39463 , n39445 , n39447 );
xor ( n39464 , n39463 , n39450 );
buf ( n39465 , n39464 );
and ( n39466 , n39271 , n39335 );
and ( n39467 , n39229 , n39333 );
nor ( n39468 , n39466 , n39467 );
xnor ( n39469 , n39468 , n39300 );
and ( n39470 , n39327 , n39258 );
and ( n39471 , n39310 , n39256 );
nor ( n39472 , n39470 , n39471 );
xnor ( n39473 , n39472 , n39215 );
and ( n39474 , n39469 , n39473 );
and ( n39475 , n39433 , n39194 );
and ( n39476 , n39397 , n39192 );
nor ( n39477 , n39475 , n39476 );
xnor ( n39478 , n39477 , n39199 );
and ( n39479 , n39473 , n39478 );
and ( n39480 , n39469 , n39478 );
or ( n39481 , n39474 , n39479 , n39480 );
not ( n39482 , n39387 );
and ( n39483 , n39481 , n39482 );
and ( n39484 , n39310 , n39258 );
and ( n39485 , n39271 , n39256 );
nor ( n39486 , n39484 , n39485 );
xnor ( n39487 , n39486 , n39215 );
and ( n39488 , n39482 , n39487 );
and ( n39489 , n39481 , n39487 );
or ( n39490 , n39483 , n39488 , n39489 );
buf ( n39491 , n1163 );
buf ( n39492 , n39491 );
buf ( n39493 , n1164 );
buf ( n39494 , n39493 );
and ( n39495 , n39492 , n39494 );
not ( n39496 , n39495 );
and ( n39497 , n39364 , n39496 );
not ( n39498 , n39497 );
and ( n39499 , n39220 , n39384 );
and ( n39500 , n39184 , n39382 );
nor ( n39501 , n39499 , n39500 );
xnor ( n39502 , n39501 , n39367 );
and ( n39503 , n39498 , n39502 );
xor ( n39504 , n31420 , n39168 );
buf ( n39505 , n39504 );
buf ( n39506 , n39505 );
buf ( n39507 , n39506 );
and ( n39508 , n39507 , n39186 );
and ( n39509 , n39502 , n39508 );
and ( n39510 , n39498 , n39508 );
or ( n39511 , n39503 , n39509 , n39510 );
and ( n39512 , n39229 , n39384 );
and ( n39513 , n39220 , n39382 );
nor ( n39514 , n39512 , n39513 );
xnor ( n39515 , n39514 , n39367 );
and ( n39516 , n39397 , n39258 );
and ( n39517 , n39327 , n39256 );
nor ( n39518 , n39516 , n39517 );
xnor ( n39519 , n39518 , n39215 );
and ( n39520 , n39515 , n39519 );
xor ( n39521 , n31421 , n39167 );
buf ( n39522 , n39521 );
buf ( n39523 , n39522 );
buf ( n39524 , n39523 );
and ( n39525 , n39524 , n39186 );
and ( n39526 , n39519 , n39525 );
and ( n39527 , n39515 , n39525 );
or ( n39528 , n39520 , n39526 , n39527 );
xor ( n39529 , n39364 , n39492 );
xor ( n39530 , n39492 , n39494 );
not ( n39531 , n39530 );
and ( n39532 , n39529 , n39531 );
and ( n39533 , n39184 , n39532 );
not ( n39534 , n39533 );
xnor ( n39535 , n39534 , n39497 );
buf ( n39536 , n39535 );
and ( n39537 , n39528 , n39536 );
xor ( n39538 , n39498 , n39502 );
xor ( n39539 , n39538 , n39508 );
and ( n39540 , n39536 , n39539 );
and ( n39541 , n39528 , n39539 );
or ( n39542 , n39537 , n39540 , n39541 );
and ( n39543 , n39511 , n39542 );
xor ( n39544 , n39424 , n39428 );
xor ( n39545 , n39544 , n39434 );
and ( n39546 , n39542 , n39545 );
and ( n39547 , n39511 , n39545 );
or ( n39548 , n39543 , n39546 , n39547 );
and ( n39549 , n39490 , n39548 );
xor ( n39550 , n39437 , n39439 );
xor ( n39551 , n39550 , n39442 );
and ( n39552 , n39548 , n39551 );
and ( n39553 , n39490 , n39551 );
or ( n39554 , n39549 , n39552 , n39553 );
and ( n39555 , n39464 , n39554 );
buf ( n39556 , n39554 );
or ( n39557 , n39465 , n39555 , n39556 );
not ( n39558 , n39453 );
xor ( n39559 , n39558 , n39456 );
and ( n39560 , n39557 , n39559 );
not ( n39561 , n39535 );
and ( n39562 , n39310 , n39335 );
and ( n39563 , n39271 , n39333 );
nor ( n39564 , n39562 , n39563 );
xnor ( n39565 , n39564 , n39300 );
and ( n39566 , n39561 , n39565 );
and ( n39567 , n39507 , n39194 );
and ( n39568 , n39433 , n39192 );
nor ( n39569 , n39567 , n39568 );
xnor ( n39570 , n39569 , n39199 );
and ( n39571 , n39565 , n39570 );
and ( n39572 , n39561 , n39570 );
or ( n39573 , n39566 , n39571 , n39572 );
xor ( n39574 , n39469 , n39473 );
xor ( n39575 , n39574 , n39478 );
and ( n39576 , n39573 , n39575 );
xor ( n39577 , n39528 , n39536 );
xor ( n39578 , n39577 , n39539 );
and ( n39579 , n39575 , n39578 );
and ( n39580 , n39573 , n39578 );
or ( n39581 , n39576 , n39579 , n39580 );
xor ( n39582 , n39481 , n39482 );
xor ( n39583 , n39582 , n39487 );
and ( n39584 , n39581 , n39583 );
xor ( n39585 , n39511 , n39542 );
xor ( n39586 , n39585 , n39545 );
and ( n39587 , n39583 , n39586 );
and ( n39588 , n39581 , n39586 );
or ( n39589 , n39584 , n39587 , n39588 );
buf ( n39590 , n39589 );
xor ( n39591 , n39490 , n39548 );
xor ( n39592 , n39591 , n39551 );
and ( n39593 , n39589 , n39592 );
buf ( n39594 , n39592 );
or ( n39595 , n39590 , n39593 , n39594 );
not ( n39596 , n39464 );
xor ( n39597 , n39596 , n39554 );
and ( n39598 , n39595 , n39597 );
xor ( n39599 , n39581 , n39583 );
xor ( n39600 , n39599 , n39586 );
buf ( n39601 , n39600 );
buf ( n39602 , n1165 );
buf ( n39603 , n39602 );
buf ( n39604 , n1166 );
buf ( n39605 , n39604 );
and ( n39606 , n39603 , n39605 );
not ( n39607 , n39606 );
and ( n39608 , n39494 , n39607 );
not ( n39609 , n39608 );
and ( n39610 , n39524 , n39194 );
and ( n39611 , n39507 , n39192 );
nor ( n39612 , n39610 , n39611 );
xnor ( n39613 , n39612 , n39199 );
and ( n39614 , n39609 , n39613 );
xor ( n39615 , n31823 , n39165 );
buf ( n39616 , n39615 );
buf ( n39617 , n39616 );
buf ( n39618 , n39617 );
and ( n39619 , n39618 , n39186 );
and ( n39620 , n39613 , n39619 );
and ( n39621 , n39609 , n39619 );
or ( n39622 , n39614 , n39620 , n39621 );
and ( n39623 , n39220 , n39532 );
and ( n39624 , n39184 , n39530 );
nor ( n39625 , n39623 , n39624 );
xnor ( n39626 , n39625 , n39497 );
and ( n39627 , n39327 , n39335 );
and ( n39628 , n39310 , n39333 );
nor ( n39629 , n39627 , n39628 );
xnor ( n39630 , n39629 , n39300 );
and ( n39631 , n39626 , n39630 );
and ( n39632 , n39433 , n39258 );
and ( n39633 , n39397 , n39256 );
nor ( n39634 , n39632 , n39633 );
xnor ( n39635 , n39634 , n39215 );
and ( n39636 , n39630 , n39635 );
and ( n39637 , n39626 , n39635 );
or ( n39638 , n39631 , n39636 , n39637 );
and ( n39639 , n39622 , n39638 );
xor ( n39640 , n39561 , n39565 );
xor ( n39641 , n39640 , n39570 );
and ( n39642 , n39638 , n39641 );
and ( n39643 , n39622 , n39641 );
or ( n39644 , n39639 , n39642 , n39643 );
and ( n39645 , n39229 , n39532 );
and ( n39646 , n39220 , n39530 );
nor ( n39647 , n39645 , n39646 );
xnor ( n39648 , n39647 , n39497 );
and ( n39649 , n39618 , n39194 );
and ( n39650 , n39524 , n39192 );
nor ( n39651 , n39649 , n39650 );
xnor ( n39652 , n39651 , n39199 );
and ( n39653 , n39648 , n39652 );
xor ( n39654 , n31826 , n39163 );
buf ( n39655 , n39654 );
buf ( n39656 , n39655 );
buf ( n39657 , n39656 );
and ( n39658 , n39657 , n39186 );
and ( n39659 , n39652 , n39658 );
and ( n39660 , n39648 , n39658 );
or ( n39661 , n39653 , n39659 , n39660 );
xor ( n39662 , n39494 , n39603 );
xor ( n39663 , n39603 , n39605 );
not ( n39664 , n39663 );
and ( n39665 , n39662 , n39664 );
and ( n39666 , n39184 , n39665 );
not ( n39667 , n39666 );
xnor ( n39668 , n39667 , n39608 );
buf ( n39669 , n39668 );
and ( n39670 , n39661 , n39669 );
and ( n39671 , n39271 , n39384 );
and ( n39672 , n39229 , n39382 );
nor ( n39673 , n39671 , n39672 );
xnor ( n39674 , n39673 , n39367 );
and ( n39675 , n39669 , n39674 );
and ( n39676 , n39661 , n39674 );
or ( n39677 , n39670 , n39675 , n39676 );
and ( n39678 , n39310 , n39384 );
and ( n39679 , n39271 , n39382 );
nor ( n39680 , n39678 , n39679 );
xnor ( n39681 , n39680 , n39367 );
and ( n39682 , n39397 , n39335 );
and ( n39683 , n39327 , n39333 );
nor ( n39684 , n39682 , n39683 );
xnor ( n39685 , n39684 , n39300 );
and ( n39686 , n39681 , n39685 );
and ( n39687 , n39507 , n39258 );
and ( n39688 , n39433 , n39256 );
nor ( n39689 , n39687 , n39688 );
xnor ( n39690 , n39689 , n39215 );
and ( n39691 , n39685 , n39690 );
and ( n39692 , n39681 , n39690 );
or ( n39693 , n39686 , n39691 , n39692 );
xor ( n39694 , n39609 , n39613 );
xor ( n39695 , n39694 , n39619 );
and ( n39696 , n39693 , n39695 );
xor ( n39697 , n39626 , n39630 );
xor ( n39698 , n39697 , n39635 );
and ( n39699 , n39695 , n39698 );
and ( n39700 , n39693 , n39698 );
or ( n39701 , n39696 , n39699 , n39700 );
and ( n39702 , n39677 , n39701 );
xor ( n39703 , n39515 , n39519 );
xor ( n39704 , n39703 , n39525 );
and ( n39705 , n39701 , n39704 );
and ( n39706 , n39677 , n39704 );
or ( n39707 , n39702 , n39705 , n39706 );
and ( n39708 , n39644 , n39707 );
xor ( n39709 , n39573 , n39575 );
xor ( n39710 , n39709 , n39578 );
and ( n39711 , n39707 , n39710 );
and ( n39712 , n39644 , n39710 );
or ( n39713 , n39708 , n39711 , n39712 );
and ( n39714 , n39600 , n39713 );
buf ( n39715 , n39713 );
or ( n39716 , n39601 , n39714 , n39715 );
not ( n39717 , n39589 );
xor ( n39718 , n39717 , n39592 );
and ( n39719 , n39716 , n39718 );
xor ( n39720 , n39644 , n39707 );
xor ( n39721 , n39720 , n39710 );
buf ( n39722 , n39721 );
buf ( n39723 , n1167 );
buf ( n39724 , n39723 );
buf ( n39725 , n1168 );
buf ( n39726 , n39725 );
and ( n39727 , n39724 , n39726 );
not ( n39728 , n39727 );
and ( n39729 , n39605 , n39728 );
not ( n39730 , n39729 );
and ( n39731 , n39524 , n39258 );
and ( n39732 , n39507 , n39256 );
nor ( n39733 , n39731 , n39732 );
xnor ( n39734 , n39733 , n39215 );
and ( n39735 , n39730 , n39734 );
xor ( n39736 , n31831 , n39161 );
buf ( n39737 , n39736 );
buf ( n39738 , n39737 );
buf ( n39739 , n39738 );
and ( n39740 , n39739 , n39186 );
and ( n39741 , n39734 , n39740 );
and ( n39742 , n39730 , n39740 );
or ( n39743 , n39735 , n39741 , n39742 );
and ( n39744 , n39220 , n39665 );
and ( n39745 , n39184 , n39663 );
nor ( n39746 , n39744 , n39745 );
xnor ( n39747 , n39746 , n39608 );
and ( n39748 , n39327 , n39384 );
and ( n39749 , n39310 , n39382 );
nor ( n39750 , n39748 , n39749 );
xnor ( n39751 , n39750 , n39367 );
and ( n39752 , n39747 , n39751 );
and ( n39753 , n39657 , n39194 );
and ( n39754 , n39618 , n39192 );
nor ( n39755 , n39753 , n39754 );
xnor ( n39756 , n39755 , n39199 );
and ( n39757 , n39751 , n39756 );
and ( n39758 , n39747 , n39756 );
or ( n39759 , n39752 , n39757 , n39758 );
and ( n39760 , n39743 , n39759 );
not ( n39761 , n39668 );
and ( n39762 , n39759 , n39761 );
and ( n39763 , n39743 , n39761 );
or ( n39764 , n39760 , n39762 , n39763 );
xor ( n39765 , n39661 , n39669 );
xor ( n39766 , n39765 , n39674 );
and ( n39767 , n39764 , n39766 );
xor ( n39768 , n39693 , n39695 );
xor ( n39769 , n39768 , n39698 );
and ( n39770 , n39766 , n39769 );
and ( n39771 , n39764 , n39769 );
or ( n39772 , n39767 , n39770 , n39771 );
xor ( n39773 , n39622 , n39638 );
xor ( n39774 , n39773 , n39641 );
and ( n39775 , n39772 , n39774 );
xor ( n39776 , n39677 , n39701 );
xor ( n39777 , n39776 , n39704 );
and ( n39778 , n39774 , n39777 );
and ( n39779 , n39772 , n39777 );
or ( n39780 , n39775 , n39778 , n39779 );
and ( n39781 , n39721 , n39780 );
buf ( n39782 , n39780 );
or ( n39783 , n39722 , n39781 , n39782 );
not ( n39784 , n39600 );
xor ( n39785 , n39784 , n39713 );
and ( n39786 , n39783 , n39785 );
not ( n39787 , n39721 );
xor ( n39788 , n39787 , n39780 );
xor ( n39789 , n39772 , n39774 );
xor ( n39790 , n39789 , n39777 );
buf ( n39791 , n39790 );
xor ( n39792 , n39605 , n39724 );
xor ( n39793 , n39724 , n39726 );
not ( n39794 , n39793 );
and ( n39795 , n39792 , n39794 );
and ( n39796 , n39184 , n39795 );
not ( n39797 , n39796 );
xnor ( n39798 , n39797 , n39729 );
buf ( n39799 , n39798 );
and ( n39800 , n39271 , n39532 );
and ( n39801 , n39229 , n39530 );
nor ( n39802 , n39800 , n39801 );
xnor ( n39803 , n39802 , n39497 );
and ( n39804 , n39799 , n39803 );
and ( n39805 , n39433 , n39335 );
and ( n39806 , n39397 , n39333 );
nor ( n39807 , n39805 , n39806 );
xnor ( n39808 , n39807 , n39300 );
and ( n39809 , n39803 , n39808 );
and ( n39810 , n39799 , n39808 );
or ( n39811 , n39804 , n39809 , n39810 );
xor ( n39812 , n39648 , n39652 );
xor ( n39813 , n39812 , n39658 );
and ( n39814 , n39811 , n39813 );
xor ( n39815 , n39681 , n39685 );
xor ( n39816 , n39815 , n39690 );
and ( n39817 , n39813 , n39816 );
and ( n39818 , n39811 , n39816 );
or ( n39819 , n39814 , n39817 , n39818 );
and ( n39820 , n39229 , n39665 );
and ( n39821 , n39220 , n39663 );
nor ( n39822 , n39820 , n39821 );
xnor ( n39823 , n39822 , n39608 );
and ( n39824 , n39397 , n39384 );
and ( n39825 , n39327 , n39382 );
nor ( n39826 , n39824 , n39825 );
xnor ( n39827 , n39826 , n39367 );
and ( n39828 , n39823 , n39827 );
and ( n39829 , n39507 , n39335 );
and ( n39830 , n39433 , n39333 );
nor ( n39831 , n39829 , n39830 );
xnor ( n39832 , n39831 , n39300 );
and ( n39833 , n39827 , n39832 );
and ( n39834 , n39823 , n39832 );
or ( n39835 , n39828 , n39833 , n39834 );
and ( n39836 , n39618 , n39258 );
and ( n39837 , n39524 , n39256 );
nor ( n39838 , n39836 , n39837 );
xnor ( n39839 , n39838 , n39215 );
and ( n39840 , n39739 , n39194 );
and ( n39841 , n39657 , n39192 );
nor ( n39842 , n39840 , n39841 );
xnor ( n39843 , n39842 , n39199 );
and ( n39844 , n39839 , n39843 );
xor ( n39845 , n32118 , n39159 );
buf ( n39846 , n39845 );
buf ( n39847 , n39846 );
buf ( n39848 , n39847 );
and ( n39849 , n39848 , n39186 );
and ( n39850 , n39843 , n39849 );
and ( n39851 , n39839 , n39849 );
or ( n39852 , n39844 , n39850 , n39851 );
and ( n39853 , n39835 , n39852 );
xor ( n39854 , n39730 , n39734 );
xor ( n39855 , n39854 , n39740 );
and ( n39856 , n39852 , n39855 );
and ( n39857 , n39835 , n39855 );
or ( n39858 , n39853 , n39856 , n39857 );
buf ( n39859 , n1169 );
buf ( n39860 , n39859 );
buf ( n39861 , n1170 );
buf ( n39862 , n39861 );
and ( n39863 , n39860 , n39862 );
not ( n39864 , n39863 );
and ( n39865 , n39726 , n39864 );
not ( n39866 , n39865 );
and ( n39867 , n39848 , n39194 );
and ( n39868 , n39739 , n39192 );
nor ( n39869 , n39867 , n39868 );
xnor ( n39870 , n39869 , n39199 );
and ( n39871 , n39866 , n39870 );
xor ( n39872 , n32471 , n39157 );
buf ( n39873 , n39872 );
buf ( n39874 , n39873 );
buf ( n39875 , n39874 );
and ( n39876 , n39875 , n39186 );
and ( n39877 , n39870 , n39876 );
and ( n39878 , n39866 , n39876 );
or ( n39879 , n39871 , n39877 , n39878 );
not ( n39880 , n39798 );
and ( n39881 , n39879 , n39880 );
and ( n39882 , n39310 , n39532 );
and ( n39883 , n39271 , n39530 );
nor ( n39884 , n39882 , n39883 );
xnor ( n39885 , n39884 , n39497 );
and ( n39886 , n39880 , n39885 );
and ( n39887 , n39879 , n39885 );
or ( n39888 , n39881 , n39886 , n39887 );
xor ( n39889 , n39747 , n39751 );
xor ( n39890 , n39889 , n39756 );
and ( n39891 , n39888 , n39890 );
xor ( n39892 , n39799 , n39803 );
xor ( n39893 , n39892 , n39808 );
and ( n39894 , n39890 , n39893 );
and ( n39895 , n39888 , n39893 );
or ( n39896 , n39891 , n39894 , n39895 );
and ( n39897 , n39858 , n39896 );
xor ( n39898 , n39743 , n39759 );
xor ( n39899 , n39898 , n39761 );
and ( n39900 , n39896 , n39899 );
and ( n39901 , n39858 , n39899 );
or ( n39902 , n39897 , n39900 , n39901 );
and ( n39903 , n39819 , n39902 );
xor ( n39904 , n39764 , n39766 );
xor ( n39905 , n39904 , n39769 );
and ( n39906 , n39902 , n39905 );
and ( n39907 , n39819 , n39905 );
or ( n39908 , n39903 , n39906 , n39907 );
and ( n39909 , n39790 , n39908 );
buf ( n39910 , n39908 );
or ( n39911 , n39791 , n39909 , n39910 );
and ( n39912 , n39788 , n39911 );
xor ( n39913 , n39819 , n39902 );
xor ( n39914 , n39913 , n39905 );
buf ( n39915 , n39914 );
and ( n39916 , n39327 , n39532 );
and ( n39917 , n39310 , n39530 );
nor ( n39918 , n39916 , n39917 );
xnor ( n39919 , n39918 , n39497 );
and ( n39920 , n39524 , n39335 );
and ( n39921 , n39507 , n39333 );
nor ( n39922 , n39920 , n39921 );
xnor ( n39923 , n39922 , n39300 );
and ( n39924 , n39919 , n39923 );
and ( n39925 , n39657 , n39258 );
and ( n39926 , n39618 , n39256 );
nor ( n39927 , n39925 , n39926 );
xnor ( n39928 , n39927 , n39215 );
and ( n39929 , n39923 , n39928 );
and ( n39930 , n39919 , n39928 );
or ( n39931 , n39924 , n39929 , n39930 );
xor ( n39932 , n33662 , n39155 );
buf ( n39933 , n39932 );
buf ( n39934 , n39933 );
buf ( n39935 , n39934 );
and ( n39936 , n39935 , n39186 );
buf ( n39937 , n39936 );
and ( n39938 , n39220 , n39795 );
and ( n39939 , n39184 , n39793 );
nor ( n39940 , n39938 , n39939 );
xnor ( n39941 , n39940 , n39729 );
and ( n39942 , n39937 , n39941 );
and ( n39943 , n39433 , n39384 );
and ( n39944 , n39397 , n39382 );
nor ( n39945 , n39943 , n39944 );
xnor ( n39946 , n39945 , n39367 );
and ( n39947 , n39941 , n39946 );
and ( n39948 , n39937 , n39946 );
or ( n39949 , n39942 , n39947 , n39948 );
and ( n39950 , n39931 , n39949 );
xor ( n39951 , n39839 , n39843 );
xor ( n39952 , n39951 , n39849 );
and ( n39953 , n39949 , n39952 );
and ( n39954 , n39931 , n39952 );
or ( n39955 , n39950 , n39953 , n39954 );
xor ( n39956 , n39835 , n39852 );
xor ( n39957 , n39956 , n39855 );
and ( n39958 , n39955 , n39957 );
xor ( n39959 , n39888 , n39890 );
xor ( n39960 , n39959 , n39893 );
and ( n39961 , n39957 , n39960 );
and ( n39962 , n39955 , n39960 );
or ( n39963 , n39958 , n39961 , n39962 );
xor ( n39964 , n39811 , n39813 );
xor ( n39965 , n39964 , n39816 );
and ( n39966 , n39963 , n39965 );
xor ( n39967 , n39858 , n39896 );
xor ( n39968 , n39967 , n39899 );
and ( n39969 , n39965 , n39968 );
and ( n39970 , n39963 , n39968 );
or ( n39971 , n39966 , n39969 , n39970 );
and ( n39972 , n39914 , n39971 );
buf ( n39973 , n39971 );
or ( n39974 , n39915 , n39972 , n39973 );
not ( n39975 , n39790 );
xor ( n39976 , n39975 , n39908 );
and ( n39977 , n39974 , n39976 );
xor ( n39978 , n39963 , n39965 );
xor ( n39979 , n39978 , n39968 );
buf ( n39980 , n39979 );
xor ( n39981 , n39726 , n39860 );
xor ( n39982 , n39860 , n39862 );
not ( n39983 , n39982 );
and ( n39984 , n39981 , n39983 );
and ( n39985 , n39184 , n39984 );
not ( n39986 , n39985 );
xnor ( n39987 , n39986 , n39865 );
and ( n39988 , n39618 , n39335 );
and ( n39989 , n39524 , n39333 );
nor ( n39990 , n39988 , n39989 );
xnor ( n39991 , n39990 , n39300 );
and ( n39992 , n39987 , n39991 );
and ( n39993 , n39875 , n39194 );
and ( n39994 , n39848 , n39192 );
nor ( n39995 , n39993 , n39994 );
xnor ( n39996 , n39995 , n39199 );
and ( n39997 , n39991 , n39996 );
and ( n39998 , n39987 , n39996 );
or ( n39999 , n39992 , n39997 , n39998 );
and ( n40000 , n39271 , n39665 );
and ( n40001 , n39229 , n39663 );
nor ( n40002 , n40000 , n40001 );
xnor ( n40003 , n40002 , n39608 );
and ( n40004 , n39999 , n40003 );
xor ( n40005 , n39866 , n39870 );
xor ( n40006 , n40005 , n39876 );
and ( n40007 , n40003 , n40006 );
and ( n40008 , n39999 , n40006 );
or ( n40009 , n40004 , n40007 , n40008 );
xor ( n40010 , n39823 , n39827 );
xor ( n40011 , n40010 , n39832 );
and ( n40012 , n40009 , n40011 );
xor ( n40013 , n39879 , n39880 );
xor ( n40014 , n40013 , n39885 );
and ( n40015 , n40011 , n40014 );
and ( n40016 , n40009 , n40014 );
or ( n40017 , n40012 , n40015 , n40016 );
and ( n40018 , n39229 , n39795 );
and ( n40019 , n39220 , n39793 );
nor ( n40020 , n40018 , n40019 );
xnor ( n40021 , n40020 , n39729 );
and ( n40022 , n39310 , n39665 );
and ( n40023 , n39271 , n39663 );
nor ( n40024 , n40022 , n40023 );
xnor ( n40025 , n40024 , n39608 );
and ( n40026 , n40021 , n40025 );
and ( n40027 , n39507 , n39384 );
and ( n40028 , n39433 , n39382 );
nor ( n40029 , n40027 , n40028 );
xnor ( n40030 , n40029 , n39367 );
and ( n40031 , n40025 , n40030 );
and ( n40032 , n40021 , n40030 );
or ( n40033 , n40026 , n40031 , n40032 );
and ( n40034 , n39397 , n39532 );
and ( n40035 , n39327 , n39530 );
nor ( n40036 , n40034 , n40035 );
xnor ( n40037 , n40036 , n39497 );
and ( n40038 , n39739 , n39258 );
and ( n40039 , n39657 , n39256 );
nor ( n40040 , n40038 , n40039 );
xnor ( n40041 , n40040 , n39215 );
and ( n40042 , n40037 , n40041 );
not ( n40043 , n39936 );
and ( n40044 , n40041 , n40043 );
and ( n40045 , n40037 , n40043 );
or ( n40046 , n40042 , n40044 , n40045 );
and ( n40047 , n40033 , n40046 );
xor ( n40048 , n39919 , n39923 );
xor ( n40049 , n40048 , n39928 );
and ( n40050 , n40046 , n40049 );
and ( n40051 , n40033 , n40049 );
or ( n40052 , n40047 , n40050 , n40051 );
buf ( n40053 , n1171 );
buf ( n40054 , n40053 );
buf ( n40055 , n1172 );
buf ( n40056 , n40055 );
and ( n40057 , n40054 , n40056 );
not ( n40058 , n40057 );
and ( n40059 , n39862 , n40058 );
not ( n40060 , n40059 );
and ( n40061 , n39935 , n39194 );
and ( n40062 , n39875 , n39192 );
nor ( n40063 , n40061 , n40062 );
xnor ( n40064 , n40063 , n39199 );
and ( n40065 , n40060 , n40064 );
xor ( n40066 , n33665 , n39153 );
buf ( n40067 , n40066 );
buf ( n40068 , n40067 );
buf ( n40069 , n40068 );
and ( n40070 , n40069 , n39186 );
and ( n40071 , n40064 , n40070 );
and ( n40072 , n40060 , n40070 );
or ( n40073 , n40065 , n40071 , n40072 );
xor ( n40074 , n33668 , n39151 );
buf ( n40075 , n40074 );
buf ( n40076 , n40075 );
buf ( n40077 , n40076 );
and ( n40078 , n40077 , n39186 );
buf ( n40079 , n40078 );
and ( n40080 , n39524 , n39384 );
and ( n40081 , n39507 , n39382 );
nor ( n40082 , n40080 , n40081 );
xnor ( n40083 , n40082 , n39367 );
and ( n40084 , n40079 , n40083 );
and ( n40085 , n39848 , n39258 );
and ( n40086 , n39739 , n39256 );
nor ( n40087 , n40085 , n40086 );
xnor ( n40088 , n40087 , n39215 );
and ( n40089 , n40083 , n40088 );
and ( n40090 , n40079 , n40088 );
or ( n40091 , n40084 , n40089 , n40090 );
and ( n40092 , n40073 , n40091 );
xor ( n40093 , n39987 , n39991 );
xor ( n40094 , n40093 , n39996 );
and ( n40095 , n40091 , n40094 );
and ( n40096 , n40073 , n40094 );
or ( n40097 , n40092 , n40095 , n40096 );
xor ( n40098 , n39937 , n39941 );
xor ( n40099 , n40098 , n39946 );
and ( n40100 , n40097 , n40099 );
xor ( n40101 , n39999 , n40003 );
xor ( n40102 , n40101 , n40006 );
and ( n40103 , n40099 , n40102 );
and ( n40104 , n40097 , n40102 );
or ( n40105 , n40100 , n40103 , n40104 );
and ( n40106 , n40052 , n40105 );
xor ( n40107 , n39931 , n39949 );
xor ( n40108 , n40107 , n39952 );
and ( n40109 , n40105 , n40108 );
and ( n40110 , n40052 , n40108 );
or ( n40111 , n40106 , n40109 , n40110 );
and ( n40112 , n40017 , n40111 );
xor ( n40113 , n39955 , n39957 );
xor ( n40114 , n40113 , n39960 );
and ( n40115 , n40111 , n40114 );
and ( n40116 , n40017 , n40114 );
or ( n40117 , n40112 , n40115 , n40116 );
and ( n40118 , n39979 , n40117 );
buf ( n40119 , n40117 );
or ( n40120 , n39980 , n40118 , n40119 );
not ( n40121 , n39914 );
xor ( n40122 , n40121 , n39971 );
and ( n40123 , n40120 , n40122 );
xor ( n40124 , n40017 , n40111 );
xor ( n40125 , n40124 , n40114 );
buf ( n40126 , n40125 );
and ( n40127 , n39220 , n39984 );
and ( n40128 , n39184 , n39982 );
nor ( n40129 , n40127 , n40128 );
xnor ( n40130 , n40129 , n39865 );
and ( n40131 , n39327 , n39665 );
and ( n40132 , n39310 , n39663 );
nor ( n40133 , n40131 , n40132 );
xnor ( n40134 , n40133 , n39608 );
and ( n40135 , n40130 , n40134 );
and ( n40136 , n39657 , n39335 );
and ( n40137 , n39618 , n39333 );
nor ( n40138 , n40136 , n40137 );
xnor ( n40139 , n40138 , n39300 );
and ( n40140 , n40134 , n40139 );
and ( n40141 , n40130 , n40139 );
or ( n40142 , n40135 , n40140 , n40141 );
xor ( n40143 , n40021 , n40025 );
xor ( n40144 , n40143 , n40030 );
and ( n40145 , n40142 , n40144 );
xor ( n40146 , n40037 , n40041 );
xor ( n40147 , n40146 , n40043 );
and ( n40148 , n40144 , n40147 );
and ( n40149 , n40142 , n40147 );
or ( n40150 , n40145 , n40148 , n40149 );
and ( n40151 , n39271 , n39795 );
and ( n40152 , n39229 , n39793 );
nor ( n40153 , n40151 , n40152 );
xnor ( n40154 , n40153 , n39729 );
and ( n40155 , n39433 , n39532 );
and ( n40156 , n39397 , n39530 );
nor ( n40157 , n40155 , n40156 );
xnor ( n40158 , n40157 , n39497 );
and ( n40159 , n40154 , n40158 );
xor ( n40160 , n40060 , n40064 );
xor ( n40161 , n40160 , n40070 );
and ( n40162 , n40158 , n40161 );
and ( n40163 , n40154 , n40161 );
or ( n40164 , n40159 , n40162 , n40163 );
xor ( n40165 , n39862 , n40054 );
xor ( n40166 , n40054 , n40056 );
not ( n40167 , n40166 );
and ( n40168 , n40165 , n40167 );
and ( n40169 , n39184 , n40168 );
not ( n40170 , n40169 );
xnor ( n40171 , n40170 , n40059 );
and ( n40172 , n39875 , n39258 );
and ( n40173 , n39848 , n39256 );
nor ( n40174 , n40172 , n40173 );
xnor ( n40175 , n40174 , n39215 );
and ( n40176 , n40171 , n40175 );
and ( n40177 , n40069 , n39194 );
and ( n40178 , n39935 , n39192 );
nor ( n40179 , n40177 , n40178 );
xnor ( n40180 , n40179 , n39199 );
and ( n40181 , n40175 , n40180 );
and ( n40182 , n40171 , n40180 );
or ( n40183 , n40176 , n40181 , n40182 );
and ( n40184 , n39618 , n39384 );
and ( n40185 , n39524 , n39382 );
nor ( n40186 , n40184 , n40185 );
xnor ( n40187 , n40186 , n39367 );
and ( n40188 , n39739 , n39335 );
and ( n40189 , n39657 , n39333 );
nor ( n40190 , n40188 , n40189 );
xnor ( n40191 , n40190 , n39300 );
and ( n40192 , n40187 , n40191 );
not ( n40193 , n40078 );
and ( n40194 , n40191 , n40193 );
and ( n40195 , n40187 , n40193 );
or ( n40196 , n40192 , n40194 , n40195 );
and ( n40197 , n40183 , n40196 );
xor ( n40198 , n40079 , n40083 );
xor ( n40199 , n40198 , n40088 );
and ( n40200 , n40196 , n40199 );
and ( n40201 , n40183 , n40199 );
or ( n40202 , n40197 , n40200 , n40201 );
and ( n40203 , n40164 , n40202 );
xor ( n40204 , n40073 , n40091 );
xor ( n40205 , n40204 , n40094 );
and ( n40206 , n40202 , n40205 );
and ( n40207 , n40164 , n40205 );
or ( n40208 , n40203 , n40206 , n40207 );
and ( n40209 , n40150 , n40208 );
xor ( n40210 , n40033 , n40046 );
xor ( n40211 , n40210 , n40049 );
and ( n40212 , n40208 , n40211 );
and ( n40213 , n40150 , n40211 );
or ( n40214 , n40209 , n40212 , n40213 );
xor ( n40215 , n40009 , n40011 );
xor ( n40216 , n40215 , n40014 );
and ( n40217 , n40214 , n40216 );
xor ( n40218 , n40052 , n40105 );
xor ( n40219 , n40218 , n40108 );
and ( n40220 , n40216 , n40219 );
and ( n40221 , n40214 , n40219 );
or ( n40222 , n40217 , n40220 , n40221 );
and ( n40223 , n40125 , n40222 );
buf ( n40224 , n40222 );
or ( n40225 , n40126 , n40223 , n40224 );
not ( n40226 , n39979 );
xor ( n40227 , n40226 , n40117 );
and ( n40228 , n40225 , n40227 );
xor ( n40229 , n40214 , n40216 );
xor ( n40230 , n40229 , n40219 );
buf ( n40231 , n40230 );
and ( n40232 , n39229 , n39984 );
and ( n40233 , n39220 , n39982 );
nor ( n40234 , n40232 , n40233 );
xnor ( n40235 , n40234 , n39865 );
and ( n40236 , n39397 , n39665 );
and ( n40237 , n39327 , n39663 );
nor ( n40238 , n40236 , n40237 );
xnor ( n40239 , n40238 , n39608 );
and ( n40240 , n40235 , n40239 );
and ( n40241 , n39507 , n39532 );
and ( n40242 , n39433 , n39530 );
nor ( n40243 , n40241 , n40242 );
xnor ( n40244 , n40243 , n39497 );
and ( n40245 , n40239 , n40244 );
and ( n40246 , n40235 , n40244 );
or ( n40247 , n40240 , n40245 , n40246 );
xor ( n40248 , n40130 , n40134 );
xor ( n40249 , n40248 , n40139 );
and ( n40250 , n40247 , n40249 );
xor ( n40251 , n40154 , n40158 );
xor ( n40252 , n40251 , n40161 );
and ( n40253 , n40249 , n40252 );
and ( n40254 , n40247 , n40252 );
or ( n40255 , n40250 , n40253 , n40254 );
buf ( n40256 , n1173 );
buf ( n40257 , n40256 );
buf ( n40258 , n1174 );
buf ( n40259 , n40258 );
and ( n40260 , n40257 , n40259 );
not ( n40261 , n40260 );
and ( n40262 , n40056 , n40261 );
not ( n40263 , n40262 );
and ( n40264 , n40077 , n39194 );
and ( n40265 , n40069 , n39192 );
nor ( n40266 , n40264 , n40265 );
xnor ( n40267 , n40266 , n39199 );
and ( n40268 , n40263 , n40267 );
xor ( n40269 , n33670 , n39150 );
buf ( n40270 , n40269 );
buf ( n40271 , n40270 );
buf ( n40272 , n40271 );
and ( n40273 , n40272 , n39186 );
and ( n40274 , n40267 , n40273 );
and ( n40275 , n40263 , n40273 );
or ( n40276 , n40268 , n40274 , n40275 );
xor ( n40277 , n33671 , n39149 );
buf ( n40278 , n40277 );
buf ( n40279 , n40278 );
buf ( n40280 , n40279 );
and ( n40281 , n40280 , n39186 );
buf ( n40282 , n40281 );
and ( n40283 , n39848 , n39335 );
and ( n40284 , n39739 , n39333 );
nor ( n40285 , n40283 , n40284 );
xnor ( n40286 , n40285 , n39300 );
and ( n40287 , n40282 , n40286 );
and ( n40288 , n39935 , n39258 );
and ( n40289 , n39875 , n39256 );
nor ( n40290 , n40288 , n40289 );
xnor ( n40291 , n40290 , n39215 );
and ( n40292 , n40286 , n40291 );
and ( n40293 , n40282 , n40291 );
or ( n40294 , n40287 , n40292 , n40293 );
and ( n40295 , n40276 , n40294 );
and ( n40296 , n39310 , n39795 );
and ( n40297 , n39271 , n39793 );
nor ( n40298 , n40296 , n40297 );
xnor ( n40299 , n40298 , n39729 );
and ( n40300 , n40294 , n40299 );
and ( n40301 , n40276 , n40299 );
or ( n40302 , n40295 , n40300 , n40301 );
and ( n40303 , n39220 , n40168 );
and ( n40304 , n39184 , n40166 );
nor ( n40305 , n40303 , n40304 );
xnor ( n40306 , n40305 , n40059 );
and ( n40307 , n39433 , n39665 );
and ( n40308 , n39397 , n39663 );
nor ( n40309 , n40307 , n40308 );
xnor ( n40310 , n40309 , n39608 );
and ( n40311 , n40306 , n40310 );
xor ( n40312 , n40263 , n40267 );
xor ( n40313 , n40312 , n40273 );
and ( n40314 , n40310 , n40313 );
and ( n40315 , n40306 , n40313 );
or ( n40316 , n40311 , n40314 , n40315 );
xor ( n40317 , n40171 , n40175 );
xor ( n40318 , n40317 , n40180 );
and ( n40319 , n40316 , n40318 );
xor ( n40320 , n40187 , n40191 );
xor ( n40321 , n40320 , n40193 );
and ( n40322 , n40318 , n40321 );
and ( n40323 , n40316 , n40321 );
or ( n40324 , n40319 , n40322 , n40323 );
and ( n40325 , n40302 , n40324 );
xor ( n40326 , n40183 , n40196 );
xor ( n40327 , n40326 , n40199 );
and ( n40328 , n40324 , n40327 );
and ( n40329 , n40302 , n40327 );
or ( n40330 , n40325 , n40328 , n40329 );
and ( n40331 , n40255 , n40330 );
xor ( n40332 , n40142 , n40144 );
xor ( n40333 , n40332 , n40147 );
and ( n40334 , n40330 , n40333 );
and ( n40335 , n40255 , n40333 );
or ( n40336 , n40331 , n40334 , n40335 );
xor ( n40337 , n40097 , n40099 );
xor ( n40338 , n40337 , n40102 );
and ( n40339 , n40336 , n40338 );
xor ( n40340 , n40150 , n40208 );
xor ( n40341 , n40340 , n40211 );
and ( n40342 , n40338 , n40341 );
and ( n40343 , n40336 , n40341 );
or ( n40344 , n40339 , n40342 , n40343 );
and ( n40345 , n40230 , n40344 );
buf ( n40346 , n40344 );
or ( n40347 , n40231 , n40345 , n40346 );
not ( n40348 , n40125 );
xor ( n40349 , n40348 , n40222 );
and ( n40350 , n40347 , n40349 );
xor ( n40351 , n40336 , n40338 );
xor ( n40352 , n40351 , n40341 );
buf ( n40353 , n40352 );
and ( n40354 , n39327 , n39795 );
and ( n40355 , n39310 , n39793 );
nor ( n40356 , n40354 , n40355 );
xnor ( n40357 , n40356 , n39729 );
and ( n40358 , n39524 , n39532 );
and ( n40359 , n39507 , n39530 );
nor ( n40360 , n40358 , n40359 );
xnor ( n40361 , n40360 , n39497 );
and ( n40362 , n40357 , n40361 );
and ( n40363 , n39657 , n39384 );
and ( n40364 , n39618 , n39382 );
nor ( n40365 , n40363 , n40364 );
xnor ( n40366 , n40365 , n39367 );
and ( n40367 , n40361 , n40366 );
and ( n40368 , n40357 , n40366 );
or ( n40369 , n40362 , n40367 , n40368 );
xor ( n40370 , n40235 , n40239 );
xor ( n40371 , n40370 , n40244 );
and ( n40372 , n40369 , n40371 );
xor ( n40373 , n40276 , n40294 );
xor ( n40374 , n40373 , n40299 );
and ( n40375 , n40371 , n40374 );
and ( n40376 , n40369 , n40374 );
or ( n40377 , n40372 , n40375 , n40376 );
xor ( n40378 , n40247 , n40249 );
xor ( n40379 , n40378 , n40252 );
and ( n40380 , n40377 , n40379 );
xor ( n40381 , n40302 , n40324 );
xor ( n40382 , n40381 , n40327 );
and ( n40383 , n40379 , n40382 );
and ( n40384 , n40377 , n40382 );
or ( n40385 , n40380 , n40383 , n40384 );
xor ( n40386 , n40164 , n40202 );
xor ( n40387 , n40386 , n40205 );
and ( n40388 , n40385 , n40387 );
xor ( n40389 , n40255 , n40330 );
xor ( n40390 , n40389 , n40333 );
and ( n40391 , n40387 , n40390 );
and ( n40392 , n40385 , n40390 );
or ( n40393 , n40388 , n40391 , n40392 );
and ( n40394 , n40352 , n40393 );
buf ( n40395 , n40393 );
or ( n40396 , n40353 , n40394 , n40395 );
not ( n40397 , n40230 );
xor ( n40398 , n40397 , n40344 );
and ( n40399 , n40396 , n40398 );
xor ( n40400 , n40385 , n40387 );
xor ( n40401 , n40400 , n40390 );
buf ( n40402 , n40401 );
xor ( n40403 , n40056 , n40257 );
xor ( n40404 , n40257 , n40259 );
not ( n40405 , n40404 );
and ( n40406 , n40403 , n40405 );
and ( n40407 , n39184 , n40406 );
not ( n40408 , n40407 );
xnor ( n40409 , n40408 , n40262 );
and ( n40410 , n39618 , n39532 );
and ( n40411 , n39524 , n39530 );
nor ( n40412 , n40410 , n40411 );
xnor ( n40413 , n40412 , n39497 );
and ( n40414 , n40409 , n40413 );
and ( n40415 , n39875 , n39335 );
and ( n40416 , n39848 , n39333 );
nor ( n40417 , n40415 , n40416 );
xnor ( n40418 , n40417 , n39300 );
and ( n40419 , n40413 , n40418 );
and ( n40420 , n40409 , n40418 );
or ( n40421 , n40414 , n40419 , n40420 );
and ( n40422 , n39229 , n40168 );
and ( n40423 , n39220 , n40166 );
nor ( n40424 , n40422 , n40423 );
xnor ( n40425 , n40424 , n40059 );
and ( n40426 , n39310 , n39984 );
and ( n40427 , n39271 , n39982 );
nor ( n40428 , n40426 , n40427 );
xnor ( n40429 , n40428 , n39865 );
and ( n40430 , n40425 , n40429 );
and ( n40431 , n39507 , n39665 );
and ( n40432 , n39433 , n39663 );
nor ( n40433 , n40431 , n40432 );
xnor ( n40434 , n40433 , n39608 );
and ( n40435 , n40429 , n40434 );
and ( n40436 , n40425 , n40434 );
or ( n40437 , n40430 , n40435 , n40436 );
and ( n40438 , n40421 , n40437 );
buf ( n40439 , n1175 );
buf ( n40440 , n40439 );
buf ( n40441 , n1176 );
buf ( n40442 , n40441 );
and ( n40443 , n40440 , n40442 );
not ( n40444 , n40443 );
and ( n40445 , n40259 , n40444 );
not ( n40446 , n40445 );
and ( n40447 , n40280 , n39194 );
and ( n40448 , n40272 , n39192 );
nor ( n40449 , n40447 , n40448 );
xnor ( n40450 , n40449 , n39199 );
and ( n40451 , n40446 , n40450 );
xor ( n40452 , n35693 , n39147 );
buf ( n40453 , n40452 );
buf ( n40454 , n40453 );
buf ( n40455 , n40454 );
and ( n40456 , n40455 , n39186 );
and ( n40457 , n40450 , n40456 );
and ( n40458 , n40446 , n40456 );
or ( n40459 , n40451 , n40457 , n40458 );
and ( n40460 , n39397 , n39795 );
and ( n40461 , n39327 , n39793 );
nor ( n40462 , n40460 , n40461 );
xnor ( n40463 , n40462 , n39729 );
and ( n40464 , n40459 , n40463 );
and ( n40465 , n39739 , n39384 );
and ( n40466 , n39657 , n39382 );
nor ( n40467 , n40465 , n40466 );
xnor ( n40468 , n40467 , n39367 );
and ( n40469 , n40463 , n40468 );
and ( n40470 , n40459 , n40468 );
or ( n40471 , n40464 , n40469 , n40470 );
and ( n40472 , n40437 , n40471 );
and ( n40473 , n40421 , n40471 );
or ( n40474 , n40438 , n40472 , n40473 );
and ( n40475 , n40069 , n39258 );
and ( n40476 , n39935 , n39256 );
nor ( n40477 , n40475 , n40476 );
xnor ( n40478 , n40477 , n39215 );
and ( n40479 , n40272 , n39194 );
and ( n40480 , n40077 , n39192 );
nor ( n40481 , n40479 , n40480 );
xnor ( n40482 , n40481 , n39199 );
and ( n40483 , n40478 , n40482 );
not ( n40484 , n40281 );
and ( n40485 , n40482 , n40484 );
and ( n40486 , n40478 , n40484 );
or ( n40487 , n40483 , n40485 , n40486 );
and ( n40488 , n39271 , n39984 );
and ( n40489 , n39229 , n39982 );
nor ( n40490 , n40488 , n40489 );
xnor ( n40491 , n40490 , n39865 );
and ( n40492 , n40487 , n40491 );
xor ( n40493 , n40282 , n40286 );
xor ( n40494 , n40493 , n40291 );
and ( n40495 , n40491 , n40494 );
and ( n40496 , n40487 , n40494 );
or ( n40497 , n40492 , n40495 , n40496 );
and ( n40498 , n40474 , n40497 );
xor ( n40499 , n40316 , n40318 );
xor ( n40500 , n40499 , n40321 );
and ( n40501 , n40497 , n40500 );
and ( n40502 , n40474 , n40500 );
or ( n40503 , n40498 , n40501 , n40502 );
and ( n40504 , n40455 , n39194 );
and ( n40505 , n40280 , n39192 );
nor ( n40506 , n40504 , n40505 );
xnor ( n40507 , n40506 , n39199 );
buf ( n40508 , n40507 );
and ( n40509 , n39935 , n39335 );
and ( n40510 , n39875 , n39333 );
nor ( n40511 , n40509 , n40510 );
xnor ( n40512 , n40511 , n39300 );
and ( n40513 , n40508 , n40512 );
and ( n40514 , n40077 , n39258 );
and ( n40515 , n40069 , n39256 );
nor ( n40516 , n40514 , n40515 );
xnor ( n40517 , n40516 , n39215 );
and ( n40518 , n40512 , n40517 );
and ( n40519 , n40508 , n40517 );
or ( n40520 , n40513 , n40518 , n40519 );
and ( n40521 , n39524 , n39665 );
and ( n40522 , n39507 , n39663 );
nor ( n40523 , n40521 , n40522 );
xnor ( n40524 , n40523 , n39608 );
and ( n40525 , n39848 , n39384 );
and ( n40526 , n39739 , n39382 );
nor ( n40527 , n40525 , n40526 );
xnor ( n40528 , n40527 , n39367 );
and ( n40529 , n40524 , n40528 );
xor ( n40530 , n40446 , n40450 );
xor ( n40531 , n40530 , n40456 );
and ( n40532 , n40528 , n40531 );
and ( n40533 , n40524 , n40531 );
or ( n40534 , n40529 , n40532 , n40533 );
and ( n40535 , n40520 , n40534 );
xor ( n40536 , n40478 , n40482 );
xor ( n40537 , n40536 , n40484 );
and ( n40538 , n40534 , n40537 );
and ( n40539 , n40520 , n40537 );
or ( n40540 , n40535 , n40538 , n40539 );
xor ( n40541 , n40357 , n40361 );
xor ( n40542 , n40541 , n40366 );
and ( n40543 , n40540 , n40542 );
xor ( n40544 , n40306 , n40310 );
xor ( n40545 , n40544 , n40313 );
and ( n40546 , n40542 , n40545 );
and ( n40547 , n40540 , n40545 );
or ( n40548 , n40543 , n40546 , n40547 );
and ( n40549 , n39220 , n40406 );
and ( n40550 , n39184 , n40404 );
nor ( n40551 , n40549 , n40550 );
xnor ( n40552 , n40551 , n40262 );
and ( n40553 , n39327 , n39984 );
and ( n40554 , n39310 , n39982 );
nor ( n40555 , n40553 , n40554 );
xnor ( n40556 , n40555 , n39865 );
and ( n40557 , n40552 , n40556 );
and ( n40558 , n39657 , n39532 );
and ( n40559 , n39618 , n39530 );
nor ( n40560 , n40558 , n40559 );
xnor ( n40561 , n40560 , n39497 );
and ( n40562 , n40556 , n40561 );
and ( n40563 , n40552 , n40561 );
or ( n40564 , n40557 , n40562 , n40563 );
and ( n40565 , n40272 , n39258 );
and ( n40566 , n40077 , n39256 );
nor ( n40567 , n40565 , n40566 );
xnor ( n40568 , n40567 , n39215 );
not ( n40569 , n40507 );
and ( n40570 , n40568 , n40569 );
xor ( n40571 , n35695 , n39146 );
buf ( n40572 , n40571 );
buf ( n40573 , n40572 );
buf ( n40574 , n40573 );
and ( n40575 , n40574 , n39186 );
and ( n40576 , n40569 , n40575 );
and ( n40577 , n40568 , n40575 );
or ( n40578 , n40570 , n40576 , n40577 );
and ( n40579 , n39271 , n40168 );
and ( n40580 , n39229 , n40166 );
nor ( n40581 , n40579 , n40580 );
xnor ( n40582 , n40581 , n40059 );
and ( n40583 , n40578 , n40582 );
and ( n40584 , n39433 , n39795 );
and ( n40585 , n39397 , n39793 );
nor ( n40586 , n40584 , n40585 );
xnor ( n40587 , n40586 , n39729 );
and ( n40588 , n40582 , n40587 );
and ( n40589 , n40578 , n40587 );
or ( n40590 , n40583 , n40588 , n40589 );
and ( n40591 , n40564 , n40590 );
xor ( n40592 , n40409 , n40413 );
xor ( n40593 , n40592 , n40418 );
and ( n40594 , n40590 , n40593 );
and ( n40595 , n40564 , n40593 );
or ( n40596 , n40591 , n40594 , n40595 );
xor ( n40597 , n40421 , n40437 );
xor ( n40598 , n40597 , n40471 );
and ( n40599 , n40596 , n40598 );
xor ( n40600 , n40487 , n40491 );
xor ( n40601 , n40600 , n40494 );
and ( n40602 , n40598 , n40601 );
and ( n40603 , n40596 , n40601 );
or ( n40604 , n40599 , n40602 , n40603 );
and ( n40605 , n40548 , n40604 );
xor ( n40606 , n40369 , n40371 );
xor ( n40607 , n40606 , n40374 );
and ( n40608 , n40604 , n40607 );
and ( n40609 , n40548 , n40607 );
or ( n40610 , n40605 , n40608 , n40609 );
and ( n40611 , n40503 , n40610 );
xor ( n40612 , n40377 , n40379 );
xor ( n40613 , n40612 , n40382 );
and ( n40614 , n40610 , n40613 );
and ( n40615 , n40503 , n40613 );
or ( n40616 , n40611 , n40614 , n40615 );
and ( n40617 , n40401 , n40616 );
buf ( n40618 , n40616 );
or ( n40619 , n40402 , n40617 , n40618 );
not ( n40620 , n40352 );
xor ( n40621 , n40620 , n40393 );
and ( n40622 , n40619 , n40621 );
xor ( n40623 , n40503 , n40610 );
xor ( n40624 , n40623 , n40613 );
buf ( n40625 , n40624 );
xor ( n40626 , n40425 , n40429 );
xor ( n40627 , n40626 , n40434 );
xor ( n40628 , n40459 , n40463 );
xor ( n40629 , n40628 , n40468 );
and ( n40630 , n40627 , n40629 );
xor ( n40631 , n40520 , n40534 );
xor ( n40632 , n40631 , n40537 );
and ( n40633 , n40629 , n40632 );
and ( n40634 , n40627 , n40632 );
or ( n40635 , n40630 , n40633 , n40634 );
xor ( n40636 , n40540 , n40542 );
xor ( n40637 , n40636 , n40545 );
and ( n40638 , n40635 , n40637 );
xor ( n40639 , n40596 , n40598 );
xor ( n40640 , n40639 , n40601 );
and ( n40641 , n40637 , n40640 );
and ( n40642 , n40635 , n40640 );
or ( n40643 , n40638 , n40641 , n40642 );
xor ( n40644 , n40474 , n40497 );
xor ( n40645 , n40644 , n40500 );
and ( n40646 , n40643 , n40645 );
xor ( n40647 , n40548 , n40604 );
xor ( n40648 , n40647 , n40607 );
and ( n40649 , n40645 , n40648 );
and ( n40650 , n40643 , n40648 );
or ( n40651 , n40646 , n40649 , n40650 );
and ( n40652 , n40624 , n40651 );
buf ( n40653 , n40651 );
or ( n40654 , n40625 , n40652 , n40653 );
not ( n40655 , n40401 );
xor ( n40656 , n40655 , n40616 );
and ( n40657 , n40654 , n40656 );
not ( n40658 , n40624 );
xor ( n40659 , n40658 , n40651 );
xor ( n40660 , n40643 , n40645 );
xor ( n40661 , n40660 , n40648 );
buf ( n40662 , n40661 );
xor ( n40663 , n40259 , n40440 );
xor ( n40664 , n40440 , n40442 );
not ( n40665 , n40664 );
and ( n40666 , n40663 , n40665 );
and ( n40667 , n39184 , n40666 );
not ( n40668 , n40667 );
xnor ( n40669 , n40668 , n40445 );
and ( n40670 , n39618 , n39665 );
and ( n40671 , n39524 , n39663 );
nor ( n40672 , n40670 , n40671 );
xnor ( n40673 , n40672 , n39608 );
and ( n40674 , n40669 , n40673 );
and ( n40675 , n39739 , n39532 );
and ( n40676 , n39657 , n39530 );
nor ( n40677 , n40675 , n40676 );
xnor ( n40678 , n40677 , n39497 );
and ( n40679 , n40673 , n40678 );
and ( n40680 , n40669 , n40678 );
or ( n40681 , n40674 , n40679 , n40680 );
buf ( n40682 , n1177 );
buf ( n40683 , n40682 );
buf ( n40684 , n1178 );
buf ( n40685 , n40684 );
and ( n40686 , n40683 , n40685 );
not ( n40687 , n40686 );
and ( n40688 , n40442 , n40687 );
not ( n40689 , n40688 );
and ( n40690 , n40574 , n39194 );
and ( n40691 , n40455 , n39192 );
nor ( n40692 , n40690 , n40691 );
xnor ( n40693 , n40692 , n39199 );
and ( n40694 , n40689 , n40693 );
xor ( n40695 , n35697 , n39145 );
buf ( n40696 , n40695 );
buf ( n40697 , n40696 );
buf ( n40698 , n40697 );
and ( n40699 , n40698 , n39186 );
and ( n40700 , n40693 , n40699 );
and ( n40701 , n40689 , n40699 );
or ( n40702 , n40694 , n40700 , n40701 );
and ( n40703 , n39875 , n39384 );
and ( n40704 , n39848 , n39382 );
nor ( n40705 , n40703 , n40704 );
xnor ( n40706 , n40705 , n39367 );
and ( n40707 , n40702 , n40706 );
and ( n40708 , n40069 , n39335 );
and ( n40709 , n39935 , n39333 );
nor ( n40710 , n40708 , n40709 );
xnor ( n40711 , n40710 , n39300 );
and ( n40712 , n40706 , n40711 );
and ( n40713 , n40702 , n40711 );
or ( n40714 , n40707 , n40712 , n40713 );
and ( n40715 , n40681 , n40714 );
xor ( n40716 , n40508 , n40512 );
xor ( n40717 , n40716 , n40517 );
and ( n40718 , n40714 , n40717 );
and ( n40719 , n40681 , n40717 );
or ( n40720 , n40715 , n40718 , n40719 );
and ( n40721 , n39229 , n40406 );
and ( n40722 , n39220 , n40404 );
nor ( n40723 , n40721 , n40722 );
xnor ( n40724 , n40723 , n40262 );
and ( n40725 , n39397 , n39984 );
and ( n40726 , n39327 , n39982 );
nor ( n40727 , n40725 , n40726 );
xnor ( n40728 , n40727 , n39865 );
and ( n40729 , n40724 , n40728 );
and ( n40730 , n39507 , n39795 );
and ( n40731 , n39433 , n39793 );
nor ( n40732 , n40730 , n40731 );
xnor ( n40733 , n40732 , n39729 );
and ( n40734 , n40728 , n40733 );
and ( n40735 , n40724 , n40733 );
or ( n40736 , n40729 , n40734 , n40735 );
xor ( n40737 , n40578 , n40582 );
xor ( n40738 , n40737 , n40587 );
and ( n40739 , n40736 , n40738 );
xor ( n40740 , n40524 , n40528 );
xor ( n40741 , n40740 , n40531 );
and ( n40742 , n40738 , n40741 );
and ( n40743 , n40736 , n40741 );
or ( n40744 , n40739 , n40742 , n40743 );
and ( n40745 , n40720 , n40744 );
xor ( n40746 , n40564 , n40590 );
xor ( n40747 , n40746 , n40593 );
and ( n40748 , n40744 , n40747 );
and ( n40749 , n40720 , n40747 );
or ( n40750 , n40745 , n40748 , n40749 );
and ( n40751 , n39524 , n39795 );
and ( n40752 , n39507 , n39793 );
nor ( n40753 , n40751 , n40752 );
xnor ( n40754 , n40753 , n39729 );
and ( n40755 , n39848 , n39532 );
and ( n40756 , n39739 , n39530 );
nor ( n40757 , n40755 , n40756 );
xnor ( n40758 , n40757 , n39497 );
and ( n40759 , n40754 , n40758 );
and ( n40760 , n39935 , n39384 );
and ( n40761 , n39875 , n39382 );
nor ( n40762 , n40760 , n40761 );
xnor ( n40763 , n40762 , n39367 );
and ( n40764 , n40758 , n40763 );
and ( n40765 , n40754 , n40763 );
or ( n40766 , n40759 , n40764 , n40765 );
and ( n40767 , n39327 , n40168 );
and ( n40768 , n39310 , n40166 );
nor ( n40769 , n40767 , n40768 );
xnor ( n40770 , n40769 , n40059 );
and ( n40771 , n39657 , n39665 );
and ( n40772 , n39618 , n39663 );
nor ( n40773 , n40771 , n40772 );
xnor ( n40774 , n40773 , n39608 );
and ( n40775 , n40770 , n40774 );
xor ( n40776 , n40689 , n40693 );
xor ( n40777 , n40776 , n40699 );
and ( n40778 , n40774 , n40777 );
and ( n40779 , n40770 , n40777 );
or ( n40780 , n40775 , n40778 , n40779 );
and ( n40781 , n40766 , n40780 );
xor ( n40782 , n40702 , n40706 );
xor ( n40783 , n40782 , n40711 );
and ( n40784 , n40780 , n40783 );
and ( n40785 , n40766 , n40783 );
or ( n40786 , n40781 , n40784 , n40785 );
and ( n40787 , n40455 , n39258 );
and ( n40788 , n40280 , n39256 );
nor ( n40789 , n40787 , n40788 );
xnor ( n40790 , n40789 , n39215 );
buf ( n40791 , n40790 );
and ( n40792 , n40077 , n39335 );
and ( n40793 , n40069 , n39333 );
nor ( n40794 , n40792 , n40793 );
xnor ( n40795 , n40794 , n39300 );
and ( n40796 , n40791 , n40795 );
and ( n40797 , n40280 , n39258 );
and ( n40798 , n40272 , n39256 );
nor ( n40799 , n40797 , n40798 );
xnor ( n40800 , n40799 , n39215 );
and ( n40801 , n40795 , n40800 );
and ( n40802 , n40791 , n40800 );
or ( n40803 , n40796 , n40801 , n40802 );
and ( n40804 , n39310 , n40168 );
and ( n40805 , n39271 , n40166 );
nor ( n40806 , n40804 , n40805 );
xnor ( n40807 , n40806 , n40059 );
and ( n40808 , n40803 , n40807 );
xor ( n40809 , n40568 , n40569 );
xor ( n40810 , n40809 , n40575 );
and ( n40811 , n40807 , n40810 );
and ( n40812 , n40803 , n40810 );
or ( n40813 , n40808 , n40811 , n40812 );
and ( n40814 , n40786 , n40813 );
xor ( n40815 , n40552 , n40556 );
xor ( n40816 , n40815 , n40561 );
and ( n40817 , n40813 , n40816 );
and ( n40818 , n40786 , n40816 );
or ( n40819 , n40814 , n40817 , n40818 );
and ( n40820 , n39220 , n40666 );
and ( n40821 , n39184 , n40664 );
nor ( n40822 , n40820 , n40821 );
xnor ( n40823 , n40822 , n40445 );
and ( n40824 , n39271 , n40406 );
and ( n40825 , n39229 , n40404 );
nor ( n40826 , n40824 , n40825 );
xnor ( n40827 , n40826 , n40262 );
and ( n40828 , n40823 , n40827 );
and ( n40829 , n39433 , n39984 );
and ( n40830 , n39397 , n39982 );
nor ( n40831 , n40829 , n40830 );
xnor ( n40832 , n40831 , n39865 );
and ( n40833 , n40827 , n40832 );
and ( n40834 , n40823 , n40832 );
or ( n40835 , n40828 , n40833 , n40834 );
xor ( n40836 , n40669 , n40673 );
xor ( n40837 , n40836 , n40678 );
and ( n40838 , n40835 , n40837 );
xor ( n40839 , n40724 , n40728 );
xor ( n40840 , n40839 , n40733 );
and ( n40841 , n40837 , n40840 );
and ( n40842 , n40835 , n40840 );
or ( n40843 , n40838 , n40841 , n40842 );
xor ( n40844 , n40681 , n40714 );
xor ( n40845 , n40844 , n40717 );
and ( n40846 , n40843 , n40845 );
xor ( n40847 , n40736 , n40738 );
xor ( n40848 , n40847 , n40741 );
and ( n40849 , n40845 , n40848 );
and ( n40850 , n40843 , n40848 );
or ( n40851 , n40846 , n40849 , n40850 );
and ( n40852 , n40819 , n40851 );
xor ( n40853 , n40627 , n40629 );
xor ( n40854 , n40853 , n40632 );
and ( n40855 , n40851 , n40854 );
and ( n40856 , n40819 , n40854 );
or ( n40857 , n40852 , n40855 , n40856 );
and ( n40858 , n40750 , n40857 );
xor ( n40859 , n40635 , n40637 );
xor ( n40860 , n40859 , n40640 );
and ( n40861 , n40857 , n40860 );
and ( n40862 , n40750 , n40860 );
or ( n40863 , n40858 , n40861 , n40862 );
and ( n40864 , n40661 , n40863 );
buf ( n40865 , n40863 );
or ( n40866 , n40662 , n40864 , n40865 );
and ( n40867 , n40659 , n40866 );
not ( n40868 , n40661 );
xor ( n40869 , n40868 , n40863 );
xor ( n40870 , n40750 , n40857 );
xor ( n40871 , n40870 , n40860 );
buf ( n40872 , n40871 );
xor ( n40873 , n40754 , n40758 );
xor ( n40874 , n40873 , n40763 );
xor ( n40875 , n40823 , n40827 );
xor ( n40876 , n40875 , n40832 );
and ( n40877 , n40874 , n40876 );
xor ( n40878 , n40770 , n40774 );
xor ( n40879 , n40878 , n40777 );
and ( n40880 , n40876 , n40879 );
and ( n40881 , n40874 , n40879 );
or ( n40882 , n40877 , n40880 , n40881 );
xor ( n40883 , n40835 , n40837 );
xor ( n40884 , n40883 , n40840 );
and ( n40885 , n40882 , n40884 );
xor ( n40886 , n40766 , n40780 );
xor ( n40887 , n40886 , n40783 );
and ( n40888 , n40884 , n40887 );
and ( n40889 , n40882 , n40887 );
or ( n40890 , n40885 , n40888 , n40889 );
and ( n40891 , n39229 , n40666 );
and ( n40892 , n39220 , n40664 );
nor ( n40893 , n40891 , n40892 );
xnor ( n40894 , n40893 , n40445 );
and ( n40895 , n39397 , n40168 );
and ( n40896 , n39327 , n40166 );
nor ( n40897 , n40895 , n40896 );
xnor ( n40898 , n40897 , n40059 );
and ( n40899 , n40894 , n40898 );
and ( n40900 , n39507 , n39984 );
and ( n40901 , n39433 , n39982 );
nor ( n40902 , n40900 , n40901 );
xnor ( n40903 , n40902 , n39865 );
and ( n40904 , n40898 , n40903 );
and ( n40905 , n40894 , n40903 );
or ( n40906 , n40899 , n40904 , n40905 );
xor ( n40907 , n35704 , n39140 );
buf ( n40908 , n40907 );
buf ( n40909 , n40908 );
buf ( n40910 , n40909 );
and ( n40911 , n40910 , n39186 );
buf ( n40912 , n40911 );
and ( n40913 , n40280 , n39335 );
and ( n40914 , n40272 , n39333 );
nor ( n40915 , n40913 , n40914 );
xnor ( n40916 , n40915 , n39300 );
and ( n40917 , n40912 , n40916 );
and ( n40918 , n40574 , n39258 );
and ( n40919 , n40455 , n39256 );
nor ( n40920 , n40918 , n40919 );
xnor ( n40921 , n40920 , n39215 );
and ( n40922 , n40916 , n40921 );
and ( n40923 , n40912 , n40921 );
or ( n40924 , n40917 , n40922 , n40923 );
xor ( n40925 , n40442 , n40683 );
xor ( n40926 , n40683 , n40685 );
not ( n40927 , n40926 );
and ( n40928 , n40925 , n40927 );
and ( n40929 , n39184 , n40928 );
not ( n40930 , n40929 );
xnor ( n40931 , n40930 , n40688 );
and ( n40932 , n40924 , n40931 );
and ( n40933 , n39875 , n39532 );
and ( n40934 , n39848 , n39530 );
nor ( n40935 , n40933 , n40934 );
xnor ( n40936 , n40935 , n39497 );
and ( n40937 , n40931 , n40936 );
and ( n40938 , n40924 , n40936 );
or ( n40939 , n40932 , n40937 , n40938 );
and ( n40940 , n40906 , n40939 );
and ( n40941 , n39618 , n39795 );
and ( n40942 , n39524 , n39793 );
nor ( n40943 , n40941 , n40942 );
xnor ( n40944 , n40943 , n39729 );
and ( n40945 , n39739 , n39665 );
and ( n40946 , n39657 , n39663 );
nor ( n40947 , n40945 , n40946 );
xnor ( n40948 , n40947 , n39608 );
and ( n40949 , n40944 , n40948 );
and ( n40950 , n40272 , n39335 );
and ( n40951 , n40077 , n39333 );
nor ( n40952 , n40950 , n40951 );
xnor ( n40953 , n40952 , n39300 );
and ( n40954 , n40698 , n39194 );
and ( n40955 , n40574 , n39192 );
nor ( n40956 , n40954 , n40955 );
xnor ( n40957 , n40956 , n39199 );
xor ( n40958 , n40953 , n40957 );
xor ( n40959 , n35700 , n39143 );
buf ( n40960 , n40959 );
buf ( n40961 , n40960 );
buf ( n40962 , n40961 );
and ( n40963 , n40962 , n39186 );
xor ( n40964 , n40958 , n40963 );
and ( n40965 , n40948 , n40964 );
and ( n40966 , n40944 , n40964 );
or ( n40967 , n40949 , n40965 , n40966 );
and ( n40968 , n40939 , n40967 );
and ( n40969 , n40906 , n40967 );
or ( n40970 , n40940 , n40968 , n40969 );
and ( n40971 , n40953 , n40957 );
and ( n40972 , n40957 , n40963 );
and ( n40973 , n40953 , n40963 );
or ( n40974 , n40971 , n40972 , n40973 );
buf ( n40975 , n1179 );
buf ( n40976 , n40975 );
buf ( n40977 , n1180 );
buf ( n40978 , n40977 );
and ( n40979 , n40976 , n40978 );
not ( n40980 , n40979 );
and ( n40981 , n40685 , n40980 );
not ( n40982 , n40981 );
and ( n40983 , n40962 , n39194 );
and ( n40984 , n40698 , n39192 );
nor ( n40985 , n40983 , n40984 );
xnor ( n40986 , n40985 , n39199 );
and ( n40987 , n40982 , n40986 );
xor ( n40988 , n35701 , n39142 );
buf ( n40989 , n40988 );
buf ( n40990 , n40989 );
buf ( n40991 , n40990 );
and ( n40992 , n40991 , n39186 );
and ( n40993 , n40986 , n40992 );
and ( n40994 , n40982 , n40992 );
or ( n40995 , n40987 , n40993 , n40994 );
and ( n40996 , n40069 , n39384 );
and ( n40997 , n39935 , n39382 );
nor ( n40998 , n40996 , n40997 );
xnor ( n40999 , n40998 , n39367 );
and ( n41000 , n40995 , n40999 );
not ( n41001 , n40790 );
and ( n41002 , n40999 , n41001 );
and ( n41003 , n40995 , n41001 );
or ( n41004 , n41000 , n41002 , n41003 );
and ( n41005 , n40974 , n41004 );
xor ( n41006 , n40791 , n40795 );
xor ( n41007 , n41006 , n40800 );
and ( n41008 , n41004 , n41007 );
and ( n41009 , n40974 , n41007 );
or ( n41010 , n41005 , n41008 , n41009 );
and ( n41011 , n40970 , n41010 );
xor ( n41012 , n40803 , n40807 );
xor ( n41013 , n41012 , n40810 );
and ( n41014 , n41010 , n41013 );
and ( n41015 , n40970 , n41013 );
or ( n41016 , n41011 , n41014 , n41015 );
and ( n41017 , n40890 , n41016 );
xor ( n41018 , n40786 , n40813 );
xor ( n41019 , n41018 , n40816 );
and ( n41020 , n41016 , n41019 );
and ( n41021 , n40890 , n41019 );
or ( n41022 , n41017 , n41020 , n41021 );
xor ( n41023 , n40720 , n40744 );
xor ( n41024 , n41023 , n40747 );
and ( n41025 , n41022 , n41024 );
xor ( n41026 , n40819 , n40851 );
xor ( n41027 , n41026 , n40854 );
and ( n41028 , n41024 , n41027 );
and ( n41029 , n41022 , n41027 );
or ( n41030 , n41025 , n41028 , n41029 );
and ( n41031 , n40871 , n41030 );
buf ( n41032 , n41030 );
or ( n41033 , n40872 , n41031 , n41032 );
and ( n41034 , n40869 , n41033 );
xor ( n41035 , n41022 , n41024 );
xor ( n41036 , n41035 , n41027 );
buf ( n41037 , n41036 );
and ( n41038 , n40455 , n39335 );
and ( n41039 , n40280 , n39333 );
nor ( n41040 , n41038 , n41039 );
xnor ( n41041 , n41040 , n39300 );
and ( n41042 , n40698 , n39258 );
and ( n41043 , n40574 , n39256 );
nor ( n41044 , n41042 , n41043 );
xnor ( n41045 , n41044 , n39215 );
and ( n41046 , n41041 , n41045 );
and ( n41047 , n40991 , n39194 );
and ( n41048 , n40962 , n39192 );
nor ( n41049 , n41047 , n41048 );
xnor ( n41050 , n41049 , n39199 );
and ( n41051 , n41045 , n41050 );
and ( n41052 , n41041 , n41050 );
or ( n41053 , n41046 , n41051 , n41052 );
and ( n41054 , n39935 , n39532 );
and ( n41055 , n39875 , n39530 );
nor ( n41056 , n41054 , n41055 );
xnor ( n41057 , n41056 , n39497 );
and ( n41058 , n41053 , n41057 );
and ( n41059 , n40077 , n39384 );
and ( n41060 , n40069 , n39382 );
nor ( n41061 , n41059 , n41060 );
xnor ( n41062 , n41061 , n39367 );
and ( n41063 , n41057 , n41062 );
and ( n41064 , n41053 , n41062 );
or ( n41065 , n41058 , n41063 , n41064 );
and ( n41066 , n39524 , n39984 );
and ( n41067 , n39507 , n39982 );
nor ( n41068 , n41066 , n41067 );
xnor ( n41069 , n41068 , n39865 );
and ( n41070 , n39848 , n39665 );
and ( n41071 , n39739 , n39663 );
nor ( n41072 , n41070 , n41071 );
xnor ( n41073 , n41072 , n39608 );
and ( n41074 , n41069 , n41073 );
xor ( n41075 , n40982 , n40986 );
xor ( n41076 , n41075 , n40992 );
and ( n41077 , n41073 , n41076 );
and ( n41078 , n41069 , n41076 );
or ( n41079 , n41074 , n41077 , n41078 );
and ( n41080 , n41065 , n41079 );
and ( n41081 , n39310 , n40406 );
and ( n41082 , n39271 , n40404 );
nor ( n41083 , n41081 , n41082 );
xnor ( n41084 , n41083 , n40262 );
and ( n41085 , n41079 , n41084 );
and ( n41086 , n41065 , n41084 );
or ( n41087 , n41080 , n41085 , n41086 );
xor ( n41088 , n36178 , n39137 );
buf ( n41089 , n41088 );
buf ( n41090 , n41089 );
buf ( n41091 , n41090 );
and ( n41092 , n41091 , n39186 );
buf ( n41093 , n41092 );
buf ( n41094 , n1181 );
buf ( n41095 , n41094 );
buf ( n41096 , n1182 );
buf ( n41097 , n41096 );
and ( n41098 , n41095 , n41097 );
not ( n41099 , n41098 );
and ( n41100 , n40978 , n41099 );
not ( n41101 , n41100 );
and ( n41102 , n41093 , n41101 );
xor ( n41103 , n35705 , n39139 );
buf ( n41104 , n41103 );
buf ( n41105 , n41104 );
buf ( n41106 , n41105 );
and ( n41107 , n41106 , n39186 );
and ( n41108 , n41101 , n41107 );
and ( n41109 , n41093 , n41107 );
or ( n41110 , n41102 , n41108 , n41109 );
and ( n41111 , n40272 , n39384 );
and ( n41112 , n40077 , n39382 );
nor ( n41113 , n41111 , n41112 );
xnor ( n41114 , n41113 , n39367 );
and ( n41115 , n41110 , n41114 );
not ( n41116 , n40911 );
and ( n41117 , n41114 , n41116 );
and ( n41118 , n41110 , n41116 );
or ( n41119 , n41115 , n41117 , n41118 );
and ( n41120 , n39220 , n40928 );
and ( n41121 , n39184 , n40926 );
nor ( n41122 , n41120 , n41121 );
xnor ( n41123 , n41122 , n40688 );
and ( n41124 , n41119 , n41123 );
and ( n41125 , n39271 , n40666 );
and ( n41126 , n39229 , n40664 );
nor ( n41127 , n41125 , n41126 );
xnor ( n41128 , n41127 , n40445 );
and ( n41129 , n41123 , n41128 );
and ( n41130 , n41119 , n41128 );
or ( n41131 , n41124 , n41129 , n41130 );
and ( n41132 , n39327 , n40406 );
and ( n41133 , n39310 , n40404 );
nor ( n41134 , n41132 , n41133 );
xnor ( n41135 , n41134 , n40262 );
and ( n41136 , n39657 , n39795 );
and ( n41137 , n39618 , n39793 );
nor ( n41138 , n41136 , n41137 );
xnor ( n41139 , n41138 , n39729 );
and ( n41140 , n41135 , n41139 );
xor ( n41141 , n40912 , n40916 );
xor ( n41142 , n41141 , n40921 );
and ( n41143 , n41139 , n41142 );
and ( n41144 , n41135 , n41142 );
or ( n41145 , n41140 , n41143 , n41144 );
and ( n41146 , n41131 , n41145 );
xor ( n41147 , n40995 , n40999 );
xor ( n41148 , n41147 , n41001 );
and ( n41149 , n41145 , n41148 );
and ( n41150 , n41131 , n41148 );
or ( n41151 , n41146 , n41149 , n41150 );
and ( n41152 , n41087 , n41151 );
xor ( n41153 , n40974 , n41004 );
xor ( n41154 , n41153 , n41007 );
and ( n41155 , n41151 , n41154 );
and ( n41156 , n41087 , n41154 );
or ( n41157 , n41152 , n41155 , n41156 );
xor ( n41158 , n40894 , n40898 );
xor ( n41159 , n41158 , n40903 );
xor ( n41160 , n40924 , n40931 );
xor ( n41161 , n41160 , n40936 );
and ( n41162 , n41159 , n41161 );
xor ( n41163 , n40944 , n40948 );
xor ( n41164 , n41163 , n40964 );
and ( n41165 , n41161 , n41164 );
and ( n41166 , n41159 , n41164 );
or ( n41167 , n41162 , n41165 , n41166 );
xor ( n41168 , n40906 , n40939 );
xor ( n41169 , n41168 , n40967 );
and ( n41170 , n41167 , n41169 );
xor ( n41171 , n40874 , n40876 );
xor ( n41172 , n41171 , n40879 );
and ( n41173 , n41169 , n41172 );
and ( n41174 , n41167 , n41172 );
or ( n41175 , n41170 , n41173 , n41174 );
and ( n41176 , n41157 , n41175 );
xor ( n41177 , n40970 , n41010 );
xor ( n41178 , n41177 , n41013 );
and ( n41179 , n41175 , n41178 );
and ( n41180 , n41157 , n41178 );
or ( n41181 , n41176 , n41179 , n41180 );
xor ( n41182 , n40890 , n41016 );
xor ( n41183 , n41182 , n41019 );
and ( n41184 , n41181 , n41183 );
xor ( n41185 , n40843 , n40845 );
xor ( n41186 , n41185 , n40848 );
and ( n41187 , n41183 , n41186 );
and ( n41188 , n41181 , n41186 );
or ( n41189 , n41184 , n41187 , n41188 );
and ( n41190 , n41036 , n41189 );
buf ( n41191 , n41189 );
or ( n41192 , n41037 , n41190 , n41191 );
not ( n41193 , n40871 );
xor ( n41194 , n41193 , n41030 );
and ( n41195 , n41192 , n41194 );
xor ( n41196 , n41181 , n41183 );
xor ( n41197 , n41196 , n41186 );
buf ( n41198 , n41197 );
and ( n41199 , n40574 , n39335 );
and ( n41200 , n40455 , n39333 );
nor ( n41201 , n41199 , n41200 );
xnor ( n41202 , n41201 , n39300 );
and ( n41203 , n40962 , n39258 );
and ( n41204 , n40698 , n39256 );
nor ( n41205 , n41203 , n41204 );
xnor ( n41206 , n41205 , n39215 );
and ( n41207 , n41202 , n41206 );
and ( n41208 , n40910 , n39194 );
and ( n41209 , n40991 , n39192 );
nor ( n41210 , n41208 , n41209 );
xnor ( n41211 , n41210 , n39199 );
and ( n41212 , n41206 , n41211 );
and ( n41213 , n41202 , n41211 );
or ( n41214 , n41207 , n41212 , n41213 );
and ( n41215 , n39875 , n39665 );
and ( n41216 , n39848 , n39663 );
nor ( n41217 , n41215 , n41216 );
xnor ( n41218 , n41217 , n39608 );
and ( n41219 , n41214 , n41218 );
and ( n41220 , n40069 , n39532 );
and ( n41221 , n39935 , n39530 );
nor ( n41222 , n41220 , n41221 );
xnor ( n41223 , n41222 , n39497 );
and ( n41224 , n41218 , n41223 );
and ( n41225 , n41214 , n41223 );
or ( n41226 , n41219 , n41224 , n41225 );
xor ( n41227 , n40685 , n40976 );
xor ( n41228 , n40976 , n40978 );
not ( n41229 , n41228 );
and ( n41230 , n41227 , n41229 );
and ( n41231 , n39184 , n41230 );
not ( n41232 , n41231 );
xnor ( n41233 , n41232 , n40981 );
and ( n41234 , n39618 , n39984 );
and ( n41235 , n39524 , n39982 );
nor ( n41236 , n41234 , n41235 );
xnor ( n41237 , n41236 , n39865 );
and ( n41238 , n41233 , n41237 );
xor ( n41239 , n41041 , n41045 );
xor ( n41240 , n41239 , n41050 );
and ( n41241 , n41237 , n41240 );
and ( n41242 , n41233 , n41240 );
or ( n41243 , n41238 , n41241 , n41242 );
and ( n41244 , n41226 , n41243 );
and ( n41245 , n39433 , n40168 );
and ( n41246 , n39397 , n40166 );
nor ( n41247 , n41245 , n41246 );
xnor ( n41248 , n41247 , n40059 );
and ( n41249 , n41243 , n41248 );
and ( n41250 , n41226 , n41248 );
or ( n41251 , n41244 , n41249 , n41250 );
xor ( n41252 , n41053 , n41057 );
xor ( n41253 , n41252 , n41062 );
xor ( n41254 , n41069 , n41073 );
xor ( n41255 , n41254 , n41076 );
and ( n41256 , n41253 , n41255 );
xor ( n41257 , n41135 , n41139 );
xor ( n41258 , n41257 , n41142 );
and ( n41259 , n41255 , n41258 );
and ( n41260 , n41253 , n41258 );
or ( n41261 , n41256 , n41259 , n41260 );
and ( n41262 , n41251 , n41261 );
xor ( n41263 , n41065 , n41079 );
xor ( n41264 , n41263 , n41084 );
and ( n41265 , n41261 , n41264 );
and ( n41266 , n41251 , n41264 );
or ( n41267 , n41262 , n41265 , n41266 );
and ( n41268 , n39229 , n40928 );
and ( n41269 , n39220 , n40926 );
nor ( n41270 , n41268 , n41269 );
xnor ( n41271 , n41270 , n40688 );
and ( n41272 , n39397 , n40406 );
and ( n41273 , n39327 , n40404 );
nor ( n41274 , n41272 , n41273 );
xnor ( n41275 , n41274 , n40262 );
and ( n41276 , n41271 , n41275 );
and ( n41277 , n39739 , n39795 );
and ( n41278 , n39657 , n39793 );
nor ( n41279 , n41277 , n41278 );
xnor ( n41280 , n41279 , n39729 );
and ( n41281 , n41275 , n41280 );
and ( n41282 , n41271 , n41280 );
or ( n41283 , n41276 , n41281 , n41282 );
and ( n41284 , n40077 , n39532 );
and ( n41285 , n40069 , n39530 );
nor ( n41286 , n41284 , n41285 );
xnor ( n41287 , n41286 , n39497 );
and ( n41288 , n40280 , n39384 );
and ( n41289 , n40272 , n39382 );
nor ( n41290 , n41288 , n41289 );
xnor ( n41291 , n41290 , n39367 );
and ( n41292 , n41287 , n41291 );
xor ( n41293 , n41093 , n41101 );
xor ( n41294 , n41293 , n41107 );
and ( n41295 , n41291 , n41294 );
and ( n41296 , n41287 , n41294 );
or ( n41297 , n41292 , n41295 , n41296 );
and ( n41298 , n39507 , n40168 );
and ( n41299 , n39433 , n40166 );
nor ( n41300 , n41298 , n41299 );
xnor ( n41301 , n41300 , n40059 );
and ( n41302 , n41297 , n41301 );
xor ( n41303 , n41110 , n41114 );
xor ( n41304 , n41303 , n41116 );
and ( n41305 , n41301 , n41304 );
and ( n41306 , n41297 , n41304 );
or ( n41307 , n41302 , n41305 , n41306 );
and ( n41308 , n41283 , n41307 );
xor ( n41309 , n41119 , n41123 );
xor ( n41310 , n41309 , n41128 );
and ( n41311 , n41307 , n41310 );
and ( n41312 , n41283 , n41310 );
or ( n41313 , n41308 , n41311 , n41312 );
xor ( n41314 , n41131 , n41145 );
xor ( n41315 , n41314 , n41148 );
and ( n41316 , n41313 , n41315 );
xor ( n41317 , n41159 , n41161 );
xor ( n41318 , n41317 , n41164 );
and ( n41319 , n41315 , n41318 );
and ( n41320 , n41313 , n41318 );
or ( n41321 , n41316 , n41319 , n41320 );
and ( n41322 , n41267 , n41321 );
xor ( n41323 , n41087 , n41151 );
xor ( n41324 , n41323 , n41154 );
and ( n41325 , n41321 , n41324 );
and ( n41326 , n41267 , n41324 );
or ( n41327 , n41322 , n41325 , n41326 );
xor ( n41328 , n40882 , n40884 );
xor ( n41329 , n41328 , n40887 );
and ( n41330 , n41327 , n41329 );
xor ( n41331 , n41157 , n41175 );
xor ( n41332 , n41331 , n41178 );
and ( n41333 , n41329 , n41332 );
and ( n41334 , n41327 , n41332 );
or ( n41335 , n41330 , n41333 , n41334 );
and ( n41336 , n41197 , n41335 );
buf ( n41337 , n41335 );
or ( n41338 , n41198 , n41336 , n41337 );
not ( n41339 , n41036 );
xor ( n41340 , n41339 , n41189 );
and ( n41341 , n41338 , n41340 );
xor ( n41342 , n41327 , n41329 );
xor ( n41343 , n41342 , n41332 );
buf ( n41344 , n41343 );
and ( n41345 , n40455 , n39384 );
and ( n41346 , n40280 , n39382 );
nor ( n41347 , n41345 , n41346 );
xnor ( n41348 , n41347 , n39367 );
and ( n41349 , n40698 , n39335 );
and ( n41350 , n40574 , n39333 );
nor ( n41351 , n41349 , n41350 );
xnor ( n41352 , n41351 , n39300 );
and ( n41353 , n41348 , n41352 );
and ( n41354 , n40991 , n39258 );
and ( n41355 , n40962 , n39256 );
nor ( n41356 , n41354 , n41355 );
xnor ( n41357 , n41356 , n39215 );
and ( n41358 , n41352 , n41357 );
and ( n41359 , n41348 , n41357 );
or ( n41360 , n41353 , n41358 , n41359 );
xor ( n41361 , n36181 , n39135 );
buf ( n41362 , n41361 );
buf ( n41363 , n41362 );
buf ( n41364 , n41363 );
and ( n41365 , n41364 , n39186 );
buf ( n41366 , n41365 );
buf ( n41367 , n1183 );
buf ( n41368 , n41367 );
buf ( n41369 , n1184 );
buf ( n41370 , n41369 );
and ( n41371 , n41368 , n41370 );
not ( n41372 , n41371 );
and ( n41373 , n41097 , n41372 );
not ( n41374 , n41373 );
and ( n41375 , n41366 , n41374 );
xor ( n41376 , n36180 , n39136 );
buf ( n41377 , n41376 );
buf ( n41378 , n41377 );
buf ( n41379 , n41378 );
and ( n41380 , n41379 , n39186 );
and ( n41381 , n41374 , n41380 );
and ( n41382 , n41366 , n41380 );
or ( n41383 , n41375 , n41381 , n41382 );
and ( n41384 , n41106 , n39194 );
and ( n41385 , n40910 , n39192 );
nor ( n41386 , n41384 , n41385 );
xnor ( n41387 , n41386 , n39199 );
and ( n41388 , n41383 , n41387 );
not ( n41389 , n41092 );
and ( n41390 , n41387 , n41389 );
and ( n41391 , n41383 , n41389 );
or ( n41392 , n41388 , n41390 , n41391 );
and ( n41393 , n41360 , n41392 );
and ( n41394 , n39935 , n39665 );
and ( n41395 , n39875 , n39663 );
nor ( n41396 , n41394 , n41395 );
xnor ( n41397 , n41396 , n39608 );
and ( n41398 , n41392 , n41397 );
and ( n41399 , n41360 , n41397 );
or ( n41400 , n41393 , n41398 , n41399 );
and ( n41401 , n39524 , n40168 );
and ( n41402 , n39507 , n40166 );
nor ( n41403 , n41401 , n41402 );
xnor ( n41404 , n41403 , n40059 );
and ( n41405 , n39848 , n39795 );
and ( n41406 , n39739 , n39793 );
nor ( n41407 , n41405 , n41406 );
xnor ( n41408 , n41407 , n39729 );
and ( n41409 , n41404 , n41408 );
xor ( n41410 , n41202 , n41206 );
xor ( n41411 , n41410 , n41211 );
and ( n41412 , n41408 , n41411 );
and ( n41413 , n41404 , n41411 );
or ( n41414 , n41409 , n41412 , n41413 );
and ( n41415 , n41400 , n41414 );
and ( n41416 , n39310 , n40666 );
and ( n41417 , n39271 , n40664 );
nor ( n41418 , n41416 , n41417 );
xnor ( n41419 , n41418 , n40445 );
and ( n41420 , n41414 , n41419 );
and ( n41421 , n41400 , n41419 );
or ( n41422 , n41415 , n41420 , n41421 );
and ( n41423 , n39271 , n40928 );
and ( n41424 , n39229 , n40926 );
nor ( n41425 , n41423 , n41424 );
xnor ( n41426 , n41425 , n40688 );
and ( n41427 , n39433 , n40406 );
and ( n41428 , n39397 , n40404 );
nor ( n41429 , n41427 , n41428 );
xnor ( n41430 , n41429 , n40262 );
and ( n41431 , n41426 , n41430 );
xor ( n41432 , n41287 , n41291 );
xor ( n41433 , n41432 , n41294 );
and ( n41434 , n41430 , n41433 );
and ( n41435 , n41426 , n41433 );
or ( n41436 , n41431 , n41434 , n41435 );
xor ( n41437 , n41214 , n41218 );
xor ( n41438 , n41437 , n41223 );
and ( n41439 , n41436 , n41438 );
xor ( n41440 , n41233 , n41237 );
xor ( n41441 , n41440 , n41240 );
and ( n41442 , n41438 , n41441 );
and ( n41443 , n41436 , n41441 );
or ( n41444 , n41439 , n41442 , n41443 );
and ( n41445 , n41422 , n41444 );
xor ( n41446 , n41226 , n41243 );
xor ( n41447 , n41446 , n41248 );
and ( n41448 , n41444 , n41447 );
and ( n41449 , n41422 , n41447 );
or ( n41450 , n41445 , n41448 , n41449 );
and ( n41451 , n39220 , n41230 );
and ( n41452 , n39184 , n41228 );
nor ( n41453 , n41451 , n41452 );
xnor ( n41454 , n41453 , n40981 );
and ( n41455 , n39327 , n40666 );
and ( n41456 , n39310 , n40664 );
nor ( n41457 , n41455 , n41456 );
xnor ( n41458 , n41457 , n40445 );
and ( n41459 , n41454 , n41458 );
and ( n41460 , n39657 , n39984 );
and ( n41461 , n39618 , n39982 );
nor ( n41462 , n41460 , n41461 );
xnor ( n41463 , n41462 , n39865 );
and ( n41464 , n41458 , n41463 );
and ( n41465 , n41454 , n41463 );
or ( n41466 , n41459 , n41464 , n41465 );
xor ( n41467 , n41271 , n41275 );
xor ( n41468 , n41467 , n41280 );
and ( n41469 , n41466 , n41468 );
xor ( n41470 , n41297 , n41301 );
xor ( n41471 , n41470 , n41304 );
and ( n41472 , n41468 , n41471 );
and ( n41473 , n41466 , n41471 );
or ( n41474 , n41469 , n41472 , n41473 );
xor ( n41475 , n41283 , n41307 );
xor ( n41476 , n41475 , n41310 );
and ( n41477 , n41474 , n41476 );
xor ( n41478 , n41253 , n41255 );
xor ( n41479 , n41478 , n41258 );
and ( n41480 , n41476 , n41479 );
and ( n41481 , n41474 , n41479 );
or ( n41482 , n41477 , n41480 , n41481 );
and ( n41483 , n41450 , n41482 );
xor ( n41484 , n41251 , n41261 );
xor ( n41485 , n41484 , n41264 );
and ( n41486 , n41482 , n41485 );
and ( n41487 , n41450 , n41485 );
or ( n41488 , n41483 , n41486 , n41487 );
xor ( n41489 , n41167 , n41169 );
xor ( n41490 , n41489 , n41172 );
and ( n41491 , n41488 , n41490 );
xor ( n41492 , n41267 , n41321 );
xor ( n41493 , n41492 , n41324 );
and ( n41494 , n41490 , n41493 );
and ( n41495 , n41488 , n41493 );
or ( n41496 , n41491 , n41494 , n41495 );
and ( n41497 , n41343 , n41496 );
buf ( n41498 , n41496 );
or ( n41499 , n41344 , n41497 , n41498 );
not ( n41500 , n41197 );
xor ( n41501 , n41500 , n41335 );
and ( n41502 , n41499 , n41501 );
and ( n41503 , n39229 , n41230 );
and ( n41504 , n39220 , n41228 );
nor ( n41505 , n41503 , n41504 );
xnor ( n41506 , n41505 , n40981 );
and ( n41507 , n39397 , n40666 );
and ( n41508 , n39327 , n40664 );
nor ( n41509 , n41507 , n41508 );
xnor ( n41510 , n41509 , n40445 );
and ( n41511 , n41506 , n41510 );
and ( n41512 , n39739 , n39984 );
and ( n41513 , n39657 , n39982 );
nor ( n41514 , n41512 , n41513 );
xnor ( n41515 , n41514 , n39865 );
and ( n41516 , n41510 , n41515 );
and ( n41517 , n41506 , n41515 );
or ( n41518 , n41511 , n41516 , n41517 );
xor ( n41519 , n40978 , n41095 );
xor ( n41520 , n41095 , n41097 );
not ( n41521 , n41520 );
and ( n41522 , n41519 , n41521 );
and ( n41523 , n39184 , n41522 );
not ( n41524 , n41523 );
xnor ( n41525 , n41524 , n41100 );
and ( n41526 , n39618 , n40168 );
and ( n41527 , n39524 , n40166 );
nor ( n41528 , n41526 , n41527 );
xnor ( n41529 , n41528 , n40059 );
and ( n41530 , n41525 , n41529 );
xor ( n41531 , n41348 , n41352 );
xor ( n41532 , n41531 , n41357 );
and ( n41533 , n41529 , n41532 );
and ( n41534 , n41525 , n41532 );
or ( n41535 , n41530 , n41533 , n41534 );
and ( n41536 , n41518 , n41535 );
xor ( n41537 , n41404 , n41408 );
xor ( n41538 , n41537 , n41411 );
and ( n41539 , n41535 , n41538 );
and ( n41540 , n41518 , n41538 );
or ( n41541 , n41536 , n41539 , n41540 );
buf ( n41542 , n41541 );
and ( n41543 , n40069 , n39665 );
and ( n41544 , n39935 , n39663 );
nor ( n41545 , n41543 , n41544 );
xnor ( n41546 , n41545 , n39608 );
buf ( n41547 , n41546 );
buf ( n41548 , n41547 );
and ( n41549 , n40962 , n39335 );
and ( n41550 , n40698 , n39333 );
nor ( n41551 , n41549 , n41550 );
xnor ( n41552 , n41551 , n39300 );
and ( n41553 , n40910 , n39258 );
and ( n41554 , n40991 , n39256 );
nor ( n41555 , n41553 , n41554 );
xnor ( n41556 , n41555 , n39215 );
and ( n41557 , n41552 , n41556 );
and ( n41558 , n41091 , n39194 );
and ( n41559 , n41106 , n39192 );
nor ( n41560 , n41558 , n41559 );
xnor ( n41561 , n41560 , n39199 );
and ( n41562 , n41556 , n41561 );
and ( n41563 , n41552 , n41561 );
or ( n41564 , n41557 , n41562 , n41563 );
not ( n41565 , n41564 );
and ( n41566 , n40272 , n39532 );
and ( n41567 , n40077 , n39530 );
nor ( n41568 , n41566 , n41567 );
xnor ( n41569 , n41568 , n39497 );
and ( n41570 , n41565 , n41569 );
and ( n41571 , n41547 , n41570 );
buf ( n41572 , n41570 );
or ( n41573 , n41548 , n41571 , n41572 );
and ( n41574 , n41541 , n41573 );
buf ( n41575 , n41573 );
or ( n41576 , n41542 , n41574 , n41575 );
buf ( n41577 , n41576 );
buf ( n41578 , n41564 );
not ( n41579 , n41546 );
xor ( n41580 , n41565 , n41569 );
and ( n41581 , n41579 , n41580 );
and ( n41582 , n41578 , n41581 );
not ( n41583 , n41547 );
xor ( n41584 , n41583 , n41570 );
and ( n41585 , n41581 , n41584 );
and ( n41586 , n41578 , n41584 );
or ( n41587 , n41582 , n41585 , n41586 );
not ( n41588 , n41541 );
xor ( n41589 , n41588 , n41573 );
and ( n41590 , n41587 , n41589 );
xor ( n41591 , n41400 , n41414 );
xor ( n41592 , n41591 , n41419 );
and ( n41593 , n41589 , n41592 );
and ( n41594 , n41587 , n41592 );
or ( n41595 , n41590 , n41593 , n41594 );
and ( n41596 , n41576 , n41595 );
buf ( n41597 , n41595 );
or ( n41598 , n41577 , n41596 , n41597 );
buf ( n41599 , n41598 );
xor ( n41600 , n41313 , n41315 );
xor ( n41601 , n41600 , n41318 );
and ( n41602 , n41598 , n41601 );
buf ( n41603 , n41601 );
or ( n41604 , n41599 , n41602 , n41603 );
buf ( n41605 , n41604 );
xor ( n41606 , n41488 , n41490 );
xor ( n41607 , n41606 , n41493 );
and ( n41608 , n41604 , n41607 );
buf ( n41609 , n41607 );
or ( n41610 , n41605 , n41608 , n41609 );
not ( n41611 , n41343 );
xor ( n41612 , n41611 , n41496 );
and ( n41613 , n41610 , n41612 );
xor ( n41614 , n41360 , n41392 );
xor ( n41615 , n41614 , n41397 );
and ( n41616 , n40280 , n39532 );
and ( n41617 , n40272 , n39530 );
nor ( n41618 , n41616 , n41617 );
xnor ( n41619 , n41618 , n39497 );
and ( n41620 , n40574 , n39384 );
and ( n41621 , n40455 , n39382 );
nor ( n41622 , n41620 , n41621 );
xnor ( n41623 , n41622 , n39367 );
and ( n41624 , n41619 , n41623 );
xor ( n41625 , n41366 , n41374 );
xor ( n41626 , n41625 , n41380 );
and ( n41627 , n41623 , n41626 );
and ( n41628 , n41619 , n41626 );
or ( n41629 , n41624 , n41627 , n41628 );
and ( n41630 , n39875 , n39795 );
and ( n41631 , n39848 , n39793 );
nor ( n41632 , n41630 , n41631 );
xnor ( n41633 , n41632 , n39729 );
and ( n41634 , n41629 , n41633 );
xor ( n41635 , n41383 , n41387 );
xor ( n41636 , n41635 , n41389 );
and ( n41637 , n41633 , n41636 );
and ( n41638 , n41629 , n41636 );
or ( n41639 , n41634 , n41637 , n41638 );
and ( n41640 , n41615 , n41639 );
xor ( n41641 , n41578 , n41581 );
xor ( n41642 , n41641 , n41584 );
and ( n41643 , n41639 , n41642 );
and ( n41644 , n41615 , n41642 );
or ( n41645 , n41640 , n41643 , n41644 );
and ( n41646 , n39220 , n41522 );
and ( n41647 , n39184 , n41520 );
nor ( n41648 , n41646 , n41647 );
xnor ( n41649 , n41648 , n41100 );
and ( n41650 , n39327 , n40928 );
and ( n41651 , n39310 , n40926 );
nor ( n41652 , n41650 , n41651 );
xnor ( n41653 , n41652 , n40688 );
and ( n41654 , n41649 , n41653 );
and ( n41655 , n39433 , n40666 );
and ( n41656 , n39397 , n40664 );
nor ( n41657 , n41655 , n41656 );
xnor ( n41658 , n41657 , n40445 );
and ( n41659 , n41653 , n41658 );
and ( n41660 , n41649 , n41658 );
or ( n41661 , n41654 , n41659 , n41660 );
xor ( n41662 , n41525 , n41529 );
xor ( n41663 , n41662 , n41532 );
and ( n41664 , n41661 , n41663 );
xor ( n41665 , n41629 , n41633 );
xor ( n41666 , n41665 , n41636 );
and ( n41667 , n41663 , n41666 );
and ( n41668 , n41661 , n41666 );
or ( n41669 , n41664 , n41667 , n41668 );
xor ( n41670 , n41579 , n41580 );
and ( n41671 , n39848 , n39984 );
and ( n41672 , n39739 , n39982 );
nor ( n41673 , n41671 , n41672 );
xnor ( n41674 , n41673 , n39865 );
and ( n41675 , n39935 , n39795 );
and ( n41676 , n39875 , n39793 );
nor ( n41677 , n41675 , n41676 );
xnor ( n41678 , n41677 , n39729 );
and ( n41679 , n41674 , n41678 );
xor ( n41680 , n41552 , n41556 );
xor ( n41681 , n41680 , n41561 );
and ( n41682 , n41678 , n41681 );
and ( n41683 , n41674 , n41681 );
or ( n41684 , n41679 , n41682 , n41683 );
and ( n41685 , n41670 , n41684 );
and ( n41686 , n39524 , n40406 );
and ( n41687 , n39507 , n40404 );
nor ( n41688 , n41686 , n41687 );
xnor ( n41689 , n41688 , n40262 );
and ( n41690 , n39657 , n40168 );
and ( n41691 , n39618 , n40166 );
nor ( n41692 , n41690 , n41691 );
xnor ( n41693 , n41692 , n40059 );
and ( n41694 , n41689 , n41693 );
xor ( n41695 , n41619 , n41623 );
xor ( n41696 , n41695 , n41626 );
and ( n41697 , n41693 , n41696 );
and ( n41698 , n41689 , n41696 );
or ( n41699 , n41694 , n41697 , n41698 );
and ( n41700 , n41684 , n41699 );
and ( n41701 , n41670 , n41699 );
or ( n41702 , n41685 , n41700 , n41701 );
and ( n41703 , n41669 , n41702 );
xor ( n41704 , n41615 , n41639 );
xor ( n41705 , n41704 , n41642 );
and ( n41706 , n41702 , n41705 );
and ( n41707 , n41669 , n41705 );
or ( n41708 , n41703 , n41706 , n41707 );
and ( n41709 , n41645 , n41708 );
xor ( n41710 , n41587 , n41589 );
xor ( n41711 , n41710 , n41592 );
and ( n41712 , n41708 , n41711 );
and ( n41713 , n41645 , n41711 );
or ( n41714 , n41709 , n41712 , n41713 );
not ( n41715 , n41576 );
xor ( n41716 , n41715 , n41595 );
and ( n41717 , n41714 , n41716 );
xor ( n41718 , n41422 , n41444 );
xor ( n41719 , n41718 , n41447 );
and ( n41720 , n41716 , n41719 );
and ( n41721 , n41714 , n41719 );
or ( n41722 , n41717 , n41720 , n41721 );
xor ( n41723 , n41450 , n41482 );
xor ( n41724 , n41723 , n41485 );
and ( n41725 , n41722 , n41724 );
not ( n41726 , n41370 );
and ( n41727 , n41364 , n39194 );
and ( n41728 , n41379 , n39192 );
nor ( n41729 , n41727 , n41728 );
xnor ( n41730 , n41729 , n39199 );
and ( n41731 , n41726 , n41730 );
xor ( n41732 , n36182 , n39134 );
buf ( n41733 , n41732 );
buf ( n41734 , n41733 );
buf ( n41735 , n41734 );
and ( n41736 , n41735 , n39186 );
and ( n41737 , n41730 , n41736 );
and ( n41738 , n41726 , n41736 );
or ( n41739 , n41731 , n41737 , n41738 );
and ( n41740 , n40455 , n39532 );
and ( n41741 , n40280 , n39530 );
nor ( n41742 , n41740 , n41741 );
xnor ( n41743 , n41742 , n39497 );
and ( n41744 , n41739 , n41743 );
and ( n41745 , n40991 , n39335 );
and ( n41746 , n40962 , n39333 );
nor ( n41747 , n41745 , n41746 );
xnor ( n41748 , n41747 , n39300 );
and ( n41749 , n41743 , n41748 );
and ( n41750 , n41739 , n41748 );
or ( n41751 , n41744 , n41749 , n41750 );
and ( n41752 , n41106 , n39258 );
and ( n41753 , n40910 , n39256 );
nor ( n41754 , n41752 , n41753 );
xnor ( n41755 , n41754 , n39215 );
and ( n41756 , n41379 , n39194 );
and ( n41757 , n41091 , n39192 );
nor ( n41758 , n41756 , n41757 );
xnor ( n41759 , n41758 , n39199 );
and ( n41760 , n41755 , n41759 );
not ( n41761 , n41365 );
and ( n41762 , n41759 , n41761 );
and ( n41763 , n41755 , n41761 );
or ( n41764 , n41760 , n41762 , n41763 );
and ( n41765 , n41751 , n41764 );
and ( n41766 , n40077 , n39665 );
and ( n41767 , n40069 , n39663 );
nor ( n41768 , n41766 , n41767 );
xnor ( n41769 , n41768 , n39608 );
and ( n41770 , n41764 , n41769 );
and ( n41771 , n41751 , n41769 );
or ( n41772 , n41765 , n41770 , n41771 );
and ( n41773 , n39310 , n40928 );
and ( n41774 , n39271 , n40926 );
nor ( n41775 , n41773 , n41774 );
xnor ( n41776 , n41775 , n40688 );
and ( n41777 , n41772 , n41776 );
and ( n41778 , n39507 , n40406 );
and ( n41779 , n39433 , n40404 );
nor ( n41780 , n41778 , n41779 );
xnor ( n41781 , n41780 , n40262 );
and ( n41782 , n41776 , n41781 );
and ( n41783 , n41772 , n41781 );
or ( n41784 , n41777 , n41782 , n41783 );
xor ( n41785 , n41454 , n41458 );
xor ( n41786 , n41785 , n41463 );
and ( n41787 , n41784 , n41786 );
xor ( n41788 , n41426 , n41430 );
xor ( n41789 , n41788 , n41433 );
and ( n41790 , n41786 , n41789 );
and ( n41791 , n41784 , n41789 );
or ( n41792 , n41787 , n41790 , n41791 );
xor ( n41793 , n41436 , n41438 );
xor ( n41794 , n41793 , n41441 );
and ( n41795 , n41792 , n41794 );
xor ( n41796 , n41466 , n41468 );
xor ( n41797 , n41796 , n41471 );
and ( n41798 , n41794 , n41797 );
and ( n41799 , n41792 , n41797 );
or ( n41800 , n41795 , n41798 , n41799 );
xor ( n41801 , n41474 , n41476 );
xor ( n41802 , n41801 , n41479 );
and ( n41803 , n41800 , n41802 );
xor ( n41804 , n41714 , n41716 );
xor ( n41805 , n41804 , n41719 );
and ( n41806 , n41802 , n41805 );
and ( n41807 , n41800 , n41805 );
or ( n41808 , n41803 , n41806 , n41807 );
and ( n41809 , n41724 , n41808 );
and ( n41810 , n41722 , n41808 );
or ( n41811 , n41725 , n41809 , n41810 );
not ( n41812 , n41604 );
xor ( n41813 , n41812 , n41607 );
and ( n41814 , n41811 , n41813 );
not ( n41815 , n41598 );
xor ( n41816 , n41815 , n41601 );
xor ( n41817 , n41722 , n41724 );
xor ( n41818 , n41817 , n41808 );
and ( n41819 , n41816 , n41818 );
xor ( n41820 , n41645 , n41708 );
xor ( n41821 , n41820 , n41711 );
xor ( n41822 , n41792 , n41794 );
xor ( n41823 , n41822 , n41797 );
and ( n41824 , n41821 , n41823 );
xor ( n41825 , n37165 , n39129 );
buf ( n41826 , n41825 );
buf ( n41827 , n41826 );
buf ( n41828 , n41827 );
and ( n41829 , n41828 , n39186 );
buf ( n41830 , n30346 );
not ( n41831 , n41830 );
and ( n41832 , n41829 , n41831 );
buf ( n41833 , n30345 );
not ( n41834 , n41833 );
and ( n41835 , n41832 , n41834 );
and ( n41836 , n41379 , n39258 );
and ( n41837 , n41091 , n39256 );
nor ( n41838 , n41836 , n41837 );
xnor ( n41839 , n41838 , n39215 );
and ( n41840 , n41835 , n41839 );
xor ( n41841 , n36616 , n39132 );
buf ( n41842 , n41841 );
buf ( n41843 , n41842 );
buf ( n41844 , n41843 );
and ( n41845 , n41844 , n39186 );
and ( n41846 , n41839 , n41845 );
and ( n41847 , n41835 , n41845 );
or ( n41848 , n41840 , n41846 , n41847 );
and ( n41849 , n41735 , n39194 );
and ( n41850 , n41364 , n39192 );
nor ( n41851 , n41849 , n41850 );
xnor ( n41852 , n41851 , n39199 );
buf ( n41853 , n41852 );
and ( n41854 , n41848 , n41853 );
and ( n41855 , n41091 , n39258 );
and ( n41856 , n41106 , n39256 );
nor ( n41857 , n41855 , n41856 );
xnor ( n41858 , n41857 , n39215 );
and ( n41859 , n41853 , n41858 );
and ( n41860 , n41848 , n41858 );
or ( n41861 , n41854 , n41859 , n41860 );
and ( n41862 , n40962 , n39384 );
and ( n41863 , n40698 , n39382 );
nor ( n41864 , n41862 , n41863 );
xnor ( n41865 , n41864 , n39367 );
and ( n41866 , n40910 , n39335 );
and ( n41867 , n40991 , n39333 );
nor ( n41868 , n41866 , n41867 );
xnor ( n41869 , n41868 , n39300 );
and ( n41870 , n41865 , n41869 );
xor ( n41871 , n41726 , n41730 );
xor ( n41872 , n41871 , n41736 );
and ( n41873 , n41869 , n41872 );
and ( n41874 , n41865 , n41872 );
or ( n41875 , n41870 , n41873 , n41874 );
and ( n41876 , n41861 , n41875 );
and ( n41877 , n40069 , n39795 );
and ( n41878 , n39935 , n39793 );
nor ( n41879 , n41877 , n41878 );
xnor ( n41880 , n41879 , n39729 );
and ( n41881 , n41875 , n41880 );
and ( n41882 , n41861 , n41880 );
or ( n41883 , n41876 , n41881 , n41882 );
and ( n41884 , n40272 , n39665 );
and ( n41885 , n40077 , n39663 );
nor ( n41886 , n41884 , n41885 );
xnor ( n41887 , n41886 , n39608 );
and ( n41888 , n40698 , n39384 );
and ( n41889 , n40574 , n39382 );
nor ( n41890 , n41888 , n41889 );
xnor ( n41891 , n41890 , n39367 );
and ( n41892 , n41887 , n41891 );
xor ( n41893 , n41755 , n41759 );
xor ( n41894 , n41893 , n41761 );
and ( n41895 , n41891 , n41894 );
and ( n41896 , n41887 , n41894 );
or ( n41897 , n41892 , n41895 , n41896 );
and ( n41898 , n41883 , n41897 );
and ( n41899 , n39271 , n41230 );
and ( n41900 , n39229 , n41228 );
nor ( n41901 , n41899 , n41900 );
xnor ( n41902 , n41901 , n40981 );
and ( n41903 , n41897 , n41902 );
and ( n41904 , n41883 , n41902 );
or ( n41905 , n41898 , n41903 , n41904 );
xor ( n41906 , n41506 , n41510 );
xor ( n41907 , n41906 , n41515 );
and ( n41908 , n41905 , n41907 );
xor ( n41909 , n41772 , n41776 );
xor ( n41910 , n41909 , n41781 );
and ( n41911 , n41907 , n41910 );
and ( n41912 , n41905 , n41910 );
or ( n41913 , n41908 , n41911 , n41912 );
xor ( n41914 , n41518 , n41535 );
xor ( n41915 , n41914 , n41538 );
and ( n41916 , n41913 , n41915 );
xor ( n41917 , n41784 , n41786 );
xor ( n41918 , n41917 , n41789 );
and ( n41919 , n41915 , n41918 );
and ( n41920 , n41913 , n41918 );
or ( n41921 , n41916 , n41919 , n41920 );
and ( n41922 , n41823 , n41921 );
and ( n41923 , n41821 , n41921 );
or ( n41924 , n41824 , n41922 , n41923 );
xor ( n41925 , n41800 , n41802 );
xor ( n41926 , n41925 , n41805 );
and ( n41927 , n41924 , n41926 );
xor ( n41928 , n41670 , n41684 );
xor ( n41929 , n41928 , n41699 );
buf ( n41930 , n41929 );
and ( n41931 , n39229 , n41522 );
and ( n41932 , n39220 , n41520 );
nor ( n41933 , n41931 , n41932 );
xnor ( n41934 , n41933 , n41100 );
and ( n41935 , n39397 , n40928 );
and ( n41936 , n39327 , n40926 );
nor ( n41937 , n41935 , n41936 );
xnor ( n41938 , n41937 , n40688 );
and ( n41939 , n41934 , n41938 );
and ( n41940 , n39507 , n40666 );
and ( n41941 , n39433 , n40664 );
nor ( n41942 , n41940 , n41941 );
xnor ( n41943 , n41942 , n40445 );
and ( n41944 , n41938 , n41943 );
and ( n41945 , n41934 , n41943 );
or ( n41946 , n41939 , n41944 , n41945 );
xor ( n41947 , n41674 , n41678 );
xor ( n41948 , n41947 , n41681 );
and ( n41949 , n41946 , n41948 );
xor ( n41950 , n41689 , n41693 );
xor ( n41951 , n41950 , n41696 );
and ( n41952 , n41948 , n41951 );
and ( n41953 , n41946 , n41951 );
or ( n41954 , n41949 , n41952 , n41953 );
and ( n41955 , n41929 , n41954 );
buf ( n41956 , n41954 );
or ( n41957 , n41930 , n41955 , n41956 );
xor ( n41958 , n41669 , n41702 );
xor ( n41959 , n41958 , n41705 );
and ( n41960 , n41957 , n41959 );
and ( n41961 , n39271 , n41522 );
and ( n41962 , n39229 , n41520 );
nor ( n41963 , n41961 , n41962 );
xnor ( n41964 , n41963 , n41100 );
and ( n41965 , n39327 , n41230 );
and ( n41966 , n39310 , n41228 );
nor ( n41967 , n41965 , n41966 );
xnor ( n41968 , n41967 , n40981 );
and ( n41969 , n41964 , n41968 );
and ( n41970 , n39433 , n40928 );
and ( n41971 , n39397 , n40926 );
nor ( n41972 , n41970 , n41971 );
xnor ( n41973 , n41972 , n40688 );
and ( n41974 , n41968 , n41973 );
and ( n41975 , n41964 , n41973 );
or ( n41976 , n41969 , n41974 , n41975 );
buf ( n41977 , n41976 );
xor ( n41978 , n41097 , n41368 );
xor ( n41979 , n41368 , n41370 );
not ( n41980 , n41979 );
and ( n41981 , n41978 , n41980 );
and ( n41982 , n39220 , n41981 );
and ( n41983 , n39184 , n41979 );
nor ( n41984 , n41982 , n41983 );
xnor ( n41985 , n41984 , n41373 );
and ( n41986 , n39524 , n40666 );
and ( n41987 , n39507 , n40664 );
nor ( n41988 , n41986 , n41987 );
xnor ( n41989 , n41988 , n40445 );
xor ( n41990 , n41985 , n41989 );
and ( n41991 , n39657 , n40406 );
and ( n41992 , n39618 , n40404 );
nor ( n41993 , n41991 , n41992 );
xnor ( n41994 , n41993 , n40262 );
xor ( n41995 , n41990 , n41994 );
buf ( n41996 , n41995 );
and ( n41997 , n39229 , n41981 );
and ( n41998 , n39220 , n41979 );
nor ( n41999 , n41997 , n41998 );
xnor ( n42000 , n41999 , n41373 );
and ( n42001 , n39397 , n41230 );
and ( n42002 , n39327 , n41228 );
nor ( n42003 , n42001 , n42002 );
xnor ( n42004 , n42003 , n40981 );
and ( n42005 , n42000 , n42004 );
and ( n42006 , n39507 , n40928 );
and ( n42007 , n39433 , n40926 );
nor ( n42008 , n42006 , n42007 );
xnor ( n42009 , n42008 , n40688 );
and ( n42010 , n42004 , n42009 );
and ( n42011 , n42000 , n42009 );
or ( n42012 , n42005 , n42010 , n42011 );
and ( n42013 , n41995 , n42012 );
buf ( n42014 , n42012 );
or ( n42015 , n41996 , n42013 , n42014 );
and ( n42016 , n41976 , n42015 );
buf ( n42017 , n42015 );
or ( n42018 , n41977 , n42016 , n42017 );
buf ( n42019 , n42018 );
and ( n42020 , n39310 , n41522 );
and ( n42021 , n39271 , n41520 );
nor ( n42022 , n42020 , n42021 );
xnor ( n42023 , n42022 , n41100 );
and ( n42024 , n40272 , n39795 );
and ( n42025 , n40077 , n39793 );
nor ( n42026 , n42024 , n42025 );
xnor ( n42027 , n42026 , n39729 );
and ( n42028 , n42023 , n42027 );
and ( n42029 , n40698 , n39532 );
and ( n42030 , n40574 , n39530 );
nor ( n42031 , n42029 , n42030 );
xnor ( n42032 , n42031 , n39497 );
and ( n42033 , n42027 , n42032 );
and ( n42034 , n42023 , n42032 );
or ( n42035 , n42028 , n42033 , n42034 );
xor ( n42036 , n41964 , n41968 );
xor ( n42037 , n42036 , n41973 );
and ( n42038 , n42035 , n42037 );
xor ( n42039 , n42000 , n42004 );
xor ( n42040 , n42039 , n42009 );
buf ( n42041 , n42040 );
and ( n42042 , n41091 , n39335 );
and ( n42043 , n41106 , n39333 );
nor ( n42044 , n42042 , n42043 );
xnor ( n42045 , n42044 , n39300 );
and ( n42046 , n41364 , n39258 );
and ( n42047 , n41379 , n39256 );
nor ( n42048 , n42046 , n42047 );
xnor ( n42049 , n42048 , n39215 );
and ( n42050 , n42045 , n42049 );
and ( n42051 , n42040 , n42050 );
buf ( n42052 , n42050 );
or ( n42053 , n42041 , n42051 , n42052 );
and ( n42054 , n42037 , n42053 );
and ( n42055 , n42035 , n42053 );
or ( n42056 , n42038 , n42054 , n42055 );
not ( n42057 , n41976 );
xor ( n42058 , n42057 , n42015 );
and ( n42059 , n42056 , n42058 );
not ( n42060 , n41995 );
xor ( n42061 , n42060 , n42012 );
and ( n42062 , n39848 , n40168 );
and ( n42063 , n39739 , n40166 );
nor ( n42064 , n42062 , n42063 );
xnor ( n42065 , n42064 , n40059 );
and ( n42066 , n39935 , n39984 );
and ( n42067 , n39875 , n39982 );
nor ( n42068 , n42066 , n42067 );
xnor ( n42069 , n42068 , n39865 );
xor ( n42070 , n42065 , n42069 );
xor ( n42071 , n41865 , n41869 );
xor ( n42072 , n42071 , n41872 );
xor ( n42073 , n42070 , n42072 );
and ( n42074 , n42061 , n42073 );
buf ( n42075 , n1185 );
buf ( n42076 , n42075 );
xor ( n42077 , n41370 , n42076 );
not ( n42078 , n42076 );
and ( n42079 , n42077 , n42078 );
and ( n42080 , n39220 , n42079 );
and ( n42081 , n39184 , n42076 );
nor ( n42082 , n42080 , n42081 );
xnor ( n42083 , n42082 , n41370 );
and ( n42084 , n39657 , n40666 );
and ( n42085 , n39618 , n40664 );
nor ( n42086 , n42084 , n42085 );
xnor ( n42087 , n42086 , n40445 );
and ( n42088 , n42083 , n42087 );
and ( n42089 , n39935 , n40168 );
and ( n42090 , n39875 , n40166 );
nor ( n42091 , n42089 , n42090 );
xnor ( n42092 , n42091 , n40059 );
and ( n42093 , n42087 , n42092 );
and ( n42094 , n42083 , n42092 );
or ( n42095 , n42088 , n42093 , n42094 );
xor ( n42096 , n42023 , n42027 );
xor ( n42097 , n42096 , n42032 );
and ( n42098 , n42095 , n42097 );
and ( n42099 , n39524 , n40928 );
and ( n42100 , n39507 , n40926 );
nor ( n42101 , n42099 , n42100 );
xnor ( n42102 , n42101 , n40688 );
and ( n42103 , n39848 , n40406 );
and ( n42104 , n39739 , n40404 );
nor ( n42105 , n42103 , n42104 );
xnor ( n42106 , n42105 , n40262 );
and ( n42107 , n42102 , n42106 );
and ( n42108 , n40280 , n39795 );
and ( n42109 , n40272 , n39793 );
nor ( n42110 , n42108 , n42109 );
xnor ( n42111 , n42110 , n39729 );
and ( n42112 , n40574 , n39665 );
and ( n42113 , n40455 , n39663 );
nor ( n42114 , n42112 , n42113 );
xnor ( n42115 , n42114 , n39608 );
xor ( n42116 , n42111 , n42115 );
and ( n42117 , n40962 , n39532 );
and ( n42118 , n40698 , n39530 );
nor ( n42119 , n42117 , n42118 );
xnor ( n42120 , n42119 , n39497 );
xor ( n42121 , n42116 , n42120 );
and ( n42122 , n42106 , n42121 );
and ( n42123 , n42102 , n42121 );
or ( n42124 , n42107 , n42122 , n42123 );
and ( n42125 , n42097 , n42124 );
and ( n42126 , n42095 , n42124 );
or ( n42127 , n42098 , n42125 , n42126 );
and ( n42128 , n42073 , n42127 );
and ( n42129 , n42061 , n42127 );
or ( n42130 , n42074 , n42128 , n42129 );
and ( n42131 , n42058 , n42130 );
and ( n42132 , n42056 , n42130 );
or ( n42133 , n42059 , n42131 , n42132 );
and ( n42134 , n42018 , n42133 );
buf ( n42135 , n42133 );
or ( n42136 , n42019 , n42134 , n42135 );
not ( n42137 , n41929 );
xor ( n42138 , n42137 , n41954 );
and ( n42139 , n42136 , n42138 );
xor ( n42140 , n41832 , n41834 );
and ( n42141 , n41844 , n39194 );
and ( n42142 , n41735 , n39192 );
nor ( n42143 , n42141 , n42142 );
xnor ( n42144 , n42143 , n39199 );
and ( n42145 , n42140 , n42144 );
xor ( n42146 , n36618 , n39131 );
buf ( n42147 , n42146 );
buf ( n42148 , n42147 );
buf ( n42149 , n42148 );
and ( n42150 , n42149 , n39186 );
and ( n42151 , n42144 , n42150 );
and ( n42152 , n42140 , n42150 );
or ( n42153 , n42145 , n42151 , n42152 );
and ( n42154 , n41106 , n39335 );
and ( n42155 , n40910 , n39333 );
nor ( n42156 , n42154 , n42155 );
xnor ( n42157 , n42156 , n39300 );
and ( n42158 , n42153 , n42157 );
not ( n42159 , n41852 );
and ( n42160 , n42157 , n42159 );
and ( n42161 , n42153 , n42159 );
or ( n42162 , n42158 , n42160 , n42161 );
and ( n42163 , n40280 , n39665 );
and ( n42164 , n40272 , n39663 );
nor ( n42165 , n42163 , n42164 );
xnor ( n42166 , n42165 , n39608 );
and ( n42167 , n42162 , n42166 );
and ( n42168 , n40574 , n39532 );
and ( n42169 , n40455 , n39530 );
nor ( n42170 , n42168 , n42169 );
xnor ( n42171 , n42170 , n39497 );
and ( n42172 , n42166 , n42171 );
and ( n42173 , n42162 , n42171 );
or ( n42174 , n42167 , n42172 , n42173 );
and ( n42175 , n39184 , n41981 );
not ( n42176 , n42175 );
xnor ( n42177 , n42176 , n41373 );
and ( n42178 , n42174 , n42177 );
and ( n42179 , n39875 , n39984 );
and ( n42180 , n39848 , n39982 );
nor ( n42181 , n42179 , n42180 );
xnor ( n42182 , n42181 , n39865 );
and ( n42183 , n42177 , n42182 );
and ( n42184 , n42174 , n42182 );
or ( n42185 , n42178 , n42183 , n42184 );
and ( n42186 , n39618 , n40406 );
and ( n42187 , n39524 , n40404 );
nor ( n42188 , n42186 , n42187 );
xnor ( n42189 , n42188 , n40262 );
and ( n42190 , n39739 , n40168 );
and ( n42191 , n39657 , n40166 );
nor ( n42192 , n42190 , n42191 );
xnor ( n42193 , n42192 , n40059 );
and ( n42194 , n42189 , n42193 );
xor ( n42195 , n41739 , n41743 );
xor ( n42196 , n42195 , n41748 );
and ( n42197 , n42193 , n42196 );
and ( n42198 , n42189 , n42196 );
or ( n42199 , n42194 , n42197 , n42198 );
and ( n42200 , n42185 , n42199 );
xor ( n42201 , n41751 , n41764 );
xor ( n42202 , n42201 , n41769 );
and ( n42203 , n42199 , n42202 );
and ( n42204 , n42185 , n42202 );
or ( n42205 , n42200 , n42203 , n42204 );
and ( n42206 , n42138 , n42205 );
and ( n42207 , n42136 , n42205 );
or ( n42208 , n42139 , n42206 , n42207 );
and ( n42209 , n41959 , n42208 );
and ( n42210 , n41957 , n42208 );
or ( n42211 , n41960 , n42209 , n42210 );
xor ( n42212 , n41913 , n41915 );
xor ( n42213 , n42212 , n41918 );
and ( n42214 , n40455 , n39665 );
and ( n42215 , n40280 , n39663 );
nor ( n42216 , n42214 , n42215 );
xnor ( n42217 , n42216 , n39608 );
and ( n42218 , n40991 , n39384 );
and ( n42219 , n40962 , n39382 );
nor ( n42220 , n42218 , n42219 );
xnor ( n42221 , n42220 , n39367 );
and ( n42222 , n42217 , n42221 );
xor ( n42223 , n41835 , n41839 );
xor ( n42224 , n42223 , n41845 );
and ( n42225 , n42221 , n42224 );
and ( n42226 , n42217 , n42224 );
or ( n42227 , n42222 , n42225 , n42226 );
and ( n42228 , n40077 , n39795 );
and ( n42229 , n40069 , n39793 );
nor ( n42230 , n42228 , n42229 );
xnor ( n42231 , n42230 , n39729 );
and ( n42232 , n42227 , n42231 );
xor ( n42233 , n41848 , n41853 );
xor ( n42234 , n42233 , n41858 );
and ( n42235 , n42231 , n42234 );
and ( n42236 , n42227 , n42234 );
or ( n42237 , n42232 , n42235 , n42236 );
and ( n42238 , n39310 , n41230 );
and ( n42239 , n39271 , n41228 );
nor ( n42240 , n42238 , n42239 );
xnor ( n42241 , n42240 , n40981 );
and ( n42242 , n42237 , n42241 );
xor ( n42243 , n41887 , n41891 );
xor ( n42244 , n42243 , n41894 );
and ( n42245 , n42241 , n42244 );
and ( n42246 , n42237 , n42244 );
or ( n42247 , n42242 , n42245 , n42246 );
xor ( n42248 , n41649 , n41653 );
xor ( n42249 , n42248 , n41658 );
and ( n42250 , n42247 , n42249 );
xor ( n42251 , n41883 , n41897 );
xor ( n42252 , n42251 , n41902 );
and ( n42253 , n42249 , n42252 );
and ( n42254 , n42247 , n42252 );
or ( n42255 , n42250 , n42253 , n42254 );
xor ( n42256 , n41905 , n41907 );
xor ( n42257 , n42256 , n41910 );
and ( n42258 , n42255 , n42257 );
xor ( n42259 , n41661 , n41663 );
xor ( n42260 , n42259 , n41666 );
and ( n42261 , n42257 , n42260 );
and ( n42262 , n42255 , n42260 );
or ( n42263 , n42258 , n42261 , n42262 );
and ( n42264 , n42213 , n42263 );
and ( n42265 , n41985 , n41989 );
and ( n42266 , n41989 , n41994 );
and ( n42267 , n41985 , n41994 );
or ( n42268 , n42265 , n42266 , n42267 );
xor ( n42269 , n42174 , n42177 );
xor ( n42270 , n42269 , n42182 );
and ( n42271 , n42268 , n42270 );
xor ( n42272 , n42189 , n42193 );
xor ( n42273 , n42272 , n42196 );
and ( n42274 , n42270 , n42273 );
and ( n42275 , n42268 , n42273 );
or ( n42276 , n42271 , n42274 , n42275 );
not ( n42277 , n42276 );
xor ( n42278 , n42185 , n42199 );
xor ( n42279 , n42278 , n42202 );
and ( n42280 , n42277 , n42279 );
buf ( n42281 , n42276 );
and ( n42282 , n42280 , n42281 );
not ( n42283 , n42018 );
xor ( n42284 , n42283 , n42133 );
and ( n42285 , n42065 , n42069 );
and ( n42286 , n42069 , n42072 );
and ( n42287 , n42065 , n42072 );
or ( n42288 , n42285 , n42286 , n42287 );
xor ( n42289 , n41861 , n41875 );
xor ( n42290 , n42289 , n41880 );
or ( n42291 , n42288 , n42290 );
and ( n42292 , n42284 , n42291 );
and ( n42293 , n40077 , n39984 );
and ( n42294 , n40069 , n39982 );
nor ( n42295 , n42293 , n42294 );
xnor ( n42296 , n42295 , n39865 );
and ( n42297 , n40910 , n39384 );
and ( n42298 , n40991 , n39382 );
nor ( n42299 , n42297 , n42298 );
xnor ( n42300 , n42299 , n39367 );
and ( n42301 , n42296 , n42300 );
and ( n42302 , n39271 , n41981 );
and ( n42303 , n39229 , n41979 );
nor ( n42304 , n42302 , n42303 );
xnor ( n42305 , n42304 , n41373 );
and ( n42306 , n39327 , n41522 );
and ( n42307 , n39310 , n41520 );
nor ( n42308 , n42306 , n42307 );
xnor ( n42309 , n42308 , n41100 );
xor ( n42310 , n42305 , n42309 );
and ( n42311 , n39433 , n41230 );
and ( n42312 , n39397 , n41228 );
nor ( n42313 , n42311 , n42312 );
xnor ( n42314 , n42313 , n40981 );
xor ( n42315 , n42310 , n42314 );
and ( n42316 , n42300 , n42315 );
and ( n42317 , n42296 , n42315 );
or ( n42318 , n42301 , n42316 , n42317 );
xor ( n42319 , n42045 , n42049 );
and ( n42320 , n39229 , n42079 );
and ( n42321 , n39220 , n42076 );
nor ( n42322 , n42320 , n42321 );
xnor ( n42323 , n42322 , n41370 );
and ( n42324 , n39618 , n40928 );
and ( n42325 , n39524 , n40926 );
nor ( n42326 , n42324 , n42325 );
xnor ( n42327 , n42326 , n40688 );
and ( n42328 , n42323 , n42327 );
and ( n42329 , n39739 , n40666 );
and ( n42330 , n39657 , n40664 );
nor ( n42331 , n42329 , n42330 );
xnor ( n42332 , n42331 , n40445 );
and ( n42333 , n42327 , n42332 );
and ( n42334 , n42323 , n42332 );
or ( n42335 , n42328 , n42333 , n42334 );
and ( n42336 , n42319 , n42335 );
and ( n42337 , n40455 , n39795 );
and ( n42338 , n40280 , n39793 );
nor ( n42339 , n42337 , n42338 );
xnor ( n42340 , n42339 , n39729 );
and ( n42341 , n40698 , n39665 );
and ( n42342 , n40574 , n39663 );
nor ( n42343 , n42341 , n42342 );
xnor ( n42344 , n42343 , n39608 );
and ( n42345 , n42340 , n42344 );
and ( n42346 , n40991 , n39532 );
and ( n42347 , n40962 , n39530 );
nor ( n42348 , n42346 , n42347 );
xnor ( n42349 , n42348 , n39497 );
and ( n42350 , n42344 , n42349 );
and ( n42351 , n42340 , n42349 );
or ( n42352 , n42345 , n42350 , n42351 );
and ( n42353 , n42335 , n42352 );
and ( n42354 , n42319 , n42352 );
or ( n42355 , n42336 , n42353 , n42354 );
and ( n42356 , n42318 , n42355 );
and ( n42357 , n39310 , n41981 );
and ( n42358 , n39271 , n41979 );
nor ( n42359 , n42357 , n42358 );
xnor ( n42360 , n42359 , n41373 );
and ( n42361 , n39397 , n41522 );
and ( n42362 , n39327 , n41520 );
nor ( n42363 , n42361 , n42362 );
xnor ( n42364 , n42363 , n41100 );
and ( n42365 , n42360 , n42364 );
and ( n42366 , n39507 , n41230 );
and ( n42367 , n39433 , n41228 );
nor ( n42368 , n42366 , n42367 );
xnor ( n42369 , n42368 , n40981 );
and ( n42370 , n42364 , n42369 );
and ( n42371 , n42360 , n42369 );
or ( n42372 , n42365 , n42370 , n42371 );
and ( n42373 , n41379 , n39335 );
and ( n42374 , n41091 , n39333 );
nor ( n42375 , n42373 , n42374 );
xnor ( n42376 , n42375 , n39300 );
and ( n42377 , n42149 , n39194 );
and ( n42378 , n41844 , n39192 );
nor ( n42379 , n42377 , n42378 );
xnor ( n42380 , n42379 , n39199 );
or ( n42381 , n42376 , n42380 );
and ( n42382 , n42372 , n42381 );
and ( n42383 , n39875 , n40406 );
and ( n42384 , n39848 , n40404 );
nor ( n42385 , n42383 , n42384 );
xnor ( n42386 , n42385 , n40262 );
and ( n42387 , n40069 , n40168 );
and ( n42388 , n39935 , n40166 );
nor ( n42389 , n42387 , n42388 );
xnor ( n42390 , n42389 , n40059 );
and ( n42391 , n42386 , n42390 );
and ( n42392 , n40272 , n39984 );
and ( n42393 , n40077 , n39982 );
nor ( n42394 , n42392 , n42393 );
xnor ( n42395 , n42394 , n39865 );
and ( n42396 , n42390 , n42395 );
and ( n42397 , n42386 , n42395 );
or ( n42398 , n42391 , n42396 , n42397 );
and ( n42399 , n42381 , n42398 );
and ( n42400 , n42372 , n42398 );
or ( n42401 , n42382 , n42399 , n42400 );
and ( n42402 , n42355 , n42401 );
and ( n42403 , n42318 , n42401 );
or ( n42404 , n42356 , n42402 , n42403 );
xor ( n42405 , n42035 , n42037 );
xor ( n42406 , n42405 , n42053 );
and ( n42407 , n42404 , n42406 );
not ( n42408 , n42040 );
xor ( n42409 , n42408 , n42050 );
xor ( n42410 , n42083 , n42087 );
xor ( n42411 , n42410 , n42092 );
xor ( n42412 , n42102 , n42106 );
xor ( n42413 , n42412 , n42121 );
and ( n42414 , n42411 , n42413 );
and ( n42415 , n41106 , n39384 );
and ( n42416 , n40910 , n39382 );
nor ( n42417 , n42415 , n42416 );
xnor ( n42418 , n42417 , n39367 );
and ( n42419 , n41735 , n39258 );
and ( n42420 , n41364 , n39256 );
nor ( n42421 , n42419 , n42420 );
xnor ( n42422 , n42421 , n39215 );
and ( n42423 , n42418 , n42422 );
xor ( n42424 , n42323 , n42327 );
xor ( n42425 , n42424 , n42332 );
and ( n42426 , n42422 , n42425 );
and ( n42427 , n42418 , n42425 );
or ( n42428 , n42423 , n42426 , n42427 );
and ( n42429 , n42413 , n42428 );
and ( n42430 , n42411 , n42428 );
or ( n42431 , n42414 , n42429 , n42430 );
and ( n42432 , n42409 , n42431 );
xor ( n42433 , n42340 , n42344 );
xor ( n42434 , n42433 , n42349 );
xor ( n42435 , n42360 , n42364 );
xor ( n42436 , n42435 , n42369 );
and ( n42437 , n42434 , n42436 );
xnor ( n42438 , n42376 , n42380 );
and ( n42439 , n42436 , n42438 );
and ( n42440 , n42434 , n42438 );
or ( n42441 , n42437 , n42439 , n42440 );
xor ( n42442 , n41829 , n41831 );
and ( n42443 , n40574 , n39795 );
and ( n42444 , n40455 , n39793 );
nor ( n42445 , n42443 , n42444 );
xnor ( n42446 , n42445 , n39729 );
and ( n42447 , n40962 , n39665 );
and ( n42448 , n40698 , n39663 );
nor ( n42449 , n42447 , n42448 );
xnor ( n42450 , n42449 , n39608 );
and ( n42451 , n42446 , n42450 );
and ( n42452 , n40910 , n39532 );
and ( n42453 , n40991 , n39530 );
nor ( n42454 , n42452 , n42453 );
xnor ( n42455 , n42454 , n39497 );
and ( n42456 , n42450 , n42455 );
and ( n42457 , n42446 , n42455 );
or ( n42458 , n42451 , n42456 , n42457 );
and ( n42459 , n42442 , n42458 );
and ( n42460 , n39271 , n42079 );
and ( n42461 , n39229 , n42076 );
nor ( n42462 , n42460 , n42461 );
xnor ( n42463 , n42462 , n41370 );
and ( n42464 , n39327 , n41981 );
and ( n42465 , n39310 , n41979 );
nor ( n42466 , n42464 , n42465 );
xnor ( n42467 , n42466 , n41373 );
and ( n42468 , n42463 , n42467 );
and ( n42469 , n39433 , n41522 );
and ( n42470 , n39397 , n41520 );
nor ( n42471 , n42469 , n42470 );
xnor ( n42472 , n42471 , n41100 );
and ( n42473 , n42467 , n42472 );
and ( n42474 , n42463 , n42472 );
or ( n42475 , n42468 , n42473 , n42474 );
and ( n42476 , n42458 , n42475 );
and ( n42477 , n42442 , n42475 );
or ( n42478 , n42459 , n42476 , n42477 );
and ( n42479 , n42441 , n42478 );
and ( n42480 , n39524 , n41230 );
and ( n42481 , n39507 , n41228 );
nor ( n42482 , n42480 , n42481 );
xnor ( n42483 , n42482 , n40981 );
and ( n42484 , n39935 , n40406 );
and ( n42485 , n39875 , n40404 );
nor ( n42486 , n42484 , n42485 );
xnor ( n42487 , n42486 , n40262 );
and ( n42488 , n42483 , n42487 );
and ( n42489 , n40077 , n40168 );
and ( n42490 , n40069 , n40166 );
nor ( n42491 , n42489 , n42490 );
xnor ( n42492 , n42491 , n40059 );
and ( n42493 , n42487 , n42492 );
and ( n42494 , n42483 , n42492 );
or ( n42495 , n42488 , n42493 , n42494 );
and ( n42496 , n40280 , n39984 );
and ( n42497 , n40272 , n39982 );
nor ( n42498 , n42496 , n42497 );
xnor ( n42499 , n42498 , n39865 );
and ( n42500 , n41091 , n39384 );
and ( n42501 , n41106 , n39382 );
nor ( n42502 , n42500 , n42501 );
xnor ( n42503 , n42502 , n39367 );
and ( n42504 , n42499 , n42503 );
and ( n42505 , n41364 , n39335 );
and ( n42506 , n41379 , n39333 );
nor ( n42507 , n42505 , n42506 );
xnor ( n42508 , n42507 , n39300 );
and ( n42509 , n42503 , n42508 );
and ( n42510 , n42499 , n42508 );
or ( n42511 , n42504 , n42509 , n42510 );
and ( n42512 , n42495 , n42511 );
and ( n42513 , n41844 , n39258 );
and ( n42514 , n41735 , n39256 );
nor ( n42515 , n42513 , n42514 );
xnor ( n42516 , n42515 , n39215 );
and ( n42517 , n41828 , n39194 );
and ( n42518 , n42149 , n39192 );
nor ( n42519 , n42517 , n42518 );
xnor ( n42520 , n42519 , n39199 );
and ( n42521 , n42516 , n42520 );
xor ( n42522 , n37166 , n39128 );
buf ( n42523 , n42522 );
buf ( n42524 , n42523 );
buf ( n42525 , n42524 );
and ( n42526 , n42525 , n39186 );
and ( n42527 , n42520 , n42526 );
and ( n42528 , n42516 , n42526 );
or ( n42529 , n42521 , n42527 , n42528 );
and ( n42530 , n42511 , n42529 );
and ( n42531 , n42495 , n42529 );
or ( n42532 , n42512 , n42530 , n42531 );
and ( n42533 , n42478 , n42532 );
and ( n42534 , n42441 , n42532 );
or ( n42535 , n42479 , n42533 , n42534 );
and ( n42536 , n42431 , n42535 );
and ( n42537 , n42409 , n42535 );
or ( n42538 , n42432 , n42536 , n42537 );
and ( n42539 , n42406 , n42538 );
and ( n42540 , n42404 , n42538 );
or ( n42541 , n42407 , n42539 , n42540 );
xor ( n42542 , n42056 , n42058 );
xor ( n42543 , n42542 , n42130 );
and ( n42544 , n42541 , n42543 );
xor ( n42545 , n42296 , n42300 );
xor ( n42546 , n42545 , n42315 );
xor ( n42547 , n42319 , n42335 );
xor ( n42548 , n42547 , n42352 );
and ( n42549 , n42546 , n42548 );
xor ( n42550 , n42372 , n42381 );
xor ( n42551 , n42550 , n42398 );
and ( n42552 , n42548 , n42551 );
and ( n42553 , n42546 , n42551 );
or ( n42554 , n42549 , n42552 , n42553 );
xor ( n42555 , n42095 , n42097 );
xor ( n42556 , n42555 , n42124 );
and ( n42557 , n42554 , n42556 );
xor ( n42558 , n42318 , n42355 );
xor ( n42559 , n42558 , n42401 );
and ( n42560 , n42556 , n42559 );
and ( n42561 , n42554 , n42559 );
or ( n42562 , n42557 , n42560 , n42561 );
xor ( n42563 , n42061 , n42073 );
xor ( n42564 , n42563 , n42127 );
and ( n42565 , n42562 , n42564 );
xor ( n42566 , n42162 , n42166 );
xor ( n42567 , n42566 , n42171 );
and ( n42568 , n42564 , n42567 );
and ( n42569 , n42562 , n42567 );
or ( n42570 , n42565 , n42568 , n42569 );
and ( n42571 , n42543 , n42570 );
and ( n42572 , n42541 , n42570 );
or ( n42573 , n42544 , n42571 , n42572 );
and ( n42574 , n42291 , n42573 );
and ( n42575 , n42284 , n42573 );
or ( n42576 , n42292 , n42574 , n42575 );
and ( n42577 , n42281 , n42576 );
and ( n42578 , n42280 , n42576 );
or ( n42579 , n42282 , n42577 , n42578 );
and ( n42580 , n42263 , n42579 );
and ( n42581 , n42213 , n42579 );
or ( n42582 , n42264 , n42580 , n42581 );
and ( n42583 , n42211 , n42582 );
xor ( n42584 , n41821 , n41823 );
xor ( n42585 , n42584 , n41921 );
and ( n42586 , n42582 , n42585 );
and ( n42587 , n42211 , n42585 );
or ( n42588 , n42583 , n42586 , n42587 );
and ( n42589 , n41926 , n42588 );
and ( n42590 , n41924 , n42588 );
or ( n42591 , n41927 , n42589 , n42590 );
and ( n42592 , n41818 , n42591 );
and ( n42593 , n41816 , n42591 );
or ( n42594 , n41819 , n42592 , n42593 );
and ( n42595 , n41813 , n42594 );
and ( n42596 , n41811 , n42594 );
or ( n42597 , n41814 , n42595 , n42596 );
and ( n42598 , n41612 , n42597 );
and ( n42599 , n41610 , n42597 );
or ( n42600 , n41613 , n42598 , n42599 );
and ( n42601 , n41501 , n42600 );
and ( n42602 , n41499 , n42600 );
or ( n42603 , n41502 , n42601 , n42602 );
and ( n42604 , n41340 , n42603 );
and ( n42605 , n41338 , n42603 );
or ( n42606 , n41341 , n42604 , n42605 );
and ( n42607 , n41194 , n42606 );
and ( n42608 , n41192 , n42606 );
or ( n42609 , n41195 , n42607 , n42608 );
and ( n42610 , n41033 , n42609 );
and ( n42611 , n40869 , n42609 );
or ( n42612 , n41034 , n42610 , n42611 );
and ( n42613 , n40866 , n42612 );
and ( n42614 , n40659 , n42612 );
or ( n42615 , n40867 , n42613 , n42614 );
and ( n42616 , n40656 , n42615 );
and ( n42617 , n40654 , n42615 );
or ( n42618 , n40657 , n42616 , n42617 );
and ( n42619 , n40621 , n42618 );
and ( n42620 , n40619 , n42618 );
or ( n42621 , n40622 , n42619 , n42620 );
and ( n42622 , n40398 , n42621 );
and ( n42623 , n40396 , n42621 );
or ( n42624 , n40399 , n42622 , n42623 );
and ( n42625 , n40349 , n42624 );
and ( n42626 , n40347 , n42624 );
or ( n42627 , n40350 , n42625 , n42626 );
and ( n42628 , n40227 , n42627 );
and ( n42629 , n40225 , n42627 );
or ( n42630 , n40228 , n42628 , n42629 );
and ( n42631 , n40122 , n42630 );
and ( n42632 , n40120 , n42630 );
or ( n42633 , n40123 , n42631 , n42632 );
and ( n42634 , n39976 , n42633 );
and ( n42635 , n39974 , n42633 );
or ( n42636 , n39977 , n42634 , n42635 );
and ( n42637 , n39911 , n42636 );
and ( n42638 , n39788 , n42636 );
or ( n42639 , n39912 , n42637 , n42638 );
and ( n42640 , n39785 , n42639 );
and ( n42641 , n39783 , n42639 );
or ( n42642 , n39786 , n42640 , n42641 );
and ( n42643 , n39718 , n42642 );
and ( n42644 , n39716 , n42642 );
or ( n42645 , n39719 , n42643 , n42644 );
and ( n42646 , n39597 , n42645 );
and ( n42647 , n39595 , n42645 );
or ( n42648 , n39598 , n42646 , n42647 );
and ( n42649 , n39559 , n42648 );
and ( n42650 , n39557 , n42648 );
or ( n42651 , n39560 , n42649 , n42650 );
and ( n42652 , n39461 , n42651 );
and ( n42653 , n39459 , n42651 );
or ( n42654 , n39462 , n42652 , n42653 );
and ( n42655 , n39419 , n42654 );
and ( n42656 , n39417 , n42654 );
or ( n42657 , n39420 , n42655 , n42656 );
and ( n42658 , n39356 , n42657 );
and ( n42659 , n39290 , n42657 );
or ( n42660 , n39357 , n42658 , n42659 );
and ( n42661 , n39287 , n42660 );
and ( n42662 , n39285 , n42660 );
or ( n42663 , n39288 , n42661 , n42662 );
and ( n42664 , n39251 , n42663 );
xor ( n42665 , n39285 , n39287 );
xor ( n42666 , n42665 , n42660 );
xor ( n42667 , n39290 , n39356 );
xor ( n42668 , n42667 , n42657 );
xor ( n42669 , n39417 , n39419 );
xor ( n42670 , n42669 , n42654 );
xor ( n42671 , n39459 , n39461 );
xor ( n42672 , n42671 , n42651 );
xor ( n42673 , n39557 , n39559 );
xor ( n42674 , n42673 , n42648 );
xor ( n42675 , n39595 , n39597 );
xor ( n42676 , n42675 , n42645 );
xor ( n42677 , n39716 , n39718 );
xor ( n42678 , n42677 , n42642 );
xor ( n42679 , n39783 , n39785 );
xor ( n42680 , n42679 , n42639 );
xor ( n42681 , n39788 , n39911 );
xor ( n42682 , n42681 , n42636 );
xor ( n42683 , n39974 , n39976 );
xor ( n42684 , n42683 , n42633 );
xor ( n42685 , n40120 , n40122 );
xor ( n42686 , n42685 , n42630 );
xor ( n42687 , n40225 , n40227 );
xor ( n42688 , n42687 , n42627 );
xor ( n42689 , n40347 , n40349 );
xor ( n42690 , n42689 , n42624 );
xor ( n42691 , n40396 , n40398 );
xor ( n42692 , n42691 , n42621 );
xor ( n42693 , n40619 , n40621 );
xor ( n42694 , n42693 , n42618 );
xor ( n42695 , n40654 , n40656 );
xor ( n42696 , n42695 , n42615 );
xor ( n42697 , n40659 , n40866 );
xor ( n42698 , n42697 , n42612 );
xor ( n42699 , n40869 , n41033 );
xor ( n42700 , n42699 , n42609 );
xor ( n42701 , n41192 , n41194 );
xor ( n42702 , n42701 , n42606 );
xor ( n42703 , n41338 , n41340 );
xor ( n42704 , n42703 , n42603 );
xor ( n42705 , n41499 , n41501 );
xor ( n42706 , n42705 , n42600 );
xor ( n42707 , n41610 , n41612 );
xor ( n42708 , n42707 , n42597 );
xor ( n42709 , n41811 , n41813 );
xor ( n42710 , n42709 , n42594 );
xor ( n42711 , n41816 , n41818 );
xor ( n42712 , n42711 , n42591 );
xor ( n42713 , n41924 , n41926 );
xor ( n42714 , n42713 , n42588 );
xor ( n42715 , n41957 , n41959 );
xor ( n42716 , n42715 , n42208 );
xor ( n42717 , n42136 , n42138 );
xor ( n42718 , n42717 , n42205 );
xor ( n42719 , n42255 , n42257 );
xor ( n42720 , n42719 , n42260 );
and ( n42721 , n42718 , n42720 );
xor ( n42722 , n42247 , n42249 );
xor ( n42723 , n42722 , n42252 );
xor ( n42724 , n41946 , n41948 );
xor ( n42725 , n42724 , n41951 );
and ( n42726 , n42723 , n42725 );
and ( n42727 , n42720 , n42726 );
and ( n42728 , n42718 , n42726 );
or ( n42729 , n42721 , n42727 , n42728 );
and ( n42730 , n42716 , n42729 );
xor ( n42731 , n42213 , n42263 );
xor ( n42732 , n42731 , n42579 );
and ( n42733 , n42729 , n42732 );
and ( n42734 , n42716 , n42732 );
or ( n42735 , n42730 , n42733 , n42734 );
xor ( n42736 , n42211 , n42582 );
xor ( n42737 , n42736 , n42585 );
and ( n42738 , n42735 , n42737 );
xor ( n42739 , n42277 , n42279 );
xor ( n42740 , n41934 , n41938 );
xor ( n42741 , n42740 , n41943 );
xor ( n42742 , n42237 , n42241 );
xor ( n42743 , n42742 , n42244 );
and ( n42744 , n42741 , n42743 );
and ( n42745 , n42739 , n42744 );
and ( n42746 , n40069 , n39984 );
and ( n42747 , n39935 , n39982 );
nor ( n42748 , n42746 , n42747 );
xnor ( n42749 , n42748 , n39865 );
xor ( n42750 , n42153 , n42157 );
xor ( n42751 , n42750 , n42159 );
and ( n42752 , n42749 , n42751 );
xor ( n42753 , n42140 , n42144 );
xor ( n42754 , n42753 , n42150 );
xor ( n42755 , n42386 , n42390 );
xor ( n42756 , n42755 , n42395 );
and ( n42757 , n39657 , n40928 );
and ( n42758 , n39618 , n40926 );
nor ( n42759 , n42757 , n42758 );
xnor ( n42760 , n42759 , n40688 );
and ( n42761 , n39848 , n40666 );
and ( n42762 , n39739 , n40664 );
nor ( n42763 , n42761 , n42762 );
xnor ( n42764 , n42763 , n40445 );
and ( n42765 , n42760 , n42764 );
xor ( n42766 , n42446 , n42450 );
xor ( n42767 , n42766 , n42455 );
and ( n42768 , n42764 , n42767 );
and ( n42769 , n42760 , n42767 );
or ( n42770 , n42765 , n42768 , n42769 );
and ( n42771 , n42756 , n42770 );
buf ( n42772 , n30347 );
not ( n42773 , n42772 );
and ( n42774 , n41735 , n39335 );
and ( n42775 , n41364 , n39333 );
nor ( n42776 , n42774 , n42775 );
xnor ( n42777 , n42776 , n39300 );
and ( n42778 , n42149 , n39258 );
and ( n42779 , n41844 , n39256 );
nor ( n42780 , n42778 , n42779 );
xnor ( n42781 , n42780 , n39215 );
or ( n42782 , n42777 , n42781 );
and ( n42783 , n42773 , n42782 );
and ( n42784 , n42525 , n39194 );
and ( n42785 , n41828 , n39192 );
nor ( n42786 , n42784 , n42785 );
xnor ( n42787 , n42786 , n39199 );
buf ( n42788 , n30348 );
not ( n42789 , n42788 );
and ( n42790 , n42787 , n42789 );
and ( n42791 , n42782 , n42790 );
and ( n42792 , n42773 , n42790 );
or ( n42793 , n42783 , n42791 , n42792 );
and ( n42794 , n42770 , n42793 );
and ( n42795 , n42756 , n42793 );
or ( n42796 , n42771 , n42794 , n42795 );
and ( n42797 , n42754 , n42796 );
and ( n42798 , n39507 , n41522 );
and ( n42799 , n39433 , n41520 );
nor ( n42800 , n42798 , n42799 );
xnor ( n42801 , n42800 , n41100 );
and ( n42802 , n39618 , n41230 );
and ( n42803 , n39524 , n41228 );
nor ( n42804 , n42802 , n42803 );
xnor ( n42805 , n42804 , n40981 );
and ( n42806 , n42801 , n42805 );
and ( n42807 , n39739 , n40928 );
and ( n42808 , n39657 , n40926 );
nor ( n42809 , n42807 , n42808 );
xnor ( n42810 , n42809 , n40688 );
and ( n42811 , n42805 , n42810 );
and ( n42812 , n42801 , n42810 );
or ( n42813 , n42806 , n42811 , n42812 );
and ( n42814 , n39875 , n40666 );
and ( n42815 , n39848 , n40664 );
nor ( n42816 , n42814 , n42815 );
xnor ( n42817 , n42816 , n40445 );
and ( n42818 , n40069 , n40406 );
and ( n42819 , n39935 , n40404 );
nor ( n42820 , n42818 , n42819 );
xnor ( n42821 , n42820 , n40262 );
and ( n42822 , n42817 , n42821 );
and ( n42823 , n40272 , n40168 );
and ( n42824 , n40077 , n40166 );
nor ( n42825 , n42823 , n42824 );
xnor ( n42826 , n42825 , n40059 );
and ( n42827 , n42821 , n42826 );
and ( n42828 , n42817 , n42826 );
or ( n42829 , n42822 , n42827 , n42828 );
and ( n42830 , n42813 , n42829 );
and ( n42831 , n40455 , n39984 );
and ( n42832 , n40280 , n39982 );
nor ( n42833 , n42831 , n42832 );
xnor ( n42834 , n42833 , n39865 );
and ( n42835 , n40698 , n39795 );
and ( n42836 , n40574 , n39793 );
nor ( n42837 , n42835 , n42836 );
xnor ( n42838 , n42837 , n39729 );
and ( n42839 , n42834 , n42838 );
and ( n42840 , n40991 , n39665 );
and ( n42841 , n40962 , n39663 );
nor ( n42842 , n42840 , n42841 );
xnor ( n42843 , n42842 , n39608 );
and ( n42844 , n42838 , n42843 );
and ( n42845 , n42834 , n42843 );
or ( n42846 , n42839 , n42844 , n42845 );
and ( n42847 , n42829 , n42846 );
and ( n42848 , n42813 , n42846 );
or ( n42849 , n42830 , n42847 , n42848 );
and ( n42850 , n41106 , n39532 );
and ( n42851 , n40910 , n39530 );
nor ( n42852 , n42850 , n42851 );
xnor ( n42853 , n42852 , n39497 );
and ( n42854 , n41379 , n39384 );
and ( n42855 , n41091 , n39382 );
nor ( n42856 , n42854 , n42855 );
xnor ( n42857 , n42856 , n39367 );
and ( n42858 , n42853 , n42857 );
xor ( n42859 , n37168 , n39127 );
buf ( n42860 , n42859 );
buf ( n42861 , n42860 );
buf ( n42862 , n42861 );
and ( n42863 , n42862 , n39186 );
and ( n42864 , n42857 , n42863 );
and ( n42865 , n42853 , n42863 );
or ( n42866 , n42858 , n42864 , n42865 );
xor ( n42867 , n42463 , n42467 );
xor ( n42868 , n42867 , n42472 );
and ( n42869 , n42866 , n42868 );
xor ( n42870 , n42483 , n42487 );
xor ( n42871 , n42870 , n42492 );
and ( n42872 , n42868 , n42871 );
and ( n42873 , n42866 , n42871 );
or ( n42874 , n42869 , n42872 , n42873 );
and ( n42875 , n42849 , n42874 );
xor ( n42876 , n42418 , n42422 );
xor ( n42877 , n42876 , n42425 );
and ( n42878 , n42874 , n42877 );
and ( n42879 , n42849 , n42877 );
or ( n42880 , n42875 , n42878 , n42879 );
and ( n42881 , n42796 , n42880 );
and ( n42882 , n42754 , n42880 );
or ( n42883 , n42797 , n42881 , n42882 );
xor ( n42884 , n42434 , n42436 );
xor ( n42885 , n42884 , n42438 );
xor ( n42886 , n42442 , n42458 );
xor ( n42887 , n42886 , n42475 );
and ( n42888 , n42885 , n42887 );
xor ( n42889 , n42495 , n42511 );
xor ( n42890 , n42889 , n42529 );
and ( n42891 , n42887 , n42890 );
and ( n42892 , n42885 , n42890 );
or ( n42893 , n42888 , n42891 , n42892 );
xor ( n42894 , n42411 , n42413 );
xor ( n42895 , n42894 , n42428 );
and ( n42896 , n42893 , n42895 );
xor ( n42897 , n42441 , n42478 );
xor ( n42898 , n42897 , n42532 );
and ( n42899 , n42895 , n42898 );
and ( n42900 , n42893 , n42898 );
or ( n42901 , n42896 , n42899 , n42900 );
and ( n42902 , n42883 , n42901 );
xor ( n42903 , n42409 , n42431 );
xor ( n42904 , n42903 , n42535 );
and ( n42905 , n42901 , n42904 );
and ( n42906 , n42883 , n42904 );
or ( n42907 , n42902 , n42905 , n42906 );
and ( n42908 , n42752 , n42907 );
xor ( n42909 , n42404 , n42406 );
xor ( n42910 , n42909 , n42538 );
and ( n42911 , n42907 , n42910 );
and ( n42912 , n42752 , n42910 );
or ( n42913 , n42908 , n42911 , n42912 );
xor ( n42914 , n42268 , n42270 );
xor ( n42915 , n42914 , n42273 );
and ( n42916 , n42913 , n42915 );
xnor ( n42917 , n42288 , n42290 );
and ( n42918 , n42915 , n42917 );
and ( n42919 , n42913 , n42917 );
or ( n42920 , n42916 , n42918 , n42919 );
and ( n42921 , n42744 , n42920 );
and ( n42922 , n42739 , n42920 );
or ( n42923 , n42745 , n42921 , n42922 );
xor ( n42924 , n42280 , n42281 );
xor ( n42925 , n42924 , n42576 );
and ( n42926 , n42923 , n42925 );
and ( n42927 , n42111 , n42115 );
and ( n42928 , n42115 , n42120 );
and ( n42929 , n42111 , n42120 );
or ( n42930 , n42927 , n42928 , n42929 );
and ( n42931 , n39184 , n42079 );
not ( n42932 , n42931 );
xnor ( n42933 , n42932 , n41370 );
and ( n42934 , n42930 , n42933 );
and ( n42935 , n39875 , n40168 );
and ( n42936 , n39848 , n40166 );
nor ( n42937 , n42935 , n42936 );
xnor ( n42938 , n42937 , n40059 );
and ( n42939 , n42933 , n42938 );
and ( n42940 , n42930 , n42938 );
or ( n42941 , n42934 , n42939 , n42940 );
and ( n42942 , n39618 , n40666 );
and ( n42943 , n39524 , n40664 );
nor ( n42944 , n42942 , n42943 );
xnor ( n42945 , n42944 , n40445 );
and ( n42946 , n39739 , n40406 );
and ( n42947 , n39657 , n40404 );
nor ( n42948 , n42946 , n42947 );
xnor ( n42949 , n42948 , n40262 );
and ( n42950 , n42945 , n42949 );
xor ( n42951 , n42217 , n42221 );
xor ( n42952 , n42951 , n42224 );
and ( n42953 , n42949 , n42952 );
and ( n42954 , n42945 , n42952 );
or ( n42955 , n42950 , n42953 , n42954 );
and ( n42956 , n42941 , n42955 );
xor ( n42957 , n42227 , n42231 );
xor ( n42958 , n42957 , n42234 );
and ( n42959 , n42955 , n42958 );
and ( n42960 , n42941 , n42958 );
or ( n42961 , n42956 , n42959 , n42960 );
and ( n42962 , n42305 , n42309 );
and ( n42963 , n42309 , n42314 );
and ( n42964 , n42305 , n42314 );
or ( n42965 , n42962 , n42963 , n42964 );
xor ( n42966 , n42930 , n42933 );
xor ( n42967 , n42966 , n42938 );
and ( n42968 , n42965 , n42967 );
xor ( n42969 , n42945 , n42949 );
xor ( n42970 , n42969 , n42952 );
and ( n42971 , n42967 , n42970 );
and ( n42972 , n42965 , n42970 );
or ( n42973 , n42968 , n42971 , n42972 );
xor ( n42974 , n42554 , n42556 );
xor ( n42975 , n42974 , n42559 );
xor ( n42976 , n42749 , n42751 );
and ( n42977 , n42975 , n42976 );
xor ( n42978 , n42546 , n42548 );
xor ( n42979 , n42978 , n42551 );
xor ( n42980 , n42499 , n42503 );
xor ( n42981 , n42980 , n42508 );
xor ( n42982 , n42516 , n42520 );
xor ( n42983 , n42982 , n42526 );
and ( n42984 , n42981 , n42983 );
xor ( n42985 , n42760 , n42764 );
xor ( n42986 , n42985 , n42767 );
and ( n42987 , n42983 , n42986 );
and ( n42988 , n42981 , n42986 );
or ( n42989 , n42984 , n42987 , n42988 );
xnor ( n42990 , n42777 , n42781 );
xor ( n42991 , n42787 , n42789 );
and ( n42992 , n42990 , n42991 );
and ( n42993 , n40574 , n39984 );
and ( n42994 , n40455 , n39982 );
nor ( n42995 , n42993 , n42994 );
xnor ( n42996 , n42995 , n39865 );
and ( n42997 , n40962 , n39795 );
and ( n42998 , n40698 , n39793 );
nor ( n42999 , n42997 , n42998 );
xnor ( n43000 , n42999 , n39729 );
and ( n43001 , n42996 , n43000 );
and ( n43002 , n40910 , n39665 );
and ( n43003 , n40991 , n39663 );
nor ( n43004 , n43002 , n43003 );
xnor ( n43005 , n43004 , n39608 );
and ( n43006 , n43000 , n43005 );
and ( n43007 , n42996 , n43005 );
or ( n43008 , n43001 , n43006 , n43007 );
and ( n43009 , n42991 , n43008 );
and ( n43010 , n42990 , n43008 );
or ( n43011 , n42992 , n43009 , n43010 );
and ( n43012 , n39327 , n42079 );
and ( n43013 , n39310 , n42076 );
nor ( n43014 , n43012 , n43013 );
xnor ( n43015 , n43014 , n41370 );
and ( n43016 , n39433 , n41981 );
and ( n43017 , n39397 , n41979 );
nor ( n43018 , n43016 , n43017 );
xnor ( n43019 , n43018 , n41373 );
and ( n43020 , n43015 , n43019 );
and ( n43021 , n40280 , n40168 );
and ( n43022 , n40272 , n40166 );
nor ( n43023 , n43021 , n43022 );
xnor ( n43024 , n43023 , n40059 );
and ( n43025 , n43019 , n43024 );
and ( n43026 , n43015 , n43024 );
or ( n43027 , n43020 , n43025 , n43026 );
and ( n43028 , n41091 , n39532 );
and ( n43029 , n41106 , n39530 );
nor ( n43030 , n43028 , n43029 );
xnor ( n43031 , n43030 , n39497 );
and ( n43032 , n41364 , n39384 );
and ( n43033 , n41379 , n39382 );
nor ( n43034 , n43032 , n43033 );
xnor ( n43035 , n43034 , n39367 );
and ( n43036 , n43031 , n43035 );
xor ( n43037 , n37477 , n39125 );
buf ( n43038 , n43037 );
buf ( n43039 , n43038 );
buf ( n43040 , n43039 );
and ( n43041 , n43040 , n39186 );
and ( n43042 , n43035 , n43041 );
and ( n43043 , n43031 , n43041 );
or ( n43044 , n43036 , n43042 , n43043 );
and ( n43045 , n43027 , n43044 );
xor ( n43046 , n42801 , n42805 );
xor ( n43047 , n43046 , n42810 );
and ( n43048 , n43044 , n43047 );
and ( n43049 , n43027 , n43047 );
or ( n43050 , n43045 , n43048 , n43049 );
and ( n43051 , n43011 , n43050 );
xor ( n43052 , n42817 , n42821 );
xor ( n43053 , n43052 , n42826 );
xor ( n43054 , n42834 , n42838 );
xor ( n43055 , n43054 , n42843 );
and ( n43056 , n43053 , n43055 );
xor ( n43057 , n42853 , n42857 );
xor ( n43058 , n43057 , n42863 );
and ( n43059 , n43055 , n43058 );
and ( n43060 , n43053 , n43058 );
or ( n43061 , n43056 , n43059 , n43060 );
and ( n43062 , n43050 , n43061 );
and ( n43063 , n43011 , n43061 );
or ( n43064 , n43051 , n43062 , n43063 );
and ( n43065 , n42989 , n43064 );
xor ( n43066 , n42773 , n42782 );
xor ( n43067 , n43066 , n42790 );
xor ( n43068 , n42813 , n42829 );
xor ( n43069 , n43068 , n42846 );
and ( n43070 , n43067 , n43069 );
xor ( n43071 , n42866 , n42868 );
xor ( n43072 , n43071 , n42871 );
and ( n43073 , n43069 , n43072 );
and ( n43074 , n43067 , n43072 );
or ( n43075 , n43070 , n43073 , n43074 );
and ( n43076 , n43064 , n43075 );
and ( n43077 , n42989 , n43075 );
or ( n43078 , n43065 , n43076 , n43077 );
and ( n43079 , n42979 , n43078 );
xor ( n43080 , n42756 , n42770 );
xor ( n43081 , n43080 , n42793 );
xor ( n43082 , n42849 , n42874 );
xor ( n43083 , n43082 , n42877 );
and ( n43084 , n43081 , n43083 );
xor ( n43085 , n42885 , n42887 );
xor ( n43086 , n43085 , n42890 );
and ( n43087 , n43083 , n43086 );
and ( n43088 , n43081 , n43086 );
or ( n43089 , n43084 , n43087 , n43088 );
and ( n43090 , n43078 , n43089 );
and ( n43091 , n42979 , n43089 );
or ( n43092 , n43079 , n43090 , n43091 );
and ( n43093 , n42976 , n43092 );
and ( n43094 , n42975 , n43092 );
or ( n43095 , n42977 , n43093 , n43094 );
and ( n43096 , n42973 , n43095 );
xor ( n43097 , n42562 , n42564 );
xor ( n43098 , n43097 , n42567 );
and ( n43099 , n43095 , n43098 );
and ( n43100 , n42973 , n43098 );
or ( n43101 , n43096 , n43099 , n43100 );
and ( n43102 , n42961 , n43101 );
xor ( n43103 , n42541 , n42543 );
xor ( n43104 , n43103 , n42570 );
and ( n43105 , n43101 , n43104 );
and ( n43106 , n42961 , n43104 );
or ( n43107 , n43102 , n43105 , n43106 );
xor ( n43108 , n42284 , n42291 );
xor ( n43109 , n43108 , n42573 );
and ( n43110 , n43107 , n43109 );
xor ( n43111 , n42723 , n42725 );
and ( n43112 , n43109 , n43111 );
and ( n43113 , n43107 , n43111 );
or ( n43114 , n43110 , n43112 , n43113 );
and ( n43115 , n42925 , n43114 );
and ( n43116 , n42923 , n43114 );
or ( n43117 , n42926 , n43115 , n43116 );
xor ( n43118 , n42716 , n42729 );
xor ( n43119 , n43118 , n42732 );
and ( n43120 , n43117 , n43119 );
xor ( n43121 , n42718 , n42720 );
xor ( n43122 , n43121 , n42726 );
xor ( n43123 , n42741 , n42743 );
xor ( n43124 , n42752 , n42907 );
xor ( n43125 , n43124 , n42910 );
xor ( n43126 , n42941 , n42955 );
xor ( n43127 , n43126 , n42958 );
and ( n43128 , n43125 , n43127 );
xor ( n43129 , n42883 , n42901 );
xor ( n43130 , n43129 , n42904 );
xor ( n43131 , n42965 , n42967 );
xor ( n43132 , n43131 , n42970 );
and ( n43133 , n43130 , n43132 );
xor ( n43134 , n42754 , n42796 );
xor ( n43135 , n43134 , n42880 );
xor ( n43136 , n42893 , n42895 );
xor ( n43137 , n43136 , n42898 );
and ( n43138 , n43135 , n43137 );
xor ( n43139 , n37480 , n39123 );
buf ( n43140 , n43139 );
buf ( n43141 , n43140 );
buf ( n43142 , n43141 );
and ( n43143 , n43142 , n39186 );
buf ( n43144 , n30350 );
not ( n43145 , n43144 );
and ( n43146 , n43143 , n43145 );
and ( n43147 , n42862 , n39194 );
and ( n43148 , n42525 , n39192 );
nor ( n43149 , n43147 , n43148 );
xnor ( n43150 , n43149 , n39199 );
and ( n43151 , n43146 , n43150 );
buf ( n43152 , n30349 );
not ( n43153 , n43152 );
xor ( n43154 , n43015 , n43019 );
xor ( n43155 , n43154 , n43024 );
and ( n43156 , n43153 , n43155 );
xor ( n43157 , n43031 , n43035 );
xor ( n43158 , n43157 , n43041 );
and ( n43159 , n43155 , n43158 );
and ( n43160 , n43153 , n43158 );
or ( n43161 , n43156 , n43159 , n43160 );
and ( n43162 , n43151 , n43161 );
xor ( n43163 , n42990 , n42991 );
xor ( n43164 , n43163 , n43008 );
and ( n43165 , n43161 , n43164 );
and ( n43166 , n43151 , n43164 );
or ( n43167 , n43162 , n43165 , n43166 );
xor ( n43168 , n42981 , n42983 );
xor ( n43169 , n43168 , n42986 );
and ( n43170 , n43167 , n43169 );
xor ( n43171 , n43011 , n43050 );
xor ( n43172 , n43171 , n43061 );
and ( n43173 , n43169 , n43172 );
and ( n43174 , n43167 , n43172 );
or ( n43175 , n43170 , n43173 , n43174 );
xor ( n43176 , n42989 , n43064 );
xor ( n43177 , n43176 , n43075 );
and ( n43178 , n43175 , n43177 );
xor ( n43179 , n43081 , n43083 );
xor ( n43180 , n43179 , n43086 );
and ( n43181 , n43177 , n43180 );
and ( n43182 , n43175 , n43180 );
or ( n43183 , n43178 , n43181 , n43182 );
and ( n43184 , n43137 , n43183 );
and ( n43185 , n43135 , n43183 );
or ( n43186 , n43138 , n43184 , n43185 );
and ( n43187 , n43132 , n43186 );
and ( n43188 , n43130 , n43186 );
or ( n43189 , n43133 , n43187 , n43188 );
and ( n43190 , n43127 , n43189 );
and ( n43191 , n43125 , n43189 );
or ( n43192 , n43128 , n43190 , n43191 );
and ( n43193 , n43123 , n43192 );
xor ( n43194 , n42913 , n42915 );
xor ( n43195 , n43194 , n42917 );
and ( n43196 , n43192 , n43195 );
and ( n43197 , n43123 , n43195 );
or ( n43198 , n43193 , n43196 , n43197 );
xor ( n43199 , n42739 , n42744 );
xor ( n43200 , n43199 , n42920 );
and ( n43201 , n43198 , n43200 );
xor ( n43202 , n43107 , n43109 );
xor ( n43203 , n43202 , n43111 );
and ( n43204 , n43200 , n43203 );
and ( n43205 , n43198 , n43203 );
or ( n43206 , n43201 , n43204 , n43205 );
or ( n43207 , n43122 , n43206 );
and ( n43208 , n43119 , n43207 );
and ( n43209 , n43117 , n43207 );
or ( n43210 , n43120 , n43208 , n43209 );
and ( n43211 , n42737 , n43210 );
and ( n43212 , n42735 , n43210 );
or ( n43213 , n42738 , n43211 , n43212 );
or ( n43214 , n42714 , n43213 );
or ( n43215 , n42712 , n43214 );
or ( n43216 , n42710 , n43215 );
or ( n43217 , n42708 , n43216 );
or ( n43218 , n42706 , n43217 );
or ( n43219 , n42704 , n43218 );
or ( n43220 , n42702 , n43219 );
or ( n43221 , n42700 , n43220 );
or ( n43222 , n42698 , n43221 );
or ( n43223 , n42696 , n43222 );
or ( n43224 , n42694 , n43223 );
or ( n43225 , n42692 , n43224 );
or ( n43226 , n42690 , n43225 );
or ( n43227 , n42688 , n43226 );
or ( n43228 , n42686 , n43227 );
or ( n43229 , n42684 , n43228 );
or ( n43230 , n42682 , n43229 );
or ( n43231 , n42680 , n43230 );
or ( n43232 , n42678 , n43231 );
or ( n43233 , n42676 , n43232 );
or ( n43234 , n42674 , n43233 );
or ( n43235 , n42672 , n43234 );
or ( n43236 , n42670 , n43235 );
or ( n43237 , n42668 , n43236 );
or ( n43238 , n42666 , n43237 );
and ( n43239 , n42663 , n43238 );
and ( n43240 , n39251 , n43238 );
or ( n43241 , n42664 , n43239 , n43240 );
and ( n43242 , n39248 , n43241 );
buf ( n43243 , n43241 );
or ( n43244 , n39249 , n43242 , n43243 );
buf ( n43245 , n43244 );
not ( n43246 , n39248 );
xor ( n43247 , n43246 , n43241 );
not ( n43248 , n43247 );
xor ( n43249 , n39251 , n42663 );
xor ( n43250 , n43249 , n43238 );
xnor ( n43251 , n42666 , n43237 );
xnor ( n43252 , n42668 , n43236 );
xnor ( n43253 , n42670 , n43235 );
xnor ( n43254 , n42672 , n43234 );
xnor ( n43255 , n42674 , n43233 );
xnor ( n43256 , n42676 , n43232 );
xnor ( n43257 , n42678 , n43231 );
xnor ( n43258 , n42680 , n43230 );
xnor ( n43259 , n42682 , n43229 );
xnor ( n43260 , n42684 , n43228 );
xnor ( n43261 , n42686 , n43227 );
xnor ( n43262 , n42688 , n43226 );
xnor ( n43263 , n42690 , n43225 );
xnor ( n43264 , n42692 , n43224 );
xnor ( n43265 , n42694 , n43223 );
xnor ( n43266 , n42696 , n43222 );
xnor ( n43267 , n42698 , n43221 );
xnor ( n43268 , n42700 , n43220 );
xnor ( n43269 , n42702 , n43219 );
xnor ( n43270 , n42704 , n43218 );
xnor ( n43271 , n42706 , n43217 );
xnor ( n43272 , n42708 , n43216 );
xnor ( n43273 , n42710 , n43215 );
xnor ( n43274 , n42712 , n43214 );
xnor ( n43275 , n42714 , n43213 );
xor ( n43276 , n42735 , n42737 );
xor ( n43277 , n43276 , n43210 );
not ( n43278 , n43277 );
xor ( n43279 , n43117 , n43119 );
xor ( n43280 , n43279 , n43207 );
xor ( n43281 , n42923 , n42925 );
xor ( n43282 , n43281 , n43114 );
xnor ( n43283 , n43122 , n43206 );
and ( n43284 , n43282 , n43283 );
xor ( n43285 , n43282 , n43283 );
xor ( n43286 , n43198 , n43200 );
xor ( n43287 , n43286 , n43203 );
xor ( n43288 , n42961 , n43101 );
xor ( n43289 , n43288 , n43104 );
xor ( n43290 , n43123 , n43192 );
xor ( n43291 , n43290 , n43195 );
and ( n43292 , n43289 , n43291 );
xor ( n43293 , n42973 , n43095 );
xor ( n43294 , n43293 , n43098 );
xor ( n43295 , n43125 , n43127 );
xor ( n43296 , n43295 , n43189 );
and ( n43297 , n43294 , n43296 );
xor ( n43298 , n42975 , n42976 );
xor ( n43299 , n43298 , n43092 );
xor ( n43300 , n43130 , n43132 );
xor ( n43301 , n43300 , n43186 );
and ( n43302 , n43299 , n43301 );
xor ( n43303 , n42979 , n43078 );
xor ( n43304 , n43303 , n43089 );
xor ( n43305 , n43135 , n43137 );
xor ( n43306 , n43305 , n43183 );
and ( n43307 , n43304 , n43306 );
xor ( n43308 , n43067 , n43069 );
xor ( n43309 , n43308 , n43072 );
xor ( n43310 , n43027 , n43044 );
xor ( n43311 , n43310 , n43047 );
xor ( n43312 , n43053 , n43055 );
xor ( n43313 , n43312 , n43058 );
and ( n43314 , n43311 , n43313 );
and ( n43315 , n43142 , n39194 );
and ( n43316 , n43040 , n39192 );
nor ( n43317 , n43315 , n43316 );
xnor ( n43318 , n43317 , n39199 );
xor ( n43319 , n37482 , n39122 );
buf ( n43320 , n43319 );
buf ( n43321 , n43320 );
buf ( n43322 , n43321 );
and ( n43323 , n43322 , n39186 );
and ( n43324 , n43318 , n43323 );
and ( n43325 , n42525 , n39258 );
and ( n43326 , n41828 , n39256 );
nor ( n43327 , n43325 , n43326 );
xnor ( n43328 , n43327 , n39215 );
and ( n43329 , n43324 , n43328 );
and ( n43330 , n43040 , n39194 );
and ( n43331 , n42862 , n39192 );
nor ( n43332 , n43330 , n43331 );
xnor ( n43333 , n43332 , n39199 );
and ( n43334 , n43328 , n43333 );
and ( n43335 , n43324 , n43333 );
or ( n43336 , n43329 , n43334 , n43335 );
and ( n43337 , n41844 , n39335 );
and ( n43338 , n41735 , n39333 );
nor ( n43339 , n43337 , n43338 );
xnor ( n43340 , n43339 , n39300 );
and ( n43341 , n43336 , n43340 );
and ( n43342 , n41828 , n39258 );
and ( n43343 , n42149 , n39256 );
nor ( n43344 , n43342 , n43343 );
xnor ( n43345 , n43344 , n39215 );
and ( n43346 , n43340 , n43345 );
and ( n43347 , n43336 , n43345 );
or ( n43348 , n43341 , n43346 , n43347 );
and ( n43349 , n43313 , n43348 );
and ( n43350 , n43311 , n43348 );
or ( n43351 , n43314 , n43349 , n43350 );
and ( n43352 , n43309 , n43351 );
xor ( n43353 , n43167 , n43169 );
xor ( n43354 , n43353 , n43172 );
and ( n43355 , n43351 , n43354 );
and ( n43356 , n43309 , n43354 );
or ( n43357 , n43352 , n43355 , n43356 );
xor ( n43358 , n43175 , n43177 );
xor ( n43359 , n43358 , n43180 );
and ( n43360 , n43357 , n43359 );
xor ( n43361 , n43151 , n43161 );
xor ( n43362 , n43361 , n43164 );
and ( n43363 , n41379 , n39532 );
and ( n43364 , n41091 , n39530 );
nor ( n43365 , n43363 , n43364 );
xnor ( n43366 , n43365 , n39497 );
and ( n43367 , n41735 , n39384 );
and ( n43368 , n41364 , n39382 );
nor ( n43369 , n43367 , n43368 );
xnor ( n43370 , n43369 , n39367 );
and ( n43371 , n43366 , n43370 );
and ( n43372 , n42149 , n39335 );
and ( n43373 , n41844 , n39333 );
nor ( n43374 , n43372 , n43373 );
xnor ( n43375 , n43374 , n39300 );
and ( n43376 , n43370 , n43375 );
and ( n43377 , n43366 , n43375 );
or ( n43378 , n43371 , n43376 , n43377 );
xor ( n43379 , n43143 , n43145 );
and ( n43380 , n43322 , n39194 );
and ( n43381 , n43142 , n39192 );
nor ( n43382 , n43380 , n43381 );
xnor ( n43383 , n43382 , n39199 );
xor ( n43384 , n37750 , n39120 );
buf ( n43385 , n43384 );
buf ( n43386 , n43385 );
buf ( n43387 , n43386 );
and ( n43388 , n43387 , n39186 );
and ( n43389 , n43383 , n43388 );
and ( n43390 , n42862 , n39258 );
and ( n43391 , n42525 , n39256 );
nor ( n43392 , n43390 , n43391 );
xnor ( n43393 , n43392 , n39215 );
and ( n43394 , n43389 , n43393 );
buf ( n43395 , n30351 );
not ( n43396 , n43395 );
and ( n43397 , n43393 , n43396 );
and ( n43398 , n43389 , n43396 );
or ( n43399 , n43394 , n43397 , n43398 );
and ( n43400 , n43379 , n43399 );
xor ( n43401 , n43324 , n43328 );
xor ( n43402 , n43401 , n43333 );
and ( n43403 , n43399 , n43402 );
and ( n43404 , n43379 , n43402 );
or ( n43405 , n43400 , n43403 , n43404 );
and ( n43406 , n43378 , n43405 );
xor ( n43407 , n43336 , n43340 );
xor ( n43408 , n43407 , n43345 );
and ( n43409 , n43405 , n43408 );
and ( n43410 , n43378 , n43408 );
or ( n43411 , n43406 , n43409 , n43410 );
and ( n43412 , n43362 , n43411 );
xor ( n43413 , n43311 , n43313 );
xor ( n43414 , n43413 , n43348 );
and ( n43415 , n43411 , n43414 );
and ( n43416 , n43362 , n43414 );
or ( n43417 , n43412 , n43415 , n43416 );
xor ( n43418 , n43309 , n43351 );
xor ( n43419 , n43418 , n43354 );
and ( n43420 , n43417 , n43419 );
and ( n43421 , n39935 , n40666 );
and ( n43422 , n39875 , n40664 );
nor ( n43423 , n43421 , n43422 );
xnor ( n43424 , n43423 , n40445 );
and ( n43425 , n40077 , n40406 );
and ( n43426 , n40069 , n40404 );
nor ( n43427 , n43425 , n43426 );
xnor ( n43428 , n43427 , n40262 );
and ( n43429 , n43424 , n43428 );
xor ( n43430 , n43378 , n43405 );
xor ( n43431 , n43430 , n43408 );
and ( n43432 , n43428 , n43431 );
and ( n43433 , n43424 , n43431 );
or ( n43434 , n43429 , n43432 , n43433 );
and ( n43435 , n39310 , n42079 );
and ( n43436 , n39271 , n42076 );
nor ( n43437 , n43435 , n43436 );
xnor ( n43438 , n43437 , n41370 );
and ( n43439 , n43434 , n43438 );
and ( n43440 , n39397 , n41981 );
and ( n43441 , n39327 , n41979 );
nor ( n43442 , n43440 , n43441 );
xnor ( n43443 , n43442 , n41373 );
and ( n43444 , n43438 , n43443 );
and ( n43445 , n43434 , n43443 );
or ( n43446 , n43439 , n43444 , n43445 );
and ( n43447 , n43419 , n43446 );
and ( n43448 , n43417 , n43446 );
or ( n43449 , n43420 , n43447 , n43448 );
and ( n43450 , n43359 , n43449 );
and ( n43451 , n43357 , n43449 );
or ( n43452 , n43360 , n43450 , n43451 );
and ( n43453 , n43306 , n43452 );
and ( n43454 , n43304 , n43452 );
or ( n43455 , n43307 , n43453 , n43454 );
and ( n43456 , n43301 , n43455 );
and ( n43457 , n43299 , n43455 );
or ( n43458 , n43302 , n43456 , n43457 );
and ( n43459 , n43296 , n43458 );
and ( n43460 , n43294 , n43458 );
or ( n43461 , n43297 , n43459 , n43460 );
and ( n43462 , n43291 , n43461 );
and ( n43463 , n43289 , n43461 );
or ( n43464 , n43292 , n43462 , n43463 );
and ( n43465 , n43287 , n43464 );
xor ( n43466 , n43287 , n43464 );
xor ( n43467 , n43289 , n43291 );
xor ( n43468 , n43467 , n43461 );
not ( n43469 , n43468 );
xor ( n43470 , n43294 , n43296 );
xor ( n43471 , n43470 , n43458 );
xor ( n43472 , n43299 , n43301 );
xor ( n43473 , n43472 , n43455 );
xor ( n43474 , n43304 , n43306 );
xor ( n43475 , n43474 , n43452 );
xor ( n43476 , n43357 , n43359 );
xor ( n43477 , n43476 , n43449 );
and ( n43478 , n40455 , n40168 );
and ( n43479 , n40280 , n40166 );
nor ( n43480 , n43478 , n43479 );
xnor ( n43481 , n43480 , n40059 );
xor ( n43482 , n43366 , n43370 );
xor ( n43483 , n43482 , n43375 );
and ( n43484 , n43481 , n43483 );
xor ( n43485 , n43379 , n43399 );
xor ( n43486 , n43485 , n43402 );
and ( n43487 , n43483 , n43486 );
and ( n43488 , n43481 , n43486 );
or ( n43489 , n43484 , n43487 , n43488 );
and ( n43490 , n39524 , n41522 );
and ( n43491 , n39507 , n41520 );
nor ( n43492 , n43490 , n43491 );
xnor ( n43493 , n43492 , n41100 );
and ( n43494 , n43489 , n43493 );
xor ( n43495 , n42996 , n43000 );
xor ( n43496 , n43495 , n43005 );
and ( n43497 , n43493 , n43496 );
and ( n43498 , n43489 , n43496 );
or ( n43499 , n43494 , n43497 , n43498 );
xor ( n43500 , n43362 , n43411 );
xor ( n43501 , n43500 , n43414 );
and ( n43502 , n43499 , n43501 );
xor ( n43503 , n43434 , n43438 );
xor ( n43504 , n43503 , n43443 );
and ( n43505 , n43501 , n43504 );
and ( n43506 , n43499 , n43504 );
or ( n43507 , n43502 , n43505 , n43506 );
xor ( n43508 , n43417 , n43419 );
xor ( n43509 , n43508 , n43446 );
and ( n43510 , n43507 , n43509 );
xor ( n43511 , n43146 , n43150 );
xor ( n43512 , n43153 , n43155 );
xor ( n43513 , n43512 , n43158 );
and ( n43514 , n43511 , n43513 );
xor ( n43515 , n43318 , n43323 );
xor ( n43516 , n43383 , n43388 );
and ( n43517 , n43387 , n39194 );
and ( n43518 , n43322 , n39192 );
nor ( n43519 , n43517 , n43518 );
xnor ( n43520 , n43519 , n39199 );
xor ( n43521 , n38367 , n39118 );
buf ( n43522 , n43521 );
buf ( n43523 , n43522 );
buf ( n43524 , n43523 );
and ( n43525 , n43524 , n39186 );
and ( n43526 , n43520 , n43525 );
and ( n43527 , n43516 , n43526 );
buf ( n43528 , n30352 );
not ( n43529 , n43528 );
and ( n43530 , n43526 , n43529 );
and ( n43531 , n43516 , n43529 );
or ( n43532 , n43527 , n43530 , n43531 );
and ( n43533 , n43515 , n43532 );
and ( n43534 , n41828 , n39335 );
and ( n43535 , n42149 , n39333 );
nor ( n43536 , n43534 , n43535 );
xnor ( n43537 , n43536 , n39300 );
and ( n43538 , n43532 , n43537 );
and ( n43539 , n43515 , n43537 );
or ( n43540 , n43533 , n43538 , n43539 );
xor ( n43541 , n43520 , n43525 );
and ( n43542 , n43524 , n39194 );
and ( n43543 , n43387 , n39192 );
nor ( n43544 , n43542 , n43543 );
xnor ( n43545 , n43544 , n39199 );
xor ( n43546 , n38369 , n39117 );
buf ( n43547 , n43546 );
buf ( n43548 , n43547 );
buf ( n43549 , n43548 );
and ( n43550 , n43549 , n39186 );
and ( n43551 , n43545 , n43550 );
and ( n43552 , n43541 , n43551 );
buf ( n43553 , n30353 );
not ( n43554 , n43553 );
and ( n43555 , n43551 , n43554 );
and ( n43556 , n43541 , n43554 );
or ( n43557 , n43552 , n43555 , n43556 );
and ( n43558 , n42525 , n39335 );
and ( n43559 , n41828 , n39333 );
nor ( n43560 , n43558 , n43559 );
xnor ( n43561 , n43560 , n39300 );
and ( n43562 , n43557 , n43561 );
and ( n43563 , n43040 , n39258 );
and ( n43564 , n42862 , n39256 );
nor ( n43565 , n43563 , n43564 );
xnor ( n43566 , n43565 , n39215 );
and ( n43567 , n43561 , n43566 );
and ( n43568 , n43557 , n43566 );
or ( n43569 , n43562 , n43567 , n43568 );
and ( n43570 , n41844 , n39384 );
and ( n43571 , n41735 , n39382 );
nor ( n43572 , n43570 , n43571 );
xnor ( n43573 , n43572 , n39367 );
and ( n43574 , n43569 , n43573 );
xor ( n43575 , n43389 , n43393 );
xor ( n43576 , n43575 , n43396 );
and ( n43577 , n43573 , n43576 );
and ( n43578 , n43569 , n43576 );
or ( n43579 , n43574 , n43577 , n43578 );
and ( n43580 , n43540 , n43579 );
and ( n43581 , n41106 , n39665 );
and ( n43582 , n40910 , n39663 );
nor ( n43583 , n43581 , n43582 );
xnor ( n43584 , n43583 , n39608 );
and ( n43585 , n43579 , n43584 );
and ( n43586 , n43540 , n43584 );
or ( n43587 , n43580 , n43585 , n43586 );
and ( n43588 , n43513 , n43587 );
and ( n43589 , n43511 , n43587 );
or ( n43590 , n43514 , n43588 , n43589 );
and ( n43591 , n41379 , n39665 );
and ( n43592 , n41091 , n39663 );
nor ( n43593 , n43591 , n43592 );
xnor ( n43594 , n43593 , n39608 );
and ( n43595 , n42149 , n39384 );
and ( n43596 , n41844 , n39382 );
nor ( n43597 , n43595 , n43596 );
xnor ( n43598 , n43597 , n39367 );
and ( n43599 , n43594 , n43598 );
xor ( n43600 , n43557 , n43561 );
xor ( n43601 , n43600 , n43566 );
and ( n43602 , n43598 , n43601 );
and ( n43603 , n43594 , n43601 );
or ( n43604 , n43599 , n43602 , n43603 );
and ( n43605 , n40910 , n39795 );
and ( n43606 , n40991 , n39793 );
nor ( n43607 , n43605 , n43606 );
xnor ( n43608 , n43607 , n39729 );
and ( n43609 , n43604 , n43608 );
xor ( n43610 , n43515 , n43532 );
xor ( n43611 , n43610 , n43537 );
and ( n43612 , n43608 , n43611 );
and ( n43613 , n43604 , n43611 );
or ( n43614 , n43609 , n43612 , n43613 );
and ( n43615 , n40272 , n40406 );
and ( n43616 , n40077 , n40404 );
nor ( n43617 , n43615 , n43616 );
xnor ( n43618 , n43617 , n40262 );
and ( n43619 , n43614 , n43618 );
xor ( n43620 , n43540 , n43579 );
xor ( n43621 , n43620 , n43584 );
and ( n43622 , n43618 , n43621 );
and ( n43623 , n43614 , n43621 );
or ( n43624 , n43619 , n43622 , n43623 );
and ( n43625 , n40574 , n40168 );
and ( n43626 , n40455 , n40166 );
nor ( n43627 , n43625 , n43626 );
xnor ( n43628 , n43627 , n40059 );
and ( n43629 , n40962 , n39984 );
and ( n43630 , n40698 , n39982 );
nor ( n43631 , n43629 , n43630 );
xnor ( n43632 , n43631 , n39865 );
and ( n43633 , n43628 , n43632 );
xor ( n43634 , n43569 , n43573 );
xor ( n43635 , n43634 , n43576 );
and ( n43636 , n43632 , n43635 );
and ( n43637 , n43628 , n43635 );
or ( n43638 , n43633 , n43636 , n43637 );
and ( n43639 , n40069 , n40666 );
and ( n43640 , n39935 , n40664 );
nor ( n43641 , n43639 , n43640 );
xnor ( n43642 , n43641 , n40445 );
and ( n43643 , n43638 , n43642 );
xor ( n43644 , n43481 , n43483 );
xor ( n43645 , n43644 , n43486 );
and ( n43646 , n43642 , n43645 );
and ( n43647 , n43638 , n43645 );
or ( n43648 , n43643 , n43646 , n43647 );
and ( n43649 , n43624 , n43648 );
xor ( n43650 , n43424 , n43428 );
xor ( n43651 , n43650 , n43431 );
and ( n43652 , n43648 , n43651 );
and ( n43653 , n43624 , n43651 );
or ( n43654 , n43649 , n43652 , n43653 );
and ( n43655 , n43590 , n43654 );
xor ( n43656 , n43499 , n43501 );
xor ( n43657 , n43656 , n43504 );
and ( n43658 , n43654 , n43657 );
and ( n43659 , n43590 , n43657 );
or ( n43660 , n43655 , n43658 , n43659 );
and ( n43661 , n43509 , n43660 );
and ( n43662 , n43507 , n43660 );
or ( n43663 , n43510 , n43661 , n43662 );
and ( n43664 , n43477 , n43663 );
xor ( n43665 , n43507 , n43509 );
xor ( n43666 , n43665 , n43660 );
xor ( n43667 , n43545 , n43550 );
xor ( n43668 , n38372 , n39115 );
buf ( n43669 , n43668 );
buf ( n43670 , n43669 );
buf ( n43671 , n43670 );
and ( n43672 , n43671 , n39194 );
and ( n43673 , n43549 , n39192 );
nor ( n43674 , n43672 , n43673 );
xnor ( n43675 , n43674 , n39199 );
xor ( n43676 , n38375 , n39113 );
buf ( n43677 , n43676 );
buf ( n43678 , n43677 );
buf ( n43679 , n43678 );
and ( n43680 , n43679 , n39186 );
and ( n43681 , n43675 , n43680 );
and ( n43682 , n43671 , n39186 );
and ( n43683 , n43681 , n43682 );
and ( n43684 , n43667 , n43683 );
and ( n43685 , n43322 , n39258 );
and ( n43686 , n43142 , n39256 );
nor ( n43687 , n43685 , n43686 );
xnor ( n43688 , n43687 , n39215 );
and ( n43689 , n43683 , n43688 );
and ( n43690 , n43667 , n43688 );
or ( n43691 , n43684 , n43689 , n43690 );
and ( n43692 , n42862 , n39335 );
and ( n43693 , n42525 , n39333 );
nor ( n43694 , n43692 , n43693 );
xnor ( n43695 , n43694 , n39300 );
and ( n43696 , n43691 , n43695 );
and ( n43697 , n43142 , n39258 );
and ( n43698 , n43040 , n39256 );
nor ( n43699 , n43697 , n43698 );
xnor ( n43700 , n43699 , n39215 );
and ( n43701 , n43695 , n43700 );
and ( n43702 , n43691 , n43700 );
or ( n43703 , n43696 , n43701 , n43702 );
and ( n43704 , n41735 , n39532 );
and ( n43705 , n41364 , n39530 );
nor ( n43706 , n43704 , n43705 );
xnor ( n43707 , n43706 , n39497 );
and ( n43708 , n43703 , n43707 );
xor ( n43709 , n43516 , n43526 );
xor ( n43710 , n43709 , n43529 );
and ( n43711 , n43707 , n43710 );
and ( n43712 , n43703 , n43710 );
or ( n43713 , n43708 , n43711 , n43712 );
and ( n43714 , n41091 , n39665 );
and ( n43715 , n41106 , n39663 );
nor ( n43716 , n43714 , n43715 );
xnor ( n43717 , n43716 , n39608 );
and ( n43718 , n43713 , n43717 );
and ( n43719 , n41364 , n39532 );
and ( n43720 , n41379 , n39530 );
nor ( n43721 , n43719 , n43720 );
xnor ( n43722 , n43721 , n39497 );
and ( n43723 , n43717 , n43722 );
and ( n43724 , n43713 , n43722 );
or ( n43725 , n43718 , n43723 , n43724 );
and ( n43726 , n40698 , n39984 );
and ( n43727 , n40574 , n39982 );
nor ( n43728 , n43726 , n43727 );
xnor ( n43729 , n43728 , n39865 );
and ( n43730 , n43725 , n43729 );
and ( n43731 , n40991 , n39795 );
and ( n43732 , n40962 , n39793 );
nor ( n43733 , n43731 , n43732 );
xnor ( n43734 , n43733 , n39729 );
and ( n43735 , n43729 , n43734 );
and ( n43736 , n43725 , n43734 );
or ( n43737 , n43730 , n43735 , n43736 );
and ( n43738 , n39657 , n41230 );
and ( n43739 , n39618 , n41228 );
nor ( n43740 , n43738 , n43739 );
xnor ( n43741 , n43740 , n40981 );
and ( n43742 , n43737 , n43741 );
and ( n43743 , n39848 , n40928 );
and ( n43744 , n39739 , n40926 );
nor ( n43745 , n43743 , n43744 );
xnor ( n43746 , n43745 , n40688 );
and ( n43747 , n43741 , n43746 );
and ( n43748 , n43737 , n43746 );
or ( n43749 , n43742 , n43747 , n43748 );
xor ( n43750 , n43590 , n43654 );
xor ( n43751 , n43750 , n43657 );
and ( n43752 , n43749 , n43751 );
and ( n43753 , n39618 , n41522 );
and ( n43754 , n39524 , n41520 );
nor ( n43755 , n43753 , n43754 );
xnor ( n43756 , n43755 , n41100 );
and ( n43757 , n39739 , n41230 );
and ( n43758 , n39657 , n41228 );
nor ( n43759 , n43757 , n43758 );
xnor ( n43760 , n43759 , n40981 );
and ( n43761 , n43756 , n43760 );
and ( n43762 , n39875 , n40928 );
and ( n43763 , n39848 , n40926 );
nor ( n43764 , n43762 , n43763 );
xnor ( n43765 , n43764 , n40688 );
and ( n43766 , n43760 , n43765 );
and ( n43767 , n43756 , n43765 );
or ( n43768 , n43761 , n43766 , n43767 );
xor ( n43769 , n43737 , n43741 );
xor ( n43770 , n43769 , n43746 );
and ( n43771 , n43768 , n43770 );
xor ( n43772 , n43489 , n43493 );
xor ( n43773 , n43772 , n43496 );
and ( n43774 , n43770 , n43773 );
and ( n43775 , n43768 , n43773 );
or ( n43776 , n43771 , n43774 , n43775 );
and ( n43777 , n43751 , n43776 );
and ( n43778 , n43749 , n43776 );
or ( n43779 , n43752 , n43777 , n43778 );
and ( n43780 , n43666 , n43779 );
xor ( n43781 , n43681 , n43682 );
and ( n43782 , n43387 , n39258 );
and ( n43783 , n43322 , n39256 );
nor ( n43784 , n43782 , n43783 );
xnor ( n43785 , n43784 , n39215 );
and ( n43786 , n43781 , n43785 );
and ( n43787 , n43549 , n39194 );
and ( n43788 , n43524 , n39192 );
nor ( n43789 , n43787 , n43788 );
xnor ( n43790 , n43789 , n39199 );
and ( n43791 , n43785 , n43790 );
and ( n43792 , n43781 , n43790 );
or ( n43793 , n43786 , n43791 , n43792 );
buf ( n43794 , n30354 );
not ( n43795 , n43794 );
and ( n43796 , n43793 , n43795 );
xor ( n43797 , n43667 , n43683 );
xor ( n43798 , n43797 , n43688 );
and ( n43799 , n43795 , n43798 );
and ( n43800 , n43793 , n43798 );
or ( n43801 , n43796 , n43799 , n43800 );
and ( n43802 , n41828 , n39384 );
and ( n43803 , n42149 , n39382 );
nor ( n43804 , n43802 , n43803 );
xnor ( n43805 , n43804 , n39367 );
and ( n43806 , n43801 , n43805 );
xor ( n43807 , n43541 , n43551 );
xor ( n43808 , n43807 , n43554 );
and ( n43809 , n43805 , n43808 );
and ( n43810 , n43801 , n43808 );
or ( n43811 , n43806 , n43809 , n43810 );
xor ( n43812 , n43675 , n43680 );
and ( n43813 , n43679 , n39194 );
and ( n43814 , n43671 , n39192 );
nor ( n43815 , n43813 , n43814 );
xnor ( n43816 , n43815 , n39199 );
xor ( n43817 , n38377 , n39112 );
buf ( n43818 , n43817 );
buf ( n43819 , n43818 );
buf ( n43820 , n43819 );
and ( n43821 , n43820 , n39186 );
and ( n43822 , n43816 , n43821 );
and ( n43823 , n43812 , n43822 );
and ( n43824 , n43524 , n39258 );
and ( n43825 , n43387 , n39256 );
nor ( n43826 , n43824 , n43825 );
xnor ( n43827 , n43826 , n39215 );
and ( n43828 , n43822 , n43827 );
and ( n43829 , n43812 , n43827 );
or ( n43830 , n43823 , n43828 , n43829 );
and ( n43831 , n43142 , n39335 );
and ( n43832 , n43040 , n39333 );
nor ( n43833 , n43831 , n43832 );
xnor ( n43834 , n43833 , n39300 );
and ( n43835 , n43830 , n43834 );
buf ( n43836 , n30355 );
not ( n43837 , n43836 );
and ( n43838 , n43834 , n43837 );
and ( n43839 , n43830 , n43837 );
or ( n43840 , n43835 , n43838 , n43839 );
and ( n43841 , n42525 , n39384 );
and ( n43842 , n41828 , n39382 );
nor ( n43843 , n43841 , n43842 );
xnor ( n43844 , n43843 , n39367 );
and ( n43845 , n43840 , n43844 );
and ( n43846 , n43040 , n39335 );
and ( n43847 , n42862 , n39333 );
nor ( n43848 , n43846 , n43847 );
xnor ( n43849 , n43848 , n39300 );
and ( n43850 , n43844 , n43849 );
and ( n43851 , n43840 , n43849 );
or ( n43852 , n43845 , n43850 , n43851 );
and ( n43853 , n41844 , n39532 );
and ( n43854 , n41735 , n39530 );
nor ( n43855 , n43853 , n43854 );
xnor ( n43856 , n43855 , n39497 );
and ( n43857 , n43852 , n43856 );
xor ( n43858 , n43691 , n43695 );
xor ( n43859 , n43858 , n43700 );
and ( n43860 , n43856 , n43859 );
and ( n43861 , n43852 , n43859 );
or ( n43862 , n43857 , n43860 , n43861 );
and ( n43863 , n43811 , n43862 );
and ( n43864 , n41106 , n39795 );
and ( n43865 , n40910 , n39793 );
nor ( n43866 , n43864 , n43865 );
xnor ( n43867 , n43866 , n39729 );
and ( n43868 , n43862 , n43867 );
and ( n43869 , n43811 , n43867 );
or ( n43870 , n43863 , n43868 , n43869 );
and ( n43871 , n40280 , n40406 );
and ( n43872 , n40272 , n40404 );
nor ( n43873 , n43871 , n43872 );
xnor ( n43874 , n43873 , n40262 );
and ( n43875 , n43870 , n43874 );
xor ( n43876 , n43713 , n43717 );
xor ( n43877 , n43876 , n43722 );
and ( n43878 , n43874 , n43877 );
and ( n43879 , n43870 , n43877 );
or ( n43880 , n43875 , n43878 , n43879 );
and ( n43881 , n39397 , n42079 );
and ( n43882 , n39327 , n42076 );
nor ( n43883 , n43881 , n43882 );
xnor ( n43884 , n43883 , n41370 );
and ( n43885 , n43880 , n43884 );
xor ( n43886 , n43725 , n43729 );
xor ( n43887 , n43886 , n43734 );
and ( n43888 , n43884 , n43887 );
and ( n43889 , n43880 , n43887 );
or ( n43890 , n43885 , n43888 , n43889 );
and ( n43891 , n40698 , n40168 );
and ( n43892 , n40574 , n40166 );
nor ( n43893 , n43891 , n43892 );
xnor ( n43894 , n43893 , n40059 );
xor ( n43895 , n43594 , n43598 );
xor ( n43896 , n43895 , n43601 );
and ( n43897 , n43894 , n43896 );
xor ( n43898 , n43703 , n43707 );
xor ( n43899 , n43898 , n43710 );
and ( n43900 , n43896 , n43899 );
and ( n43901 , n43894 , n43899 );
or ( n43902 , n43897 , n43900 , n43901 );
and ( n43903 , n40077 , n40666 );
and ( n43904 , n40069 , n40664 );
nor ( n43905 , n43903 , n43904 );
xnor ( n43906 , n43905 , n40445 );
and ( n43907 , n43902 , n43906 );
xor ( n43908 , n43604 , n43608 );
xor ( n43909 , n43908 , n43611 );
and ( n43910 , n43906 , n43909 );
and ( n43911 , n43902 , n43909 );
or ( n43912 , n43907 , n43910 , n43911 );
and ( n43913 , n39507 , n41981 );
and ( n43914 , n39433 , n41979 );
nor ( n43915 , n43913 , n43914 );
xnor ( n43916 , n43915 , n41373 );
and ( n43917 , n43912 , n43916 );
xor ( n43918 , n43614 , n43618 );
xor ( n43919 , n43918 , n43621 );
and ( n43920 , n43916 , n43919 );
and ( n43921 , n43912 , n43919 );
or ( n43922 , n43917 , n43920 , n43921 );
and ( n43923 , n43890 , n43922 );
and ( n43924 , n41379 , n39795 );
and ( n43925 , n41091 , n39793 );
nor ( n43926 , n43924 , n43925 );
xnor ( n43927 , n43926 , n39729 );
and ( n43928 , n41735 , n39665 );
and ( n43929 , n41364 , n39663 );
nor ( n43930 , n43928 , n43929 );
xnor ( n43931 , n43930 , n39608 );
and ( n43932 , n43927 , n43931 );
xor ( n43933 , n43840 , n43844 );
xor ( n43934 , n43933 , n43849 );
and ( n43935 , n43931 , n43934 );
and ( n43936 , n43927 , n43934 );
or ( n43937 , n43932 , n43935 , n43936 );
and ( n43938 , n40910 , n39984 );
and ( n43939 , n40991 , n39982 );
nor ( n43940 , n43938 , n43939 );
xnor ( n43941 , n43940 , n39865 );
and ( n43942 , n43937 , n43941 );
xor ( n43943 , n43801 , n43805 );
xor ( n43944 , n43943 , n43808 );
and ( n43945 , n43941 , n43944 );
and ( n43946 , n43937 , n43944 );
or ( n43947 , n43942 , n43945 , n43946 );
and ( n43948 , n40272 , n40666 );
and ( n43949 , n40077 , n40664 );
nor ( n43950 , n43948 , n43949 );
xnor ( n43951 , n43950 , n40445 );
and ( n43952 , n43947 , n43951 );
xor ( n43953 , n43811 , n43862 );
xor ( n43954 , n43953 , n43867 );
and ( n43955 , n43951 , n43954 );
and ( n43956 , n43947 , n43954 );
or ( n43957 , n43952 , n43955 , n43956 );
and ( n43958 , n39433 , n42079 );
and ( n43959 , n39397 , n42076 );
nor ( n43960 , n43958 , n43959 );
xnor ( n43961 , n43960 , n41370 );
and ( n43962 , n43957 , n43961 );
xor ( n43963 , n43870 , n43874 );
xor ( n43964 , n43963 , n43877 );
and ( n43965 , n43961 , n43964 );
and ( n43966 , n43957 , n43964 );
or ( n43967 , n43962 , n43965 , n43966 );
xor ( n43968 , n43756 , n43760 );
xor ( n43969 , n43968 , n43765 );
and ( n43970 , n43967 , n43969 );
xor ( n43971 , n43880 , n43884 );
xor ( n43972 , n43971 , n43887 );
and ( n43973 , n43969 , n43972 );
and ( n43974 , n43967 , n43972 );
or ( n43975 , n43970 , n43973 , n43974 );
and ( n43976 , n39657 , n41522 );
and ( n43977 , n39618 , n41520 );
nor ( n43978 , n43976 , n43977 );
xnor ( n43979 , n43978 , n41100 );
and ( n43980 , n39848 , n41230 );
and ( n43981 , n39739 , n41228 );
nor ( n43982 , n43980 , n43981 );
xnor ( n43983 , n43982 , n40981 );
and ( n43984 , n43979 , n43983 );
and ( n43985 , n39935 , n40928 );
and ( n43986 , n39875 , n40926 );
nor ( n43987 , n43985 , n43986 );
xnor ( n43988 , n43987 , n40688 );
and ( n43989 , n43983 , n43988 );
and ( n43990 , n43979 , n43988 );
or ( n43991 , n43984 , n43989 , n43990 );
xor ( n43992 , n43816 , n43821 );
and ( n43993 , n43820 , n39194 );
and ( n43994 , n43679 , n39192 );
nor ( n43995 , n43993 , n43994 );
xnor ( n43996 , n43995 , n39199 );
xor ( n43997 , n39025 , n39110 );
buf ( n43998 , n43997 );
buf ( n43999 , n43998 );
buf ( n44000 , n43999 );
and ( n44001 , n44000 , n39186 );
and ( n44002 , n43996 , n44001 );
and ( n44003 , n43992 , n44002 );
and ( n44004 , n43387 , n39335 );
and ( n44005 , n43322 , n39333 );
nor ( n44006 , n44004 , n44005 );
xnor ( n44007 , n44006 , n39300 );
and ( n44008 , n44002 , n44007 );
and ( n44009 , n43992 , n44007 );
or ( n44010 , n44003 , n44008 , n44009 );
and ( n44011 , n43322 , n39335 );
and ( n44012 , n43142 , n39333 );
nor ( n44013 , n44011 , n44012 );
xnor ( n44014 , n44013 , n39300 );
and ( n44015 , n44010 , n44014 );
buf ( n44016 , n30356 );
not ( n44017 , n44016 );
and ( n44018 , n44014 , n44017 );
and ( n44019 , n44010 , n44017 );
or ( n44020 , n44015 , n44018 , n44019 );
and ( n44021 , n42862 , n39384 );
and ( n44022 , n42525 , n39382 );
nor ( n44023 , n44021 , n44022 );
xnor ( n44024 , n44023 , n39367 );
and ( n44025 , n44020 , n44024 );
xor ( n44026 , n43781 , n43785 );
xor ( n44027 , n44026 , n43790 );
and ( n44028 , n44024 , n44027 );
and ( n44029 , n44020 , n44027 );
or ( n44030 , n44025 , n44028 , n44029 );
and ( n44031 , n42149 , n39532 );
and ( n44032 , n41844 , n39530 );
nor ( n44033 , n44031 , n44032 );
xnor ( n44034 , n44033 , n39497 );
and ( n44035 , n44030 , n44034 );
xor ( n44036 , n43793 , n43795 );
xor ( n44037 , n44036 , n43798 );
and ( n44038 , n44034 , n44037 );
and ( n44039 , n44030 , n44037 );
or ( n44040 , n44035 , n44038 , n44039 );
and ( n44041 , n41091 , n39795 );
and ( n44042 , n41106 , n39793 );
nor ( n44043 , n44041 , n44042 );
xnor ( n44044 , n44043 , n39729 );
and ( n44045 , n44040 , n44044 );
and ( n44046 , n41364 , n39665 );
and ( n44047 , n41379 , n39663 );
nor ( n44048 , n44046 , n44047 );
xnor ( n44049 , n44048 , n39608 );
and ( n44050 , n44044 , n44049 );
and ( n44051 , n44040 , n44049 );
or ( n44052 , n44045 , n44050 , n44051 );
and ( n44053 , n40455 , n40406 );
and ( n44054 , n40280 , n40404 );
nor ( n44055 , n44053 , n44054 );
xnor ( n44056 , n44055 , n40262 );
and ( n44057 , n44052 , n44056 );
and ( n44058 , n40991 , n39984 );
and ( n44059 , n40962 , n39982 );
nor ( n44060 , n44058 , n44059 );
xnor ( n44061 , n44060 , n39865 );
and ( n44062 , n44056 , n44061 );
and ( n44063 , n44052 , n44061 );
or ( n44064 , n44057 , n44062 , n44063 );
and ( n44065 , n39524 , n41981 );
and ( n44066 , n39507 , n41979 );
nor ( n44067 , n44065 , n44066 );
xnor ( n44068 , n44067 , n41373 );
and ( n44069 , n44064 , n44068 );
xor ( n44070 , n43628 , n43632 );
xor ( n44071 , n44070 , n43635 );
and ( n44072 , n44068 , n44071 );
and ( n44073 , n44064 , n44071 );
or ( n44074 , n44069 , n44072 , n44073 );
and ( n44075 , n43991 , n44074 );
xor ( n44076 , n43638 , n43642 );
xor ( n44077 , n44076 , n43645 );
and ( n44078 , n44074 , n44077 );
and ( n44079 , n43991 , n44077 );
or ( n44080 , n44075 , n44078 , n44079 );
and ( n44081 , n43975 , n44080 );
xor ( n44082 , n43624 , n43648 );
xor ( n44083 , n44082 , n43651 );
and ( n44084 , n44080 , n44083 );
and ( n44085 , n43975 , n44083 );
or ( n44086 , n44081 , n44084 , n44085 );
and ( n44087 , n43923 , n44086 );
xor ( n44088 , n43511 , n43513 );
xor ( n44089 , n44088 , n43587 );
xor ( n44090 , n43768 , n43770 );
xor ( n44091 , n44090 , n43773 );
and ( n44092 , n44089 , n44091 );
xor ( n44093 , n43890 , n43922 );
and ( n44094 , n44091 , n44093 );
and ( n44095 , n44089 , n44093 );
or ( n44096 , n44092 , n44094 , n44095 );
and ( n44097 , n44086 , n44096 );
and ( n44098 , n43923 , n44096 );
or ( n44099 , n44087 , n44097 , n44098 );
and ( n44100 , n43779 , n44099 );
and ( n44101 , n43666 , n44099 );
or ( n44102 , n43780 , n44100 , n44101 );
and ( n44103 , n43663 , n44102 );
and ( n44104 , n43477 , n44102 );
or ( n44105 , n43664 , n44103 , n44104 );
or ( n44106 , n43475 , n44105 );
and ( n44107 , n43473 , n44106 );
xor ( n44108 , n43473 , n44106 );
xnor ( n44109 , n43475 , n44105 );
xor ( n44110 , n43477 , n43663 );
xor ( n44111 , n44110 , n44102 );
xor ( n44112 , n43749 , n43751 );
xor ( n44113 , n44112 , n43776 );
xor ( n44114 , n43975 , n44080 );
xor ( n44115 , n44114 , n44083 );
xor ( n44116 , n43967 , n43969 );
xor ( n44117 , n44116 , n43972 );
xor ( n44118 , n43991 , n44074 );
xor ( n44119 , n44118 , n44077 );
or ( n44120 , n44117 , n44119 );
and ( n44121 , n44115 , n44120 );
and ( n44122 , n39739 , n41522 );
and ( n44123 , n39657 , n41520 );
nor ( n44124 , n44122 , n44123 );
xnor ( n44125 , n44124 , n41100 );
and ( n44126 , n39875 , n41230 );
and ( n44127 , n39848 , n41228 );
nor ( n44128 , n44126 , n44127 );
xnor ( n44129 , n44128 , n40981 );
and ( n44130 , n44125 , n44129 );
xor ( n44131 , n44052 , n44056 );
xor ( n44132 , n44131 , n44061 );
and ( n44133 , n44129 , n44132 );
and ( n44134 , n44125 , n44132 );
or ( n44135 , n44130 , n44133 , n44134 );
and ( n44136 , n40574 , n40406 );
and ( n44137 , n40455 , n40404 );
nor ( n44138 , n44136 , n44137 );
xnor ( n44139 , n44138 , n40262 );
and ( n44140 , n40962 , n40168 );
and ( n44141 , n40698 , n40166 );
nor ( n44142 , n44140 , n44141 );
xnor ( n44143 , n44142 , n40059 );
and ( n44144 , n44139 , n44143 );
xor ( n44145 , n43852 , n43856 );
xor ( n44146 , n44145 , n43859 );
and ( n44147 , n44143 , n44146 );
and ( n44148 , n44139 , n44146 );
or ( n44149 , n44144 , n44147 , n44148 );
and ( n44150 , n40069 , n40928 );
and ( n44151 , n39935 , n40926 );
nor ( n44152 , n44150 , n44151 );
xnor ( n44153 , n44152 , n40688 );
and ( n44154 , n44149 , n44153 );
xor ( n44155 , n43894 , n43896 );
xor ( n44156 , n44155 , n43899 );
and ( n44157 , n44153 , n44156 );
and ( n44158 , n44149 , n44156 );
or ( n44159 , n44154 , n44157 , n44158 );
and ( n44160 , n44135 , n44159 );
xor ( n44161 , n43902 , n43906 );
xor ( n44162 , n44161 , n43909 );
and ( n44163 , n44159 , n44162 );
and ( n44164 , n44135 , n44162 );
or ( n44165 , n44160 , n44163 , n44164 );
xor ( n44166 , n43912 , n43916 );
xor ( n44167 , n44166 , n43919 );
and ( n44168 , n44165 , n44167 );
and ( n44169 , n44120 , n44168 );
and ( n44170 , n44115 , n44168 );
or ( n44171 , n44121 , n44169 , n44170 );
and ( n44172 , n44113 , n44171 );
xor ( n44173 , n43923 , n44086 );
xor ( n44174 , n44173 , n44096 );
and ( n44175 , n44171 , n44174 );
and ( n44176 , n44113 , n44174 );
or ( n44177 , n44172 , n44175 , n44176 );
xor ( n44178 , n43666 , n43779 );
xor ( n44179 , n44178 , n44099 );
and ( n44180 , n44177 , n44179 );
xor ( n44181 , n44089 , n44091 );
xor ( n44182 , n44181 , n44093 );
xor ( n44183 , n43979 , n43983 );
xor ( n44184 , n44183 , n43988 );
xor ( n44185 , n44064 , n44068 );
xor ( n44186 , n44185 , n44071 );
or ( n44187 , n44184 , n44186 );
xnor ( n44188 , n44117 , n44119 );
and ( n44189 , n44187 , n44188 );
xor ( n44190 , n44165 , n44167 );
and ( n44191 , n44188 , n44190 );
and ( n44192 , n44187 , n44190 );
or ( n44193 , n44189 , n44191 , n44192 );
and ( n44194 , n44182 , n44193 );
xor ( n44195 , n44115 , n44120 );
xor ( n44196 , n44195 , n44168 );
and ( n44197 , n44193 , n44196 );
and ( n44198 , n44182 , n44196 );
or ( n44199 , n44194 , n44197 , n44198 );
xor ( n44200 , n44113 , n44171 );
xor ( n44201 , n44200 , n44174 );
and ( n44202 , n44199 , n44201 );
and ( n44203 , n39507 , n42079 );
and ( n44204 , n39433 , n42076 );
nor ( n44205 , n44203 , n44204 );
xnor ( n44206 , n44205 , n41370 );
and ( n44207 , n39618 , n41981 );
and ( n44208 , n39524 , n41979 );
nor ( n44209 , n44207 , n44208 );
xnor ( n44210 , n44209 , n41373 );
and ( n44211 , n44206 , n44210 );
and ( n44212 , n40280 , n40666 );
and ( n44213 , n40272 , n40664 );
nor ( n44214 , n44212 , n44213 );
xnor ( n44215 , n44214 , n40445 );
and ( n44216 , n39618 , n42079 );
and ( n44217 , n39524 , n42076 );
nor ( n44218 , n44216 , n44217 );
xnor ( n44219 , n44218 , n41370 );
and ( n44220 , n40272 , n40928 );
and ( n44221 , n40077 , n40926 );
nor ( n44222 , n44220 , n44221 );
xnor ( n44223 , n44222 , n40688 );
and ( n44224 , n44219 , n44223 );
and ( n44225 , n41106 , n39984 );
and ( n44226 , n40910 , n39982 );
nor ( n44227 , n44225 , n44226 );
xnor ( n44228 , n44227 , n39865 );
and ( n44229 , n44223 , n44228 );
and ( n44230 , n44219 , n44228 );
or ( n44231 , n44224 , n44229 , n44230 );
and ( n44232 , n44215 , n44231 );
and ( n44233 , n39657 , n42079 );
and ( n44234 , n39618 , n42076 );
nor ( n44235 , n44233 , n44234 );
xnor ( n44236 , n44235 , n41370 );
and ( n44237 , n39935 , n41522 );
and ( n44238 , n39875 , n41520 );
nor ( n44239 , n44237 , n44238 );
xnor ( n44240 , n44239 , n41100 );
and ( n44241 , n44236 , n44240 );
and ( n44242 , n40077 , n41230 );
and ( n44243 , n40069 , n41228 );
nor ( n44244 , n44242 , n44243 );
xnor ( n44245 , n44244 , n40981 );
and ( n44246 , n44240 , n44245 );
and ( n44247 , n44236 , n44245 );
or ( n44248 , n44241 , n44246 , n44247 );
and ( n44249 , n40574 , n40666 );
and ( n44250 , n40455 , n40664 );
nor ( n44251 , n44249 , n44250 );
xnor ( n44252 , n44251 , n40445 );
and ( n44253 , n40962 , n40406 );
and ( n44254 , n40698 , n40404 );
nor ( n44255 , n44253 , n44254 );
xnor ( n44256 , n44255 , n40262 );
and ( n44257 , n44252 , n44256 );
and ( n44258 , n40910 , n40168 );
and ( n44259 , n40991 , n40166 );
nor ( n44260 , n44258 , n44259 );
xnor ( n44261 , n44260 , n40059 );
and ( n44262 , n44256 , n44261 );
and ( n44263 , n44252 , n44261 );
or ( n44264 , n44257 , n44262 , n44263 );
and ( n44265 , n44248 , n44264 );
xor ( n44266 , n44219 , n44223 );
xor ( n44267 , n44266 , n44228 );
and ( n44268 , n44264 , n44267 );
and ( n44269 , n44248 , n44267 );
or ( n44270 , n44265 , n44268 , n44269 );
and ( n44271 , n44231 , n44270 );
and ( n44272 , n44215 , n44270 );
or ( n44273 , n44232 , n44271 , n44272 );
and ( n44274 , n44210 , n44273 );
and ( n44275 , n44206 , n44273 );
or ( n44276 , n44211 , n44274 , n44275 );
and ( n44277 , n40991 , n40168 );
and ( n44278 , n40962 , n40166 );
nor ( n44279 , n44277 , n44278 );
xnor ( n44280 , n44279 , n40059 );
xor ( n44281 , n43927 , n43931 );
xor ( n44282 , n44281 , n43934 );
and ( n44283 , n44280 , n44282 );
xor ( n44284 , n44030 , n44034 );
xor ( n44285 , n44284 , n44037 );
and ( n44286 , n44282 , n44285 );
and ( n44287 , n44280 , n44285 );
or ( n44288 , n44283 , n44286 , n44287 );
and ( n44289 , n39848 , n41522 );
and ( n44290 , n39739 , n41520 );
nor ( n44291 , n44289 , n44290 );
xnor ( n44292 , n44291 , n41100 );
and ( n44293 , n44288 , n44292 );
xor ( n44294 , n44139 , n44143 );
xor ( n44295 , n44294 , n44146 );
and ( n44296 , n44292 , n44295 );
and ( n44297 , n44288 , n44295 );
or ( n44298 , n44293 , n44296 , n44297 );
xor ( n44299 , n44149 , n44153 );
xor ( n44300 , n44299 , n44156 );
or ( n44301 , n44298 , n44300 );
and ( n44302 , n44276 , n44301 );
xor ( n44303 , n44135 , n44159 );
xor ( n44304 , n44303 , n44162 );
and ( n44305 , n44301 , n44304 );
and ( n44306 , n44276 , n44304 );
or ( n44307 , n44302 , n44305 , n44306 );
buf ( n44308 , n30357 );
not ( n44309 , n44308 );
xor ( n44310 , n43996 , n44001 );
and ( n44311 , n44000 , n39194 );
and ( n44312 , n43820 , n39192 );
nor ( n44313 , n44311 , n44312 );
xnor ( n44314 , n44313 , n39199 );
xor ( n44315 , n39026 , n39109 );
buf ( n44316 , n44315 );
buf ( n44317 , n44316 );
buf ( n44318 , n44317 );
and ( n44319 , n44318 , n39186 );
and ( n44320 , n44314 , n44319 );
and ( n44321 , n44310 , n44320 );
and ( n44322 , n43671 , n39258 );
and ( n44323 , n43549 , n39256 );
nor ( n44324 , n44322 , n44323 );
xnor ( n44325 , n44324 , n39215 );
and ( n44326 , n44320 , n44325 );
and ( n44327 , n44310 , n44325 );
or ( n44328 , n44321 , n44326 , n44327 );
not ( n44329 , n44328 );
and ( n44330 , n43549 , n39258 );
and ( n44331 , n43524 , n39256 );
nor ( n44332 , n44330 , n44331 );
xnor ( n44333 , n44332 , n39215 );
xor ( n44334 , n44329 , n44333 );
xnor ( n44335 , n44309 , n44334 );
and ( n44336 , n43820 , n39258 );
and ( n44337 , n43679 , n39256 );
nor ( n44338 , n44336 , n44337 );
xnor ( n44339 , n44338 , n39215 );
and ( n44340 , n44318 , n39194 );
and ( n44341 , n44000 , n39192 );
nor ( n44342 , n44340 , n44341 );
xnor ( n44343 , n44342 , n39199 );
xor ( n44344 , n39029 , n39107 );
buf ( n44345 , n44344 );
buf ( n44346 , n44345 );
buf ( n44347 , n44346 );
and ( n44348 , n44347 , n39186 );
xor ( n44349 , n44343 , n44348 );
and ( n44350 , n44339 , n44349 );
and ( n44351 , n43387 , n39384 );
and ( n44352 , n43322 , n39382 );
nor ( n44353 , n44351 , n44352 );
xnor ( n44354 , n44353 , n39367 );
and ( n44355 , n44350 , n44354 );
xor ( n44356 , n44314 , n44319 );
and ( n44357 , n44343 , n44348 );
xor ( n44358 , n44356 , n44357 );
and ( n44359 , n43679 , n39258 );
and ( n44360 , n43671 , n39256 );
nor ( n44361 , n44359 , n44360 );
xnor ( n44362 , n44361 , n39215 );
xor ( n44363 , n44358 , n44362 );
and ( n44364 , n44354 , n44363 );
and ( n44365 , n44350 , n44363 );
or ( n44366 , n44355 , n44364 , n44365 );
and ( n44367 , n43322 , n39384 );
and ( n44368 , n43142 , n39382 );
nor ( n44369 , n44367 , n44368 );
xnor ( n44370 , n44369 , n39367 );
and ( n44371 , n44366 , n44370 );
buf ( n44372 , n30358 );
not ( n44373 , n44372 );
and ( n44374 , n44370 , n44373 );
and ( n44375 , n44366 , n44373 );
or ( n44376 , n44371 , n44374 , n44375 );
and ( n44377 , n44335 , n44376 );
and ( n44378 , n42862 , n39532 );
and ( n44379 , n42525 , n39530 );
nor ( n44380 , n44378 , n44379 );
xnor ( n44381 , n44380 , n39497 );
and ( n44382 , n44376 , n44381 );
and ( n44383 , n44335 , n44381 );
or ( n44384 , n44377 , n44382 , n44383 );
and ( n44385 , n41735 , n39795 );
and ( n44386 , n41364 , n39793 );
nor ( n44387 , n44385 , n44386 );
xnor ( n44388 , n44387 , n39729 );
and ( n44389 , n44384 , n44388 );
and ( n44390 , n42149 , n39665 );
and ( n44391 , n41844 , n39663 );
nor ( n44392 , n44390 , n44391 );
xnor ( n44393 , n44392 , n39608 );
and ( n44394 , n44388 , n44393 );
and ( n44395 , n44384 , n44393 );
or ( n44396 , n44389 , n44394 , n44395 );
and ( n44397 , n41091 , n39984 );
and ( n44398 , n41106 , n39982 );
nor ( n44399 , n44397 , n44398 );
xnor ( n44400 , n44399 , n39865 );
and ( n44401 , n44396 , n44400 );
and ( n44402 , n41364 , n39795 );
and ( n44403 , n41379 , n39793 );
nor ( n44404 , n44402 , n44403 );
xnor ( n44405 , n44404 , n39729 );
and ( n44406 , n44400 , n44405 );
and ( n44407 , n44396 , n44405 );
or ( n44408 , n44401 , n44406 , n44407 );
and ( n44409 , n40455 , n40666 );
and ( n44410 , n40280 , n40664 );
nor ( n44411 , n44409 , n44410 );
xnor ( n44412 , n44411 , n40445 );
and ( n44413 , n44408 , n44412 );
and ( n44414 , n40698 , n40406 );
and ( n44415 , n40574 , n40404 );
nor ( n44416 , n44414 , n44415 );
xnor ( n44417 , n44416 , n40262 );
and ( n44418 , n44412 , n44417 );
and ( n44419 , n44408 , n44417 );
or ( n44420 , n44413 , n44418 , n44419 );
and ( n44421 , n39524 , n42079 );
and ( n44422 , n39507 , n42076 );
nor ( n44423 , n44421 , n44422 );
xnor ( n44424 , n44423 , n41370 );
and ( n44425 , n44420 , n44424 );
and ( n44426 , n39657 , n41981 );
and ( n44427 , n39618 , n41979 );
nor ( n44428 , n44426 , n44427 );
xnor ( n44429 , n44428 , n41373 );
and ( n44430 , n44424 , n44429 );
and ( n44431 , n44420 , n44429 );
or ( n44432 , n44425 , n44430 , n44431 );
and ( n44433 , n39935 , n41230 );
and ( n44434 , n39875 , n41228 );
nor ( n44435 , n44433 , n44434 );
xnor ( n44436 , n44435 , n40981 );
and ( n44437 , n40077 , n40928 );
and ( n44438 , n40069 , n40926 );
nor ( n44439 , n44437 , n44438 );
xnor ( n44440 , n44439 , n40688 );
and ( n44441 , n44436 , n44440 );
xor ( n44442 , n43937 , n43941 );
xor ( n44443 , n44442 , n43944 );
and ( n44444 , n44440 , n44443 );
and ( n44445 , n44436 , n44443 );
or ( n44446 , n44441 , n44444 , n44445 );
and ( n44447 , n44432 , n44446 );
xor ( n44448 , n43947 , n43951 );
xor ( n44449 , n44448 , n43954 );
and ( n44450 , n44446 , n44449 );
and ( n44451 , n44432 , n44449 );
or ( n44452 , n44447 , n44450 , n44451 );
xor ( n44453 , n43957 , n43961 );
xor ( n44454 , n44453 , n43964 );
or ( n44455 , n44452 , n44454 );
and ( n44456 , n44307 , n44455 );
xnor ( n44457 , n44184 , n44186 );
xor ( n44458 , n44206 , n44210 );
xor ( n44459 , n44458 , n44273 );
xor ( n44460 , n44215 , n44231 );
xor ( n44461 , n44460 , n44270 );
and ( n44462 , n39739 , n42079 );
and ( n44463 , n39657 , n42076 );
nor ( n44464 , n44462 , n44463 );
xnor ( n44465 , n44464 , n41370 );
and ( n44466 , n39875 , n41981 );
and ( n44467 , n39848 , n41979 );
nor ( n44468 , n44466 , n44467 );
xnor ( n44469 , n44468 , n41373 );
or ( n44470 , n44465 , n44469 );
and ( n44471 , n40991 , n40406 );
and ( n44472 , n40962 , n40404 );
nor ( n44473 , n44471 , n44472 );
xnor ( n44474 , n44473 , n40262 );
and ( n44475 , n41379 , n39984 );
and ( n44476 , n41091 , n39982 );
nor ( n44477 , n44475 , n44476 );
xnor ( n44478 , n44477 , n39865 );
and ( n44479 , n44474 , n44478 );
and ( n44480 , n42525 , n39532 );
and ( n44481 , n41828 , n39530 );
nor ( n44482 , n44480 , n44481 );
xnor ( n44483 , n44482 , n39497 );
and ( n44484 , n44478 , n44483 );
and ( n44485 , n44474 , n44483 );
or ( n44486 , n44479 , n44484 , n44485 );
and ( n44487 , n44470 , n44486 );
xor ( n44488 , n44236 , n44240 );
xor ( n44489 , n44488 , n44245 );
and ( n44490 , n44486 , n44489 );
and ( n44491 , n44470 , n44489 );
or ( n44492 , n44487 , n44490 , n44491 );
xor ( n44493 , n44248 , n44264 );
xor ( n44494 , n44493 , n44267 );
and ( n44495 , n44492 , n44494 );
and ( n44496 , n41828 , n39532 );
and ( n44497 , n42149 , n39530 );
nor ( n44498 , n44496 , n44497 );
xnor ( n44499 , n44498 , n39497 );
xor ( n44500 , n43830 , n43834 );
xor ( n44501 , n44500 , n43837 );
and ( n44502 , n44499 , n44501 );
and ( n44503 , n44494 , n44502 );
and ( n44504 , n44492 , n44502 );
or ( n44505 , n44495 , n44503 , n44504 );
and ( n44506 , n44461 , n44505 );
xor ( n44507 , n44040 , n44044 );
xor ( n44508 , n44507 , n44049 );
and ( n44509 , n44505 , n44508 );
and ( n44510 , n44461 , n44508 );
or ( n44511 , n44506 , n44509 , n44510 );
and ( n44512 , n44459 , n44511 );
xor ( n44513 , n44125 , n44129 );
xor ( n44514 , n44513 , n44132 );
and ( n44515 , n44511 , n44514 );
and ( n44516 , n44459 , n44514 );
or ( n44517 , n44512 , n44515 , n44516 );
and ( n44518 , n44457 , n44517 );
xnor ( n44519 , n44298 , n44300 );
xor ( n44520 , n44252 , n44256 );
xor ( n44521 , n44520 , n44261 );
xor ( n44522 , n44470 , n44486 );
xor ( n44523 , n44522 , n44489 );
and ( n44524 , n44521 , n44523 );
xnor ( n44525 , n44465 , n44469 );
xor ( n44526 , n44474 , n44478 );
xor ( n44527 , n44526 , n44483 );
and ( n44528 , n44525 , n44527 );
xor ( n44529 , n43812 , n43822 );
xor ( n44530 , n44529 , n43827 );
and ( n44531 , n44527 , n44530 );
and ( n44532 , n44525 , n44530 );
or ( n44533 , n44528 , n44531 , n44532 );
and ( n44534 , n44523 , n44533 );
and ( n44535 , n44521 , n44533 );
or ( n44536 , n44524 , n44534 , n44535 );
xor ( n44537 , n44499 , n44501 );
and ( n44538 , n39848 , n42079 );
and ( n44539 , n39739 , n42076 );
nor ( n44540 , n44538 , n44539 );
xnor ( n44541 , n44540 , n41370 );
and ( n44542 , n39935 , n41981 );
and ( n44543 , n39875 , n41979 );
nor ( n44544 , n44542 , n44543 );
xnor ( n44545 , n44544 , n41373 );
and ( n44546 , n44541 , n44545 );
and ( n44547 , n40272 , n41522 );
and ( n44548 , n40077 , n41520 );
nor ( n44549 , n44547 , n44548 );
xnor ( n44550 , n44549 , n41100 );
and ( n44551 , n40455 , n41230 );
and ( n44552 , n40280 , n41228 );
nor ( n44553 , n44551 , n44552 );
xnor ( n44554 , n44553 , n40981 );
and ( n44555 , n44550 , n44554 );
and ( n44556 , n40698 , n40928 );
and ( n44557 , n40574 , n40926 );
nor ( n44558 , n44556 , n44557 );
xnor ( n44559 , n44558 , n40688 );
and ( n44560 , n44554 , n44559 );
and ( n44561 , n44550 , n44559 );
or ( n44562 , n44555 , n44560 , n44561 );
and ( n44563 , n44545 , n44562 );
and ( n44564 , n44541 , n44562 );
or ( n44565 , n44546 , n44563 , n44564 );
and ( n44566 , n44329 , n44333 );
and ( n44567 , n44565 , n44566 );
buf ( n44568 , n44328 );
and ( n44569 , n44566 , n44568 );
and ( n44570 , n44565 , n44568 );
or ( n44571 , n44567 , n44569 , n44570 );
and ( n44572 , n44537 , n44571 );
xor ( n44573 , n44521 , n44523 );
xor ( n44574 , n44573 , n44533 );
and ( n44575 , n44571 , n44574 );
and ( n44576 , n44537 , n44574 );
or ( n44577 , n44572 , n44575 , n44576 );
and ( n44578 , n44536 , n44577 );
xor ( n44579 , n44492 , n44494 );
xor ( n44580 , n44579 , n44502 );
and ( n44581 , n44577 , n44580 );
and ( n44582 , n44536 , n44580 );
or ( n44583 , n44578 , n44581 , n44582 );
xor ( n44584 , n44288 , n44292 );
xor ( n44585 , n44584 , n44295 );
and ( n44586 , n44583 , n44585 );
and ( n44587 , n40069 , n41230 );
and ( n44588 , n39935 , n41228 );
nor ( n44589 , n44587 , n44588 );
xnor ( n44590 , n44589 , n40981 );
xor ( n44591 , n44280 , n44282 );
xor ( n44592 , n44591 , n44285 );
or ( n44593 , n44590 , n44592 );
and ( n44594 , n44585 , n44593 );
and ( n44595 , n44583 , n44593 );
or ( n44596 , n44586 , n44594 , n44595 );
and ( n44597 , n44519 , n44596 );
xor ( n44598 , n44461 , n44505 );
xor ( n44599 , n44598 , n44508 );
and ( n44600 , n44356 , n44357 );
and ( n44601 , n44357 , n44362 );
and ( n44602 , n44356 , n44362 );
or ( n44603 , n44600 , n44601 , n44602 );
and ( n44604 , n43524 , n39335 );
and ( n44605 , n43387 , n39333 );
nor ( n44606 , n44604 , n44605 );
xnor ( n44607 , n44606 , n39300 );
and ( n44608 , n44603 , n44607 );
xor ( n44609 , n44310 , n44320 );
xor ( n44610 , n44609 , n44325 );
and ( n44611 , n44607 , n44610 );
and ( n44612 , n44603 , n44610 );
or ( n44613 , n44608 , n44611 , n44612 );
and ( n44614 , n43142 , n39384 );
and ( n44615 , n43040 , n39382 );
nor ( n44616 , n44614 , n44615 );
xnor ( n44617 , n44616 , n39367 );
and ( n44618 , n44613 , n44617 );
xor ( n44619 , n43992 , n44002 );
xor ( n44620 , n44619 , n44007 );
and ( n44621 , n44617 , n44620 );
and ( n44622 , n44613 , n44620 );
or ( n44623 , n44618 , n44621 , n44622 );
and ( n44624 , n43040 , n39384 );
and ( n44625 , n42862 , n39382 );
nor ( n44626 , n44624 , n44625 );
xnor ( n44627 , n44626 , n39367 );
and ( n44628 , n44623 , n44627 );
xor ( n44629 , n44010 , n44014 );
xor ( n44630 , n44629 , n44017 );
and ( n44631 , n44627 , n44630 );
and ( n44632 , n44623 , n44630 );
or ( n44633 , n44628 , n44631 , n44632 );
and ( n44634 , n41844 , n39665 );
and ( n44635 , n41735 , n39663 );
nor ( n44636 , n44634 , n44635 );
xnor ( n44637 , n44636 , n39608 );
and ( n44638 , n44633 , n44637 );
xor ( n44639 , n44020 , n44024 );
xor ( n44640 , n44639 , n44027 );
and ( n44641 , n44637 , n44640 );
and ( n44642 , n44633 , n44640 );
or ( n44643 , n44638 , n44641 , n44642 );
xor ( n44644 , n44536 , n44577 );
xor ( n44645 , n44644 , n44580 );
and ( n44646 , n44643 , n44645 );
xnor ( n44647 , n44590 , n44592 );
and ( n44648 , n44645 , n44647 );
and ( n44649 , n44643 , n44647 );
or ( n44650 , n44646 , n44648 , n44649 );
and ( n44651 , n44599 , n44650 );
xor ( n44652 , n44583 , n44585 );
xor ( n44653 , n44652 , n44593 );
and ( n44654 , n44650 , n44653 );
and ( n44655 , n44599 , n44653 );
or ( n44656 , n44651 , n44654 , n44655 );
and ( n44657 , n44596 , n44656 );
and ( n44658 , n44519 , n44656 );
or ( n44659 , n44597 , n44657 , n44658 );
and ( n44660 , n44517 , n44659 );
and ( n44661 , n44457 , n44659 );
or ( n44662 , n44518 , n44660 , n44661 );
and ( n44663 , n44455 , n44662 );
and ( n44664 , n44307 , n44662 );
or ( n44665 , n44456 , n44663 , n44664 );
xor ( n44666 , n44182 , n44193 );
xor ( n44667 , n44666 , n44196 );
and ( n44668 , n44665 , n44667 );
xor ( n44669 , n44187 , n44188 );
xor ( n44670 , n44669 , n44190 );
xor ( n44671 , n44276 , n44301 );
xor ( n44672 , n44671 , n44304 );
xnor ( n44673 , n44452 , n44454 );
and ( n44674 , n44672 , n44673 );
xor ( n44675 , n44459 , n44511 );
xor ( n44676 , n44675 , n44514 );
xor ( n44677 , n44432 , n44446 );
xor ( n44678 , n44677 , n44449 );
and ( n44679 , n44676 , n44678 );
and ( n44680 , n39739 , n41981 );
and ( n44681 , n39657 , n41979 );
nor ( n44682 , n44680 , n44681 );
xnor ( n44683 , n44682 , n41373 );
and ( n44684 , n39875 , n41522 );
and ( n44685 , n39848 , n41520 );
nor ( n44686 , n44684 , n44685 );
xnor ( n44687 , n44686 , n41100 );
and ( n44688 , n44683 , n44687 );
xor ( n44689 , n44408 , n44412 );
xor ( n44690 , n44689 , n44417 );
and ( n44691 , n44687 , n44690 );
and ( n44692 , n44683 , n44690 );
or ( n44693 , n44688 , n44691 , n44692 );
xor ( n44694 , n44420 , n44424 );
xor ( n44695 , n44694 , n44429 );
and ( n44696 , n44693 , n44695 );
xor ( n44697 , n44436 , n44440 );
xor ( n44698 , n44697 , n44443 );
and ( n44699 , n44695 , n44698 );
and ( n44700 , n44693 , n44698 );
or ( n44701 , n44696 , n44699 , n44700 );
and ( n44702 , n44678 , n44701 );
and ( n44703 , n44676 , n44701 );
or ( n44704 , n44679 , n44702 , n44703 );
and ( n44705 , n44673 , n44704 );
and ( n44706 , n44672 , n44704 );
or ( n44707 , n44674 , n44705 , n44706 );
and ( n44708 , n44670 , n44707 );
xor ( n44709 , n44307 , n44455 );
xor ( n44710 , n44709 , n44662 );
and ( n44711 , n44707 , n44710 );
and ( n44712 , n44670 , n44710 );
or ( n44713 , n44708 , n44711 , n44712 );
and ( n44714 , n44667 , n44713 );
and ( n44715 , n44665 , n44713 );
or ( n44716 , n44668 , n44714 , n44715 );
and ( n44717 , n44201 , n44716 );
and ( n44718 , n44199 , n44716 );
or ( n44719 , n44202 , n44717 , n44718 );
and ( n44720 , n44179 , n44719 );
and ( n44721 , n44177 , n44719 );
or ( n44722 , n44180 , n44720 , n44721 );
and ( n44723 , n44111 , n44722 );
xor ( n44724 , n44111 , n44722 );
xor ( n44725 , n44177 , n44179 );
xor ( n44726 , n44725 , n44719 );
not ( n44727 , n44726 );
xor ( n44728 , n44199 , n44201 );
xor ( n44729 , n44728 , n44716 );
xor ( n44730 , n44665 , n44667 );
xor ( n44731 , n44730 , n44713 );
xor ( n44732 , n44457 , n44517 );
xor ( n44733 , n44732 , n44659 );
xor ( n44734 , n44519 , n44596 );
xor ( n44735 , n44734 , n44656 );
and ( n44736 , n40574 , n41230 );
and ( n44737 , n40455 , n41228 );
nor ( n44738 , n44736 , n44737 );
xnor ( n44739 , n44738 , n40981 );
and ( n44740 , n40962 , n40928 );
and ( n44741 , n40698 , n40926 );
nor ( n44742 , n44740 , n44741 );
xnor ( n44743 , n44742 , n40688 );
and ( n44744 , n44739 , n44743 );
and ( n44745 , n40910 , n40666 );
and ( n44746 , n40991 , n40664 );
nor ( n44747 , n44745 , n44746 );
xnor ( n44748 , n44747 , n40445 );
and ( n44749 , n44743 , n44748 );
and ( n44750 , n44739 , n44748 );
or ( n44751 , n44744 , n44749 , n44750 );
and ( n44752 , n39875 , n42079 );
and ( n44753 , n39848 , n42076 );
nor ( n44754 , n44752 , n44753 );
xnor ( n44755 , n44754 , n41370 );
and ( n44756 , n44751 , n44755 );
and ( n44757 , n40069 , n41981 );
and ( n44758 , n39935 , n41979 );
nor ( n44759 , n44757 , n44758 );
xnor ( n44760 , n44759 , n41373 );
and ( n44761 , n44755 , n44760 );
and ( n44762 , n44751 , n44760 );
or ( n44763 , n44756 , n44761 , n44762 );
and ( n44764 , n40991 , n40666 );
and ( n44765 , n40962 , n40664 );
nor ( n44766 , n44764 , n44765 );
xnor ( n44767 , n44766 , n40445 );
and ( n44768 , n41106 , n40406 );
and ( n44769 , n40910 , n40404 );
nor ( n44770 , n44768 , n44769 );
xnor ( n44771 , n44770 , n40262 );
and ( n44772 , n44767 , n44771 );
and ( n44773 , n39935 , n42079 );
and ( n44774 , n39875 , n42076 );
nor ( n44775 , n44773 , n44774 );
xnor ( n44776 , n44775 , n41370 );
and ( n44777 , n40077 , n41981 );
and ( n44778 , n40069 , n41979 );
nor ( n44779 , n44777 , n44778 );
xnor ( n44780 , n44779 , n41373 );
and ( n44781 , n44776 , n44780 );
and ( n44782 , n40280 , n41522 );
and ( n44783 , n40272 , n41520 );
nor ( n44784 , n44782 , n44783 );
xnor ( n44785 , n44784 , n41100 );
and ( n44786 , n44780 , n44785 );
and ( n44787 , n44776 , n44785 );
or ( n44788 , n44781 , n44786 , n44787 );
and ( n44789 , n44771 , n44788 );
and ( n44790 , n44767 , n44788 );
or ( n44791 , n44772 , n44789 , n44790 );
and ( n44792 , n44763 , n44791 );
xor ( n44793 , n44541 , n44545 );
xor ( n44794 , n44793 , n44562 );
and ( n44795 , n44791 , n44794 );
and ( n44796 , n44763 , n44794 );
or ( n44797 , n44792 , n44795 , n44796 );
xor ( n44798 , n44525 , n44527 );
xor ( n44799 , n44798 , n44530 );
and ( n44800 , n44797 , n44799 );
or ( n44801 , n44309 , n44334 );
and ( n44802 , n44799 , n44801 );
and ( n44803 , n44797 , n44801 );
or ( n44804 , n44800 , n44802 , n44803 );
xor ( n44805 , n44537 , n44571 );
xor ( n44806 , n44805 , n44574 );
and ( n44807 , n44804 , n44806 );
xor ( n44808 , n44633 , n44637 );
xor ( n44809 , n44808 , n44640 );
and ( n44810 , n44806 , n44809 );
and ( n44811 , n44804 , n44809 );
or ( n44812 , n44807 , n44810 , n44811 );
xor ( n44813 , n44339 , n44349 );
and ( n44814 , n44000 , n39258 );
and ( n44815 , n43820 , n39256 );
nor ( n44816 , n44814 , n44815 );
xnor ( n44817 , n44816 , n39215 );
and ( n44818 , n44347 , n39194 );
and ( n44819 , n44318 , n39192 );
nor ( n44820 , n44818 , n44819 );
xnor ( n44821 , n44820 , n39199 );
and ( n44822 , n44817 , n44821 );
xor ( n44823 , n39030 , n39106 );
buf ( n44824 , n44823 );
buf ( n44825 , n44824 );
buf ( n44826 , n44825 );
and ( n44827 , n44826 , n39186 );
and ( n44828 , n44821 , n44827 );
and ( n44829 , n44817 , n44827 );
or ( n44830 , n44822 , n44828 , n44829 );
and ( n44831 , n44813 , n44830 );
and ( n44832 , n43671 , n39335 );
and ( n44833 , n43549 , n39333 );
nor ( n44834 , n44832 , n44833 );
xnor ( n44835 , n44834 , n39300 );
and ( n44836 , n44830 , n44835 );
and ( n44837 , n44813 , n44835 );
or ( n44838 , n44831 , n44836 , n44837 );
and ( n44839 , n43549 , n39335 );
and ( n44840 , n43524 , n39333 );
nor ( n44841 , n44839 , n44840 );
xnor ( n44842 , n44841 , n39300 );
and ( n44843 , n44838 , n44842 );
buf ( n44844 , n30359 );
not ( n44845 , n44844 );
and ( n44846 , n44842 , n44845 );
and ( n44847 , n44838 , n44845 );
or ( n44848 , n44843 , n44846 , n44847 );
and ( n44849 , n43040 , n39532 );
and ( n44850 , n42862 , n39530 );
nor ( n44851 , n44849 , n44850 );
xnor ( n44852 , n44851 , n39497 );
and ( n44853 , n44848 , n44852 );
xor ( n44854 , n44603 , n44607 );
xor ( n44855 , n44854 , n44610 );
and ( n44856 , n44852 , n44855 );
and ( n44857 , n44848 , n44855 );
or ( n44858 , n44853 , n44856 , n44857 );
and ( n44859 , n41828 , n39665 );
and ( n44860 , n42149 , n39663 );
nor ( n44861 , n44859 , n44860 );
xnor ( n44862 , n44861 , n39608 );
and ( n44863 , n44858 , n44862 );
xor ( n44864 , n44613 , n44617 );
xor ( n44865 , n44864 , n44620 );
and ( n44866 , n44862 , n44865 );
and ( n44867 , n44858 , n44865 );
or ( n44868 , n44863 , n44866 , n44867 );
and ( n44869 , n41106 , n40168 );
and ( n44870 , n40910 , n40166 );
nor ( n44871 , n44869 , n44870 );
xnor ( n44872 , n44871 , n40059 );
and ( n44873 , n44868 , n44872 );
xor ( n44874 , n44384 , n44388 );
xor ( n44875 , n44874 , n44393 );
and ( n44876 , n44872 , n44875 );
and ( n44877 , n44868 , n44875 );
or ( n44878 , n44873 , n44876 , n44877 );
and ( n44879 , n40280 , n40928 );
and ( n44880 , n40272 , n40926 );
nor ( n44881 , n44879 , n44880 );
xnor ( n44882 , n44881 , n40688 );
and ( n44883 , n44878 , n44882 );
xor ( n44884 , n44396 , n44400 );
xor ( n44885 , n44884 , n44405 );
and ( n44886 , n44882 , n44885 );
and ( n44887 , n44878 , n44885 );
or ( n44888 , n44883 , n44886 , n44887 );
and ( n44889 , n44812 , n44888 );
and ( n44890 , n41091 , n40406 );
and ( n44891 , n41106 , n40404 );
nor ( n44892 , n44890 , n44891 );
xnor ( n44893 , n44892 , n40262 );
and ( n44894 , n41364 , n40168 );
and ( n44895 , n41379 , n40166 );
nor ( n44896 , n44894 , n44895 );
xnor ( n44897 , n44896 , n40059 );
and ( n44898 , n44893 , n44897 );
and ( n44899 , n41844 , n39984 );
and ( n44900 , n41735 , n39982 );
nor ( n44901 , n44899 , n44900 );
xnor ( n44902 , n44901 , n39865 );
and ( n44903 , n44897 , n44902 );
and ( n44904 , n44893 , n44902 );
or ( n44905 , n44898 , n44903 , n44904 );
xor ( n44906 , n44550 , n44554 );
xor ( n44907 , n44906 , n44559 );
and ( n44908 , n44905 , n44907 );
xor ( n44909 , n44751 , n44755 );
xor ( n44910 , n44909 , n44760 );
and ( n44911 , n44907 , n44910 );
and ( n44912 , n44905 , n44910 );
or ( n44913 , n44908 , n44911 , n44912 );
xor ( n44914 , n44739 , n44743 );
xor ( n44915 , n44914 , n44748 );
and ( n44916 , n40698 , n41230 );
and ( n44917 , n40574 , n41228 );
nor ( n44918 , n44916 , n44917 );
xnor ( n44919 , n44918 , n40981 );
and ( n44920 , n40991 , n40928 );
and ( n44921 , n40962 , n40926 );
nor ( n44922 , n44920 , n44921 );
xnor ( n44923 , n44922 , n40688 );
or ( n44924 , n44919 , n44923 );
and ( n44925 , n44915 , n44924 );
and ( n44926 , n40069 , n42079 );
and ( n44927 , n39935 , n42076 );
nor ( n44928 , n44926 , n44927 );
xnor ( n44929 , n44928 , n41370 );
and ( n44930 , n40272 , n41981 );
and ( n44931 , n40077 , n41979 );
nor ( n44932 , n44930 , n44931 );
xnor ( n44933 , n44932 , n41373 );
and ( n44934 , n44929 , n44933 );
and ( n44935 , n40455 , n41522 );
and ( n44936 , n40280 , n41520 );
nor ( n44937 , n44935 , n44936 );
xnor ( n44938 , n44937 , n41100 );
and ( n44939 , n44933 , n44938 );
and ( n44940 , n44929 , n44938 );
or ( n44941 , n44934 , n44939 , n44940 );
and ( n44942 , n44924 , n44941 );
and ( n44943 , n44915 , n44941 );
or ( n44944 , n44925 , n44942 , n44943 );
and ( n44945 , n41106 , n40666 );
and ( n44946 , n40910 , n40664 );
nor ( n44947 , n44945 , n44946 );
xnor ( n44948 , n44947 , n40445 );
and ( n44949 , n41379 , n40406 );
and ( n44950 , n41091 , n40404 );
nor ( n44951 , n44949 , n44950 );
xnor ( n44952 , n44951 , n40262 );
and ( n44953 , n44948 , n44952 );
and ( n44954 , n41735 , n40168 );
and ( n44955 , n41364 , n40166 );
nor ( n44956 , n44954 , n44955 );
xnor ( n44957 , n44956 , n40059 );
and ( n44958 , n44952 , n44957 );
and ( n44959 , n44948 , n44957 );
or ( n44960 , n44953 , n44958 , n44959 );
xor ( n44961 , n44776 , n44780 );
xor ( n44962 , n44961 , n44785 );
and ( n44963 , n44960 , n44962 );
xor ( n44964 , n44893 , n44897 );
xor ( n44965 , n44964 , n44902 );
and ( n44966 , n44962 , n44965 );
and ( n44967 , n44960 , n44965 );
or ( n44968 , n44963 , n44966 , n44967 );
and ( n44969 , n44944 , n44968 );
xor ( n44970 , n44767 , n44771 );
xor ( n44971 , n44970 , n44788 );
and ( n44972 , n44968 , n44971 );
and ( n44973 , n44944 , n44971 );
or ( n44974 , n44969 , n44972 , n44973 );
and ( n44975 , n44913 , n44974 );
xor ( n44976 , n44763 , n44791 );
xor ( n44977 , n44976 , n44794 );
and ( n44978 , n44974 , n44977 );
and ( n44979 , n44913 , n44977 );
or ( n44980 , n44975 , n44978 , n44979 );
xor ( n44981 , n44565 , n44566 );
xor ( n44982 , n44981 , n44568 );
and ( n44983 , n44980 , n44982 );
xor ( n44984 , n44623 , n44627 );
xor ( n44985 , n44984 , n44630 );
and ( n44986 , n44982 , n44985 );
and ( n44987 , n44980 , n44985 );
or ( n44988 , n44983 , n44986 , n44987 );
xor ( n44989 , n44797 , n44799 );
xor ( n44990 , n44989 , n44801 );
and ( n44991 , n41364 , n39984 );
and ( n44992 , n41379 , n39982 );
nor ( n44993 , n44991 , n44992 );
xnor ( n44994 , n44993 , n39865 );
and ( n44995 , n41844 , n39795 );
and ( n44996 , n41735 , n39793 );
nor ( n44997 , n44995 , n44996 );
xnor ( n44998 , n44997 , n39729 );
and ( n44999 , n44994 , n44998 );
xor ( n45000 , n44335 , n44376 );
xor ( n45001 , n45000 , n44381 );
and ( n45002 , n44998 , n45001 );
and ( n45003 , n44994 , n45001 );
or ( n45004 , n44999 , n45002 , n45003 );
and ( n45005 , n44990 , n45004 );
xor ( n45006 , n44980 , n44982 );
xor ( n45007 , n45006 , n44985 );
and ( n45008 , n45004 , n45007 );
and ( n45009 , n44990 , n45007 );
or ( n45010 , n45005 , n45008 , n45009 );
and ( n45011 , n44988 , n45010 );
xor ( n45012 , n44804 , n44806 );
xor ( n45013 , n45012 , n44809 );
and ( n45014 , n45010 , n45013 );
and ( n45015 , n44988 , n45013 );
or ( n45016 , n45011 , n45014 , n45015 );
and ( n45017 , n44888 , n45016 );
and ( n45018 , n44812 , n45016 );
or ( n45019 , n44889 , n45017 , n45018 );
xor ( n45020 , n44599 , n44650 );
xor ( n45021 , n45020 , n44653 );
and ( n45022 , n45019 , n45021 );
xor ( n45023 , n44693 , n44695 );
xor ( n45024 , n45023 , n44698 );
and ( n45025 , n45021 , n45024 );
and ( n45026 , n45019 , n45024 );
or ( n45027 , n45022 , n45025 , n45026 );
and ( n45028 , n44735 , n45027 );
xor ( n45029 , n44676 , n44678 );
xor ( n45030 , n45029 , n44701 );
and ( n45031 , n45027 , n45030 );
and ( n45032 , n44735 , n45030 );
or ( n45033 , n45028 , n45031 , n45032 );
and ( n45034 , n44733 , n45033 );
xor ( n45035 , n44672 , n44673 );
xor ( n45036 , n45035 , n44704 );
and ( n45037 , n45033 , n45036 );
and ( n45038 , n44733 , n45036 );
or ( n45039 , n45034 , n45037 , n45038 );
xor ( n45040 , n44670 , n44707 );
xor ( n45041 , n45040 , n44710 );
and ( n45042 , n45039 , n45041 );
xor ( n45043 , n44733 , n45033 );
xor ( n45044 , n45043 , n45036 );
and ( n45045 , n44318 , n39258 );
and ( n45046 , n44000 , n39256 );
nor ( n45047 , n45045 , n45046 );
xnor ( n45048 , n45047 , n39215 );
and ( n45049 , n44826 , n39194 );
and ( n45050 , n44347 , n39192 );
nor ( n45051 , n45049 , n45050 );
xnor ( n45052 , n45051 , n39199 );
and ( n45053 , n45048 , n45052 );
xor ( n45054 , n39032 , n39105 );
buf ( n45055 , n45054 );
buf ( n45056 , n45055 );
buf ( n45057 , n45056 );
and ( n45058 , n45057 , n39186 );
and ( n45059 , n45052 , n45058 );
and ( n45060 , n45048 , n45058 );
or ( n45061 , n45053 , n45059 , n45060 );
and ( n45062 , n43679 , n39335 );
and ( n45063 , n43671 , n39333 );
nor ( n45064 , n45062 , n45063 );
xnor ( n45065 , n45064 , n39300 );
and ( n45066 , n45061 , n45065 );
xor ( n45067 , n44817 , n44821 );
xor ( n45068 , n45067 , n44827 );
and ( n45069 , n45065 , n45068 );
and ( n45070 , n45061 , n45068 );
or ( n45071 , n45066 , n45069 , n45070 );
and ( n45072 , n43322 , n39532 );
and ( n45073 , n43142 , n39530 );
nor ( n45074 , n45072 , n45073 );
xnor ( n45075 , n45074 , n39497 );
and ( n45076 , n45071 , n45075 );
and ( n45077 , n43524 , n39384 );
and ( n45078 , n43387 , n39382 );
nor ( n45079 , n45077 , n45078 );
xnor ( n45080 , n45079 , n39367 );
and ( n45081 , n45075 , n45080 );
and ( n45082 , n45071 , n45080 );
or ( n45083 , n45076 , n45081 , n45082 );
and ( n45084 , n43142 , n39532 );
and ( n45085 , n43040 , n39530 );
nor ( n45086 , n45084 , n45085 );
xnor ( n45087 , n45086 , n39497 );
and ( n45088 , n45083 , n45087 );
xor ( n45089 , n44350 , n44354 );
xor ( n45090 , n45089 , n44363 );
and ( n45091 , n45087 , n45090 );
and ( n45092 , n45083 , n45090 );
or ( n45093 , n45088 , n45091 , n45092 );
and ( n45094 , n42525 , n39665 );
and ( n45095 , n41828 , n39663 );
nor ( n45096 , n45094 , n45095 );
xnor ( n45097 , n45096 , n39608 );
and ( n45098 , n45093 , n45097 );
xor ( n45099 , n44366 , n44370 );
xor ( n45100 , n45099 , n44373 );
and ( n45101 , n45097 , n45100 );
and ( n45102 , n45093 , n45100 );
or ( n45103 , n45098 , n45101 , n45102 );
and ( n45104 , n41091 , n40168 );
and ( n45105 , n41106 , n40166 );
nor ( n45106 , n45104 , n45105 );
xnor ( n45107 , n45106 , n40059 );
and ( n45108 , n45103 , n45107 );
xor ( n45109 , n44858 , n44862 );
xor ( n45110 , n45109 , n44865 );
and ( n45111 , n45107 , n45110 );
and ( n45112 , n45103 , n45110 );
or ( n45113 , n45108 , n45111 , n45112 );
and ( n45114 , n40455 , n40928 );
and ( n45115 , n40280 , n40926 );
nor ( n45116 , n45114 , n45115 );
xnor ( n45117 , n45116 , n40688 );
and ( n45118 , n45113 , n45117 );
and ( n45119 , n40698 , n40666 );
and ( n45120 , n40574 , n40664 );
nor ( n45121 , n45119 , n45120 );
xnor ( n45122 , n45121 , n40445 );
and ( n45123 , n45117 , n45122 );
and ( n45124 , n45113 , n45122 );
or ( n45125 , n45118 , n45123 , n45124 );
and ( n45126 , n39848 , n41981 );
and ( n45127 , n39739 , n41979 );
nor ( n45128 , n45126 , n45127 );
xnor ( n45129 , n45128 , n41373 );
and ( n45130 , n45125 , n45129 );
xor ( n45131 , n44878 , n44882 );
xor ( n45132 , n45131 , n44885 );
and ( n45133 , n45129 , n45132 );
and ( n45134 , n45125 , n45132 );
or ( n45135 , n45130 , n45133 , n45134 );
not ( n45136 , n45135 );
xor ( n45137 , n44683 , n44687 );
xor ( n45138 , n45137 , n44690 );
and ( n45139 , n45136 , n45138 );
buf ( n45140 , n45135 );
and ( n45141 , n45139 , n45140 );
xor ( n45142 , n44643 , n44645 );
xor ( n45143 , n45142 , n44647 );
xor ( n45144 , n44812 , n44888 );
xor ( n45145 , n45144 , n45016 );
and ( n45146 , n45143 , n45145 );
xor ( n45147 , n45136 , n45138 );
and ( n45148 , n45145 , n45147 );
and ( n45149 , n45143 , n45147 );
or ( n45150 , n45146 , n45148 , n45149 );
and ( n45151 , n45140 , n45150 );
and ( n45152 , n45139 , n45150 );
or ( n45153 , n45141 , n45151 , n45152 );
xor ( n45154 , n44735 , n45027 );
xor ( n45155 , n45154 , n45030 );
and ( n45156 , n45153 , n45155 );
xor ( n45157 , n45019 , n45021 );
xor ( n45158 , n45157 , n45024 );
and ( n45159 , n44347 , n39258 );
and ( n45160 , n44318 , n39256 );
nor ( n45161 , n45159 , n45160 );
xnor ( n45162 , n45161 , n39215 );
and ( n45163 , n45057 , n39194 );
and ( n45164 , n44826 , n39192 );
nor ( n45165 , n45163 , n45164 );
xnor ( n45166 , n45165 , n39199 );
and ( n45167 , n45162 , n45166 );
xor ( n45168 , n39035 , n39103 );
buf ( n45169 , n45168 );
buf ( n45170 , n45169 );
buf ( n45171 , n45170 );
and ( n45172 , n45171 , n39186 );
and ( n45173 , n45166 , n45172 );
and ( n45174 , n45162 , n45172 );
or ( n45175 , n45167 , n45173 , n45174 );
and ( n45176 , n43820 , n39335 );
and ( n45177 , n43679 , n39333 );
nor ( n45178 , n45176 , n45177 );
xnor ( n45179 , n45178 , n39300 );
and ( n45180 , n45175 , n45179 );
xor ( n45181 , n45048 , n45052 );
xor ( n45182 , n45181 , n45058 );
and ( n45183 , n45179 , n45182 );
and ( n45184 , n45175 , n45182 );
or ( n45185 , n45180 , n45183 , n45184 );
and ( n45186 , n43387 , n39532 );
and ( n45187 , n43322 , n39530 );
nor ( n45188 , n45186 , n45187 );
xnor ( n45189 , n45188 , n39497 );
and ( n45190 , n45185 , n45189 );
xor ( n45191 , n45061 , n45065 );
xor ( n45192 , n45191 , n45068 );
and ( n45193 , n45189 , n45192 );
and ( n45194 , n45185 , n45192 );
or ( n45195 , n45190 , n45193 , n45194 );
buf ( n45196 , n30360 );
not ( n45197 , n45196 );
and ( n45198 , n45195 , n45197 );
xor ( n45199 , n44813 , n44830 );
xor ( n45200 , n45199 , n44835 );
and ( n45201 , n45197 , n45200 );
and ( n45202 , n45195 , n45200 );
or ( n45203 , n45198 , n45201 , n45202 );
and ( n45204 , n42862 , n39665 );
and ( n45205 , n42525 , n39663 );
nor ( n45206 , n45204 , n45205 );
xnor ( n45207 , n45206 , n39608 );
and ( n45208 , n45203 , n45207 );
xor ( n45209 , n44838 , n44842 );
xor ( n45210 , n45209 , n44845 );
and ( n45211 , n45207 , n45210 );
and ( n45212 , n45203 , n45210 );
or ( n45213 , n45208 , n45211 , n45212 );
and ( n45214 , n41735 , n39984 );
and ( n45215 , n41364 , n39982 );
nor ( n45216 , n45214 , n45215 );
xnor ( n45217 , n45216 , n39865 );
and ( n45218 , n45213 , n45217 );
and ( n45219 , n42149 , n39795 );
and ( n45220 , n41844 , n39793 );
nor ( n45221 , n45219 , n45220 );
xnor ( n45222 , n45221 , n39729 );
and ( n45223 , n45217 , n45222 );
and ( n45224 , n45213 , n45222 );
or ( n45225 , n45218 , n45223 , n45224 );
and ( n45226 , n41379 , n40168 );
and ( n45227 , n41091 , n40166 );
nor ( n45228 , n45226 , n45227 );
xnor ( n45229 , n45228 , n40059 );
xor ( n45230 , n45093 , n45097 );
xor ( n45231 , n45230 , n45100 );
and ( n45232 , n45229 , n45231 );
xor ( n45233 , n44848 , n44852 );
xor ( n45234 , n45233 , n44855 );
and ( n45235 , n45231 , n45234 );
and ( n45236 , n45229 , n45234 );
or ( n45237 , n45232 , n45235 , n45236 );
and ( n45238 , n45225 , n45237 );
and ( n45239 , n40910 , n40406 );
and ( n45240 , n40991 , n40404 );
nor ( n45241 , n45239 , n45240 );
xnor ( n45242 , n45241 , n40262 );
and ( n45243 , n45237 , n45242 );
and ( n45244 , n45225 , n45242 );
or ( n45245 , n45238 , n45243 , n45244 );
and ( n45246 , n40272 , n41230 );
and ( n45247 , n40077 , n41228 );
nor ( n45248 , n45246 , n45247 );
xnor ( n45249 , n45248 , n40981 );
and ( n45250 , n45245 , n45249 );
xor ( n45251 , n44868 , n44872 );
xor ( n45252 , n45251 , n44875 );
and ( n45253 , n45249 , n45252 );
and ( n45254 , n45245 , n45252 );
or ( n45255 , n45250 , n45253 , n45254 );
xor ( n45256 , n44988 , n45010 );
xor ( n45257 , n45256 , n45013 );
and ( n45258 , n45255 , n45257 );
xor ( n45259 , n45125 , n45129 );
xor ( n45260 , n45259 , n45132 );
and ( n45261 , n45257 , n45260 );
and ( n45262 , n45255 , n45260 );
or ( n45263 , n45258 , n45261 , n45262 );
and ( n45264 , n40574 , n40928 );
and ( n45265 , n40455 , n40926 );
nor ( n45266 , n45264 , n45265 );
xnor ( n45267 , n45266 , n40688 );
and ( n45268 , n40962 , n40666 );
and ( n45269 , n40698 , n40664 );
nor ( n45270 , n45268 , n45269 );
xnor ( n45271 , n45270 , n40445 );
and ( n45272 , n45267 , n45271 );
xor ( n45273 , n44994 , n44998 );
xor ( n45274 , n45273 , n45001 );
and ( n45275 , n45271 , n45274 );
and ( n45276 , n45267 , n45274 );
or ( n45277 , n45272 , n45275 , n45276 );
and ( n45278 , n40069 , n41522 );
and ( n45279 , n39935 , n41520 );
nor ( n45280 , n45278 , n45279 );
xnor ( n45281 , n45280 , n41100 );
and ( n45282 , n45277 , n45281 );
xor ( n45283 , n45113 , n45117 );
xor ( n45284 , n45283 , n45122 );
and ( n45285 , n45281 , n45284 );
and ( n45286 , n45277 , n45284 );
or ( n45287 , n45282 , n45285 , n45286 );
and ( n45288 , n42149 , n39984 );
and ( n45289 , n41844 , n39982 );
nor ( n45290 , n45288 , n45289 );
xnor ( n45291 , n45290 , n39865 );
and ( n45292 , n42525 , n39795 );
and ( n45293 , n41828 , n39793 );
nor ( n45294 , n45292 , n45293 );
xnor ( n45295 , n45294 , n39729 );
and ( n45296 , n45291 , n45295 );
xnor ( n45297 , n44919 , n44923 );
and ( n45298 , n45295 , n45297 );
and ( n45299 , n45291 , n45297 );
or ( n45300 , n45296 , n45298 , n45299 );
and ( n45301 , n40077 , n42079 );
and ( n45302 , n40069 , n42076 );
nor ( n45303 , n45301 , n45302 );
xnor ( n45304 , n45303 , n41370 );
and ( n45305 , n40280 , n41981 );
and ( n45306 , n40272 , n41979 );
nor ( n45307 , n45305 , n45306 );
xnor ( n45308 , n45307 , n41373 );
and ( n45309 , n45304 , n45308 );
and ( n45310 , n40574 , n41522 );
and ( n45311 , n40455 , n41520 );
nor ( n45312 , n45310 , n45311 );
xnor ( n45313 , n45312 , n41100 );
and ( n45314 , n45308 , n45313 );
and ( n45315 , n45304 , n45313 );
or ( n45316 , n45309 , n45314 , n45315 );
and ( n45317 , n40962 , n41230 );
and ( n45318 , n40698 , n41228 );
nor ( n45319 , n45317 , n45318 );
xnor ( n45320 , n45319 , n40981 );
and ( n45321 , n40910 , n40928 );
and ( n45322 , n40991 , n40926 );
nor ( n45323 , n45321 , n45322 );
xnor ( n45324 , n45323 , n40688 );
and ( n45325 , n45320 , n45324 );
and ( n45326 , n41091 , n40666 );
and ( n45327 , n41106 , n40664 );
nor ( n45328 , n45326 , n45327 );
xnor ( n45329 , n45328 , n40445 );
and ( n45330 , n45324 , n45329 );
and ( n45331 , n45320 , n45329 );
or ( n45332 , n45325 , n45330 , n45331 );
and ( n45333 , n45316 , n45332 );
and ( n45334 , n41364 , n40406 );
and ( n45335 , n41379 , n40404 );
nor ( n45336 , n45334 , n45335 );
xnor ( n45337 , n45336 , n40262 );
and ( n45338 , n41844 , n40168 );
and ( n45339 , n41735 , n40166 );
nor ( n45340 , n45338 , n45339 );
xnor ( n45341 , n45340 , n40059 );
and ( n45342 , n45337 , n45341 );
and ( n45343 , n41828 , n39984 );
and ( n45344 , n42149 , n39982 );
nor ( n45345 , n45343 , n45344 );
xnor ( n45346 , n45345 , n39865 );
and ( n45347 , n45341 , n45346 );
and ( n45348 , n45337 , n45346 );
or ( n45349 , n45342 , n45347 , n45348 );
and ( n45350 , n45332 , n45349 );
and ( n45351 , n45316 , n45349 );
or ( n45352 , n45333 , n45350 , n45351 );
and ( n45353 , n45300 , n45352 );
and ( n45354 , n42862 , n39795 );
and ( n45355 , n42525 , n39793 );
nor ( n45356 , n45354 , n45355 );
xnor ( n45357 , n45356 , n39729 );
and ( n45358 , n43549 , n39384 );
and ( n45359 , n43524 , n39382 );
nor ( n45360 , n45358 , n45359 );
xnor ( n45361 , n45360 , n39367 );
and ( n45362 , n45357 , n45361 );
buf ( n45363 , n30361 );
not ( n45364 , n45363 );
and ( n45365 , n45361 , n45364 );
and ( n45366 , n45357 , n45364 );
or ( n45367 , n45362 , n45365 , n45366 );
xor ( n45368 , n44929 , n44933 );
xor ( n45369 , n45368 , n44938 );
and ( n45370 , n45367 , n45369 );
xor ( n45371 , n44948 , n44952 );
xor ( n45372 , n45371 , n44957 );
and ( n45373 , n45369 , n45372 );
and ( n45374 , n45367 , n45372 );
or ( n45375 , n45370 , n45373 , n45374 );
and ( n45376 , n45352 , n45375 );
and ( n45377 , n45300 , n45375 );
or ( n45378 , n45353 , n45376 , n45377 );
xor ( n45379 , n44905 , n44907 );
xor ( n45380 , n45379 , n44910 );
and ( n45381 , n45378 , n45380 );
xor ( n45382 , n44944 , n44968 );
xor ( n45383 , n45382 , n44971 );
and ( n45384 , n45380 , n45383 );
and ( n45385 , n45378 , n45383 );
or ( n45386 , n45381 , n45384 , n45385 );
xor ( n45387 , n44913 , n44974 );
xor ( n45388 , n45387 , n44977 );
and ( n45389 , n45386 , n45388 );
xor ( n45390 , n44915 , n44924 );
xor ( n45391 , n45390 , n44941 );
xor ( n45392 , n44960 , n44962 );
xor ( n45393 , n45392 , n44965 );
and ( n45394 , n45391 , n45393 );
and ( n45395 , n40272 , n42079 );
and ( n45396 , n40077 , n42076 );
nor ( n45397 , n45395 , n45396 );
xnor ( n45398 , n45397 , n41370 );
and ( n45399 , n40455 , n41981 );
and ( n45400 , n40280 , n41979 );
nor ( n45401 , n45399 , n45400 );
xnor ( n45402 , n45401 , n41373 );
and ( n45403 , n45398 , n45402 );
and ( n45404 , n40698 , n41522 );
and ( n45405 , n40574 , n41520 );
nor ( n45406 , n45404 , n45405 );
xnor ( n45407 , n45406 , n41100 );
and ( n45408 , n45402 , n45407 );
and ( n45409 , n45398 , n45407 );
or ( n45410 , n45403 , n45408 , n45409 );
and ( n45411 , n40991 , n41230 );
and ( n45412 , n40962 , n41228 );
nor ( n45413 , n45411 , n45412 );
xnor ( n45414 , n45413 , n40981 );
and ( n45415 , n41106 , n40928 );
and ( n45416 , n40910 , n40926 );
nor ( n45417 , n45415 , n45416 );
xnor ( n45418 , n45417 , n40688 );
and ( n45419 , n45414 , n45418 );
and ( n45420 , n41379 , n40666 );
and ( n45421 , n41091 , n40664 );
nor ( n45422 , n45420 , n45421 );
xnor ( n45423 , n45422 , n40445 );
and ( n45424 , n45418 , n45423 );
and ( n45425 , n45414 , n45423 );
or ( n45426 , n45419 , n45424 , n45425 );
and ( n45427 , n45410 , n45426 );
and ( n45428 , n41735 , n40406 );
and ( n45429 , n41364 , n40404 );
nor ( n45430 , n45428 , n45429 );
xnor ( n45431 , n45430 , n40262 );
and ( n45432 , n42149 , n40168 );
and ( n45433 , n41844 , n40166 );
nor ( n45434 , n45432 , n45433 );
xnor ( n45435 , n45434 , n40059 );
and ( n45436 , n45431 , n45435 );
and ( n45437 , n42525 , n39984 );
and ( n45438 , n41828 , n39982 );
nor ( n45439 , n45437 , n45438 );
xnor ( n45440 , n45439 , n39865 );
and ( n45441 , n45435 , n45440 );
and ( n45442 , n45431 , n45440 );
or ( n45443 , n45436 , n45441 , n45442 );
and ( n45444 , n45426 , n45443 );
and ( n45445 , n45410 , n45443 );
or ( n45446 , n45427 , n45444 , n45445 );
and ( n45447 , n43040 , n39795 );
and ( n45448 , n42862 , n39793 );
nor ( n45449 , n45447 , n45448 );
xnor ( n45450 , n45449 , n39729 );
and ( n45451 , n43322 , n39665 );
and ( n45452 , n43142 , n39663 );
nor ( n45453 , n45451 , n45452 );
xnor ( n45454 , n45453 , n39608 );
and ( n45455 , n45450 , n45454 );
and ( n45456 , n43671 , n39384 );
and ( n45457 , n43549 , n39382 );
nor ( n45458 , n45456 , n45457 );
xnor ( n45459 , n45458 , n39367 );
and ( n45460 , n45454 , n45459 );
and ( n45461 , n45450 , n45459 );
or ( n45462 , n45455 , n45460 , n45461 );
xor ( n45463 , n45304 , n45308 );
xor ( n45464 , n45463 , n45313 );
and ( n45465 , n45462 , n45464 );
xor ( n45466 , n45320 , n45324 );
xor ( n45467 , n45466 , n45329 );
and ( n45468 , n45464 , n45467 );
and ( n45469 , n45462 , n45467 );
or ( n45470 , n45465 , n45468 , n45469 );
and ( n45471 , n45446 , n45470 );
xor ( n45472 , n45291 , n45295 );
xor ( n45473 , n45472 , n45297 );
and ( n45474 , n45470 , n45473 );
and ( n45475 , n45446 , n45473 );
or ( n45476 , n45471 , n45474 , n45475 );
and ( n45477 , n45393 , n45476 );
and ( n45478 , n45391 , n45476 );
or ( n45479 , n45394 , n45477 , n45478 );
xor ( n45480 , n45378 , n45380 );
xor ( n45481 , n45480 , n45383 );
and ( n45482 , n45479 , n45481 );
and ( n45483 , n41828 , n39795 );
and ( n45484 , n42149 , n39793 );
nor ( n45485 , n45483 , n45484 );
xnor ( n45486 , n45485 , n39729 );
xor ( n45487 , n45083 , n45087 );
xor ( n45488 , n45487 , n45090 );
and ( n45489 , n45486 , n45488 );
and ( n45490 , n45481 , n45489 );
and ( n45491 , n45479 , n45489 );
or ( n45492 , n45482 , n45490 , n45491 );
and ( n45493 , n45388 , n45492 );
and ( n45494 , n45386 , n45492 );
or ( n45495 , n45389 , n45493 , n45494 );
xor ( n45496 , n44990 , n45004 );
xor ( n45497 , n45496 , n45007 );
and ( n45498 , n45495 , n45497 );
xor ( n45499 , n45245 , n45249 );
xor ( n45500 , n45499 , n45252 );
and ( n45501 , n45497 , n45500 );
and ( n45502 , n45495 , n45500 );
or ( n45503 , n45498 , n45501 , n45502 );
and ( n45504 , n45287 , n45503 );
and ( n45505 , n40077 , n41522 );
and ( n45506 , n40069 , n41520 );
nor ( n45507 , n45505 , n45506 );
xnor ( n45508 , n45507 , n41100 );
and ( n45509 , n40280 , n41230 );
and ( n45510 , n40272 , n41228 );
nor ( n45511 , n45509 , n45510 );
xnor ( n45512 , n45511 , n40981 );
and ( n45513 , n45508 , n45512 );
xor ( n45514 , n45103 , n45107 );
xor ( n45515 , n45514 , n45110 );
and ( n45516 , n45512 , n45515 );
and ( n45517 , n45508 , n45515 );
or ( n45518 , n45513 , n45516 , n45517 );
xor ( n45519 , n45225 , n45237 );
xor ( n45520 , n45519 , n45242 );
xor ( n45521 , n45267 , n45271 );
xor ( n45522 , n45521 , n45274 );
and ( n45523 , n45520 , n45522 );
xor ( n45524 , n45300 , n45352 );
xor ( n45525 , n45524 , n45375 );
xor ( n45526 , n45316 , n45332 );
xor ( n45527 , n45526 , n45349 );
xor ( n45528 , n45367 , n45369 );
xor ( n45529 , n45528 , n45372 );
and ( n45530 , n45527 , n45529 );
xor ( n45531 , n45071 , n45075 );
xor ( n45532 , n45531 , n45080 );
and ( n45533 , n45529 , n45532 );
and ( n45534 , n45527 , n45532 );
or ( n45535 , n45530 , n45533 , n45534 );
and ( n45536 , n45525 , n45535 );
xor ( n45537 , n45337 , n45341 );
xor ( n45538 , n45537 , n45346 );
xor ( n45539 , n45357 , n45361 );
xor ( n45540 , n45539 , n45364 );
and ( n45541 , n45538 , n45540 );
buf ( n45542 , n30362 );
not ( n45543 , n45542 );
and ( n45544 , n41091 , n40928 );
and ( n45545 , n41106 , n40926 );
nor ( n45546 , n45544 , n45545 );
xnor ( n45547 , n45546 , n40688 );
and ( n45548 , n41364 , n40666 );
and ( n45549 , n41379 , n40664 );
nor ( n45550 , n45548 , n45549 );
xnor ( n45551 , n45550 , n40445 );
or ( n45552 , n45547 , n45551 );
and ( n45553 , n45543 , n45552 );
and ( n45554 , n40280 , n42079 );
and ( n45555 , n40272 , n42076 );
nor ( n45556 , n45554 , n45555 );
xnor ( n45557 , n45556 , n41370 );
and ( n45558 , n40574 , n41981 );
and ( n45559 , n40455 , n41979 );
nor ( n45560 , n45558 , n45559 );
xnor ( n45561 , n45560 , n41373 );
and ( n45562 , n45557 , n45561 );
and ( n45563 , n40962 , n41522 );
and ( n45564 , n40698 , n41520 );
nor ( n45565 , n45563 , n45564 );
xnor ( n45566 , n45565 , n41100 );
and ( n45567 , n45561 , n45566 );
and ( n45568 , n45557 , n45566 );
or ( n45569 , n45562 , n45567 , n45568 );
and ( n45570 , n45552 , n45569 );
and ( n45571 , n45543 , n45569 );
or ( n45572 , n45553 , n45570 , n45571 );
and ( n45573 , n45540 , n45572 );
and ( n45574 , n45538 , n45572 );
or ( n45575 , n45541 , n45573 , n45574 );
and ( n45576 , n40910 , n41230 );
and ( n45577 , n40991 , n41228 );
nor ( n45578 , n45576 , n45577 );
xnor ( n45579 , n45578 , n40981 );
and ( n45580 , n41844 , n40406 );
and ( n45581 , n41735 , n40404 );
nor ( n45582 , n45580 , n45581 );
xnor ( n45583 , n45582 , n40262 );
and ( n45584 , n45579 , n45583 );
and ( n45585 , n41828 , n40168 );
and ( n45586 , n42149 , n40166 );
nor ( n45587 , n45585 , n45586 );
xnor ( n45588 , n45587 , n40059 );
and ( n45589 , n45583 , n45588 );
and ( n45590 , n45579 , n45588 );
or ( n45591 , n45584 , n45589 , n45590 );
and ( n45592 , n42862 , n39984 );
and ( n45593 , n42525 , n39982 );
nor ( n45594 , n45592 , n45593 );
xnor ( n45595 , n45594 , n39865 );
and ( n45596 , n43142 , n39795 );
and ( n45597 , n43040 , n39793 );
nor ( n45598 , n45596 , n45597 );
xnor ( n45599 , n45598 , n39729 );
and ( n45600 , n45595 , n45599 );
and ( n45601 , n43387 , n39665 );
and ( n45602 , n43322 , n39663 );
nor ( n45603 , n45601 , n45602 );
xnor ( n45604 , n45603 , n39608 );
and ( n45605 , n45599 , n45604 );
and ( n45606 , n45595 , n45604 );
or ( n45607 , n45600 , n45605 , n45606 );
and ( n45608 , n45591 , n45607 );
and ( n45609 , n43549 , n39532 );
and ( n45610 , n43524 , n39530 );
nor ( n45611 , n45609 , n45610 );
xnor ( n45612 , n45611 , n39497 );
and ( n45613 , n43679 , n39384 );
and ( n45614 , n43671 , n39382 );
nor ( n45615 , n45613 , n45614 );
xnor ( n45616 , n45615 , n39367 );
and ( n45617 , n45612 , n45616 );
and ( n45618 , n44000 , n39335 );
and ( n45619 , n43820 , n39333 );
nor ( n45620 , n45618 , n45619 );
xnor ( n45621 , n45620 , n39300 );
and ( n45622 , n45616 , n45621 );
and ( n45623 , n45612 , n45621 );
or ( n45624 , n45617 , n45622 , n45623 );
and ( n45625 , n45607 , n45624 );
and ( n45626 , n45591 , n45624 );
or ( n45627 , n45608 , n45625 , n45626 );
xor ( n45628 , n45398 , n45402 );
xor ( n45629 , n45628 , n45407 );
xor ( n45630 , n45414 , n45418 );
xor ( n45631 , n45630 , n45423 );
and ( n45632 , n45629 , n45631 );
xor ( n45633 , n45431 , n45435 );
xor ( n45634 , n45633 , n45440 );
and ( n45635 , n45631 , n45634 );
and ( n45636 , n45629 , n45634 );
or ( n45637 , n45632 , n45635 , n45636 );
and ( n45638 , n45627 , n45637 );
xor ( n45639 , n45410 , n45426 );
xor ( n45640 , n45639 , n45443 );
and ( n45641 , n45637 , n45640 );
and ( n45642 , n45627 , n45640 );
or ( n45643 , n45638 , n45641 , n45642 );
and ( n45644 , n45575 , n45643 );
xor ( n45645 , n45446 , n45470 );
xor ( n45646 , n45645 , n45473 );
and ( n45647 , n45643 , n45646 );
and ( n45648 , n45575 , n45646 );
or ( n45649 , n45644 , n45647 , n45648 );
and ( n45650 , n45535 , n45649 );
and ( n45651 , n45525 , n45649 );
or ( n45652 , n45536 , n45650 , n45651 );
xor ( n45653 , n45213 , n45217 );
xor ( n45654 , n45653 , n45222 );
and ( n45655 , n45652 , n45654 );
xor ( n45656 , n45229 , n45231 );
xor ( n45657 , n45656 , n45234 );
and ( n45658 , n45654 , n45657 );
and ( n45659 , n45652 , n45657 );
or ( n45660 , n45655 , n45658 , n45659 );
and ( n45661 , n45522 , n45660 );
and ( n45662 , n45520 , n45660 );
or ( n45663 , n45523 , n45661 , n45662 );
and ( n45664 , n45518 , n45663 );
xor ( n45665 , n45277 , n45281 );
xor ( n45666 , n45665 , n45284 );
and ( n45667 , n45663 , n45666 );
and ( n45668 , n45518 , n45666 );
or ( n45669 , n45664 , n45667 , n45668 );
and ( n45670 , n45503 , n45669 );
and ( n45671 , n45287 , n45669 );
or ( n45672 , n45504 , n45670 , n45671 );
and ( n45673 , n45263 , n45672 );
xor ( n45674 , n45143 , n45145 );
xor ( n45675 , n45674 , n45147 );
and ( n45676 , n45672 , n45675 );
and ( n45677 , n45263 , n45675 );
or ( n45678 , n45673 , n45676 , n45677 );
and ( n45679 , n45158 , n45678 );
xor ( n45680 , n45139 , n45140 );
xor ( n45681 , n45680 , n45150 );
and ( n45682 , n45678 , n45681 );
and ( n45683 , n45158 , n45681 );
or ( n45684 , n45679 , n45682 , n45683 );
and ( n45685 , n45155 , n45684 );
and ( n45686 , n45153 , n45684 );
or ( n45687 , n45156 , n45685 , n45686 );
or ( n45688 , n45044 , n45687 );
and ( n45689 , n45041 , n45688 );
and ( n45690 , n45039 , n45688 );
or ( n45691 , n45042 , n45689 , n45690 );
and ( n45692 , n44731 , n45691 );
xor ( n45693 , n44731 , n45691 );
xor ( n45694 , n45039 , n45041 );
xor ( n45695 , n45694 , n45688 );
not ( n45696 , n45695 );
xnor ( n45697 , n45044 , n45687 );
xor ( n45698 , n45153 , n45155 );
xor ( n45699 , n45698 , n45684 );
xor ( n45700 , n45255 , n45257 );
xor ( n45701 , n45700 , n45260 );
xor ( n45702 , n45391 , n45393 );
xor ( n45703 , n45702 , n45476 );
xor ( n45704 , n45203 , n45207 );
xor ( n45705 , n45704 , n45210 );
and ( n45706 , n45703 , n45705 );
xor ( n45707 , n45486 , n45488 );
and ( n45708 , n45705 , n45707 );
and ( n45709 , n45703 , n45707 );
or ( n45710 , n45706 , n45708 , n45709 );
and ( n45711 , n43040 , n39665 );
and ( n45712 , n42862 , n39663 );
nor ( n45713 , n45711 , n45712 );
xnor ( n45714 , n45713 , n39608 );
xor ( n45715 , n45195 , n45197 );
xor ( n45716 , n45715 , n45200 );
and ( n45717 , n45714 , n45716 );
and ( n45718 , n43142 , n39665 );
and ( n45719 , n43040 , n39663 );
nor ( n45720 , n45718 , n45719 );
xnor ( n45721 , n45720 , n39608 );
xor ( n45722 , n45185 , n45189 );
xor ( n45723 , n45722 , n45192 );
or ( n45724 , n45721 , n45723 );
xor ( n45725 , n45462 , n45464 );
xor ( n45726 , n45725 , n45467 );
and ( n45727 , n43524 , n39532 );
and ( n45728 , n43387 , n39530 );
nor ( n45729 , n45727 , n45728 );
xnor ( n45730 , n45729 , n39497 );
xor ( n45731 , n45175 , n45179 );
xor ( n45732 , n45731 , n45182 );
and ( n45733 , n45730 , n45732 );
and ( n45734 , n45726 , n45733 );
xor ( n45735 , n45450 , n45454 );
xor ( n45736 , n45735 , n45459 );
buf ( n45737 , n30363 );
not ( n45738 , n45737 );
xor ( n45739 , n45162 , n45166 );
xor ( n45740 , n45739 , n45172 );
and ( n45741 , n45738 , n45740 );
xnor ( n45742 , n45547 , n45551 );
and ( n45743 , n45740 , n45742 );
and ( n45744 , n45738 , n45742 );
or ( n45745 , n45741 , n45743 , n45744 );
and ( n45746 , n45736 , n45745 );
and ( n45747 , n45171 , n39194 );
and ( n45748 , n45057 , n39192 );
nor ( n45749 , n45747 , n45748 );
xnor ( n45750 , n45749 , n39199 );
xor ( n45751 , n39036 , n39102 );
buf ( n45752 , n45751 );
buf ( n45753 , n45752 );
buf ( n45754 , n45753 );
and ( n45755 , n45754 , n39186 );
and ( n45756 , n45750 , n45755 );
and ( n45757 , n40455 , n42079 );
and ( n45758 , n40280 , n42076 );
nor ( n45759 , n45757 , n45758 );
xnor ( n45760 , n45759 , n41370 );
and ( n45761 , n40698 , n41981 );
and ( n45762 , n40574 , n41979 );
nor ( n45763 , n45761 , n45762 );
xnor ( n45764 , n45763 , n41373 );
and ( n45765 , n45760 , n45764 );
and ( n45766 , n40991 , n41522 );
and ( n45767 , n40962 , n41520 );
nor ( n45768 , n45766 , n45767 );
xnor ( n45769 , n45768 , n41100 );
and ( n45770 , n45764 , n45769 );
and ( n45771 , n45760 , n45769 );
or ( n45772 , n45765 , n45770 , n45771 );
and ( n45773 , n45756 , n45772 );
and ( n45774 , n41106 , n41230 );
and ( n45775 , n40910 , n41228 );
nor ( n45776 , n45774 , n45775 );
xnor ( n45777 , n45776 , n40981 );
and ( n45778 , n41379 , n40928 );
and ( n45779 , n41091 , n40926 );
nor ( n45780 , n45778 , n45779 );
xnor ( n45781 , n45780 , n40688 );
and ( n45782 , n45777 , n45781 );
and ( n45783 , n41735 , n40666 );
and ( n45784 , n41364 , n40664 );
nor ( n45785 , n45783 , n45784 );
xnor ( n45786 , n45785 , n40445 );
and ( n45787 , n45781 , n45786 );
and ( n45788 , n45777 , n45786 );
or ( n45789 , n45782 , n45787 , n45788 );
and ( n45790 , n45772 , n45789 );
and ( n45791 , n45756 , n45789 );
or ( n45792 , n45773 , n45790 , n45791 );
and ( n45793 , n45745 , n45792 );
and ( n45794 , n45736 , n45792 );
or ( n45795 , n45746 , n45793 , n45794 );
and ( n45796 , n45733 , n45795 );
and ( n45797 , n45726 , n45795 );
or ( n45798 , n45734 , n45796 , n45797 );
and ( n45799 , n45724 , n45798 );
and ( n45800 , n42149 , n40406 );
and ( n45801 , n41844 , n40404 );
nor ( n45802 , n45800 , n45801 );
xnor ( n45803 , n45802 , n40262 );
and ( n45804 , n42525 , n40168 );
and ( n45805 , n41828 , n40166 );
nor ( n45806 , n45804 , n45805 );
xnor ( n45807 , n45806 , n40059 );
and ( n45808 , n45803 , n45807 );
and ( n45809 , n43040 , n39984 );
and ( n45810 , n42862 , n39982 );
nor ( n45811 , n45809 , n45810 );
xnor ( n45812 , n45811 , n39865 );
and ( n45813 , n45807 , n45812 );
and ( n45814 , n45803 , n45812 );
or ( n45815 , n45808 , n45813 , n45814 );
and ( n45816 , n43322 , n39795 );
and ( n45817 , n43142 , n39793 );
nor ( n45818 , n45816 , n45817 );
xnor ( n45819 , n45818 , n39729 );
and ( n45820 , n43524 , n39665 );
and ( n45821 , n43387 , n39663 );
nor ( n45822 , n45820 , n45821 );
xnor ( n45823 , n45822 , n39608 );
and ( n45824 , n45819 , n45823 );
and ( n45825 , n43671 , n39532 );
and ( n45826 , n43549 , n39530 );
nor ( n45827 , n45825 , n45826 );
xnor ( n45828 , n45827 , n39497 );
and ( n45829 , n45823 , n45828 );
and ( n45830 , n45819 , n45828 );
or ( n45831 , n45824 , n45829 , n45830 );
and ( n45832 , n45815 , n45831 );
and ( n45833 , n43820 , n39384 );
and ( n45834 , n43679 , n39382 );
nor ( n45835 , n45833 , n45834 );
xnor ( n45836 , n45835 , n39367 );
and ( n45837 , n44318 , n39335 );
and ( n45838 , n44000 , n39333 );
nor ( n45839 , n45837 , n45838 );
xnor ( n45840 , n45839 , n39300 );
and ( n45841 , n45836 , n45840 );
and ( n45842 , n44826 , n39258 );
and ( n45843 , n44347 , n39256 );
nor ( n45844 , n45842 , n45843 );
xnor ( n45845 , n45844 , n39215 );
and ( n45846 , n45840 , n45845 );
and ( n45847 , n45836 , n45845 );
or ( n45848 , n45841 , n45846 , n45847 );
and ( n45849 , n45831 , n45848 );
and ( n45850 , n45815 , n45848 );
or ( n45851 , n45832 , n45849 , n45850 );
xor ( n45852 , n45557 , n45561 );
xor ( n45853 , n45852 , n45566 );
xor ( n45854 , n45579 , n45583 );
xor ( n45855 , n45854 , n45588 );
and ( n45856 , n45853 , n45855 );
xor ( n45857 , n45595 , n45599 );
xor ( n45858 , n45857 , n45604 );
and ( n45859 , n45855 , n45858 );
and ( n45860 , n45853 , n45858 );
or ( n45861 , n45856 , n45859 , n45860 );
and ( n45862 , n45851 , n45861 );
xor ( n45863 , n45543 , n45552 );
xor ( n45864 , n45863 , n45569 );
and ( n45865 , n45861 , n45864 );
and ( n45866 , n45851 , n45864 );
or ( n45867 , n45862 , n45865 , n45866 );
xor ( n45868 , n45538 , n45540 );
xor ( n45869 , n45868 , n45572 );
and ( n45870 , n45867 , n45869 );
xor ( n45871 , n45627 , n45637 );
xor ( n45872 , n45871 , n45640 );
and ( n45873 , n45869 , n45872 );
and ( n45874 , n45867 , n45872 );
or ( n45875 , n45870 , n45873 , n45874 );
and ( n45876 , n45798 , n45875 );
and ( n45877 , n45724 , n45875 );
or ( n45878 , n45799 , n45876 , n45877 );
and ( n45879 , n45717 , n45878 );
xor ( n45880 , n45525 , n45535 );
xor ( n45881 , n45880 , n45649 );
and ( n45882 , n45878 , n45881 );
and ( n45883 , n45717 , n45881 );
or ( n45884 , n45879 , n45882 , n45883 );
and ( n45885 , n45710 , n45884 );
xor ( n45886 , n45479 , n45481 );
xor ( n45887 , n45886 , n45489 );
and ( n45888 , n45884 , n45887 );
and ( n45889 , n45710 , n45887 );
or ( n45890 , n45885 , n45888 , n45889 );
xor ( n45891 , n45386 , n45388 );
xor ( n45892 , n45891 , n45492 );
and ( n45893 , n45890 , n45892 );
xor ( n45894 , n45508 , n45512 );
xor ( n45895 , n45894 , n45515 );
and ( n45896 , n45892 , n45895 );
and ( n45897 , n45890 , n45895 );
or ( n45898 , n45893 , n45896 , n45897 );
xor ( n45899 , n45495 , n45497 );
xor ( n45900 , n45899 , n45500 );
and ( n45901 , n45898 , n45900 );
xor ( n45902 , n45527 , n45529 );
xor ( n45903 , n45902 , n45532 );
xor ( n45904 , n45575 , n45643 );
xor ( n45905 , n45904 , n45646 );
and ( n45906 , n45903 , n45905 );
xor ( n45907 , n45714 , n45716 );
and ( n45908 , n45905 , n45907 );
and ( n45909 , n45903 , n45907 );
or ( n45910 , n45906 , n45908 , n45909 );
xor ( n45911 , n45703 , n45705 );
xor ( n45912 , n45911 , n45707 );
and ( n45913 , n45910 , n45912 );
xor ( n45914 , n45717 , n45878 );
xor ( n45915 , n45914 , n45881 );
and ( n45916 , n45912 , n45915 );
and ( n45917 , n45910 , n45915 );
or ( n45918 , n45913 , n45916 , n45917 );
xor ( n45919 , n45652 , n45654 );
xor ( n45920 , n45919 , n45657 );
and ( n45921 , n45918 , n45920 );
xor ( n45922 , n45710 , n45884 );
xor ( n45923 , n45922 , n45887 );
and ( n45924 , n45920 , n45923 );
and ( n45925 , n45918 , n45923 );
or ( n45926 , n45921 , n45924 , n45925 );
xor ( n45927 , n45520 , n45522 );
xor ( n45928 , n45927 , n45660 );
and ( n45929 , n45926 , n45928 );
xor ( n45930 , n45890 , n45892 );
xor ( n45931 , n45930 , n45895 );
and ( n45932 , n45928 , n45931 );
and ( n45933 , n45926 , n45931 );
or ( n45934 , n45929 , n45932 , n45933 );
and ( n45935 , n45900 , n45934 );
and ( n45936 , n45898 , n45934 );
or ( n45937 , n45901 , n45935 , n45936 );
and ( n45938 , n45701 , n45937 );
xor ( n45939 , n45287 , n45503 );
xor ( n45940 , n45939 , n45669 );
and ( n45941 , n45937 , n45940 );
and ( n45942 , n45701 , n45940 );
or ( n45943 , n45938 , n45941 , n45942 );
xor ( n45944 , n45263 , n45672 );
xor ( n45945 , n45944 , n45675 );
or ( n45946 , n45943 , n45945 );
xor ( n45947 , n45158 , n45678 );
xor ( n45948 , n45947 , n45681 );
and ( n45949 , n45946 , n45948 );
xor ( n45950 , n45946 , n45948 );
xnor ( n45951 , n45943 , n45945 );
xor ( n45952 , n45518 , n45663 );
xor ( n45953 , n45952 , n45666 );
xor ( n45954 , n45918 , n45920 );
xor ( n45955 , n45954 , n45923 );
xnor ( n45956 , n45721 , n45723 );
xor ( n45957 , n45591 , n45607 );
xor ( n45958 , n45957 , n45624 );
xor ( n45959 , n45629 , n45631 );
xor ( n45960 , n45959 , n45634 );
and ( n45961 , n45958 , n45960 );
xor ( n45962 , n45730 , n45732 );
and ( n45963 , n45960 , n45962 );
and ( n45964 , n45958 , n45962 );
or ( n45965 , n45961 , n45963 , n45964 );
and ( n45966 , n45956 , n45965 );
xor ( n45967 , n45612 , n45616 );
xor ( n45968 , n45967 , n45621 );
buf ( n45969 , n30364 );
not ( n45970 , n45969 );
xor ( n45971 , n45750 , n45755 );
and ( n45972 , n45970 , n45971 );
and ( n45973 , n41091 , n41230 );
and ( n45974 , n41106 , n41228 );
nor ( n45975 , n45973 , n45974 );
xnor ( n45976 , n45975 , n40981 );
and ( n45977 , n41364 , n40928 );
and ( n45978 , n41379 , n40926 );
nor ( n45979 , n45977 , n45978 );
xnor ( n45980 , n45979 , n40688 );
or ( n45981 , n45976 , n45980 );
and ( n45982 , n45971 , n45981 );
and ( n45983 , n45970 , n45981 );
or ( n45984 , n45972 , n45982 , n45983 );
and ( n45985 , n45968 , n45984 );
and ( n45986 , n40574 , n42079 );
and ( n45987 , n40455 , n42076 );
nor ( n45988 , n45986 , n45987 );
xnor ( n45989 , n45988 , n41370 );
and ( n45990 , n40962 , n41981 );
and ( n45991 , n40698 , n41979 );
nor ( n45992 , n45990 , n45991 );
xnor ( n45993 , n45992 , n41373 );
and ( n45994 , n45989 , n45993 );
and ( n45995 , n40910 , n41522 );
and ( n45996 , n40991 , n41520 );
nor ( n45997 , n45995 , n45996 );
xnor ( n45998 , n45997 , n41100 );
and ( n45999 , n45993 , n45998 );
and ( n46000 , n45989 , n45998 );
or ( n46001 , n45994 , n45999 , n46000 );
and ( n46002 , n41844 , n40666 );
and ( n46003 , n41735 , n40664 );
nor ( n46004 , n46002 , n46003 );
xnor ( n46005 , n46004 , n40445 );
and ( n46006 , n41828 , n40406 );
and ( n46007 , n42149 , n40404 );
nor ( n46008 , n46006 , n46007 );
xnor ( n46009 , n46008 , n40262 );
and ( n46010 , n46005 , n46009 );
and ( n46011 , n42862 , n40168 );
and ( n46012 , n42525 , n40166 );
nor ( n46013 , n46011 , n46012 );
xnor ( n46014 , n46013 , n40059 );
and ( n46015 , n46009 , n46014 );
and ( n46016 , n46005 , n46014 );
or ( n46017 , n46010 , n46015 , n46016 );
and ( n46018 , n46001 , n46017 );
and ( n46019 , n43142 , n39984 );
and ( n46020 , n43040 , n39982 );
nor ( n46021 , n46019 , n46020 );
xnor ( n46022 , n46021 , n39865 );
and ( n46023 , n43387 , n39795 );
and ( n46024 , n43322 , n39793 );
nor ( n46025 , n46023 , n46024 );
xnor ( n46026 , n46025 , n39729 );
and ( n46027 , n46022 , n46026 );
and ( n46028 , n43549 , n39665 );
and ( n46029 , n43524 , n39663 );
nor ( n46030 , n46028 , n46029 );
xnor ( n46031 , n46030 , n39608 );
and ( n46032 , n46026 , n46031 );
and ( n46033 , n46022 , n46031 );
or ( n46034 , n46027 , n46032 , n46033 );
and ( n46035 , n46017 , n46034 );
and ( n46036 , n46001 , n46034 );
or ( n46037 , n46018 , n46035 , n46036 );
and ( n46038 , n45984 , n46037 );
and ( n46039 , n45968 , n46037 );
or ( n46040 , n45985 , n46038 , n46039 );
and ( n46041 , n43679 , n39532 );
and ( n46042 , n43671 , n39530 );
nor ( n46043 , n46041 , n46042 );
xnor ( n46044 , n46043 , n39497 );
and ( n46045 , n44000 , n39384 );
and ( n46046 , n43820 , n39382 );
nor ( n46047 , n46045 , n46046 );
xnor ( n46048 , n46047 , n39367 );
and ( n46049 , n46044 , n46048 );
and ( n46050 , n44347 , n39335 );
and ( n46051 , n44318 , n39333 );
nor ( n46052 , n46050 , n46051 );
xnor ( n46053 , n46052 , n39300 );
and ( n46054 , n46048 , n46053 );
and ( n46055 , n46044 , n46053 );
or ( n46056 , n46049 , n46054 , n46055 );
and ( n46057 , n45057 , n39258 );
and ( n46058 , n44826 , n39256 );
nor ( n46059 , n46057 , n46058 );
xnor ( n46060 , n46059 , n39215 );
and ( n46061 , n45754 , n39194 );
and ( n46062 , n45171 , n39192 );
nor ( n46063 , n46061 , n46062 );
xnor ( n46064 , n46063 , n39199 );
and ( n46065 , n46060 , n46064 );
xor ( n46066 , n39037 , n39101 );
buf ( n46067 , n46066 );
buf ( n46068 , n46067 );
buf ( n46069 , n46068 );
and ( n46070 , n46069 , n39186 );
and ( n46071 , n46064 , n46070 );
and ( n46072 , n46060 , n46070 );
or ( n46073 , n46065 , n46071 , n46072 );
and ( n46074 , n46056 , n46073 );
xor ( n46075 , n45760 , n45764 );
xor ( n46076 , n46075 , n45769 );
and ( n46077 , n46073 , n46076 );
and ( n46078 , n46056 , n46076 );
or ( n46079 , n46074 , n46077 , n46078 );
xor ( n46080 , n45777 , n45781 );
xor ( n46081 , n46080 , n45786 );
xor ( n46082 , n45803 , n45807 );
xor ( n46083 , n46082 , n45812 );
and ( n46084 , n46081 , n46083 );
xor ( n46085 , n45819 , n45823 );
xor ( n46086 , n46085 , n45828 );
and ( n46087 , n46083 , n46086 );
and ( n46088 , n46081 , n46086 );
or ( n46089 , n46084 , n46087 , n46088 );
and ( n46090 , n46079 , n46089 );
xor ( n46091 , n45738 , n45740 );
xor ( n46092 , n46091 , n45742 );
and ( n46093 , n46089 , n46092 );
and ( n46094 , n46079 , n46092 );
or ( n46095 , n46090 , n46093 , n46094 );
and ( n46096 , n46040 , n46095 );
xor ( n46097 , n45756 , n45772 );
xor ( n46098 , n46097 , n45789 );
xor ( n46099 , n45815 , n45831 );
xor ( n46100 , n46099 , n45848 );
and ( n46101 , n46098 , n46100 );
xor ( n46102 , n45853 , n45855 );
xor ( n46103 , n46102 , n45858 );
and ( n46104 , n46100 , n46103 );
and ( n46105 , n46098 , n46103 );
or ( n46106 , n46101 , n46104 , n46105 );
and ( n46107 , n46095 , n46106 );
and ( n46108 , n46040 , n46106 );
or ( n46109 , n46096 , n46107 , n46108 );
and ( n46110 , n45965 , n46109 );
and ( n46111 , n45956 , n46109 );
or ( n46112 , n45966 , n46110 , n46111 );
xor ( n46113 , n45724 , n45798 );
xor ( n46114 , n46113 , n45875 );
and ( n46115 , n46112 , n46114 );
xor ( n46116 , n45726 , n45733 );
xor ( n46117 , n46116 , n45795 );
xor ( n46118 , n45867 , n45869 );
xor ( n46119 , n46118 , n45872 );
and ( n46120 , n46117 , n46119 );
xor ( n46121 , n45736 , n45745 );
xor ( n46122 , n46121 , n45792 );
xor ( n46123 , n45851 , n45861 );
xor ( n46124 , n46123 , n45864 );
and ( n46125 , n46122 , n46124 );
xor ( n46126 , n45836 , n45840 );
xor ( n46127 , n46126 , n45845 );
buf ( n46128 , n30365 );
not ( n46129 , n46128 );
xnor ( n46130 , n45976 , n45980 );
and ( n46131 , n46129 , n46130 );
and ( n46132 , n43820 , n39532 );
and ( n46133 , n43679 , n39530 );
nor ( n46134 , n46132 , n46133 );
xnor ( n46135 , n46134 , n39497 );
and ( n46136 , n44318 , n39384 );
and ( n46137 , n44000 , n39382 );
nor ( n46138 , n46136 , n46137 );
xnor ( n46139 , n46138 , n39367 );
and ( n46140 , n46135 , n46139 );
and ( n46141 , n44826 , n39335 );
and ( n46142 , n44347 , n39333 );
nor ( n46143 , n46141 , n46142 );
xnor ( n46144 , n46143 , n39300 );
and ( n46145 , n46139 , n46144 );
and ( n46146 , n46135 , n46144 );
or ( n46147 , n46140 , n46145 , n46146 );
and ( n46148 , n46130 , n46147 );
and ( n46149 , n46129 , n46147 );
or ( n46150 , n46131 , n46148 , n46149 );
and ( n46151 , n46127 , n46150 );
and ( n46152 , n46069 , n39194 );
and ( n46153 , n45754 , n39192 );
nor ( n46154 , n46152 , n46153 );
xnor ( n46155 , n46154 , n39199 );
xor ( n46156 , n39040 , n39099 );
buf ( n46157 , n46156 );
buf ( n46158 , n46157 );
buf ( n46159 , n46158 );
and ( n46160 , n46159 , n39186 );
or ( n46161 , n46155 , n46160 );
and ( n46162 , n40698 , n42079 );
and ( n46163 , n40574 , n42076 );
nor ( n46164 , n46162 , n46163 );
xnor ( n46165 , n46164 , n41370 );
and ( n46166 , n40991 , n41981 );
and ( n46167 , n40962 , n41979 );
nor ( n46168 , n46166 , n46167 );
xnor ( n46169 , n46168 , n41373 );
and ( n46170 , n46165 , n46169 );
and ( n46171 , n41106 , n41522 );
and ( n46172 , n40910 , n41520 );
nor ( n46173 , n46171 , n46172 );
xnor ( n46174 , n46173 , n41100 );
and ( n46175 , n46169 , n46174 );
and ( n46176 , n46165 , n46174 );
or ( n46177 , n46170 , n46175 , n46176 );
and ( n46178 , n46161 , n46177 );
and ( n46179 , n41379 , n41230 );
and ( n46180 , n41091 , n41228 );
nor ( n46181 , n46179 , n46180 );
xnor ( n46182 , n46181 , n40981 );
and ( n46183 , n41735 , n40928 );
and ( n46184 , n41364 , n40926 );
nor ( n46185 , n46183 , n46184 );
xnor ( n46186 , n46185 , n40688 );
and ( n46187 , n46182 , n46186 );
and ( n46188 , n42149 , n40666 );
and ( n46189 , n41844 , n40664 );
nor ( n46190 , n46188 , n46189 );
xnor ( n46191 , n46190 , n40445 );
and ( n46192 , n46186 , n46191 );
and ( n46193 , n46182 , n46191 );
or ( n46194 , n46187 , n46192 , n46193 );
and ( n46195 , n46177 , n46194 );
and ( n46196 , n46161 , n46194 );
or ( n46197 , n46178 , n46195 , n46196 );
and ( n46198 , n46150 , n46197 );
and ( n46199 , n46127 , n46197 );
or ( n46200 , n46151 , n46198 , n46199 );
and ( n46201 , n42525 , n40406 );
and ( n46202 , n41828 , n40404 );
nor ( n46203 , n46201 , n46202 );
xnor ( n46204 , n46203 , n40262 );
and ( n46205 , n43040 , n40168 );
and ( n46206 , n42862 , n40166 );
nor ( n46207 , n46205 , n46206 );
xnor ( n46208 , n46207 , n40059 );
and ( n46209 , n46204 , n46208 );
and ( n46210 , n43322 , n39984 );
and ( n46211 , n43142 , n39982 );
nor ( n46212 , n46210 , n46211 );
xnor ( n46213 , n46212 , n39865 );
and ( n46214 , n46208 , n46213 );
and ( n46215 , n46204 , n46213 );
or ( n46216 , n46209 , n46214 , n46215 );
and ( n46217 , n43524 , n39795 );
and ( n46218 , n43387 , n39793 );
nor ( n46219 , n46217 , n46218 );
xnor ( n46220 , n46219 , n39729 );
and ( n46221 , n45171 , n39258 );
and ( n46222 , n45057 , n39256 );
nor ( n46223 , n46221 , n46222 );
xnor ( n46224 , n46223 , n39215 );
and ( n46225 , n46220 , n46224 );
buf ( n46226 , n30366 );
not ( n46227 , n46226 );
and ( n46228 , n46224 , n46227 );
and ( n46229 , n46220 , n46227 );
or ( n46230 , n46225 , n46228 , n46229 );
and ( n46231 , n46216 , n46230 );
xor ( n46232 , n45989 , n45993 );
xor ( n46233 , n46232 , n45998 );
and ( n46234 , n46230 , n46233 );
and ( n46235 , n46216 , n46233 );
or ( n46236 , n46231 , n46234 , n46235 );
xor ( n46237 , n46005 , n46009 );
xor ( n46238 , n46237 , n46014 );
xor ( n46239 , n46022 , n46026 );
xor ( n46240 , n46239 , n46031 );
and ( n46241 , n46238 , n46240 );
xor ( n46242 , n46044 , n46048 );
xor ( n46243 , n46242 , n46053 );
and ( n46244 , n46240 , n46243 );
and ( n46245 , n46238 , n46243 );
or ( n46246 , n46241 , n46244 , n46245 );
and ( n46247 , n46236 , n46246 );
xor ( n46248 , n45970 , n45971 );
xor ( n46249 , n46248 , n45981 );
and ( n46250 , n46246 , n46249 );
and ( n46251 , n46236 , n46249 );
or ( n46252 , n46247 , n46250 , n46251 );
and ( n46253 , n46200 , n46252 );
xor ( n46254 , n46001 , n46017 );
xor ( n46255 , n46254 , n46034 );
xor ( n46256 , n46056 , n46073 );
xor ( n46257 , n46256 , n46076 );
and ( n46258 , n46255 , n46257 );
xor ( n46259 , n46081 , n46083 );
xor ( n46260 , n46259 , n46086 );
and ( n46261 , n46257 , n46260 );
and ( n46262 , n46255 , n46260 );
or ( n46263 , n46258 , n46261 , n46262 );
and ( n46264 , n46252 , n46263 );
and ( n46265 , n46200 , n46263 );
or ( n46266 , n46253 , n46264 , n46265 );
and ( n46267 , n46124 , n46266 );
and ( n46268 , n46122 , n46266 );
or ( n46269 , n46125 , n46267 , n46268 );
and ( n46270 , n46119 , n46269 );
and ( n46271 , n46117 , n46269 );
or ( n46272 , n46120 , n46270 , n46271 );
and ( n46273 , n46114 , n46272 );
and ( n46274 , n46112 , n46272 );
or ( n46275 , n46115 , n46273 , n46274 );
xor ( n46276 , n45910 , n45912 );
xor ( n46277 , n46276 , n45915 );
and ( n46278 , n46275 , n46277 );
xor ( n46279 , n45903 , n45905 );
xor ( n46280 , n46279 , n45907 );
xor ( n46281 , n45968 , n45984 );
xor ( n46282 , n46281 , n46037 );
xor ( n46283 , n46079 , n46089 );
xor ( n46284 , n46283 , n46092 );
and ( n46285 , n46282 , n46284 );
xor ( n46286 , n46098 , n46100 );
xor ( n46287 , n46286 , n46103 );
and ( n46288 , n46284 , n46287 );
and ( n46289 , n46282 , n46287 );
or ( n46290 , n46285 , n46288 , n46289 );
xor ( n46291 , n45958 , n45960 );
xor ( n46292 , n46291 , n45962 );
and ( n46293 , n46290 , n46292 );
xor ( n46294 , n46040 , n46095 );
xor ( n46295 , n46294 , n46106 );
and ( n46296 , n46292 , n46295 );
and ( n46297 , n46290 , n46295 );
or ( n46298 , n46293 , n46296 , n46297 );
xor ( n46299 , n45956 , n45965 );
xor ( n46300 , n46299 , n46109 );
and ( n46301 , n46298 , n46300 );
xor ( n46302 , n46060 , n46064 );
xor ( n46303 , n46302 , n46070 );
and ( n46304 , n43671 , n39665 );
and ( n46305 , n43549 , n39663 );
nor ( n46306 , n46304 , n46305 );
xnor ( n46307 , n46306 , n39608 );
xor ( n46308 , n46135 , n46139 );
xor ( n46309 , n46308 , n46144 );
or ( n46310 , n46307 , n46309 );
and ( n46311 , n46303 , n46310 );
xnor ( n46312 , n46155 , n46160 );
and ( n46313 , n40962 , n42079 );
and ( n46314 , n40698 , n42076 );
nor ( n46315 , n46313 , n46314 );
xnor ( n46316 , n46315 , n41370 );
and ( n46317 , n40910 , n41981 );
and ( n46318 , n40991 , n41979 );
nor ( n46319 , n46317 , n46318 );
xnor ( n46320 , n46319 , n41373 );
or ( n46321 , n46316 , n46320 );
and ( n46322 , n46312 , n46321 );
and ( n46323 , n41091 , n41522 );
and ( n46324 , n41106 , n41520 );
nor ( n46325 , n46323 , n46324 );
xnor ( n46326 , n46325 , n41100 );
and ( n46327 , n41364 , n41230 );
and ( n46328 , n41379 , n41228 );
nor ( n46329 , n46327 , n46328 );
xnor ( n46330 , n46329 , n40981 );
and ( n46331 , n46326 , n46330 );
and ( n46332 , n46321 , n46331 );
and ( n46333 , n46312 , n46331 );
or ( n46334 , n46322 , n46332 , n46333 );
and ( n46335 , n46310 , n46334 );
and ( n46336 , n46303 , n46334 );
or ( n46337 , n46311 , n46335 , n46336 );
and ( n46338 , n41844 , n40928 );
and ( n46339 , n41735 , n40926 );
nor ( n46340 , n46338 , n46339 );
xnor ( n46341 , n46340 , n40688 );
and ( n46342 , n41828 , n40666 );
and ( n46343 , n42149 , n40664 );
nor ( n46344 , n46342 , n46343 );
xnor ( n46345 , n46344 , n40445 );
and ( n46346 , n46341 , n46345 );
and ( n46347 , n42862 , n40406 );
and ( n46348 , n42525 , n40404 );
nor ( n46349 , n46347 , n46348 );
xnor ( n46350 , n46349 , n40262 );
and ( n46351 , n46345 , n46350 );
and ( n46352 , n46341 , n46350 );
or ( n46353 , n46346 , n46351 , n46352 );
and ( n46354 , n43142 , n40168 );
and ( n46355 , n43040 , n40166 );
nor ( n46356 , n46354 , n46355 );
xnor ( n46357 , n46356 , n40059 );
and ( n46358 , n43387 , n39984 );
and ( n46359 , n43322 , n39982 );
nor ( n46360 , n46358 , n46359 );
xnor ( n46361 , n46360 , n39865 );
and ( n46362 , n46357 , n46361 );
and ( n46363 , n43549 , n39795 );
and ( n46364 , n43524 , n39793 );
nor ( n46365 , n46363 , n46364 );
xnor ( n46366 , n46365 , n39729 );
and ( n46367 , n46361 , n46366 );
and ( n46368 , n46357 , n46366 );
or ( n46369 , n46362 , n46367 , n46368 );
and ( n46370 , n46353 , n46369 );
and ( n46371 , n43679 , n39665 );
and ( n46372 , n43671 , n39663 );
nor ( n46373 , n46371 , n46372 );
xnor ( n46374 , n46373 , n39608 );
and ( n46375 , n44000 , n39532 );
and ( n46376 , n43820 , n39530 );
nor ( n46377 , n46375 , n46376 );
xnor ( n46378 , n46377 , n39497 );
and ( n46379 , n46374 , n46378 );
and ( n46380 , n44347 , n39384 );
and ( n46381 , n44318 , n39382 );
nor ( n46382 , n46380 , n46381 );
xnor ( n46383 , n46382 , n39367 );
and ( n46384 , n46378 , n46383 );
and ( n46385 , n46374 , n46383 );
or ( n46386 , n46379 , n46384 , n46385 );
and ( n46387 , n46369 , n46386 );
and ( n46388 , n46353 , n46386 );
or ( n46389 , n46370 , n46387 , n46388 );
and ( n46390 , n45057 , n39335 );
and ( n46391 , n44826 , n39333 );
nor ( n46392 , n46390 , n46391 );
xnor ( n46393 , n46392 , n39300 );
and ( n46394 , n45754 , n39258 );
and ( n46395 , n45171 , n39256 );
nor ( n46396 , n46394 , n46395 );
xnor ( n46397 , n46396 , n39215 );
and ( n46398 , n46393 , n46397 );
and ( n46399 , n46159 , n39194 );
and ( n46400 , n46069 , n39192 );
nor ( n46401 , n46399 , n46400 );
xnor ( n46402 , n46401 , n39199 );
and ( n46403 , n46397 , n46402 );
and ( n46404 , n46393 , n46402 );
or ( n46405 , n46398 , n46403 , n46404 );
xor ( n46406 , n46165 , n46169 );
xor ( n46407 , n46406 , n46174 );
and ( n46408 , n46405 , n46407 );
xor ( n46409 , n46182 , n46186 );
xor ( n46410 , n46409 , n46191 );
and ( n46411 , n46407 , n46410 );
and ( n46412 , n46405 , n46410 );
or ( n46413 , n46408 , n46411 , n46412 );
and ( n46414 , n46389 , n46413 );
xor ( n46415 , n46129 , n46130 );
xor ( n46416 , n46415 , n46147 );
and ( n46417 , n46413 , n46416 );
and ( n46418 , n46389 , n46416 );
or ( n46419 , n46414 , n46417 , n46418 );
and ( n46420 , n46337 , n46419 );
xor ( n46421 , n46161 , n46177 );
xor ( n46422 , n46421 , n46194 );
xor ( n46423 , n46216 , n46230 );
xor ( n46424 , n46423 , n46233 );
and ( n46425 , n46422 , n46424 );
xor ( n46426 , n46238 , n46240 );
xor ( n46427 , n46426 , n46243 );
and ( n46428 , n46424 , n46427 );
and ( n46429 , n46422 , n46427 );
or ( n46430 , n46425 , n46428 , n46429 );
and ( n46431 , n46419 , n46430 );
and ( n46432 , n46337 , n46430 );
or ( n46433 , n46420 , n46431 , n46432 );
xor ( n46434 , n46127 , n46150 );
xor ( n46435 , n46434 , n46197 );
xor ( n46436 , n46236 , n46246 );
xor ( n46437 , n46436 , n46249 );
and ( n46438 , n46435 , n46437 );
xor ( n46439 , n46255 , n46257 );
xor ( n46440 , n46439 , n46260 );
and ( n46441 , n46437 , n46440 );
and ( n46442 , n46435 , n46440 );
or ( n46443 , n46438 , n46441 , n46442 );
and ( n46444 , n46433 , n46443 );
xor ( n46445 , n46200 , n46252 );
xor ( n46446 , n46445 , n46263 );
and ( n46447 , n46443 , n46446 );
and ( n46448 , n46433 , n46446 );
or ( n46449 , n46444 , n46447 , n46448 );
xor ( n46450 , n46122 , n46124 );
xor ( n46451 , n46450 , n46266 );
and ( n46452 , n46449 , n46451 );
xor ( n46453 , n46290 , n46292 );
xor ( n46454 , n46453 , n46295 );
and ( n46455 , n46451 , n46454 );
and ( n46456 , n46449 , n46454 );
or ( n46457 , n46452 , n46455 , n46456 );
and ( n46458 , n46300 , n46457 );
and ( n46459 , n46298 , n46457 );
or ( n46460 , n46301 , n46458 , n46459 );
and ( n46461 , n46280 , n46460 );
xor ( n46462 , n46112 , n46114 );
xor ( n46463 , n46462 , n46272 );
and ( n46464 , n46460 , n46463 );
and ( n46465 , n46280 , n46463 );
or ( n46466 , n46461 , n46464 , n46465 );
and ( n46467 , n46277 , n46466 );
and ( n46468 , n46275 , n46466 );
or ( n46469 , n46278 , n46467 , n46468 );
or ( n46470 , n45955 , n46469 );
xor ( n46471 , n45926 , n45928 );
xor ( n46472 , n46471 , n45931 );
or ( n46473 , n46470 , n46472 );
or ( n46474 , n45953 , n46473 );
xor ( n46475 , n45701 , n45937 );
xor ( n46476 , n46475 , n45940 );
and ( n46477 , n46474 , n46476 );
xor ( n46478 , n46474 , n46476 );
xor ( n46479 , n45898 , n45900 );
xor ( n46480 , n46479 , n45934 );
xnor ( n46481 , n45953 , n46473 );
and ( n46482 , n46480 , n46481 );
xor ( n46483 , n46480 , n46481 );
xnor ( n46484 , n46470 , n46472 );
xnor ( n46485 , n45955 , n46469 );
xor ( n46486 , n46275 , n46277 );
xor ( n46487 , n46486 , n46466 );
not ( n46488 , n46487 );
xor ( n46489 , n46280 , n46460 );
xor ( n46490 , n46489 , n46463 );
xor ( n46491 , n46117 , n46119 );
xor ( n46492 , n46491 , n46269 );
xor ( n46493 , n46298 , n46300 );
xor ( n46494 , n46493 , n46457 );
and ( n46495 , n46492 , n46494 );
xor ( n46496 , n46282 , n46284 );
xor ( n46497 , n46496 , n46287 );
xor ( n46498 , n46204 , n46208 );
xor ( n46499 , n46498 , n46213 );
xor ( n46500 , n46220 , n46224 );
xor ( n46501 , n46500 , n46227 );
and ( n46502 , n46499 , n46501 );
xnor ( n46503 , n46307 , n46309 );
and ( n46504 , n46501 , n46503 );
and ( n46505 , n46499 , n46503 );
or ( n46506 , n46502 , n46504 , n46505 );
xor ( n46507 , n39043 , n39097 );
buf ( n46508 , n46507 );
buf ( n46509 , n46508 );
buf ( n46510 , n46509 );
and ( n46511 , n46510 , n39186 );
buf ( n46512 , n30367 );
not ( n46513 , n46512 );
and ( n46514 , n46511 , n46513 );
xnor ( n46515 , n46316 , n46320 );
and ( n46516 , n46513 , n46515 );
and ( n46517 , n46511 , n46515 );
or ( n46518 , n46514 , n46516 , n46517 );
xor ( n46519 , n46326 , n46330 );
and ( n46520 , n43820 , n39665 );
and ( n46521 , n43679 , n39663 );
nor ( n46522 , n46520 , n46521 );
xnor ( n46523 , n46522 , n39608 );
and ( n46524 , n44318 , n39532 );
and ( n46525 , n44000 , n39530 );
nor ( n46526 , n46524 , n46525 );
xnor ( n46527 , n46526 , n39497 );
and ( n46528 , n46523 , n46527 );
and ( n46529 , n44826 , n39384 );
and ( n46530 , n44347 , n39382 );
nor ( n46531 , n46529 , n46530 );
xnor ( n46532 , n46531 , n39367 );
and ( n46533 , n46527 , n46532 );
and ( n46534 , n46523 , n46532 );
or ( n46535 , n46528 , n46533 , n46534 );
and ( n46536 , n46519 , n46535 );
and ( n46537 , n40991 , n42079 );
and ( n46538 , n40962 , n42076 );
nor ( n46539 , n46537 , n46538 );
xnor ( n46540 , n46539 , n41370 );
and ( n46541 , n41106 , n41981 );
and ( n46542 , n40910 , n41979 );
nor ( n46543 , n46541 , n46542 );
xnor ( n46544 , n46543 , n41373 );
and ( n46545 , n46540 , n46544 );
and ( n46546 , n41379 , n41522 );
and ( n46547 , n41091 , n41520 );
nor ( n46548 , n46546 , n46547 );
xnor ( n46549 , n46548 , n41100 );
and ( n46550 , n46544 , n46549 );
and ( n46551 , n46540 , n46549 );
or ( n46552 , n46545 , n46550 , n46551 );
and ( n46553 , n46535 , n46552 );
and ( n46554 , n46519 , n46552 );
or ( n46555 , n46536 , n46553 , n46554 );
and ( n46556 , n46518 , n46555 );
and ( n46557 , n41735 , n41230 );
and ( n46558 , n41364 , n41228 );
nor ( n46559 , n46557 , n46558 );
xnor ( n46560 , n46559 , n40981 );
and ( n46561 , n42149 , n40928 );
and ( n46562 , n41844 , n40926 );
nor ( n46563 , n46561 , n46562 );
xnor ( n46564 , n46563 , n40688 );
and ( n46565 , n46560 , n46564 );
and ( n46566 , n42525 , n40666 );
and ( n46567 , n41828 , n40664 );
nor ( n46568 , n46566 , n46567 );
xnor ( n46569 , n46568 , n40445 );
and ( n46570 , n46564 , n46569 );
and ( n46571 , n46560 , n46569 );
or ( n46572 , n46565 , n46570 , n46571 );
and ( n46573 , n43040 , n40406 );
and ( n46574 , n42862 , n40404 );
nor ( n46575 , n46573 , n46574 );
xnor ( n46576 , n46575 , n40262 );
and ( n46577 , n43322 , n40168 );
and ( n46578 , n43142 , n40166 );
nor ( n46579 , n46577 , n46578 );
xnor ( n46580 , n46579 , n40059 );
and ( n46581 , n46576 , n46580 );
and ( n46582 , n43524 , n39984 );
and ( n46583 , n43387 , n39982 );
nor ( n46584 , n46582 , n46583 );
xnor ( n46585 , n46584 , n39865 );
and ( n46586 , n46580 , n46585 );
and ( n46587 , n46576 , n46585 );
or ( n46588 , n46581 , n46586 , n46587 );
and ( n46589 , n46572 , n46588 );
and ( n46590 , n45171 , n39335 );
and ( n46591 , n45057 , n39333 );
nor ( n46592 , n46590 , n46591 );
xnor ( n46593 , n46592 , n39300 );
and ( n46594 , n46069 , n39258 );
and ( n46595 , n45754 , n39256 );
nor ( n46596 , n46594 , n46595 );
xnor ( n46597 , n46596 , n39215 );
and ( n46598 , n46593 , n46597 );
and ( n46599 , n46510 , n39194 );
and ( n46600 , n46159 , n39192 );
nor ( n46601 , n46599 , n46600 );
xnor ( n46602 , n46601 , n39199 );
and ( n46603 , n46597 , n46602 );
and ( n46604 , n46593 , n46602 );
or ( n46605 , n46598 , n46603 , n46604 );
and ( n46606 , n46588 , n46605 );
and ( n46607 , n46572 , n46605 );
or ( n46608 , n46589 , n46606 , n46607 );
and ( n46609 , n46555 , n46608 );
and ( n46610 , n46518 , n46608 );
or ( n46611 , n46556 , n46609 , n46610 );
and ( n46612 , n46506 , n46611 );
xor ( n46613 , n46341 , n46345 );
xor ( n46614 , n46613 , n46350 );
xor ( n46615 , n46357 , n46361 );
xor ( n46616 , n46615 , n46366 );
and ( n46617 , n46614 , n46616 );
xor ( n46618 , n46374 , n46378 );
xor ( n46619 , n46618 , n46383 );
and ( n46620 , n46616 , n46619 );
and ( n46621 , n46614 , n46619 );
or ( n46622 , n46617 , n46620 , n46621 );
xor ( n46623 , n46312 , n46321 );
xor ( n46624 , n46623 , n46331 );
and ( n46625 , n46622 , n46624 );
xor ( n46626 , n46353 , n46369 );
xor ( n46627 , n46626 , n46386 );
and ( n46628 , n46624 , n46627 );
and ( n46629 , n46622 , n46627 );
or ( n46630 , n46625 , n46628 , n46629 );
and ( n46631 , n46611 , n46630 );
and ( n46632 , n46506 , n46630 );
or ( n46633 , n46612 , n46631 , n46632 );
xor ( n46634 , n46303 , n46310 );
xor ( n46635 , n46634 , n46334 );
xor ( n46636 , n46389 , n46413 );
xor ( n46637 , n46636 , n46416 );
and ( n46638 , n46635 , n46637 );
xor ( n46639 , n46422 , n46424 );
xor ( n46640 , n46639 , n46427 );
and ( n46641 , n46637 , n46640 );
and ( n46642 , n46635 , n46640 );
or ( n46643 , n46638 , n46641 , n46642 );
and ( n46644 , n46633 , n46643 );
xor ( n46645 , n46337 , n46419 );
xor ( n46646 , n46645 , n46430 );
and ( n46647 , n46643 , n46646 );
and ( n46648 , n46633 , n46646 );
or ( n46649 , n46644 , n46647 , n46648 );
and ( n46650 , n46497 , n46649 );
xor ( n46651 , n46433 , n46443 );
xor ( n46652 , n46651 , n46446 );
and ( n46653 , n46649 , n46652 );
and ( n46654 , n46497 , n46652 );
or ( n46655 , n46650 , n46653 , n46654 );
xor ( n46656 , n46449 , n46451 );
xor ( n46657 , n46656 , n46454 );
and ( n46658 , n46655 , n46657 );
xor ( n46659 , n46435 , n46437 );
xor ( n46660 , n46659 , n46440 );
xor ( n46661 , n46405 , n46407 );
xor ( n46662 , n46661 , n46410 );
xor ( n46663 , n46393 , n46397 );
xor ( n46664 , n46663 , n46402 );
and ( n46665 , n43671 , n39795 );
and ( n46666 , n43549 , n39793 );
nor ( n46667 , n46665 , n46666 );
xnor ( n46668 , n46667 , n39729 );
xor ( n46669 , n46523 , n46527 );
xor ( n46670 , n46669 , n46532 );
or ( n46671 , n46668 , n46670 );
and ( n46672 , n46664 , n46671 );
xor ( n46673 , n39044 , n39096 );
buf ( n46674 , n46673 );
buf ( n46675 , n46674 );
buf ( n46676 , n46675 );
and ( n46677 , n46676 , n39186 );
buf ( n46678 , n30368 );
not ( n46679 , n46678 );
and ( n46680 , n46677 , n46679 );
and ( n46681 , n41091 , n41981 );
and ( n46682 , n41106 , n41979 );
nor ( n46683 , n46681 , n46682 );
xnor ( n46684 , n46683 , n41373 );
and ( n46685 , n41364 , n41522 );
and ( n46686 , n41379 , n41520 );
nor ( n46687 , n46685 , n46686 );
xnor ( n46688 , n46687 , n41100 );
and ( n46689 , n46684 , n46688 );
and ( n46690 , n46679 , n46689 );
and ( n46691 , n46677 , n46689 );
or ( n46692 , n46680 , n46690 , n46691 );
and ( n46693 , n46671 , n46692 );
and ( n46694 , n46664 , n46692 );
or ( n46695 , n46672 , n46693 , n46694 );
and ( n46696 , n46662 , n46695 );
and ( n46697 , n40910 , n42079 );
and ( n46698 , n40991 , n42076 );
nor ( n46699 , n46697 , n46698 );
xnor ( n46700 , n46699 , n41370 );
and ( n46701 , n41844 , n41230 );
and ( n46702 , n41735 , n41228 );
nor ( n46703 , n46701 , n46702 );
xnor ( n46704 , n46703 , n40981 );
and ( n46705 , n46700 , n46704 );
and ( n46706 , n41828 , n40928 );
and ( n46707 , n42149 , n40926 );
nor ( n46708 , n46706 , n46707 );
xnor ( n46709 , n46708 , n40688 );
and ( n46710 , n46704 , n46709 );
and ( n46711 , n46700 , n46709 );
or ( n46712 , n46705 , n46710 , n46711 );
and ( n46713 , n42862 , n40666 );
and ( n46714 , n42525 , n40664 );
nor ( n46715 , n46713 , n46714 );
xnor ( n46716 , n46715 , n40445 );
and ( n46717 , n43142 , n40406 );
and ( n46718 , n43040 , n40404 );
nor ( n46719 , n46717 , n46718 );
xnor ( n46720 , n46719 , n40262 );
and ( n46721 , n46716 , n46720 );
and ( n46722 , n43387 , n40168 );
and ( n46723 , n43322 , n40166 );
nor ( n46724 , n46722 , n46723 );
xnor ( n46725 , n46724 , n40059 );
and ( n46726 , n46720 , n46725 );
and ( n46727 , n46716 , n46725 );
or ( n46728 , n46721 , n46726 , n46727 );
and ( n46729 , n46712 , n46728 );
and ( n46730 , n43549 , n39984 );
and ( n46731 , n43524 , n39982 );
nor ( n46732 , n46730 , n46731 );
xnor ( n46733 , n46732 , n39865 );
and ( n46734 , n43679 , n39795 );
and ( n46735 , n43671 , n39793 );
nor ( n46736 , n46734 , n46735 );
xnor ( n46737 , n46736 , n39729 );
and ( n46738 , n46733 , n46737 );
and ( n46739 , n44000 , n39665 );
and ( n46740 , n43820 , n39663 );
nor ( n46741 , n46739 , n46740 );
xnor ( n46742 , n46741 , n39608 );
and ( n46743 , n46737 , n46742 );
and ( n46744 , n46733 , n46742 );
or ( n46745 , n46738 , n46743 , n46744 );
and ( n46746 , n46728 , n46745 );
and ( n46747 , n46712 , n46745 );
or ( n46748 , n46729 , n46746 , n46747 );
and ( n46749 , n44347 , n39532 );
and ( n46750 , n44318 , n39530 );
nor ( n46751 , n46749 , n46750 );
xnor ( n46752 , n46751 , n39497 );
and ( n46753 , n45057 , n39384 );
and ( n46754 , n44826 , n39382 );
nor ( n46755 , n46753 , n46754 );
xnor ( n46756 , n46755 , n39367 );
and ( n46757 , n46752 , n46756 );
and ( n46758 , n45754 , n39335 );
and ( n46759 , n45171 , n39333 );
nor ( n46760 , n46758 , n46759 );
xnor ( n46761 , n46760 , n39300 );
and ( n46762 , n46756 , n46761 );
and ( n46763 , n46752 , n46761 );
or ( n46764 , n46757 , n46762 , n46763 );
and ( n46765 , n46159 , n39258 );
and ( n46766 , n46069 , n39256 );
nor ( n46767 , n46765 , n46766 );
xnor ( n46768 , n46767 , n39215 );
and ( n46769 , n46676 , n39194 );
and ( n46770 , n46510 , n39192 );
nor ( n46771 , n46769 , n46770 );
xnor ( n46772 , n46771 , n39199 );
and ( n46773 , n46768 , n46772 );
xor ( n46774 , n39046 , n39095 );
buf ( n46775 , n46774 );
buf ( n46776 , n46775 );
buf ( n46777 , n46776 );
and ( n46778 , n46777 , n39186 );
and ( n46779 , n46772 , n46778 );
and ( n46780 , n46768 , n46778 );
or ( n46781 , n46773 , n46779 , n46780 );
and ( n46782 , n46764 , n46781 );
xor ( n46783 , n46540 , n46544 );
xor ( n46784 , n46783 , n46549 );
and ( n46785 , n46781 , n46784 );
and ( n46786 , n46764 , n46784 );
or ( n46787 , n46782 , n46785 , n46786 );
and ( n46788 , n46748 , n46787 );
xor ( n46789 , n46560 , n46564 );
xor ( n46790 , n46789 , n46569 );
xor ( n46791 , n46576 , n46580 );
xor ( n46792 , n46791 , n46585 );
and ( n46793 , n46790 , n46792 );
xor ( n46794 , n46593 , n46597 );
xor ( n46795 , n46794 , n46602 );
and ( n46796 , n46792 , n46795 );
and ( n46797 , n46790 , n46795 );
or ( n46798 , n46793 , n46796 , n46797 );
and ( n46799 , n46787 , n46798 );
and ( n46800 , n46748 , n46798 );
or ( n46801 , n46788 , n46799 , n46800 );
and ( n46802 , n46695 , n46801 );
and ( n46803 , n46662 , n46801 );
or ( n46804 , n46696 , n46802 , n46803 );
xor ( n46805 , n46511 , n46513 );
xor ( n46806 , n46805 , n46515 );
xor ( n46807 , n46519 , n46535 );
xor ( n46808 , n46807 , n46552 );
and ( n46809 , n46806 , n46808 );
xor ( n46810 , n46572 , n46588 );
xor ( n46811 , n46810 , n46605 );
and ( n46812 , n46808 , n46811 );
and ( n46813 , n46806 , n46811 );
or ( n46814 , n46809 , n46812 , n46813 );
xor ( n46815 , n46499 , n46501 );
xor ( n46816 , n46815 , n46503 );
and ( n46817 , n46814 , n46816 );
xor ( n46818 , n46518 , n46555 );
xor ( n46819 , n46818 , n46608 );
and ( n46820 , n46816 , n46819 );
and ( n46821 , n46814 , n46819 );
or ( n46822 , n46817 , n46820 , n46821 );
and ( n46823 , n46804 , n46822 );
xor ( n46824 , n46506 , n46611 );
xor ( n46825 , n46824 , n46630 );
and ( n46826 , n46822 , n46825 );
and ( n46827 , n46804 , n46825 );
or ( n46828 , n46823 , n46826 , n46827 );
and ( n46829 , n46660 , n46828 );
xor ( n46830 , n46633 , n46643 );
xor ( n46831 , n46830 , n46646 );
and ( n46832 , n46828 , n46831 );
and ( n46833 , n46660 , n46831 );
or ( n46834 , n46829 , n46832 , n46833 );
xor ( n46835 , n46497 , n46649 );
xor ( n46836 , n46835 , n46652 );
and ( n46837 , n46834 , n46836 );
xor ( n46838 , n46635 , n46637 );
xor ( n46839 , n46838 , n46640 );
xor ( n46840 , n46622 , n46624 );
xor ( n46841 , n46840 , n46627 );
xor ( n46842 , n46614 , n46616 );
xor ( n46843 , n46842 , n46619 );
xnor ( n46844 , n46668 , n46670 );
buf ( n46845 , n30369 );
not ( n46846 , n46845 );
xor ( n46847 , n46684 , n46688 );
and ( n46848 , n46846 , n46847 );
and ( n46849 , n43820 , n39795 );
and ( n46850 , n43679 , n39793 );
nor ( n46851 , n46849 , n46850 );
xnor ( n46852 , n46851 , n39729 );
and ( n46853 , n44318 , n39665 );
and ( n46854 , n44000 , n39663 );
nor ( n46855 , n46853 , n46854 );
xnor ( n46856 , n46855 , n39608 );
and ( n46857 , n46852 , n46856 );
and ( n46858 , n44826 , n39532 );
and ( n46859 , n44347 , n39530 );
nor ( n46860 , n46858 , n46859 );
xnor ( n46861 , n46860 , n39497 );
and ( n46862 , n46856 , n46861 );
and ( n46863 , n46852 , n46861 );
or ( n46864 , n46857 , n46862 , n46863 );
and ( n46865 , n46847 , n46864 );
and ( n46866 , n46846 , n46864 );
or ( n46867 , n46848 , n46865 , n46866 );
and ( n46868 , n46844 , n46867 );
and ( n46869 , n41106 , n42079 );
and ( n46870 , n40910 , n42076 );
nor ( n46871 , n46869 , n46870 );
xnor ( n46872 , n46871 , n41370 );
and ( n46873 , n41379 , n41981 );
and ( n46874 , n41091 , n41979 );
nor ( n46875 , n46873 , n46874 );
xnor ( n46876 , n46875 , n41373 );
and ( n46877 , n46872 , n46876 );
and ( n46878 , n41735 , n41522 );
and ( n46879 , n41364 , n41520 );
nor ( n46880 , n46878 , n46879 );
xnor ( n46881 , n46880 , n41100 );
and ( n46882 , n46876 , n46881 );
and ( n46883 , n46872 , n46881 );
or ( n46884 , n46877 , n46882 , n46883 );
and ( n46885 , n42149 , n41230 );
and ( n46886 , n41844 , n41228 );
nor ( n46887 , n46885 , n46886 );
xnor ( n46888 , n46887 , n40981 );
and ( n46889 , n42525 , n40928 );
and ( n46890 , n41828 , n40926 );
nor ( n46891 , n46889 , n46890 );
xnor ( n46892 , n46891 , n40688 );
and ( n46893 , n46888 , n46892 );
and ( n46894 , n43040 , n40666 );
and ( n46895 , n42862 , n40664 );
nor ( n46896 , n46894 , n46895 );
xnor ( n46897 , n46896 , n40445 );
and ( n46898 , n46892 , n46897 );
and ( n46899 , n46888 , n46897 );
or ( n46900 , n46893 , n46898 , n46899 );
and ( n46901 , n46884 , n46900 );
and ( n46902 , n43322 , n40406 );
and ( n46903 , n43142 , n40404 );
nor ( n46904 , n46902 , n46903 );
xnor ( n46905 , n46904 , n40262 );
and ( n46906 , n43524 , n40168 );
and ( n46907 , n43387 , n40166 );
nor ( n46908 , n46906 , n46907 );
xnor ( n46909 , n46908 , n40059 );
and ( n46910 , n46905 , n46909 );
and ( n46911 , n43671 , n39984 );
and ( n46912 , n43549 , n39982 );
nor ( n46913 , n46911 , n46912 );
xnor ( n46914 , n46913 , n39865 );
and ( n46915 , n46909 , n46914 );
and ( n46916 , n46905 , n46914 );
or ( n46917 , n46910 , n46915 , n46916 );
and ( n46918 , n46900 , n46917 );
and ( n46919 , n46884 , n46917 );
or ( n46920 , n46901 , n46918 , n46919 );
and ( n46921 , n46867 , n46920 );
and ( n46922 , n46844 , n46920 );
or ( n46923 , n46868 , n46921 , n46922 );
and ( n46924 , n46843 , n46923 );
and ( n46925 , n45171 , n39384 );
and ( n46926 , n45057 , n39382 );
nor ( n46927 , n46925 , n46926 );
xnor ( n46928 , n46927 , n39367 );
and ( n46929 , n46069 , n39335 );
and ( n46930 , n45754 , n39333 );
nor ( n46931 , n46929 , n46930 );
xnor ( n46932 , n46931 , n39300 );
and ( n46933 , n46928 , n46932 );
and ( n46934 , n46510 , n39258 );
and ( n46935 , n46159 , n39256 );
nor ( n46936 , n46934 , n46935 );
xnor ( n46937 , n46936 , n39215 );
and ( n46938 , n46932 , n46937 );
and ( n46939 , n46928 , n46937 );
or ( n46940 , n46933 , n46938 , n46939 );
and ( n46941 , n46777 , n39194 );
and ( n46942 , n46676 , n39192 );
nor ( n46943 , n46941 , n46942 );
xnor ( n46944 , n46943 , n39199 );
xor ( n46945 , n39049 , n39093 );
buf ( n46946 , n46945 );
buf ( n46947 , n46946 );
buf ( n46948 , n46947 );
and ( n46949 , n46948 , n39186 );
and ( n46950 , n46944 , n46949 );
buf ( n46951 , n30370 );
not ( n46952 , n46951 );
and ( n46953 , n46949 , n46952 );
and ( n46954 , n46944 , n46952 );
or ( n46955 , n46950 , n46953 , n46954 );
and ( n46956 , n46940 , n46955 );
xor ( n46957 , n46700 , n46704 );
xor ( n46958 , n46957 , n46709 );
and ( n46959 , n46955 , n46958 );
and ( n46960 , n46940 , n46958 );
or ( n46961 , n46956 , n46959 , n46960 );
xor ( n46962 , n46716 , n46720 );
xor ( n46963 , n46962 , n46725 );
xor ( n46964 , n46733 , n46737 );
xor ( n46965 , n46964 , n46742 );
and ( n46966 , n46963 , n46965 );
xor ( n46967 , n46752 , n46756 );
xor ( n46968 , n46967 , n46761 );
and ( n46969 , n46965 , n46968 );
and ( n46970 , n46963 , n46968 );
or ( n46971 , n46966 , n46969 , n46970 );
and ( n46972 , n46961 , n46971 );
xor ( n46973 , n46677 , n46679 );
xor ( n46974 , n46973 , n46689 );
and ( n46975 , n46971 , n46974 );
and ( n46976 , n46961 , n46974 );
or ( n46977 , n46972 , n46975 , n46976 );
and ( n46978 , n46923 , n46977 );
and ( n46979 , n46843 , n46977 );
or ( n46980 , n46924 , n46978 , n46979 );
and ( n46981 , n46841 , n46980 );
xor ( n46982 , n46712 , n46728 );
xor ( n46983 , n46982 , n46745 );
xor ( n46984 , n46764 , n46781 );
xor ( n46985 , n46984 , n46784 );
and ( n46986 , n46983 , n46985 );
xor ( n46987 , n46790 , n46792 );
xor ( n46988 , n46987 , n46795 );
and ( n46989 , n46985 , n46988 );
and ( n46990 , n46983 , n46988 );
or ( n46991 , n46986 , n46989 , n46990 );
xor ( n46992 , n46664 , n46671 );
xor ( n46993 , n46992 , n46692 );
and ( n46994 , n46991 , n46993 );
xor ( n46995 , n46748 , n46787 );
xor ( n46996 , n46995 , n46798 );
and ( n46997 , n46993 , n46996 );
and ( n46998 , n46991 , n46996 );
or ( n46999 , n46994 , n46997 , n46998 );
and ( n47000 , n46980 , n46999 );
and ( n47001 , n46841 , n46999 );
or ( n47002 , n46981 , n47000 , n47001 );
and ( n47003 , n46839 , n47002 );
xor ( n47004 , n46804 , n46822 );
xor ( n47005 , n47004 , n46825 );
and ( n47006 , n47002 , n47005 );
and ( n47007 , n46839 , n47005 );
or ( n47008 , n47003 , n47006 , n47007 );
xor ( n47009 , n46660 , n46828 );
xor ( n47010 , n47009 , n46831 );
and ( n47011 , n47008 , n47010 );
xor ( n47012 , n46662 , n46695 );
xor ( n47013 , n47012 , n46801 );
xor ( n47014 , n46814 , n46816 );
xor ( n47015 , n47014 , n46819 );
and ( n47016 , n47013 , n47015 );
xor ( n47017 , n46806 , n46808 );
xor ( n47018 , n47017 , n46811 );
xor ( n47019 , n46768 , n46772 );
xor ( n47020 , n47019 , n46778 );
xor ( n47021 , n46852 , n46856 );
xor ( n47022 , n47021 , n46861 );
and ( n47023 , n41091 , n42079 );
and ( n47024 , n41106 , n42076 );
nor ( n47025 , n47023 , n47024 );
xnor ( n47026 , n47025 , n41370 );
and ( n47027 , n41364 , n41981 );
and ( n47028 , n41379 , n41979 );
nor ( n47029 , n47027 , n47028 );
xnor ( n47030 , n47029 , n41373 );
or ( n47031 , n47026 , n47030 );
and ( n47032 , n47022 , n47031 );
and ( n47033 , n41844 , n41522 );
and ( n47034 , n41735 , n41520 );
nor ( n47035 , n47033 , n47034 );
xnor ( n47036 , n47035 , n41100 );
and ( n47037 , n41828 , n41230 );
and ( n47038 , n42149 , n41228 );
nor ( n47039 , n47037 , n47038 );
xnor ( n47040 , n47039 , n40981 );
and ( n47041 , n47036 , n47040 );
and ( n47042 , n42862 , n40928 );
and ( n47043 , n42525 , n40926 );
nor ( n47044 , n47042 , n47043 );
xnor ( n47045 , n47044 , n40688 );
and ( n47046 , n47040 , n47045 );
and ( n47047 , n47036 , n47045 );
or ( n47048 , n47041 , n47046 , n47047 );
and ( n47049 , n47031 , n47048 );
and ( n47050 , n47022 , n47048 );
or ( n47051 , n47032 , n47049 , n47050 );
and ( n47052 , n47020 , n47051 );
and ( n47053 , n43142 , n40666 );
and ( n47054 , n43040 , n40664 );
nor ( n47055 , n47053 , n47054 );
xnor ( n47056 , n47055 , n40445 );
and ( n47057 , n43387 , n40406 );
and ( n47058 , n43322 , n40404 );
nor ( n47059 , n47057 , n47058 );
xnor ( n47060 , n47059 , n40262 );
and ( n47061 , n47056 , n47060 );
and ( n47062 , n43549 , n40168 );
and ( n47063 , n43524 , n40166 );
nor ( n47064 , n47062 , n47063 );
xnor ( n47065 , n47064 , n40059 );
and ( n47066 , n47060 , n47065 );
and ( n47067 , n47056 , n47065 );
or ( n47068 , n47061 , n47066 , n47067 );
and ( n47069 , n43679 , n39984 );
and ( n47070 , n43671 , n39982 );
nor ( n47071 , n47069 , n47070 );
xnor ( n47072 , n47071 , n39865 );
and ( n47073 , n44000 , n39795 );
and ( n47074 , n43820 , n39793 );
nor ( n47075 , n47073 , n47074 );
xnor ( n47076 , n47075 , n39729 );
and ( n47077 , n47072 , n47076 );
and ( n47078 , n44347 , n39665 );
and ( n47079 , n44318 , n39663 );
nor ( n47080 , n47078 , n47079 );
xnor ( n47081 , n47080 , n39608 );
and ( n47082 , n47076 , n47081 );
and ( n47083 , n47072 , n47081 );
or ( n47084 , n47077 , n47082 , n47083 );
and ( n47085 , n47068 , n47084 );
and ( n47086 , n45057 , n39532 );
and ( n47087 , n44826 , n39530 );
nor ( n47088 , n47086 , n47087 );
xnor ( n47089 , n47088 , n39497 );
and ( n47090 , n45754 , n39384 );
and ( n47091 , n45171 , n39382 );
nor ( n47092 , n47090 , n47091 );
xnor ( n47093 , n47092 , n39367 );
and ( n47094 , n47089 , n47093 );
and ( n47095 , n46159 , n39335 );
and ( n47096 , n46069 , n39333 );
nor ( n47097 , n47095 , n47096 );
xnor ( n47098 , n47097 , n39300 );
and ( n47099 , n47093 , n47098 );
and ( n47100 , n47089 , n47098 );
or ( n47101 , n47094 , n47099 , n47100 );
and ( n47102 , n47084 , n47101 );
and ( n47103 , n47068 , n47101 );
or ( n47104 , n47085 , n47102 , n47103 );
and ( n47105 , n47051 , n47104 );
and ( n47106 , n47020 , n47104 );
or ( n47107 , n47052 , n47105 , n47106 );
xor ( n47108 , n46872 , n46876 );
xor ( n47109 , n47108 , n46881 );
xor ( n47110 , n46888 , n46892 );
xor ( n47111 , n47110 , n46897 );
and ( n47112 , n47109 , n47111 );
xor ( n47113 , n46905 , n46909 );
xor ( n47114 , n47113 , n46914 );
and ( n47115 , n47111 , n47114 );
and ( n47116 , n47109 , n47114 );
or ( n47117 , n47112 , n47115 , n47116 );
xor ( n47118 , n46846 , n46847 );
xor ( n47119 , n47118 , n46864 );
and ( n47120 , n47117 , n47119 );
xor ( n47121 , n46884 , n46900 );
xor ( n47122 , n47121 , n46917 );
and ( n47123 , n47119 , n47122 );
and ( n47124 , n47117 , n47122 );
or ( n47125 , n47120 , n47123 , n47124 );
and ( n47126 , n47107 , n47125 );
xor ( n47127 , n46844 , n46867 );
xor ( n47128 , n47127 , n46920 );
and ( n47129 , n47125 , n47128 );
and ( n47130 , n47107 , n47128 );
or ( n47131 , n47126 , n47129 , n47130 );
and ( n47132 , n47018 , n47131 );
xor ( n47133 , n46843 , n46923 );
xor ( n47134 , n47133 , n46977 );
and ( n47135 , n47131 , n47134 );
and ( n47136 , n47018 , n47134 );
or ( n47137 , n47132 , n47135 , n47136 );
and ( n47138 , n47015 , n47137 );
and ( n47139 , n47013 , n47137 );
or ( n47140 , n47016 , n47138 , n47139 );
xor ( n47141 , n46839 , n47002 );
xor ( n47142 , n47141 , n47005 );
and ( n47143 , n47140 , n47142 );
xor ( n47144 , n46841 , n46980 );
xor ( n47145 , n47144 , n46999 );
xor ( n47146 , n46991 , n46993 );
xor ( n47147 , n47146 , n46996 );
xor ( n47148 , n46961 , n46971 );
xor ( n47149 , n47148 , n46974 );
xor ( n47150 , n46983 , n46985 );
xor ( n47151 , n47150 , n46988 );
and ( n47152 , n47149 , n47151 );
xor ( n47153 , n46940 , n46955 );
xor ( n47154 , n47153 , n46958 );
xor ( n47155 , n46963 , n46965 );
xor ( n47156 , n47155 , n46968 );
and ( n47157 , n47154 , n47156 );
xor ( n47158 , n46928 , n46932 );
xor ( n47159 , n47158 , n46937 );
xor ( n47160 , n46944 , n46949 );
xor ( n47161 , n47160 , n46952 );
and ( n47162 , n47159 , n47161 );
buf ( n47163 , n30371 );
not ( n47164 , n47163 );
xnor ( n47165 , n47026 , n47030 );
and ( n47166 , n47164 , n47165 );
and ( n47167 , n44318 , n39795 );
and ( n47168 , n44000 , n39793 );
nor ( n47169 , n47167 , n47168 );
xnor ( n47170 , n47169 , n39729 );
and ( n47171 , n44826 , n39665 );
and ( n47172 , n44347 , n39663 );
nor ( n47173 , n47171 , n47172 );
xnor ( n47174 , n47173 , n39608 );
and ( n47175 , n47170 , n47174 );
buf ( n47176 , n30372 );
not ( n47177 , n47176 );
and ( n47178 , n47174 , n47177 );
and ( n47179 , n47170 , n47177 );
or ( n47180 , n47175 , n47178 , n47179 );
and ( n47181 , n47165 , n47180 );
and ( n47182 , n47164 , n47180 );
or ( n47183 , n47166 , n47181 , n47182 );
and ( n47184 , n47161 , n47183 );
and ( n47185 , n47159 , n47183 );
or ( n47186 , n47162 , n47184 , n47185 );
and ( n47187 , n47156 , n47186 );
and ( n47188 , n47154 , n47186 );
or ( n47189 , n47157 , n47187 , n47188 );
and ( n47190 , n47151 , n47189 );
and ( n47191 , n47149 , n47189 );
or ( n47192 , n47152 , n47190 , n47191 );
and ( n47193 , n47147 , n47192 );
xor ( n47194 , n47018 , n47131 );
xor ( n47195 , n47194 , n47134 );
and ( n47196 , n47192 , n47195 );
and ( n47197 , n47147 , n47195 );
or ( n47198 , n47193 , n47196 , n47197 );
and ( n47199 , n47145 , n47198 );
xor ( n47200 , n47013 , n47015 );
xor ( n47201 , n47200 , n47137 );
and ( n47202 , n47198 , n47201 );
and ( n47203 , n47145 , n47201 );
or ( n47204 , n47199 , n47202 , n47203 );
and ( n47205 , n47142 , n47204 );
and ( n47206 , n47140 , n47204 );
or ( n47207 , n47143 , n47205 , n47206 );
and ( n47208 , n47010 , n47207 );
and ( n47209 , n47008 , n47207 );
or ( n47210 , n47011 , n47208 , n47209 );
and ( n47211 , n46836 , n47210 );
and ( n47212 , n46834 , n47210 );
or ( n47213 , n46837 , n47211 , n47212 );
and ( n47214 , n46657 , n47213 );
and ( n47215 , n46655 , n47213 );
or ( n47216 , n46658 , n47214 , n47215 );
and ( n47217 , n46494 , n47216 );
and ( n47218 , n46492 , n47216 );
or ( n47219 , n46495 , n47217 , n47218 );
and ( n47220 , n46490 , n47219 );
xor ( n47221 , n46490 , n47219 );
xor ( n47222 , n46492 , n46494 );
xor ( n47223 , n47222 , n47216 );
xor ( n47224 , n46655 , n46657 );
xor ( n47225 , n47224 , n47213 );
not ( n47226 , n47225 );
xor ( n47227 , n46834 , n46836 );
xor ( n47228 , n47227 , n47210 );
xor ( n47229 , n47008 , n47010 );
xor ( n47230 , n47229 , n47207 );
xor ( n47231 , n47140 , n47142 );
xor ( n47232 , n47231 , n47204 );
xor ( n47233 , n47145 , n47198 );
xor ( n47234 , n47233 , n47201 );
and ( n47235 , n41379 , n42079 );
and ( n47236 , n41091 , n42076 );
nor ( n47237 , n47235 , n47236 );
xnor ( n47238 , n47237 , n41370 );
and ( n47239 , n41735 , n41981 );
and ( n47240 , n41364 , n41979 );
nor ( n47241 , n47239 , n47240 );
xnor ( n47242 , n47241 , n41373 );
and ( n47243 , n47238 , n47242 );
and ( n47244 , n42149 , n41522 );
and ( n47245 , n41844 , n41520 );
nor ( n47246 , n47244 , n47245 );
xnor ( n47247 , n47246 , n41100 );
and ( n47248 , n47242 , n47247 );
and ( n47249 , n47238 , n47247 );
or ( n47250 , n47243 , n47248 , n47249 );
and ( n47251 , n42525 , n41230 );
and ( n47252 , n41828 , n41228 );
nor ( n47253 , n47251 , n47252 );
xnor ( n47254 , n47253 , n40981 );
and ( n47255 , n43040 , n40928 );
and ( n47256 , n42862 , n40926 );
nor ( n47257 , n47255 , n47256 );
xnor ( n47258 , n47257 , n40688 );
and ( n47259 , n47254 , n47258 );
and ( n47260 , n43322 , n40666 );
and ( n47261 , n43142 , n40664 );
nor ( n47262 , n47260 , n47261 );
xnor ( n47263 , n47262 , n40445 );
and ( n47264 , n47258 , n47263 );
and ( n47265 , n47254 , n47263 );
or ( n47266 , n47259 , n47264 , n47265 );
and ( n47267 , n47250 , n47266 );
and ( n47268 , n43524 , n40406 );
and ( n47269 , n43387 , n40404 );
nor ( n47270 , n47268 , n47269 );
xnor ( n47271 , n47270 , n40262 );
and ( n47272 , n43671 , n40168 );
and ( n47273 , n43549 , n40166 );
nor ( n47274 , n47272 , n47273 );
xnor ( n47275 , n47274 , n40059 );
and ( n47276 , n47271 , n47275 );
and ( n47277 , n43820 , n39984 );
and ( n47278 , n43679 , n39982 );
nor ( n47279 , n47277 , n47278 );
xnor ( n47280 , n47279 , n39865 );
and ( n47281 , n47275 , n47280 );
and ( n47282 , n47271 , n47280 );
or ( n47283 , n47276 , n47281 , n47282 );
and ( n47284 , n47266 , n47283 );
and ( n47285 , n47250 , n47283 );
or ( n47286 , n47267 , n47284 , n47285 );
and ( n47287 , n45171 , n39532 );
and ( n47288 , n45057 , n39530 );
nor ( n47289 , n47287 , n47288 );
xnor ( n47290 , n47289 , n39497 );
and ( n47291 , n46069 , n39384 );
and ( n47292 , n45754 , n39382 );
nor ( n47293 , n47291 , n47292 );
xnor ( n47294 , n47293 , n39367 );
and ( n47295 , n47290 , n47294 );
and ( n47296 , n46510 , n39335 );
and ( n47297 , n46159 , n39333 );
nor ( n47298 , n47296 , n47297 );
xnor ( n47299 , n47298 , n39300 );
and ( n47300 , n47294 , n47299 );
and ( n47301 , n47290 , n47299 );
or ( n47302 , n47295 , n47300 , n47301 );
xor ( n47303 , n47036 , n47040 );
xor ( n47304 , n47303 , n47045 );
and ( n47305 , n47302 , n47304 );
xor ( n47306 , n47056 , n47060 );
xor ( n47307 , n47306 , n47065 );
and ( n47308 , n47304 , n47307 );
and ( n47309 , n47302 , n47307 );
or ( n47310 , n47305 , n47308 , n47309 );
and ( n47311 , n47286 , n47310 );
xor ( n47312 , n47022 , n47031 );
xor ( n47313 , n47312 , n47048 );
and ( n47314 , n47310 , n47313 );
and ( n47315 , n47286 , n47313 );
or ( n47316 , n47311 , n47314 , n47315 );
xor ( n47317 , n47020 , n47051 );
xor ( n47318 , n47317 , n47104 );
and ( n47319 , n47316 , n47318 );
xor ( n47320 , n47117 , n47119 );
xor ( n47321 , n47320 , n47122 );
and ( n47322 , n47318 , n47321 );
and ( n47323 , n47316 , n47321 );
or ( n47324 , n47319 , n47322 , n47323 );
xor ( n47325 , n47107 , n47125 );
xor ( n47326 , n47325 , n47128 );
and ( n47327 , n47324 , n47326 );
xor ( n47328 , n47068 , n47084 );
xor ( n47329 , n47328 , n47101 );
xor ( n47330 , n47109 , n47111 );
xor ( n47331 , n47330 , n47114 );
and ( n47332 , n47329 , n47331 );
xor ( n47333 , n47072 , n47076 );
xor ( n47334 , n47333 , n47081 );
xor ( n47335 , n47089 , n47093 );
xor ( n47336 , n47335 , n47098 );
and ( n47337 , n47334 , n47336 );
xor ( n47338 , n47170 , n47174 );
xor ( n47339 , n47338 , n47177 );
and ( n47340 , n41364 , n42079 );
and ( n47341 , n41379 , n42076 );
nor ( n47342 , n47340 , n47341 );
xnor ( n47343 , n47342 , n41370 );
and ( n47344 , n41844 , n41981 );
and ( n47345 , n41735 , n41979 );
nor ( n47346 , n47344 , n47345 );
xnor ( n47347 , n47346 , n41373 );
and ( n47348 , n47343 , n47347 );
and ( n47349 , n41828 , n41522 );
and ( n47350 , n42149 , n41520 );
nor ( n47351 , n47349 , n47350 );
xnor ( n47352 , n47351 , n41100 );
and ( n47353 , n47347 , n47352 );
and ( n47354 , n47343 , n47352 );
or ( n47355 , n47348 , n47353 , n47354 );
and ( n47356 , n47339 , n47355 );
and ( n47357 , n42862 , n41230 );
and ( n47358 , n42525 , n41228 );
nor ( n47359 , n47357 , n47358 );
xnor ( n47360 , n47359 , n40981 );
and ( n47361 , n43142 , n40928 );
and ( n47362 , n43040 , n40926 );
nor ( n47363 , n47361 , n47362 );
xnor ( n47364 , n47363 , n40688 );
and ( n47365 , n47360 , n47364 );
and ( n47366 , n43387 , n40666 );
and ( n47367 , n43322 , n40664 );
nor ( n47368 , n47366 , n47367 );
xnor ( n47369 , n47368 , n40445 );
and ( n47370 , n47364 , n47369 );
and ( n47371 , n47360 , n47369 );
or ( n47372 , n47365 , n47370 , n47371 );
and ( n47373 , n47355 , n47372 );
and ( n47374 , n47339 , n47372 );
or ( n47375 , n47356 , n47373 , n47374 );
and ( n47376 , n47336 , n47375 );
and ( n47377 , n47334 , n47375 );
or ( n47378 , n47337 , n47376 , n47377 );
and ( n47379 , n47331 , n47378 );
and ( n47380 , n47329 , n47378 );
or ( n47381 , n47332 , n47379 , n47380 );
and ( n47382 , n43549 , n40406 );
and ( n47383 , n43524 , n40404 );
nor ( n47384 , n47382 , n47383 );
xnor ( n47385 , n47384 , n40262 );
and ( n47386 , n43679 , n40168 );
and ( n47387 , n43671 , n40166 );
nor ( n47388 , n47386 , n47387 );
xnor ( n47389 , n47388 , n40059 );
and ( n47390 , n47385 , n47389 );
and ( n47391 , n44000 , n39984 );
and ( n47392 , n43820 , n39982 );
nor ( n47393 , n47391 , n47392 );
xnor ( n47394 , n47393 , n39865 );
and ( n47395 , n47389 , n47394 );
and ( n47396 , n47385 , n47394 );
or ( n47397 , n47390 , n47395 , n47396 );
and ( n47398 , n44347 , n39795 );
and ( n47399 , n44318 , n39793 );
nor ( n47400 , n47398 , n47399 );
xnor ( n47401 , n47400 , n39729 );
and ( n47402 , n45057 , n39665 );
and ( n47403 , n44826 , n39663 );
nor ( n47404 , n47402 , n47403 );
xnor ( n47405 , n47404 , n39608 );
and ( n47406 , n47401 , n47405 );
and ( n47407 , n45754 , n39532 );
and ( n47408 , n45171 , n39530 );
nor ( n47409 , n47407 , n47408 );
xnor ( n47410 , n47409 , n39497 );
and ( n47411 , n47405 , n47410 );
and ( n47412 , n47401 , n47410 );
or ( n47413 , n47406 , n47411 , n47412 );
and ( n47414 , n47397 , n47413 );
and ( n47415 , n46159 , n39384 );
and ( n47416 , n46069 , n39382 );
nor ( n47417 , n47415 , n47416 );
xnor ( n47418 , n47417 , n39367 );
and ( n47419 , n46676 , n39335 );
and ( n47420 , n46510 , n39333 );
nor ( n47421 , n47419 , n47420 );
xnor ( n47422 , n47421 , n39300 );
and ( n47423 , n47418 , n47422 );
and ( n47424 , n46948 , n39258 );
and ( n47425 , n46777 , n39256 );
nor ( n47426 , n47424 , n47425 );
xnor ( n47427 , n47426 , n39215 );
and ( n47428 , n47422 , n47427 );
and ( n47429 , n47418 , n47427 );
or ( n47430 , n47423 , n47428 , n47429 );
and ( n47431 , n47413 , n47430 );
and ( n47432 , n47397 , n47430 );
or ( n47433 , n47414 , n47431 , n47432 );
xor ( n47434 , n47238 , n47242 );
xor ( n47435 , n47434 , n47247 );
xor ( n47436 , n47254 , n47258 );
xor ( n47437 , n47436 , n47263 );
and ( n47438 , n47435 , n47437 );
xor ( n47439 , n47271 , n47275 );
xor ( n47440 , n47439 , n47280 );
and ( n47441 , n47437 , n47440 );
and ( n47442 , n47435 , n47440 );
or ( n47443 , n47438 , n47441 , n47442 );
and ( n47444 , n47433 , n47443 );
xor ( n47445 , n47164 , n47165 );
xor ( n47446 , n47445 , n47180 );
and ( n47447 , n47443 , n47446 );
and ( n47448 , n47433 , n47446 );
or ( n47449 , n47444 , n47447 , n47448 );
xor ( n47450 , n47159 , n47161 );
xor ( n47451 , n47450 , n47183 );
and ( n47452 , n47449 , n47451 );
xor ( n47453 , n47286 , n47310 );
xor ( n47454 , n47453 , n47313 );
and ( n47455 , n47451 , n47454 );
and ( n47456 , n47449 , n47454 );
or ( n47457 , n47452 , n47455 , n47456 );
and ( n47458 , n47381 , n47457 );
xor ( n47459 , n47154 , n47156 );
xor ( n47460 , n47459 , n47186 );
and ( n47461 , n47457 , n47460 );
and ( n47462 , n47381 , n47460 );
or ( n47463 , n47458 , n47461 , n47462 );
and ( n47464 , n47326 , n47463 );
and ( n47465 , n47324 , n47463 );
or ( n47466 , n47327 , n47464 , n47465 );
xor ( n47467 , n47147 , n47192 );
xor ( n47468 , n47467 , n47195 );
and ( n47469 , n47466 , n47468 );
xor ( n47470 , n47149 , n47151 );
xor ( n47471 , n47470 , n47189 );
xor ( n47472 , n47316 , n47318 );
xor ( n47473 , n47472 , n47321 );
xor ( n47474 , n47250 , n47266 );
xor ( n47475 , n47474 , n47283 );
xor ( n47476 , n47302 , n47304 );
xor ( n47477 , n47476 , n47307 );
and ( n47478 , n47475 , n47477 );
xor ( n47479 , n47290 , n47294 );
xor ( n47480 , n47479 , n47299 );
buf ( n47481 , n30373 );
not ( n47482 , n47481 );
and ( n47483 , n44318 , n39984 );
and ( n47484 , n44000 , n39982 );
nor ( n47485 , n47483 , n47484 );
xnor ( n47486 , n47485 , n39865 );
and ( n47487 , n44826 , n39795 );
and ( n47488 , n44347 , n39793 );
nor ( n47489 , n47487 , n47488 );
xnor ( n47490 , n47489 , n39729 );
and ( n47491 , n47486 , n47490 );
buf ( n47492 , n30374 );
not ( n47493 , n47492 );
and ( n47494 , n47490 , n47493 );
and ( n47495 , n47486 , n47493 );
or ( n47496 , n47491 , n47494 , n47495 );
and ( n47497 , n47482 , n47496 );
and ( n47498 , n41735 , n42079 );
and ( n47499 , n41364 , n42076 );
nor ( n47500 , n47498 , n47499 );
xnor ( n47501 , n47500 , n41370 );
and ( n47502 , n42149 , n41981 );
and ( n47503 , n41844 , n41979 );
nor ( n47504 , n47502 , n47503 );
xnor ( n47505 , n47504 , n41373 );
and ( n47506 , n47501 , n47505 );
and ( n47507 , n42525 , n41522 );
and ( n47508 , n41828 , n41520 );
nor ( n47509 , n47507 , n47508 );
xnor ( n47510 , n47509 , n41100 );
and ( n47511 , n47505 , n47510 );
and ( n47512 , n47501 , n47510 );
or ( n47513 , n47506 , n47511 , n47512 );
and ( n47514 , n47496 , n47513 );
and ( n47515 , n47482 , n47513 );
or ( n47516 , n47497 , n47514 , n47515 );
and ( n47517 , n47480 , n47516 );
and ( n47518 , n43040 , n41230 );
and ( n47519 , n42862 , n41228 );
nor ( n47520 , n47518 , n47519 );
xnor ( n47521 , n47520 , n40981 );
and ( n47522 , n43322 , n40928 );
and ( n47523 , n43142 , n40926 );
nor ( n47524 , n47522 , n47523 );
xnor ( n47525 , n47524 , n40688 );
and ( n47526 , n47521 , n47525 );
and ( n47527 , n43524 , n40666 );
and ( n47528 , n43387 , n40664 );
nor ( n47529 , n47527 , n47528 );
xnor ( n47530 , n47529 , n40445 );
and ( n47531 , n47525 , n47530 );
and ( n47532 , n47521 , n47530 );
or ( n47533 , n47526 , n47531 , n47532 );
and ( n47534 , n43671 , n40406 );
and ( n47535 , n43549 , n40404 );
nor ( n47536 , n47534 , n47535 );
xnor ( n47537 , n47536 , n40262 );
and ( n47538 , n43820 , n40168 );
and ( n47539 , n43679 , n40166 );
nor ( n47540 , n47538 , n47539 );
xnor ( n47541 , n47540 , n40059 );
and ( n47542 , n47537 , n47541 );
and ( n47543 , n45171 , n39665 );
and ( n47544 , n45057 , n39663 );
nor ( n47545 , n47543 , n47544 );
xnor ( n47546 , n47545 , n39608 );
and ( n47547 , n47541 , n47546 );
and ( n47548 , n47537 , n47546 );
or ( n47549 , n47542 , n47547 , n47548 );
and ( n47550 , n47533 , n47549 );
and ( n47551 , n46069 , n39532 );
and ( n47552 , n45754 , n39530 );
nor ( n47553 , n47551 , n47552 );
xnor ( n47554 , n47553 , n39497 );
and ( n47555 , n46510 , n39384 );
and ( n47556 , n46159 , n39382 );
nor ( n47557 , n47555 , n47556 );
xnor ( n47558 , n47557 , n39367 );
and ( n47559 , n47554 , n47558 );
and ( n47560 , n46777 , n39335 );
and ( n47561 , n46676 , n39333 );
nor ( n47562 , n47560 , n47561 );
xnor ( n47563 , n47562 , n39300 );
and ( n47564 , n47558 , n47563 );
and ( n47565 , n47554 , n47563 );
or ( n47566 , n47559 , n47564 , n47565 );
and ( n47567 , n47549 , n47566 );
and ( n47568 , n47533 , n47566 );
or ( n47569 , n47550 , n47567 , n47568 );
and ( n47570 , n47516 , n47569 );
and ( n47571 , n47480 , n47569 );
or ( n47572 , n47517 , n47570 , n47571 );
and ( n47573 , n47477 , n47572 );
and ( n47574 , n47475 , n47572 );
or ( n47575 , n47478 , n47573 , n47574 );
xor ( n47576 , n47343 , n47347 );
xor ( n47577 , n47576 , n47352 );
xor ( n47578 , n47360 , n47364 );
xor ( n47579 , n47578 , n47369 );
and ( n47580 , n47577 , n47579 );
xor ( n47581 , n47385 , n47389 );
xor ( n47582 , n47581 , n47394 );
and ( n47583 , n47579 , n47582 );
and ( n47584 , n47577 , n47582 );
or ( n47585 , n47580 , n47583 , n47584 );
xor ( n47586 , n47339 , n47355 );
xor ( n47587 , n47586 , n47372 );
and ( n47588 , n47585 , n47587 );
xor ( n47589 , n47397 , n47413 );
xor ( n47590 , n47589 , n47430 );
and ( n47591 , n47587 , n47590 );
and ( n47592 , n47585 , n47590 );
or ( n47593 , n47588 , n47591 , n47592 );
xor ( n47594 , n47334 , n47336 );
xor ( n47595 , n47594 , n47375 );
and ( n47596 , n47593 , n47595 );
xor ( n47597 , n47433 , n47443 );
xor ( n47598 , n47597 , n47446 );
and ( n47599 , n47595 , n47598 );
and ( n47600 , n47593 , n47598 );
or ( n47601 , n47596 , n47599 , n47600 );
and ( n47602 , n47575 , n47601 );
xor ( n47603 , n47329 , n47331 );
xor ( n47604 , n47603 , n47378 );
and ( n47605 , n47601 , n47604 );
and ( n47606 , n47575 , n47604 );
or ( n47607 , n47602 , n47605 , n47606 );
and ( n47608 , n47473 , n47607 );
xor ( n47609 , n47381 , n47457 );
xor ( n47610 , n47609 , n47460 );
and ( n47611 , n47607 , n47610 );
and ( n47612 , n47473 , n47610 );
or ( n47613 , n47608 , n47611 , n47612 );
and ( n47614 , n47471 , n47613 );
xor ( n47615 , n47324 , n47326 );
xor ( n47616 , n47615 , n47463 );
and ( n47617 , n47613 , n47616 );
and ( n47618 , n47471 , n47616 );
or ( n47619 , n47614 , n47617 , n47618 );
and ( n47620 , n47468 , n47619 );
and ( n47621 , n47466 , n47619 );
or ( n47622 , n47469 , n47620 , n47621 );
or ( n47623 , n47234 , n47622 );
or ( n47624 , n47232 , n47623 );
and ( n47625 , n47230 , n47624 );
xor ( n47626 , n47230 , n47624 );
xnor ( n47627 , n47232 , n47623 );
xnor ( n47628 , n47234 , n47622 );
xor ( n47629 , n47466 , n47468 );
xor ( n47630 , n47629 , n47619 );
xor ( n47631 , n47471 , n47613 );
xor ( n47632 , n47631 , n47616 );
xor ( n47633 , n47449 , n47451 );
xor ( n47634 , n47633 , n47454 );
xor ( n47635 , n47435 , n47437 );
xor ( n47636 , n47635 , n47440 );
xor ( n47637 , n47401 , n47405 );
xor ( n47638 , n47637 , n47410 );
xor ( n47639 , n47418 , n47422 );
xor ( n47640 , n47639 , n47427 );
and ( n47641 , n47638 , n47640 );
xor ( n47642 , n39050 , n39092 );
buf ( n47643 , n47642 );
buf ( n47644 , n47643 );
buf ( n47645 , n47644 );
and ( n47646 , n47645 , n39258 );
and ( n47647 , n46948 , n39256 );
nor ( n47648 , n47646 , n47647 );
xnor ( n47649 , n47648 , n39215 );
xor ( n47650 , n47486 , n47490 );
xor ( n47651 , n47650 , n47493 );
and ( n47652 , n47649 , n47651 );
and ( n47653 , n41844 , n42079 );
and ( n47654 , n41735 , n42076 );
nor ( n47655 , n47653 , n47654 );
xnor ( n47656 , n47655 , n41370 );
and ( n47657 , n41828 , n41981 );
and ( n47658 , n42149 , n41979 );
nor ( n47659 , n47657 , n47658 );
xnor ( n47660 , n47659 , n41373 );
and ( n47661 , n47656 , n47660 );
and ( n47662 , n42862 , n41522 );
and ( n47663 , n42525 , n41520 );
nor ( n47664 , n47662 , n47663 );
xnor ( n47665 , n47664 , n41100 );
and ( n47666 , n47660 , n47665 );
and ( n47667 , n47656 , n47665 );
or ( n47668 , n47661 , n47666 , n47667 );
and ( n47669 , n47651 , n47668 );
and ( n47670 , n47649 , n47668 );
or ( n47671 , n47652 , n47669 , n47670 );
and ( n47672 , n47640 , n47671 );
and ( n47673 , n47638 , n47671 );
or ( n47674 , n47641 , n47672 , n47673 );
and ( n47675 , n47636 , n47674 );
and ( n47676 , n43142 , n41230 );
and ( n47677 , n43040 , n41228 );
nor ( n47678 , n47676 , n47677 );
xnor ( n47679 , n47678 , n40981 );
and ( n47680 , n43387 , n40928 );
and ( n47681 , n43322 , n40926 );
nor ( n47682 , n47680 , n47681 );
xnor ( n47683 , n47682 , n40688 );
and ( n47684 , n47679 , n47683 );
and ( n47685 , n43549 , n40666 );
and ( n47686 , n43524 , n40664 );
nor ( n47687 , n47685 , n47686 );
xnor ( n47688 , n47687 , n40445 );
and ( n47689 , n47683 , n47688 );
and ( n47690 , n47679 , n47688 );
or ( n47691 , n47684 , n47689 , n47690 );
and ( n47692 , n43679 , n40406 );
and ( n47693 , n43671 , n40404 );
nor ( n47694 , n47692 , n47693 );
xnor ( n47695 , n47694 , n40262 );
and ( n47696 , n44000 , n40168 );
and ( n47697 , n43820 , n40166 );
nor ( n47698 , n47696 , n47697 );
xnor ( n47699 , n47698 , n40059 );
and ( n47700 , n47695 , n47699 );
and ( n47701 , n44347 , n39984 );
and ( n47702 , n44318 , n39982 );
nor ( n47703 , n47701 , n47702 );
xnor ( n47704 , n47703 , n39865 );
and ( n47705 , n47699 , n47704 );
and ( n47706 , n47695 , n47704 );
or ( n47707 , n47700 , n47705 , n47706 );
and ( n47708 , n47691 , n47707 );
and ( n47709 , n45057 , n39795 );
and ( n47710 , n44826 , n39793 );
nor ( n47711 , n47709 , n47710 );
xnor ( n47712 , n47711 , n39729 );
and ( n47713 , n45754 , n39665 );
and ( n47714 , n45171 , n39663 );
nor ( n47715 , n47713 , n47714 );
xnor ( n47716 , n47715 , n39608 );
and ( n47717 , n47712 , n47716 );
and ( n47718 , n46159 , n39532 );
and ( n47719 , n46069 , n39530 );
nor ( n47720 , n47718 , n47719 );
xnor ( n47721 , n47720 , n39497 );
and ( n47722 , n47716 , n47721 );
and ( n47723 , n47712 , n47721 );
or ( n47724 , n47717 , n47722 , n47723 );
and ( n47725 , n47707 , n47724 );
and ( n47726 , n47691 , n47724 );
or ( n47727 , n47708 , n47725 , n47726 );
and ( n47728 , n46676 , n39384 );
and ( n47729 , n46510 , n39382 );
nor ( n47730 , n47728 , n47729 );
xnor ( n47731 , n47730 , n39367 );
and ( n47732 , n46948 , n39335 );
and ( n47733 , n46777 , n39333 );
nor ( n47734 , n47732 , n47733 );
xnor ( n47735 , n47734 , n39300 );
and ( n47736 , n47731 , n47735 );
buf ( n47737 , n30375 );
not ( n47738 , n47737 );
and ( n47739 , n47735 , n47738 );
and ( n47740 , n47731 , n47738 );
or ( n47741 , n47736 , n47739 , n47740 );
xor ( n47742 , n47501 , n47505 );
xor ( n47743 , n47742 , n47510 );
and ( n47744 , n47741 , n47743 );
xor ( n47745 , n47521 , n47525 );
xor ( n47746 , n47745 , n47530 );
and ( n47747 , n47743 , n47746 );
and ( n47748 , n47741 , n47746 );
or ( n47749 , n47744 , n47747 , n47748 );
and ( n47750 , n47727 , n47749 );
xor ( n47751 , n47482 , n47496 );
xor ( n47752 , n47751 , n47513 );
and ( n47753 , n47749 , n47752 );
and ( n47754 , n47727 , n47752 );
or ( n47755 , n47750 , n47753 , n47754 );
and ( n47756 , n47674 , n47755 );
and ( n47757 , n47636 , n47755 );
or ( n47758 , n47675 , n47756 , n47757 );
xor ( n47759 , n47475 , n47477 );
xor ( n47760 , n47759 , n47572 );
and ( n47761 , n47758 , n47760 );
xor ( n47762 , n47593 , n47595 );
xor ( n47763 , n47762 , n47598 );
and ( n47764 , n47760 , n47763 );
and ( n47765 , n47758 , n47763 );
or ( n47766 , n47761 , n47764 , n47765 );
and ( n47767 , n47634 , n47766 );
xor ( n47768 , n47575 , n47601 );
xor ( n47769 , n47768 , n47604 );
and ( n47770 , n47766 , n47769 );
and ( n47771 , n47634 , n47769 );
or ( n47772 , n47767 , n47770 , n47771 );
xor ( n47773 , n47473 , n47607 );
xor ( n47774 , n47773 , n47610 );
and ( n47775 , n47772 , n47774 );
xor ( n47776 , n47634 , n47766 );
xor ( n47777 , n47776 , n47769 );
xor ( n47778 , n47480 , n47516 );
xor ( n47779 , n47778 , n47569 );
xor ( n47780 , n47585 , n47587 );
xor ( n47781 , n47780 , n47590 );
and ( n47782 , n47779 , n47781 );
xor ( n47783 , n47533 , n47549 );
xor ( n47784 , n47783 , n47566 );
xor ( n47785 , n47577 , n47579 );
xor ( n47786 , n47785 , n47582 );
and ( n47787 , n47784 , n47786 );
xor ( n47788 , n47537 , n47541 );
xor ( n47789 , n47788 , n47546 );
xor ( n47790 , n47554 , n47558 );
xor ( n47791 , n47790 , n47563 );
and ( n47792 , n47789 , n47791 );
and ( n47793 , n44318 , n40168 );
and ( n47794 , n44000 , n40166 );
nor ( n47795 , n47793 , n47794 );
xnor ( n47796 , n47795 , n40059 );
and ( n47797 , n44826 , n39984 );
and ( n47798 , n44347 , n39982 );
nor ( n47799 , n47797 , n47798 );
xnor ( n47800 , n47799 , n39865 );
and ( n47801 , n47796 , n47800 );
buf ( n47802 , n30376 );
not ( n47803 , n47802 );
and ( n47804 , n47800 , n47803 );
and ( n47805 , n47796 , n47803 );
or ( n47806 , n47801 , n47804 , n47805 );
and ( n47807 , n43322 , n41230 );
and ( n47808 , n43142 , n41228 );
nor ( n47809 , n47807 , n47808 );
xnor ( n47810 , n47809 , n40981 );
and ( n47811 , n43524 , n40928 );
and ( n47812 , n43387 , n40926 );
nor ( n47813 , n47811 , n47812 );
xnor ( n47814 , n47813 , n40688 );
or ( n47815 , n47810 , n47814 );
and ( n47816 , n47806 , n47815 );
and ( n47817 , n42149 , n42079 );
and ( n47818 , n41844 , n42076 );
nor ( n47819 , n47817 , n47818 );
xnor ( n47820 , n47819 , n41370 );
and ( n47821 , n42525 , n41981 );
and ( n47822 , n41828 , n41979 );
nor ( n47823 , n47821 , n47822 );
xnor ( n47824 , n47823 , n41373 );
and ( n47825 , n47820 , n47824 );
and ( n47826 , n43040 , n41522 );
and ( n47827 , n42862 , n41520 );
nor ( n47828 , n47826 , n47827 );
xnor ( n47829 , n47828 , n41100 );
and ( n47830 , n47824 , n47829 );
and ( n47831 , n47820 , n47829 );
or ( n47832 , n47825 , n47830 , n47831 );
and ( n47833 , n47815 , n47832 );
and ( n47834 , n47806 , n47832 );
or ( n47835 , n47816 , n47833 , n47834 );
and ( n47836 , n47791 , n47835 );
and ( n47837 , n47789 , n47835 );
or ( n47838 , n47792 , n47836 , n47837 );
and ( n47839 , n47786 , n47838 );
and ( n47840 , n47784 , n47838 );
or ( n47841 , n47787 , n47839 , n47840 );
and ( n47842 , n47781 , n47841 );
and ( n47843 , n47779 , n47841 );
or ( n47844 , n47782 , n47842 , n47843 );
xor ( n47845 , n47758 , n47760 );
xor ( n47846 , n47845 , n47763 );
and ( n47847 , n47844 , n47846 );
and ( n47848 , n43671 , n40666 );
and ( n47849 , n43549 , n40664 );
nor ( n47850 , n47848 , n47849 );
xnor ( n47851 , n47850 , n40445 );
and ( n47852 , n43820 , n40406 );
and ( n47853 , n43679 , n40404 );
nor ( n47854 , n47852 , n47853 );
xnor ( n47855 , n47854 , n40262 );
and ( n47856 , n47851 , n47855 );
and ( n47857 , n45171 , n39795 );
and ( n47858 , n45057 , n39793 );
nor ( n47859 , n47857 , n47858 );
xnor ( n47860 , n47859 , n39729 );
and ( n47861 , n47855 , n47860 );
and ( n47862 , n47851 , n47860 );
or ( n47863 , n47856 , n47861 , n47862 );
and ( n47864 , n46069 , n39665 );
and ( n47865 , n45754 , n39663 );
nor ( n47866 , n47864 , n47865 );
xnor ( n47867 , n47866 , n39608 );
and ( n47868 , n46510 , n39532 );
and ( n47869 , n46159 , n39530 );
nor ( n47870 , n47868 , n47869 );
xnor ( n47871 , n47870 , n39497 );
and ( n47872 , n47867 , n47871 );
and ( n47873 , n46777 , n39384 );
and ( n47874 , n46676 , n39382 );
nor ( n47875 , n47873 , n47874 );
xnor ( n47876 , n47875 , n39367 );
and ( n47877 , n47871 , n47876 );
and ( n47878 , n47867 , n47876 );
or ( n47879 , n47872 , n47877 , n47878 );
and ( n47880 , n47863 , n47879 );
xor ( n47881 , n47656 , n47660 );
xor ( n47882 , n47881 , n47665 );
and ( n47883 , n47879 , n47882 );
and ( n47884 , n47863 , n47882 );
or ( n47885 , n47880 , n47883 , n47884 );
xor ( n47886 , n47679 , n47683 );
xor ( n47887 , n47886 , n47688 );
xor ( n47888 , n47695 , n47699 );
xor ( n47889 , n47888 , n47704 );
and ( n47890 , n47887 , n47889 );
xor ( n47891 , n47712 , n47716 );
xor ( n47892 , n47891 , n47721 );
and ( n47893 , n47889 , n47892 );
and ( n47894 , n47887 , n47892 );
or ( n47895 , n47890 , n47893 , n47894 );
and ( n47896 , n47885 , n47895 );
xor ( n47897 , n47649 , n47651 );
xor ( n47898 , n47897 , n47668 );
and ( n47899 , n47895 , n47898 );
and ( n47900 , n47885 , n47898 );
or ( n47901 , n47896 , n47899 , n47900 );
xor ( n47902 , n47638 , n47640 );
xor ( n47903 , n47902 , n47671 );
and ( n47904 , n47901 , n47903 );
xor ( n47905 , n47727 , n47749 );
xor ( n47906 , n47905 , n47752 );
and ( n47907 , n47903 , n47906 );
and ( n47908 , n47901 , n47906 );
or ( n47909 , n47904 , n47907 , n47908 );
xor ( n47910 , n47636 , n47674 );
xor ( n47911 , n47910 , n47755 );
and ( n47912 , n47909 , n47911 );
xor ( n47913 , n47691 , n47707 );
xor ( n47914 , n47913 , n47724 );
xor ( n47915 , n47741 , n47743 );
xor ( n47916 , n47915 , n47746 );
and ( n47917 , n47914 , n47916 );
xor ( n47918 , n47731 , n47735 );
xor ( n47919 , n47918 , n47738 );
and ( n47920 , n47645 , n39335 );
and ( n47921 , n46948 , n39333 );
nor ( n47922 , n47920 , n47921 );
xnor ( n47923 , n47922 , n39300 );
xor ( n47924 , n39067 , n39089 );
buf ( n47925 , n47924 );
buf ( n47926 , n47925 );
buf ( n47927 , n47926 );
and ( n47928 , n47927 , n39258 );
xor ( n47929 , n39052 , n39091 );
buf ( n47930 , n47929 );
buf ( n47931 , n47930 );
buf ( n47932 , n47931 );
and ( n47933 , n47932 , n39256 );
nor ( n47934 , n47928 , n47933 );
xnor ( n47935 , n47934 , n39215 );
and ( n47936 , n47923 , n47935 );
xor ( n47937 , n47796 , n47800 );
xor ( n47938 , n47937 , n47803 );
and ( n47939 , n47935 , n47938 );
and ( n47940 , n47923 , n47938 );
or ( n47941 , n47936 , n47939 , n47940 );
and ( n47942 , n47919 , n47941 );
xnor ( n47943 , n47810 , n47814 );
and ( n47944 , n45057 , n39984 );
and ( n47945 , n44826 , n39982 );
nor ( n47946 , n47944 , n47945 );
xnor ( n47947 , n47946 , n39865 );
buf ( n47948 , n30377 );
not ( n47949 , n47948 );
and ( n47950 , n47947 , n47949 );
and ( n47951 , n47943 , n47950 );
and ( n47952 , n41828 , n42079 );
and ( n47953 , n42149 , n42076 );
nor ( n47954 , n47952 , n47953 );
xnor ( n47955 , n47954 , n41370 );
and ( n47956 , n42862 , n41981 );
and ( n47957 , n42525 , n41979 );
nor ( n47958 , n47956 , n47957 );
xnor ( n47959 , n47958 , n41373 );
and ( n47960 , n47955 , n47959 );
and ( n47961 , n43142 , n41522 );
and ( n47962 , n43040 , n41520 );
nor ( n47963 , n47961 , n47962 );
xnor ( n47964 , n47963 , n41100 );
and ( n47965 , n47959 , n47964 );
and ( n47966 , n47955 , n47964 );
or ( n47967 , n47960 , n47965 , n47966 );
and ( n47968 , n47950 , n47967 );
and ( n47969 , n47943 , n47967 );
or ( n47970 , n47951 , n47968 , n47969 );
and ( n47971 , n47941 , n47970 );
and ( n47972 , n47919 , n47970 );
or ( n47973 , n47942 , n47971 , n47972 );
and ( n47974 , n47916 , n47973 );
and ( n47975 , n47914 , n47973 );
or ( n47976 , n47917 , n47974 , n47975 );
and ( n47977 , n43387 , n41230 );
and ( n47978 , n43322 , n41228 );
nor ( n47979 , n47977 , n47978 );
xnor ( n47980 , n47979 , n40981 );
and ( n47981 , n43549 , n40928 );
and ( n47982 , n43524 , n40926 );
nor ( n47983 , n47981 , n47982 );
xnor ( n47984 , n47983 , n40688 );
and ( n47985 , n47980 , n47984 );
and ( n47986 , n43679 , n40666 );
and ( n47987 , n43671 , n40664 );
nor ( n47988 , n47986 , n47987 );
xnor ( n47989 , n47988 , n40445 );
and ( n47990 , n47984 , n47989 );
and ( n47991 , n47980 , n47989 );
or ( n47992 , n47985 , n47990 , n47991 );
and ( n47993 , n44000 , n40406 );
and ( n47994 , n43820 , n40404 );
nor ( n47995 , n47993 , n47994 );
xnor ( n47996 , n47995 , n40262 );
and ( n47997 , n44347 , n40168 );
and ( n47998 , n44318 , n40166 );
nor ( n47999 , n47997 , n47998 );
xnor ( n48000 , n47999 , n40059 );
and ( n48001 , n47996 , n48000 );
and ( n48002 , n45754 , n39795 );
and ( n48003 , n45171 , n39793 );
nor ( n48004 , n48002 , n48003 );
xnor ( n48005 , n48004 , n39729 );
and ( n48006 , n48000 , n48005 );
and ( n48007 , n47996 , n48005 );
or ( n48008 , n48001 , n48006 , n48007 );
and ( n48009 , n47992 , n48008 );
and ( n48010 , n46159 , n39665 );
and ( n48011 , n46069 , n39663 );
nor ( n48012 , n48010 , n48011 );
xnor ( n48013 , n48012 , n39608 );
and ( n48014 , n46676 , n39532 );
and ( n48015 , n46510 , n39530 );
nor ( n48016 , n48014 , n48015 );
xnor ( n48017 , n48016 , n39497 );
and ( n48018 , n48013 , n48017 );
and ( n48019 , n46948 , n39384 );
and ( n48020 , n46777 , n39382 );
nor ( n48021 , n48019 , n48020 );
xnor ( n48022 , n48021 , n39367 );
and ( n48023 , n48017 , n48022 );
and ( n48024 , n48013 , n48022 );
or ( n48025 , n48018 , n48023 , n48024 );
and ( n48026 , n48008 , n48025 );
and ( n48027 , n47992 , n48025 );
or ( n48028 , n48009 , n48026 , n48027 );
xor ( n48029 , n47820 , n47824 );
xor ( n48030 , n48029 , n47829 );
xor ( n48031 , n47851 , n47855 );
xor ( n48032 , n48031 , n47860 );
and ( n48033 , n48030 , n48032 );
xor ( n48034 , n47867 , n47871 );
xor ( n48035 , n48034 , n47876 );
and ( n48036 , n48032 , n48035 );
and ( n48037 , n48030 , n48035 );
or ( n48038 , n48033 , n48036 , n48037 );
and ( n48039 , n48028 , n48038 );
xor ( n48040 , n47806 , n47815 );
xor ( n48041 , n48040 , n47832 );
and ( n48042 , n48038 , n48041 );
and ( n48043 , n48028 , n48041 );
or ( n48044 , n48039 , n48042 , n48043 );
xor ( n48045 , n47789 , n47791 );
xor ( n48046 , n48045 , n47835 );
and ( n48047 , n48044 , n48046 );
xor ( n48048 , n47885 , n47895 );
xor ( n48049 , n48048 , n47898 );
and ( n48050 , n48046 , n48049 );
and ( n48051 , n48044 , n48049 );
or ( n48052 , n48047 , n48050 , n48051 );
and ( n48053 , n47976 , n48052 );
xor ( n48054 , n47784 , n47786 );
xor ( n48055 , n48054 , n47838 );
and ( n48056 , n48052 , n48055 );
and ( n48057 , n47976 , n48055 );
or ( n48058 , n48053 , n48056 , n48057 );
and ( n48059 , n47911 , n48058 );
and ( n48060 , n47909 , n48058 );
or ( n48061 , n47912 , n48059 , n48060 );
and ( n48062 , n47846 , n48061 );
and ( n48063 , n47844 , n48061 );
or ( n48064 , n47847 , n48062 , n48063 );
and ( n48065 , n47777 , n48064 );
xor ( n48066 , n39081 , n39083 );
buf ( n48067 , n48066 );
buf ( n48068 , n48067 );
buf ( n48069 , n48068 );
and ( n48070 , n48069 , n39192 );
not ( n48071 , n48070 );
and ( n48072 , n48071 , n39199 );
and ( n48073 , n48069 , n39194 );
xor ( n48074 , n39080 , n39084 );
buf ( n48075 , n48074 );
buf ( n48076 , n48075 );
buf ( n48077 , n48076 );
and ( n48078 , n48077 , n39192 );
nor ( n48079 , n48073 , n48078 );
xnor ( n48080 , n48079 , n39199 );
and ( n48081 , n48072 , n48080 );
and ( n48082 , n48077 , n39194 );
xor ( n48083 , n39075 , n39086 );
buf ( n48084 , n48083 );
buf ( n48085 , n48084 );
buf ( n48086 , n48085 );
and ( n48087 , n48086 , n39192 );
nor ( n48088 , n48082 , n48087 );
xnor ( n48089 , n48088 , n39199 );
and ( n48090 , n48081 , n48089 );
and ( n48091 , n48069 , n39186 );
and ( n48092 , n48089 , n48091 );
and ( n48093 , n48081 , n48091 );
or ( n48094 , n48090 , n48092 , n48093 );
and ( n48095 , n48086 , n39194 );
xor ( n48096 , n39074 , n39087 );
buf ( n48097 , n48096 );
buf ( n48098 , n48097 );
buf ( n48099 , n48098 );
and ( n48100 , n48099 , n39192 );
nor ( n48101 , n48095 , n48100 );
xnor ( n48102 , n48101 , n39199 );
and ( n48103 , n48094 , n48102 );
and ( n48104 , n48077 , n39186 );
and ( n48105 , n48102 , n48104 );
and ( n48106 , n48094 , n48104 );
or ( n48107 , n48103 , n48105 , n48106 );
and ( n48108 , n48099 , n39194 );
and ( n48109 , n47927 , n39192 );
nor ( n48110 , n48108 , n48109 );
xnor ( n48111 , n48110 , n39199 );
and ( n48112 , n48107 , n48111 );
and ( n48113 , n48086 , n39186 );
and ( n48114 , n48111 , n48113 );
and ( n48115 , n48107 , n48113 );
or ( n48116 , n48112 , n48114 , n48115 );
and ( n48117 , n47927 , n39194 );
and ( n48118 , n47932 , n39192 );
nor ( n48119 , n48117 , n48118 );
xnor ( n48120 , n48119 , n39199 );
and ( n48121 , n48116 , n48120 );
and ( n48122 , n48099 , n39186 );
and ( n48123 , n48120 , n48122 );
and ( n48124 , n48116 , n48122 );
or ( n48125 , n48121 , n48123 , n48124 );
and ( n48126 , n47932 , n39194 );
and ( n48127 , n47645 , n39192 );
nor ( n48128 , n48126 , n48127 );
xnor ( n48129 , n48128 , n39199 );
and ( n48130 , n48125 , n48129 );
and ( n48131 , n47927 , n39186 );
and ( n48132 , n48129 , n48131 );
and ( n48133 , n48125 , n48131 );
or ( n48134 , n48130 , n48132 , n48133 );
and ( n48135 , n47645 , n39194 );
and ( n48136 , n46948 , n39192 );
nor ( n48137 , n48135 , n48136 );
xnor ( n48138 , n48137 , n39199 );
and ( n48139 , n48134 , n48138 );
and ( n48140 , n47932 , n39186 );
and ( n48141 , n48138 , n48140 );
and ( n48142 , n48134 , n48140 );
or ( n48143 , n48139 , n48141 , n48142 );
and ( n48144 , n46948 , n39194 );
and ( n48145 , n46777 , n39192 );
nor ( n48146 , n48144 , n48145 );
xnor ( n48147 , n48146 , n39199 );
and ( n48148 , n48143 , n48147 );
and ( n48149 , n47645 , n39186 );
and ( n48150 , n48147 , n48149 );
and ( n48151 , n48143 , n48149 );
or ( n48152 , n48148 , n48150 , n48151 );
and ( n48153 , n48064 , n48152 );
and ( n48154 , n47777 , n48152 );
or ( n48155 , n48065 , n48153 , n48154 );
and ( n48156 , n47774 , n48155 );
and ( n48157 , n47772 , n48155 );
or ( n48158 , n47775 , n48156 , n48157 );
and ( n48159 , n47632 , n48158 );
and ( n48160 , n46676 , n39258 );
and ( n48161 , n46510 , n39256 );
nor ( n48162 , n48160 , n48161 );
xnor ( n48163 , n48162 , n39215 );
xor ( n48164 , n48143 , n48147 );
xor ( n48165 , n48164 , n48149 );
and ( n48166 , n48163 , n48165 );
xor ( n48167 , n47779 , n47781 );
xor ( n48168 , n48167 , n47841 );
xor ( n48169 , n47901 , n47903 );
xor ( n48170 , n48169 , n47906 );
xor ( n48171 , n47863 , n47879 );
xor ( n48172 , n48171 , n47882 );
xor ( n48173 , n47887 , n47889 );
xor ( n48174 , n48173 , n47892 );
and ( n48175 , n48172 , n48174 );
and ( n48176 , n47932 , n39335 );
and ( n48177 , n47645 , n39333 );
nor ( n48178 , n48176 , n48177 );
xnor ( n48179 , n48178 , n39300 );
and ( n48180 , n48099 , n39258 );
and ( n48181 , n47927 , n39256 );
nor ( n48182 , n48180 , n48181 );
xnor ( n48183 , n48182 , n39215 );
and ( n48184 , n48179 , n48183 );
xor ( n48185 , n47947 , n47949 );
and ( n48186 , n48183 , n48185 );
and ( n48187 , n48179 , n48185 );
or ( n48188 , n48184 , n48186 , n48187 );
and ( n48189 , n43820 , n40666 );
and ( n48190 , n43679 , n40664 );
nor ( n48191 , n48189 , n48190 );
xnor ( n48192 , n48191 , n40445 );
and ( n48193 , n44318 , n40406 );
and ( n48194 , n44000 , n40404 );
nor ( n48195 , n48193 , n48194 );
xnor ( n48196 , n48195 , n40262 );
and ( n48197 , n48192 , n48196 );
and ( n48198 , n42525 , n42079 );
and ( n48199 , n41828 , n42076 );
nor ( n48200 , n48198 , n48199 );
xnor ( n48201 , n48200 , n41370 );
and ( n48202 , n43040 , n41981 );
and ( n48203 , n42862 , n41979 );
nor ( n48204 , n48202 , n48203 );
xnor ( n48205 , n48204 , n41373 );
and ( n48206 , n48201 , n48205 );
and ( n48207 , n43322 , n41522 );
and ( n48208 , n43142 , n41520 );
nor ( n48209 , n48207 , n48208 );
xnor ( n48210 , n48209 , n41100 );
and ( n48211 , n48205 , n48210 );
and ( n48212 , n48201 , n48210 );
or ( n48213 , n48206 , n48211 , n48212 );
and ( n48214 , n48197 , n48213 );
and ( n48215 , n43524 , n41230 );
and ( n48216 , n43387 , n41228 );
nor ( n48217 , n48215 , n48216 );
xnor ( n48218 , n48217 , n40981 );
and ( n48219 , n43671 , n40928 );
and ( n48220 , n43549 , n40926 );
nor ( n48221 , n48219 , n48220 );
xnor ( n48222 , n48221 , n40688 );
and ( n48223 , n48218 , n48222 );
and ( n48224 , n44826 , n40168 );
and ( n48225 , n44347 , n40166 );
nor ( n48226 , n48224 , n48225 );
xnor ( n48227 , n48226 , n40059 );
and ( n48228 , n48222 , n48227 );
and ( n48229 , n48218 , n48227 );
or ( n48230 , n48223 , n48228 , n48229 );
and ( n48231 , n48213 , n48230 );
and ( n48232 , n48197 , n48230 );
or ( n48233 , n48214 , n48231 , n48232 );
and ( n48234 , n48188 , n48233 );
and ( n48235 , n45171 , n39984 );
and ( n48236 , n45057 , n39982 );
nor ( n48237 , n48235 , n48236 );
xnor ( n48238 , n48237 , n39865 );
and ( n48239 , n46069 , n39795 );
and ( n48240 , n45754 , n39793 );
nor ( n48241 , n48239 , n48240 );
xnor ( n48242 , n48241 , n39729 );
and ( n48243 , n48238 , n48242 );
and ( n48244 , n46510 , n39665 );
and ( n48245 , n46159 , n39663 );
nor ( n48246 , n48244 , n48245 );
xnor ( n48247 , n48246 , n39608 );
and ( n48248 , n48242 , n48247 );
and ( n48249 , n48238 , n48247 );
or ( n48250 , n48243 , n48248 , n48249 );
and ( n48251 , n46777 , n39532 );
and ( n48252 , n46676 , n39530 );
nor ( n48253 , n48251 , n48252 );
xnor ( n48254 , n48253 , n39497 );
and ( n48255 , n47645 , n39384 );
and ( n48256 , n46948 , n39382 );
nor ( n48257 , n48255 , n48256 );
xnor ( n48258 , n48257 , n39367 );
and ( n48259 , n48254 , n48258 );
and ( n48260 , n47927 , n39335 );
and ( n48261 , n47932 , n39333 );
nor ( n48262 , n48260 , n48261 );
xnor ( n48263 , n48262 , n39300 );
and ( n48264 , n48258 , n48263 );
and ( n48265 , n48254 , n48263 );
or ( n48266 , n48259 , n48264 , n48265 );
and ( n48267 , n48250 , n48266 );
xor ( n48268 , n47955 , n47959 );
xor ( n48269 , n48268 , n47964 );
and ( n48270 , n48266 , n48269 );
and ( n48271 , n48250 , n48269 );
or ( n48272 , n48267 , n48270 , n48271 );
and ( n48273 , n48233 , n48272 );
and ( n48274 , n48188 , n48272 );
or ( n48275 , n48234 , n48273 , n48274 );
and ( n48276 , n48174 , n48275 );
and ( n48277 , n48172 , n48275 );
or ( n48278 , n48175 , n48276 , n48277 );
xor ( n48279 , n47980 , n47984 );
xor ( n48280 , n48279 , n47989 );
xor ( n48281 , n47996 , n48000 );
xor ( n48282 , n48281 , n48005 );
and ( n48283 , n48280 , n48282 );
xor ( n48284 , n48013 , n48017 );
xor ( n48285 , n48284 , n48022 );
and ( n48286 , n48282 , n48285 );
and ( n48287 , n48280 , n48285 );
or ( n48288 , n48283 , n48286 , n48287 );
xor ( n48289 , n47923 , n47935 );
xor ( n48290 , n48289 , n47938 );
and ( n48291 , n48288 , n48290 );
xor ( n48292 , n47943 , n47950 );
xor ( n48293 , n48292 , n47967 );
and ( n48294 , n48290 , n48293 );
and ( n48295 , n48288 , n48293 );
or ( n48296 , n48291 , n48294 , n48295 );
xor ( n48297 , n47919 , n47941 );
xor ( n48298 , n48297 , n47970 );
and ( n48299 , n48296 , n48298 );
xor ( n48300 , n48028 , n48038 );
xor ( n48301 , n48300 , n48041 );
and ( n48302 , n48298 , n48301 );
and ( n48303 , n48296 , n48301 );
or ( n48304 , n48299 , n48302 , n48303 );
and ( n48305 , n48278 , n48304 );
xor ( n48306 , n47914 , n47916 );
xor ( n48307 , n48306 , n47973 );
and ( n48308 , n48304 , n48307 );
and ( n48309 , n48278 , n48307 );
or ( n48310 , n48305 , n48308 , n48309 );
and ( n48311 , n48170 , n48310 );
xor ( n48312 , n47976 , n48052 );
xor ( n48313 , n48312 , n48055 );
and ( n48314 , n48310 , n48313 );
and ( n48315 , n48170 , n48313 );
or ( n48316 , n48311 , n48314 , n48315 );
and ( n48317 , n48168 , n48316 );
xor ( n48318 , n47909 , n47911 );
xor ( n48319 , n48318 , n48058 );
and ( n48320 , n48316 , n48319 );
and ( n48321 , n48168 , n48319 );
or ( n48322 , n48317 , n48320 , n48321 );
xor ( n48323 , n47844 , n47846 );
xor ( n48324 , n48323 , n48061 );
and ( n48325 , n48322 , n48324 );
and ( n48326 , n46777 , n39258 );
and ( n48327 , n46676 , n39256 );
nor ( n48328 , n48326 , n48327 );
xnor ( n48329 , n48328 , n39215 );
xor ( n48330 , n48134 , n48138 );
xor ( n48331 , n48330 , n48140 );
and ( n48332 , n48329 , n48331 );
and ( n48333 , n48324 , n48332 );
and ( n48334 , n48322 , n48332 );
or ( n48335 , n48325 , n48333 , n48334 );
and ( n48336 , n48166 , n48335 );
xor ( n48337 , n47777 , n48064 );
xor ( n48338 , n48337 , n48152 );
and ( n48339 , n48335 , n48338 );
and ( n48340 , n48166 , n48338 );
or ( n48341 , n48336 , n48339 , n48340 );
xor ( n48342 , n47772 , n47774 );
xor ( n48343 , n48342 , n48155 );
and ( n48344 , n48341 , n48343 );
xor ( n48345 , n48163 , n48165 );
xor ( n48346 , n48125 , n48129 );
xor ( n48347 , n48346 , n48131 );
xor ( n48348 , n48044 , n48046 );
xor ( n48349 , n48348 , n48049 );
xor ( n48350 , n48116 , n48120 );
xor ( n48351 , n48350 , n48122 );
and ( n48352 , n48349 , n48351 );
and ( n48353 , n47932 , n39258 );
and ( n48354 , n47645 , n39256 );
nor ( n48355 , n48353 , n48354 );
xnor ( n48356 , n48355 , n39215 );
xor ( n48357 , n48107 , n48111 );
xor ( n48358 , n48357 , n48113 );
or ( n48359 , n48356 , n48358 );
and ( n48360 , n48351 , n48359 );
and ( n48361 , n48349 , n48359 );
or ( n48362 , n48352 , n48360 , n48361 );
and ( n48363 , n48347 , n48362 );
xor ( n48364 , n48170 , n48310 );
xor ( n48365 , n48364 , n48313 );
and ( n48366 , n48362 , n48365 );
and ( n48367 , n48347 , n48365 );
or ( n48368 , n48363 , n48366 , n48367 );
xor ( n48369 , n48168 , n48316 );
xor ( n48370 , n48369 , n48319 );
and ( n48371 , n48368 , n48370 );
xor ( n48372 , n48329 , n48331 );
and ( n48373 , n48370 , n48372 );
and ( n48374 , n48368 , n48372 );
or ( n48375 , n48371 , n48373 , n48374 );
and ( n48376 , n48345 , n48375 );
xor ( n48377 , n48322 , n48324 );
xor ( n48378 , n48377 , n48332 );
and ( n48379 , n48375 , n48378 );
and ( n48380 , n48345 , n48378 );
or ( n48381 , n48376 , n48379 , n48380 );
xor ( n48382 , n48166 , n48335 );
xor ( n48383 , n48382 , n48338 );
or ( n48384 , n48381 , n48383 );
and ( n48385 , n48343 , n48384 );
and ( n48386 , n48341 , n48384 );
or ( n48387 , n48344 , n48385 , n48386 );
and ( n48388 , n48158 , n48387 );
and ( n48389 , n47632 , n48387 );
or ( n48390 , n48159 , n48388 , n48389 );
and ( n48391 , n47630 , n48390 );
xor ( n48392 , n47630 , n48390 );
xor ( n48393 , n47632 , n48158 );
xor ( n48394 , n48393 , n48387 );
xor ( n48395 , n48341 , n48343 );
xor ( n48396 , n48395 , n48384 );
not ( n48397 , n48396 );
xnor ( n48398 , n48381 , n48383 );
xor ( n48399 , n48345 , n48375 );
xor ( n48400 , n48399 , n48378 );
xor ( n48401 , n47992 , n48008 );
xor ( n48402 , n48401 , n48025 );
xor ( n48403 , n48030 , n48032 );
xor ( n48404 , n48403 , n48035 );
and ( n48405 , n48402 , n48404 );
xor ( n48406 , n48094 , n48102 );
xor ( n48407 , n48406 , n48104 );
and ( n48408 , n48404 , n48407 );
and ( n48409 , n48402 , n48407 );
or ( n48410 , n48405 , n48408 , n48409 );
xor ( n48411 , n48081 , n48089 );
xor ( n48412 , n48411 , n48091 );
and ( n48413 , n48086 , n39258 );
and ( n48414 , n48099 , n39256 );
nor ( n48415 , n48413 , n48414 );
xnor ( n48416 , n48415 , n39215 );
xor ( n48417 , n48072 , n48080 );
and ( n48418 , n48416 , n48417 );
and ( n48419 , n48412 , n48418 );
buf ( n48420 , n30378 );
not ( n48421 , n48420 );
xor ( n48422 , n48192 , n48196 );
and ( n48423 , n48421 , n48422 );
and ( n48424 , n42862 , n42079 );
and ( n48425 , n42525 , n42076 );
nor ( n48426 , n48424 , n48425 );
xnor ( n48427 , n48426 , n41370 );
and ( n48428 , n43142 , n41981 );
and ( n48429 , n43040 , n41979 );
nor ( n48430 , n48428 , n48429 );
xnor ( n48431 , n48430 , n41373 );
and ( n48432 , n48427 , n48431 );
and ( n48433 , n43387 , n41522 );
and ( n48434 , n43322 , n41520 );
nor ( n48435 , n48433 , n48434 );
xnor ( n48436 , n48435 , n41100 );
and ( n48437 , n48431 , n48436 );
and ( n48438 , n48427 , n48436 );
or ( n48439 , n48432 , n48437 , n48438 );
and ( n48440 , n48422 , n48439 );
and ( n48441 , n48421 , n48439 );
or ( n48442 , n48423 , n48440 , n48441 );
and ( n48443 , n48418 , n48442 );
and ( n48444 , n48412 , n48442 );
or ( n48445 , n48419 , n48443 , n48444 );
and ( n48446 , n43549 , n41230 );
and ( n48447 , n43524 , n41228 );
nor ( n48448 , n48446 , n48447 );
xnor ( n48449 , n48448 , n40981 );
and ( n48450 , n43679 , n40928 );
and ( n48451 , n43671 , n40926 );
nor ( n48452 , n48450 , n48451 );
xnor ( n48453 , n48452 , n40688 );
and ( n48454 , n48449 , n48453 );
and ( n48455 , n44000 , n40666 );
and ( n48456 , n43820 , n40664 );
nor ( n48457 , n48455 , n48456 );
xnor ( n48458 , n48457 , n40445 );
and ( n48459 , n48453 , n48458 );
and ( n48460 , n48449 , n48458 );
or ( n48461 , n48454 , n48459 , n48460 );
and ( n48462 , n44347 , n40406 );
and ( n48463 , n44318 , n40404 );
nor ( n48464 , n48462 , n48463 );
xnor ( n48465 , n48464 , n40262 );
and ( n48466 , n45057 , n40168 );
and ( n48467 , n44826 , n40166 );
nor ( n48468 , n48466 , n48467 );
xnor ( n48469 , n48468 , n40059 );
and ( n48470 , n48465 , n48469 );
and ( n48471 , n45754 , n39984 );
and ( n48472 , n45171 , n39982 );
nor ( n48473 , n48471 , n48472 );
xnor ( n48474 , n48473 , n39865 );
and ( n48475 , n48469 , n48474 );
and ( n48476 , n48465 , n48474 );
or ( n48477 , n48470 , n48475 , n48476 );
and ( n48478 , n48461 , n48477 );
and ( n48479 , n46159 , n39795 );
and ( n48480 , n46069 , n39793 );
nor ( n48481 , n48479 , n48480 );
xnor ( n48482 , n48481 , n39729 );
and ( n48483 , n46676 , n39665 );
and ( n48484 , n46510 , n39663 );
nor ( n48485 , n48483 , n48484 );
xnor ( n48486 , n48485 , n39608 );
and ( n48487 , n48482 , n48486 );
and ( n48488 , n46948 , n39532 );
and ( n48489 , n46777 , n39530 );
nor ( n48490 , n48488 , n48489 );
xnor ( n48491 , n48490 , n39497 );
and ( n48492 , n48486 , n48491 );
and ( n48493 , n48482 , n48491 );
or ( n48494 , n48487 , n48492 , n48493 );
and ( n48495 , n48477 , n48494 );
and ( n48496 , n48461 , n48494 );
or ( n48497 , n48478 , n48495 , n48496 );
xor ( n48498 , n48201 , n48205 );
xor ( n48499 , n48498 , n48210 );
xor ( n48500 , n48218 , n48222 );
xor ( n48501 , n48500 , n48227 );
and ( n48502 , n48499 , n48501 );
xor ( n48503 , n48238 , n48242 );
xor ( n48504 , n48503 , n48247 );
and ( n48505 , n48501 , n48504 );
and ( n48506 , n48499 , n48504 );
or ( n48507 , n48502 , n48505 , n48506 );
and ( n48508 , n48497 , n48507 );
xor ( n48509 , n48179 , n48183 );
xor ( n48510 , n48509 , n48185 );
and ( n48511 , n48507 , n48510 );
and ( n48512 , n48497 , n48510 );
or ( n48513 , n48508 , n48511 , n48512 );
and ( n48514 , n48445 , n48513 );
xor ( n48515 , n48197 , n48213 );
xor ( n48516 , n48515 , n48230 );
xor ( n48517 , n48250 , n48266 );
xor ( n48518 , n48517 , n48269 );
and ( n48519 , n48516 , n48518 );
xor ( n48520 , n48280 , n48282 );
xor ( n48521 , n48520 , n48285 );
and ( n48522 , n48518 , n48521 );
and ( n48523 , n48516 , n48521 );
or ( n48524 , n48519 , n48522 , n48523 );
and ( n48525 , n48513 , n48524 );
and ( n48526 , n48445 , n48524 );
or ( n48527 , n48514 , n48525 , n48526 );
and ( n48528 , n48410 , n48527 );
xor ( n48529 , n48172 , n48174 );
xor ( n48530 , n48529 , n48275 );
and ( n48531 , n48527 , n48530 );
and ( n48532 , n48410 , n48530 );
or ( n48533 , n48528 , n48531 , n48532 );
xor ( n48534 , n48278 , n48304 );
xor ( n48535 , n48534 , n48307 );
and ( n48536 , n48533 , n48535 );
xor ( n48537 , n48296 , n48298 );
xor ( n48538 , n48537 , n48301 );
xnor ( n48539 , n48356 , n48358 );
and ( n48540 , n48538 , n48539 );
xor ( n48541 , n48188 , n48233 );
xor ( n48542 , n48541 , n48272 );
xor ( n48543 , n48288 , n48290 );
xor ( n48544 , n48543 , n48293 );
and ( n48545 , n48542 , n48544 );
xor ( n48546 , n48254 , n48258 );
xor ( n48547 , n48546 , n48263 );
xor ( n48548 , n48416 , n48417 );
and ( n48549 , n48547 , n48548 );
and ( n48550 , n48069 , n39256 );
not ( n48551 , n48550 );
and ( n48552 , n48551 , n39215 );
and ( n48553 , n48069 , n39258 );
and ( n48554 , n48077 , n39256 );
nor ( n48555 , n48553 , n48554 );
xnor ( n48556 , n48555 , n39215 );
and ( n48557 , n48552 , n48556 );
or ( n48558 , n48557 , n48070 );
and ( n48559 , n48548 , n48558 );
and ( n48560 , n48547 , n48558 );
or ( n48561 , n48549 , n48559 , n48560 );
and ( n48562 , n47932 , n39384 );
and ( n48563 , n47645 , n39382 );
nor ( n48564 , n48562 , n48563 );
xnor ( n48565 , n48564 , n39367 );
buf ( n48566 , n30379 );
not ( n48567 , n48566 );
and ( n48568 , n48565 , n48567 );
and ( n48569 , n45171 , n40168 );
and ( n48570 , n45057 , n40166 );
nor ( n48571 , n48569 , n48570 );
xnor ( n48572 , n48571 , n40059 );
buf ( n48573 , n30380 );
not ( n48574 , n48573 );
and ( n48575 , n48572 , n48574 );
and ( n48576 , n48567 , n48575 );
and ( n48577 , n48565 , n48575 );
or ( n48578 , n48568 , n48576 , n48577 );
and ( n48579 , n43040 , n42079 );
and ( n48580 , n42862 , n42076 );
nor ( n48581 , n48579 , n48580 );
xnor ( n48582 , n48581 , n41370 );
and ( n48583 , n43322 , n41981 );
and ( n48584 , n43142 , n41979 );
nor ( n48585 , n48583 , n48584 );
xnor ( n48586 , n48585 , n41373 );
and ( n48587 , n48582 , n48586 );
and ( n48588 , n43524 , n41522 );
and ( n48589 , n43387 , n41520 );
nor ( n48590 , n48588 , n48589 );
xnor ( n48591 , n48590 , n41100 );
and ( n48592 , n48586 , n48591 );
and ( n48593 , n48582 , n48591 );
or ( n48594 , n48587 , n48592 , n48593 );
and ( n48595 , n43671 , n41230 );
and ( n48596 , n43549 , n41228 );
nor ( n48597 , n48595 , n48596 );
xnor ( n48598 , n48597 , n40981 );
and ( n48599 , n43820 , n40928 );
and ( n48600 , n43679 , n40926 );
nor ( n48601 , n48599 , n48600 );
xnor ( n48602 , n48601 , n40688 );
and ( n48603 , n48598 , n48602 );
and ( n48604 , n44318 , n40666 );
and ( n48605 , n44000 , n40664 );
nor ( n48606 , n48604 , n48605 );
xnor ( n48607 , n48606 , n40445 );
and ( n48608 , n48602 , n48607 );
and ( n48609 , n48598 , n48607 );
or ( n48610 , n48603 , n48608 , n48609 );
and ( n48611 , n48594 , n48610 );
and ( n48612 , n44826 , n40406 );
and ( n48613 , n44347 , n40404 );
nor ( n48614 , n48612 , n48613 );
xnor ( n48615 , n48614 , n40262 );
and ( n48616 , n46069 , n39984 );
and ( n48617 , n45754 , n39982 );
nor ( n48618 , n48616 , n48617 );
xnor ( n48619 , n48618 , n39865 );
and ( n48620 , n48615 , n48619 );
and ( n48621 , n46510 , n39795 );
and ( n48622 , n46159 , n39793 );
nor ( n48623 , n48621 , n48622 );
xnor ( n48624 , n48623 , n39729 );
and ( n48625 , n48619 , n48624 );
and ( n48626 , n48615 , n48624 );
or ( n48627 , n48620 , n48625 , n48626 );
and ( n48628 , n48610 , n48627 );
and ( n48629 , n48594 , n48627 );
or ( n48630 , n48611 , n48628 , n48629 );
and ( n48631 , n48578 , n48630 );
and ( n48632 , n46777 , n39665 );
and ( n48633 , n46676 , n39663 );
nor ( n48634 , n48632 , n48633 );
xnor ( n48635 , n48634 , n39608 );
and ( n48636 , n47645 , n39532 );
and ( n48637 , n46948 , n39530 );
nor ( n48638 , n48636 , n48637 );
xnor ( n48639 , n48638 , n39497 );
and ( n48640 , n48635 , n48639 );
and ( n48641 , n47927 , n39384 );
and ( n48642 , n47932 , n39382 );
nor ( n48643 , n48641 , n48642 );
xnor ( n48644 , n48643 , n39367 );
and ( n48645 , n48639 , n48644 );
and ( n48646 , n48635 , n48644 );
or ( n48647 , n48640 , n48645 , n48646 );
xor ( n48648 , n48427 , n48431 );
xor ( n48649 , n48648 , n48436 );
and ( n48650 , n48647 , n48649 );
xor ( n48651 , n48449 , n48453 );
xor ( n48652 , n48651 , n48458 );
and ( n48653 , n48649 , n48652 );
and ( n48654 , n48647 , n48652 );
or ( n48655 , n48650 , n48653 , n48654 );
and ( n48656 , n48630 , n48655 );
and ( n48657 , n48578 , n48655 );
or ( n48658 , n48631 , n48656 , n48657 );
and ( n48659 , n48561 , n48658 );
xor ( n48660 , n48421 , n48422 );
xor ( n48661 , n48660 , n48439 );
xor ( n48662 , n48461 , n48477 );
xor ( n48663 , n48662 , n48494 );
and ( n48664 , n48661 , n48663 );
xor ( n48665 , n48499 , n48501 );
xor ( n48666 , n48665 , n48504 );
and ( n48667 , n48663 , n48666 );
and ( n48668 , n48661 , n48666 );
or ( n48669 , n48664 , n48667 , n48668 );
and ( n48670 , n48658 , n48669 );
and ( n48671 , n48561 , n48669 );
or ( n48672 , n48659 , n48670 , n48671 );
and ( n48673 , n48544 , n48672 );
and ( n48674 , n48542 , n48672 );
or ( n48675 , n48545 , n48673 , n48674 );
and ( n48676 , n48539 , n48675 );
and ( n48677 , n48538 , n48675 );
or ( n48678 , n48540 , n48676 , n48677 );
and ( n48679 , n48535 , n48678 );
and ( n48680 , n48533 , n48678 );
or ( n48681 , n48536 , n48679 , n48680 );
xor ( n48682 , n48347 , n48362 );
xor ( n48683 , n48682 , n48365 );
and ( n48684 , n48681 , n48683 );
xor ( n48685 , n48349 , n48351 );
xor ( n48686 , n48685 , n48359 );
xor ( n48687 , n48412 , n48418 );
xor ( n48688 , n48687 , n48442 );
xor ( n48689 , n48497 , n48507 );
xor ( n48690 , n48689 , n48510 );
and ( n48691 , n48688 , n48690 );
xor ( n48692 , n48516 , n48518 );
xor ( n48693 , n48692 , n48521 );
and ( n48694 , n48690 , n48693 );
and ( n48695 , n48688 , n48693 );
or ( n48696 , n48691 , n48694 , n48695 );
xor ( n48697 , n48402 , n48404 );
xor ( n48698 , n48697 , n48407 );
and ( n48699 , n48696 , n48698 );
xor ( n48700 , n48445 , n48513 );
xor ( n48701 , n48700 , n48524 );
and ( n48702 , n48698 , n48701 );
and ( n48703 , n48696 , n48701 );
or ( n48704 , n48699 , n48702 , n48703 );
xor ( n48705 , n48410 , n48527 );
xor ( n48706 , n48705 , n48530 );
and ( n48707 , n48704 , n48706 );
and ( n48708 , n48077 , n39258 );
and ( n48709 , n48086 , n39256 );
nor ( n48710 , n48708 , n48709 );
xnor ( n48711 , n48710 , n39215 );
xnor ( n48712 , n48557 , n48070 );
or ( n48713 , n48711 , n48712 );
xor ( n48714 , n48465 , n48469 );
xor ( n48715 , n48714 , n48474 );
xor ( n48716 , n48482 , n48486 );
xor ( n48717 , n48716 , n48491 );
and ( n48718 , n48715 , n48717 );
and ( n48719 , n48086 , n39335 );
and ( n48720 , n48099 , n39333 );
nor ( n48721 , n48719 , n48720 );
xnor ( n48722 , n48721 , n39300 );
xor ( n48723 , n48552 , n48556 );
or ( n48724 , n48722 , n48723 );
and ( n48725 , n48717 , n48724 );
and ( n48726 , n48715 , n48724 );
or ( n48727 , n48718 , n48725 , n48726 );
and ( n48728 , n48713 , n48727 );
xor ( n48729 , n48572 , n48574 );
and ( n48730 , n43387 , n41981 );
and ( n48731 , n43322 , n41979 );
nor ( n48732 , n48730 , n48731 );
xnor ( n48733 , n48732 , n41373 );
and ( n48734 , n43549 , n41522 );
and ( n48735 , n43524 , n41520 );
nor ( n48736 , n48734 , n48735 );
xnor ( n48737 , n48736 , n41100 );
or ( n48738 , n48733 , n48737 );
and ( n48739 , n48729 , n48738 );
and ( n48740 , n43142 , n42079 );
and ( n48741 , n43040 , n42076 );
nor ( n48742 , n48740 , n48741 );
xnor ( n48743 , n48742 , n41370 );
and ( n48744 , n43679 , n41230 );
and ( n48745 , n43671 , n41228 );
nor ( n48746 , n48744 , n48745 );
xnor ( n48747 , n48746 , n40981 );
and ( n48748 , n48743 , n48747 );
and ( n48749 , n44000 , n40928 );
and ( n48750 , n43820 , n40926 );
nor ( n48751 , n48749 , n48750 );
xnor ( n48752 , n48751 , n40688 );
and ( n48753 , n48747 , n48752 );
and ( n48754 , n48743 , n48752 );
or ( n48755 , n48748 , n48753 , n48754 );
and ( n48756 , n48738 , n48755 );
and ( n48757 , n48729 , n48755 );
or ( n48758 , n48739 , n48756 , n48757 );
and ( n48759 , n44347 , n40666 );
and ( n48760 , n44318 , n40664 );
nor ( n48761 , n48759 , n48760 );
xnor ( n48762 , n48761 , n40445 );
and ( n48763 , n45057 , n40406 );
and ( n48764 , n44826 , n40404 );
nor ( n48765 , n48763 , n48764 );
xnor ( n48766 , n48765 , n40262 );
and ( n48767 , n48762 , n48766 );
and ( n48768 , n45754 , n40168 );
and ( n48769 , n45171 , n40166 );
nor ( n48770 , n48768 , n48769 );
xnor ( n48771 , n48770 , n40059 );
and ( n48772 , n48766 , n48771 );
and ( n48773 , n48762 , n48771 );
or ( n48774 , n48767 , n48772 , n48773 );
and ( n48775 , n46159 , n39984 );
and ( n48776 , n46069 , n39982 );
nor ( n48777 , n48775 , n48776 );
xnor ( n48778 , n48777 , n39865 );
and ( n48779 , n46676 , n39795 );
and ( n48780 , n46510 , n39793 );
nor ( n48781 , n48779 , n48780 );
xnor ( n48782 , n48781 , n39729 );
and ( n48783 , n48778 , n48782 );
and ( n48784 , n46948 , n39665 );
and ( n48785 , n46777 , n39663 );
nor ( n48786 , n48784 , n48785 );
xnor ( n48787 , n48786 , n39608 );
and ( n48788 , n48782 , n48787 );
and ( n48789 , n48778 , n48787 );
or ( n48790 , n48783 , n48788 , n48789 );
and ( n48791 , n48774 , n48790 );
and ( n48792 , n47932 , n39532 );
and ( n48793 , n47645 , n39530 );
nor ( n48794 , n48792 , n48793 );
xnor ( n48795 , n48794 , n39497 );
and ( n48796 , n48099 , n39384 );
and ( n48797 , n47927 , n39382 );
nor ( n48798 , n48796 , n48797 );
xnor ( n48799 , n48798 , n39367 );
and ( n48800 , n48795 , n48799 );
and ( n48801 , n48077 , n39335 );
and ( n48802 , n48086 , n39333 );
nor ( n48803 , n48801 , n48802 );
xnor ( n48804 , n48803 , n39300 );
and ( n48805 , n48799 , n48804 );
and ( n48806 , n48795 , n48804 );
or ( n48807 , n48800 , n48805 , n48806 );
and ( n48808 , n48790 , n48807 );
and ( n48809 , n48774 , n48807 );
or ( n48810 , n48791 , n48808 , n48809 );
and ( n48811 , n48758 , n48810 );
xor ( n48812 , n48582 , n48586 );
xor ( n48813 , n48812 , n48591 );
xor ( n48814 , n48598 , n48602 );
xor ( n48815 , n48814 , n48607 );
and ( n48816 , n48813 , n48815 );
xor ( n48817 , n48615 , n48619 );
xor ( n48818 , n48817 , n48624 );
and ( n48819 , n48815 , n48818 );
and ( n48820 , n48813 , n48818 );
or ( n48821 , n48816 , n48819 , n48820 );
and ( n48822 , n48810 , n48821 );
and ( n48823 , n48758 , n48821 );
or ( n48824 , n48811 , n48822 , n48823 );
and ( n48825 , n48727 , n48824 );
and ( n48826 , n48713 , n48824 );
or ( n48827 , n48728 , n48825 , n48826 );
xor ( n48828 , n48565 , n48567 );
xor ( n48829 , n48828 , n48575 );
xor ( n48830 , n48594 , n48610 );
xor ( n48831 , n48830 , n48627 );
and ( n48832 , n48829 , n48831 );
xor ( n48833 , n48647 , n48649 );
xor ( n48834 , n48833 , n48652 );
and ( n48835 , n48831 , n48834 );
and ( n48836 , n48829 , n48834 );
or ( n48837 , n48832 , n48835 , n48836 );
xor ( n48838 , n48547 , n48548 );
xor ( n48839 , n48838 , n48558 );
and ( n48840 , n48837 , n48839 );
xor ( n48841 , n48578 , n48630 );
xor ( n48842 , n48841 , n48655 );
and ( n48843 , n48839 , n48842 );
and ( n48844 , n48837 , n48842 );
or ( n48845 , n48840 , n48843 , n48844 );
and ( n48846 , n48827 , n48845 );
xor ( n48847 , n48561 , n48658 );
xor ( n48848 , n48847 , n48669 );
and ( n48849 , n48845 , n48848 );
and ( n48850 , n48827 , n48848 );
or ( n48851 , n48846 , n48849 , n48850 );
xor ( n48852 , n48542 , n48544 );
xor ( n48853 , n48852 , n48672 );
and ( n48854 , n48851 , n48853 );
xor ( n48855 , n48696 , n48698 );
xor ( n48856 , n48855 , n48701 );
and ( n48857 , n48853 , n48856 );
and ( n48858 , n48851 , n48856 );
or ( n48859 , n48854 , n48857 , n48858 );
and ( n48860 , n48706 , n48859 );
and ( n48861 , n48704 , n48859 );
or ( n48862 , n48707 , n48860 , n48861 );
and ( n48863 , n48686 , n48862 );
xor ( n48864 , n48533 , n48535 );
xor ( n48865 , n48864 , n48678 );
and ( n48866 , n48862 , n48865 );
and ( n48867 , n48686 , n48865 );
or ( n48868 , n48863 , n48866 , n48867 );
and ( n48869 , n48683 , n48868 );
and ( n48870 , n48681 , n48868 );
or ( n48871 , n48684 , n48869 , n48870 );
xor ( n48872 , n48368 , n48370 );
xor ( n48873 , n48872 , n48372 );
and ( n48874 , n48871 , n48873 );
xor ( n48875 , n48681 , n48683 );
xor ( n48876 , n48875 , n48868 );
xor ( n48877 , n48686 , n48862 );
xor ( n48878 , n48877 , n48865 );
xor ( n48879 , n48538 , n48539 );
xor ( n48880 , n48879 , n48675 );
xor ( n48881 , n48704 , n48706 );
xor ( n48882 , n48881 , n48859 );
and ( n48883 , n48880 , n48882 );
xor ( n48884 , n48688 , n48690 );
xor ( n48885 , n48884 , n48693 );
xor ( n48886 , n48661 , n48663 );
xor ( n48887 , n48886 , n48666 );
and ( n48888 , n48099 , n39335 );
and ( n48889 , n47927 , n39333 );
nor ( n48890 , n48888 , n48889 );
xnor ( n48891 , n48890 , n39300 );
xnor ( n48892 , n48711 , n48712 );
or ( n48893 , n48891 , n48892 );
and ( n48894 , n48887 , n48893 );
xor ( n48895 , n48635 , n48639 );
xor ( n48896 , n48895 , n48644 );
xnor ( n48897 , n48722 , n48723 );
and ( n48898 , n48896 , n48897 );
buf ( n48899 , n30381 );
not ( n48900 , n48899 );
and ( n48901 , n48550 , n48900 );
xnor ( n48902 , n48733 , n48737 );
and ( n48903 , n48900 , n48902 );
and ( n48904 , n48550 , n48902 );
or ( n48905 , n48901 , n48903 , n48904 );
and ( n48906 , n48897 , n48905 );
and ( n48907 , n48896 , n48905 );
or ( n48908 , n48898 , n48906 , n48907 );
and ( n48909 , n48069 , n39333 );
not ( n48910 , n48909 );
and ( n48911 , n48910 , n39300 );
and ( n48912 , n48069 , n39335 );
and ( n48913 , n48077 , n39333 );
nor ( n48914 , n48912 , n48913 );
xnor ( n48915 , n48914 , n39300 );
and ( n48916 , n48911 , n48915 );
and ( n48917 , n43820 , n41230 );
and ( n48918 , n43679 , n41228 );
nor ( n48919 , n48917 , n48918 );
xnor ( n48920 , n48919 , n40981 );
and ( n48921 , n44318 , n40928 );
and ( n48922 , n44000 , n40926 );
nor ( n48923 , n48921 , n48922 );
xnor ( n48924 , n48923 , n40688 );
or ( n48925 , n48920 , n48924 );
and ( n48926 , n48916 , n48925 );
and ( n48927 , n43322 , n42079 );
and ( n48928 , n43142 , n42076 );
nor ( n48929 , n48927 , n48928 );
xnor ( n48930 , n48929 , n41370 );
and ( n48931 , n43524 , n41981 );
and ( n48932 , n43387 , n41979 );
nor ( n48933 , n48931 , n48932 );
xnor ( n48934 , n48933 , n41373 );
and ( n48935 , n48930 , n48934 );
and ( n48936 , n43671 , n41522 );
and ( n48937 , n43549 , n41520 );
nor ( n48938 , n48936 , n48937 );
xnor ( n48939 , n48938 , n41100 );
and ( n48940 , n48934 , n48939 );
and ( n48941 , n48930 , n48939 );
or ( n48942 , n48935 , n48940 , n48941 );
and ( n48943 , n48925 , n48942 );
and ( n48944 , n48916 , n48942 );
or ( n48945 , n48926 , n48943 , n48944 );
and ( n48946 , n44826 , n40666 );
and ( n48947 , n44347 , n40664 );
nor ( n48948 , n48946 , n48947 );
xnor ( n48949 , n48948 , n40445 );
and ( n48950 , n45171 , n40406 );
and ( n48951 , n45057 , n40404 );
nor ( n48952 , n48950 , n48951 );
xnor ( n48953 , n48952 , n40262 );
and ( n48954 , n48949 , n48953 );
and ( n48955 , n46069 , n40168 );
and ( n48956 , n45754 , n40166 );
nor ( n48957 , n48955 , n48956 );
xnor ( n48958 , n48957 , n40059 );
and ( n48959 , n48953 , n48958 );
and ( n48960 , n48949 , n48958 );
or ( n48961 , n48954 , n48959 , n48960 );
xor ( n48962 , n48743 , n48747 );
xor ( n48963 , n48962 , n48752 );
and ( n48964 , n48961 , n48963 );
xor ( n48965 , n48762 , n48766 );
xor ( n48966 , n48965 , n48771 );
and ( n48967 , n48963 , n48966 );
and ( n48968 , n48961 , n48966 );
or ( n48969 , n48964 , n48967 , n48968 );
and ( n48970 , n48945 , n48969 );
xor ( n48971 , n48729 , n48738 );
xor ( n48972 , n48971 , n48755 );
and ( n48973 , n48969 , n48972 );
and ( n48974 , n48945 , n48972 );
or ( n48975 , n48970 , n48973 , n48974 );
and ( n48976 , n48908 , n48975 );
xor ( n48977 , n48715 , n48717 );
xor ( n48978 , n48977 , n48724 );
and ( n48979 , n48975 , n48978 );
and ( n48980 , n48908 , n48978 );
or ( n48981 , n48976 , n48979 , n48980 );
and ( n48982 , n48893 , n48981 );
and ( n48983 , n48887 , n48981 );
or ( n48984 , n48894 , n48982 , n48983 );
and ( n48985 , n48885 , n48984 );
xor ( n48986 , n48827 , n48845 );
xor ( n48987 , n48986 , n48848 );
and ( n48988 , n48984 , n48987 );
and ( n48989 , n48885 , n48987 );
or ( n48990 , n48985 , n48988 , n48989 );
xor ( n48991 , n48851 , n48853 );
xor ( n48992 , n48991 , n48856 );
and ( n48993 , n48990 , n48992 );
xor ( n48994 , n48713 , n48727 );
xor ( n48995 , n48994 , n48824 );
xor ( n48996 , n48837 , n48839 );
xor ( n48997 , n48996 , n48842 );
and ( n48998 , n48995 , n48997 );
xor ( n48999 , n48758 , n48810 );
xor ( n49000 , n48999 , n48821 );
xor ( n49001 , n48829 , n48831 );
xor ( n49002 , n49001 , n48834 );
and ( n49003 , n49000 , n49002 );
xnor ( n49004 , n48891 , n48892 );
and ( n49005 , n49002 , n49004 );
and ( n49006 , n49000 , n49004 );
or ( n49007 , n49003 , n49005 , n49006 );
and ( n49008 , n48997 , n49007 );
and ( n49009 , n48995 , n49007 );
or ( n49010 , n48998 , n49008 , n49009 );
xor ( n49011 , n48885 , n48984 );
xor ( n49012 , n49011 , n48987 );
and ( n49013 , n49010 , n49012 );
xor ( n49014 , n48774 , n48790 );
xor ( n49015 , n49014 , n48807 );
xor ( n49016 , n48813 , n48815 );
xor ( n49017 , n49016 , n48818 );
and ( n49018 , n49015 , n49017 );
xor ( n49019 , n48778 , n48782 );
xor ( n49020 , n49019 , n48787 );
xor ( n49021 , n48795 , n48799 );
xor ( n49022 , n49021 , n48804 );
and ( n49023 , n49020 , n49022 );
and ( n49024 , n46510 , n39984 );
and ( n49025 , n46159 , n39982 );
nor ( n49026 , n49024 , n49025 );
xnor ( n49027 , n49026 , n39865 );
buf ( n49028 , n30382 );
not ( n49029 , n49028 );
and ( n49030 , n49027 , n49029 );
xnor ( n49031 , n48920 , n48924 );
and ( n49032 , n49029 , n49031 );
and ( n49033 , n49027 , n49031 );
or ( n49034 , n49030 , n49032 , n49033 );
and ( n49035 , n49022 , n49034 );
and ( n49036 , n49020 , n49034 );
or ( n49037 , n49023 , n49035 , n49036 );
and ( n49038 , n49017 , n49037 );
and ( n49039 , n49015 , n49037 );
or ( n49040 , n49018 , n49038 , n49039 );
and ( n49041 , n43387 , n42079 );
and ( n49042 , n43322 , n42076 );
nor ( n49043 , n49041 , n49042 );
xnor ( n49044 , n49043 , n41370 );
and ( n49045 , n43549 , n41981 );
and ( n49046 , n43524 , n41979 );
nor ( n49047 , n49045 , n49046 );
xnor ( n49048 , n49047 , n41373 );
and ( n49049 , n49044 , n49048 );
and ( n49050 , n43679 , n41522 );
and ( n49051 , n43671 , n41520 );
nor ( n49052 , n49050 , n49051 );
xnor ( n49053 , n49052 , n41100 );
and ( n49054 , n49048 , n49053 );
and ( n49055 , n49044 , n49053 );
or ( n49056 , n49049 , n49054 , n49055 );
and ( n49057 , n44000 , n41230 );
and ( n49058 , n43820 , n41228 );
nor ( n49059 , n49057 , n49058 );
xnor ( n49060 , n49059 , n40981 );
and ( n49061 , n44347 , n40928 );
and ( n49062 , n44318 , n40926 );
nor ( n49063 , n49061 , n49062 );
xnor ( n49064 , n49063 , n40688 );
and ( n49065 , n49060 , n49064 );
and ( n49066 , n45057 , n40666 );
and ( n49067 , n44826 , n40664 );
nor ( n49068 , n49066 , n49067 );
xnor ( n49069 , n49068 , n40445 );
and ( n49070 , n49064 , n49069 );
and ( n49071 , n49060 , n49069 );
or ( n49072 , n49065 , n49070 , n49071 );
and ( n49073 , n49056 , n49072 );
and ( n49074 , n45754 , n40406 );
and ( n49075 , n45171 , n40404 );
nor ( n49076 , n49074 , n49075 );
xnor ( n49077 , n49076 , n40262 );
and ( n49078 , n46159 , n40168 );
and ( n49079 , n46069 , n40166 );
nor ( n49080 , n49078 , n49079 );
xnor ( n49081 , n49080 , n40059 );
and ( n49082 , n49077 , n49081 );
buf ( n49083 , n30383 );
not ( n49084 , n49083 );
and ( n49085 , n49081 , n49084 );
and ( n49086 , n49077 , n49084 );
or ( n49087 , n49082 , n49085 , n49086 );
and ( n49088 , n49072 , n49087 );
and ( n49089 , n49056 , n49087 );
or ( n49090 , n49073 , n49088 , n49089 );
xor ( n49091 , n48550 , n48900 );
xor ( n49092 , n49091 , n48902 );
and ( n49093 , n49090 , n49092 );
xor ( n49094 , n48916 , n48925 );
xor ( n49095 , n49094 , n48942 );
and ( n49096 , n49092 , n49095 );
and ( n49097 , n49090 , n49095 );
or ( n49098 , n49093 , n49096 , n49097 );
xor ( n49099 , n48896 , n48897 );
xor ( n49100 , n49099 , n48905 );
and ( n49101 , n49098 , n49100 );
xor ( n49102 , n48945 , n48969 );
xor ( n49103 , n49102 , n48972 );
and ( n49104 , n49100 , n49103 );
and ( n49105 , n49098 , n49103 );
or ( n49106 , n49101 , n49104 , n49105 );
and ( n49107 , n49040 , n49106 );
xor ( n49108 , n48908 , n48975 );
xor ( n49109 , n49108 , n48978 );
and ( n49110 , n49106 , n49109 );
and ( n49111 , n49040 , n49109 );
or ( n49112 , n49107 , n49110 , n49111 );
xor ( n49113 , n48887 , n48893 );
xor ( n49114 , n49113 , n48981 );
and ( n49115 , n49112 , n49114 );
xor ( n49116 , n48961 , n48963 );
xor ( n49117 , n49116 , n48966 );
xor ( n49118 , n48911 , n48915 );
and ( n49119 , n48069 , n39382 );
not ( n49120 , n49119 );
and ( n49121 , n49120 , n39367 );
and ( n49122 , n48069 , n39384 );
and ( n49123 , n48077 , n39382 );
nor ( n49124 , n49122 , n49123 );
xnor ( n49125 , n49124 , n39367 );
and ( n49126 , n49121 , n49125 );
and ( n49127 , n48077 , n39384 );
and ( n49128 , n48086 , n39382 );
nor ( n49129 , n49127 , n49128 );
xnor ( n49130 , n49129 , n39367 );
and ( n49131 , n49126 , n49130 );
and ( n49132 , n49130 , n48909 );
and ( n49133 , n49126 , n48909 );
or ( n49134 , n49131 , n49132 , n49133 );
and ( n49135 , n49118 , n49134 );
and ( n49136 , n48086 , n39384 );
and ( n49137 , n48099 , n39382 );
nor ( n49138 , n49136 , n49137 );
xnor ( n49139 , n49138 , n39367 );
and ( n49140 , n49134 , n49139 );
and ( n49141 , n49118 , n49139 );
or ( n49142 , n49135 , n49140 , n49141 );
and ( n49143 , n49117 , n49142 );
xor ( n49144 , n48930 , n48934 );
xor ( n49145 , n49144 , n48939 );
xor ( n49146 , n48949 , n48953 );
xor ( n49147 , n49146 , n48958 );
and ( n49148 , n49145 , n49147 );
and ( n49149 , n46069 , n40406 );
and ( n49150 , n45754 , n40404 );
nor ( n49151 , n49149 , n49150 );
xnor ( n49152 , n49151 , n40262 );
buf ( n49153 , n30384 );
not ( n49154 , n49153 );
and ( n49155 , n49152 , n49154 );
and ( n49156 , n43524 , n42079 );
and ( n49157 , n43387 , n42076 );
nor ( n49158 , n49156 , n49157 );
xnor ( n49159 , n49158 , n41370 );
and ( n49160 , n43671 , n41981 );
and ( n49161 , n43549 , n41979 );
nor ( n49162 , n49160 , n49161 );
xnor ( n49163 , n49162 , n41373 );
and ( n49164 , n49159 , n49163 );
and ( n49165 , n43820 , n41522 );
and ( n49166 , n43679 , n41520 );
nor ( n49167 , n49165 , n49166 );
xnor ( n49168 , n49167 , n41100 );
and ( n49169 , n49163 , n49168 );
and ( n49170 , n49159 , n49168 );
or ( n49171 , n49164 , n49169 , n49170 );
and ( n49172 , n49155 , n49171 );
and ( n49173 , n44318 , n41230 );
and ( n49174 , n44000 , n41228 );
nor ( n49175 , n49173 , n49174 );
xnor ( n49176 , n49175 , n40981 );
and ( n49177 , n44826 , n40928 );
and ( n49178 , n44347 , n40926 );
nor ( n49179 , n49177 , n49178 );
xnor ( n49180 , n49179 , n40688 );
and ( n49181 , n49176 , n49180 );
and ( n49182 , n45171 , n40666 );
and ( n49183 , n45057 , n40664 );
nor ( n49184 , n49182 , n49183 );
xnor ( n49185 , n49184 , n40445 );
and ( n49186 , n49180 , n49185 );
and ( n49187 , n49176 , n49185 );
or ( n49188 , n49181 , n49186 , n49187 );
and ( n49189 , n49171 , n49188 );
and ( n49190 , n49155 , n49188 );
or ( n49191 , n49172 , n49189 , n49190 );
and ( n49192 , n49147 , n49191 );
and ( n49193 , n49145 , n49191 );
or ( n49194 , n49148 , n49192 , n49193 );
and ( n49195 , n49142 , n49194 );
and ( n49196 , n49117 , n49194 );
or ( n49197 , n49143 , n49195 , n49196 );
xor ( n49198 , n49044 , n49048 );
xor ( n49199 , n49198 , n49053 );
xor ( n49200 , n49060 , n49064 );
xor ( n49201 , n49200 , n49069 );
and ( n49202 , n49199 , n49201 );
xor ( n49203 , n49077 , n49081 );
xor ( n49204 , n49203 , n49084 );
and ( n49205 , n49201 , n49204 );
and ( n49206 , n49199 , n49204 );
or ( n49207 , n49202 , n49205 , n49206 );
xor ( n49208 , n49027 , n49029 );
xor ( n49209 , n49208 , n49031 );
and ( n49210 , n49207 , n49209 );
xor ( n49211 , n49056 , n49072 );
xor ( n49212 , n49211 , n49087 );
and ( n49213 , n49209 , n49212 );
and ( n49214 , n49207 , n49212 );
or ( n49215 , n49210 , n49213 , n49214 );
xor ( n49216 , n49020 , n49022 );
xor ( n49217 , n49216 , n49034 );
and ( n49218 , n49215 , n49217 );
xor ( n49219 , n49090 , n49092 );
xor ( n49220 , n49219 , n49095 );
and ( n49221 , n49217 , n49220 );
and ( n49222 , n49215 , n49220 );
or ( n49223 , n49218 , n49221 , n49222 );
and ( n49224 , n49197 , n49223 );
xor ( n49225 , n49015 , n49017 );
xor ( n49226 , n49225 , n49037 );
and ( n49227 , n49223 , n49226 );
and ( n49228 , n49197 , n49226 );
or ( n49229 , n49224 , n49227 , n49228 );
xor ( n49230 , n49000 , n49002 );
xor ( n49231 , n49230 , n49004 );
and ( n49232 , n49229 , n49231 );
xor ( n49233 , n49040 , n49106 );
xor ( n49234 , n49233 , n49109 );
and ( n49235 , n49231 , n49234 );
and ( n49236 , n49229 , n49234 );
or ( n49237 , n49232 , n49235 , n49236 );
and ( n49238 , n49114 , n49237 );
and ( n49239 , n49112 , n49237 );
or ( n49240 , n49115 , n49238 , n49239 );
and ( n49241 , n49012 , n49240 );
and ( n49242 , n49010 , n49240 );
or ( n49243 , n49013 , n49241 , n49242 );
and ( n49244 , n48992 , n49243 );
and ( n49245 , n48990 , n49243 );
or ( n49246 , n48993 , n49244 , n49245 );
and ( n49247 , n48882 , n49246 );
and ( n49248 , n48880 , n49246 );
or ( n49249 , n48883 , n49247 , n49248 );
or ( n49250 , n48878 , n49249 );
or ( n49251 , n48876 , n49250 );
and ( n49252 , n48873 , n49251 );
and ( n49253 , n48871 , n49251 );
or ( n49254 , n48874 , n49252 , n49253 );
and ( n49255 , n48400 , n49254 );
xor ( n49256 , n48400 , n49254 );
xor ( n49257 , n48871 , n48873 );
xor ( n49258 , n49257 , n49251 );
not ( n49259 , n49258 );
xnor ( n49260 , n48876 , n49250 );
xnor ( n49261 , n48878 , n49249 );
xor ( n49262 , n48880 , n48882 );
xor ( n49263 , n49262 , n49246 );
xor ( n49264 , n48990 , n48992 );
xor ( n49265 , n49264 , n49243 );
xor ( n49266 , n49010 , n49012 );
xor ( n49267 , n49266 , n49240 );
xor ( n49268 , n48995 , n48997 );
xor ( n49269 , n49268 , n49007 );
xor ( n49270 , n49112 , n49114 );
xor ( n49271 , n49270 , n49237 );
and ( n49272 , n49269 , n49271 );
xor ( n49273 , n49098 , n49100 );
xor ( n49274 , n49273 , n49103 );
and ( n49275 , n46510 , n40168 );
and ( n49276 , n46159 , n40166 );
nor ( n49277 , n49275 , n49276 );
xnor ( n49278 , n49277 , n40059 );
xor ( n49279 , n49152 , n49154 );
and ( n49280 , n49278 , n49279 );
and ( n49281 , n43549 , n42079 );
and ( n49282 , n43524 , n42076 );
nor ( n49283 , n49281 , n49282 );
xnor ( n49284 , n49283 , n41370 );
and ( n49285 , n43679 , n41981 );
and ( n49286 , n43671 , n41979 );
nor ( n49287 , n49285 , n49286 );
xnor ( n49288 , n49287 , n41373 );
and ( n49289 , n49284 , n49288 );
and ( n49290 , n44000 , n41522 );
and ( n49291 , n43820 , n41520 );
nor ( n49292 , n49290 , n49291 );
xnor ( n49293 , n49292 , n41100 );
and ( n49294 , n49288 , n49293 );
and ( n49295 , n49284 , n49293 );
or ( n49296 , n49289 , n49294 , n49295 );
and ( n49297 , n49279 , n49296 );
and ( n49298 , n49278 , n49296 );
or ( n49299 , n49280 , n49297 , n49298 );
and ( n49300 , n44347 , n41230 );
and ( n49301 , n44318 , n41228 );
nor ( n49302 , n49300 , n49301 );
xnor ( n49303 , n49302 , n40981 );
and ( n49304 , n45057 , n40928 );
and ( n49305 , n44826 , n40926 );
nor ( n49306 , n49304 , n49305 );
xnor ( n49307 , n49306 , n40688 );
and ( n49308 , n49303 , n49307 );
and ( n49309 , n45754 , n40666 );
and ( n49310 , n45171 , n40664 );
nor ( n49311 , n49309 , n49310 );
xnor ( n49312 , n49311 , n40445 );
and ( n49313 , n49307 , n49312 );
and ( n49314 , n49303 , n49312 );
or ( n49315 , n49308 , n49313 , n49314 );
and ( n49316 , n46159 , n40406 );
and ( n49317 , n46069 , n40404 );
nor ( n49318 , n49316 , n49317 );
xnor ( n49319 , n49318 , n40262 );
and ( n49320 , n46676 , n40168 );
and ( n49321 , n46510 , n40166 );
nor ( n49322 , n49320 , n49321 );
xnor ( n49323 , n49322 , n40059 );
and ( n49324 , n49319 , n49323 );
and ( n49325 , n46948 , n39984 );
and ( n49326 , n46777 , n39982 );
nor ( n49327 , n49325 , n49326 );
xnor ( n49328 , n49327 , n39865 );
and ( n49329 , n49323 , n49328 );
and ( n49330 , n49319 , n49328 );
or ( n49331 , n49324 , n49329 , n49330 );
and ( n49332 , n49315 , n49331 );
xor ( n49333 , n49159 , n49163 );
xor ( n49334 , n49333 , n49168 );
and ( n49335 , n49331 , n49334 );
and ( n49336 , n49315 , n49334 );
or ( n49337 , n49332 , n49335 , n49336 );
and ( n49338 , n49299 , n49337 );
xor ( n49339 , n49155 , n49171 );
xor ( n49340 , n49339 , n49188 );
and ( n49341 , n49337 , n49340 );
and ( n49342 , n49299 , n49340 );
or ( n49343 , n49338 , n49341 , n49342 );
xor ( n49344 , n49145 , n49147 );
xor ( n49345 , n49344 , n49191 );
and ( n49346 , n49343 , n49345 );
xor ( n49347 , n49207 , n49209 );
xor ( n49348 , n49347 , n49212 );
and ( n49349 , n49345 , n49348 );
and ( n49350 , n49343 , n49348 );
or ( n49351 , n49346 , n49349 , n49350 );
xor ( n49352 , n49117 , n49142 );
xor ( n49353 , n49352 , n49194 );
and ( n49354 , n49351 , n49353 );
xor ( n49355 , n49215 , n49217 );
xor ( n49356 , n49355 , n49220 );
and ( n49357 , n49353 , n49356 );
and ( n49358 , n49351 , n49356 );
or ( n49359 , n49354 , n49357 , n49358 );
and ( n49360 , n49274 , n49359 );
xor ( n49361 , n49197 , n49223 );
xor ( n49362 , n49361 , n49226 );
and ( n49363 , n49359 , n49362 );
and ( n49364 , n49274 , n49362 );
or ( n49365 , n49360 , n49363 , n49364 );
xor ( n49366 , n49229 , n49231 );
xor ( n49367 , n49366 , n49234 );
and ( n49368 , n49365 , n49367 );
xor ( n49369 , n49274 , n49359 );
xor ( n49370 , n49369 , n49362 );
xor ( n49371 , n49121 , n49125 );
and ( n49372 , n48069 , n39530 );
not ( n49373 , n49372 );
and ( n49374 , n49373 , n39497 );
and ( n49375 , n48069 , n39532 );
and ( n49376 , n48077 , n39530 );
nor ( n49377 , n49375 , n49376 );
xnor ( n49378 , n49377 , n39497 );
and ( n49379 , n49374 , n49378 );
and ( n49380 , n48077 , n39532 );
and ( n49381 , n48086 , n39530 );
nor ( n49382 , n49380 , n49381 );
xnor ( n49383 , n49382 , n39497 );
and ( n49384 , n49379 , n49383 );
and ( n49385 , n49383 , n49119 );
and ( n49386 , n49379 , n49119 );
or ( n49387 , n49384 , n49385 , n49386 );
and ( n49388 , n49371 , n49387 );
and ( n49389 , n48086 , n39532 );
and ( n49390 , n48099 , n39530 );
nor ( n49391 , n49389 , n49390 );
xnor ( n49392 , n49391 , n39497 );
and ( n49393 , n49387 , n49392 );
and ( n49394 , n49371 , n49392 );
or ( n49395 , n49388 , n49393 , n49394 );
and ( n49396 , n48099 , n39532 );
and ( n49397 , n47927 , n39530 );
nor ( n49398 , n49396 , n49397 );
xnor ( n49399 , n49398 , n39497 );
and ( n49400 , n49395 , n49399 );
xor ( n49401 , n49126 , n49130 );
xor ( n49402 , n49401 , n48909 );
and ( n49403 , n49399 , n49402 );
and ( n49404 , n49395 , n49402 );
or ( n49405 , n49400 , n49403 , n49404 );
and ( n49406 , n47927 , n39532 );
and ( n49407 , n47932 , n39530 );
nor ( n49408 , n49406 , n49407 );
xnor ( n49409 , n49408 , n39497 );
and ( n49410 , n49405 , n49409 );
xor ( n49411 , n49118 , n49134 );
xor ( n49412 , n49411 , n49139 );
and ( n49413 , n49409 , n49412 );
and ( n49414 , n49405 , n49412 );
or ( n49415 , n49410 , n49413 , n49414 );
xor ( n49416 , n49351 , n49353 );
xor ( n49417 , n49416 , n49356 );
and ( n49418 , n49415 , n49417 );
xor ( n49419 , n49374 , n49378 );
and ( n49420 , n48069 , n39663 );
not ( n49421 , n49420 );
and ( n49422 , n49421 , n39608 );
and ( n49423 , n48069 , n39665 );
and ( n49424 , n48077 , n39663 );
nor ( n49425 , n49423 , n49424 );
xnor ( n49426 , n49425 , n39608 );
and ( n49427 , n49422 , n49426 );
and ( n49428 , n48077 , n39665 );
and ( n49429 , n48086 , n39663 );
nor ( n49430 , n49428 , n49429 );
xnor ( n49431 , n49430 , n39608 );
and ( n49432 , n49427 , n49431 );
and ( n49433 , n49431 , n49372 );
and ( n49434 , n49427 , n49372 );
or ( n49435 , n49432 , n49433 , n49434 );
and ( n49436 , n49419 , n49435 );
and ( n49437 , n48086 , n39665 );
and ( n49438 , n48099 , n39663 );
nor ( n49439 , n49437 , n49438 );
xnor ( n49440 , n49439 , n39608 );
and ( n49441 , n49435 , n49440 );
and ( n49442 , n49419 , n49440 );
or ( n49443 , n49436 , n49441 , n49442 );
and ( n49444 , n48099 , n39665 );
and ( n49445 , n47927 , n39663 );
nor ( n49446 , n49444 , n49445 );
xnor ( n49447 , n49446 , n39608 );
and ( n49448 , n49443 , n49447 );
xor ( n49449 , n49379 , n49383 );
xor ( n49450 , n49449 , n49119 );
and ( n49451 , n49447 , n49450 );
and ( n49452 , n49443 , n49450 );
or ( n49453 , n49448 , n49451 , n49452 );
and ( n49454 , n47927 , n39665 );
and ( n49455 , n47932 , n39663 );
nor ( n49456 , n49454 , n49455 );
xnor ( n49457 , n49456 , n39608 );
and ( n49458 , n49453 , n49457 );
xor ( n49459 , n49371 , n49387 );
xor ( n49460 , n49459 , n49392 );
and ( n49461 , n49457 , n49460 );
and ( n49462 , n49453 , n49460 );
or ( n49463 , n49458 , n49461 , n49462 );
and ( n49464 , n47932 , n39665 );
and ( n49465 , n47645 , n39663 );
nor ( n49466 , n49464 , n49465 );
xnor ( n49467 , n49466 , n39608 );
and ( n49468 , n49463 , n49467 );
xor ( n49469 , n49395 , n49399 );
xor ( n49470 , n49469 , n49402 );
and ( n49471 , n49467 , n49470 );
and ( n49472 , n49463 , n49470 );
or ( n49473 , n49468 , n49471 , n49472 );
and ( n49474 , n47645 , n39665 );
and ( n49475 , n46948 , n39663 );
nor ( n49476 , n49474 , n49475 );
xnor ( n49477 , n49476 , n39608 );
and ( n49478 , n49473 , n49477 );
xor ( n49479 , n49405 , n49409 );
xor ( n49480 , n49479 , n49412 );
and ( n49481 , n49477 , n49480 );
and ( n49482 , n49473 , n49480 );
or ( n49483 , n49478 , n49481 , n49482 );
and ( n49484 , n49417 , n49483 );
and ( n49485 , n49415 , n49483 );
or ( n49486 , n49418 , n49484 , n49485 );
and ( n49487 , n49370 , n49486 );
xor ( n49488 , n49415 , n49417 );
xor ( n49489 , n49488 , n49483 );
xor ( n49490 , n49422 , n49426 );
and ( n49491 , n48069 , n39793 );
not ( n49492 , n49491 );
and ( n49493 , n49492 , n39729 );
and ( n49494 , n48069 , n39795 );
and ( n49495 , n48077 , n39793 );
nor ( n49496 , n49494 , n49495 );
xnor ( n49497 , n49496 , n39729 );
and ( n49498 , n49493 , n49497 );
and ( n49499 , n48077 , n39795 );
and ( n49500 , n48086 , n39793 );
nor ( n49501 , n49499 , n49500 );
xnor ( n49502 , n49501 , n39729 );
and ( n49503 , n49498 , n49502 );
and ( n49504 , n49502 , n49420 );
and ( n49505 , n49498 , n49420 );
or ( n49506 , n49503 , n49504 , n49505 );
and ( n49507 , n49490 , n49506 );
and ( n49508 , n48086 , n39795 );
and ( n49509 , n48099 , n39793 );
nor ( n49510 , n49508 , n49509 );
xnor ( n49511 , n49510 , n39729 );
and ( n49512 , n49506 , n49511 );
and ( n49513 , n49490 , n49511 );
or ( n49514 , n49507 , n49512 , n49513 );
and ( n49515 , n48099 , n39795 );
and ( n49516 , n47927 , n39793 );
nor ( n49517 , n49515 , n49516 );
xnor ( n49518 , n49517 , n39729 );
and ( n49519 , n49514 , n49518 );
xor ( n49520 , n49427 , n49431 );
xor ( n49521 , n49520 , n49372 );
and ( n49522 , n49518 , n49521 );
and ( n49523 , n49514 , n49521 );
or ( n49524 , n49519 , n49522 , n49523 );
and ( n49525 , n47927 , n39795 );
and ( n49526 , n47932 , n39793 );
nor ( n49527 , n49525 , n49526 );
xnor ( n49528 , n49527 , n39729 );
and ( n49529 , n49524 , n49528 );
xor ( n49530 , n49419 , n49435 );
xor ( n49531 , n49530 , n49440 );
and ( n49532 , n49528 , n49531 );
and ( n49533 , n49524 , n49531 );
or ( n49534 , n49529 , n49532 , n49533 );
and ( n49535 , n47932 , n39795 );
and ( n49536 , n47645 , n39793 );
nor ( n49537 , n49535 , n49536 );
xnor ( n49538 , n49537 , n39729 );
and ( n49539 , n49534 , n49538 );
xor ( n49540 , n49443 , n49447 );
xor ( n49541 , n49540 , n49450 );
and ( n49542 , n49538 , n49541 );
and ( n49543 , n49534 , n49541 );
or ( n49544 , n49539 , n49542 , n49543 );
and ( n49545 , n47645 , n39795 );
and ( n49546 , n46948 , n39793 );
nor ( n49547 , n49545 , n49546 );
xnor ( n49548 , n49547 , n39729 );
and ( n49549 , n49544 , n49548 );
xor ( n49550 , n49453 , n49457 );
xor ( n49551 , n49550 , n49460 );
and ( n49552 , n49548 , n49551 );
and ( n49553 , n49544 , n49551 );
or ( n49554 , n49549 , n49552 , n49553 );
and ( n49555 , n46948 , n39795 );
and ( n49556 , n46777 , n39793 );
nor ( n49557 , n49555 , n49556 );
xnor ( n49558 , n49557 , n39729 );
and ( n49559 , n49554 , n49558 );
xor ( n49560 , n49463 , n49467 );
xor ( n49561 , n49560 , n49470 );
and ( n49562 , n49558 , n49561 );
and ( n49563 , n49554 , n49561 );
or ( n49564 , n49559 , n49562 , n49563 );
and ( n49565 , n46777 , n39795 );
and ( n49566 , n46676 , n39793 );
nor ( n49567 , n49565 , n49566 );
xnor ( n49568 , n49567 , n39729 );
and ( n49569 , n49564 , n49568 );
xor ( n49570 , n49473 , n49477 );
xor ( n49571 , n49570 , n49480 );
and ( n49572 , n49568 , n49571 );
and ( n49573 , n49564 , n49571 );
or ( n49574 , n49569 , n49572 , n49573 );
and ( n49575 , n49489 , n49574 );
xor ( n49576 , n49199 , n49201 );
xor ( n49577 , n49576 , n49204 );
xor ( n49578 , n49176 , n49180 );
xor ( n49579 , n49578 , n49185 );
buf ( n49580 , n30385 );
not ( n49581 , n49580 );
and ( n49582 , n43671 , n42079 );
and ( n49583 , n43549 , n42076 );
nor ( n49584 , n49582 , n49583 );
xnor ( n49585 , n49584 , n41370 );
and ( n49586 , n45171 , n40928 );
and ( n49587 , n45057 , n40926 );
nor ( n49588 , n49586 , n49587 );
xnor ( n49589 , n49588 , n40688 );
and ( n49590 , n49585 , n49589 );
and ( n49591 , n46069 , n40666 );
and ( n49592 , n45754 , n40664 );
nor ( n49593 , n49591 , n49592 );
xnor ( n49594 , n49593 , n40445 );
and ( n49595 , n49589 , n49594 );
and ( n49596 , n49585 , n49594 );
or ( n49597 , n49590 , n49595 , n49596 );
and ( n49598 , n49581 , n49597 );
and ( n49599 , n46510 , n40406 );
and ( n49600 , n46159 , n40404 );
nor ( n49601 , n49599 , n49600 );
xnor ( n49602 , n49601 , n40262 );
and ( n49603 , n46777 , n40168 );
and ( n49604 , n46676 , n40166 );
nor ( n49605 , n49603 , n49604 );
xnor ( n49606 , n49605 , n40059 );
and ( n49607 , n49602 , n49606 );
and ( n49608 , n47645 , n39984 );
and ( n49609 , n46948 , n39982 );
nor ( n49610 , n49608 , n49609 );
xnor ( n49611 , n49610 , n39865 );
and ( n49612 , n49606 , n49611 );
and ( n49613 , n49602 , n49611 );
or ( n49614 , n49607 , n49612 , n49613 );
and ( n49615 , n49597 , n49614 );
and ( n49616 , n49581 , n49614 );
or ( n49617 , n49598 , n49615 , n49616 );
and ( n49618 , n49579 , n49617 );
xor ( n49619 , n49284 , n49288 );
xor ( n49620 , n49619 , n49293 );
xor ( n49621 , n49303 , n49307 );
xor ( n49622 , n49621 , n49312 );
and ( n49623 , n49620 , n49622 );
xor ( n49624 , n49319 , n49323 );
xor ( n49625 , n49624 , n49328 );
and ( n49626 , n49622 , n49625 );
and ( n49627 , n49620 , n49625 );
or ( n49628 , n49623 , n49626 , n49627 );
and ( n49629 , n49617 , n49628 );
and ( n49630 , n49579 , n49628 );
or ( n49631 , n49618 , n49629 , n49630 );
and ( n49632 , n49577 , n49631 );
xor ( n49633 , n49299 , n49337 );
xor ( n49634 , n49633 , n49340 );
and ( n49635 , n49631 , n49634 );
and ( n49636 , n49577 , n49634 );
or ( n49637 , n49632 , n49635 , n49636 );
xor ( n49638 , n49343 , n49345 );
xor ( n49639 , n49638 , n49348 );
and ( n49640 , n49637 , n49639 );
xor ( n49641 , n49564 , n49568 );
xor ( n49642 , n49641 , n49571 );
and ( n49643 , n49639 , n49642 );
and ( n49644 , n49637 , n49642 );
or ( n49645 , n49640 , n49643 , n49644 );
and ( n49646 , n49574 , n49645 );
and ( n49647 , n49489 , n49645 );
or ( n49648 , n49575 , n49646 , n49647 );
and ( n49649 , n49486 , n49648 );
and ( n49650 , n49370 , n49648 );
or ( n49651 , n49487 , n49649 , n49650 );
and ( n49652 , n49367 , n49651 );
and ( n49653 , n49365 , n49651 );
or ( n49654 , n49368 , n49652 , n49653 );
and ( n49655 , n49271 , n49654 );
and ( n49656 , n49269 , n49654 );
or ( n49657 , n49272 , n49655 , n49656 );
or ( n49658 , n49267 , n49657 );
and ( n49659 , n49265 , n49658 );
xor ( n49660 , n49265 , n49658 );
xnor ( n49661 , n49267 , n49657 );
xor ( n49662 , n49269 , n49271 );
xor ( n49663 , n49662 , n49654 );
xor ( n49664 , n49365 , n49367 );
xor ( n49665 , n49664 , n49651 );
xor ( n49666 , n49370 , n49486 );
xor ( n49667 , n49666 , n49648 );
and ( n49668 , n46676 , n39984 );
and ( n49669 , n46510 , n39982 );
nor ( n49670 , n49668 , n49669 );
xnor ( n49671 , n49670 , n39865 );
xor ( n49672 , n49554 , n49558 );
xor ( n49673 , n49672 , n49561 );
and ( n49674 , n49671 , n49673 );
xor ( n49675 , n49278 , n49279 );
xor ( n49676 , n49675 , n49296 );
xor ( n49677 , n49315 , n49331 );
xor ( n49678 , n49677 , n49334 );
and ( n49679 , n49676 , n49678 );
buf ( n49680 , n30386 );
not ( n49681 , n49680 );
xor ( n49682 , n49585 , n49589 );
xor ( n49683 , n49682 , n49594 );
and ( n49684 , n49681 , n49683 );
xor ( n49685 , n49602 , n49606 );
xor ( n49686 , n49685 , n49611 );
and ( n49687 , n49683 , n49686 );
and ( n49688 , n49681 , n49686 );
or ( n49689 , n49684 , n49687 , n49688 );
xor ( n49690 , n49581 , n49597 );
xor ( n49691 , n49690 , n49614 );
and ( n49692 , n49689 , n49691 );
xor ( n49693 , n49620 , n49622 );
xor ( n49694 , n49693 , n49625 );
and ( n49695 , n49691 , n49694 );
and ( n49696 , n49689 , n49694 );
or ( n49697 , n49692 , n49695 , n49696 );
and ( n49698 , n49678 , n49697 );
and ( n49699 , n49676 , n49697 );
or ( n49700 , n49679 , n49698 , n49699 );
xor ( n49701 , n49577 , n49631 );
xor ( n49702 , n49701 , n49634 );
and ( n49703 , n49700 , n49702 );
and ( n49704 , n46777 , n39984 );
and ( n49705 , n46676 , n39982 );
nor ( n49706 , n49704 , n49705 );
xnor ( n49707 , n49706 , n39865 );
xor ( n49708 , n49544 , n49548 );
xor ( n49709 , n49708 , n49551 );
and ( n49710 , n49707 , n49709 );
and ( n49711 , n49702 , n49710 );
and ( n49712 , n49700 , n49710 );
or ( n49713 , n49703 , n49711 , n49712 );
and ( n49714 , n49674 , n49713 );
xor ( n49715 , n49671 , n49673 );
xor ( n49716 , n49579 , n49617 );
xor ( n49717 , n49716 , n49628 );
xor ( n49718 , n49676 , n49678 );
xor ( n49719 , n49718 , n49697 );
and ( n49720 , n49717 , n49719 );
xor ( n49721 , n49707 , n49709 );
and ( n49722 , n49719 , n49721 );
and ( n49723 , n49717 , n49721 );
or ( n49724 , n49720 , n49722 , n49723 );
and ( n49725 , n49715 , n49724 );
xor ( n49726 , n49700 , n49702 );
xor ( n49727 , n49726 , n49710 );
and ( n49728 , n49724 , n49727 );
and ( n49729 , n49715 , n49727 );
or ( n49730 , n49725 , n49728 , n49729 );
and ( n49731 , n49713 , n49730 );
and ( n49732 , n49674 , n49730 );
or ( n49733 , n49714 , n49731 , n49732 );
xor ( n49734 , n49489 , n49574 );
xor ( n49735 , n49734 , n49645 );
and ( n49736 , n49733 , n49735 );
xor ( n49737 , n49637 , n49639 );
xor ( n49738 , n49737 , n49642 );
xor ( n49739 , n49674 , n49713 );
xor ( n49740 , n49739 , n49730 );
and ( n49741 , n49738 , n49740 );
xor ( n49742 , n49715 , n49724 );
xor ( n49743 , n49742 , n49727 );
xor ( n49744 , n49689 , n49691 );
xor ( n49745 , n49744 , n49694 );
xor ( n49746 , n49534 , n49538 );
xor ( n49747 , n49746 , n49541 );
and ( n49748 , n49745 , n49747 );
xor ( n49749 , n49493 , n49497 );
and ( n49750 , n48069 , n39982 );
not ( n49751 , n49750 );
and ( n49752 , n49751 , n39865 );
and ( n49753 , n48069 , n39984 );
and ( n49754 , n48077 , n39982 );
nor ( n49755 , n49753 , n49754 );
xnor ( n49756 , n49755 , n39865 );
and ( n49757 , n49752 , n49756 );
and ( n49758 , n48077 , n39984 );
and ( n49759 , n48086 , n39982 );
nor ( n49760 , n49758 , n49759 );
xnor ( n49761 , n49760 , n39865 );
and ( n49762 , n49757 , n49761 );
and ( n49763 , n49761 , n49491 );
and ( n49764 , n49757 , n49491 );
or ( n49765 , n49762 , n49763 , n49764 );
and ( n49766 , n49749 , n49765 );
and ( n49767 , n48086 , n39984 );
and ( n49768 , n48099 , n39982 );
nor ( n49769 , n49767 , n49768 );
xnor ( n49770 , n49769 , n39865 );
and ( n49771 , n49765 , n49770 );
and ( n49772 , n49749 , n49770 );
or ( n49773 , n49766 , n49771 , n49772 );
and ( n49774 , n48099 , n39984 );
and ( n49775 , n47927 , n39982 );
nor ( n49776 , n49774 , n49775 );
xnor ( n49777 , n49776 , n39865 );
and ( n49778 , n49773 , n49777 );
xor ( n49779 , n49498 , n49502 );
xor ( n49780 , n49779 , n49420 );
and ( n49781 , n49777 , n49780 );
and ( n49782 , n49773 , n49780 );
or ( n49783 , n49778 , n49781 , n49782 );
and ( n49784 , n47927 , n39984 );
and ( n49785 , n47932 , n39982 );
nor ( n49786 , n49784 , n49785 );
xnor ( n49787 , n49786 , n39865 );
and ( n49788 , n49783 , n49787 );
xor ( n49789 , n49490 , n49506 );
xor ( n49790 , n49789 , n49511 );
and ( n49791 , n49787 , n49790 );
and ( n49792 , n49783 , n49790 );
or ( n49793 , n49788 , n49791 , n49792 );
and ( n49794 , n47932 , n39984 );
and ( n49795 , n47645 , n39982 );
nor ( n49796 , n49794 , n49795 );
xnor ( n49797 , n49796 , n39865 );
and ( n49798 , n49793 , n49797 );
xor ( n49799 , n49514 , n49518 );
xor ( n49800 , n49799 , n49521 );
and ( n49801 , n49797 , n49800 );
and ( n49802 , n49793 , n49800 );
or ( n49803 , n49798 , n49801 , n49802 );
xor ( n49804 , n49524 , n49528 );
xor ( n49805 , n49804 , n49531 );
and ( n49806 , n49803 , n49805 );
and ( n49807 , n49747 , n49806 );
and ( n49808 , n49745 , n49806 );
or ( n49809 , n49748 , n49807 , n49808 );
xor ( n49810 , n49717 , n49719 );
xor ( n49811 , n49810 , n49721 );
and ( n49812 , n49809 , n49811 );
xor ( n49813 , n49745 , n49747 );
xor ( n49814 , n49813 , n49806 );
xor ( n49815 , n49681 , n49683 );
xor ( n49816 , n49815 , n49686 );
xor ( n49817 , n49803 , n49805 );
and ( n49818 , n49816 , n49817 );
xor ( n49819 , n49752 , n49756 );
and ( n49820 , n48069 , n40166 );
not ( n49821 , n49820 );
and ( n49822 , n49821 , n40059 );
and ( n49823 , n48069 , n40168 );
and ( n49824 , n48077 , n40166 );
nor ( n49825 , n49823 , n49824 );
xnor ( n49826 , n49825 , n40059 );
and ( n49827 , n49822 , n49826 );
and ( n49828 , n48077 , n40168 );
and ( n49829 , n48086 , n40166 );
nor ( n49830 , n49828 , n49829 );
xnor ( n49831 , n49830 , n40059 );
and ( n49832 , n49827 , n49831 );
and ( n49833 , n49831 , n49750 );
and ( n49834 , n49827 , n49750 );
or ( n49835 , n49832 , n49833 , n49834 );
and ( n49836 , n49819 , n49835 );
and ( n49837 , n48086 , n40168 );
and ( n49838 , n48099 , n40166 );
nor ( n49839 , n49837 , n49838 );
xnor ( n49840 , n49839 , n40059 );
and ( n49841 , n49835 , n49840 );
and ( n49842 , n49819 , n49840 );
or ( n49843 , n49836 , n49841 , n49842 );
and ( n49844 , n48099 , n40168 );
and ( n49845 , n47927 , n40166 );
nor ( n49846 , n49844 , n49845 );
xnor ( n49847 , n49846 , n40059 );
and ( n49848 , n49843 , n49847 );
xor ( n49849 , n49757 , n49761 );
xor ( n49850 , n49849 , n49491 );
and ( n49851 , n49847 , n49850 );
and ( n49852 , n49843 , n49850 );
or ( n49853 , n49848 , n49851 , n49852 );
and ( n49854 , n47927 , n40168 );
and ( n49855 , n47932 , n40166 );
nor ( n49856 , n49854 , n49855 );
xnor ( n49857 , n49856 , n40059 );
and ( n49858 , n49853 , n49857 );
xor ( n49859 , n49749 , n49765 );
xor ( n49860 , n49859 , n49770 );
and ( n49861 , n49857 , n49860 );
and ( n49862 , n49853 , n49860 );
or ( n49863 , n49858 , n49861 , n49862 );
and ( n49864 , n47932 , n40168 );
and ( n49865 , n47645 , n40166 );
nor ( n49866 , n49864 , n49865 );
xnor ( n49867 , n49866 , n40059 );
and ( n49868 , n49863 , n49867 );
xor ( n49869 , n49773 , n49777 );
xor ( n49870 , n49869 , n49780 );
and ( n49871 , n49867 , n49870 );
and ( n49872 , n49863 , n49870 );
or ( n49873 , n49868 , n49871 , n49872 );
and ( n49874 , n47645 , n40168 );
and ( n49875 , n46948 , n40166 );
nor ( n49876 , n49874 , n49875 );
xnor ( n49877 , n49876 , n40059 );
and ( n49878 , n49873 , n49877 );
xor ( n49879 , n49783 , n49787 );
xor ( n49880 , n49879 , n49790 );
and ( n49881 , n49877 , n49880 );
and ( n49882 , n49873 , n49880 );
or ( n49883 , n49878 , n49881 , n49882 );
and ( n49884 , n46948 , n40168 );
and ( n49885 , n46777 , n40166 );
nor ( n49886 , n49884 , n49885 );
xnor ( n49887 , n49886 , n40059 );
and ( n49888 , n49883 , n49887 );
xor ( n49889 , n49793 , n49797 );
xor ( n49890 , n49889 , n49800 );
and ( n49891 , n49887 , n49890 );
and ( n49892 , n49883 , n49890 );
or ( n49893 , n49888 , n49891 , n49892 );
and ( n49894 , n49817 , n49893 );
and ( n49895 , n49816 , n49893 );
or ( n49896 , n49818 , n49894 , n49895 );
and ( n49897 , n49814 , n49896 );
xor ( n49898 , n49816 , n49817 );
xor ( n49899 , n49898 , n49893 );
xor ( n49900 , n49822 , n49826 );
and ( n49901 , n48069 , n40404 );
not ( n49902 , n49901 );
and ( n49903 , n49902 , n40262 );
and ( n49904 , n48069 , n40406 );
and ( n49905 , n48077 , n40404 );
nor ( n49906 , n49904 , n49905 );
xnor ( n49907 , n49906 , n40262 );
and ( n49908 , n49903 , n49907 );
and ( n49909 , n48077 , n40406 );
and ( n49910 , n48086 , n40404 );
nor ( n49911 , n49909 , n49910 );
xnor ( n49912 , n49911 , n40262 );
and ( n49913 , n49908 , n49912 );
and ( n49914 , n49912 , n49820 );
and ( n49915 , n49908 , n49820 );
or ( n49916 , n49913 , n49914 , n49915 );
and ( n49917 , n49900 , n49916 );
and ( n49918 , n48086 , n40406 );
and ( n49919 , n48099 , n40404 );
nor ( n49920 , n49918 , n49919 );
xnor ( n49921 , n49920 , n40262 );
and ( n49922 , n49916 , n49921 );
and ( n49923 , n49900 , n49921 );
or ( n49924 , n49917 , n49922 , n49923 );
and ( n49925 , n48099 , n40406 );
and ( n49926 , n47927 , n40404 );
nor ( n49927 , n49925 , n49926 );
xnor ( n49928 , n49927 , n40262 );
and ( n49929 , n49924 , n49928 );
xor ( n49930 , n49827 , n49831 );
xor ( n49931 , n49930 , n49750 );
and ( n49932 , n49928 , n49931 );
and ( n49933 , n49924 , n49931 );
or ( n49934 , n49929 , n49932 , n49933 );
and ( n49935 , n47927 , n40406 );
and ( n49936 , n47932 , n40404 );
nor ( n49937 , n49935 , n49936 );
xnor ( n49938 , n49937 , n40262 );
and ( n49939 , n49934 , n49938 );
xor ( n49940 , n49819 , n49835 );
xor ( n49941 , n49940 , n49840 );
and ( n49942 , n49938 , n49941 );
and ( n49943 , n49934 , n49941 );
or ( n49944 , n49939 , n49942 , n49943 );
and ( n49945 , n47932 , n40406 );
and ( n49946 , n47645 , n40404 );
nor ( n49947 , n49945 , n49946 );
xnor ( n49948 , n49947 , n40262 );
and ( n49949 , n49944 , n49948 );
xor ( n49950 , n49843 , n49847 );
xor ( n49951 , n49950 , n49850 );
and ( n49952 , n49948 , n49951 );
and ( n49953 , n49944 , n49951 );
or ( n49954 , n49949 , n49952 , n49953 );
and ( n49955 , n47645 , n40406 );
and ( n49956 , n46948 , n40404 );
nor ( n49957 , n49955 , n49956 );
xnor ( n49958 , n49957 , n40262 );
and ( n49959 , n49954 , n49958 );
xor ( n49960 , n49853 , n49857 );
xor ( n49961 , n49960 , n49860 );
and ( n49962 , n49958 , n49961 );
and ( n49963 , n49954 , n49961 );
or ( n49964 , n49959 , n49962 , n49963 );
and ( n49965 , n46948 , n40406 );
and ( n49966 , n46777 , n40404 );
nor ( n49967 , n49965 , n49966 );
xnor ( n49968 , n49967 , n40262 );
and ( n49969 , n49964 , n49968 );
xor ( n49970 , n49863 , n49867 );
xor ( n49971 , n49970 , n49870 );
and ( n49972 , n49968 , n49971 );
and ( n49973 , n49964 , n49971 );
or ( n49974 , n49969 , n49972 , n49973 );
and ( n49975 , n46777 , n40406 );
and ( n49976 , n46676 , n40404 );
nor ( n49977 , n49975 , n49976 );
xnor ( n49978 , n49977 , n40262 );
and ( n49979 , n49974 , n49978 );
xor ( n49980 , n49873 , n49877 );
xor ( n49981 , n49980 , n49880 );
and ( n49982 , n49978 , n49981 );
and ( n49983 , n49974 , n49981 );
or ( n49984 , n49979 , n49982 , n49983 );
and ( n49985 , n46676 , n40406 );
and ( n49986 , n46510 , n40404 );
nor ( n49987 , n49985 , n49986 );
xnor ( n49988 , n49987 , n40262 );
and ( n49989 , n49984 , n49988 );
xor ( n49990 , n49883 , n49887 );
xor ( n49991 , n49990 , n49890 );
and ( n49992 , n49988 , n49991 );
and ( n49993 , n49984 , n49991 );
or ( n49994 , n49989 , n49992 , n49993 );
and ( n49995 , n49899 , n49994 );
and ( n49996 , n46159 , n40666 );
and ( n49997 , n46069 , n40664 );
nor ( n49998 , n49996 , n49997 );
xnor ( n49999 , n49998 , n40445 );
buf ( n50000 , n30387 );
not ( n50001 , n50000 );
and ( n50002 , n49999 , n50001 );
xor ( n50003 , n49984 , n49988 );
xor ( n50004 , n50003 , n49991 );
and ( n50005 , n50001 , n50004 );
and ( n50006 , n49999 , n50004 );
or ( n50007 , n50002 , n50005 , n50006 );
and ( n50008 , n49994 , n50007 );
and ( n50009 , n49899 , n50007 );
or ( n50010 , n49995 , n50008 , n50009 );
and ( n50011 , n49896 , n50010 );
and ( n50012 , n49814 , n50010 );
or ( n50013 , n49897 , n50011 , n50012 );
and ( n50014 , n49811 , n50013 );
and ( n50015 , n49809 , n50013 );
or ( n50016 , n49812 , n50014 , n50015 );
and ( n50017 , n49743 , n50016 );
xor ( n50018 , n49809 , n49811 );
xor ( n50019 , n50018 , n50013 );
xor ( n50020 , n49814 , n49896 );
xor ( n50021 , n50020 , n50010 );
xor ( n50022 , n49903 , n49907 );
and ( n50023 , n48069 , n40664 );
not ( n50024 , n50023 );
and ( n50025 , n50024 , n40445 );
and ( n50026 , n48069 , n40666 );
and ( n50027 , n48077 , n40664 );
nor ( n50028 , n50026 , n50027 );
xnor ( n50029 , n50028 , n40445 );
and ( n50030 , n50025 , n50029 );
and ( n50031 , n48077 , n40666 );
and ( n50032 , n48086 , n40664 );
nor ( n50033 , n50031 , n50032 );
xnor ( n50034 , n50033 , n40445 );
and ( n50035 , n50030 , n50034 );
and ( n50036 , n50034 , n49901 );
and ( n50037 , n50030 , n49901 );
or ( n50038 , n50035 , n50036 , n50037 );
and ( n50039 , n50022 , n50038 );
and ( n50040 , n48086 , n40666 );
and ( n50041 , n48099 , n40664 );
nor ( n50042 , n50040 , n50041 );
xnor ( n50043 , n50042 , n40445 );
and ( n50044 , n50038 , n50043 );
and ( n50045 , n50022 , n50043 );
or ( n50046 , n50039 , n50044 , n50045 );
and ( n50047 , n48099 , n40666 );
and ( n50048 , n47927 , n40664 );
nor ( n50049 , n50047 , n50048 );
xnor ( n50050 , n50049 , n40445 );
and ( n50051 , n50046 , n50050 );
xor ( n50052 , n49908 , n49912 );
xor ( n50053 , n50052 , n49820 );
and ( n50054 , n50050 , n50053 );
and ( n50055 , n50046 , n50053 );
or ( n50056 , n50051 , n50054 , n50055 );
and ( n50057 , n47927 , n40666 );
and ( n50058 , n47932 , n40664 );
nor ( n50059 , n50057 , n50058 );
xnor ( n50060 , n50059 , n40445 );
and ( n50061 , n50056 , n50060 );
xor ( n50062 , n49900 , n49916 );
xor ( n50063 , n50062 , n49921 );
and ( n50064 , n50060 , n50063 );
and ( n50065 , n50056 , n50063 );
or ( n50066 , n50061 , n50064 , n50065 );
and ( n50067 , n47932 , n40666 );
and ( n50068 , n47645 , n40664 );
nor ( n50069 , n50067 , n50068 );
xnor ( n50070 , n50069 , n40445 );
and ( n50071 , n50066 , n50070 );
xor ( n50072 , n49924 , n49928 );
xor ( n50073 , n50072 , n49931 );
and ( n50074 , n50070 , n50073 );
and ( n50075 , n50066 , n50073 );
or ( n50076 , n50071 , n50074 , n50075 );
and ( n50077 , n47645 , n40666 );
and ( n50078 , n46948 , n40664 );
nor ( n50079 , n50077 , n50078 );
xnor ( n50080 , n50079 , n40445 );
and ( n50081 , n50076 , n50080 );
xor ( n50082 , n49934 , n49938 );
xor ( n50083 , n50082 , n49941 );
and ( n50084 , n50080 , n50083 );
and ( n50085 , n50076 , n50083 );
or ( n50086 , n50081 , n50084 , n50085 );
and ( n50087 , n46948 , n40666 );
and ( n50088 , n46777 , n40664 );
nor ( n50089 , n50087 , n50088 );
xnor ( n50090 , n50089 , n40445 );
and ( n50091 , n50086 , n50090 );
xor ( n50092 , n49944 , n49948 );
xor ( n50093 , n50092 , n49951 );
and ( n50094 , n50090 , n50093 );
and ( n50095 , n50086 , n50093 );
or ( n50096 , n50091 , n50094 , n50095 );
and ( n50097 , n46777 , n40666 );
and ( n50098 , n46676 , n40664 );
nor ( n50099 , n50097 , n50098 );
xnor ( n50100 , n50099 , n40445 );
and ( n50101 , n50096 , n50100 );
xor ( n50102 , n49954 , n49958 );
xor ( n50103 , n50102 , n49961 );
and ( n50104 , n50100 , n50103 );
and ( n50105 , n50096 , n50103 );
or ( n50106 , n50101 , n50104 , n50105 );
and ( n50107 , n46676 , n40666 );
and ( n50108 , n46510 , n40664 );
nor ( n50109 , n50107 , n50108 );
xnor ( n50110 , n50109 , n40445 );
and ( n50111 , n50106 , n50110 );
xor ( n50112 , n49964 , n49968 );
xor ( n50113 , n50112 , n49971 );
and ( n50114 , n50110 , n50113 );
and ( n50115 , n50106 , n50113 );
or ( n50116 , n50111 , n50114 , n50115 );
and ( n50117 , n46510 , n40666 );
and ( n50118 , n46159 , n40664 );
nor ( n50119 , n50117 , n50118 );
xnor ( n50120 , n50119 , n40445 );
and ( n50121 , n50116 , n50120 );
xor ( n50122 , n49974 , n49978 );
xor ( n50123 , n50122 , n49981 );
and ( n50124 , n50120 , n50123 );
and ( n50125 , n50116 , n50123 );
or ( n50126 , n50121 , n50124 , n50125 );
and ( n50127 , n46069 , n40928 );
and ( n50128 , n45754 , n40926 );
nor ( n50129 , n50127 , n50128 );
xnor ( n50130 , n50129 , n40688 );
buf ( n50131 , n30388 );
not ( n50132 , n50131 );
and ( n50133 , n50130 , n50132 );
xor ( n50134 , n50116 , n50120 );
xor ( n50135 , n50134 , n50123 );
and ( n50136 , n50132 , n50135 );
and ( n50137 , n50130 , n50135 );
or ( n50138 , n50133 , n50136 , n50137 );
and ( n50139 , n50126 , n50138 );
xor ( n50140 , n49999 , n50001 );
xor ( n50141 , n50140 , n50004 );
and ( n50142 , n50138 , n50141 );
and ( n50143 , n50126 , n50141 );
or ( n50144 , n50139 , n50142 , n50143 );
and ( n50145 , n44826 , n41230 );
and ( n50146 , n44347 , n41228 );
nor ( n50147 , n50145 , n50146 );
xnor ( n50148 , n50147 , n40981 );
and ( n50149 , n50144 , n50148 );
and ( n50150 , n50021 , n50149 );
and ( n50151 , n45057 , n41230 );
and ( n50152 , n44826 , n41228 );
nor ( n50153 , n50151 , n50152 );
xnor ( n50154 , n50153 , n40981 );
and ( n50155 , n45754 , n40928 );
and ( n50156 , n45171 , n40926 );
nor ( n50157 , n50155 , n50156 );
xnor ( n50158 , n50157 , n40688 );
and ( n50159 , n50154 , n50158 );
xor ( n50160 , n50126 , n50138 );
xor ( n50161 , n50160 , n50141 );
and ( n50162 , n50158 , n50161 );
and ( n50163 , n50154 , n50161 );
or ( n50164 , n50159 , n50162 , n50163 );
and ( n50165 , n43820 , n41981 );
and ( n50166 , n43679 , n41979 );
nor ( n50167 , n50165 , n50166 );
xnor ( n50168 , n50167 , n41373 );
and ( n50169 , n50164 , n50168 );
and ( n50170 , n44318 , n41522 );
and ( n50171 , n44000 , n41520 );
nor ( n50172 , n50170 , n50171 );
xnor ( n50173 , n50172 , n41100 );
and ( n50174 , n50168 , n50173 );
and ( n50175 , n50164 , n50173 );
or ( n50176 , n50169 , n50174 , n50175 );
and ( n50177 , n50149 , n50176 );
and ( n50178 , n50021 , n50176 );
or ( n50179 , n50150 , n50177 , n50178 );
and ( n50180 , n50019 , n50179 );
xor ( n50181 , n49899 , n49994 );
xor ( n50182 , n50181 , n50007 );
xor ( n50183 , n50144 , n50148 );
and ( n50184 , n50182 , n50183 );
and ( n50185 , n43679 , n42079 );
and ( n50186 , n43671 , n42076 );
nor ( n50187 , n50185 , n50186 );
xnor ( n50188 , n50187 , n41370 );
and ( n50189 , n44000 , n41981 );
and ( n50190 , n43820 , n41979 );
nor ( n50191 , n50189 , n50190 );
xnor ( n50192 , n50191 , n41373 );
and ( n50193 , n50188 , n50192 );
and ( n50194 , n44318 , n41981 );
and ( n50195 , n44000 , n41979 );
nor ( n50196 , n50194 , n50195 );
xnor ( n50197 , n50196 , n41373 );
and ( n50198 , n44000 , n42079 );
and ( n50199 , n43820 , n42076 );
nor ( n50200 , n50198 , n50199 );
xnor ( n50201 , n50200 , n41370 );
and ( n50202 , n44347 , n41981 );
and ( n50203 , n44318 , n41979 );
nor ( n50204 , n50202 , n50203 );
xnor ( n50205 , n50204 , n41373 );
and ( n50206 , n50201 , n50205 );
and ( n50207 , n45057 , n41522 );
and ( n50208 , n44826 , n41520 );
nor ( n50209 , n50207 , n50208 );
xnor ( n50210 , n50209 , n41100 );
and ( n50211 , n50205 , n50210 );
and ( n50212 , n50201 , n50210 );
or ( n50213 , n50206 , n50211 , n50212 );
and ( n50214 , n50197 , n50213 );
xor ( n50215 , n50025 , n50029 );
and ( n50216 , n48069 , n40926 );
not ( n50217 , n50216 );
and ( n50218 , n50217 , n40688 );
and ( n50219 , n48069 , n40928 );
and ( n50220 , n48077 , n40926 );
nor ( n50221 , n50219 , n50220 );
xnor ( n50222 , n50221 , n40688 );
and ( n50223 , n50218 , n50222 );
and ( n50224 , n48077 , n40928 );
and ( n50225 , n48086 , n40926 );
nor ( n50226 , n50224 , n50225 );
xnor ( n50227 , n50226 , n40688 );
and ( n50228 , n50223 , n50227 );
and ( n50229 , n50227 , n50023 );
and ( n50230 , n50223 , n50023 );
or ( n50231 , n50228 , n50229 , n50230 );
and ( n50232 , n50215 , n50231 );
and ( n50233 , n48086 , n40928 );
and ( n50234 , n48099 , n40926 );
nor ( n50235 , n50233 , n50234 );
xnor ( n50236 , n50235 , n40688 );
and ( n50237 , n50231 , n50236 );
and ( n50238 , n50215 , n50236 );
or ( n50239 , n50232 , n50237 , n50238 );
and ( n50240 , n48099 , n40928 );
and ( n50241 , n47927 , n40926 );
nor ( n50242 , n50240 , n50241 );
xnor ( n50243 , n50242 , n40688 );
and ( n50244 , n50239 , n50243 );
xor ( n50245 , n50030 , n50034 );
xor ( n50246 , n50245 , n49901 );
and ( n50247 , n50243 , n50246 );
and ( n50248 , n50239 , n50246 );
or ( n50249 , n50244 , n50247 , n50248 );
and ( n50250 , n47927 , n40928 );
and ( n50251 , n47932 , n40926 );
nor ( n50252 , n50250 , n50251 );
xnor ( n50253 , n50252 , n40688 );
and ( n50254 , n50249 , n50253 );
xor ( n50255 , n50022 , n50038 );
xor ( n50256 , n50255 , n50043 );
and ( n50257 , n50253 , n50256 );
and ( n50258 , n50249 , n50256 );
or ( n50259 , n50254 , n50257 , n50258 );
and ( n50260 , n47932 , n40928 );
and ( n50261 , n47645 , n40926 );
nor ( n50262 , n50260 , n50261 );
xnor ( n50263 , n50262 , n40688 );
and ( n50264 , n50259 , n50263 );
xor ( n50265 , n50046 , n50050 );
xor ( n50266 , n50265 , n50053 );
and ( n50267 , n50263 , n50266 );
and ( n50268 , n50259 , n50266 );
or ( n50269 , n50264 , n50267 , n50268 );
and ( n50270 , n47645 , n40928 );
and ( n50271 , n46948 , n40926 );
nor ( n50272 , n50270 , n50271 );
xnor ( n50273 , n50272 , n40688 );
and ( n50274 , n50269 , n50273 );
xor ( n50275 , n50056 , n50060 );
xor ( n50276 , n50275 , n50063 );
and ( n50277 , n50273 , n50276 );
and ( n50278 , n50269 , n50276 );
or ( n50279 , n50274 , n50277 , n50278 );
and ( n50280 , n46948 , n40928 );
and ( n50281 , n46777 , n40926 );
nor ( n50282 , n50280 , n50281 );
xnor ( n50283 , n50282 , n40688 );
and ( n50284 , n50279 , n50283 );
xor ( n50285 , n50066 , n50070 );
xor ( n50286 , n50285 , n50073 );
and ( n50287 , n50283 , n50286 );
and ( n50288 , n50279 , n50286 );
or ( n50289 , n50284 , n50287 , n50288 );
and ( n50290 , n46777 , n40928 );
and ( n50291 , n46676 , n40926 );
nor ( n50292 , n50290 , n50291 );
xnor ( n50293 , n50292 , n40688 );
and ( n50294 , n50289 , n50293 );
xor ( n50295 , n50076 , n50080 );
xor ( n50296 , n50295 , n50083 );
and ( n50297 , n50293 , n50296 );
and ( n50298 , n50289 , n50296 );
or ( n50299 , n50294 , n50297 , n50298 );
and ( n50300 , n46676 , n40928 );
and ( n50301 , n46510 , n40926 );
nor ( n50302 , n50300 , n50301 );
xnor ( n50303 , n50302 , n40688 );
and ( n50304 , n50299 , n50303 );
xor ( n50305 , n50086 , n50090 );
xor ( n50306 , n50305 , n50093 );
and ( n50307 , n50303 , n50306 );
and ( n50308 , n50299 , n50306 );
or ( n50309 , n50304 , n50307 , n50308 );
and ( n50310 , n46069 , n41230 );
and ( n50311 , n45754 , n41228 );
nor ( n50312 , n50310 , n50311 );
xnor ( n50313 , n50312 , n40981 );
and ( n50314 , n50309 , n50313 );
and ( n50315 , n46510 , n40928 );
and ( n50316 , n46159 , n40926 );
nor ( n50317 , n50315 , n50316 );
xnor ( n50318 , n50317 , n40688 );
buf ( n50319 , n30390 );
not ( n50320 , n50319 );
xor ( n50321 , n50318 , n50320 );
xor ( n50322 , n50096 , n50100 );
xor ( n50323 , n50322 , n50103 );
xor ( n50324 , n50321 , n50323 );
and ( n50325 , n50313 , n50324 );
and ( n50326 , n50309 , n50324 );
or ( n50327 , n50314 , n50325 , n50326 );
and ( n50328 , n46159 , n40928 );
and ( n50329 , n46069 , n40926 );
nor ( n50330 , n50328 , n50329 );
xnor ( n50331 , n50330 , n40688 );
and ( n50332 , n50327 , n50331 );
and ( n50333 , n50318 , n50320 );
and ( n50334 , n50320 , n50323 );
and ( n50335 , n50318 , n50323 );
or ( n50336 , n50333 , n50334 , n50335 );
buf ( n50337 , n30389 );
not ( n50338 , n50337 );
xor ( n50339 , n50336 , n50338 );
xor ( n50340 , n50106 , n50110 );
xor ( n50341 , n50340 , n50113 );
xor ( n50342 , n50339 , n50341 );
and ( n50343 , n50331 , n50342 );
and ( n50344 , n50327 , n50342 );
or ( n50345 , n50332 , n50343 , n50344 );
and ( n50346 , n50213 , n50345 );
and ( n50347 , n50197 , n50345 );
or ( n50348 , n50214 , n50346 , n50347 );
and ( n50349 , n50192 , n50348 );
and ( n50350 , n50188 , n50348 );
or ( n50351 , n50193 , n50349 , n50350 );
and ( n50352 , n50183 , n50351 );
and ( n50353 , n50182 , n50351 );
or ( n50354 , n50184 , n50352 , n50353 );
xor ( n50355 , n50164 , n50168 );
xor ( n50356 , n50355 , n50173 );
and ( n50357 , n50336 , n50338 );
and ( n50358 , n50338 , n50341 );
and ( n50359 , n50336 , n50341 );
or ( n50360 , n50357 , n50358 , n50359 );
and ( n50361 , n45171 , n41230 );
and ( n50362 , n45057 , n41228 );
nor ( n50363 , n50361 , n50362 );
xnor ( n50364 , n50363 , n40981 );
and ( n50365 , n50360 , n50364 );
xor ( n50366 , n50130 , n50132 );
xor ( n50367 , n50366 , n50135 );
and ( n50368 , n50364 , n50367 );
and ( n50369 , n50360 , n50367 );
or ( n50370 , n50365 , n50368 , n50369 );
and ( n50371 , n44347 , n41522 );
and ( n50372 , n44318 , n41520 );
nor ( n50373 , n50371 , n50372 );
xnor ( n50374 , n50373 , n41100 );
and ( n50375 , n50370 , n50374 );
xor ( n50376 , n50154 , n50158 );
xor ( n50377 , n50376 , n50161 );
and ( n50378 , n50374 , n50377 );
and ( n50379 , n50370 , n50377 );
or ( n50380 , n50375 , n50378 , n50379 );
and ( n50381 , n50356 , n50380 );
xor ( n50382 , n50182 , n50183 );
xor ( n50383 , n50382 , n50351 );
and ( n50384 , n50380 , n50383 );
and ( n50385 , n50356 , n50383 );
or ( n50386 , n50381 , n50384 , n50385 );
and ( n50387 , n50354 , n50386 );
xor ( n50388 , n50021 , n50149 );
xor ( n50389 , n50388 , n50176 );
and ( n50390 , n50386 , n50389 );
and ( n50391 , n50354 , n50389 );
or ( n50392 , n50387 , n50390 , n50391 );
and ( n50393 , n50179 , n50392 );
and ( n50394 , n50019 , n50392 );
or ( n50395 , n50180 , n50393 , n50394 );
and ( n50396 , n50016 , n50395 );
and ( n50397 , n49743 , n50395 );
or ( n50398 , n50017 , n50396 , n50397 );
and ( n50399 , n49740 , n50398 );
and ( n50400 , n49738 , n50398 );
or ( n50401 , n49741 , n50399 , n50400 );
and ( n50402 , n49735 , n50401 );
and ( n50403 , n49733 , n50401 );
or ( n50404 , n49736 , n50402 , n50403 );
and ( n50405 , n49667 , n50404 );
xor ( n50406 , n49667 , n50404 );
xor ( n50407 , n49733 , n49735 );
xor ( n50408 , n50407 , n50401 );
xor ( n50409 , n49738 , n49740 );
xor ( n50410 , n50409 , n50398 );
xor ( n50411 , n49743 , n50016 );
xor ( n50412 , n50411 , n50395 );
xor ( n50413 , n50019 , n50179 );
xor ( n50414 , n50413 , n50392 );
xor ( n50415 , n50354 , n50386 );
xor ( n50416 , n50415 , n50389 );
and ( n50417 , n46159 , n41230 );
and ( n50418 , n46069 , n41228 );
nor ( n50419 , n50417 , n50418 );
xnor ( n50420 , n50419 , n40981 );
buf ( n50421 , n30391 );
not ( n50422 , n50421 );
and ( n50423 , n50420 , n50422 );
xor ( n50424 , n50299 , n50303 );
xor ( n50425 , n50424 , n50306 );
and ( n50426 , n50422 , n50425 );
and ( n50427 , n50420 , n50425 );
or ( n50428 , n50423 , n50426 , n50427 );
and ( n50429 , n45171 , n41522 );
and ( n50430 , n45057 , n41520 );
nor ( n50431 , n50429 , n50430 );
xnor ( n50432 , n50431 , n41100 );
and ( n50433 , n50428 , n50432 );
xor ( n50434 , n50309 , n50313 );
xor ( n50435 , n50434 , n50324 );
and ( n50436 , n50432 , n50435 );
and ( n50437 , n50428 , n50435 );
or ( n50438 , n50433 , n50436 , n50437 );
and ( n50439 , n45754 , n41230 );
and ( n50440 , n45171 , n41228 );
nor ( n50441 , n50439 , n50440 );
xnor ( n50442 , n50441 , n40981 );
and ( n50443 , n50438 , n50442 );
xor ( n50444 , n50327 , n50331 );
xor ( n50445 , n50444 , n50342 );
and ( n50446 , n50442 , n50445 );
and ( n50447 , n50438 , n50445 );
or ( n50448 , n50443 , n50446 , n50447 );
and ( n50449 , n43820 , n42079 );
and ( n50450 , n43679 , n42076 );
nor ( n50451 , n50449 , n50450 );
xnor ( n50452 , n50451 , n41370 );
and ( n50453 , n50448 , n50452 );
and ( n50454 , n44826 , n41522 );
and ( n50455 , n44347 , n41520 );
nor ( n50456 , n50454 , n50455 );
xnor ( n50457 , n50456 , n41100 );
and ( n50458 , n50452 , n50457 );
and ( n50459 , n50448 , n50457 );
or ( n50460 , n50453 , n50458 , n50459 );
xor ( n50461 , n50370 , n50374 );
xor ( n50462 , n50461 , n50377 );
or ( n50463 , n50460 , n50462 );
xor ( n50464 , n50356 , n50380 );
xor ( n50465 , n50464 , n50383 );
and ( n50466 , n50463 , n50465 );
xor ( n50467 , n50188 , n50192 );
xor ( n50468 , n50467 , n50348 );
xor ( n50469 , n50360 , n50364 );
xor ( n50470 , n50469 , n50367 );
xor ( n50471 , n50197 , n50213 );
xor ( n50472 , n50471 , n50345 );
and ( n50473 , n50470 , n50472 );
xor ( n50474 , n50448 , n50452 );
xor ( n50475 , n50474 , n50457 );
and ( n50476 , n50472 , n50475 );
and ( n50477 , n50470 , n50475 );
or ( n50478 , n50473 , n50476 , n50477 );
and ( n50479 , n50468 , n50478 );
xnor ( n50480 , n50460 , n50462 );
and ( n50481 , n50478 , n50480 );
and ( n50482 , n50468 , n50480 );
or ( n50483 , n50479 , n50481 , n50482 );
and ( n50484 , n50465 , n50483 );
and ( n50485 , n50463 , n50483 );
or ( n50486 , n50466 , n50484 , n50485 );
and ( n50487 , n50416 , n50486 );
xor ( n50488 , n50463 , n50465 );
xor ( n50489 , n50488 , n50483 );
xor ( n50490 , n50468 , n50478 );
xor ( n50491 , n50490 , n50480 );
and ( n50492 , n46510 , n41230 );
and ( n50493 , n46159 , n41228 );
nor ( n50494 , n50492 , n50493 );
xnor ( n50495 , n50494 , n40981 );
buf ( n50496 , n30392 );
not ( n50497 , n50496 );
and ( n50498 , n50495 , n50497 );
xor ( n50499 , n50289 , n50293 );
xor ( n50500 , n50499 , n50296 );
and ( n50501 , n50497 , n50500 );
and ( n50502 , n50495 , n50500 );
or ( n50503 , n50498 , n50501 , n50502 );
and ( n50504 , n46777 , n41230 );
and ( n50505 , n46676 , n41228 );
nor ( n50506 , n50504 , n50505 );
xnor ( n50507 , n50506 , n40981 );
buf ( n50508 , n30394 );
not ( n50509 , n50508 );
and ( n50510 , n50507 , n50509 );
xor ( n50511 , n50269 , n50273 );
xor ( n50512 , n50511 , n50276 );
and ( n50513 , n50509 , n50512 );
and ( n50514 , n50507 , n50512 );
or ( n50515 , n50510 , n50513 , n50514 );
and ( n50516 , n46676 , n41230 );
and ( n50517 , n46510 , n41228 );
nor ( n50518 , n50516 , n50517 );
xnor ( n50519 , n50518 , n40981 );
and ( n50520 , n50515 , n50519 );
xor ( n50521 , n50279 , n50283 );
xor ( n50522 , n50521 , n50286 );
and ( n50523 , n50519 , n50522 );
and ( n50524 , n50515 , n50522 );
or ( n50525 , n50520 , n50523 , n50524 );
and ( n50526 , n46069 , n41522 );
and ( n50527 , n45754 , n41520 );
nor ( n50528 , n50526 , n50527 );
xnor ( n50529 , n50528 , n41100 );
and ( n50530 , n50525 , n50529 );
xor ( n50531 , n50495 , n50497 );
xor ( n50532 , n50531 , n50500 );
and ( n50533 , n50529 , n50532 );
and ( n50534 , n50525 , n50532 );
or ( n50535 , n50530 , n50533 , n50534 );
and ( n50536 , n50503 , n50535 );
xor ( n50537 , n50420 , n50422 );
xor ( n50538 , n50537 , n50425 );
and ( n50539 , n50535 , n50538 );
and ( n50540 , n50503 , n50538 );
or ( n50541 , n50536 , n50539 , n50540 );
and ( n50542 , n44826 , n41981 );
and ( n50543 , n44347 , n41979 );
nor ( n50544 , n50542 , n50543 );
xnor ( n50545 , n50544 , n41373 );
and ( n50546 , n50541 , n50545 );
xor ( n50547 , n50428 , n50432 );
xor ( n50548 , n50547 , n50435 );
and ( n50549 , n50545 , n50548 );
and ( n50550 , n50541 , n50548 );
or ( n50551 , n50546 , n50549 , n50550 );
xor ( n50552 , n50201 , n50205 );
xor ( n50553 , n50552 , n50210 );
and ( n50554 , n50551 , n50553 );
xor ( n50555 , n50438 , n50442 );
xor ( n50556 , n50555 , n50445 );
and ( n50557 , n50553 , n50556 );
and ( n50558 , n50551 , n50556 );
or ( n50559 , n50554 , n50557 , n50558 );
xor ( n50560 , n50470 , n50472 );
xor ( n50561 , n50560 , n50475 );
and ( n50562 , n50559 , n50561 );
xor ( n50563 , n50551 , n50553 );
xor ( n50564 , n50563 , n50556 );
and ( n50565 , n45057 , n41981 );
and ( n50566 , n44826 , n41979 );
nor ( n50567 , n50565 , n50566 );
xnor ( n50568 , n50567 , n41373 );
and ( n50569 , n45754 , n41522 );
and ( n50570 , n45171 , n41520 );
nor ( n50571 , n50569 , n50570 );
xnor ( n50572 , n50571 , n41100 );
and ( n50573 , n50568 , n50572 );
xor ( n50574 , n50503 , n50535 );
xor ( n50575 , n50574 , n50538 );
and ( n50576 , n50572 , n50575 );
and ( n50577 , n50568 , n50575 );
or ( n50578 , n50573 , n50576 , n50577 );
and ( n50579 , n44318 , n42079 );
and ( n50580 , n44000 , n42076 );
nor ( n50581 , n50579 , n50580 );
xnor ( n50582 , n50581 , n41370 );
and ( n50583 , n50578 , n50582 );
xor ( n50584 , n50541 , n50545 );
xor ( n50585 , n50584 , n50548 );
and ( n50586 , n50582 , n50585 );
and ( n50587 , n50578 , n50585 );
or ( n50588 , n50583 , n50586 , n50587 );
and ( n50589 , n50564 , n50588 );
xor ( n50590 , n50578 , n50582 );
xor ( n50591 , n50590 , n50585 );
xor ( n50592 , n50218 , n50222 );
and ( n50593 , n48069 , n41228 );
not ( n50594 , n50593 );
and ( n50595 , n50594 , n40981 );
and ( n50596 , n48069 , n41230 );
and ( n50597 , n48077 , n41228 );
nor ( n50598 , n50596 , n50597 );
xnor ( n50599 , n50598 , n40981 );
and ( n50600 , n50595 , n50599 );
and ( n50601 , n48077 , n41230 );
and ( n50602 , n48086 , n41228 );
nor ( n50603 , n50601 , n50602 );
xnor ( n50604 , n50603 , n40981 );
and ( n50605 , n50600 , n50604 );
and ( n50606 , n50604 , n50216 );
and ( n50607 , n50600 , n50216 );
or ( n50608 , n50605 , n50606 , n50607 );
and ( n50609 , n50592 , n50608 );
and ( n50610 , n48086 , n41230 );
and ( n50611 , n48099 , n41228 );
nor ( n50612 , n50610 , n50611 );
xnor ( n50613 , n50612 , n40981 );
and ( n50614 , n50608 , n50613 );
and ( n50615 , n50592 , n50613 );
or ( n50616 , n50609 , n50614 , n50615 );
and ( n50617 , n48099 , n41230 );
and ( n50618 , n47927 , n41228 );
nor ( n50619 , n50617 , n50618 );
xnor ( n50620 , n50619 , n40981 );
and ( n50621 , n50616 , n50620 );
xor ( n50622 , n50223 , n50227 );
xor ( n50623 , n50622 , n50023 );
and ( n50624 , n50620 , n50623 );
and ( n50625 , n50616 , n50623 );
or ( n50626 , n50621 , n50624 , n50625 );
and ( n50627 , n47927 , n41230 );
and ( n50628 , n47932 , n41228 );
nor ( n50629 , n50627 , n50628 );
xnor ( n50630 , n50629 , n40981 );
and ( n50631 , n50626 , n50630 );
xor ( n50632 , n50215 , n50231 );
xor ( n50633 , n50632 , n50236 );
and ( n50634 , n50630 , n50633 );
and ( n50635 , n50626 , n50633 );
or ( n50636 , n50631 , n50634 , n50635 );
and ( n50637 , n47932 , n41230 );
and ( n50638 , n47645 , n41228 );
nor ( n50639 , n50637 , n50638 );
xnor ( n50640 , n50639 , n40981 );
and ( n50641 , n50636 , n50640 );
xor ( n50642 , n50239 , n50243 );
xor ( n50643 , n50642 , n50246 );
and ( n50644 , n50640 , n50643 );
and ( n50645 , n50636 , n50643 );
or ( n50646 , n50641 , n50644 , n50645 );
and ( n50647 , n47645 , n41230 );
and ( n50648 , n46948 , n41228 );
nor ( n50649 , n50647 , n50648 );
xnor ( n50650 , n50649 , n40981 );
and ( n50651 , n50646 , n50650 );
xor ( n50652 , n50249 , n50253 );
xor ( n50653 , n50652 , n50256 );
and ( n50654 , n50650 , n50653 );
and ( n50655 , n50646 , n50653 );
or ( n50656 , n50651 , n50654 , n50655 );
and ( n50657 , n46948 , n41230 );
and ( n50658 , n46777 , n41228 );
nor ( n50659 , n50657 , n50658 );
xnor ( n50660 , n50659 , n40981 );
and ( n50661 , n50656 , n50660 );
xor ( n50662 , n50259 , n50263 );
xor ( n50663 , n50662 , n50266 );
and ( n50664 , n50660 , n50663 );
and ( n50665 , n50656 , n50663 );
or ( n50666 , n50661 , n50664 , n50665 );
and ( n50667 , n46676 , n41522 );
and ( n50668 , n46510 , n41520 );
nor ( n50669 , n50667 , n50668 );
xnor ( n50670 , n50669 , n41100 );
buf ( n50671 , n30395 );
not ( n50672 , n50671 );
and ( n50673 , n50670 , n50672 );
xor ( n50674 , n50656 , n50660 );
xor ( n50675 , n50674 , n50663 );
and ( n50676 , n50672 , n50675 );
and ( n50677 , n50670 , n50675 );
or ( n50678 , n50673 , n50676 , n50677 );
and ( n50679 , n50666 , n50678 );
xor ( n50680 , n50507 , n50509 );
xor ( n50681 , n50680 , n50512 );
and ( n50682 , n50678 , n50681 );
and ( n50683 , n50666 , n50681 );
or ( n50684 , n50679 , n50682 , n50683 );
buf ( n50685 , n30393 );
not ( n50686 , n50685 );
and ( n50687 , n50684 , n50686 );
xor ( n50688 , n50515 , n50519 );
xor ( n50689 , n50688 , n50522 );
and ( n50690 , n50686 , n50689 );
and ( n50691 , n50684 , n50689 );
or ( n50692 , n50687 , n50690 , n50691 );
and ( n50693 , n46069 , n41981 );
and ( n50694 , n45754 , n41979 );
nor ( n50695 , n50693 , n50694 );
xnor ( n50696 , n50695 , n41373 );
and ( n50697 , n46510 , n41522 );
and ( n50698 , n46159 , n41520 );
nor ( n50699 , n50697 , n50698 );
xnor ( n50700 , n50699 , n41100 );
and ( n50701 , n50696 , n50700 );
xor ( n50702 , n50666 , n50678 );
xor ( n50703 , n50702 , n50681 );
and ( n50704 , n50700 , n50703 );
and ( n50705 , n50696 , n50703 );
or ( n50706 , n50701 , n50704 , n50705 );
and ( n50707 , n46159 , n41522 );
and ( n50708 , n46069 , n41520 );
nor ( n50709 , n50707 , n50708 );
xnor ( n50710 , n50709 , n41100 );
and ( n50711 , n50706 , n50710 );
xor ( n50712 , n50684 , n50686 );
xor ( n50713 , n50712 , n50689 );
and ( n50714 , n50710 , n50713 );
and ( n50715 , n50706 , n50713 );
or ( n50716 , n50711 , n50714 , n50715 );
and ( n50717 , n50692 , n50716 );
xor ( n50718 , n50525 , n50529 );
xor ( n50719 , n50718 , n50532 );
and ( n50720 , n50716 , n50719 );
and ( n50721 , n50692 , n50719 );
or ( n50722 , n50717 , n50720 , n50721 );
and ( n50723 , n44347 , n42079 );
and ( n50724 , n44318 , n42076 );
nor ( n50725 , n50723 , n50724 );
xnor ( n50726 , n50725 , n41370 );
and ( n50727 , n50722 , n50726 );
xor ( n50728 , n50568 , n50572 );
xor ( n50729 , n50728 , n50575 );
and ( n50730 , n50726 , n50729 );
and ( n50731 , n50722 , n50729 );
or ( n50732 , n50727 , n50730 , n50731 );
and ( n50733 , n50591 , n50732 );
xor ( n50734 , n50722 , n50726 );
xor ( n50735 , n50734 , n50729 );
and ( n50736 , n46777 , n41522 );
and ( n50737 , n46676 , n41520 );
nor ( n50738 , n50736 , n50737 );
xnor ( n50739 , n50738 , n41100 );
buf ( n50740 , n30396 );
not ( n50741 , n50740 );
and ( n50742 , n50739 , n50741 );
xor ( n50743 , n50646 , n50650 );
xor ( n50744 , n50743 , n50653 );
and ( n50745 , n50741 , n50744 );
and ( n50746 , n50739 , n50744 );
or ( n50747 , n50742 , n50745 , n50746 );
xor ( n50748 , n50595 , n50599 );
and ( n50749 , n48069 , n41520 );
not ( n50750 , n50749 );
and ( n50751 , n50750 , n41100 );
and ( n50752 , n48069 , n41522 );
and ( n50753 , n48077 , n41520 );
nor ( n50754 , n50752 , n50753 );
xnor ( n50755 , n50754 , n41100 );
and ( n50756 , n50751 , n50755 );
and ( n50757 , n48077 , n41522 );
and ( n50758 , n48086 , n41520 );
nor ( n50759 , n50757 , n50758 );
xnor ( n50760 , n50759 , n41100 );
and ( n50761 , n50756 , n50760 );
and ( n50762 , n50760 , n50593 );
and ( n50763 , n50756 , n50593 );
or ( n50764 , n50761 , n50762 , n50763 );
and ( n50765 , n50748 , n50764 );
and ( n50766 , n48086 , n41522 );
and ( n50767 , n48099 , n41520 );
nor ( n50768 , n50766 , n50767 );
xnor ( n50769 , n50768 , n41100 );
and ( n50770 , n50764 , n50769 );
and ( n50771 , n50748 , n50769 );
or ( n50772 , n50765 , n50770 , n50771 );
and ( n50773 , n48099 , n41522 );
and ( n50774 , n47927 , n41520 );
nor ( n50775 , n50773 , n50774 );
xnor ( n50776 , n50775 , n41100 );
and ( n50777 , n50772 , n50776 );
xor ( n50778 , n50600 , n50604 );
xor ( n50779 , n50778 , n50216 );
and ( n50780 , n50776 , n50779 );
and ( n50781 , n50772 , n50779 );
or ( n50782 , n50777 , n50780 , n50781 );
and ( n50783 , n47927 , n41522 );
and ( n50784 , n47932 , n41520 );
nor ( n50785 , n50783 , n50784 );
xnor ( n50786 , n50785 , n41100 );
and ( n50787 , n50782 , n50786 );
xor ( n50788 , n50592 , n50608 );
xor ( n50789 , n50788 , n50613 );
and ( n50790 , n50786 , n50789 );
and ( n50791 , n50782 , n50789 );
or ( n50792 , n50787 , n50790 , n50791 );
and ( n50793 , n47932 , n41522 );
and ( n50794 , n47645 , n41520 );
nor ( n50795 , n50793 , n50794 );
xnor ( n50796 , n50795 , n41100 );
and ( n50797 , n50792 , n50796 );
xor ( n50798 , n50616 , n50620 );
xor ( n50799 , n50798 , n50623 );
and ( n50800 , n50796 , n50799 );
and ( n50801 , n50792 , n50799 );
or ( n50802 , n50797 , n50800 , n50801 );
buf ( n50803 , n30398 );
not ( n50804 , n50803 );
and ( n50805 , n50802 , n50804 );
xor ( n50806 , n50626 , n50630 );
xor ( n50807 , n50806 , n50633 );
and ( n50808 , n50804 , n50807 );
and ( n50809 , n50802 , n50807 );
or ( n50810 , n50805 , n50808 , n50809 );
buf ( n50811 , n30397 );
not ( n50812 , n50811 );
and ( n50813 , n50810 , n50812 );
xor ( n50814 , n50636 , n50640 );
xor ( n50815 , n50814 , n50643 );
and ( n50816 , n50812 , n50815 );
and ( n50817 , n50810 , n50815 );
or ( n50818 , n50813 , n50816 , n50817 );
xor ( n50819 , n50751 , n50755 );
and ( n50820 , n48069 , n41979 );
not ( n50821 , n50820 );
and ( n50822 , n50821 , n41373 );
and ( n50823 , n48069 , n41981 );
and ( n50824 , n48077 , n41979 );
nor ( n50825 , n50823 , n50824 );
xnor ( n50826 , n50825 , n41373 );
and ( n50827 , n50822 , n50826 );
and ( n50828 , n50827 , n50749 );
buf ( n50829 , n30405 );
not ( n50830 , n50829 );
and ( n50831 , n50749 , n50830 );
and ( n50832 , n50827 , n50830 );
or ( n50833 , n50828 , n50831 , n50832 );
and ( n50834 , n50819 , n50833 );
buf ( n50835 , n30404 );
not ( n50836 , n50835 );
and ( n50837 , n50833 , n50836 );
and ( n50838 , n50819 , n50836 );
or ( n50839 , n50834 , n50837 , n50838 );
buf ( n50840 , n30403 );
not ( n50841 , n50840 );
and ( n50842 , n50839 , n50841 );
xor ( n50843 , n50756 , n50760 );
xor ( n50844 , n50843 , n50593 );
and ( n50845 , n50841 , n50844 );
and ( n50846 , n50839 , n50844 );
or ( n50847 , n50842 , n50845 , n50846 );
buf ( n50848 , n30402 );
not ( n50849 , n50848 );
and ( n50850 , n50847 , n50849 );
xor ( n50851 , n50748 , n50764 );
xor ( n50852 , n50851 , n50769 );
and ( n50853 , n50849 , n50852 );
and ( n50854 , n50847 , n50852 );
or ( n50855 , n50850 , n50853 , n50854 );
buf ( n50856 , n30401 );
not ( n50857 , n50856 );
and ( n50858 , n50855 , n50857 );
xor ( n50859 , n50772 , n50776 );
xor ( n50860 , n50859 , n50779 );
and ( n50861 , n50857 , n50860 );
and ( n50862 , n50855 , n50860 );
or ( n50863 , n50858 , n50861 , n50862 );
buf ( n50864 , n30400 );
not ( n50865 , n50864 );
and ( n50866 , n50863 , n50865 );
xor ( n50867 , n50782 , n50786 );
xor ( n50868 , n50867 , n50789 );
and ( n50869 , n50865 , n50868 );
and ( n50870 , n50863 , n50868 );
or ( n50871 , n50866 , n50869 , n50870 );
buf ( n50872 , n30399 );
not ( n50873 , n50872 );
and ( n50874 , n50871 , n50873 );
xor ( n50875 , n50792 , n50796 );
xor ( n50876 , n50875 , n50799 );
and ( n50877 , n50873 , n50876 );
and ( n50878 , n50871 , n50876 );
or ( n50879 , n50874 , n50877 , n50878 );
and ( n50880 , n47645 , n41522 );
and ( n50881 , n46948 , n41520 );
nor ( n50882 , n50880 , n50881 );
xnor ( n50883 , n50882 , n41100 );
and ( n50884 , n50879 , n50883 );
xor ( n50885 , n50802 , n50804 );
xor ( n50886 , n50885 , n50807 );
and ( n50887 , n50883 , n50886 );
and ( n50888 , n50879 , n50886 );
or ( n50889 , n50884 , n50887 , n50888 );
and ( n50890 , n46948 , n41522 );
and ( n50891 , n46777 , n41520 );
nor ( n50892 , n50890 , n50891 );
xnor ( n50893 , n50892 , n41100 );
and ( n50894 , n50889 , n50893 );
xor ( n50895 , n50810 , n50812 );
xor ( n50896 , n50895 , n50815 );
and ( n50897 , n50893 , n50896 );
and ( n50898 , n50889 , n50896 );
or ( n50899 , n50894 , n50897 , n50898 );
and ( n50900 , n50818 , n50899 );
xor ( n50901 , n50739 , n50741 );
xor ( n50902 , n50901 , n50744 );
and ( n50903 , n50899 , n50902 );
and ( n50904 , n50818 , n50902 );
or ( n50905 , n50900 , n50903 , n50904 );
and ( n50906 , n50747 , n50905 );
xor ( n50907 , n50670 , n50672 );
xor ( n50908 , n50907 , n50675 );
and ( n50909 , n50905 , n50908 );
and ( n50910 , n50747 , n50908 );
or ( n50911 , n50906 , n50909 , n50910 );
xor ( n50912 , n50822 , n50826 );
and ( n50913 , n48069 , n42076 );
not ( n50914 , n50913 );
and ( n50915 , n50914 , n41370 );
buf ( n50916 , n30408 );
not ( n50917 , n50916 );
and ( n50918 , n50915 , n50917 );
and ( n50919 , n50918 , n50820 );
buf ( n50920 , n30407 );
not ( n50921 , n50920 );
and ( n50922 , n50820 , n50921 );
and ( n50923 , n50918 , n50921 );
or ( n50924 , n50919 , n50922 , n50923 );
and ( n50925 , n50912 , n50924 );
buf ( n50926 , n30406 );
not ( n50927 , n50926 );
and ( n50928 , n50924 , n50927 );
and ( n50929 , n50912 , n50927 );
or ( n50930 , n50925 , n50928 , n50929 );
and ( n50931 , n48077 , n41981 );
and ( n50932 , n48086 , n41979 );
nor ( n50933 , n50931 , n50932 );
xnor ( n50934 , n50933 , n41373 );
and ( n50935 , n50930 , n50934 );
xor ( n50936 , n50827 , n50749 );
xor ( n50937 , n50936 , n50830 );
and ( n50938 , n50934 , n50937 );
and ( n50939 , n50930 , n50937 );
or ( n50940 , n50935 , n50938 , n50939 );
and ( n50941 , n48086 , n41981 );
and ( n50942 , n48099 , n41979 );
nor ( n50943 , n50941 , n50942 );
xnor ( n50944 , n50943 , n41373 );
and ( n50945 , n50940 , n50944 );
xor ( n50946 , n50819 , n50833 );
xor ( n50947 , n50946 , n50836 );
and ( n50948 , n50944 , n50947 );
and ( n50949 , n50940 , n50947 );
or ( n50950 , n50945 , n50948 , n50949 );
and ( n50951 , n48099 , n41981 );
and ( n50952 , n47927 , n41979 );
nor ( n50953 , n50951 , n50952 );
xnor ( n50954 , n50953 , n41373 );
and ( n50955 , n50950 , n50954 );
xor ( n50956 , n50839 , n50841 );
xor ( n50957 , n50956 , n50844 );
and ( n50958 , n50954 , n50957 );
and ( n50959 , n50950 , n50957 );
or ( n50960 , n50955 , n50958 , n50959 );
and ( n50961 , n47927 , n41981 );
and ( n50962 , n47932 , n41979 );
nor ( n50963 , n50961 , n50962 );
xnor ( n50964 , n50963 , n41373 );
and ( n50965 , n50960 , n50964 );
xor ( n50966 , n50847 , n50849 );
xor ( n50967 , n50966 , n50852 );
and ( n50968 , n50964 , n50967 );
and ( n50969 , n50960 , n50967 );
or ( n50970 , n50965 , n50968 , n50969 );
and ( n50971 , n47932 , n41981 );
and ( n50972 , n47645 , n41979 );
nor ( n50973 , n50971 , n50972 );
xnor ( n50974 , n50973 , n41373 );
and ( n50975 , n50970 , n50974 );
xor ( n50976 , n50855 , n50857 );
xor ( n50977 , n50976 , n50860 );
and ( n50978 , n50974 , n50977 );
and ( n50979 , n50970 , n50977 );
or ( n50980 , n50975 , n50978 , n50979 );
and ( n50981 , n47645 , n41981 );
and ( n50982 , n46948 , n41979 );
nor ( n50983 , n50981 , n50982 );
xnor ( n50984 , n50983 , n41373 );
and ( n50985 , n50980 , n50984 );
xor ( n50986 , n50863 , n50865 );
xor ( n50987 , n50986 , n50868 );
and ( n50988 , n50984 , n50987 );
and ( n50989 , n50980 , n50987 );
or ( n50990 , n50985 , n50988 , n50989 );
and ( n50991 , n46948 , n41981 );
and ( n50992 , n46777 , n41979 );
nor ( n50993 , n50991 , n50992 );
xnor ( n50994 , n50993 , n41373 );
and ( n50995 , n50990 , n50994 );
xor ( n50996 , n50871 , n50873 );
xor ( n50997 , n50996 , n50876 );
and ( n50998 , n50994 , n50997 );
and ( n50999 , n50990 , n50997 );
or ( n51000 , n50995 , n50998 , n50999 );
and ( n51001 , n46777 , n41981 );
and ( n51002 , n46676 , n41979 );
nor ( n51003 , n51001 , n51002 );
xnor ( n51004 , n51003 , n41373 );
and ( n51005 , n51000 , n51004 );
xor ( n51006 , n50879 , n50883 );
xor ( n51007 , n51006 , n50886 );
and ( n51008 , n51004 , n51007 );
and ( n51009 , n51000 , n51007 );
or ( n51010 , n51005 , n51008 , n51009 );
and ( n51011 , n46676 , n41981 );
and ( n51012 , n46510 , n41979 );
nor ( n51013 , n51011 , n51012 );
xnor ( n51014 , n51013 , n41373 );
and ( n51015 , n51010 , n51014 );
xor ( n51016 , n50889 , n50893 );
xor ( n51017 , n51016 , n50896 );
and ( n51018 , n51014 , n51017 );
and ( n51019 , n51010 , n51017 );
or ( n51020 , n51015 , n51018 , n51019 );
and ( n51021 , n46510 , n41981 );
and ( n51022 , n46159 , n41979 );
nor ( n51023 , n51021 , n51022 );
xnor ( n51024 , n51023 , n41373 );
and ( n51025 , n51020 , n51024 );
xor ( n51026 , n50818 , n50899 );
xor ( n51027 , n51026 , n50902 );
and ( n51028 , n51024 , n51027 );
and ( n51029 , n51020 , n51027 );
or ( n51030 , n51025 , n51028 , n51029 );
and ( n51031 , n46159 , n41981 );
and ( n51032 , n46069 , n41979 );
nor ( n51033 , n51031 , n51032 );
xnor ( n51034 , n51033 , n41373 );
and ( n51035 , n51030 , n51034 );
xor ( n51036 , n50747 , n50905 );
xor ( n51037 , n51036 , n50908 );
and ( n51038 , n51034 , n51037 );
and ( n51039 , n51030 , n51037 );
or ( n51040 , n51035 , n51038 , n51039 );
and ( n51041 , n50911 , n51040 );
xor ( n51042 , n50696 , n50700 );
xor ( n51043 , n51042 , n50703 );
and ( n51044 , n51040 , n51043 );
and ( n51045 , n50911 , n51043 );
or ( n51046 , n51041 , n51044 , n51045 );
and ( n51047 , n45754 , n41981 );
and ( n51048 , n45171 , n41979 );
nor ( n51049 , n51047 , n51048 );
xnor ( n51050 , n51049 , n41373 );
and ( n51051 , n51046 , n51050 );
xor ( n51052 , n50706 , n50710 );
xor ( n51053 , n51052 , n50713 );
and ( n51054 , n51050 , n51053 );
and ( n51055 , n51046 , n51053 );
or ( n51056 , n51051 , n51054 , n51055 );
and ( n51057 , n45171 , n41981 );
and ( n51058 , n45057 , n41979 );
nor ( n51059 , n51057 , n51058 );
xnor ( n51060 , n51059 , n41373 );
and ( n51061 , n51056 , n51060 );
xor ( n51062 , n50692 , n50716 );
xor ( n51063 , n51062 , n50719 );
and ( n51064 , n51060 , n51063 );
and ( n51065 , n51056 , n51063 );
or ( n51066 , n51061 , n51064 , n51065 );
and ( n51067 , n50735 , n51066 );
and ( n51068 , n44826 , n42079 );
and ( n51069 , n44347 , n42076 );
nor ( n51070 , n51068 , n51069 );
xnor ( n51071 , n51070 , n41370 );
xor ( n51072 , n51056 , n51060 );
xor ( n51073 , n51072 , n51063 );
and ( n51074 , n51071 , n51073 );
and ( n51075 , n45057 , n42079 );
and ( n51076 , n44826 , n42076 );
nor ( n51077 , n51075 , n51076 );
xnor ( n51078 , n51077 , n41370 );
xor ( n51079 , n51046 , n51050 );
xor ( n51080 , n51079 , n51053 );
and ( n51081 , n51078 , n51080 );
and ( n51082 , n45171 , n42079 );
and ( n51083 , n45057 , n42076 );
nor ( n51084 , n51082 , n51083 );
xnor ( n51085 , n51084 , n41370 );
xor ( n51086 , n50911 , n51040 );
xor ( n51087 , n51086 , n51043 );
and ( n51088 , n51085 , n51087 );
and ( n51089 , n45754 , n42079 );
and ( n51090 , n45171 , n42076 );
nor ( n51091 , n51089 , n51090 );
xnor ( n51092 , n51091 , n41370 );
xor ( n51093 , n51030 , n51034 );
xor ( n51094 , n51093 , n51037 );
and ( n51095 , n51092 , n51094 );
and ( n51096 , n46069 , n42079 );
and ( n51097 , n45754 , n42076 );
nor ( n51098 , n51096 , n51097 );
xnor ( n51099 , n51098 , n41370 );
xor ( n51100 , n51020 , n51024 );
xor ( n51101 , n51100 , n51027 );
and ( n51102 , n51099 , n51101 );
and ( n51103 , n46159 , n42079 );
and ( n51104 , n46069 , n42076 );
nor ( n51105 , n51103 , n51104 );
xnor ( n51106 , n51105 , n41370 );
xor ( n51107 , n51010 , n51014 );
xor ( n51108 , n51107 , n51017 );
and ( n51109 , n51106 , n51108 );
and ( n51110 , n46510 , n42079 );
and ( n51111 , n46159 , n42076 );
nor ( n51112 , n51110 , n51111 );
xnor ( n51113 , n51112 , n41370 );
xor ( n51114 , n51000 , n51004 );
xor ( n51115 , n51114 , n51007 );
and ( n51116 , n51113 , n51115 );
and ( n51117 , n46676 , n42079 );
and ( n51118 , n46510 , n42076 );
nor ( n51119 , n51117 , n51118 );
xnor ( n51120 , n51119 , n41370 );
xor ( n51121 , n50990 , n50994 );
xor ( n51122 , n51121 , n50997 );
and ( n51123 , n51120 , n51122 );
and ( n51124 , n46777 , n42079 );
and ( n51125 , n46676 , n42076 );
nor ( n51126 , n51124 , n51125 );
xnor ( n51127 , n51126 , n41370 );
xor ( n51128 , n50980 , n50984 );
xor ( n51129 , n51128 , n50987 );
and ( n51130 , n51127 , n51129 );
and ( n51131 , n46948 , n42079 );
and ( n51132 , n46777 , n42076 );
nor ( n51133 , n51131 , n51132 );
xnor ( n51134 , n51133 , n41370 );
xor ( n51135 , n50970 , n50974 );
xor ( n51136 , n51135 , n50977 );
and ( n51137 , n51134 , n51136 );
and ( n51138 , n47645 , n42079 );
and ( n51139 , n46948 , n42076 );
nor ( n51140 , n51138 , n51139 );
xnor ( n51141 , n51140 , n41370 );
xor ( n51142 , n50960 , n50964 );
xor ( n51143 , n51142 , n50967 );
and ( n51144 , n51141 , n51143 );
and ( n51145 , n47932 , n42079 );
and ( n51146 , n47645 , n42076 );
nor ( n51147 , n51145 , n51146 );
xnor ( n51148 , n51147 , n41370 );
xor ( n51149 , n50950 , n50954 );
xor ( n51150 , n51149 , n50957 );
and ( n51151 , n51148 , n51150 );
and ( n51152 , n47927 , n42079 );
and ( n51153 , n47932 , n42076 );
nor ( n51154 , n51152 , n51153 );
xnor ( n51155 , n51154 , n41370 );
xor ( n51156 , n50940 , n50944 );
xor ( n51157 , n51156 , n50947 );
and ( n51158 , n51155 , n51157 );
and ( n51159 , n48099 , n42079 );
and ( n51160 , n47927 , n42076 );
nor ( n51161 , n51159 , n51160 );
xnor ( n51162 , n51161 , n41370 );
xor ( n51163 , n50930 , n50934 );
xor ( n51164 , n51163 , n50937 );
and ( n51165 , n51162 , n51164 );
and ( n51166 , n48086 , n42079 );
and ( n51167 , n48099 , n42076 );
nor ( n51168 , n51166 , n51167 );
xnor ( n51169 , n51168 , n41370 );
xor ( n51170 , n50912 , n50924 );
xor ( n51171 , n51170 , n50927 );
and ( n51172 , n51169 , n51171 );
and ( n51173 , n48077 , n42079 );
and ( n51174 , n48086 , n42076 );
nor ( n51175 , n51173 , n51174 );
xnor ( n51176 , n51175 , n41370 );
xor ( n51177 , n50918 , n50820 );
xor ( n51178 , n51177 , n50921 );
and ( n51179 , n51176 , n51178 );
and ( n51180 , n48069 , n42079 );
and ( n51181 , n48077 , n42076 );
nor ( n51182 , n51180 , n51181 );
xnor ( n51183 , n51182 , n41370 );
xor ( n51184 , n50915 , n50917 );
and ( n51185 , n51183 , n51184 );
buf ( n51186 , n30409 );
not ( n51187 , n51186 );
or ( n51188 , n50913 , n51187 );
and ( n51189 , n51184 , n51188 );
and ( n51190 , n51183 , n51188 );
or ( n51191 , n51185 , n51189 , n51190 );
and ( n51192 , n51178 , n51191 );
and ( n51193 , n51176 , n51191 );
or ( n51194 , n51179 , n51192 , n51193 );
and ( n51195 , n51171 , n51194 );
and ( n51196 , n51169 , n51194 );
or ( n51197 , n51172 , n51195 , n51196 );
and ( n51198 , n51164 , n51197 );
and ( n51199 , n51162 , n51197 );
or ( n51200 , n51165 , n51198 , n51199 );
and ( n51201 , n51157 , n51200 );
and ( n51202 , n51155 , n51200 );
or ( n51203 , n51158 , n51201 , n51202 );
and ( n51204 , n51150 , n51203 );
and ( n51205 , n51148 , n51203 );
or ( n51206 , n51151 , n51204 , n51205 );
and ( n51207 , n51143 , n51206 );
and ( n51208 , n51141 , n51206 );
or ( n51209 , n51144 , n51207 , n51208 );
and ( n51210 , n51136 , n51209 );
and ( n51211 , n51134 , n51209 );
or ( n51212 , n51137 , n51210 , n51211 );
and ( n51213 , n51129 , n51212 );
and ( n51214 , n51127 , n51212 );
or ( n51215 , n51130 , n51213 , n51214 );
and ( n51216 , n51122 , n51215 );
and ( n51217 , n51120 , n51215 );
or ( n51218 , n51123 , n51216 , n51217 );
and ( n51219 , n51115 , n51218 );
and ( n51220 , n51113 , n51218 );
or ( n51221 , n51116 , n51219 , n51220 );
and ( n51222 , n51108 , n51221 );
and ( n51223 , n51106 , n51221 );
or ( n51224 , n51109 , n51222 , n51223 );
and ( n51225 , n51101 , n51224 );
and ( n51226 , n51099 , n51224 );
or ( n51227 , n51102 , n51225 , n51226 );
and ( n51228 , n51094 , n51227 );
and ( n51229 , n51092 , n51227 );
or ( n51230 , n51095 , n51228 , n51229 );
and ( n51231 , n51087 , n51230 );
and ( n51232 , n51085 , n51230 );
or ( n51233 , n51088 , n51231 , n51232 );
and ( n51234 , n51080 , n51233 );
and ( n51235 , n51078 , n51233 );
or ( n51236 , n51081 , n51234 , n51235 );
and ( n51237 , n51073 , n51236 );
and ( n51238 , n51071 , n51236 );
or ( n51239 , n51074 , n51237 , n51238 );
and ( n51240 , n51066 , n51239 );
and ( n51241 , n50735 , n51239 );
or ( n51242 , n51067 , n51240 , n51241 );
and ( n51243 , n50732 , n51242 );
and ( n51244 , n50591 , n51242 );
or ( n51245 , n50733 , n51243 , n51244 );
and ( n51246 , n50588 , n51245 );
and ( n51247 , n50564 , n51245 );
or ( n51248 , n50589 , n51246 , n51247 );
and ( n51249 , n50561 , n51248 );
and ( n51250 , n50559 , n51248 );
or ( n51251 , n50562 , n51249 , n51250 );
or ( n51252 , n50491 , n51251 );
or ( n51253 , n50489 , n51252 );
and ( n51254 , n50486 , n51253 );
and ( n51255 , n50416 , n51253 );
or ( n51256 , n50487 , n51254 , n51255 );
or ( n51257 , n50414 , n51256 );
or ( n51258 , n50412 , n51257 );
and ( n51259 , n50410 , n51258 );
xor ( n51260 , n50410 , n51258 );
xnor ( n51261 , n50412 , n51257 );
xnor ( n51262 , n50414 , n51256 );
xor ( n51263 , n50416 , n50486 );
xor ( n51264 , n51263 , n51253 );
and ( n51265 , n51262 , n51264 );
and ( n51266 , n51261 , n51265 );
and ( n51267 , n51260 , n51266 );
or ( n51268 , n51259 , n51267 );
and ( n51269 , n50408 , n51268 );
and ( n51270 , n50406 , n51269 );
or ( n51271 , n50405 , n51270 );
and ( n51272 , n49665 , n51271 );
and ( n51273 , n49663 , n51272 );
and ( n51274 , n49661 , n51273 );
and ( n51275 , n49660 , n51274 );
or ( n51276 , n49659 , n51275 );
and ( n51277 , n49263 , n51276 );
and ( n51278 , n49261 , n51277 );
and ( n51279 , n49260 , n51278 );
and ( n51280 , n49259 , n51279 );
or ( n51281 , n49258 , n51280 );
and ( n51282 , n49256 , n51281 );
or ( n51283 , n49255 , n51282 );
and ( n51284 , n48398 , n51283 );
and ( n51285 , n48397 , n51284 );
or ( n51286 , n48396 , n51285 );
and ( n51287 , n48394 , n51286 );
and ( n51288 , n48392 , n51287 );
or ( n51289 , n48391 , n51288 );
and ( n51290 , n47628 , n51289 );
and ( n51291 , n47627 , n51290 );
and ( n51292 , n47626 , n51291 );
or ( n51293 , n47625 , n51292 );
and ( n51294 , n47228 , n51293 );
and ( n51295 , n47226 , n51294 );
or ( n51296 , n47225 , n51295 );
and ( n51297 , n47223 , n51296 );
and ( n51298 , n47221 , n51297 );
or ( n51299 , n47220 , n51298 );
and ( n51300 , n46488 , n51299 );
or ( n51301 , n46487 , n51300 );
and ( n51302 , n46485 , n51301 );
and ( n51303 , n46484 , n51302 );
and ( n51304 , n46483 , n51303 );
or ( n51305 , n46482 , n51304 );
and ( n51306 , n46478 , n51305 );
or ( n51307 , n46477 , n51306 );
and ( n51308 , n45951 , n51307 );
and ( n51309 , n45950 , n51308 );
or ( n51310 , n45949 , n51309 );
and ( n51311 , n45699 , n51310 );
and ( n51312 , n45697 , n51311 );
and ( n51313 , n45696 , n51312 );
or ( n51314 , n45695 , n51313 );
and ( n51315 , n45693 , n51314 );
or ( n51316 , n45692 , n51315 );
and ( n51317 , n44729 , n51316 );
and ( n51318 , n44727 , n51317 );
or ( n51319 , n44726 , n51318 );
and ( n51320 , n44724 , n51319 );
or ( n51321 , n44723 , n51320 );
and ( n51322 , n44109 , n51321 );
and ( n51323 , n44108 , n51322 );
or ( n51324 , n44107 , n51323 );
and ( n51325 , n43471 , n51324 );
and ( n51326 , n43469 , n51325 );
or ( n51327 , n43468 , n51326 );
and ( n51328 , n43466 , n51327 );
or ( n51329 , n43465 , n51328 );
and ( n51330 , n43285 , n51329 );
or ( n51331 , n43284 , n51330 );
and ( n51332 , n43280 , n51331 );
and ( n51333 , n43278 , n51332 );
or ( n51334 , n43277 , n51333 );
and ( n51335 , n43275 , n51334 );
and ( n51336 , n43274 , n51335 );
and ( n51337 , n43273 , n51336 );
and ( n51338 , n43272 , n51337 );
and ( n51339 , n43271 , n51338 );
and ( n51340 , n43270 , n51339 );
and ( n51341 , n43269 , n51340 );
and ( n51342 , n43268 , n51341 );
and ( n51343 , n43267 , n51342 );
and ( n51344 , n43266 , n51343 );
and ( n51345 , n43265 , n51344 );
and ( n51346 , n43264 , n51345 );
and ( n51347 , n43263 , n51346 );
and ( n51348 , n43262 , n51347 );
and ( n51349 , n43261 , n51348 );
and ( n51350 , n43260 , n51349 );
and ( n51351 , n43259 , n51350 );
and ( n51352 , n43258 , n51351 );
and ( n51353 , n43257 , n51352 );
and ( n51354 , n43256 , n51353 );
and ( n51355 , n43255 , n51354 );
and ( n51356 , n43254 , n51355 );
and ( n51357 , n43253 , n51356 );
and ( n51358 , n43252 , n51357 );
and ( n51359 , n43251 , n51358 );
and ( n51360 , n43250 , n51359 );
and ( n51361 , n43248 , n51360 );
or ( n51362 , n43247 , n51361 );
and ( n51363 , n43245 , n51362 );
buf ( n51364 , n51363 );
buf ( n51365 , n51364 );
buf ( n51366 , n51365 );
buf ( n51367 , n51366 );
buf ( n51368 , n51367 );
buf ( n51369 , n51368 );
buf ( n51370 , n51369 );
buf ( n51371 , n51370 );
buf ( n51372 , n51371 );
buf ( n51373 , n51372 );
buf ( n51374 , n51373 );
buf ( n51375 , n51374 );
buf ( n51376 , n51375 );
buf ( n51377 , n51376 );
buf ( n51378 , n51377 );
buf ( n51379 , n51378 );
buf ( n51380 , n51379 );
buf ( n51381 , n51380 );
buf ( n51382 , n51381 );
buf ( n51383 , n51382 );
buf ( n51384 , n51383 );
buf ( n51385 , n51384 );
buf ( n51386 , n51385 );
buf ( n51387 , n51386 );
buf ( n51388 , n51387 );
buf ( n51389 , n51388 );
buf ( n51390 , n51389 );
buf ( n51391 , n51390 );
not ( n51392 , n51391 );
buf ( n51393 , n51392 );
not ( n51394 , n51390 );
buf ( n51395 , n51394 );
not ( n51396 , n51389 );
buf ( n51397 , n51396 );
not ( n51398 , n51388 );
buf ( n51399 , n51398 );
not ( n51400 , n51387 );
buf ( n51401 , n51400 );
not ( n51402 , n51386 );
buf ( n51403 , n51402 );
not ( n51404 , n51385 );
buf ( n51405 , n51404 );
not ( n51406 , n51384 );
buf ( n51407 , n51406 );
not ( n51408 , n51383 );
buf ( n51409 , n51408 );
not ( n51410 , n51382 );
buf ( n51411 , n51410 );
not ( n51412 , n51381 );
buf ( n51413 , n51412 );
not ( n51414 , n51380 );
buf ( n51415 , n51414 );
not ( n51416 , n51379 );
buf ( n51417 , n51416 );
not ( n51418 , n51378 );
buf ( n51419 , n51418 );
not ( n51420 , n51377 );
buf ( n51421 , n51420 );
not ( n51422 , n51376 );
buf ( n51423 , n51422 );
not ( n51424 , n51375 );
buf ( n51425 , n51424 );
not ( n51426 , n51374 );
buf ( n51427 , n51426 );
not ( n51428 , n51373 );
buf ( n51429 , n51428 );
not ( n51430 , n51372 );
buf ( n51431 , n51430 );
not ( n51432 , n51371 );
buf ( n51433 , n51432 );
not ( n51434 , n51370 );
buf ( n51435 , n51434 );
not ( n51436 , n51369 );
buf ( n51437 , n51436 );
not ( n51438 , n51368 );
buf ( n51439 , n51438 );
not ( n51440 , n51367 );
buf ( n51441 , n51440 );
not ( n51442 , n51366 );
buf ( n51443 , n51442 );
not ( n51444 , n51365 );
buf ( n51445 , n51444 );
not ( n51446 , n51364 );
buf ( n51447 , n51446 );
not ( n51448 , n51363 );
buf ( n51449 , n51448 );
xor ( n51450 , n43245 , n51362 );
buf ( n51451 , n51450 );
xor ( n51452 , n43248 , n51360 );
buf ( n51453 , n51452 );
xor ( n51454 , n43250 , n51359 );
buf ( n51455 , n51454 );
xor ( n51456 , n43251 , n51358 );
buf ( n51457 , n51456 );
xor ( n51458 , n43252 , n51357 );
buf ( n51459 , n51458 );
xor ( n51460 , n43253 , n51356 );
buf ( n51461 , n51460 );
xor ( n51462 , n43254 , n51355 );
buf ( n51463 , n51462 );
xor ( n51464 , n43255 , n51354 );
buf ( n51465 , n51464 );
xor ( n51466 , n43256 , n51353 );
buf ( n51467 , n51466 );
xor ( n51468 , n43257 , n51352 );
buf ( n51469 , n51468 );
xor ( n51470 , n43258 , n51351 );
buf ( n51471 , n51470 );
xor ( n51472 , n43259 , n51350 );
buf ( n51473 , n51472 );
xor ( n51474 , n43260 , n51349 );
buf ( n51475 , n51474 );
xor ( n51476 , n43261 , n51348 );
buf ( n51477 , n51476 );
xor ( n51478 , n43262 , n51347 );
buf ( n51479 , n51478 );
xor ( n51480 , n43263 , n51346 );
buf ( n51481 , n51480 );
xor ( n51482 , n43264 , n51345 );
buf ( n51483 , n51482 );
xor ( n51484 , n43265 , n51344 );
buf ( n51485 , n51484 );
xor ( n51486 , n43266 , n51343 );
buf ( n51487 , n51486 );
xor ( n51488 , n43267 , n51342 );
buf ( n51489 , n51488 );
xor ( n51490 , n43268 , n51341 );
buf ( n51491 , n51490 );
xor ( n51492 , n43269 , n51340 );
buf ( n51493 , n51492 );
xor ( n51494 , n43270 , n51339 );
buf ( n51495 , n51494 );
xor ( n51496 , n43271 , n51338 );
buf ( n51497 , n51496 );
xor ( n51498 , n43272 , n51337 );
buf ( n51499 , n51498 );
xor ( n51500 , n43273 , n51336 );
buf ( n51501 , n51500 );
xor ( n51502 , n43274 , n51335 );
buf ( n51503 , n51502 );
xor ( n51504 , n43275 , n51334 );
buf ( n51505 , n51504 );
xor ( n51506 , n43278 , n51332 );
buf ( n51507 , n51506 );
xor ( n51508 , n43280 , n51331 );
buf ( n51509 , n51508 );
xor ( n51510 , n43285 , n51329 );
buf ( n51511 , n51510 );
xor ( n51512 , n43466 , n51327 );
buf ( n51513 , n51512 );
xor ( n51514 , n43469 , n51325 );
buf ( n51515 , n51514 );
xor ( n51516 , n43471 , n51324 );
buf ( n51517 , n51516 );
xor ( n51518 , n44108 , n51322 );
buf ( n51519 , n51518 );
xor ( n51520 , n44109 , n51321 );
buf ( n51521 , n51520 );
xor ( n51522 , n44724 , n51319 );
buf ( n51523 , n51522 );
xor ( n51524 , n44727 , n51317 );
buf ( n51525 , n51524 );
xor ( n51526 , n44729 , n51316 );
buf ( n51527 , n51526 );
xor ( n51528 , n45693 , n51314 );
buf ( n51529 , n51528 );
xor ( n51530 , n45696 , n51312 );
buf ( n51531 , n51530 );
xor ( n51532 , n45697 , n51311 );
buf ( n51533 , n51532 );
xor ( n51534 , n45699 , n51310 );
buf ( n51535 , n51534 );
xor ( n51536 , n45950 , n51308 );
buf ( n51537 , n51536 );
xor ( n51538 , n45951 , n51307 );
buf ( n51539 , n51538 );
xor ( n51540 , n46478 , n51305 );
buf ( n51541 , n51540 );
xor ( n51542 , n46483 , n51303 );
buf ( n51543 , n51542 );
xor ( n51544 , n46484 , n51302 );
buf ( n51545 , n51544 );
xor ( n51546 , n46485 , n51301 );
buf ( n51547 , n51546 );
xor ( n51548 , n46488 , n51299 );
buf ( n51549 , n51548 );
xor ( n51550 , n47221 , n51297 );
buf ( n51551 , n51550 );
xor ( n51552 , n47223 , n51296 );
buf ( n51553 , n51552 );
xor ( n51554 , n47226 , n51294 );
buf ( n51555 , n51554 );
xor ( n51556 , n47228 , n51293 );
buf ( n51557 , n51556 );
xor ( n51558 , n47626 , n51291 );
buf ( n51559 , n51558 );
xor ( n51560 , n47627 , n51290 );
buf ( n51561 , n51560 );
xor ( n51562 , n47628 , n51289 );
buf ( n51563 , n51562 );
xor ( n51564 , n48392 , n51287 );
buf ( n51565 , n51564 );
xor ( n51566 , n48394 , n51286 );
buf ( n51567 , n51566 );
xor ( n51568 , n48397 , n51284 );
buf ( n51569 , n51568 );
xor ( n51570 , n48398 , n51283 );
buf ( n51571 , n51570 );
xor ( n51572 , n49256 , n51281 );
buf ( n51573 , n51572 );
xor ( n51574 , n49259 , n51279 );
buf ( n51575 , n51574 );
xor ( n51576 , n49260 , n51278 );
buf ( n51577 , n51576 );
xor ( n51578 , n49261 , n51277 );
buf ( n51579 , n51578 );
xor ( n51580 , n49263 , n51276 );
buf ( n51581 , n51580 );
xor ( n51582 , n49660 , n51274 );
buf ( n51583 , n51582 );
xor ( n51584 , n49661 , n51273 );
buf ( n51585 , n51584 );
xor ( n51586 , n49663 , n51272 );
buf ( n51587 , n51586 );
xor ( n51588 , n49665 , n51271 );
buf ( n51589 , n51588 );
xor ( n51590 , n50406 , n51269 );
buf ( n51591 , n51590 );
xor ( n51592 , n50408 , n51268 );
buf ( n51593 , n51592 );
xor ( n51594 , n51260 , n51266 );
buf ( n51595 , n51594 );
xor ( n51596 , n51261 , n51265 );
buf ( n51597 , n51596 );
xor ( n51598 , n51262 , n51264 );
buf ( n51599 , n51598 );
not ( n51600 , n51264 );
buf ( n51601 , n51600 );
xnor ( n51602 , n50489 , n51252 );
buf ( n51603 , n51602 );
xnor ( n51604 , n50491 , n51251 );
buf ( n51605 , n51604 );
xor ( n51606 , n50559 , n50561 );
xor ( n51607 , n51606 , n51248 );
buf ( n51608 , n51607 );
xor ( n51609 , n50564 , n50588 );
xor ( n51610 , n51609 , n51245 );
buf ( n51611 , n51610 );
xor ( n51612 , n50591 , n50732 );
xor ( n51613 , n51612 , n51242 );
buf ( n51614 , n51613 );
xor ( n51615 , n50735 , n51066 );
xor ( n51616 , n51615 , n51239 );
buf ( n51617 , n51616 );
xor ( n51618 , n51071 , n51073 );
xor ( n51619 , n51618 , n51236 );
buf ( n51620 , n51619 );
xor ( n51621 , n51078 , n51080 );
xor ( n51622 , n51621 , n51233 );
buf ( n51623 , n51622 );
xor ( n51624 , n51085 , n51087 );
xor ( n51625 , n51624 , n51230 );
buf ( n51626 , n51625 );
xor ( n51627 , n51092 , n51094 );
xor ( n51628 , n51627 , n51227 );
buf ( n51629 , n51628 );
xor ( n51630 , n51099 , n51101 );
xor ( n51631 , n51630 , n51224 );
buf ( n51632 , n51631 );
xor ( n51633 , n51106 , n51108 );
xor ( n51634 , n51633 , n51221 );
buf ( n51635 , n51634 );
xor ( n51636 , n51113 , n51115 );
xor ( n51637 , n51636 , n51218 );
buf ( n51638 , n51637 );
xor ( n51639 , n51120 , n51122 );
xor ( n51640 , n51639 , n51215 );
buf ( n51641 , n51640 );
xor ( n51642 , n51127 , n51129 );
xor ( n51643 , n51642 , n51212 );
buf ( n51644 , n51643 );
xor ( n51645 , n51134 , n51136 );
xor ( n51646 , n51645 , n51209 );
buf ( n51647 , n51646 );
xor ( n51648 , n51141 , n51143 );
xor ( n51649 , n51648 , n51206 );
buf ( n51650 , n51649 );
xor ( n51651 , n51148 , n51150 );
xor ( n51652 , n51651 , n51203 );
buf ( n51653 , n51652 );
xor ( n51654 , n51155 , n51157 );
xor ( n51655 , n51654 , n51200 );
buf ( n51656 , n51655 );
xor ( n51657 , n51162 , n51164 );
xor ( n51658 , n51657 , n51197 );
buf ( n51659 , n51658 );
xor ( n51660 , n51169 , n51171 );
xor ( n51661 , n51660 , n51194 );
buf ( n51662 , n51661 );
xor ( n51663 , n51176 , n51178 );
xor ( n51664 , n51663 , n51191 );
buf ( n51665 , n51664 );
xor ( n51666 , n51183 , n51184 );
xor ( n51667 , n51666 , n51188 );
buf ( n51668 , n51667 );
xnor ( n51669 , n50913 , n51187 );
buf ( n51670 , n51669 );
buf ( n51671 , n30153 );
buf ( n51672 , n30156 );
buf ( n51673 , n30159 );
buf ( n51674 , n30162 );
buf ( n51675 , n30165 );
buf ( n51676 , n30168 );
buf ( n51677 , n30171 );
buf ( n51678 , n30174 );
buf ( n51679 , n30177 );
buf ( n51680 , n30180 );
buf ( n51681 , n30183 );
buf ( n51682 , n30186 );
buf ( n51683 , n30189 );
buf ( n51684 , n30192 );
buf ( n51685 , n30195 );
buf ( n51686 , n30198 );
buf ( n51687 , n30201 );
buf ( n51688 , n30204 );
buf ( n51689 , n30207 );
buf ( n51690 , n30210 );
buf ( n51691 , n30213 );
buf ( n51692 , n30216 );
buf ( n51693 , n30219 );
buf ( n51694 , n30222 );
buf ( n51695 , n30225 );
buf ( n51696 , n30228 );
buf ( n51697 , n30231 );
buf ( n51698 , n30234 );
buf ( n51699 , n30237 );
buf ( n51700 , n30240 );
buf ( n51701 , n30243 );
buf ( n51702 , n30246 );
buf ( n51703 , n30249 );
buf ( n51704 , n30252 );
buf ( n51705 , n30255 );
buf ( n51706 , n30258 );
buf ( n51707 , n30261 );
buf ( n51708 , n30264 );
buf ( n51709 , n30267 );
buf ( n51710 , n30270 );
buf ( n51711 , n30273 );
buf ( n51712 , n30276 );
buf ( n51713 , n30279 );
buf ( n51714 , n30282 );
buf ( n51715 , n30285 );
buf ( n51716 , n30288 );
buf ( n51717 , n30291 );
buf ( n51718 , n30294 );
buf ( n51719 , n30297 );
buf ( n51720 , n30300 );
buf ( n51721 , n30303 );
buf ( n51722 , n30306 );
buf ( n51723 , n30309 );
buf ( n51724 , n30312 );
buf ( n51725 , n30315 );
buf ( n51726 , n30318 );
buf ( n51727 , n30321 );
buf ( n51728 , n30324 );
buf ( n51729 , n30327 );
buf ( n51730 , n30330 );
buf ( n51731 , n30333 );
buf ( n51732 , n30336 );
buf ( n51733 , n30339 );
buf ( n51734 , n30342 );
buf ( n51735 , n30344 );
buf ( n51736 , n1218 );
buf ( n51737 , n1186 );
and ( n51738 , n51736 , n51737 );
buf ( n51739 , n1219 );
buf ( n51740 , n1187 );
and ( n51741 , n51739 , n51740 );
buf ( n51742 , n1220 );
buf ( n51743 , n1188 );
and ( n51744 , n51742 , n51743 );
buf ( n51745 , n1221 );
buf ( n51746 , n1189 );
and ( n51747 , n51745 , n51746 );
buf ( n51748 , n1222 );
buf ( n51749 , n1190 );
and ( n51750 , n51748 , n51749 );
buf ( n51751 , n1223 );
buf ( n51752 , n1191 );
and ( n51753 , n51751 , n51752 );
buf ( n51754 , n1224 );
buf ( n51755 , n1192 );
and ( n51756 , n51754 , n51755 );
buf ( n51757 , n1225 );
buf ( n51758 , n1193 );
and ( n51759 , n51757 , n51758 );
buf ( n51760 , n1226 );
buf ( n51761 , n1194 );
and ( n51762 , n51760 , n51761 );
buf ( n51763 , n1227 );
buf ( n51764 , n1195 );
and ( n51765 , n51763 , n51764 );
buf ( n51766 , n1228 );
buf ( n51767 , n1196 );
and ( n51768 , n51766 , n51767 );
buf ( n51769 , n1229 );
buf ( n51770 , n1197 );
and ( n51771 , n51769 , n51770 );
buf ( n51772 , n1230 );
buf ( n51773 , n1198 );
and ( n51774 , n51772 , n51773 );
buf ( n51775 , n1231 );
buf ( n51776 , n1199 );
and ( n51777 , n51775 , n51776 );
buf ( n51778 , n1232 );
buf ( n51779 , n1200 );
and ( n51780 , n51778 , n51779 );
buf ( n51781 , n1233 );
buf ( n51782 , n1201 );
and ( n51783 , n51781 , n51782 );
buf ( n51784 , n1234 );
buf ( n51785 , n1202 );
and ( n51786 , n51784 , n51785 );
buf ( n51787 , n1235 );
buf ( n51788 , n1203 );
and ( n51789 , n51787 , n51788 );
buf ( n51790 , n1236 );
buf ( n51791 , n1204 );
and ( n51792 , n51790 , n51791 );
buf ( n51793 , n1237 );
buf ( n51794 , n1205 );
and ( n51795 , n51793 , n51794 );
buf ( n51796 , n1238 );
buf ( n51797 , n1206 );
and ( n51798 , n51796 , n51797 );
buf ( n51799 , n1239 );
buf ( n51800 , n1207 );
and ( n51801 , n51799 , n51800 );
buf ( n51802 , n1240 );
buf ( n51803 , n1208 );
and ( n51804 , n51802 , n51803 );
buf ( n51805 , n1241 );
buf ( n51806 , n1209 );
and ( n51807 , n51805 , n51806 );
buf ( n51808 , n1242 );
buf ( n51809 , n1210 );
and ( n51810 , n51808 , n51809 );
buf ( n51811 , n1243 );
buf ( n51812 , n1211 );
and ( n51813 , n51811 , n51812 );
buf ( n51814 , n1244 );
buf ( n51815 , n1212 );
and ( n51816 , n51814 , n51815 );
buf ( n51817 , n1245 );
buf ( n51818 , n1213 );
and ( n51819 , n51817 , n51818 );
buf ( n51820 , n1246 );
buf ( n51821 , n1214 );
and ( n51822 , n51820 , n51821 );
buf ( n51823 , n1247 );
buf ( n51824 , n1215 );
and ( n51825 , n51823 , n51824 );
buf ( n51826 , n1248 );
buf ( n51827 , n1216 );
and ( n51828 , n51826 , n51827 );
buf ( n51829 , n1249 );
buf ( n51830 , n1217 );
and ( n51831 , n51829 , n51830 );
and ( n51832 , n51827 , n51831 );
and ( n51833 , n51826 , n51831 );
or ( n51834 , n51828 , n51832 , n51833 );
and ( n51835 , n51824 , n51834 );
and ( n51836 , n51823 , n51834 );
or ( n51837 , n51825 , n51835 , n51836 );
and ( n51838 , n51821 , n51837 );
and ( n51839 , n51820 , n51837 );
or ( n51840 , n51822 , n51838 , n51839 );
and ( n51841 , n51818 , n51840 );
and ( n51842 , n51817 , n51840 );
or ( n51843 , n51819 , n51841 , n51842 );
and ( n51844 , n51815 , n51843 );
and ( n51845 , n51814 , n51843 );
or ( n51846 , n51816 , n51844 , n51845 );
and ( n51847 , n51812 , n51846 );
and ( n51848 , n51811 , n51846 );
or ( n51849 , n51813 , n51847 , n51848 );
and ( n51850 , n51809 , n51849 );
and ( n51851 , n51808 , n51849 );
or ( n51852 , n51810 , n51850 , n51851 );
and ( n51853 , n51806 , n51852 );
and ( n51854 , n51805 , n51852 );
or ( n51855 , n51807 , n51853 , n51854 );
and ( n51856 , n51803 , n51855 );
and ( n51857 , n51802 , n51855 );
or ( n51858 , n51804 , n51856 , n51857 );
and ( n51859 , n51800 , n51858 );
and ( n51860 , n51799 , n51858 );
or ( n51861 , n51801 , n51859 , n51860 );
and ( n51862 , n51797 , n51861 );
and ( n51863 , n51796 , n51861 );
or ( n51864 , n51798 , n51862 , n51863 );
and ( n51865 , n51794 , n51864 );
and ( n51866 , n51793 , n51864 );
or ( n51867 , n51795 , n51865 , n51866 );
and ( n51868 , n51791 , n51867 );
and ( n51869 , n51790 , n51867 );
or ( n51870 , n51792 , n51868 , n51869 );
and ( n51871 , n51788 , n51870 );
and ( n51872 , n51787 , n51870 );
or ( n51873 , n51789 , n51871 , n51872 );
and ( n51874 , n51785 , n51873 );
and ( n51875 , n51784 , n51873 );
or ( n51876 , n51786 , n51874 , n51875 );
and ( n51877 , n51782 , n51876 );
and ( n51878 , n51781 , n51876 );
or ( n51879 , n51783 , n51877 , n51878 );
and ( n51880 , n51779 , n51879 );
and ( n51881 , n51778 , n51879 );
or ( n51882 , n51780 , n51880 , n51881 );
and ( n51883 , n51776 , n51882 );
and ( n51884 , n51775 , n51882 );
or ( n51885 , n51777 , n51883 , n51884 );
and ( n51886 , n51773 , n51885 );
and ( n51887 , n51772 , n51885 );
or ( n51888 , n51774 , n51886 , n51887 );
and ( n51889 , n51770 , n51888 );
and ( n51890 , n51769 , n51888 );
or ( n51891 , n51771 , n51889 , n51890 );
and ( n51892 , n51767 , n51891 );
and ( n51893 , n51766 , n51891 );
or ( n51894 , n51768 , n51892 , n51893 );
and ( n51895 , n51764 , n51894 );
and ( n51896 , n51763 , n51894 );
or ( n51897 , n51765 , n51895 , n51896 );
and ( n51898 , n51761 , n51897 );
and ( n51899 , n51760 , n51897 );
or ( n51900 , n51762 , n51898 , n51899 );
and ( n51901 , n51758 , n51900 );
and ( n51902 , n51757 , n51900 );
or ( n51903 , n51759 , n51901 , n51902 );
and ( n51904 , n51755 , n51903 );
and ( n51905 , n51754 , n51903 );
or ( n51906 , n51756 , n51904 , n51905 );
and ( n51907 , n51752 , n51906 );
and ( n51908 , n51751 , n51906 );
or ( n51909 , n51753 , n51907 , n51908 );
and ( n51910 , n51749 , n51909 );
and ( n51911 , n51748 , n51909 );
or ( n51912 , n51750 , n51910 , n51911 );
and ( n51913 , n51746 , n51912 );
and ( n51914 , n51745 , n51912 );
or ( n51915 , n51747 , n51913 , n51914 );
and ( n51916 , n51743 , n51915 );
and ( n51917 , n51742 , n51915 );
or ( n51918 , n51744 , n51916 , n51917 );
and ( n51919 , n51740 , n51918 );
and ( n51920 , n51739 , n51918 );
or ( n51921 , n51741 , n51919 , n51920 );
and ( n51922 , n51737 , n51921 );
and ( n51923 , n51736 , n51921 );
or ( n51924 , n51738 , n51922 , n51923 );
buf ( n51925 , n51924 );
buf ( n51926 , n51925 );
xor ( n51927 , n51736 , n51737 );
xor ( n51928 , n51927 , n51921 );
buf ( n51929 , n51928 );
buf ( n51930 , n51929 );
xor ( n51931 , n51739 , n51740 );
xor ( n51932 , n51931 , n51918 );
buf ( n51933 , n51932 );
buf ( n51934 , n51933 );
xor ( n51935 , n51742 , n51743 );
xor ( n51936 , n51935 , n51915 );
buf ( n51937 , n51936 );
buf ( n51938 , n51937 );
xor ( n51939 , n51745 , n51746 );
xor ( n51940 , n51939 , n51912 );
buf ( n51941 , n51940 );
buf ( n51942 , n51941 );
xor ( n51943 , n51748 , n51749 );
xor ( n51944 , n51943 , n51909 );
buf ( n51945 , n51944 );
buf ( n51946 , n51945 );
xor ( n51947 , n51751 , n51752 );
xor ( n51948 , n51947 , n51906 );
buf ( n51949 , n51948 );
buf ( n51950 , n51949 );
xor ( n51951 , n51754 , n51755 );
xor ( n51952 , n51951 , n51903 );
buf ( n51953 , n51952 );
buf ( n51954 , n51953 );
xor ( n51955 , n51757 , n51758 );
xor ( n51956 , n51955 , n51900 );
buf ( n51957 , n51956 );
buf ( n51958 , n51957 );
xor ( n51959 , n51760 , n51761 );
xor ( n51960 , n51959 , n51897 );
buf ( n51961 , n51960 );
buf ( n51962 , n51961 );
xor ( n51963 , n51763 , n51764 );
xor ( n51964 , n51963 , n51894 );
buf ( n51965 , n51964 );
buf ( n51966 , n51965 );
xor ( n51967 , n51766 , n51767 );
xor ( n51968 , n51967 , n51891 );
buf ( n51969 , n51968 );
buf ( n51970 , n51969 );
xor ( n51971 , n51769 , n51770 );
xor ( n51972 , n51971 , n51888 );
buf ( n51973 , n51972 );
buf ( n51974 , n51973 );
xor ( n51975 , n51772 , n51773 );
xor ( n51976 , n51975 , n51885 );
buf ( n51977 , n51976 );
buf ( n51978 , n51977 );
xor ( n51979 , n51775 , n51776 );
xor ( n51980 , n51979 , n51882 );
buf ( n51981 , n51980 );
buf ( n51982 , n51981 );
xor ( n51983 , n51778 , n51779 );
xor ( n51984 , n51983 , n51879 );
buf ( n51985 , n51984 );
buf ( n51986 , n51985 );
xor ( n51987 , n51781 , n51782 );
xor ( n51988 , n51987 , n51876 );
buf ( n51989 , n51988 );
buf ( n51990 , n51989 );
xor ( n51991 , n51784 , n51785 );
xor ( n51992 , n51991 , n51873 );
buf ( n51993 , n51992 );
buf ( n51994 , n51993 );
xor ( n51995 , n51787 , n51788 );
xor ( n51996 , n51995 , n51870 );
buf ( n51997 , n51996 );
buf ( n51998 , n51997 );
xor ( n51999 , n51790 , n51791 );
xor ( n52000 , n51999 , n51867 );
buf ( n52001 , n52000 );
buf ( n52002 , n52001 );
xor ( n52003 , n51793 , n51794 );
xor ( n52004 , n52003 , n51864 );
buf ( n52005 , n52004 );
buf ( n52006 , n52005 );
xor ( n52007 , n51796 , n51797 );
xor ( n52008 , n52007 , n51861 );
buf ( n52009 , n52008 );
buf ( n52010 , n52009 );
xor ( n52011 , n51799 , n51800 );
xor ( n52012 , n52011 , n51858 );
buf ( n52013 , n52012 );
buf ( n52014 , n52013 );
xor ( n52015 , n51802 , n51803 );
xor ( n52016 , n52015 , n51855 );
buf ( n52017 , n52016 );
buf ( n52018 , n52017 );
xor ( n52019 , n51805 , n51806 );
xor ( n52020 , n52019 , n51852 );
buf ( n52021 , n52020 );
buf ( n52022 , n52021 );
xor ( n52023 , n51808 , n51809 );
xor ( n52024 , n52023 , n51849 );
buf ( n52025 , n52024 );
buf ( n52026 , n52025 );
xor ( n52027 , n51811 , n51812 );
xor ( n52028 , n52027 , n51846 );
buf ( n52029 , n52028 );
buf ( n52030 , n52029 );
xor ( n52031 , n51814 , n51815 );
xor ( n52032 , n52031 , n51843 );
buf ( n52033 , n52032 );
buf ( n52034 , n52033 );
xor ( n52035 , n51817 , n51818 );
xor ( n52036 , n52035 , n51840 );
buf ( n52037 , n52036 );
buf ( n52038 , n52037 );
xor ( n52039 , n51820 , n51821 );
xor ( n52040 , n52039 , n51837 );
buf ( n52041 , n52040 );
buf ( n52042 , n52041 );
xor ( n52043 , n51823 , n51824 );
xor ( n52044 , n52043 , n51834 );
buf ( n52045 , n52044 );
buf ( n52046 , n52045 );
xor ( n52047 , n51826 , n51827 );
xor ( n52048 , n52047 , n51831 );
buf ( n52049 , n52048 );
buf ( n52050 , n52049 );
xor ( n52051 , n51829 , n51830 );
buf ( n52052 , n52051 );
buf ( n52053 , n52052 );
buf ( n52054 , n51671 );
buf ( n52055 , n51926 );
buf ( n52056 , n51930 );
xor ( n52057 , n52055 , n52056 );
not ( n52058 , n52057 );
and ( n52059 , n52055 , n52058 );
and ( n52060 , n52054 , n52059 );
buf ( n52061 , n51673 );
and ( n52062 , n52061 , n52059 );
buf ( n52063 , n51672 );
and ( n52064 , n52063 , n52057 );
nor ( n52065 , n52062 , n52064 );
not ( n52066 , n52065 );
buf ( n52067 , n52066 );
buf ( n52068 , n51934 );
buf ( n52069 , n51938 );
and ( n52070 , n52068 , n52069 );
not ( n52071 , n52070 );
and ( n52072 , n52056 , n52071 );
not ( n52073 , n52072 );
and ( n52074 , n52067 , n52073 );
and ( n52075 , n52063 , n52059 );
and ( n52076 , n52054 , n52057 );
nor ( n52077 , n52075 , n52076 );
not ( n52078 , n52077 );
and ( n52079 , n52073 , n52078 );
and ( n52080 , n52067 , n52078 );
or ( n52081 , n52074 , n52079 , n52080 );
xor ( n52082 , n52060 , n52081 );
buf ( n52083 , n51942 );
buf ( n52084 , n51946 );
and ( n52085 , n52083 , n52084 );
not ( n52086 , n52085 );
and ( n52087 , n52069 , n52086 );
not ( n52088 , n52087 );
xor ( n52089 , n52056 , n52068 );
xor ( n52090 , n52068 , n52069 );
not ( n52091 , n52090 );
and ( n52092 , n52089 , n52091 );
and ( n52093 , n52063 , n52092 );
and ( n52094 , n52054 , n52090 );
nor ( n52095 , n52093 , n52094 );
xnor ( n52096 , n52095 , n52072 );
and ( n52097 , n52088 , n52096 );
buf ( n52098 , n51674 );
and ( n52099 , n52098 , n52059 );
and ( n52100 , n52061 , n52057 );
nor ( n52101 , n52099 , n52100 );
not ( n52102 , n52101 );
and ( n52103 , n52096 , n52102 );
and ( n52104 , n52088 , n52102 );
or ( n52105 , n52097 , n52103 , n52104 );
and ( n52106 , n52054 , n52092 );
not ( n52107 , n52106 );
xnor ( n52108 , n52107 , n52072 );
and ( n52109 , n52105 , n52108 );
and ( n52110 , n52108 , n52065 );
and ( n52111 , n52105 , n52065 );
or ( n52112 , n52109 , n52110 , n52111 );
xor ( n52113 , n52067 , n52073 );
xor ( n52114 , n52113 , n52078 );
and ( n52115 , n52112 , n52114 );
xor ( n52116 , n52105 , n52108 );
xor ( n52117 , n52116 , n52065 );
xor ( n52118 , n52069 , n52083 );
xor ( n52119 , n52083 , n52084 );
not ( n52120 , n52119 );
and ( n52121 , n52118 , n52120 );
and ( n52122 , n52054 , n52121 );
not ( n52123 , n52122 );
xnor ( n52124 , n52123 , n52087 );
and ( n52125 , n52061 , n52092 );
and ( n52126 , n52063 , n52090 );
nor ( n52127 , n52125 , n52126 );
xnor ( n52128 , n52127 , n52072 );
and ( n52129 , n52124 , n52128 );
buf ( n52130 , n51675 );
and ( n52131 , n52130 , n52059 );
and ( n52132 , n52098 , n52057 );
nor ( n52133 , n52131 , n52132 );
and ( n52134 , n52128 , n52133 );
and ( n52135 , n52124 , n52133 );
or ( n52136 , n52129 , n52134 , n52135 );
not ( n52137 , n52133 );
buf ( n52138 , n52137 );
and ( n52139 , n52136 , n52138 );
xor ( n52140 , n52088 , n52096 );
xor ( n52141 , n52140 , n52102 );
and ( n52142 , n52138 , n52141 );
and ( n52143 , n52136 , n52141 );
or ( n52144 , n52139 , n52142 , n52143 );
and ( n52145 , n52117 , n52144 );
xor ( n52146 , n52136 , n52138 );
xor ( n52147 , n52146 , n52141 );
buf ( n52148 , n51950 );
buf ( n52149 , n51954 );
and ( n52150 , n52148 , n52149 );
not ( n52151 , n52150 );
and ( n52152 , n52084 , n52151 );
not ( n52153 , n52152 );
and ( n52154 , n52098 , n52092 );
and ( n52155 , n52061 , n52090 );
nor ( n52156 , n52154 , n52155 );
xnor ( n52157 , n52156 , n52072 );
and ( n52158 , n52153 , n52157 );
buf ( n52159 , n51676 );
and ( n52160 , n52159 , n52059 );
and ( n52161 , n52130 , n52057 );
nor ( n52162 , n52160 , n52161 );
not ( n52163 , n52162 );
and ( n52164 , n52157 , n52163 );
and ( n52165 , n52153 , n52163 );
or ( n52166 , n52158 , n52164 , n52165 );
xor ( n52167 , n52084 , n52148 );
xor ( n52168 , n52148 , n52149 );
not ( n52169 , n52168 );
and ( n52170 , n52167 , n52169 );
and ( n52171 , n52054 , n52170 );
not ( n52172 , n52171 );
xnor ( n52173 , n52172 , n52152 );
and ( n52174 , n52061 , n52121 );
and ( n52175 , n52063 , n52119 );
nor ( n52176 , n52174 , n52175 );
xnor ( n52177 , n52176 , n52087 );
and ( n52178 , n52173 , n52177 );
and ( n52179 , n52130 , n52092 );
and ( n52180 , n52098 , n52090 );
nor ( n52181 , n52179 , n52180 );
xnor ( n52182 , n52181 , n52072 );
and ( n52183 , n52177 , n52182 );
and ( n52184 , n52173 , n52182 );
or ( n52185 , n52178 , n52183 , n52184 );
buf ( n52186 , n51677 );
and ( n52187 , n52186 , n52059 );
and ( n52188 , n52159 , n52057 );
nor ( n52189 , n52187 , n52188 );
not ( n52190 , n52189 );
buf ( n52191 , n52190 );
and ( n52192 , n52185 , n52191 );
and ( n52193 , n52063 , n52121 );
and ( n52194 , n52054 , n52119 );
nor ( n52195 , n52193 , n52194 );
xnor ( n52196 , n52195 , n52087 );
and ( n52197 , n52191 , n52196 );
and ( n52198 , n52185 , n52196 );
or ( n52199 , n52192 , n52197 , n52198 );
and ( n52200 , n52166 , n52199 );
xor ( n52201 , n52124 , n52128 );
xor ( n52202 , n52201 , n52133 );
and ( n52203 , n52199 , n52202 );
and ( n52204 , n52166 , n52202 );
or ( n52205 , n52200 , n52203 , n52204 );
and ( n52206 , n52147 , n52205 );
xor ( n52207 , n52166 , n52199 );
xor ( n52208 , n52207 , n52202 );
buf ( n52209 , n51958 );
buf ( n52210 , n51962 );
and ( n52211 , n52209 , n52210 );
not ( n52212 , n52211 );
and ( n52213 , n52149 , n52212 );
not ( n52214 , n52213 );
and ( n52215 , n52063 , n52170 );
and ( n52216 , n52054 , n52168 );
nor ( n52217 , n52215 , n52216 );
xnor ( n52218 , n52217 , n52152 );
and ( n52219 , n52214 , n52218 );
buf ( n52220 , n51678 );
and ( n52221 , n52220 , n52059 );
and ( n52222 , n52186 , n52057 );
nor ( n52223 , n52221 , n52222 );
not ( n52224 , n52223 );
and ( n52225 , n52218 , n52224 );
and ( n52226 , n52214 , n52224 );
or ( n52227 , n52219 , n52225 , n52226 );
and ( n52228 , n52227 , n52189 );
xor ( n52229 , n52173 , n52177 );
xor ( n52230 , n52229 , n52182 );
and ( n52231 , n52189 , n52230 );
and ( n52232 , n52227 , n52230 );
or ( n52233 , n52228 , n52231 , n52232 );
xor ( n52234 , n52153 , n52157 );
xor ( n52235 , n52234 , n52163 );
and ( n52236 , n52233 , n52235 );
xor ( n52237 , n52185 , n52191 );
xor ( n52238 , n52237 , n52196 );
and ( n52239 , n52235 , n52238 );
and ( n52240 , n52233 , n52238 );
or ( n52241 , n52236 , n52239 , n52240 );
and ( n52242 , n52208 , n52241 );
xor ( n52243 , n52233 , n52235 );
xor ( n52244 , n52243 , n52238 );
and ( n52245 , n52061 , n52170 );
and ( n52246 , n52063 , n52168 );
nor ( n52247 , n52245 , n52246 );
xnor ( n52248 , n52247 , n52152 );
buf ( n52249 , n52248 );
and ( n52250 , n52098 , n52121 );
and ( n52251 , n52061 , n52119 );
nor ( n52252 , n52250 , n52251 );
xnor ( n52253 , n52252 , n52087 );
and ( n52254 , n52249 , n52253 );
and ( n52255 , n52159 , n52092 );
and ( n52256 , n52130 , n52090 );
nor ( n52257 , n52255 , n52256 );
xnor ( n52258 , n52257 , n52072 );
and ( n52259 , n52253 , n52258 );
and ( n52260 , n52249 , n52258 );
or ( n52261 , n52254 , n52259 , n52260 );
and ( n52262 , n52130 , n52121 );
and ( n52263 , n52098 , n52119 );
nor ( n52264 , n52262 , n52263 );
xnor ( n52265 , n52264 , n52087 );
and ( n52266 , n52186 , n52092 );
and ( n52267 , n52159 , n52090 );
nor ( n52268 , n52266 , n52267 );
xnor ( n52269 , n52268 , n52072 );
and ( n52270 , n52265 , n52269 );
buf ( n52271 , n51679 );
and ( n52272 , n52271 , n52059 );
and ( n52273 , n52220 , n52057 );
nor ( n52274 , n52272 , n52273 );
not ( n52275 , n52274 );
and ( n52276 , n52269 , n52275 );
and ( n52277 , n52265 , n52275 );
or ( n52278 , n52270 , n52276 , n52277 );
xor ( n52279 , n52214 , n52218 );
xor ( n52280 , n52279 , n52224 );
and ( n52281 , n52278 , n52280 );
xor ( n52282 , n52249 , n52253 );
xor ( n52283 , n52282 , n52258 );
and ( n52284 , n52280 , n52283 );
and ( n52285 , n52278 , n52283 );
or ( n52286 , n52281 , n52284 , n52285 );
and ( n52287 , n52261 , n52286 );
xor ( n52288 , n52227 , n52189 );
xor ( n52289 , n52288 , n52230 );
and ( n52290 , n52286 , n52289 );
and ( n52291 , n52261 , n52289 );
or ( n52292 , n52287 , n52290 , n52291 );
and ( n52293 , n52244 , n52292 );
xor ( n52294 , n52261 , n52286 );
xor ( n52295 , n52294 , n52289 );
buf ( n52296 , n51966 );
buf ( n52297 , n51970 );
and ( n52298 , n52296 , n52297 );
not ( n52299 , n52298 );
and ( n52300 , n52210 , n52299 );
not ( n52301 , n52300 );
and ( n52302 , n52098 , n52170 );
and ( n52303 , n52061 , n52168 );
nor ( n52304 , n52302 , n52303 );
xnor ( n52305 , n52304 , n52152 );
and ( n52306 , n52301 , n52305 );
buf ( n52307 , n51680 );
and ( n52308 , n52307 , n52059 );
and ( n52309 , n52271 , n52057 );
nor ( n52310 , n52308 , n52309 );
not ( n52311 , n52310 );
and ( n52312 , n52305 , n52311 );
and ( n52313 , n52301 , n52311 );
or ( n52314 , n52306 , n52312 , n52313 );
xor ( n52315 , n52149 , n52209 );
xor ( n52316 , n52209 , n52210 );
not ( n52317 , n52316 );
and ( n52318 , n52315 , n52317 );
and ( n52319 , n52054 , n52318 );
not ( n52320 , n52319 );
xnor ( n52321 , n52320 , n52213 );
and ( n52322 , n52314 , n52321 );
not ( n52323 , n52248 );
and ( n52324 , n52321 , n52323 );
and ( n52325 , n52314 , n52323 );
or ( n52326 , n52322 , n52324 , n52325 );
and ( n52327 , n52063 , n52318 );
and ( n52328 , n52054 , n52316 );
nor ( n52329 , n52327 , n52328 );
xnor ( n52330 , n52329 , n52213 );
and ( n52331 , n52159 , n52121 );
and ( n52332 , n52130 , n52119 );
nor ( n52333 , n52331 , n52332 );
xnor ( n52334 , n52333 , n52087 );
and ( n52335 , n52330 , n52334 );
and ( n52336 , n52220 , n52092 );
and ( n52337 , n52186 , n52090 );
nor ( n52338 , n52336 , n52337 );
xnor ( n52339 , n52338 , n52072 );
and ( n52340 , n52334 , n52339 );
and ( n52341 , n52330 , n52339 );
or ( n52342 , n52335 , n52340 , n52341 );
xor ( n52343 , n52210 , n52296 );
xor ( n52344 , n52296 , n52297 );
not ( n52345 , n52344 );
and ( n52346 , n52343 , n52345 );
and ( n52347 , n52054 , n52346 );
not ( n52348 , n52347 );
xnor ( n52349 , n52348 , n52300 );
and ( n52350 , n52061 , n52318 );
and ( n52351 , n52063 , n52316 );
nor ( n52352 , n52350 , n52351 );
xnor ( n52353 , n52352 , n52213 );
and ( n52354 , n52349 , n52353 );
and ( n52355 , n52186 , n52121 );
and ( n52356 , n52159 , n52119 );
nor ( n52357 , n52355 , n52356 );
xnor ( n52358 , n52357 , n52087 );
and ( n52359 , n52353 , n52358 );
and ( n52360 , n52349 , n52358 );
or ( n52361 , n52354 , n52359 , n52360 );
and ( n52362 , n52130 , n52170 );
and ( n52363 , n52098 , n52168 );
nor ( n52364 , n52362 , n52363 );
xnor ( n52365 , n52364 , n52152 );
and ( n52366 , n52271 , n52092 );
and ( n52367 , n52220 , n52090 );
nor ( n52368 , n52366 , n52367 );
xnor ( n52369 , n52368 , n52072 );
and ( n52370 , n52365 , n52369 );
buf ( n52371 , n51681 );
and ( n52372 , n52371 , n52059 );
and ( n52373 , n52307 , n52057 );
nor ( n52374 , n52372 , n52373 );
and ( n52375 , n52369 , n52374 );
and ( n52376 , n52365 , n52374 );
or ( n52377 , n52370 , n52375 , n52376 );
and ( n52378 , n52361 , n52377 );
not ( n52379 , n52374 );
buf ( n52380 , n52379 );
and ( n52381 , n52377 , n52380 );
and ( n52382 , n52361 , n52380 );
or ( n52383 , n52378 , n52381 , n52382 );
and ( n52384 , n52342 , n52383 );
xor ( n52385 , n52265 , n52269 );
xor ( n52386 , n52385 , n52275 );
and ( n52387 , n52383 , n52386 );
and ( n52388 , n52342 , n52386 );
or ( n52389 , n52384 , n52387 , n52388 );
and ( n52390 , n52326 , n52389 );
xor ( n52391 , n52278 , n52280 );
xor ( n52392 , n52391 , n52283 );
and ( n52393 , n52389 , n52392 );
and ( n52394 , n52326 , n52392 );
or ( n52395 , n52390 , n52393 , n52394 );
and ( n52396 , n52295 , n52395 );
xor ( n52397 , n52301 , n52305 );
xor ( n52398 , n52397 , n52311 );
xor ( n52399 , n52330 , n52334 );
xor ( n52400 , n52399 , n52339 );
and ( n52401 , n52398 , n52400 );
xor ( n52402 , n52361 , n52377 );
xor ( n52403 , n52402 , n52380 );
and ( n52404 , n52400 , n52403 );
and ( n52405 , n52398 , n52403 );
or ( n52406 , n52401 , n52404 , n52405 );
xor ( n52407 , n52314 , n52321 );
xor ( n52408 , n52407 , n52323 );
and ( n52409 , n52406 , n52408 );
xor ( n52410 , n52342 , n52383 );
xor ( n52411 , n52410 , n52386 );
and ( n52412 , n52408 , n52411 );
and ( n52413 , n52406 , n52411 );
or ( n52414 , n52409 , n52412 , n52413 );
xor ( n52415 , n52326 , n52389 );
xor ( n52416 , n52415 , n52392 );
and ( n52417 , n52414 , n52416 );
xor ( n52418 , n52406 , n52408 );
xor ( n52419 , n52418 , n52411 );
buf ( n52420 , n51974 );
buf ( n52421 , n51978 );
and ( n52422 , n52420 , n52421 );
not ( n52423 , n52422 );
and ( n52424 , n52297 , n52423 );
not ( n52425 , n52424 );
and ( n52426 , n52307 , n52092 );
and ( n52427 , n52271 , n52090 );
nor ( n52428 , n52426 , n52427 );
xnor ( n52429 , n52428 , n52072 );
and ( n52430 , n52425 , n52429 );
buf ( n52431 , n51682 );
and ( n52432 , n52431 , n52059 );
and ( n52433 , n52371 , n52057 );
nor ( n52434 , n52432 , n52433 );
not ( n52435 , n52434 );
and ( n52436 , n52429 , n52435 );
and ( n52437 , n52425 , n52435 );
or ( n52438 , n52430 , n52436 , n52437 );
buf ( n52439 , n51683 );
and ( n52440 , n52439 , n52059 );
and ( n52441 , n52431 , n52057 );
nor ( n52442 , n52440 , n52441 );
not ( n52443 , n52442 );
buf ( n52444 , n52443 );
and ( n52445 , n52063 , n52346 );
and ( n52446 , n52054 , n52344 );
nor ( n52447 , n52445 , n52446 );
xnor ( n52448 , n52447 , n52300 );
and ( n52449 , n52444 , n52448 );
and ( n52450 , n52220 , n52121 );
and ( n52451 , n52186 , n52119 );
nor ( n52452 , n52450 , n52451 );
xnor ( n52453 , n52452 , n52087 );
and ( n52454 , n52448 , n52453 );
and ( n52455 , n52444 , n52453 );
or ( n52456 , n52449 , n52454 , n52455 );
and ( n52457 , n52438 , n52456 );
xor ( n52458 , n52349 , n52353 );
xor ( n52459 , n52458 , n52358 );
and ( n52460 , n52456 , n52459 );
and ( n52461 , n52438 , n52459 );
or ( n52462 , n52457 , n52460 , n52461 );
and ( n52463 , n52098 , n52318 );
and ( n52464 , n52061 , n52316 );
nor ( n52465 , n52463 , n52464 );
xnor ( n52466 , n52465 , n52213 );
and ( n52467 , n52159 , n52170 );
and ( n52468 , n52130 , n52168 );
nor ( n52469 , n52467 , n52468 );
xnor ( n52470 , n52469 , n52152 );
and ( n52471 , n52466 , n52470 );
xor ( n52472 , n52425 , n52429 );
xor ( n52473 , n52472 , n52435 );
and ( n52474 , n52470 , n52473 );
and ( n52475 , n52466 , n52473 );
or ( n52476 , n52471 , n52474 , n52475 );
xor ( n52477 , n52365 , n52369 );
xor ( n52478 , n52477 , n52374 );
and ( n52479 , n52476 , n52478 );
xor ( n52480 , n52438 , n52456 );
xor ( n52481 , n52480 , n52459 );
and ( n52482 , n52478 , n52481 );
and ( n52483 , n52476 , n52481 );
or ( n52484 , n52479 , n52482 , n52483 );
and ( n52485 , n52462 , n52484 );
xor ( n52486 , n52398 , n52400 );
xor ( n52487 , n52486 , n52403 );
and ( n52488 , n52484 , n52487 );
and ( n52489 , n52462 , n52487 );
or ( n52490 , n52485 , n52488 , n52489 );
and ( n52491 , n52419 , n52490 );
xor ( n52492 , n52462 , n52484 );
xor ( n52493 , n52492 , n52487 );
and ( n52494 , n52061 , n52346 );
and ( n52495 , n52063 , n52344 );
nor ( n52496 , n52494 , n52495 );
xnor ( n52497 , n52496 , n52300 );
and ( n52498 , n52271 , n52121 );
and ( n52499 , n52220 , n52119 );
nor ( n52500 , n52498 , n52499 );
xnor ( n52501 , n52500 , n52087 );
and ( n52502 , n52497 , n52501 );
and ( n52503 , n52186 , n52170 );
and ( n52504 , n52159 , n52168 );
nor ( n52505 , n52503 , n52504 );
xnor ( n52506 , n52505 , n52152 );
and ( n52507 , n52371 , n52092 );
and ( n52508 , n52307 , n52090 );
nor ( n52509 , n52507 , n52508 );
xnor ( n52510 , n52509 , n52072 );
xor ( n52511 , n52506 , n52510 );
xor ( n52512 , n52511 , n52442 );
and ( n52513 , n52501 , n52512 );
and ( n52514 , n52497 , n52512 );
or ( n52515 , n52502 , n52513 , n52514 );
and ( n52516 , n52098 , n52346 );
and ( n52517 , n52061 , n52344 );
nor ( n52518 , n52516 , n52517 );
xnor ( n52519 , n52518 , n52300 );
and ( n52520 , n52159 , n52318 );
and ( n52521 , n52130 , n52316 );
nor ( n52522 , n52520 , n52521 );
xnor ( n52523 , n52522 , n52213 );
and ( n52524 , n52519 , n52523 );
and ( n52525 , n52220 , n52170 );
and ( n52526 , n52186 , n52168 );
nor ( n52527 , n52525 , n52526 );
xnor ( n52528 , n52527 , n52152 );
and ( n52529 , n52523 , n52528 );
and ( n52530 , n52519 , n52528 );
or ( n52531 , n52524 , n52529 , n52530 );
and ( n52532 , n52439 , n52092 );
and ( n52533 , n52431 , n52090 );
nor ( n52534 , n52532 , n52533 );
xnor ( n52535 , n52534 , n52072 );
buf ( n52536 , n52535 );
xor ( n52537 , n52297 , n52420 );
xor ( n52538 , n52420 , n52421 );
not ( n52539 , n52538 );
and ( n52540 , n52537 , n52539 );
and ( n52541 , n52063 , n52540 );
and ( n52542 , n52054 , n52538 );
nor ( n52543 , n52541 , n52542 );
xnor ( n52544 , n52543 , n52424 );
and ( n52545 , n52536 , n52544 );
and ( n52546 , n52307 , n52121 );
and ( n52547 , n52271 , n52119 );
nor ( n52548 , n52546 , n52547 );
xnor ( n52549 , n52548 , n52087 );
and ( n52550 , n52544 , n52549 );
and ( n52551 , n52536 , n52549 );
or ( n52552 , n52545 , n52550 , n52551 );
and ( n52553 , n52531 , n52552 );
buf ( n52554 , n51982 );
buf ( n52555 , n51986 );
and ( n52556 , n52554 , n52555 );
not ( n52557 , n52556 );
and ( n52558 , n52421 , n52557 );
not ( n52559 , n52558 );
and ( n52560 , n52431 , n52092 );
and ( n52561 , n52371 , n52090 );
nor ( n52562 , n52560 , n52561 );
xnor ( n52563 , n52562 , n52072 );
and ( n52564 , n52559 , n52563 );
buf ( n52565 , n51684 );
and ( n52566 , n52565 , n52059 );
and ( n52567 , n52439 , n52057 );
nor ( n52568 , n52566 , n52567 );
not ( n52569 , n52568 );
and ( n52570 , n52563 , n52569 );
and ( n52571 , n52559 , n52569 );
or ( n52572 , n52564 , n52570 , n52571 );
and ( n52573 , n52054 , n52540 );
not ( n52574 , n52573 );
xnor ( n52575 , n52574 , n52424 );
xor ( n52576 , n52572 , n52575 );
and ( n52577 , n52130 , n52318 );
and ( n52578 , n52098 , n52316 );
nor ( n52579 , n52577 , n52578 );
xnor ( n52580 , n52579 , n52213 );
xor ( n52581 , n52576 , n52580 );
and ( n52582 , n52552 , n52581 );
and ( n52583 , n52531 , n52581 );
or ( n52584 , n52553 , n52582 , n52583 );
and ( n52585 , n52515 , n52584 );
xor ( n52586 , n52444 , n52448 );
xor ( n52587 , n52586 , n52453 );
and ( n52588 , n52584 , n52587 );
and ( n52589 , n52515 , n52587 );
or ( n52590 , n52585 , n52588 , n52589 );
and ( n52591 , n52572 , n52575 );
and ( n52592 , n52575 , n52580 );
and ( n52593 , n52572 , n52580 );
or ( n52594 , n52591 , n52592 , n52593 );
and ( n52595 , n52506 , n52510 );
and ( n52596 , n52510 , n52442 );
and ( n52597 , n52506 , n52442 );
or ( n52598 , n52595 , n52596 , n52597 );
and ( n52599 , n52594 , n52598 );
xor ( n52600 , n52466 , n52470 );
xor ( n52601 , n52600 , n52473 );
and ( n52602 , n52598 , n52601 );
and ( n52603 , n52594 , n52601 );
or ( n52604 , n52599 , n52602 , n52603 );
and ( n52605 , n52590 , n52604 );
xor ( n52606 , n52476 , n52478 );
xor ( n52607 , n52606 , n52481 );
and ( n52608 , n52604 , n52607 );
and ( n52609 , n52590 , n52607 );
or ( n52610 , n52605 , n52608 , n52609 );
and ( n52611 , n52493 , n52610 );
xor ( n52612 , n52590 , n52604 );
xor ( n52613 , n52612 , n52607 );
xor ( n52614 , n52421 , n52554 );
xor ( n52615 , n52554 , n52555 );
not ( n52616 , n52615 );
and ( n52617 , n52614 , n52616 );
and ( n52618 , n52054 , n52617 );
not ( n52619 , n52618 );
xnor ( n52620 , n52619 , n52558 );
and ( n52621 , n52061 , n52540 );
and ( n52622 , n52063 , n52538 );
nor ( n52623 , n52621 , n52622 );
xnor ( n52624 , n52623 , n52424 );
and ( n52625 , n52620 , n52624 );
and ( n52626 , n52271 , n52170 );
and ( n52627 , n52220 , n52168 );
nor ( n52628 , n52626 , n52627 );
xnor ( n52629 , n52628 , n52152 );
and ( n52630 , n52624 , n52629 );
and ( n52631 , n52620 , n52629 );
or ( n52632 , n52625 , n52630 , n52631 );
and ( n52633 , n52371 , n52121 );
and ( n52634 , n52307 , n52119 );
nor ( n52635 , n52633 , n52634 );
xnor ( n52636 , n52635 , n52087 );
not ( n52637 , n52535 );
and ( n52638 , n52636 , n52637 );
buf ( n52639 , n51685 );
and ( n52640 , n52639 , n52059 );
and ( n52641 , n52565 , n52057 );
nor ( n52642 , n52640 , n52641 );
not ( n52643 , n52642 );
and ( n52644 , n52637 , n52643 );
and ( n52645 , n52636 , n52643 );
or ( n52646 , n52638 , n52644 , n52645 );
and ( n52647 , n52632 , n52646 );
xor ( n52648 , n52559 , n52563 );
xor ( n52649 , n52648 , n52569 );
and ( n52650 , n52646 , n52649 );
and ( n52651 , n52632 , n52649 );
or ( n52652 , n52647 , n52650 , n52651 );
buf ( n52653 , n51990 );
buf ( n52654 , n51994 );
and ( n52655 , n52653 , n52654 );
not ( n52656 , n52655 );
and ( n52657 , n52555 , n52656 );
not ( n52658 , n52657 );
and ( n52659 , n52565 , n52092 );
and ( n52660 , n52439 , n52090 );
nor ( n52661 , n52659 , n52660 );
xnor ( n52662 , n52661 , n52072 );
and ( n52663 , n52658 , n52662 );
buf ( n52664 , n51686 );
and ( n52665 , n52664 , n52059 );
and ( n52666 , n52639 , n52057 );
nor ( n52667 , n52665 , n52666 );
not ( n52668 , n52667 );
and ( n52669 , n52662 , n52668 );
and ( n52670 , n52658 , n52668 );
or ( n52671 , n52663 , n52669 , n52670 );
and ( n52672 , n52130 , n52346 );
and ( n52673 , n52098 , n52344 );
nor ( n52674 , n52672 , n52673 );
xnor ( n52675 , n52674 , n52300 );
and ( n52676 , n52671 , n52675 );
and ( n52677 , n52186 , n52318 );
and ( n52678 , n52159 , n52316 );
nor ( n52679 , n52677 , n52678 );
xnor ( n52680 , n52679 , n52213 );
and ( n52681 , n52675 , n52680 );
and ( n52682 , n52671 , n52680 );
or ( n52683 , n52676 , n52681 , n52682 );
xor ( n52684 , n52519 , n52523 );
xor ( n52685 , n52684 , n52528 );
and ( n52686 , n52683 , n52685 );
xor ( n52687 , n52536 , n52544 );
xor ( n52688 , n52687 , n52549 );
and ( n52689 , n52685 , n52688 );
and ( n52690 , n52683 , n52688 );
or ( n52691 , n52686 , n52689 , n52690 );
and ( n52692 , n52652 , n52691 );
xor ( n52693 , n52497 , n52501 );
xor ( n52694 , n52693 , n52512 );
and ( n52695 , n52691 , n52694 );
and ( n52696 , n52652 , n52694 );
or ( n52697 , n52692 , n52695 , n52696 );
xor ( n52698 , n52515 , n52584 );
xor ( n52699 , n52698 , n52587 );
and ( n52700 , n52697 , n52699 );
xor ( n52701 , n52594 , n52598 );
xor ( n52702 , n52701 , n52601 );
and ( n52703 , n52699 , n52702 );
and ( n52704 , n52697 , n52702 );
or ( n52705 , n52700 , n52703 , n52704 );
and ( n52706 , n52613 , n52705 );
xor ( n52707 , n52697 , n52699 );
xor ( n52708 , n52707 , n52702 );
and ( n52709 , n52371 , n52170 );
and ( n52710 , n52307 , n52168 );
nor ( n52711 , n52709 , n52710 );
xnor ( n52712 , n52711 , n52152 );
and ( n52713 , n52639 , n52092 );
and ( n52714 , n52565 , n52090 );
nor ( n52715 , n52713 , n52714 );
xnor ( n52716 , n52715 , n52072 );
and ( n52717 , n52712 , n52716 );
buf ( n52718 , n51687 );
and ( n52719 , n52718 , n52059 );
and ( n52720 , n52664 , n52057 );
nor ( n52721 , n52719 , n52720 );
not ( n52722 , n52721 );
and ( n52723 , n52716 , n52722 );
and ( n52724 , n52712 , n52722 );
or ( n52725 , n52717 , n52723 , n52724 );
and ( n52726 , n52098 , n52540 );
and ( n52727 , n52061 , n52538 );
nor ( n52728 , n52726 , n52727 );
xnor ( n52729 , n52728 , n52424 );
and ( n52730 , n52725 , n52729 );
xor ( n52731 , n52658 , n52662 );
xor ( n52732 , n52731 , n52668 );
and ( n52733 , n52729 , n52732 );
and ( n52734 , n52725 , n52732 );
or ( n52735 , n52730 , n52733 , n52734 );
xor ( n52736 , n52620 , n52624 );
xor ( n52737 , n52736 , n52629 );
and ( n52738 , n52735 , n52737 );
xor ( n52739 , n52671 , n52675 );
xor ( n52740 , n52739 , n52680 );
and ( n52741 , n52737 , n52740 );
and ( n52742 , n52735 , n52740 );
or ( n52743 , n52738 , n52741 , n52742 );
and ( n52744 , n52063 , n52617 );
and ( n52745 , n52054 , n52615 );
nor ( n52746 , n52744 , n52745 );
xnor ( n52747 , n52746 , n52558 );
and ( n52748 , n52159 , n52346 );
and ( n52749 , n52130 , n52344 );
nor ( n52750 , n52748 , n52749 );
xnor ( n52751 , n52750 , n52300 );
and ( n52752 , n52747 , n52751 );
and ( n52753 , n52220 , n52318 );
and ( n52754 , n52186 , n52316 );
nor ( n52755 , n52753 , n52754 );
xnor ( n52756 , n52755 , n52213 );
and ( n52757 , n52751 , n52756 );
and ( n52758 , n52747 , n52756 );
or ( n52759 , n52752 , n52757 , n52758 );
and ( n52760 , n52439 , n52121 );
and ( n52761 , n52431 , n52119 );
nor ( n52762 , n52760 , n52761 );
xnor ( n52763 , n52762 , n52087 );
buf ( n52764 , n52763 );
and ( n52765 , n52307 , n52170 );
and ( n52766 , n52271 , n52168 );
nor ( n52767 , n52765 , n52766 );
xnor ( n52768 , n52767 , n52152 );
and ( n52769 , n52764 , n52768 );
and ( n52770 , n52431 , n52121 );
and ( n52771 , n52371 , n52119 );
nor ( n52772 , n52770 , n52771 );
xnor ( n52773 , n52772 , n52087 );
and ( n52774 , n52768 , n52773 );
and ( n52775 , n52764 , n52773 );
or ( n52776 , n52769 , n52774 , n52775 );
and ( n52777 , n52759 , n52776 );
xor ( n52778 , n52636 , n52637 );
xor ( n52779 , n52778 , n52643 );
and ( n52780 , n52776 , n52779 );
and ( n52781 , n52759 , n52779 );
or ( n52782 , n52777 , n52780 , n52781 );
and ( n52783 , n52743 , n52782 );
xor ( n52784 , n52632 , n52646 );
xor ( n52785 , n52784 , n52649 );
and ( n52786 , n52782 , n52785 );
and ( n52787 , n52743 , n52785 );
or ( n52788 , n52783 , n52786 , n52787 );
xor ( n52789 , n52531 , n52552 );
xor ( n52790 , n52789 , n52581 );
and ( n52791 , n52788 , n52790 );
xor ( n52792 , n52652 , n52691 );
xor ( n52793 , n52792 , n52694 );
and ( n52794 , n52790 , n52793 );
and ( n52795 , n52788 , n52793 );
or ( n52796 , n52791 , n52794 , n52795 );
and ( n52797 , n52708 , n52796 );
xor ( n52798 , n52788 , n52790 );
xor ( n52799 , n52798 , n52793 );
and ( n52800 , n52431 , n52170 );
and ( n52801 , n52371 , n52168 );
nor ( n52802 , n52800 , n52801 );
xnor ( n52803 , n52802 , n52152 );
and ( n52804 , n52664 , n52092 );
and ( n52805 , n52639 , n52090 );
nor ( n52806 , n52804 , n52805 );
xnor ( n52807 , n52806 , n52072 );
and ( n52808 , n52803 , n52807 );
buf ( n52809 , n51688 );
and ( n52810 , n52809 , n52059 );
and ( n52811 , n52718 , n52057 );
nor ( n52812 , n52810 , n52811 );
not ( n52813 , n52812 );
and ( n52814 , n52807 , n52813 );
and ( n52815 , n52803 , n52813 );
or ( n52816 , n52808 , n52814 , n52815 );
and ( n52817 , n52061 , n52617 );
and ( n52818 , n52063 , n52615 );
nor ( n52819 , n52817 , n52818 );
xnor ( n52820 , n52819 , n52558 );
and ( n52821 , n52816 , n52820 );
and ( n52822 , n52130 , n52540 );
and ( n52823 , n52098 , n52538 );
nor ( n52824 , n52822 , n52823 );
xnor ( n52825 , n52824 , n52424 );
and ( n52826 , n52820 , n52825 );
and ( n52827 , n52816 , n52825 );
or ( n52828 , n52821 , n52826 , n52827 );
buf ( n52829 , n51689 );
and ( n52830 , n52829 , n52059 );
and ( n52831 , n52809 , n52057 );
nor ( n52832 , n52830 , n52831 );
not ( n52833 , n52832 );
buf ( n52834 , n52833 );
buf ( n52835 , n51998 );
buf ( n52836 , n52002 );
and ( n52837 , n52835 , n52836 );
not ( n52838 , n52837 );
and ( n52839 , n52654 , n52838 );
not ( n52840 , n52839 );
and ( n52841 , n52834 , n52840 );
and ( n52842 , n52565 , n52121 );
and ( n52843 , n52439 , n52119 );
nor ( n52844 , n52842 , n52843 );
xnor ( n52845 , n52844 , n52087 );
and ( n52846 , n52840 , n52845 );
and ( n52847 , n52834 , n52845 );
or ( n52848 , n52841 , n52846 , n52847 );
and ( n52849 , n52271 , n52318 );
and ( n52850 , n52220 , n52316 );
nor ( n52851 , n52849 , n52850 );
xnor ( n52852 , n52851 , n52213 );
and ( n52853 , n52848 , n52852 );
not ( n52854 , n52763 );
and ( n52855 , n52852 , n52854 );
and ( n52856 , n52848 , n52854 );
or ( n52857 , n52853 , n52855 , n52856 );
and ( n52858 , n52828 , n52857 );
xor ( n52859 , n52764 , n52768 );
xor ( n52860 , n52859 , n52773 );
and ( n52861 , n52857 , n52860 );
and ( n52862 , n52828 , n52860 );
or ( n52863 , n52858 , n52861 , n52862 );
xor ( n52864 , n52735 , n52737 );
xor ( n52865 , n52864 , n52740 );
and ( n52866 , n52863 , n52865 );
xor ( n52867 , n52759 , n52776 );
xor ( n52868 , n52867 , n52779 );
and ( n52869 , n52865 , n52868 );
and ( n52870 , n52863 , n52868 );
or ( n52871 , n52866 , n52869 , n52870 );
xor ( n52872 , n52683 , n52685 );
xor ( n52873 , n52872 , n52688 );
and ( n52874 , n52871 , n52873 );
xor ( n52875 , n52743 , n52782 );
xor ( n52876 , n52875 , n52785 );
and ( n52877 , n52873 , n52876 );
and ( n52878 , n52871 , n52876 );
or ( n52879 , n52874 , n52877 , n52878 );
and ( n52880 , n52799 , n52879 );
xor ( n52881 , n52871 , n52873 );
xor ( n52882 , n52881 , n52876 );
xor ( n52883 , n52555 , n52653 );
xor ( n52884 , n52653 , n52654 );
not ( n52885 , n52884 );
and ( n52886 , n52883 , n52885 );
and ( n52887 , n52054 , n52886 );
not ( n52888 , n52887 );
xnor ( n52889 , n52888 , n52657 );
and ( n52890 , n52186 , n52346 );
and ( n52891 , n52159 , n52344 );
nor ( n52892 , n52890 , n52891 );
xnor ( n52893 , n52892 , n52300 );
and ( n52894 , n52889 , n52893 );
xor ( n52895 , n52712 , n52716 );
xor ( n52896 , n52895 , n52722 );
and ( n52897 , n52893 , n52896 );
and ( n52898 , n52889 , n52896 );
or ( n52899 , n52894 , n52897 , n52898 );
xor ( n52900 , n52747 , n52751 );
xor ( n52901 , n52900 , n52756 );
and ( n52902 , n52899 , n52901 );
xor ( n52903 , n52725 , n52729 );
xor ( n52904 , n52903 , n52732 );
and ( n52905 , n52901 , n52904 );
and ( n52906 , n52899 , n52904 );
or ( n52907 , n52902 , n52905 , n52906 );
and ( n52908 , n52098 , n52617 );
and ( n52909 , n52061 , n52615 );
nor ( n52910 , n52908 , n52909 );
xnor ( n52911 , n52910 , n52558 );
and ( n52912 , n52220 , n52346 );
and ( n52913 , n52186 , n52344 );
nor ( n52914 , n52912 , n52913 );
xnor ( n52915 , n52914 , n52300 );
and ( n52916 , n52911 , n52915 );
and ( n52917 , n52307 , n52318 );
and ( n52918 , n52271 , n52316 );
nor ( n52919 , n52917 , n52918 );
xnor ( n52920 , n52919 , n52213 );
and ( n52921 , n52915 , n52920 );
and ( n52922 , n52911 , n52920 );
or ( n52923 , n52916 , n52921 , n52922 );
and ( n52924 , n52639 , n52121 );
and ( n52925 , n52565 , n52119 );
nor ( n52926 , n52924 , n52925 );
xnor ( n52927 , n52926 , n52087 );
and ( n52928 , n52718 , n52092 );
and ( n52929 , n52664 , n52090 );
nor ( n52930 , n52928 , n52929 );
xnor ( n52931 , n52930 , n52072 );
and ( n52932 , n52927 , n52931 );
and ( n52933 , n52931 , n52832 );
and ( n52934 , n52927 , n52832 );
or ( n52935 , n52932 , n52933 , n52934 );
and ( n52936 , n52159 , n52540 );
and ( n52937 , n52130 , n52538 );
nor ( n52938 , n52936 , n52937 );
xnor ( n52939 , n52938 , n52424 );
and ( n52940 , n52935 , n52939 );
xor ( n52941 , n52834 , n52840 );
xor ( n52942 , n52941 , n52845 );
and ( n52943 , n52939 , n52942 );
and ( n52944 , n52935 , n52942 );
or ( n52945 , n52940 , n52943 , n52944 );
and ( n52946 , n52923 , n52945 );
xor ( n52947 , n52848 , n52852 );
xor ( n52948 , n52947 , n52854 );
and ( n52949 , n52945 , n52948 );
and ( n52950 , n52923 , n52948 );
or ( n52951 , n52946 , n52949 , n52950 );
buf ( n52952 , n51691 );
and ( n52953 , n52952 , n52059 );
buf ( n52954 , n51690 );
and ( n52955 , n52954 , n52057 );
nor ( n52956 , n52953 , n52955 );
not ( n52957 , n52956 );
buf ( n52958 , n52957 );
buf ( n52959 , n52006 );
buf ( n52960 , n52010 );
and ( n52961 , n52959 , n52960 );
not ( n52962 , n52961 );
and ( n52963 , n52836 , n52962 );
not ( n52964 , n52963 );
and ( n52965 , n52958 , n52964 );
and ( n52966 , n52954 , n52059 );
and ( n52967 , n52829 , n52057 );
nor ( n52968 , n52966 , n52967 );
not ( n52969 , n52968 );
and ( n52970 , n52964 , n52969 );
and ( n52971 , n52958 , n52969 );
or ( n52972 , n52965 , n52970 , n52971 );
and ( n52973 , n52371 , n52318 );
and ( n52974 , n52307 , n52316 );
nor ( n52975 , n52973 , n52974 );
xnor ( n52976 , n52975 , n52213 );
and ( n52977 , n52972 , n52976 );
and ( n52978 , n52439 , n52170 );
and ( n52979 , n52431 , n52168 );
nor ( n52980 , n52978 , n52979 );
xnor ( n52981 , n52980 , n52152 );
and ( n52982 , n52976 , n52981 );
and ( n52983 , n52972 , n52981 );
or ( n52984 , n52977 , n52982 , n52983 );
and ( n52985 , n52063 , n52886 );
and ( n52986 , n52054 , n52884 );
nor ( n52987 , n52985 , n52986 );
xnor ( n52988 , n52987 , n52657 );
and ( n52989 , n52984 , n52988 );
xor ( n52990 , n52803 , n52807 );
xor ( n52991 , n52990 , n52813 );
and ( n52992 , n52988 , n52991 );
and ( n52993 , n52984 , n52991 );
or ( n52994 , n52989 , n52992 , n52993 );
xor ( n52995 , n52816 , n52820 );
xor ( n52996 , n52995 , n52825 );
and ( n52997 , n52994 , n52996 );
xor ( n52998 , n52889 , n52893 );
xor ( n52999 , n52998 , n52896 );
and ( n53000 , n52996 , n52999 );
and ( n53001 , n52994 , n52999 );
or ( n53002 , n52997 , n53000 , n53001 );
and ( n53003 , n52951 , n53002 );
xor ( n53004 , n52828 , n52857 );
xor ( n53005 , n53004 , n52860 );
and ( n53006 , n53002 , n53005 );
and ( n53007 , n52951 , n53005 );
or ( n53008 , n53003 , n53006 , n53007 );
and ( n53009 , n52907 , n53008 );
xor ( n53010 , n52863 , n52865 );
xor ( n53011 , n53010 , n52868 );
and ( n53012 , n53008 , n53011 );
and ( n53013 , n52907 , n53011 );
or ( n53014 , n53009 , n53012 , n53013 );
and ( n53015 , n52882 , n53014 );
xor ( n53016 , n52907 , n53008 );
xor ( n53017 , n53016 , n53011 );
xor ( n53018 , n52654 , n52835 );
xor ( n53019 , n52835 , n52836 );
not ( n53020 , n53019 );
and ( n53021 , n53018 , n53020 );
and ( n53022 , n52054 , n53021 );
not ( n53023 , n53022 );
xnor ( n53024 , n53023 , n52839 );
and ( n53025 , n52186 , n52540 );
and ( n53026 , n52159 , n52538 );
nor ( n53027 , n53025 , n53026 );
xnor ( n53028 , n53027 , n52424 );
and ( n53029 , n53024 , n53028 );
and ( n53030 , n52271 , n52346 );
and ( n53031 , n52220 , n52344 );
nor ( n53032 , n53030 , n53031 );
xnor ( n53033 , n53032 , n52300 );
and ( n53034 , n53028 , n53033 );
and ( n53035 , n53024 , n53033 );
or ( n53036 , n53029 , n53034 , n53035 );
and ( n53037 , n52565 , n52170 );
and ( n53038 , n52439 , n52168 );
nor ( n53039 , n53037 , n53038 );
xnor ( n53040 , n53039 , n52152 );
and ( n53041 , n52664 , n52121 );
and ( n53042 , n52639 , n52119 );
nor ( n53043 , n53041 , n53042 );
xnor ( n53044 , n53043 , n52087 );
and ( n53045 , n53040 , n53044 );
and ( n53046 , n52809 , n52092 );
and ( n53047 , n52718 , n52090 );
nor ( n53048 , n53046 , n53047 );
xnor ( n53049 , n53048 , n52072 );
and ( n53050 , n53044 , n53049 );
and ( n53051 , n53040 , n53049 );
or ( n53052 , n53045 , n53050 , n53051 );
and ( n53053 , n52061 , n52886 );
and ( n53054 , n52063 , n52884 );
nor ( n53055 , n53053 , n53054 );
xnor ( n53056 , n53055 , n52657 );
and ( n53057 , n53052 , n53056 );
and ( n53058 , n52130 , n52617 );
and ( n53059 , n52098 , n52615 );
nor ( n53060 , n53058 , n53059 );
xnor ( n53061 , n53060 , n52558 );
and ( n53062 , n53056 , n53061 );
and ( n53063 , n53052 , n53061 );
or ( n53064 , n53057 , n53062 , n53063 );
and ( n53065 , n53036 , n53064 );
xor ( n53066 , n52911 , n52915 );
xor ( n53067 , n53066 , n52920 );
and ( n53068 , n53064 , n53067 );
and ( n53069 , n53036 , n53067 );
or ( n53070 , n53065 , n53068 , n53069 );
xor ( n53071 , n52923 , n52945 );
xor ( n53072 , n53071 , n52948 );
and ( n53073 , n53070 , n53072 );
xor ( n53074 , n52994 , n52996 );
xor ( n53075 , n53074 , n52999 );
and ( n53076 , n53072 , n53075 );
and ( n53077 , n53070 , n53075 );
or ( n53078 , n53073 , n53076 , n53077 );
xor ( n53079 , n52899 , n52901 );
xor ( n53080 , n53079 , n52904 );
and ( n53081 , n53078 , n53080 );
xor ( n53082 , n52951 , n53002 );
xor ( n53083 , n53082 , n53005 );
and ( n53084 , n53080 , n53083 );
and ( n53085 , n53078 , n53083 );
or ( n53086 , n53081 , n53084 , n53085 );
and ( n53087 , n53017 , n53086 );
xor ( n53088 , n53078 , n53080 );
xor ( n53089 , n53088 , n53083 );
and ( n53090 , n52307 , n52346 );
and ( n53091 , n52271 , n52344 );
nor ( n53092 , n53090 , n53091 );
xnor ( n53093 , n53092 , n52300 );
and ( n53094 , n52431 , n52318 );
and ( n53095 , n52371 , n52316 );
nor ( n53096 , n53094 , n53095 );
xnor ( n53097 , n53096 , n52213 );
and ( n53098 , n53093 , n53097 );
xor ( n53099 , n52958 , n52964 );
xor ( n53100 , n53099 , n52969 );
and ( n53101 , n53097 , n53100 );
and ( n53102 , n53093 , n53100 );
or ( n53103 , n53098 , n53101 , n53102 );
xor ( n53104 , n52972 , n52976 );
xor ( n53105 , n53104 , n52981 );
and ( n53106 , n53103 , n53105 );
xor ( n53107 , n52927 , n52931 );
xor ( n53108 , n53107 , n52832 );
and ( n53109 , n53105 , n53108 );
and ( n53110 , n53103 , n53108 );
or ( n53111 , n53106 , n53109 , n53110 );
xor ( n53112 , n52935 , n52939 );
xor ( n53113 , n53112 , n52942 );
and ( n53114 , n53111 , n53113 );
xor ( n53115 , n52984 , n52988 );
xor ( n53116 , n53115 , n52991 );
and ( n53117 , n53113 , n53116 );
and ( n53118 , n53111 , n53116 );
or ( n53119 , n53114 , n53117 , n53118 );
and ( n53120 , n52439 , n52318 );
and ( n53121 , n52431 , n52316 );
nor ( n53122 , n53120 , n53121 );
xnor ( n53123 , n53122 , n52213 );
and ( n53124 , n52639 , n52170 );
and ( n53125 , n52565 , n52168 );
nor ( n53126 , n53124 , n53125 );
xnor ( n53127 , n53126 , n52152 );
and ( n53128 , n53123 , n53127 );
and ( n53129 , n52718 , n52121 );
and ( n53130 , n52664 , n52119 );
nor ( n53131 , n53129 , n53130 );
xnor ( n53132 , n53131 , n52087 );
and ( n53133 , n53127 , n53132 );
and ( n53134 , n53123 , n53132 );
or ( n53135 , n53128 , n53133 , n53134 );
and ( n53136 , n52098 , n52886 );
and ( n53137 , n52061 , n52884 );
nor ( n53138 , n53136 , n53137 );
xnor ( n53139 , n53138 , n52657 );
and ( n53140 , n53135 , n53139 );
and ( n53141 , n52159 , n52617 );
and ( n53142 , n52130 , n52615 );
nor ( n53143 , n53141 , n53142 );
xnor ( n53144 , n53143 , n52558 );
and ( n53145 , n53139 , n53144 );
and ( n53146 , n53135 , n53144 );
or ( n53147 , n53140 , n53145 , n53146 );
buf ( n53148 , n51693 );
and ( n53149 , n53148 , n52059 );
buf ( n53150 , n51692 );
and ( n53151 , n53150 , n52057 );
nor ( n53152 , n53149 , n53151 );
not ( n53153 , n53152 );
buf ( n53154 , n53153 );
buf ( n53155 , n52014 );
buf ( n53156 , n52018 );
and ( n53157 , n53155 , n53156 );
not ( n53158 , n53157 );
and ( n53159 , n52960 , n53158 );
not ( n53160 , n53159 );
and ( n53161 , n53154 , n53160 );
and ( n53162 , n53150 , n52059 );
and ( n53163 , n52952 , n52057 );
nor ( n53164 , n53162 , n53163 );
not ( n53165 , n53164 );
and ( n53166 , n53160 , n53165 );
and ( n53167 , n53154 , n53165 );
or ( n53168 , n53161 , n53166 , n53167 );
and ( n53169 , n52829 , n52092 );
and ( n53170 , n52809 , n52090 );
nor ( n53171 , n53169 , n53170 );
xnor ( n53172 , n53171 , n52072 );
and ( n53173 , n53168 , n53172 );
and ( n53174 , n53172 , n52956 );
and ( n53175 , n53168 , n52956 );
or ( n53176 , n53173 , n53174 , n53175 );
and ( n53177 , n52063 , n53021 );
and ( n53178 , n52054 , n53019 );
nor ( n53179 , n53177 , n53178 );
xnor ( n53180 , n53179 , n52839 );
and ( n53181 , n53176 , n53180 );
and ( n53182 , n52220 , n52540 );
and ( n53183 , n52186 , n52538 );
nor ( n53184 , n53182 , n53183 );
xnor ( n53185 , n53184 , n52424 );
and ( n53186 , n53180 , n53185 );
and ( n53187 , n53176 , n53185 );
or ( n53188 , n53181 , n53186 , n53187 );
and ( n53189 , n53147 , n53188 );
xor ( n53190 , n53052 , n53056 );
xor ( n53191 , n53190 , n53061 );
and ( n53192 , n53188 , n53191 );
and ( n53193 , n53147 , n53191 );
or ( n53194 , n53189 , n53192 , n53193 );
and ( n53195 , n52829 , n52121 );
and ( n53196 , n52809 , n52119 );
nor ( n53197 , n53195 , n53196 );
xnor ( n53198 , n53197 , n52087 );
and ( n53199 , n52952 , n52092 );
and ( n53200 , n52954 , n52090 );
nor ( n53201 , n53199 , n53200 );
xnor ( n53202 , n53201 , n52072 );
and ( n53203 , n53198 , n53202 );
and ( n53204 , n53202 , n53152 );
and ( n53205 , n53198 , n53152 );
or ( n53206 , n53203 , n53204 , n53205 );
and ( n53207 , n52954 , n52092 );
and ( n53208 , n52829 , n52090 );
nor ( n53209 , n53207 , n53208 );
xnor ( n53210 , n53209 , n52072 );
and ( n53211 , n53206 , n53210 );
xor ( n53212 , n53154 , n53160 );
xor ( n53213 , n53212 , n53165 );
and ( n53214 , n53210 , n53213 );
and ( n53215 , n53206 , n53213 );
or ( n53216 , n53211 , n53214 , n53215 );
and ( n53217 , n52371 , n52346 );
and ( n53218 , n52307 , n52344 );
nor ( n53219 , n53217 , n53218 );
xnor ( n53220 , n53219 , n52300 );
and ( n53221 , n53216 , n53220 );
xor ( n53222 , n53168 , n53172 );
xor ( n53223 , n53222 , n52956 );
and ( n53224 , n53220 , n53223 );
and ( n53225 , n53216 , n53223 );
or ( n53226 , n53221 , n53224 , n53225 );
xor ( n53227 , n53040 , n53044 );
xor ( n53228 , n53227 , n53049 );
and ( n53229 , n53226 , n53228 );
xor ( n53230 , n53093 , n53097 );
xor ( n53231 , n53230 , n53100 );
and ( n53232 , n53228 , n53231 );
and ( n53233 , n53226 , n53231 );
or ( n53234 , n53229 , n53232 , n53233 );
xor ( n53235 , n53024 , n53028 );
xor ( n53236 , n53235 , n53033 );
and ( n53237 , n53234 , n53236 );
xor ( n53238 , n53103 , n53105 );
xor ( n53239 , n53238 , n53108 );
and ( n53240 , n53236 , n53239 );
and ( n53241 , n53234 , n53239 );
or ( n53242 , n53237 , n53240 , n53241 );
and ( n53243 , n53194 , n53242 );
xor ( n53244 , n53036 , n53064 );
xor ( n53245 , n53244 , n53067 );
and ( n53246 , n53242 , n53245 );
and ( n53247 , n53194 , n53245 );
or ( n53248 , n53243 , n53246 , n53247 );
and ( n53249 , n53119 , n53248 );
xor ( n53250 , n53070 , n53072 );
xor ( n53251 , n53250 , n53075 );
and ( n53252 , n53248 , n53251 );
and ( n53253 , n53119 , n53251 );
or ( n53254 , n53249 , n53252 , n53253 );
and ( n53255 , n53089 , n53254 );
xor ( n53256 , n53119 , n53248 );
xor ( n53257 , n53256 , n53251 );
and ( n53258 , n52130 , n52886 );
and ( n53259 , n52098 , n52884 );
nor ( n53260 , n53258 , n53259 );
xnor ( n53261 , n53260 , n52657 );
and ( n53262 , n52186 , n52617 );
and ( n53263 , n52159 , n52615 );
nor ( n53264 , n53262 , n53263 );
xnor ( n53265 , n53264 , n52558 );
and ( n53266 , n53261 , n53265 );
and ( n53267 , n52271 , n52540 );
and ( n53268 , n52220 , n52538 );
nor ( n53269 , n53267 , n53268 );
xnor ( n53270 , n53269 , n52424 );
and ( n53271 , n53265 , n53270 );
and ( n53272 , n53261 , n53270 );
or ( n53273 , n53266 , n53271 , n53272 );
and ( n53274 , n52431 , n52346 );
and ( n53275 , n52371 , n52344 );
nor ( n53276 , n53274 , n53275 );
xnor ( n53277 , n53276 , n52300 );
and ( n53278 , n52565 , n52318 );
and ( n53279 , n52439 , n52316 );
nor ( n53280 , n53278 , n53279 );
xnor ( n53281 , n53280 , n52213 );
and ( n53282 , n53277 , n53281 );
and ( n53283 , n52809 , n52121 );
and ( n53284 , n52718 , n52119 );
nor ( n53285 , n53283 , n53284 );
xnor ( n53286 , n53285 , n52087 );
and ( n53287 , n53281 , n53286 );
and ( n53288 , n53277 , n53286 );
or ( n53289 , n53282 , n53287 , n53288 );
xor ( n53290 , n52836 , n52959 );
xor ( n53291 , n52959 , n52960 );
not ( n53292 , n53291 );
and ( n53293 , n53290 , n53292 );
and ( n53294 , n52054 , n53293 );
not ( n53295 , n53294 );
xnor ( n53296 , n53295 , n52963 );
and ( n53297 , n53289 , n53296 );
and ( n53298 , n52061 , n53021 );
and ( n53299 , n52063 , n53019 );
nor ( n53300 , n53298 , n53299 );
xnor ( n53301 , n53300 , n52839 );
and ( n53302 , n53296 , n53301 );
and ( n53303 , n53289 , n53301 );
or ( n53304 , n53297 , n53302 , n53303 );
and ( n53305 , n53273 , n53304 );
xor ( n53306 , n53176 , n53180 );
xor ( n53307 , n53306 , n53185 );
and ( n53308 , n53304 , n53307 );
and ( n53309 , n53273 , n53307 );
or ( n53310 , n53305 , n53308 , n53309 );
buf ( n53311 , n52022 );
buf ( n53312 , n52026 );
and ( n53313 , n53311 , n53312 );
not ( n53314 , n53313 );
and ( n53315 , n53156 , n53314 );
not ( n53316 , n53315 );
and ( n53317 , n53150 , n52092 );
and ( n53318 , n52952 , n52090 );
nor ( n53319 , n53317 , n53318 );
xnor ( n53320 , n53319 , n52072 );
and ( n53321 , n53316 , n53320 );
buf ( n53322 , n51694 );
and ( n53323 , n53322 , n52059 );
and ( n53324 , n53148 , n52057 );
nor ( n53325 , n53323 , n53324 );
not ( n53326 , n53325 );
and ( n53327 , n53320 , n53326 );
and ( n53328 , n53316 , n53326 );
or ( n53329 , n53321 , n53327 , n53328 );
and ( n53330 , n52718 , n52170 );
and ( n53331 , n52664 , n52168 );
nor ( n53332 , n53330 , n53331 );
xnor ( n53333 , n53332 , n52152 );
and ( n53334 , n53329 , n53333 );
xor ( n53335 , n53198 , n53202 );
xor ( n53336 , n53335 , n53152 );
and ( n53337 , n53333 , n53336 );
and ( n53338 , n53329 , n53336 );
or ( n53339 , n53334 , n53337 , n53338 );
and ( n53340 , n52063 , n53293 );
and ( n53341 , n52054 , n53291 );
nor ( n53342 , n53340 , n53341 );
xnor ( n53343 , n53342 , n52963 );
and ( n53344 , n53339 , n53343 );
and ( n53345 , n52220 , n52617 );
and ( n53346 , n52186 , n52615 );
nor ( n53347 , n53345 , n53346 );
xnor ( n53348 , n53347 , n52558 );
and ( n53349 , n53343 , n53348 );
and ( n53350 , n53339 , n53348 );
or ( n53351 , n53344 , n53349 , n53350 );
and ( n53352 , n52307 , n52540 );
and ( n53353 , n52271 , n52538 );
nor ( n53354 , n53352 , n53353 );
xnor ( n53355 , n53354 , n52424 );
and ( n53356 , n52664 , n52170 );
and ( n53357 , n52639 , n52168 );
nor ( n53358 , n53356 , n53357 );
xnor ( n53359 , n53358 , n52152 );
and ( n53360 , n53355 , n53359 );
xor ( n53361 , n53206 , n53210 );
xor ( n53362 , n53361 , n53213 );
and ( n53363 , n53359 , n53362 );
and ( n53364 , n53355 , n53362 );
or ( n53365 , n53360 , n53363 , n53364 );
and ( n53366 , n53351 , n53365 );
xor ( n53367 , n53123 , n53127 );
xor ( n53368 , n53367 , n53132 );
and ( n53369 , n53365 , n53368 );
and ( n53370 , n53351 , n53368 );
or ( n53371 , n53366 , n53369 , n53370 );
xor ( n53372 , n53135 , n53139 );
xor ( n53373 , n53372 , n53144 );
and ( n53374 , n53371 , n53373 );
xor ( n53375 , n53226 , n53228 );
xor ( n53376 , n53375 , n53231 );
and ( n53377 , n53373 , n53376 );
and ( n53378 , n53371 , n53376 );
or ( n53379 , n53374 , n53377 , n53378 );
and ( n53380 , n53310 , n53379 );
xor ( n53381 , n53147 , n53188 );
xor ( n53382 , n53381 , n53191 );
and ( n53383 , n53379 , n53382 );
and ( n53384 , n53310 , n53382 );
or ( n53385 , n53380 , n53383 , n53384 );
xor ( n53386 , n53111 , n53113 );
xor ( n53387 , n53386 , n53116 );
and ( n53388 , n53385 , n53387 );
xor ( n53389 , n53194 , n53242 );
xor ( n53390 , n53389 , n53245 );
and ( n53391 , n53387 , n53390 );
and ( n53392 , n53385 , n53390 );
or ( n53393 , n53388 , n53391 , n53392 );
and ( n53394 , n53257 , n53393 );
xor ( n53395 , n53385 , n53387 );
xor ( n53396 , n53395 , n53390 );
and ( n53397 , n52371 , n52540 );
and ( n53398 , n52307 , n52538 );
nor ( n53399 , n53397 , n53398 );
xnor ( n53400 , n53399 , n52424 );
and ( n53401 , n52439 , n52346 );
and ( n53402 , n52431 , n52344 );
nor ( n53403 , n53401 , n53402 );
xnor ( n53404 , n53403 , n52300 );
and ( n53405 , n53400 , n53404 );
and ( n53406 , n52639 , n52318 );
and ( n53407 , n52565 , n52316 );
nor ( n53408 , n53406 , n53407 );
xnor ( n53409 , n53408 , n52213 );
and ( n53410 , n53404 , n53409 );
and ( n53411 , n53400 , n53409 );
or ( n53412 , n53405 , n53410 , n53411 );
and ( n53413 , n52098 , n53021 );
and ( n53414 , n52061 , n53019 );
nor ( n53415 , n53413 , n53414 );
xnor ( n53416 , n53415 , n52839 );
and ( n53417 , n53412 , n53416 );
and ( n53418 , n52159 , n52886 );
and ( n53419 , n52130 , n52884 );
nor ( n53420 , n53418 , n53419 );
xnor ( n53421 , n53420 , n52657 );
and ( n53422 , n53416 , n53421 );
and ( n53423 , n53412 , n53421 );
or ( n53424 , n53417 , n53422 , n53423 );
xor ( n53425 , n53261 , n53265 );
xor ( n53426 , n53425 , n53270 );
and ( n53427 , n53424 , n53426 );
xor ( n53428 , n53216 , n53220 );
xor ( n53429 , n53428 , n53223 );
and ( n53430 , n53426 , n53429 );
and ( n53431 , n53424 , n53429 );
or ( n53432 , n53427 , n53430 , n53431 );
xor ( n53433 , n53273 , n53304 );
xor ( n53434 , n53433 , n53307 );
and ( n53435 , n53432 , n53434 );
xor ( n53436 , n53371 , n53373 );
xor ( n53437 , n53436 , n53376 );
and ( n53438 , n53434 , n53437 );
and ( n53439 , n53432 , n53437 );
or ( n53440 , n53435 , n53438 , n53439 );
xor ( n53441 , n53234 , n53236 );
xor ( n53442 , n53441 , n53239 );
and ( n53443 , n53440 , n53442 );
xor ( n53444 , n53310 , n53379 );
xor ( n53445 , n53444 , n53382 );
and ( n53446 , n53442 , n53445 );
and ( n53447 , n53440 , n53445 );
or ( n53448 , n53443 , n53446 , n53447 );
and ( n53449 , n53396 , n53448 );
xor ( n53450 , n53440 , n53442 );
xor ( n53451 , n53450 , n53445 );
xor ( n53452 , n52960 , n53155 );
xor ( n53453 , n53155 , n53156 );
not ( n53454 , n53453 );
and ( n53455 , n53452 , n53454 );
and ( n53456 , n52054 , n53455 );
not ( n53457 , n53456 );
xnor ( n53458 , n53457 , n53159 );
and ( n53459 , n52130 , n53021 );
and ( n53460 , n52098 , n53019 );
nor ( n53461 , n53459 , n53460 );
xnor ( n53462 , n53461 , n52839 );
and ( n53463 , n53458 , n53462 );
and ( n53464 , n52271 , n52617 );
and ( n53465 , n52220 , n52615 );
nor ( n53466 , n53464 , n53465 );
xnor ( n53467 , n53466 , n52558 );
and ( n53468 , n53462 , n53467 );
and ( n53469 , n53458 , n53467 );
or ( n53470 , n53463 , n53468 , n53469 );
and ( n53471 , n52829 , n52170 );
and ( n53472 , n52809 , n52168 );
nor ( n53473 , n53471 , n53472 );
xnor ( n53474 , n53473 , n52152 );
and ( n53475 , n52952 , n52121 );
and ( n53476 , n52954 , n52119 );
nor ( n53477 , n53475 , n53476 );
xnor ( n53478 , n53477 , n52087 );
and ( n53479 , n53474 , n53478 );
and ( n53480 , n53148 , n52092 );
and ( n53481 , n53150 , n52090 );
nor ( n53482 , n53480 , n53481 );
xnor ( n53483 , n53482 , n52072 );
and ( n53484 , n53478 , n53483 );
and ( n53485 , n53474 , n53483 );
or ( n53486 , n53479 , n53484 , n53485 );
and ( n53487 , n52664 , n52318 );
and ( n53488 , n52639 , n52316 );
nor ( n53489 , n53487 , n53488 );
xnor ( n53490 , n53489 , n52213 );
and ( n53491 , n53486 , n53490 );
and ( n53492 , n52809 , n52170 );
and ( n53493 , n52718 , n52168 );
nor ( n53494 , n53492 , n53493 );
xnor ( n53495 , n53494 , n52152 );
and ( n53496 , n53490 , n53495 );
and ( n53497 , n53486 , n53495 );
or ( n53498 , n53491 , n53496 , n53497 );
buf ( n53499 , n51695 );
and ( n53500 , n53499 , n52059 );
and ( n53501 , n53322 , n52057 );
nor ( n53502 , n53500 , n53501 );
not ( n53503 , n53502 );
buf ( n53504 , n53503 );
and ( n53505 , n52954 , n52121 );
and ( n53506 , n52829 , n52119 );
nor ( n53507 , n53505 , n53506 );
xnor ( n53508 , n53507 , n52087 );
and ( n53509 , n53504 , n53508 );
xor ( n53510 , n53316 , n53320 );
xor ( n53511 , n53510 , n53326 );
and ( n53512 , n53508 , n53511 );
and ( n53513 , n53504 , n53511 );
or ( n53514 , n53509 , n53512 , n53513 );
and ( n53515 , n53498 , n53514 );
and ( n53516 , n52186 , n52886 );
and ( n53517 , n52159 , n52884 );
nor ( n53518 , n53516 , n53517 );
xnor ( n53519 , n53518 , n52657 );
and ( n53520 , n53514 , n53519 );
and ( n53521 , n53498 , n53519 );
or ( n53522 , n53515 , n53520 , n53521 );
and ( n53523 , n53470 , n53522 );
xor ( n53524 , n53277 , n53281 );
xor ( n53525 , n53524 , n53286 );
and ( n53526 , n53522 , n53525 );
and ( n53527 , n53470 , n53525 );
or ( n53528 , n53523 , n53526 , n53527 );
xor ( n53529 , n53412 , n53416 );
xor ( n53530 , n53529 , n53421 );
xor ( n53531 , n53339 , n53343 );
xor ( n53532 , n53531 , n53348 );
and ( n53533 , n53530 , n53532 );
xor ( n53534 , n53355 , n53359 );
xor ( n53535 , n53534 , n53362 );
and ( n53536 , n53532 , n53535 );
and ( n53537 , n53530 , n53535 );
or ( n53538 , n53533 , n53536 , n53537 );
and ( n53539 , n53528 , n53538 );
xor ( n53540 , n53289 , n53296 );
xor ( n53541 , n53540 , n53301 );
and ( n53542 , n53538 , n53541 );
and ( n53543 , n53528 , n53541 );
or ( n53544 , n53539 , n53542 , n53543 );
xor ( n53545 , n53351 , n53365 );
xor ( n53546 , n53545 , n53368 );
xor ( n53547 , n53528 , n53538 );
xor ( n53548 , n53547 , n53541 );
and ( n53549 , n53546 , n53548 );
xor ( n53550 , n53424 , n53426 );
xor ( n53551 , n53550 , n53429 );
and ( n53552 , n53548 , n53551 );
and ( n53553 , n53546 , n53551 );
or ( n53554 , n53549 , n53552 , n53553 );
and ( n53555 , n53544 , n53554 );
xor ( n53556 , n53432 , n53434 );
xor ( n53557 , n53556 , n53437 );
and ( n53558 , n53554 , n53557 );
and ( n53559 , n53544 , n53557 );
or ( n53560 , n53555 , n53558 , n53559 );
and ( n53561 , n53451 , n53560 );
xor ( n53562 , n53544 , n53554 );
xor ( n53563 , n53562 , n53557 );
and ( n53564 , n52431 , n52540 );
and ( n53565 , n52371 , n52538 );
nor ( n53566 , n53564 , n53565 );
xnor ( n53567 , n53566 , n52424 );
and ( n53568 , n52565 , n52346 );
and ( n53569 , n52439 , n52344 );
nor ( n53570 , n53568 , n53569 );
xnor ( n53571 , n53570 , n52300 );
and ( n53572 , n53567 , n53571 );
xor ( n53573 , n53504 , n53508 );
xor ( n53574 , n53573 , n53511 );
and ( n53575 , n53571 , n53574 );
and ( n53576 , n53567 , n53574 );
or ( n53577 , n53572 , n53575 , n53576 );
and ( n53578 , n52061 , n53293 );
and ( n53579 , n52063 , n53291 );
nor ( n53580 , n53578 , n53579 );
xnor ( n53581 , n53580 , n52963 );
and ( n53582 , n53577 , n53581 );
xor ( n53583 , n53400 , n53404 );
xor ( n53584 , n53583 , n53409 );
and ( n53585 , n53581 , n53584 );
and ( n53586 , n53577 , n53584 );
or ( n53587 , n53582 , n53585 , n53586 );
and ( n53588 , n52220 , n52886 );
and ( n53589 , n52186 , n52884 );
nor ( n53590 , n53588 , n53589 );
xnor ( n53591 , n53590 , n52657 );
xor ( n53592 , n53486 , n53490 );
xor ( n53593 , n53592 , n53495 );
and ( n53594 , n53591 , n53593 );
xor ( n53595 , n53567 , n53571 );
xor ( n53596 , n53595 , n53574 );
and ( n53597 , n53593 , n53596 );
and ( n53598 , n53591 , n53596 );
or ( n53599 , n53594 , n53597 , n53598 );
xor ( n53600 , n53458 , n53462 );
xor ( n53601 , n53600 , n53467 );
and ( n53602 , n53599 , n53601 );
xor ( n53603 , n53498 , n53514 );
xor ( n53604 , n53603 , n53519 );
and ( n53605 , n53601 , n53604 );
and ( n53606 , n53599 , n53604 );
or ( n53607 , n53602 , n53605 , n53606 );
and ( n53608 , n53587 , n53607 );
and ( n53609 , n52439 , n52540 );
and ( n53610 , n52431 , n52538 );
nor ( n53611 , n53609 , n53610 );
xnor ( n53612 , n53611 , n52424 );
and ( n53613 , n52718 , n52318 );
and ( n53614 , n52664 , n52316 );
nor ( n53615 , n53613 , n53614 );
xnor ( n53616 , n53615 , n52213 );
and ( n53617 , n53612 , n53616 );
xor ( n53618 , n53474 , n53478 );
xor ( n53619 , n53618 , n53483 );
and ( n53620 , n53616 , n53619 );
and ( n53621 , n53612 , n53619 );
or ( n53622 , n53617 , n53620 , n53621 );
and ( n53623 , n52063 , n53455 );
and ( n53624 , n52054 , n53453 );
nor ( n53625 , n53623 , n53624 );
xnor ( n53626 , n53625 , n53159 );
and ( n53627 , n53622 , n53626 );
and ( n53628 , n52159 , n53021 );
and ( n53629 , n52130 , n53019 );
nor ( n53630 , n53628 , n53629 );
xnor ( n53631 , n53630 , n52839 );
and ( n53632 , n53626 , n53631 );
and ( n53633 , n53622 , n53631 );
or ( n53634 , n53627 , n53632 , n53633 );
and ( n53635 , n52954 , n52170 );
and ( n53636 , n52829 , n52168 );
nor ( n53637 , n53635 , n53636 );
xnor ( n53638 , n53637 , n52152 );
and ( n53639 , n53150 , n52121 );
and ( n53640 , n52952 , n52119 );
nor ( n53641 , n53639 , n53640 );
xnor ( n53642 , n53641 , n52087 );
and ( n53643 , n53638 , n53642 );
buf ( n53644 , n51696 );
and ( n53645 , n53644 , n52059 );
and ( n53646 , n53499 , n52057 );
nor ( n53647 , n53645 , n53646 );
not ( n53648 , n53647 );
and ( n53649 , n53642 , n53648 );
and ( n53650 , n53638 , n53648 );
or ( n53651 , n53643 , n53649 , n53650 );
buf ( n53652 , n51697 );
and ( n53653 , n53652 , n52059 );
and ( n53654 , n53644 , n52057 );
nor ( n53655 , n53653 , n53654 );
not ( n53656 , n53655 );
buf ( n53657 , n53656 );
buf ( n53658 , n52030 );
buf ( n53659 , n52034 );
and ( n53660 , n53658 , n53659 );
not ( n53661 , n53660 );
and ( n53662 , n53312 , n53661 );
not ( n53663 , n53662 );
and ( n53664 , n53657 , n53663 );
and ( n53665 , n53322 , n52092 );
and ( n53666 , n53148 , n52090 );
nor ( n53667 , n53665 , n53666 );
xnor ( n53668 , n53667 , n52072 );
and ( n53669 , n53663 , n53668 );
and ( n53670 , n53657 , n53668 );
or ( n53671 , n53664 , n53669 , n53670 );
and ( n53672 , n53651 , n53671 );
and ( n53673 , n53671 , n53502 );
and ( n53674 , n53651 , n53502 );
or ( n53675 , n53672 , n53673 , n53674 );
and ( n53676 , n52098 , n53293 );
and ( n53677 , n52061 , n53291 );
nor ( n53678 , n53676 , n53677 );
xnor ( n53679 , n53678 , n52963 );
and ( n53680 , n53675 , n53679 );
and ( n53681 , n52307 , n52617 );
and ( n53682 , n52271 , n52615 );
nor ( n53683 , n53681 , n53682 );
xnor ( n53684 , n53683 , n52558 );
and ( n53685 , n53679 , n53684 );
and ( n53686 , n53675 , n53684 );
or ( n53687 , n53680 , n53685 , n53686 );
and ( n53688 , n53634 , n53687 );
xor ( n53689 , n53329 , n53333 );
xor ( n53690 , n53689 , n53336 );
and ( n53691 , n53687 , n53690 );
and ( n53692 , n53634 , n53690 );
or ( n53693 , n53688 , n53691 , n53692 );
and ( n53694 , n53607 , n53693 );
and ( n53695 , n53587 , n53693 );
or ( n53696 , n53608 , n53694 , n53695 );
xor ( n53697 , n53587 , n53607 );
xor ( n53698 , n53697 , n53693 );
xor ( n53699 , n53470 , n53522 );
xor ( n53700 , n53699 , n53525 );
and ( n53701 , n53698 , n53700 );
xor ( n53702 , n53530 , n53532 );
xor ( n53703 , n53702 , n53535 );
and ( n53704 , n53700 , n53703 );
and ( n53705 , n53698 , n53703 );
or ( n53706 , n53701 , n53704 , n53705 );
and ( n53707 , n53696 , n53706 );
xor ( n53708 , n53546 , n53548 );
xor ( n53709 , n53708 , n53551 );
and ( n53710 , n53706 , n53709 );
and ( n53711 , n53696 , n53709 );
or ( n53712 , n53707 , n53710 , n53711 );
and ( n53713 , n53563 , n53712 );
xor ( n53714 , n53696 , n53706 );
xor ( n53715 , n53714 , n53709 );
and ( n53716 , n53148 , n52121 );
and ( n53717 , n53150 , n52119 );
nor ( n53718 , n53716 , n53717 );
xnor ( n53719 , n53718 , n52087 );
and ( n53720 , n53499 , n52092 );
and ( n53721 , n53322 , n52090 );
nor ( n53722 , n53720 , n53721 );
xnor ( n53723 , n53722 , n52072 );
and ( n53724 , n53719 , n53723 );
and ( n53725 , n53723 , n53655 );
and ( n53726 , n53719 , n53655 );
or ( n53727 , n53724 , n53725 , n53726 );
xor ( n53728 , n53638 , n53642 );
xor ( n53729 , n53728 , n53648 );
and ( n53730 , n53727 , n53729 );
xor ( n53731 , n53657 , n53663 );
xor ( n53732 , n53731 , n53668 );
and ( n53733 , n53729 , n53732 );
and ( n53734 , n53727 , n53732 );
or ( n53735 , n53730 , n53733 , n53734 );
xor ( n53736 , n53156 , n53311 );
xor ( n53737 , n53311 , n53312 );
not ( n53738 , n53737 );
and ( n53739 , n53736 , n53738 );
and ( n53740 , n52054 , n53739 );
not ( n53741 , n53740 );
xnor ( n53742 , n53741 , n53315 );
and ( n53743 , n53735 , n53742 );
and ( n53744 , n52186 , n53021 );
and ( n53745 , n52159 , n53019 );
nor ( n53746 , n53744 , n53745 );
xnor ( n53747 , n53746 , n52839 );
and ( n53748 , n53742 , n53747 );
and ( n53749 , n53735 , n53747 );
or ( n53750 , n53743 , n53748 , n53749 );
and ( n53751 , n52307 , n52886 );
and ( n53752 , n52271 , n52884 );
nor ( n53753 , n53751 , n53752 );
xnor ( n53754 , n53753 , n52657 );
and ( n53755 , n52664 , n52346 );
and ( n53756 , n52639 , n52344 );
nor ( n53757 , n53755 , n53756 );
xnor ( n53758 , n53757 , n52300 );
and ( n53759 , n53754 , n53758 );
and ( n53760 , n52809 , n52318 );
and ( n53761 , n52718 , n52316 );
nor ( n53762 , n53760 , n53761 );
xnor ( n53763 , n53762 , n52213 );
and ( n53764 , n53758 , n53763 );
and ( n53765 , n53754 , n53763 );
or ( n53766 , n53759 , n53764 , n53765 );
and ( n53767 , n52130 , n53293 );
and ( n53768 , n52098 , n53291 );
nor ( n53769 , n53767 , n53768 );
xnor ( n53770 , n53769 , n52963 );
and ( n53771 , n53766 , n53770 );
xor ( n53772 , n53612 , n53616 );
xor ( n53773 , n53772 , n53619 );
and ( n53774 , n53770 , n53773 );
and ( n53775 , n53766 , n53773 );
or ( n53776 , n53771 , n53774 , n53775 );
and ( n53777 , n53750 , n53776 );
xor ( n53778 , n53622 , n53626 );
xor ( n53779 , n53778 , n53631 );
and ( n53780 , n53776 , n53779 );
and ( n53781 , n53750 , n53779 );
or ( n53782 , n53777 , n53780 , n53781 );
buf ( n53783 , n51699 );
and ( n53784 , n53783 , n52059 );
buf ( n53785 , n51698 );
and ( n53786 , n53785 , n52057 );
nor ( n53787 , n53784 , n53786 );
not ( n53788 , n53787 );
buf ( n53789 , n53788 );
buf ( n53790 , n52038 );
buf ( n53791 , n52042 );
and ( n53792 , n53790 , n53791 );
not ( n53793 , n53792 );
and ( n53794 , n53659 , n53793 );
not ( n53795 , n53794 );
and ( n53796 , n53789 , n53795 );
and ( n53797 , n53785 , n52059 );
and ( n53798 , n53652 , n52057 );
nor ( n53799 , n53797 , n53798 );
not ( n53800 , n53799 );
and ( n53801 , n53795 , n53800 );
and ( n53802 , n53789 , n53800 );
or ( n53803 , n53796 , n53801 , n53802 );
and ( n53804 , n52829 , n52318 );
and ( n53805 , n52809 , n52316 );
nor ( n53806 , n53804 , n53805 );
xnor ( n53807 , n53806 , n52213 );
and ( n53808 , n53803 , n53807 );
and ( n53809 , n52952 , n52170 );
and ( n53810 , n52954 , n52168 );
nor ( n53811 , n53809 , n53810 );
xnor ( n53812 , n53811 , n52152 );
and ( n53813 , n53807 , n53812 );
and ( n53814 , n53803 , n53812 );
or ( n53815 , n53808 , n53813 , n53814 );
and ( n53816 , n52431 , n52617 );
and ( n53817 , n52371 , n52615 );
nor ( n53818 , n53816 , n53817 );
xnor ( n53819 , n53818 , n52558 );
and ( n53820 , n53815 , n53819 );
and ( n53821 , n52565 , n52540 );
and ( n53822 , n52439 , n52538 );
nor ( n53823 , n53821 , n53822 );
xnor ( n53824 , n53823 , n52424 );
and ( n53825 , n53819 , n53824 );
and ( n53826 , n53815 , n53824 );
or ( n53827 , n53820 , n53825 , n53826 );
and ( n53828 , n52061 , n53455 );
and ( n53829 , n52063 , n53453 );
nor ( n53830 , n53828 , n53829 );
xnor ( n53831 , n53830 , n53159 );
and ( n53832 , n53827 , n53831 );
and ( n53833 , n52271 , n52886 );
and ( n53834 , n52220 , n52884 );
nor ( n53835 , n53833 , n53834 );
xnor ( n53836 , n53835 , n52657 );
and ( n53837 , n53831 , n53836 );
and ( n53838 , n53827 , n53836 );
or ( n53839 , n53832 , n53837 , n53838 );
and ( n53840 , n52371 , n52617 );
and ( n53841 , n52307 , n52615 );
nor ( n53842 , n53840 , n53841 );
xnor ( n53843 , n53842 , n52558 );
and ( n53844 , n52639 , n52346 );
and ( n53845 , n52565 , n52344 );
nor ( n53846 , n53844 , n53845 );
xnor ( n53847 , n53846 , n52300 );
and ( n53848 , n53843 , n53847 );
xor ( n53849 , n53651 , n53671 );
xor ( n53850 , n53849 , n53502 );
and ( n53851 , n53847 , n53850 );
and ( n53852 , n53843 , n53850 );
or ( n53853 , n53848 , n53851 , n53852 );
and ( n53854 , n53839 , n53853 );
xor ( n53855 , n53675 , n53679 );
xor ( n53856 , n53855 , n53684 );
and ( n53857 , n53853 , n53856 );
and ( n53858 , n53839 , n53856 );
or ( n53859 , n53854 , n53857 , n53858 );
and ( n53860 , n53782 , n53859 );
xor ( n53861 , n53577 , n53581 );
xor ( n53862 , n53861 , n53584 );
and ( n53863 , n53859 , n53862 );
and ( n53864 , n53782 , n53862 );
or ( n53865 , n53860 , n53863 , n53864 );
xor ( n53866 , n53599 , n53601 );
xor ( n53867 , n53866 , n53604 );
xor ( n53868 , n53634 , n53687 );
xor ( n53869 , n53868 , n53690 );
and ( n53870 , n53867 , n53869 );
xor ( n53871 , n53782 , n53859 );
xor ( n53872 , n53871 , n53862 );
and ( n53873 , n53869 , n53872 );
and ( n53874 , n53867 , n53872 );
or ( n53875 , n53870 , n53873 , n53874 );
and ( n53876 , n53865 , n53875 );
xor ( n53877 , n53698 , n53700 );
xor ( n53878 , n53877 , n53703 );
and ( n53879 , n53875 , n53878 );
and ( n53880 , n53865 , n53878 );
or ( n53881 , n53876 , n53879 , n53880 );
and ( n53882 , n53715 , n53881 );
xor ( n53883 , n53865 , n53875 );
xor ( n53884 , n53883 , n53878 );
buf ( n53885 , n52050 );
not ( n53886 , n53885 );
buf ( n53887 , n53886 );
buf ( n53888 , n53887 );
buf ( n53889 , n52046 );
and ( n53890 , n53889 , n53885 );
not ( n53891 , n53890 );
and ( n53892 , n53791 , n53891 );
not ( n53893 , n53892 );
and ( n53894 , n53888 , n53893 );
buf ( n53895 , n51700 );
and ( n53896 , n53895 , n52059 );
and ( n53897 , n53783 , n52057 );
nor ( n53898 , n53896 , n53897 );
not ( n53899 , n53898 );
and ( n53900 , n53893 , n53899 );
and ( n53901 , n53888 , n53899 );
or ( n53902 , n53894 , n53900 , n53901 );
and ( n53903 , n53148 , n52170 );
and ( n53904 , n53150 , n52168 );
nor ( n53905 , n53903 , n53904 );
xnor ( n53906 , n53905 , n52152 );
and ( n53907 , n53902 , n53906 );
and ( n53908 , n53652 , n52092 );
and ( n53909 , n53644 , n52090 );
nor ( n53910 , n53908 , n53909 );
xnor ( n53911 , n53910 , n52072 );
and ( n53912 , n53906 , n53911 );
and ( n53913 , n53902 , n53911 );
or ( n53914 , n53907 , n53912 , n53913 );
and ( n53915 , n52954 , n52318 );
and ( n53916 , n52829 , n52316 );
nor ( n53917 , n53915 , n53916 );
xnor ( n53918 , n53917 , n52213 );
and ( n53919 , n53914 , n53918 );
xor ( n53920 , n53789 , n53795 );
xor ( n53921 , n53920 , n53800 );
and ( n53922 , n53918 , n53921 );
and ( n53923 , n53914 , n53921 );
or ( n53924 , n53919 , n53922 , n53923 );
and ( n53925 , n52639 , n52540 );
and ( n53926 , n52565 , n52538 );
nor ( n53927 , n53925 , n53926 );
xnor ( n53928 , n53927 , n52424 );
and ( n53929 , n53924 , n53928 );
and ( n53930 , n52718 , n52346 );
and ( n53931 , n52664 , n52344 );
nor ( n53932 , n53930 , n53931 );
xnor ( n53933 , n53932 , n52300 );
and ( n53934 , n53928 , n53933 );
and ( n53935 , n53924 , n53933 );
or ( n53936 , n53929 , n53934 , n53935 );
xor ( n53937 , n53754 , n53758 );
xor ( n53938 , n53937 , n53763 );
and ( n53939 , n53936 , n53938 );
xor ( n53940 , n53815 , n53819 );
xor ( n53941 , n53940 , n53824 );
and ( n53942 , n53938 , n53941 );
and ( n53943 , n53936 , n53941 );
or ( n53944 , n53939 , n53942 , n53943 );
xor ( n53945 , n53735 , n53742 );
xor ( n53946 , n53945 , n53747 );
and ( n53947 , n53944 , n53946 );
xor ( n53948 , n53827 , n53831 );
xor ( n53949 , n53948 , n53836 );
and ( n53950 , n53946 , n53949 );
and ( n53951 , n53944 , n53949 );
or ( n53952 , n53947 , n53950 , n53951 );
and ( n53953 , n52130 , n53455 );
and ( n53954 , n52098 , n53453 );
nor ( n53955 , n53953 , n53954 );
xnor ( n53956 , n53955 , n53159 );
and ( n53957 , n52186 , n53293 );
and ( n53958 , n52159 , n53291 );
nor ( n53959 , n53957 , n53958 );
xnor ( n53960 , n53959 , n52963 );
and ( n53961 , n53956 , n53960 );
and ( n53962 , n52271 , n53021 );
and ( n53963 , n52220 , n53019 );
nor ( n53964 , n53962 , n53963 );
xnor ( n53965 , n53964 , n52839 );
and ( n53966 , n53960 , n53965 );
and ( n53967 , n53956 , n53965 );
or ( n53968 , n53961 , n53966 , n53967 );
xor ( n53969 , n53312 , n53658 );
xor ( n53970 , n53658 , n53659 );
not ( n53971 , n53970 );
and ( n53972 , n53969 , n53971 );
and ( n53973 , n52054 , n53972 );
not ( n53974 , n53973 );
xnor ( n53975 , n53974 , n53662 );
and ( n53976 , n52371 , n52886 );
and ( n53977 , n52307 , n52884 );
nor ( n53978 , n53976 , n53977 );
xnor ( n53979 , n53978 , n52657 );
and ( n53980 , n53975 , n53979 );
xor ( n53981 , n53803 , n53807 );
xor ( n53982 , n53981 , n53812 );
and ( n53983 , n53979 , n53982 );
and ( n53984 , n53975 , n53982 );
or ( n53985 , n53980 , n53983 , n53984 );
and ( n53986 , n53968 , n53985 );
and ( n53987 , n52431 , n52886 );
and ( n53988 , n52371 , n52884 );
nor ( n53989 , n53987 , n53988 );
xnor ( n53990 , n53989 , n52657 );
and ( n53991 , n52565 , n52617 );
and ( n53992 , n52439 , n52615 );
nor ( n53993 , n53991 , n53992 );
xnor ( n53994 , n53993 , n52558 );
and ( n53995 , n53990 , n53994 );
and ( n53996 , n52664 , n52540 );
and ( n53997 , n52639 , n52538 );
nor ( n53998 , n53996 , n53997 );
xnor ( n53999 , n53998 , n52424 );
and ( n54000 , n53994 , n53999 );
and ( n54001 , n53990 , n53999 );
or ( n54002 , n53995 , n54000 , n54001 );
and ( n54003 , n52952 , n52318 );
and ( n54004 , n52954 , n52316 );
nor ( n54005 , n54003 , n54004 );
xnor ( n54006 , n54005 , n52213 );
and ( n54007 , n53499 , n52121 );
and ( n54008 , n53322 , n52119 );
nor ( n54009 , n54007 , n54008 );
xnor ( n54010 , n54009 , n52087 );
and ( n54011 , n54006 , n54010 );
and ( n54012 , n54010 , n53787 );
and ( n54013 , n54006 , n53787 );
or ( n54014 , n54011 , n54012 , n54013 );
and ( n54015 , n52809 , n52346 );
and ( n54016 , n52718 , n52344 );
nor ( n54017 , n54015 , n54016 );
xnor ( n54018 , n54017 , n52300 );
and ( n54019 , n54014 , n54018 );
and ( n54020 , n53150 , n52170 );
and ( n54021 , n52952 , n52168 );
nor ( n54022 , n54020 , n54021 );
xnor ( n54023 , n54022 , n52152 );
and ( n54024 , n53322 , n52121 );
and ( n54025 , n53148 , n52119 );
nor ( n54026 , n54024 , n54025 );
xnor ( n54027 , n54026 , n52087 );
xor ( n54028 , n54023 , n54027 );
and ( n54029 , n53644 , n52092 );
and ( n54030 , n53499 , n52090 );
nor ( n54031 , n54029 , n54030 );
xnor ( n54032 , n54031 , n52072 );
xor ( n54033 , n54028 , n54032 );
and ( n54034 , n54018 , n54033 );
and ( n54035 , n54014 , n54033 );
or ( n54036 , n54019 , n54034 , n54035 );
and ( n54037 , n54002 , n54036 );
and ( n54038 , n54023 , n54027 );
and ( n54039 , n54027 , n54032 );
and ( n54040 , n54023 , n54032 );
or ( n54041 , n54038 , n54039 , n54040 );
and ( n54042 , n52439 , n52617 );
and ( n54043 , n52431 , n52615 );
nor ( n54044 , n54042 , n54043 );
xnor ( n54045 , n54044 , n52558 );
xor ( n54046 , n54041 , n54045 );
xor ( n54047 , n53719 , n53723 );
xor ( n54048 , n54047 , n53655 );
xor ( n54049 , n54046 , n54048 );
and ( n54050 , n54036 , n54049 );
and ( n54051 , n54002 , n54049 );
or ( n54052 , n54037 , n54050 , n54051 );
and ( n54053 , n53985 , n54052 );
and ( n54054 , n53968 , n54052 );
or ( n54055 , n53986 , n54053 , n54054 );
and ( n54056 , n53322 , n52170 );
and ( n54057 , n53148 , n52168 );
nor ( n54058 , n54056 , n54057 );
xnor ( n54059 , n54058 , n52152 );
and ( n54060 , n53644 , n52121 );
and ( n54061 , n53499 , n52119 );
nor ( n54062 , n54060 , n54061 );
xnor ( n54063 , n54062 , n52087 );
and ( n54064 , n54059 , n54063 );
and ( n54065 , n53785 , n52092 );
and ( n54066 , n53652 , n52090 );
nor ( n54067 , n54065 , n54066 );
xnor ( n54068 , n54067 , n52072 );
and ( n54069 , n54063 , n54068 );
and ( n54070 , n54059 , n54068 );
or ( n54071 , n54064 , n54069 , n54070 );
not ( n54072 , n53887 );
and ( n54073 , n53652 , n52121 );
and ( n54074 , n53644 , n52119 );
nor ( n54075 , n54073 , n54074 );
xnor ( n54076 , n54075 , n52087 );
and ( n54077 , n54072 , n54076 );
buf ( n54078 , n51701 );
and ( n54079 , n54078 , n52059 );
and ( n54080 , n53895 , n52057 );
nor ( n54081 , n54079 , n54080 );
not ( n54082 , n54081 );
and ( n54083 , n54076 , n54082 );
and ( n54084 , n54072 , n54082 );
or ( n54085 , n54077 , n54083 , n54084 );
and ( n54086 , n53150 , n52318 );
and ( n54087 , n52952 , n52316 );
nor ( n54088 , n54086 , n54087 );
xnor ( n54089 , n54088 , n52213 );
and ( n54090 , n54085 , n54089 );
xor ( n54091 , n53888 , n53893 );
xor ( n54092 , n54091 , n53899 );
and ( n54093 , n54089 , n54092 );
and ( n54094 , n54085 , n54092 );
or ( n54095 , n54090 , n54093 , n54094 );
and ( n54096 , n54071 , n54095 );
and ( n54097 , n52829 , n52346 );
and ( n54098 , n52809 , n52344 );
nor ( n54099 , n54097 , n54098 );
xnor ( n54100 , n54099 , n52300 );
and ( n54101 , n54095 , n54100 );
and ( n54102 , n54071 , n54100 );
or ( n54103 , n54096 , n54101 , n54102 );
and ( n54104 , n52307 , n53021 );
and ( n54105 , n52271 , n53019 );
nor ( n54106 , n54104 , n54105 );
xnor ( n54107 , n54106 , n52839 );
and ( n54108 , n54103 , n54107 );
xor ( n54109 , n53914 , n53918 );
xor ( n54110 , n54109 , n53921 );
and ( n54111 , n54107 , n54110 );
and ( n54112 , n54103 , n54110 );
or ( n54113 , n54108 , n54111 , n54112 );
and ( n54114 , n52061 , n53739 );
and ( n54115 , n52063 , n53737 );
nor ( n54116 , n54114 , n54115 );
xnor ( n54117 , n54116 , n53315 );
and ( n54118 , n54113 , n54117 );
xor ( n54119 , n53924 , n53928 );
xor ( n54120 , n54119 , n53933 );
and ( n54121 , n54117 , n54120 );
and ( n54122 , n54113 , n54120 );
or ( n54123 , n54118 , n54121 , n54122 );
and ( n54124 , n54041 , n54045 );
and ( n54125 , n54045 , n54048 );
and ( n54126 , n54041 , n54048 );
or ( n54127 , n54124 , n54125 , n54126 );
and ( n54128 , n52098 , n53455 );
and ( n54129 , n52061 , n53453 );
nor ( n54130 , n54128 , n54129 );
xnor ( n54131 , n54130 , n53159 );
xor ( n54132 , n54127 , n54131 );
and ( n54133 , n52159 , n53293 );
and ( n54134 , n52130 , n53291 );
nor ( n54135 , n54133 , n54134 );
xnor ( n54136 , n54135 , n52963 );
xor ( n54137 , n54132 , n54136 );
and ( n54138 , n54123 , n54137 );
and ( n54139 , n52063 , n53739 );
and ( n54140 , n52054 , n53737 );
nor ( n54141 , n54139 , n54140 );
xnor ( n54142 , n54141 , n53315 );
and ( n54143 , n52220 , n53021 );
and ( n54144 , n52186 , n53019 );
nor ( n54145 , n54143 , n54144 );
xnor ( n54146 , n54145 , n52839 );
xor ( n54147 , n54142 , n54146 );
xor ( n54148 , n53727 , n53729 );
xor ( n54149 , n54148 , n53732 );
xor ( n54150 , n54147 , n54149 );
and ( n54151 , n54137 , n54150 );
and ( n54152 , n54123 , n54150 );
or ( n54153 , n54138 , n54151 , n54152 );
and ( n54154 , n54055 , n54153 );
xor ( n54155 , n53766 , n53770 );
xor ( n54156 , n54155 , n53773 );
and ( n54157 , n54153 , n54156 );
and ( n54158 , n54055 , n54156 );
or ( n54159 , n54154 , n54157 , n54158 );
and ( n54160 , n53952 , n54159 );
xor ( n54161 , n53750 , n53776 );
xor ( n54162 , n54161 , n53779 );
and ( n54163 , n54159 , n54162 );
and ( n54164 , n53952 , n54162 );
or ( n54165 , n54160 , n54163 , n54164 );
and ( n54166 , n54127 , n54131 );
and ( n54167 , n54131 , n54136 );
and ( n54168 , n54127 , n54136 );
or ( n54169 , n54166 , n54167 , n54168 );
and ( n54170 , n54142 , n54146 );
and ( n54171 , n54146 , n54149 );
and ( n54172 , n54142 , n54149 );
or ( n54173 , n54170 , n54171 , n54172 );
and ( n54174 , n54169 , n54173 );
xor ( n54175 , n53843 , n53847 );
xor ( n54176 , n54175 , n53850 );
and ( n54177 , n54173 , n54176 );
and ( n54178 , n54169 , n54176 );
or ( n54179 , n54174 , n54177 , n54178 );
xor ( n54180 , n53839 , n53853 );
xor ( n54181 , n54180 , n53856 );
and ( n54182 , n54179 , n54181 );
xor ( n54183 , n53591 , n53593 );
xor ( n54184 , n54183 , n53596 );
and ( n54185 , n54181 , n54184 );
and ( n54186 , n54179 , n54184 );
or ( n54187 , n54182 , n54185 , n54186 );
and ( n54188 , n54165 , n54187 );
xor ( n54189 , n53867 , n53869 );
xor ( n54190 , n54189 , n53872 );
and ( n54191 , n54187 , n54190 );
and ( n54192 , n54165 , n54190 );
or ( n54193 , n54188 , n54191 , n54192 );
and ( n54194 , n53884 , n54193 );
xor ( n54195 , n54165 , n54187 );
xor ( n54196 , n54195 , n54190 );
and ( n54197 , n52718 , n52540 );
and ( n54198 , n52664 , n52538 );
nor ( n54199 , n54197 , n54198 );
xnor ( n54200 , n54199 , n52424 );
xor ( n54201 , n53902 , n53906 );
xor ( n54202 , n54201 , n53911 );
and ( n54203 , n54200 , n54202 );
xor ( n54204 , n54006 , n54010 );
xor ( n54205 , n54204 , n53787 );
and ( n54206 , n54202 , n54205 );
and ( n54207 , n54200 , n54205 );
or ( n54208 , n54203 , n54206 , n54207 );
and ( n54209 , n52063 , n53972 );
and ( n54210 , n52054 , n53970 );
nor ( n54211 , n54209 , n54210 );
xnor ( n54212 , n54211 , n53662 );
and ( n54213 , n54208 , n54212 );
and ( n54214 , n52159 , n53455 );
and ( n54215 , n52130 , n53453 );
nor ( n54216 , n54214 , n54215 );
xnor ( n54217 , n54216 , n53159 );
and ( n54218 , n54212 , n54217 );
and ( n54219 , n54208 , n54217 );
or ( n54220 , n54213 , n54218 , n54219 );
and ( n54221 , n52098 , n53739 );
and ( n54222 , n52061 , n53737 );
nor ( n54223 , n54221 , n54222 );
xnor ( n54224 , n54223 , n53315 );
and ( n54225 , n52220 , n53293 );
and ( n54226 , n52186 , n53291 );
nor ( n54227 , n54225 , n54226 );
xnor ( n54228 , n54227 , n52963 );
and ( n54229 , n54224 , n54228 );
xor ( n54230 , n54014 , n54018 );
xor ( n54231 , n54230 , n54033 );
and ( n54232 , n54228 , n54231 );
and ( n54233 , n54224 , n54231 );
or ( n54234 , n54229 , n54232 , n54233 );
and ( n54235 , n54220 , n54234 );
xor ( n54236 , n53975 , n53979 );
xor ( n54237 , n54236 , n53982 );
and ( n54238 , n54234 , n54237 );
and ( n54239 , n54220 , n54237 );
or ( n54240 , n54235 , n54238 , n54239 );
xor ( n54241 , n53968 , n53985 );
xor ( n54242 , n54241 , n54052 );
and ( n54243 , n54240 , n54242 );
xor ( n54244 , n53936 , n53938 );
xor ( n54245 , n54244 , n53941 );
and ( n54246 , n54242 , n54245 );
and ( n54247 , n54240 , n54245 );
or ( n54248 , n54243 , n54246 , n54247 );
xor ( n54249 , n53944 , n53946 );
xor ( n54250 , n54249 , n53949 );
and ( n54251 , n54248 , n54250 );
xor ( n54252 , n54169 , n54173 );
xor ( n54253 , n54252 , n54176 );
and ( n54254 , n54250 , n54253 );
and ( n54255 , n54248 , n54253 );
or ( n54256 , n54251 , n54254 , n54255 );
xor ( n54257 , n53952 , n54159 );
xor ( n54258 , n54257 , n54162 );
and ( n54259 , n54256 , n54258 );
xor ( n54260 , n54179 , n54181 );
xor ( n54261 , n54260 , n54184 );
and ( n54262 , n54258 , n54261 );
and ( n54263 , n54256 , n54261 );
or ( n54264 , n54259 , n54262 , n54263 );
and ( n54265 , n54196 , n54264 );
and ( n54266 , n52565 , n52886 );
and ( n54267 , n52439 , n52884 );
nor ( n54268 , n54266 , n54267 );
xnor ( n54269 , n54268 , n52657 );
and ( n54270 , n52664 , n52617 );
and ( n54271 , n52639 , n52615 );
nor ( n54272 , n54270 , n54271 );
xnor ( n54273 , n54272 , n52558 );
and ( n54274 , n54269 , n54273 );
and ( n54275 , n52809 , n52540 );
and ( n54276 , n52718 , n52538 );
nor ( n54277 , n54275 , n54276 );
xnor ( n54278 , n54277 , n52424 );
and ( n54279 , n54273 , n54278 );
and ( n54280 , n54269 , n54278 );
or ( n54281 , n54274 , n54279 , n54280 );
xor ( n54282 , n53659 , n53790 );
xor ( n54283 , n53790 , n53791 );
not ( n54284 , n54283 );
and ( n54285 , n54282 , n54284 );
and ( n54286 , n52054 , n54285 );
not ( n54287 , n54286 );
xnor ( n54288 , n54287 , n53794 );
and ( n54289 , n54281 , n54288 );
and ( n54290 , n52061 , n53972 );
and ( n54291 , n52063 , n53970 );
nor ( n54292 , n54290 , n54291 );
xnor ( n54293 , n54292 , n53662 );
and ( n54294 , n54288 , n54293 );
and ( n54295 , n54281 , n54293 );
or ( n54296 , n54289 , n54294 , n54295 );
and ( n54297 , n52829 , n52540 );
and ( n54298 , n52809 , n52538 );
nor ( n54299 , n54297 , n54298 );
xnor ( n54300 , n54299 , n52424 );
and ( n54301 , n53148 , n52318 );
and ( n54302 , n53150 , n52316 );
nor ( n54303 , n54301 , n54302 );
xnor ( n54304 , n54303 , n52213 );
and ( n54305 , n54300 , n54304 );
xor ( n54306 , n54072 , n54076 );
xor ( n54307 , n54306 , n54082 );
and ( n54308 , n54304 , n54307 );
and ( n54309 , n54300 , n54307 );
or ( n54310 , n54305 , n54308 , n54309 );
and ( n54311 , n52431 , n53021 );
and ( n54312 , n52371 , n53019 );
nor ( n54313 , n54311 , n54312 );
xnor ( n54314 , n54313 , n52839 );
and ( n54315 , n54310 , n54314 );
xor ( n54316 , n54085 , n54089 );
xor ( n54317 , n54316 , n54092 );
and ( n54318 , n54314 , n54317 );
and ( n54319 , n54310 , n54317 );
or ( n54320 , n54315 , n54318 , n54319 );
and ( n54321 , n52130 , n53739 );
and ( n54322 , n52098 , n53737 );
nor ( n54323 , n54321 , n54322 );
xnor ( n54324 , n54323 , n53315 );
and ( n54325 , n54320 , n54324 );
and ( n54326 , n52271 , n53293 );
and ( n54327 , n52220 , n53291 );
nor ( n54328 , n54326 , n54327 );
xnor ( n54329 , n54328 , n52963 );
and ( n54330 , n54324 , n54329 );
and ( n54331 , n54320 , n54329 );
or ( n54332 , n54325 , n54330 , n54331 );
and ( n54333 , n54296 , n54332 );
and ( n54334 , n52186 , n53455 );
and ( n54335 , n52159 , n53453 );
nor ( n54336 , n54334 , n54335 );
xnor ( n54337 , n54336 , n53159 );
and ( n54338 , n52371 , n53021 );
and ( n54339 , n52307 , n53019 );
nor ( n54340 , n54338 , n54339 );
xnor ( n54341 , n54340 , n52839 );
and ( n54342 , n54337 , n54341 );
xor ( n54343 , n54071 , n54095 );
xor ( n54344 , n54343 , n54100 );
and ( n54345 , n54341 , n54344 );
and ( n54346 , n54337 , n54344 );
or ( n54347 , n54342 , n54345 , n54346 );
and ( n54348 , n54332 , n54347 );
and ( n54349 , n54296 , n54347 );
or ( n54350 , n54333 , n54348 , n54349 );
xor ( n54351 , n54113 , n54117 );
xor ( n54352 , n54351 , n54120 );
and ( n54353 , n54350 , n54352 );
xor ( n54354 , n54220 , n54234 );
xor ( n54355 , n54354 , n54237 );
and ( n54356 , n54352 , n54355 );
and ( n54357 , n54350 , n54355 );
or ( n54358 , n54353 , n54356 , n54357 );
and ( n54359 , n53895 , n52092 );
and ( n54360 , n53783 , n52090 );
nor ( n54361 , n54359 , n54360 );
xnor ( n54362 , n54361 , n52072 );
and ( n54363 , n53885 , n54362 );
buf ( n54364 , n51702 );
and ( n54365 , n54364 , n52059 );
and ( n54366 , n54078 , n52057 );
nor ( n54367 , n54365 , n54366 );
not ( n54368 , n54367 );
and ( n54369 , n54362 , n54368 );
and ( n54370 , n53885 , n54368 );
or ( n54371 , n54363 , n54369 , n54370 );
and ( n54372 , n53499 , n52170 );
and ( n54373 , n53322 , n52168 );
nor ( n54374 , n54372 , n54373 );
xnor ( n54375 , n54374 , n52152 );
and ( n54376 , n54371 , n54375 );
and ( n54377 , n53783 , n52092 );
and ( n54378 , n53785 , n52090 );
nor ( n54379 , n54377 , n54378 );
xnor ( n54380 , n54379 , n52072 );
and ( n54381 , n54375 , n54380 );
and ( n54382 , n54371 , n54380 );
or ( n54383 , n54376 , n54381 , n54382 );
and ( n54384 , n52954 , n52346 );
and ( n54385 , n52829 , n52344 );
nor ( n54386 , n54384 , n54385 );
xnor ( n54387 , n54386 , n52300 );
and ( n54388 , n54383 , n54387 );
xor ( n54389 , n54059 , n54063 );
xor ( n54390 , n54389 , n54068 );
and ( n54391 , n54387 , n54390 );
and ( n54392 , n54383 , n54390 );
or ( n54393 , n54388 , n54391 , n54392 );
and ( n54394 , n52439 , n52886 );
and ( n54395 , n52431 , n52884 );
nor ( n54396 , n54394 , n54395 );
xnor ( n54397 , n54396 , n52657 );
and ( n54398 , n54393 , n54397 );
and ( n54399 , n52639 , n52617 );
and ( n54400 , n52565 , n52615 );
nor ( n54401 , n54399 , n54400 );
xnor ( n54402 , n54401 , n52558 );
and ( n54403 , n54397 , n54402 );
and ( n54404 , n54393 , n54402 );
or ( n54405 , n54398 , n54403 , n54404 );
xor ( n54406 , n53990 , n53994 );
xor ( n54407 , n54406 , n53999 );
and ( n54408 , n54405 , n54407 );
xor ( n54409 , n54103 , n54107 );
xor ( n54410 , n54409 , n54110 );
and ( n54411 , n54407 , n54410 );
and ( n54412 , n54405 , n54410 );
or ( n54413 , n54408 , n54411 , n54412 );
xor ( n54414 , n53956 , n53960 );
xor ( n54415 , n54414 , n53965 );
and ( n54416 , n54413 , n54415 );
xor ( n54417 , n54002 , n54036 );
xor ( n54418 , n54417 , n54049 );
and ( n54419 , n54415 , n54418 );
and ( n54420 , n54413 , n54418 );
or ( n54421 , n54416 , n54419 , n54420 );
and ( n54422 , n54358 , n54421 );
xor ( n54423 , n54123 , n54137 );
xor ( n54424 , n54423 , n54150 );
and ( n54425 , n54421 , n54424 );
and ( n54426 , n54358 , n54424 );
or ( n54427 , n54422 , n54425 , n54426 );
xor ( n54428 , n54248 , n54250 );
xor ( n54429 , n54428 , n54253 );
and ( n54430 , n54427 , n54429 );
xor ( n54431 , n54055 , n54153 );
xor ( n54432 , n54431 , n54156 );
and ( n54433 , n54429 , n54432 );
and ( n54434 , n54427 , n54432 );
or ( n54435 , n54430 , n54433 , n54434 );
xor ( n54436 , n54256 , n54258 );
xor ( n54437 , n54436 , n54261 );
and ( n54438 , n54435 , n54437 );
xor ( n54439 , n54427 , n54429 );
xor ( n54440 , n54439 , n54432 );
and ( n54441 , n53322 , n52318 );
and ( n54442 , n53148 , n52316 );
nor ( n54443 , n54441 , n54442 );
xnor ( n54444 , n54443 , n52213 );
and ( n54445 , n53644 , n52170 );
and ( n54446 , n53499 , n52168 );
nor ( n54447 , n54445 , n54446 );
xnor ( n54448 , n54447 , n52152 );
and ( n54449 , n54444 , n54448 );
and ( n54450 , n53785 , n52121 );
and ( n54451 , n53652 , n52119 );
nor ( n54452 , n54450 , n54451 );
xnor ( n54453 , n54452 , n52087 );
and ( n54454 , n54448 , n54453 );
and ( n54455 , n54444 , n54453 );
or ( n54456 , n54449 , n54454 , n54455 );
and ( n54457 , n53652 , n52170 );
and ( n54458 , n53644 , n52168 );
nor ( n54459 , n54457 , n54458 );
xnor ( n54460 , n54459 , n52152 );
and ( n54461 , n54078 , n52092 );
and ( n54462 , n53895 , n52090 );
nor ( n54463 , n54461 , n54462 );
xnor ( n54464 , n54463 , n52072 );
and ( n54465 , n54460 , n54464 );
buf ( n54466 , n51703 );
and ( n54467 , n54466 , n52059 );
and ( n54468 , n54364 , n52057 );
nor ( n54469 , n54467 , n54468 );
not ( n54470 , n54469 );
and ( n54471 , n54464 , n54470 );
and ( n54472 , n54460 , n54470 );
or ( n54473 , n54465 , n54471 , n54472 );
and ( n54474 , n53150 , n52346 );
and ( n54475 , n52952 , n52344 );
nor ( n54476 , n54474 , n54475 );
xnor ( n54477 , n54476 , n52300 );
and ( n54478 , n54473 , n54477 );
xor ( n54479 , n53885 , n54362 );
xor ( n54480 , n54479 , n54368 );
and ( n54481 , n54477 , n54480 );
and ( n54482 , n54473 , n54480 );
or ( n54483 , n54478 , n54481 , n54482 );
and ( n54484 , n54456 , n54483 );
and ( n54485 , n52952 , n52346 );
and ( n54486 , n52954 , n52344 );
nor ( n54487 , n54485 , n54486 );
xnor ( n54488 , n54487 , n52300 );
and ( n54489 , n54483 , n54488 );
and ( n54490 , n54456 , n54488 );
or ( n54491 , n54484 , n54489 , n54490 );
and ( n54492 , n52307 , n53293 );
and ( n54493 , n52271 , n53291 );
nor ( n54494 , n54492 , n54493 );
xnor ( n54495 , n54494 , n52963 );
and ( n54496 , n54491 , n54495 );
xor ( n54497 , n54383 , n54387 );
xor ( n54498 , n54497 , n54390 );
and ( n54499 , n54495 , n54498 );
and ( n54500 , n54491 , n54498 );
or ( n54501 , n54496 , n54499 , n54500 );
xor ( n54502 , n54393 , n54397 );
xor ( n54503 , n54502 , n54402 );
and ( n54504 , n54501 , n54503 );
xor ( n54505 , n54200 , n54202 );
xor ( n54506 , n54505 , n54205 );
and ( n54507 , n54503 , n54506 );
and ( n54508 , n54501 , n54506 );
or ( n54509 , n54504 , n54507 , n54508 );
xor ( n54510 , n54208 , n54212 );
xor ( n54511 , n54510 , n54217 );
and ( n54512 , n54509 , n54511 );
xor ( n54513 , n54224 , n54228 );
xor ( n54514 , n54513 , n54231 );
and ( n54515 , n54511 , n54514 );
and ( n54516 , n54509 , n54514 );
or ( n54517 , n54512 , n54515 , n54516 );
and ( n54518 , n52439 , n53021 );
and ( n54519 , n52431 , n53019 );
nor ( n54520 , n54518 , n54519 );
xnor ( n54521 , n54520 , n52839 );
xor ( n54522 , n54371 , n54375 );
xor ( n54523 , n54522 , n54380 );
and ( n54524 , n54521 , n54523 );
xor ( n54525 , n54300 , n54304 );
xor ( n54526 , n54525 , n54307 );
and ( n54527 , n54523 , n54526 );
and ( n54528 , n54521 , n54526 );
or ( n54529 , n54524 , n54527 , n54528 );
and ( n54530 , n52098 , n53972 );
and ( n54531 , n52061 , n53970 );
nor ( n54532 , n54530 , n54531 );
xnor ( n54533 , n54532 , n53662 );
and ( n54534 , n54529 , n54533 );
and ( n54535 , n52159 , n53739 );
and ( n54536 , n52130 , n53737 );
nor ( n54537 , n54535 , n54536 );
xnor ( n54538 , n54537 , n53315 );
and ( n54539 , n54533 , n54538 );
and ( n54540 , n54529 , n54538 );
or ( n54541 , n54534 , n54539 , n54540 );
and ( n54542 , n52063 , n54285 );
and ( n54543 , n52054 , n54283 );
nor ( n54544 , n54542 , n54543 );
xnor ( n54545 , n54544 , n53794 );
and ( n54546 , n52220 , n53455 );
and ( n54547 , n52186 , n53453 );
nor ( n54548 , n54546 , n54547 );
xnor ( n54549 , n54548 , n53159 );
and ( n54550 , n54545 , n54549 );
xor ( n54551 , n54310 , n54314 );
xor ( n54552 , n54551 , n54317 );
and ( n54553 , n54549 , n54552 );
and ( n54554 , n54545 , n54552 );
or ( n54555 , n54550 , n54553 , n54554 );
and ( n54556 , n54541 , n54555 );
xor ( n54557 , n54337 , n54341 );
xor ( n54558 , n54557 , n54344 );
and ( n54559 , n54555 , n54558 );
and ( n54560 , n54541 , n54558 );
or ( n54561 , n54556 , n54559 , n54560 );
xor ( n54562 , n54296 , n54332 );
xor ( n54563 , n54562 , n54347 );
and ( n54564 , n54561 , n54563 );
xor ( n54565 , n54405 , n54407 );
xor ( n54566 , n54565 , n54410 );
and ( n54567 , n54563 , n54566 );
and ( n54568 , n54561 , n54566 );
or ( n54569 , n54564 , n54567 , n54568 );
and ( n54570 , n54517 , n54569 );
xor ( n54571 , n54413 , n54415 );
xor ( n54572 , n54571 , n54418 );
and ( n54573 , n54569 , n54572 );
and ( n54574 , n54517 , n54572 );
or ( n54575 , n54570 , n54573 , n54574 );
xor ( n54576 , n54240 , n54242 );
xor ( n54577 , n54576 , n54245 );
and ( n54578 , n54575 , n54577 );
xor ( n54579 , n54358 , n54421 );
xor ( n54580 , n54579 , n54424 );
and ( n54581 , n54577 , n54580 );
and ( n54582 , n54575 , n54580 );
or ( n54583 , n54578 , n54581 , n54582 );
and ( n54584 , n54440 , n54583 );
xor ( n54585 , n54575 , n54577 );
xor ( n54586 , n54585 , n54580 );
and ( n54587 , n52371 , n53293 );
and ( n54588 , n52307 , n53291 );
nor ( n54589 , n54587 , n54588 );
xnor ( n54590 , n54589 , n52963 );
and ( n54591 , n52639 , n52886 );
and ( n54592 , n52565 , n52884 );
nor ( n54593 , n54591 , n54592 );
xnor ( n54594 , n54593 , n52657 );
and ( n54595 , n54590 , n54594 );
and ( n54596 , n52718 , n52617 );
and ( n54597 , n52664 , n52615 );
nor ( n54598 , n54596 , n54597 );
xnor ( n54599 , n54598 , n52558 );
and ( n54600 , n54594 , n54599 );
and ( n54601 , n54590 , n54599 );
or ( n54602 , n54595 , n54600 , n54601 );
xor ( n54603 , n54269 , n54273 );
xor ( n54604 , n54603 , n54278 );
and ( n54605 , n54602 , n54604 );
xor ( n54606 , n54491 , n54495 );
xor ( n54607 , n54606 , n54498 );
and ( n54608 , n54604 , n54607 );
and ( n54609 , n54602 , n54607 );
or ( n54610 , n54605 , n54608 , n54609 );
xor ( n54611 , n54281 , n54288 );
xor ( n54612 , n54611 , n54293 );
and ( n54613 , n54610 , n54612 );
xor ( n54614 , n54320 , n54324 );
xor ( n54615 , n54614 , n54329 );
and ( n54616 , n54612 , n54615 );
and ( n54617 , n54610 , n54615 );
or ( n54618 , n54613 , n54616 , n54617 );
xor ( n54619 , n54509 , n54511 );
xor ( n54620 , n54619 , n54514 );
and ( n54621 , n54618 , n54620 );
xor ( n54622 , n54561 , n54563 );
xor ( n54623 , n54622 , n54566 );
and ( n54624 , n54620 , n54623 );
and ( n54625 , n54618 , n54623 );
or ( n54626 , n54621 , n54624 , n54625 );
xor ( n54627 , n54350 , n54352 );
xor ( n54628 , n54627 , n54355 );
and ( n54629 , n54626 , n54628 );
xor ( n54630 , n54517 , n54569 );
xor ( n54631 , n54630 , n54572 );
and ( n54632 , n54628 , n54631 );
and ( n54633 , n54626 , n54631 );
or ( n54634 , n54629 , n54632 , n54633 );
and ( n54635 , n54586 , n54634 );
xor ( n54636 , n54626 , n54628 );
xor ( n54637 , n54636 , n54631 );
and ( n54638 , n52565 , n53021 );
and ( n54639 , n52439 , n53019 );
nor ( n54640 , n54638 , n54639 );
xnor ( n54641 , n54640 , n52839 );
and ( n54642 , n52664 , n52886 );
and ( n54643 , n52639 , n52884 );
nor ( n54644 , n54642 , n54643 );
xnor ( n54645 , n54644 , n52657 );
and ( n54646 , n54641 , n54645 );
and ( n54647 , n52809 , n52617 );
and ( n54648 , n52718 , n52615 );
nor ( n54649 , n54647 , n54648 );
xnor ( n54650 , n54649 , n52558 );
and ( n54651 , n54645 , n54650 );
and ( n54652 , n54641 , n54650 );
or ( n54653 , n54646 , n54651 , n54652 );
and ( n54654 , n52061 , n54285 );
and ( n54655 , n52063 , n54283 );
nor ( n54656 , n54654 , n54655 );
xnor ( n54657 , n54656 , n53794 );
and ( n54658 , n54653 , n54657 );
and ( n54659 , n52186 , n53739 );
and ( n54660 , n52159 , n53737 );
nor ( n54661 , n54659 , n54660 );
xnor ( n54662 , n54661 , n53315 );
and ( n54663 , n54657 , n54662 );
and ( n54664 , n54653 , n54662 );
or ( n54665 , n54658 , n54663 , n54664 );
and ( n54666 , n52829 , n52617 );
and ( n54667 , n52809 , n52615 );
nor ( n54668 , n54666 , n54667 );
xnor ( n54669 , n54668 , n52558 );
and ( n54670 , n53148 , n52346 );
and ( n54671 , n53150 , n52344 );
nor ( n54672 , n54670 , n54671 );
xnor ( n54673 , n54672 , n52300 );
and ( n54674 , n54669 , n54673 );
xor ( n54675 , n54460 , n54464 );
xor ( n54676 , n54675 , n54470 );
and ( n54677 , n54673 , n54676 );
and ( n54678 , n54669 , n54676 );
or ( n54679 , n54674 , n54677 , n54678 );
and ( n54680 , n52431 , n53293 );
and ( n54681 , n52371 , n53291 );
nor ( n54682 , n54680 , n54681 );
xnor ( n54683 , n54682 , n52963 );
and ( n54684 , n54679 , n54683 );
xor ( n54685 , n54473 , n54477 );
xor ( n54686 , n54685 , n54480 );
and ( n54687 , n54683 , n54686 );
and ( n54688 , n54679 , n54686 );
or ( n54689 , n54684 , n54687 , n54688 );
xor ( n54690 , n53791 , n53889 );
xor ( n54691 , n53889 , n53885 );
not ( n54692 , n54691 );
and ( n54693 , n54690 , n54692 );
and ( n54694 , n52054 , n54693 );
not ( n54695 , n54694 );
xnor ( n54696 , n54695 , n53892 );
and ( n54697 , n54689 , n54696 );
and ( n54698 , n52271 , n53455 );
and ( n54699 , n52220 , n53453 );
nor ( n54700 , n54698 , n54699 );
xnor ( n54701 , n54700 , n53159 );
and ( n54702 , n54696 , n54701 );
and ( n54703 , n54689 , n54701 );
or ( n54704 , n54697 , n54702 , n54703 );
and ( n54705 , n54665 , n54704 );
and ( n54706 , n53895 , n52121 );
and ( n54707 , n53783 , n52119 );
nor ( n54708 , n54706 , n54707 );
xnor ( n54709 , n54708 , n52087 );
and ( n54710 , n54364 , n52092 );
and ( n54711 , n54078 , n52090 );
nor ( n54712 , n54710 , n54711 );
xnor ( n54713 , n54712 , n52072 );
and ( n54714 , n54709 , n54713 );
buf ( n54715 , n51704 );
and ( n54716 , n54715 , n52059 );
and ( n54717 , n54466 , n52057 );
nor ( n54718 , n54716 , n54717 );
not ( n54719 , n54718 );
and ( n54720 , n54713 , n54719 );
and ( n54721 , n54709 , n54719 );
or ( n54722 , n54714 , n54720 , n54721 );
and ( n54723 , n53499 , n52318 );
and ( n54724 , n53322 , n52316 );
nor ( n54725 , n54723 , n54724 );
xnor ( n54726 , n54725 , n52213 );
and ( n54727 , n54722 , n54726 );
and ( n54728 , n53783 , n52121 );
and ( n54729 , n53785 , n52119 );
nor ( n54730 , n54728 , n54729 );
xnor ( n54731 , n54730 , n52087 );
and ( n54732 , n54726 , n54731 );
and ( n54733 , n54722 , n54731 );
or ( n54734 , n54727 , n54732 , n54733 );
and ( n54735 , n52954 , n52540 );
and ( n54736 , n52829 , n52538 );
nor ( n54737 , n54735 , n54736 );
xnor ( n54738 , n54737 , n52424 );
and ( n54739 , n54734 , n54738 );
xor ( n54740 , n54444 , n54448 );
xor ( n54741 , n54740 , n54453 );
and ( n54742 , n54738 , n54741 );
and ( n54743 , n54734 , n54741 );
or ( n54744 , n54739 , n54742 , n54743 );
and ( n54745 , n52130 , n53972 );
and ( n54746 , n52098 , n53970 );
nor ( n54747 , n54745 , n54746 );
xnor ( n54748 , n54747 , n53662 );
and ( n54749 , n54744 , n54748 );
xor ( n54750 , n54456 , n54483 );
xor ( n54751 , n54750 , n54488 );
and ( n54752 , n54748 , n54751 );
and ( n54753 , n54744 , n54751 );
or ( n54754 , n54749 , n54752 , n54753 );
and ( n54755 , n54704 , n54754 );
and ( n54756 , n54665 , n54754 );
or ( n54757 , n54705 , n54755 , n54756 );
and ( n54758 , n54078 , n52121 );
and ( n54759 , n53895 , n52119 );
nor ( n54760 , n54758 , n54759 );
xnor ( n54761 , n54760 , n52087 );
and ( n54762 , n54466 , n52092 );
and ( n54763 , n54364 , n52090 );
nor ( n54764 , n54762 , n54763 );
xnor ( n54765 , n54764 , n52072 );
and ( n54766 , n54761 , n54765 );
buf ( n54767 , n51705 );
and ( n54768 , n54767 , n52059 );
and ( n54769 , n54715 , n52057 );
nor ( n54770 , n54768 , n54769 );
not ( n54771 , n54770 );
and ( n54772 , n54765 , n54771 );
and ( n54773 , n54761 , n54771 );
or ( n54774 , n54766 , n54772 , n54773 );
and ( n54775 , n53644 , n52318 );
and ( n54776 , n53499 , n52316 );
nor ( n54777 , n54775 , n54776 );
xnor ( n54778 , n54777 , n52213 );
and ( n54779 , n54774 , n54778 );
and ( n54780 , n53785 , n52170 );
and ( n54781 , n53652 , n52168 );
nor ( n54782 , n54780 , n54781 );
xnor ( n54783 , n54782 , n52152 );
and ( n54784 , n54778 , n54783 );
and ( n54785 , n54774 , n54783 );
or ( n54786 , n54779 , n54784 , n54785 );
and ( n54787 , n53150 , n52540 );
and ( n54788 , n52952 , n52538 );
nor ( n54789 , n54787 , n54788 );
xnor ( n54790 , n54789 , n52424 );
and ( n54791 , n53322 , n52346 );
and ( n54792 , n53148 , n52344 );
nor ( n54793 , n54791 , n54792 );
xnor ( n54794 , n54793 , n52300 );
and ( n54795 , n54790 , n54794 );
xor ( n54796 , n54709 , n54713 );
xor ( n54797 , n54796 , n54719 );
and ( n54798 , n54794 , n54797 );
and ( n54799 , n54790 , n54797 );
or ( n54800 , n54795 , n54798 , n54799 );
and ( n54801 , n54786 , n54800 );
and ( n54802 , n52952 , n52540 );
and ( n54803 , n52954 , n52538 );
nor ( n54804 , n54802 , n54803 );
xnor ( n54805 , n54804 , n52424 );
and ( n54806 , n54800 , n54805 );
and ( n54807 , n54786 , n54805 );
or ( n54808 , n54801 , n54806 , n54807 );
and ( n54809 , n52307 , n53455 );
and ( n54810 , n52271 , n53453 );
nor ( n54811 , n54809 , n54810 );
xnor ( n54812 , n54811 , n53159 );
and ( n54813 , n54808 , n54812 );
xor ( n54814 , n54734 , n54738 );
xor ( n54815 , n54814 , n54741 );
and ( n54816 , n54812 , n54815 );
and ( n54817 , n54808 , n54815 );
or ( n54818 , n54813 , n54816 , n54817 );
xor ( n54819 , n54590 , n54594 );
xor ( n54820 , n54819 , n54599 );
and ( n54821 , n54818 , n54820 );
xor ( n54822 , n54521 , n54523 );
xor ( n54823 , n54822 , n54526 );
and ( n54824 , n54820 , n54823 );
and ( n54825 , n54818 , n54823 );
or ( n54826 , n54821 , n54824 , n54825 );
xor ( n54827 , n54529 , n54533 );
xor ( n54828 , n54827 , n54538 );
and ( n54829 , n54826 , n54828 );
xor ( n54830 , n54545 , n54549 );
xor ( n54831 , n54830 , n54552 );
and ( n54832 , n54828 , n54831 );
and ( n54833 , n54826 , n54831 );
or ( n54834 , n54829 , n54832 , n54833 );
and ( n54835 , n54757 , n54834 );
xor ( n54836 , n54501 , n54503 );
xor ( n54837 , n54836 , n54506 );
and ( n54838 , n54834 , n54837 );
and ( n54839 , n54757 , n54837 );
or ( n54840 , n54835 , n54838 , n54839 );
xor ( n54841 , n54610 , n54612 );
xor ( n54842 , n54841 , n54615 );
xor ( n54843 , n54541 , n54555 );
xor ( n54844 , n54843 , n54558 );
and ( n54845 , n54842 , n54844 );
xor ( n54846 , n54757 , n54834 );
xor ( n54847 , n54846 , n54837 );
and ( n54848 , n54844 , n54847 );
and ( n54849 , n54842 , n54847 );
or ( n54850 , n54845 , n54848 , n54849 );
and ( n54851 , n54840 , n54850 );
xor ( n54852 , n54618 , n54620 );
xor ( n54853 , n54852 , n54623 );
and ( n54854 , n54850 , n54853 );
and ( n54855 , n54840 , n54853 );
or ( n54856 , n54851 , n54854 , n54855 );
and ( n54857 , n54637 , n54856 );
xor ( n54858 , n54840 , n54850 );
xor ( n54859 , n54858 , n54853 );
and ( n54860 , n52063 , n54693 );
and ( n54861 , n52054 , n54691 );
nor ( n54862 , n54860 , n54861 );
xnor ( n54863 , n54862 , n53892 );
and ( n54864 , n52098 , n54285 );
and ( n54865 , n52061 , n54283 );
nor ( n54866 , n54864 , n54865 );
xnor ( n54867 , n54866 , n53794 );
and ( n54868 , n54863 , n54867 );
and ( n54869 , n52220 , n53739 );
and ( n54870 , n52186 , n53737 );
nor ( n54871 , n54869 , n54870 );
xnor ( n54872 , n54871 , n53315 );
and ( n54873 , n54867 , n54872 );
and ( n54874 , n54863 , n54872 );
or ( n54875 , n54868 , n54873 , n54874 );
and ( n54876 , n54364 , n52121 );
and ( n54877 , n54078 , n52119 );
nor ( n54878 , n54876 , n54877 );
xnor ( n54879 , n54878 , n52087 );
and ( n54880 , n54715 , n52092 );
and ( n54881 , n54466 , n52090 );
nor ( n54882 , n54880 , n54881 );
xnor ( n54883 , n54882 , n52072 );
and ( n54884 , n54879 , n54883 );
buf ( n54885 , n51706 );
and ( n54886 , n54885 , n52059 );
and ( n54887 , n54767 , n52057 );
nor ( n54888 , n54886 , n54887 );
not ( n54889 , n54888 );
and ( n54890 , n54883 , n54889 );
and ( n54891 , n54879 , n54889 );
or ( n54892 , n54884 , n54890 , n54891 );
and ( n54893 , n53652 , n52318 );
and ( n54894 , n53644 , n52316 );
nor ( n54895 , n54893 , n54894 );
xnor ( n54896 , n54895 , n52213 );
and ( n54897 , n54892 , n54896 );
and ( n54898 , n53783 , n52170 );
and ( n54899 , n53785 , n52168 );
nor ( n54900 , n54898 , n54899 );
xnor ( n54901 , n54900 , n52152 );
and ( n54902 , n54896 , n54901 );
and ( n54903 , n54892 , n54901 );
or ( n54904 , n54897 , n54902 , n54903 );
and ( n54905 , n53148 , n52540 );
and ( n54906 , n53150 , n52538 );
nor ( n54907 , n54905 , n54906 );
xnor ( n54908 , n54907 , n52424 );
and ( n54909 , n53499 , n52346 );
and ( n54910 , n53322 , n52344 );
nor ( n54911 , n54909 , n54910 );
xnor ( n54912 , n54911 , n52300 );
and ( n54913 , n54908 , n54912 );
xor ( n54914 , n54761 , n54765 );
xor ( n54915 , n54914 , n54771 );
and ( n54916 , n54912 , n54915 );
and ( n54917 , n54908 , n54915 );
or ( n54918 , n54913 , n54916 , n54917 );
and ( n54919 , n54904 , n54918 );
and ( n54920 , n52954 , n52617 );
and ( n54921 , n52829 , n52615 );
nor ( n54922 , n54920 , n54921 );
xnor ( n54923 , n54922 , n52558 );
and ( n54924 , n54918 , n54923 );
and ( n54925 , n54904 , n54923 );
or ( n54926 , n54919 , n54924 , n54925 );
and ( n54927 , n52439 , n53293 );
and ( n54928 , n52431 , n53291 );
nor ( n54929 , n54927 , n54928 );
xnor ( n54930 , n54929 , n52963 );
and ( n54931 , n54926 , n54930 );
and ( n54932 , n52718 , n52886 );
and ( n54933 , n52664 , n52884 );
nor ( n54934 , n54932 , n54933 );
xnor ( n54935 , n54934 , n52657 );
and ( n54936 , n54930 , n54935 );
and ( n54937 , n54926 , n54935 );
or ( n54938 , n54931 , n54936 , n54937 );
and ( n54939 , n52639 , n53021 );
and ( n54940 , n52565 , n53019 );
nor ( n54941 , n54939 , n54940 );
xnor ( n54942 , n54941 , n52839 );
xor ( n54943 , n54722 , n54726 );
xor ( n54944 , n54943 , n54731 );
and ( n54945 , n54942 , n54944 );
xor ( n54946 , n54669 , n54673 );
xor ( n54947 , n54946 , n54676 );
and ( n54948 , n54944 , n54947 );
and ( n54949 , n54942 , n54947 );
or ( n54950 , n54945 , n54948 , n54949 );
and ( n54951 , n54938 , n54950 );
and ( n54952 , n52159 , n53972 );
and ( n54953 , n52130 , n53970 );
nor ( n54954 , n54952 , n54953 );
xnor ( n54955 , n54954 , n53662 );
and ( n54956 , n54950 , n54955 );
and ( n54957 , n54938 , n54955 );
or ( n54958 , n54951 , n54956 , n54957 );
and ( n54959 , n54875 , n54958 );
xor ( n54960 , n54744 , n54748 );
xor ( n54961 , n54960 , n54751 );
and ( n54962 , n54958 , n54961 );
and ( n54963 , n54875 , n54961 );
or ( n54964 , n54959 , n54962 , n54963 );
xor ( n54965 , n54665 , n54704 );
xor ( n54966 , n54965 , n54754 );
and ( n54967 , n54964 , n54966 );
xor ( n54968 , n54602 , n54604 );
xor ( n54969 , n54968 , n54607 );
and ( n54970 , n54966 , n54969 );
and ( n54971 , n54964 , n54969 );
or ( n54972 , n54967 , n54970 , n54971 );
xor ( n54973 , n54653 , n54657 );
xor ( n54974 , n54973 , n54662 );
xor ( n54975 , n54689 , n54696 );
xor ( n54976 , n54975 , n54701 );
and ( n54977 , n54974 , n54976 );
xor ( n54978 , n54818 , n54820 );
xor ( n54979 , n54978 , n54823 );
and ( n54980 , n54976 , n54979 );
and ( n54981 , n54974 , n54979 );
or ( n54982 , n54977 , n54980 , n54981 );
xor ( n54983 , n54826 , n54828 );
xor ( n54984 , n54983 , n54831 );
and ( n54985 , n54982 , n54984 );
xor ( n54986 , n54964 , n54966 );
xor ( n54987 , n54986 , n54969 );
and ( n54988 , n54984 , n54987 );
and ( n54989 , n54982 , n54987 );
or ( n54990 , n54985 , n54988 , n54989 );
and ( n54991 , n54972 , n54990 );
xor ( n54992 , n54842 , n54844 );
xor ( n54993 , n54992 , n54847 );
and ( n54994 , n54990 , n54993 );
and ( n54995 , n54972 , n54993 );
or ( n54996 , n54991 , n54994 , n54995 );
and ( n54997 , n54859 , n54996 );
and ( n54998 , n52061 , n54693 );
and ( n54999 , n52063 , n54691 );
nor ( n55000 , n54998 , n54999 );
xnor ( n55001 , n55000 , n53892 );
and ( n55002 , n52130 , n54285 );
and ( n55003 , n52098 , n54283 );
nor ( n55004 , n55002 , n55003 );
xnor ( n55005 , n55004 , n53794 );
and ( n55006 , n55001 , n55005 );
and ( n55007 , n52271 , n53739 );
and ( n55008 , n52220 , n53737 );
nor ( n55009 , n55007 , n55008 );
xnor ( n55010 , n55009 , n53315 );
and ( n55011 , n55005 , n55010 );
and ( n55012 , n55001 , n55010 );
or ( n55013 , n55006 , n55011 , n55012 );
and ( n55014 , n52431 , n53455 );
and ( n55015 , n52371 , n53453 );
nor ( n55016 , n55014 , n55015 );
xnor ( n55017 , n55016 , n53159 );
and ( n55018 , n52565 , n53293 );
and ( n55019 , n52439 , n53291 );
nor ( n55020 , n55018 , n55019 );
xnor ( n55021 , n55020 , n52963 );
and ( n55022 , n55017 , n55021 );
and ( n55023 , n52664 , n53021 );
and ( n55024 , n52639 , n53019 );
nor ( n55025 , n55023 , n55024 );
xnor ( n55026 , n55025 , n52839 );
and ( n55027 , n55021 , n55026 );
and ( n55028 , n55017 , n55026 );
or ( n55029 , n55022 , n55027 , n55028 );
buf ( n55030 , n52053 );
xor ( n55031 , n53885 , n55030 );
not ( n55032 , n55030 );
and ( n55033 , n55031 , n55032 );
and ( n55034 , n52054 , n55033 );
not ( n55035 , n55034 );
xnor ( n55036 , n55035 , n53885 );
and ( n55037 , n55029 , n55036 );
and ( n55038 , n52186 , n53972 );
and ( n55039 , n52159 , n53970 );
nor ( n55040 , n55038 , n55039 );
xnor ( n55041 , n55040 , n53662 );
and ( n55042 , n55036 , n55041 );
and ( n55043 , n55029 , n55041 );
or ( n55044 , n55037 , n55042 , n55043 );
and ( n55045 , n55013 , n55044 );
and ( n55046 , n54078 , n52170 );
and ( n55047 , n53895 , n52168 );
nor ( n55048 , n55046 , n55047 );
xnor ( n55049 , n55048 , n52152 );
and ( n55050 , n54767 , n52092 );
and ( n55051 , n54715 , n52090 );
nor ( n55052 , n55050 , n55051 );
xnor ( n55053 , n55052 , n52072 );
and ( n55054 , n55049 , n55053 );
buf ( n55055 , n51707 );
and ( n55056 , n55055 , n52059 );
and ( n55057 , n54885 , n52057 );
nor ( n55058 , n55056 , n55057 );
not ( n55059 , n55058 );
and ( n55060 , n55053 , n55059 );
and ( n55061 , n55049 , n55059 );
or ( n55062 , n55054 , n55060 , n55061 );
and ( n55063 , n53785 , n52318 );
and ( n55064 , n53652 , n52316 );
nor ( n55065 , n55063 , n55064 );
xnor ( n55066 , n55065 , n52213 );
and ( n55067 , n55062 , n55066 );
and ( n55068 , n53895 , n52170 );
and ( n55069 , n53783 , n52168 );
nor ( n55070 , n55068 , n55069 );
xnor ( n55071 , n55070 , n52152 );
and ( n55072 , n55066 , n55071 );
and ( n55073 , n55062 , n55071 );
or ( n55074 , n55067 , n55072 , n55073 );
and ( n55075 , n52829 , n52886 );
and ( n55076 , n52809 , n52884 );
nor ( n55077 , n55075 , n55076 );
xnor ( n55078 , n55077 , n52657 );
and ( n55079 , n55074 , n55078 );
and ( n55080 , n52952 , n52617 );
and ( n55081 , n52954 , n52615 );
nor ( n55082 , n55080 , n55081 );
xnor ( n55083 , n55082 , n52558 );
and ( n55084 , n55078 , n55083 );
and ( n55085 , n55074 , n55083 );
or ( n55086 , n55079 , n55084 , n55085 );
xor ( n55087 , n54774 , n54778 );
xor ( n55088 , n55087 , n54783 );
and ( n55089 , n55086 , n55088 );
xor ( n55090 , n54790 , n54794 );
xor ( n55091 , n55090 , n54797 );
and ( n55092 , n55088 , n55091 );
and ( n55093 , n55086 , n55091 );
or ( n55094 , n55089 , n55092 , n55093 );
and ( n55095 , n52371 , n53455 );
and ( n55096 , n52307 , n53453 );
nor ( n55097 , n55095 , n55096 );
xnor ( n55098 , n55097 , n53159 );
and ( n55099 , n55094 , n55098 );
xor ( n55100 , n54786 , n54800 );
xor ( n55101 , n55100 , n54805 );
and ( n55102 , n55098 , n55101 );
and ( n55103 , n55094 , n55101 );
or ( n55104 , n55099 , n55102 , n55103 );
and ( n55105 , n55044 , n55104 );
and ( n55106 , n55013 , n55104 );
or ( n55107 , n55045 , n55105 , n55106 );
and ( n55108 , n53322 , n52540 );
and ( n55109 , n53148 , n52538 );
nor ( n55110 , n55108 , n55109 );
xnor ( n55111 , n55110 , n52424 );
and ( n55112 , n53644 , n52346 );
and ( n55113 , n53499 , n52344 );
nor ( n55114 , n55112 , n55113 );
xnor ( n55115 , n55114 , n52300 );
and ( n55116 , n55111 , n55115 );
xor ( n55117 , n54879 , n54883 );
xor ( n55118 , n55117 , n54889 );
and ( n55119 , n55115 , n55118 );
and ( n55120 , n55111 , n55118 );
or ( n55121 , n55116 , n55119 , n55120 );
xor ( n55122 , n54892 , n54896 );
xor ( n55123 , n55122 , n54901 );
and ( n55124 , n55121 , n55123 );
xor ( n55125 , n54908 , n54912 );
xor ( n55126 , n55125 , n54915 );
and ( n55127 , n55123 , n55126 );
and ( n55128 , n55121 , n55126 );
or ( n55129 , n55124 , n55127 , n55128 );
and ( n55130 , n52809 , n52886 );
and ( n55131 , n52718 , n52884 );
nor ( n55132 , n55130 , n55131 );
xnor ( n55133 , n55132 , n52657 );
and ( n55134 , n55129 , n55133 );
xor ( n55135 , n54904 , n54918 );
xor ( n55136 , n55135 , n54923 );
and ( n55137 , n55133 , n55136 );
and ( n55138 , n55129 , n55136 );
or ( n55139 , n55134 , n55137 , n55138 );
xor ( n55140 , n54926 , n54930 );
xor ( n55141 , n55140 , n54935 );
and ( n55142 , n55139 , n55141 );
xor ( n55143 , n54942 , n54944 );
xor ( n55144 , n55143 , n54947 );
and ( n55145 , n55141 , n55144 );
and ( n55146 , n55139 , n55144 );
or ( n55147 , n55142 , n55145 , n55146 );
xor ( n55148 , n54863 , n54867 );
xor ( n55149 , n55148 , n54872 );
and ( n55150 , n55147 , n55149 );
xor ( n55151 , n54938 , n54950 );
xor ( n55152 , n55151 , n54955 );
and ( n55153 , n55149 , n55152 );
and ( n55154 , n55147 , n55152 );
or ( n55155 , n55150 , n55153 , n55154 );
and ( n55156 , n55107 , n55155 );
xor ( n55157 , n54641 , n54645 );
xor ( n55158 , n55157 , n54650 );
xor ( n55159 , n54679 , n54683 );
xor ( n55160 , n55159 , n54686 );
and ( n55161 , n55158 , n55160 );
xor ( n55162 , n54808 , n54812 );
xor ( n55163 , n55162 , n54815 );
and ( n55164 , n55160 , n55163 );
and ( n55165 , n55158 , n55163 );
or ( n55166 , n55161 , n55164 , n55165 );
and ( n55167 , n55155 , n55166 );
and ( n55168 , n55107 , n55166 );
or ( n55169 , n55156 , n55167 , n55168 );
and ( n55170 , n52098 , n54693 );
and ( n55171 , n52061 , n54691 );
nor ( n55172 , n55170 , n55171 );
xnor ( n55173 , n55172 , n53892 );
xor ( n55174 , n55017 , n55021 );
xor ( n55175 , n55174 , n55026 );
and ( n55176 , n55173 , n55175 );
xor ( n55177 , n55129 , n55133 );
xor ( n55178 , n55177 , n55136 );
and ( n55179 , n55175 , n55178 );
and ( n55180 , n55173 , n55178 );
or ( n55181 , n55176 , n55179 , n55180 );
xor ( n55182 , n55001 , n55005 );
xor ( n55183 , n55182 , n55010 );
and ( n55184 , n55181 , n55183 );
xor ( n55185 , n55029 , n55036 );
xor ( n55186 , n55185 , n55041 );
and ( n55187 , n55183 , n55186 );
and ( n55188 , n55181 , n55186 );
or ( n55189 , n55184 , n55187 , n55188 );
and ( n55190 , n54715 , n52121 );
and ( n55191 , n54466 , n52119 );
nor ( n55192 , n55190 , n55191 );
xnor ( n55193 , n55192 , n52087 );
and ( n55194 , n54885 , n52092 );
and ( n55195 , n54767 , n52090 );
nor ( n55196 , n55194 , n55195 );
xnor ( n55197 , n55196 , n52072 );
and ( n55198 , n55193 , n55197 );
buf ( n55199 , n51708 );
and ( n55200 , n55199 , n52059 );
and ( n55201 , n55055 , n52057 );
nor ( n55202 , n55200 , n55201 );
not ( n55203 , n55202 );
and ( n55204 , n55197 , n55203 );
and ( n55205 , n55193 , n55203 );
or ( n55206 , n55198 , n55204 , n55205 );
and ( n55207 , n53783 , n52318 );
and ( n55208 , n53785 , n52316 );
nor ( n55209 , n55207 , n55208 );
xnor ( n55210 , n55209 , n52213 );
and ( n55211 , n55206 , n55210 );
and ( n55212 , n54466 , n52121 );
and ( n55213 , n54364 , n52119 );
nor ( n55214 , n55212 , n55213 );
xnor ( n55215 , n55214 , n52087 );
and ( n55216 , n55210 , n55215 );
and ( n55217 , n55206 , n55215 );
or ( n55218 , n55211 , n55216 , n55217 );
and ( n55219 , n52954 , n52886 );
and ( n55220 , n52829 , n52884 );
nor ( n55221 , n55219 , n55220 );
xnor ( n55222 , n55221 , n52657 );
and ( n55223 , n55218 , n55222 );
and ( n55224 , n53150 , n52617 );
and ( n55225 , n52952 , n52615 );
nor ( n55226 , n55224 , n55225 );
xnor ( n55227 , n55226 , n52558 );
and ( n55228 , n55222 , n55227 );
and ( n55229 , n55218 , n55227 );
or ( n55230 , n55223 , n55228 , n55229 );
and ( n55231 , n52439 , n53455 );
and ( n55232 , n52431 , n53453 );
nor ( n55233 , n55231 , n55232 );
xnor ( n55234 , n55233 , n53159 );
and ( n55235 , n55230 , n55234 );
and ( n55236 , n52639 , n53293 );
and ( n55237 , n52565 , n53291 );
nor ( n55238 , n55236 , n55237 );
xnor ( n55239 , n55238 , n52963 );
and ( n55240 , n55234 , n55239 );
and ( n55241 , n55230 , n55239 );
or ( n55242 , n55235 , n55240 , n55241 );
and ( n55243 , n52063 , n55033 );
and ( n55244 , n52054 , n55030 );
nor ( n55245 , n55243 , n55244 );
xnor ( n55246 , n55245 , n53885 );
and ( n55247 , n55242 , n55246 );
and ( n55248 , n52220 , n53972 );
and ( n55249 , n52186 , n53970 );
nor ( n55250 , n55248 , n55249 );
xnor ( n55251 , n55250 , n53662 );
and ( n55252 , n55246 , n55251 );
and ( n55253 , n55242 , n55251 );
or ( n55254 , n55247 , n55252 , n55253 );
and ( n55255 , n52159 , n54285 );
and ( n55256 , n52130 , n54283 );
nor ( n55257 , n55255 , n55256 );
xnor ( n55258 , n55257 , n53794 );
and ( n55259 , n52307 , n53739 );
and ( n55260 , n52271 , n53737 );
nor ( n55261 , n55259 , n55260 );
xnor ( n55262 , n55261 , n53315 );
and ( n55263 , n55258 , n55262 );
xor ( n55264 , n55086 , n55088 );
xor ( n55265 , n55264 , n55091 );
and ( n55266 , n55262 , n55265 );
and ( n55267 , n55258 , n55265 );
or ( n55268 , n55263 , n55266 , n55267 );
and ( n55269 , n55254 , n55268 );
xor ( n55270 , n55094 , n55098 );
xor ( n55271 , n55270 , n55101 );
and ( n55272 , n55268 , n55271 );
and ( n55273 , n55254 , n55271 );
or ( n55274 , n55269 , n55272 , n55273 );
and ( n55275 , n55189 , n55274 );
xor ( n55276 , n55158 , n55160 );
xor ( n55277 , n55276 , n55163 );
and ( n55278 , n55274 , n55277 );
and ( n55279 , n55189 , n55277 );
or ( n55280 , n55275 , n55278 , n55279 );
xor ( n55281 , n54875 , n54958 );
xor ( n55282 , n55281 , n54961 );
and ( n55283 , n55280 , n55282 );
xor ( n55284 , n54974 , n54976 );
xor ( n55285 , n55284 , n54979 );
and ( n55286 , n55282 , n55285 );
and ( n55287 , n55280 , n55285 );
or ( n55288 , n55283 , n55286 , n55287 );
and ( n55289 , n55169 , n55288 );
xor ( n55290 , n54982 , n54984 );
xor ( n55291 , n55290 , n54987 );
and ( n55292 , n55288 , n55291 );
and ( n55293 , n55169 , n55291 );
or ( n55294 , n55289 , n55292 , n55293 );
xor ( n55295 , n54972 , n54990 );
xor ( n55296 , n55295 , n54993 );
and ( n55297 , n55294 , n55296 );
xor ( n55298 , n55169 , n55288 );
xor ( n55299 , n55298 , n55291 );
xor ( n55300 , n55013 , n55044 );
xor ( n55301 , n55300 , n55104 );
xor ( n55302 , n55147 , n55149 );
xor ( n55303 , n55302 , n55152 );
and ( n55304 , n55301 , n55303 );
xor ( n55305 , n55189 , n55274 );
xor ( n55306 , n55305 , n55277 );
and ( n55307 , n55303 , n55306 );
and ( n55308 , n55301 , n55306 );
or ( n55309 , n55304 , n55307 , n55308 );
xor ( n55310 , n55107 , n55155 );
xor ( n55311 , n55310 , n55166 );
and ( n55312 , n55309 , n55311 );
xor ( n55313 , n55280 , n55282 );
xor ( n55314 , n55313 , n55285 );
and ( n55315 , n55311 , n55314 );
and ( n55316 , n55309 , n55314 );
or ( n55317 , n55312 , n55315 , n55316 );
and ( n55318 , n55299 , n55317 );
xor ( n55319 , n55309 , n55311 );
xor ( n55320 , n55319 , n55314 );
and ( n55321 , n52307 , n53972 );
and ( n55322 , n52271 , n53970 );
nor ( n55323 , n55321 , n55322 );
xnor ( n55324 , n55323 , n53662 );
and ( n55325 , n52664 , n53293 );
and ( n55326 , n52639 , n53291 );
nor ( n55327 , n55325 , n55326 );
xnor ( n55328 , n55327 , n52963 );
and ( n55329 , n55324 , n55328 );
and ( n55330 , n53148 , n52617 );
and ( n55331 , n53150 , n52615 );
nor ( n55332 , n55330 , n55331 );
xnor ( n55333 , n55332 , n52558 );
and ( n55334 , n53652 , n52346 );
and ( n55335 , n53644 , n52344 );
nor ( n55336 , n55334 , n55335 );
xnor ( n55337 , n55336 , n52300 );
and ( n55338 , n55333 , n55337 );
xor ( n55339 , n55049 , n55053 );
xor ( n55340 , n55339 , n55059 );
and ( n55341 , n55337 , n55340 );
and ( n55342 , n55333 , n55340 );
or ( n55343 , n55338 , n55341 , n55342 );
xor ( n55344 , n55062 , n55066 );
xor ( n55345 , n55344 , n55071 );
xor ( n55346 , n55343 , n55345 );
xor ( n55347 , n55111 , n55115 );
xor ( n55348 , n55347 , n55118 );
xor ( n55349 , n55346 , n55348 );
and ( n55350 , n55328 , n55349 );
and ( n55351 , n55324 , n55349 );
or ( n55352 , n55329 , n55350 , n55351 );
xor ( n55353 , n55230 , n55234 );
xor ( n55354 , n55353 , n55239 );
and ( n55355 , n55352 , n55354 );
and ( n55356 , n54767 , n52121 );
and ( n55357 , n54715 , n52119 );
nor ( n55358 , n55356 , n55357 );
xnor ( n55359 , n55358 , n52087 );
and ( n55360 , n55055 , n52092 );
and ( n55361 , n54885 , n52090 );
nor ( n55362 , n55360 , n55361 );
xnor ( n55363 , n55362 , n52072 );
and ( n55364 , n55359 , n55363 );
buf ( n55365 , n51709 );
and ( n55366 , n55365 , n52059 );
and ( n55367 , n55199 , n52057 );
nor ( n55368 , n55366 , n55367 );
not ( n55369 , n55368 );
and ( n55370 , n55363 , n55369 );
and ( n55371 , n55359 , n55369 );
or ( n55372 , n55364 , n55370 , n55371 );
and ( n55373 , n53895 , n52318 );
and ( n55374 , n53783 , n52316 );
nor ( n55375 , n55373 , n55374 );
xnor ( n55376 , n55375 , n52213 );
and ( n55377 , n55372 , n55376 );
and ( n55378 , n54364 , n52170 );
and ( n55379 , n54078 , n52168 );
nor ( n55380 , n55378 , n55379 );
xnor ( n55381 , n55380 , n52152 );
and ( n55382 , n55376 , n55381 );
and ( n55383 , n55372 , n55381 );
or ( n55384 , n55377 , n55382 , n55383 );
and ( n55385 , n52829 , n53021 );
and ( n55386 , n52809 , n53019 );
nor ( n55387 , n55385 , n55386 );
xnor ( n55388 , n55387 , n52839 );
and ( n55389 , n55384 , n55388 );
and ( n55390 , n53499 , n52540 );
and ( n55391 , n53322 , n52538 );
nor ( n55392 , n55390 , n55391 );
xnor ( n55393 , n55392 , n52424 );
and ( n55394 , n55388 , n55393 );
and ( n55395 , n55384 , n55393 );
or ( n55396 , n55389 , n55394 , n55395 );
and ( n55397 , n54885 , n52121 );
and ( n55398 , n54767 , n52119 );
nor ( n55399 , n55397 , n55398 );
xnor ( n55400 , n55399 , n52087 );
and ( n55401 , n55199 , n52092 );
and ( n55402 , n55055 , n52090 );
nor ( n55403 , n55401 , n55402 );
xnor ( n55404 , n55403 , n52072 );
and ( n55405 , n55400 , n55404 );
buf ( n55406 , n51710 );
and ( n55407 , n55406 , n52059 );
and ( n55408 , n55365 , n52057 );
nor ( n55409 , n55407 , n55408 );
not ( n55410 , n55409 );
and ( n55411 , n55404 , n55410 );
and ( n55412 , n55400 , n55410 );
or ( n55413 , n55405 , n55411 , n55412 );
and ( n55414 , n54078 , n52318 );
and ( n55415 , n53895 , n52316 );
nor ( n55416 , n55414 , n55415 );
xnor ( n55417 , n55416 , n52213 );
and ( n55418 , n55413 , n55417 );
and ( n55419 , n54466 , n52170 );
and ( n55420 , n54364 , n52168 );
nor ( n55421 , n55419 , n55420 );
xnor ( n55422 , n55421 , n52152 );
and ( n55423 , n55417 , n55422 );
and ( n55424 , n55413 , n55422 );
or ( n55425 , n55418 , n55423 , n55424 );
and ( n55426 , n53785 , n52346 );
and ( n55427 , n53652 , n52344 );
nor ( n55428 , n55426 , n55427 );
xnor ( n55429 , n55428 , n52300 );
and ( n55430 , n55425 , n55429 );
xor ( n55431 , n55193 , n55197 );
xor ( n55432 , n55431 , n55203 );
and ( n55433 , n55429 , n55432 );
and ( n55434 , n55425 , n55432 );
or ( n55435 , n55430 , n55433 , n55434 );
and ( n55436 , n52952 , n52886 );
and ( n55437 , n52954 , n52884 );
nor ( n55438 , n55436 , n55437 );
xnor ( n55439 , n55438 , n52657 );
and ( n55440 , n55435 , n55439 );
xor ( n55441 , n55206 , n55210 );
xor ( n55442 , n55441 , n55215 );
and ( n55443 , n55439 , n55442 );
and ( n55444 , n55435 , n55442 );
or ( n55445 , n55440 , n55443 , n55444 );
and ( n55446 , n55396 , n55445 );
xor ( n55447 , n55218 , n55222 );
xor ( n55448 , n55447 , n55227 );
and ( n55449 , n55445 , n55448 );
and ( n55450 , n55396 , n55448 );
or ( n55451 , n55446 , n55449 , n55450 );
and ( n55452 , n52371 , n53739 );
and ( n55453 , n52307 , n53737 );
nor ( n55454 , n55452 , n55453 );
xnor ( n55455 , n55454 , n53315 );
xor ( n55456 , n55451 , n55455 );
xor ( n55457 , n55121 , n55123 );
xor ( n55458 , n55457 , n55126 );
xor ( n55459 , n55456 , n55458 );
and ( n55460 , n55354 , n55459 );
and ( n55461 , n55352 , n55459 );
or ( n55462 , n55355 , n55460 , n55461 );
and ( n55463 , n52130 , n54693 );
and ( n55464 , n52098 , n54691 );
nor ( n55465 , n55463 , n55464 );
xnor ( n55466 , n55465 , n53892 );
and ( n55467 , n52186 , n54285 );
and ( n55468 , n52159 , n54283 );
nor ( n55469 , n55467 , n55468 );
xnor ( n55470 , n55469 , n53794 );
and ( n55471 , n55466 , n55470 );
and ( n55472 , n52271 , n53972 );
and ( n55473 , n52220 , n53970 );
nor ( n55474 , n55472 , n55473 );
xnor ( n55475 , n55474 , n53662 );
and ( n55476 , n55470 , n55475 );
and ( n55477 , n55466 , n55475 );
or ( n55478 , n55471 , n55476 , n55477 );
and ( n55479 , n55343 , n55345 );
and ( n55480 , n55345 , n55348 );
and ( n55481 , n55343 , n55348 );
or ( n55482 , n55479 , n55480 , n55481 );
and ( n55483 , n52718 , n53021 );
and ( n55484 , n52664 , n53019 );
nor ( n55485 , n55483 , n55484 );
xnor ( n55486 , n55485 , n52839 );
and ( n55487 , n55482 , n55486 );
xor ( n55488 , n55074 , n55078 );
xor ( n55489 , n55488 , n55083 );
and ( n55490 , n55486 , n55489 );
and ( n55491 , n55482 , n55489 );
or ( n55492 , n55487 , n55490 , n55491 );
xor ( n55493 , n55478 , n55492 );
and ( n55494 , n55451 , n55455 );
and ( n55495 , n55455 , n55458 );
and ( n55496 , n55451 , n55458 );
or ( n55497 , n55494 , n55495 , n55496 );
xor ( n55498 , n55493 , n55497 );
and ( n55499 , n55462 , n55498 );
xor ( n55500 , n55173 , n55175 );
xor ( n55501 , n55500 , n55178 );
and ( n55502 , n55498 , n55501 );
and ( n55503 , n55462 , n55501 );
or ( n55504 , n55499 , n55502 , n55503 );
xor ( n55505 , n55181 , n55183 );
xor ( n55506 , n55505 , n55186 );
and ( n55507 , n55504 , n55506 );
xor ( n55508 , n55254 , n55268 );
xor ( n55509 , n55508 , n55271 );
and ( n55510 , n55506 , n55509 );
and ( n55511 , n55504 , n55509 );
or ( n55512 , n55507 , n55510 , n55511 );
and ( n55513 , n55478 , n55492 );
and ( n55514 , n55492 , n55497 );
and ( n55515 , n55478 , n55497 );
or ( n55516 , n55513 , n55514 , n55515 );
and ( n55517 , n52431 , n53739 );
and ( n55518 , n52371 , n53737 );
nor ( n55519 , n55517 , n55518 );
xnor ( n55520 , n55519 , n53315 );
and ( n55521 , n52565 , n53455 );
and ( n55522 , n52439 , n53453 );
nor ( n55523 , n55521 , n55522 );
xnor ( n55524 , n55523 , n53159 );
and ( n55525 , n55520 , n55524 );
and ( n55526 , n52809 , n53021 );
and ( n55527 , n52718 , n53019 );
nor ( n55528 , n55526 , n55527 );
xnor ( n55529 , n55528 , n52839 );
and ( n55530 , n55524 , n55529 );
and ( n55531 , n55520 , n55529 );
or ( n55532 , n55525 , n55530 , n55531 );
and ( n55533 , n52061 , n55033 );
and ( n55534 , n52063 , n55030 );
nor ( n55535 , n55533 , n55534 );
xnor ( n55536 , n55535 , n53885 );
and ( n55537 , n55532 , n55536 );
xor ( n55538 , n55482 , n55486 );
xor ( n55539 , n55538 , n55489 );
and ( n55540 , n55536 , n55539 );
and ( n55541 , n55532 , n55539 );
or ( n55542 , n55537 , n55540 , n55541 );
xor ( n55543 , n55242 , n55246 );
xor ( n55544 , n55543 , n55251 );
and ( n55545 , n55542 , n55544 );
xor ( n55546 , n55258 , n55262 );
xor ( n55547 , n55546 , n55265 );
and ( n55548 , n55544 , n55547 );
and ( n55549 , n55542 , n55547 );
or ( n55550 , n55545 , n55548 , n55549 );
and ( n55551 , n55516 , n55550 );
xor ( n55552 , n55139 , n55141 );
xor ( n55553 , n55552 , n55144 );
and ( n55554 , n55550 , n55553 );
and ( n55555 , n55516 , n55553 );
or ( n55556 , n55551 , n55554 , n55555 );
and ( n55557 , n55512 , n55556 );
xor ( n55558 , n55301 , n55303 );
xor ( n55559 , n55558 , n55306 );
and ( n55560 , n55556 , n55559 );
and ( n55561 , n55512 , n55559 );
or ( n55562 , n55557 , n55560 , n55561 );
and ( n55563 , n55320 , n55562 );
xor ( n55564 , n55512 , n55556 );
xor ( n55565 , n55564 , n55559 );
and ( n55566 , n52439 , n53739 );
and ( n55567 , n52431 , n53737 );
nor ( n55568 , n55566 , n55567 );
xnor ( n55569 , n55568 , n53315 );
and ( n55570 , n52718 , n53293 );
and ( n55571 , n52664 , n53291 );
nor ( n55572 , n55570 , n55571 );
xnor ( n55573 , n55572 , n52963 );
and ( n55574 , n55569 , n55573 );
xor ( n55575 , n55384 , n55388 );
xor ( n55576 , n55575 , n55393 );
and ( n55577 , n55573 , n55576 );
and ( n55578 , n55569 , n55576 );
or ( n55579 , n55574 , n55577 , n55578 );
and ( n55580 , n52098 , n55033 );
and ( n55581 , n52061 , n55030 );
nor ( n55582 , n55580 , n55581 );
xnor ( n55583 , n55582 , n53885 );
and ( n55584 , n55579 , n55583 );
and ( n55585 , n52159 , n54693 );
and ( n55586 , n52130 , n54691 );
nor ( n55587 , n55585 , n55586 );
xnor ( n55588 , n55587 , n53892 );
and ( n55589 , n55583 , n55588 );
and ( n55590 , n55579 , n55588 );
or ( n55591 , n55584 , n55589 , n55590 );
and ( n55592 , n53322 , n52617 );
and ( n55593 , n53148 , n52615 );
nor ( n55594 , n55592 , n55593 );
xnor ( n55595 , n55594 , n52558 );
and ( n55596 , n53644 , n52540 );
and ( n55597 , n53499 , n52538 );
nor ( n55598 , n55596 , n55597 );
xnor ( n55599 , n55598 , n52424 );
and ( n55600 , n55595 , n55599 );
xor ( n55601 , n55372 , n55376 );
xor ( n55602 , n55601 , n55381 );
and ( n55603 , n55599 , n55602 );
and ( n55604 , n55595 , n55602 );
or ( n55605 , n55600 , n55603 , n55604 );
and ( n55606 , n53652 , n52540 );
and ( n55607 , n53644 , n52538 );
nor ( n55608 , n55606 , n55607 );
xnor ( n55609 , n55608 , n52424 );
and ( n55610 , n53783 , n52346 );
and ( n55611 , n53785 , n52344 );
nor ( n55612 , n55610 , n55611 );
xnor ( n55613 , n55612 , n52300 );
and ( n55614 , n55609 , n55613 );
xor ( n55615 , n55359 , n55363 );
xor ( n55616 , n55615 , n55369 );
and ( n55617 , n55613 , n55616 );
and ( n55618 , n55609 , n55616 );
or ( n55619 , n55614 , n55617 , n55618 );
and ( n55620 , n53150 , n52886 );
and ( n55621 , n52952 , n52884 );
nor ( n55622 , n55620 , n55621 );
xnor ( n55623 , n55622 , n52657 );
and ( n55624 , n55619 , n55623 );
xor ( n55625 , n55425 , n55429 );
xor ( n55626 , n55625 , n55432 );
and ( n55627 , n55623 , n55626 );
and ( n55628 , n55619 , n55626 );
or ( n55629 , n55624 , n55627 , n55628 );
and ( n55630 , n55605 , n55629 );
xor ( n55631 , n55333 , n55337 );
xor ( n55632 , n55631 , n55340 );
and ( n55633 , n55629 , n55632 );
and ( n55634 , n55605 , n55632 );
or ( n55635 , n55630 , n55633 , n55634 );
and ( n55636 , n52220 , n54285 );
and ( n55637 , n52186 , n54283 );
nor ( n55638 , n55636 , n55637 );
xnor ( n55639 , n55638 , n53794 );
and ( n55640 , n55635 , n55639 );
xor ( n55641 , n55396 , n55445 );
xor ( n55642 , n55641 , n55448 );
and ( n55643 , n55639 , n55642 );
and ( n55644 , n55635 , n55642 );
or ( n55645 , n55640 , n55643 , n55644 );
and ( n55646 , n55591 , n55645 );
xor ( n55647 , n55466 , n55470 );
xor ( n55648 , n55647 , n55475 );
and ( n55649 , n55645 , n55648 );
and ( n55650 , n55591 , n55648 );
or ( n55651 , n55646 , n55649 , n55650 );
and ( n55652 , n54767 , n52170 );
and ( n55653 , n54715 , n52168 );
nor ( n55654 , n55652 , n55653 );
xnor ( n55655 , n55654 , n52152 );
and ( n55656 , n55365 , n52092 );
and ( n55657 , n55199 , n52090 );
nor ( n55658 , n55656 , n55657 );
xnor ( n55659 , n55658 , n52072 );
and ( n55660 , n55655 , n55659 );
buf ( n55661 , n51711 );
and ( n55662 , n55661 , n52059 );
and ( n55663 , n55406 , n52057 );
nor ( n55664 , n55662 , n55663 );
not ( n55665 , n55664 );
and ( n55666 , n55659 , n55665 );
and ( n55667 , n55655 , n55665 );
or ( n55668 , n55660 , n55666 , n55667 );
and ( n55669 , n54715 , n52170 );
and ( n55670 , n54466 , n52168 );
nor ( n55671 , n55669 , n55670 );
xnor ( n55672 , n55671 , n52152 );
and ( n55673 , n55668 , n55672 );
xor ( n55674 , n55400 , n55404 );
xor ( n55675 , n55674 , n55410 );
and ( n55676 , n55672 , n55675 );
and ( n55677 , n55668 , n55675 );
or ( n55678 , n55673 , n55676 , n55677 );
and ( n55679 , n53148 , n52886 );
and ( n55680 , n53150 , n52884 );
nor ( n55681 , n55679 , n55680 );
xnor ( n55682 , n55681 , n52657 );
and ( n55683 , n55678 , n55682 );
and ( n55684 , n53499 , n52617 );
and ( n55685 , n53322 , n52615 );
nor ( n55686 , n55684 , n55685 );
xnor ( n55687 , n55686 , n52558 );
and ( n55688 , n55682 , n55687 );
and ( n55689 , n55678 , n55687 );
or ( n55690 , n55683 , n55688 , n55689 );
and ( n55691 , n52954 , n53021 );
and ( n55692 , n52829 , n53019 );
nor ( n55693 , n55691 , n55692 );
xnor ( n55694 , n55693 , n52839 );
and ( n55695 , n55690 , n55694 );
xor ( n55696 , n55595 , n55599 );
xor ( n55697 , n55696 , n55602 );
and ( n55698 , n55694 , n55697 );
and ( n55699 , n55690 , n55697 );
or ( n55700 , n55695 , n55698 , n55699 );
and ( n55701 , n52639 , n53455 );
and ( n55702 , n52565 , n53453 );
nor ( n55703 , n55701 , n55702 );
xnor ( n55704 , n55703 , n53159 );
and ( n55705 , n55700 , n55704 );
xor ( n55706 , n55435 , n55439 );
xor ( n55707 , n55706 , n55442 );
and ( n55708 , n55704 , n55707 );
and ( n55709 , n55700 , n55707 );
or ( n55710 , n55705 , n55708 , n55709 );
and ( n55711 , n55199 , n52121 );
and ( n55712 , n55055 , n52119 );
nor ( n55713 , n55711 , n55712 );
xnor ( n55714 , n55713 , n52087 );
and ( n55715 , n55406 , n52092 );
and ( n55716 , n55365 , n52090 );
nor ( n55717 , n55715 , n55716 );
xnor ( n55718 , n55717 , n52072 );
and ( n55719 , n55714 , n55718 );
buf ( n55720 , n51712 );
and ( n55721 , n55720 , n52059 );
and ( n55722 , n55661 , n52057 );
nor ( n55723 , n55721 , n55722 );
not ( n55724 , n55723 );
and ( n55725 , n55718 , n55724 );
and ( n55726 , n55714 , n55724 );
or ( n55727 , n55719 , n55725 , n55726 );
and ( n55728 , n55055 , n52121 );
and ( n55729 , n54885 , n52119 );
nor ( n55730 , n55728 , n55729 );
xnor ( n55731 , n55730 , n52087 );
and ( n55732 , n55727 , n55731 );
xor ( n55733 , n55655 , n55659 );
xor ( n55734 , n55733 , n55665 );
and ( n55735 , n55731 , n55734 );
and ( n55736 , n55727 , n55734 );
or ( n55737 , n55732 , n55735 , n55736 );
and ( n55738 , n53895 , n52346 );
and ( n55739 , n53783 , n52344 );
nor ( n55740 , n55738 , n55739 );
xnor ( n55741 , n55740 , n52300 );
and ( n55742 , n55737 , n55741 );
and ( n55743 , n54364 , n52318 );
and ( n55744 , n54078 , n52316 );
nor ( n55745 , n55743 , n55744 );
xnor ( n55746 , n55745 , n52213 );
and ( n55747 , n55741 , n55746 );
and ( n55748 , n55737 , n55746 );
or ( n55749 , n55742 , n55747 , n55748 );
and ( n55750 , n52829 , n53293 );
and ( n55751 , n52809 , n53291 );
nor ( n55752 , n55750 , n55751 );
xnor ( n55753 , n55752 , n52963 );
and ( n55754 , n55749 , n55753 );
xor ( n55755 , n55413 , n55417 );
xor ( n55756 , n55755 , n55422 );
and ( n55757 , n55753 , n55756 );
and ( n55758 , n55749 , n55756 );
or ( n55759 , n55754 , n55757 , n55758 );
and ( n55760 , n55365 , n52121 );
and ( n55761 , n55199 , n52119 );
nor ( n55762 , n55760 , n55761 );
xnor ( n55763 , n55762 , n52087 );
and ( n55764 , n55661 , n52092 );
and ( n55765 , n55406 , n52090 );
nor ( n55766 , n55764 , n55765 );
xnor ( n55767 , n55766 , n52072 );
and ( n55768 , n55763 , n55767 );
buf ( n55769 , n51713 );
and ( n55770 , n55769 , n52059 );
and ( n55771 , n55720 , n52057 );
nor ( n55772 , n55770 , n55771 );
not ( n55773 , n55772 );
and ( n55774 , n55767 , n55773 );
and ( n55775 , n55763 , n55773 );
or ( n55776 , n55768 , n55774 , n55775 );
and ( n55777 , n54885 , n52170 );
and ( n55778 , n54767 , n52168 );
nor ( n55779 , n55777 , n55778 );
xnor ( n55780 , n55779 , n52152 );
and ( n55781 , n55776 , n55780 );
xor ( n55782 , n55714 , n55718 );
xor ( n55783 , n55782 , n55724 );
and ( n55784 , n55780 , n55783 );
and ( n55785 , n55776 , n55783 );
or ( n55786 , n55781 , n55784 , n55785 );
and ( n55787 , n54078 , n52346 );
and ( n55788 , n53895 , n52344 );
nor ( n55789 , n55787 , n55788 );
xnor ( n55790 , n55789 , n52300 );
and ( n55791 , n55786 , n55790 );
and ( n55792 , n54466 , n52318 );
and ( n55793 , n54364 , n52316 );
nor ( n55794 , n55792 , n55793 );
xnor ( n55795 , n55794 , n52213 );
and ( n55796 , n55790 , n55795 );
and ( n55797 , n55786 , n55795 );
or ( n55798 , n55791 , n55796 , n55797 );
and ( n55799 , n53785 , n52540 );
and ( n55800 , n53652 , n52538 );
nor ( n55801 , n55799 , n55800 );
xnor ( n55802 , n55801 , n52424 );
and ( n55803 , n55798 , n55802 );
xor ( n55804 , n55668 , n55672 );
xor ( n55805 , n55804 , n55675 );
and ( n55806 , n55802 , n55805 );
and ( n55807 , n55798 , n55805 );
or ( n55808 , n55803 , n55806 , n55807 );
and ( n55809 , n52952 , n53021 );
and ( n55810 , n52954 , n53019 );
nor ( n55811 , n55809 , n55810 );
xnor ( n55812 , n55811 , n52839 );
and ( n55813 , n55808 , n55812 );
xor ( n55814 , n55609 , n55613 );
xor ( n55815 , n55814 , n55616 );
and ( n55816 , n55812 , n55815 );
and ( n55817 , n55808 , n55815 );
or ( n55818 , n55813 , n55816 , n55817 );
and ( n55819 , n55759 , n55818 );
xor ( n55820 , n55619 , n55623 );
xor ( n55821 , n55820 , n55626 );
and ( n55822 , n55818 , n55821 );
and ( n55823 , n55759 , n55821 );
or ( n55824 , n55819 , n55822 , n55823 );
and ( n55825 , n52371 , n53972 );
and ( n55826 , n52307 , n53970 );
nor ( n55827 , n55825 , n55826 );
xnor ( n55828 , n55827 , n53662 );
and ( n55829 , n55824 , n55828 );
xor ( n55830 , n55605 , n55629 );
xor ( n55831 , n55830 , n55632 );
and ( n55832 , n55828 , n55831 );
and ( n55833 , n55824 , n55831 );
or ( n55834 , n55829 , n55832 , n55833 );
and ( n55835 , n55710 , n55834 );
xor ( n55836 , n55520 , n55524 );
xor ( n55837 , n55836 , n55529 );
and ( n55838 , n55834 , n55837 );
and ( n55839 , n55710 , n55837 );
or ( n55840 , n55835 , n55838 , n55839 );
xor ( n55841 , n55532 , n55536 );
xor ( n55842 , n55841 , n55539 );
and ( n55843 , n55840 , n55842 );
xor ( n55844 , n55352 , n55354 );
xor ( n55845 , n55844 , n55459 );
and ( n55846 , n55842 , n55845 );
and ( n55847 , n55840 , n55845 );
or ( n55848 , n55843 , n55846 , n55847 );
and ( n55849 , n55651 , n55848 );
xor ( n55850 , n55542 , n55544 );
xor ( n55851 , n55850 , n55547 );
and ( n55852 , n55848 , n55851 );
and ( n55853 , n55651 , n55851 );
or ( n55854 , n55849 , n55852 , n55853 );
xor ( n55855 , n55504 , n55506 );
xor ( n55856 , n55855 , n55509 );
and ( n55857 , n55854 , n55856 );
xor ( n55858 , n55516 , n55550 );
xor ( n55859 , n55858 , n55553 );
and ( n55860 , n55856 , n55859 );
and ( n55861 , n55854 , n55859 );
or ( n55862 , n55857 , n55860 , n55861 );
and ( n55863 , n55565 , n55862 );
xor ( n55864 , n55854 , n55856 );
xor ( n55865 , n55864 , n55859 );
xor ( n55866 , n55579 , n55583 );
xor ( n55867 , n55866 , n55588 );
xor ( n55868 , n55710 , n55834 );
xor ( n55869 , n55868 , n55837 );
and ( n55870 , n55867 , n55869 );
xor ( n55871 , n55635 , n55639 );
xor ( n55872 , n55871 , n55642 );
and ( n55873 , n55869 , n55872 );
and ( n55874 , n55867 , n55872 );
or ( n55875 , n55870 , n55873 , n55874 );
and ( n55876 , n52431 , n53972 );
and ( n55877 , n52371 , n53970 );
nor ( n55878 , n55876 , n55877 );
xnor ( n55879 , n55878 , n53662 );
and ( n55880 , n52565 , n53739 );
and ( n55881 , n52439 , n53737 );
nor ( n55882 , n55880 , n55881 );
xnor ( n55883 , n55882 , n53315 );
and ( n55884 , n55879 , n55883 );
and ( n55885 , n52809 , n53293 );
and ( n55886 , n52718 , n53291 );
nor ( n55887 , n55885 , n55886 );
xnor ( n55888 , n55887 , n52963 );
and ( n55889 , n55883 , n55888 );
and ( n55890 , n55879 , n55888 );
or ( n55891 , n55884 , n55889 , n55890 );
and ( n55892 , n52186 , n54693 );
and ( n55893 , n52159 , n54691 );
nor ( n55894 , n55892 , n55893 );
xnor ( n55895 , n55894 , n53892 );
and ( n55896 , n55891 , n55895 );
and ( n55897 , n52271 , n54285 );
and ( n55898 , n52220 , n54283 );
nor ( n55899 , n55897 , n55898 );
xnor ( n55900 , n55899 , n53794 );
and ( n55901 , n55895 , n55900 );
and ( n55902 , n55891 , n55900 );
or ( n55903 , n55896 , n55901 , n55902 );
and ( n55904 , n52130 , n55033 );
and ( n55905 , n52098 , n55030 );
nor ( n55906 , n55904 , n55905 );
xnor ( n55907 , n55906 , n53885 );
xor ( n55908 , n55569 , n55573 );
xor ( n55909 , n55908 , n55576 );
and ( n55910 , n55907 , n55909 );
xor ( n55911 , n55700 , n55704 );
xor ( n55912 , n55911 , n55707 );
and ( n55913 , n55909 , n55912 );
and ( n55914 , n55907 , n55912 );
or ( n55915 , n55910 , n55913 , n55914 );
and ( n55916 , n55903 , n55915 );
xor ( n55917 , n55324 , n55328 );
xor ( n55918 , n55917 , n55349 );
and ( n55919 , n55915 , n55918 );
and ( n55920 , n55903 , n55918 );
or ( n55921 , n55916 , n55919 , n55920 );
and ( n55922 , n55875 , n55921 );
xor ( n55923 , n55591 , n55645 );
xor ( n55924 , n55923 , n55648 );
and ( n55925 , n55921 , n55924 );
and ( n55926 , n55875 , n55924 );
or ( n55927 , n55922 , n55925 , n55926 );
xor ( n55928 , n55462 , n55498 );
xor ( n55929 , n55928 , n55501 );
and ( n55930 , n55927 , n55929 );
xor ( n55931 , n55651 , n55848 );
xor ( n55932 , n55931 , n55851 );
and ( n55933 , n55929 , n55932 );
and ( n55934 , n55927 , n55932 );
or ( n55935 , n55930 , n55933 , n55934 );
and ( n55936 , n55865 , n55935 );
xor ( n55937 , n55927 , n55929 );
xor ( n55938 , n55937 , n55932 );
and ( n55939 , n52439 , n53972 );
and ( n55940 , n52431 , n53970 );
nor ( n55941 , n55939 , n55940 );
xnor ( n55942 , n55941 , n53662 );
and ( n55943 , n52639 , n53739 );
and ( n55944 , n52565 , n53737 );
nor ( n55945 , n55943 , n55944 );
xnor ( n55946 , n55945 , n53315 );
and ( n55947 , n55942 , n55946 );
xor ( n55948 , n55749 , n55753 );
xor ( n55949 , n55948 , n55756 );
and ( n55950 , n55946 , n55949 );
and ( n55951 , n55942 , n55949 );
or ( n55952 , n55947 , n55950 , n55951 );
and ( n55953 , n52159 , n55033 );
and ( n55954 , n52130 , n55030 );
nor ( n55955 , n55953 , n55954 );
xnor ( n55956 , n55955 , n53885 );
and ( n55957 , n55952 , n55956 );
xor ( n55958 , n55879 , n55883 );
xor ( n55959 , n55958 , n55888 );
and ( n55960 , n55956 , n55959 );
and ( n55961 , n55952 , n55959 );
or ( n55962 , n55957 , n55960 , n55961 );
xor ( n55963 , n55891 , n55895 );
xor ( n55964 , n55963 , n55900 );
and ( n55965 , n55962 , n55964 );
xor ( n55966 , n55907 , n55909 );
xor ( n55967 , n55966 , n55912 );
and ( n55968 , n55964 , n55967 );
and ( n55969 , n55962 , n55967 );
or ( n55970 , n55965 , n55968 , n55969 );
and ( n55971 , n52307 , n54285 );
and ( n55972 , n52271 , n54283 );
nor ( n55973 , n55971 , n55972 );
xnor ( n55974 , n55973 , n53794 );
and ( n55975 , n52664 , n53455 );
and ( n55976 , n52639 , n53453 );
nor ( n55977 , n55975 , n55976 );
xnor ( n55978 , n55977 , n53159 );
and ( n55979 , n55974 , n55978 );
xor ( n55980 , n55690 , n55694 );
xor ( n55981 , n55980 , n55697 );
and ( n55982 , n55978 , n55981 );
and ( n55983 , n55974 , n55981 );
or ( n55984 , n55979 , n55982 , n55983 );
and ( n55985 , n53652 , n52617 );
and ( n55986 , n53644 , n52615 );
nor ( n55987 , n55985 , n55986 );
xnor ( n55988 , n55987 , n52558 );
and ( n55989 , n53783 , n52540 );
and ( n55990 , n53785 , n52538 );
nor ( n55991 , n55989 , n55990 );
xnor ( n55992 , n55991 , n52424 );
and ( n55993 , n55988 , n55992 );
xor ( n55994 , n55727 , n55731 );
xor ( n55995 , n55994 , n55734 );
and ( n55996 , n55992 , n55995 );
and ( n55997 , n55988 , n55995 );
or ( n55998 , n55993 , n55996 , n55997 );
and ( n55999 , n52954 , n53293 );
and ( n56000 , n52829 , n53291 );
nor ( n56001 , n55999 , n56000 );
xnor ( n56002 , n56001 , n52963 );
and ( n56003 , n55998 , n56002 );
and ( n56004 , n53150 , n53021 );
and ( n56005 , n52952 , n53019 );
nor ( n56006 , n56004 , n56005 );
xnor ( n56007 , n56006 , n52839 );
and ( n56008 , n56002 , n56007 );
and ( n56009 , n55998 , n56007 );
or ( n56010 , n56003 , n56008 , n56009 );
and ( n56011 , n53322 , n52886 );
and ( n56012 , n53148 , n52884 );
nor ( n56013 , n56011 , n56012 );
xnor ( n56014 , n56013 , n52657 );
and ( n56015 , n53644 , n52617 );
and ( n56016 , n53499 , n52615 );
nor ( n56017 , n56015 , n56016 );
xnor ( n56018 , n56017 , n52558 );
and ( n56019 , n56014 , n56018 );
xor ( n56020 , n55737 , n55741 );
xor ( n56021 , n56020 , n55746 );
and ( n56022 , n56018 , n56021 );
and ( n56023 , n56014 , n56021 );
or ( n56024 , n56019 , n56022 , n56023 );
and ( n56025 , n56010 , n56024 );
xor ( n56026 , n55678 , n55682 );
xor ( n56027 , n56026 , n55687 );
and ( n56028 , n56024 , n56027 );
and ( n56029 , n56010 , n56027 );
or ( n56030 , n56025 , n56028 , n56029 );
and ( n56031 , n52220 , n54693 );
and ( n56032 , n52186 , n54691 );
nor ( n56033 , n56031 , n56032 );
xnor ( n56034 , n56033 , n53892 );
and ( n56035 , n56030 , n56034 );
xor ( n56036 , n55759 , n55818 );
xor ( n56037 , n56036 , n55821 );
and ( n56038 , n56034 , n56037 );
and ( n56039 , n56030 , n56037 );
or ( n56040 , n56035 , n56038 , n56039 );
and ( n56041 , n55984 , n56040 );
xor ( n56042 , n55824 , n55828 );
xor ( n56043 , n56042 , n55831 );
and ( n56044 , n56040 , n56043 );
and ( n56045 , n55984 , n56043 );
or ( n56046 , n56041 , n56044 , n56045 );
and ( n56047 , n55970 , n56046 );
xor ( n56048 , n55903 , n55915 );
xor ( n56049 , n56048 , n55918 );
and ( n56050 , n56046 , n56049 );
and ( n56051 , n55970 , n56049 );
or ( n56052 , n56047 , n56050 , n56051 );
xor ( n56053 , n55875 , n55921 );
xor ( n56054 , n56053 , n55924 );
and ( n56055 , n56052 , n56054 );
xor ( n56056 , n55840 , n55842 );
xor ( n56057 , n56056 , n55845 );
and ( n56058 , n56054 , n56057 );
and ( n56059 , n56052 , n56057 );
or ( n56060 , n56055 , n56058 , n56059 );
and ( n56061 , n55938 , n56060 );
and ( n56062 , n55365 , n52170 );
and ( n56063 , n55199 , n52168 );
nor ( n56064 , n56062 , n56063 );
xnor ( n56065 , n56064 , n52152 );
and ( n56066 , n55769 , n52092 );
and ( n56067 , n55720 , n52090 );
nor ( n56068 , n56066 , n56067 );
xnor ( n56069 , n56068 , n52072 );
and ( n56070 , n56065 , n56069 );
buf ( n56071 , n51715 );
and ( n56072 , n56071 , n52059 );
buf ( n56073 , n51714 );
and ( n56074 , n56073 , n52057 );
nor ( n56075 , n56072 , n56074 );
not ( n56076 , n56075 );
and ( n56077 , n56069 , n56076 );
and ( n56078 , n56065 , n56076 );
or ( n56079 , n56070 , n56077 , n56078 );
and ( n56080 , n54885 , n52318 );
and ( n56081 , n54767 , n52316 );
nor ( n56082 , n56080 , n56081 );
xnor ( n56083 , n56082 , n52213 );
and ( n56084 , n56079 , n56083 );
and ( n56085 , n55199 , n52170 );
and ( n56086 , n55055 , n52168 );
nor ( n56087 , n56085 , n56086 );
xnor ( n56088 , n56087 , n52152 );
and ( n56089 , n56083 , n56088 );
and ( n56090 , n56079 , n56088 );
or ( n56091 , n56084 , n56089 , n56090 );
and ( n56092 , n54466 , n52346 );
and ( n56093 , n54364 , n52344 );
nor ( n56094 , n56092 , n56093 );
xnor ( n56095 , n56094 , n52300 );
and ( n56096 , n56091 , n56095 );
xor ( n56097 , n55763 , n55767 );
xor ( n56098 , n56097 , n55773 );
and ( n56099 , n56095 , n56098 );
and ( n56100 , n56091 , n56098 );
or ( n56101 , n56096 , n56099 , n56100 );
and ( n56102 , n53644 , n52886 );
and ( n56103 , n53499 , n52884 );
nor ( n56104 , n56102 , n56103 );
xnor ( n56105 , n56104 , n52657 );
and ( n56106 , n56101 , n56105 );
and ( n56107 , n55406 , n52121 );
and ( n56108 , n55365 , n52119 );
nor ( n56109 , n56107 , n56108 );
xnor ( n56110 , n56109 , n52087 );
and ( n56111 , n55720 , n52092 );
and ( n56112 , n55661 , n52090 );
nor ( n56113 , n56111 , n56112 );
xnor ( n56114 , n56113 , n52072 );
and ( n56115 , n56110 , n56114 );
and ( n56116 , n56073 , n52059 );
and ( n56117 , n55769 , n52057 );
nor ( n56118 , n56116 , n56117 );
not ( n56119 , n56118 );
and ( n56120 , n56114 , n56119 );
and ( n56121 , n56110 , n56119 );
or ( n56122 , n56115 , n56120 , n56121 );
and ( n56123 , n54767 , n52318 );
and ( n56124 , n54715 , n52316 );
nor ( n56125 , n56123 , n56124 );
xnor ( n56126 , n56125 , n52213 );
and ( n56127 , n56122 , n56126 );
and ( n56128 , n55055 , n52170 );
and ( n56129 , n54885 , n52168 );
nor ( n56130 , n56128 , n56129 );
xnor ( n56131 , n56130 , n52152 );
and ( n56132 , n56126 , n56131 );
and ( n56133 , n56122 , n56131 );
or ( n56134 , n56127 , n56132 , n56133 );
and ( n56135 , n54364 , n52346 );
and ( n56136 , n54078 , n52344 );
nor ( n56137 , n56135 , n56136 );
xnor ( n56138 , n56137 , n52300 );
xor ( n56139 , n56134 , n56138 );
and ( n56140 , n54715 , n52318 );
and ( n56141 , n54466 , n52316 );
nor ( n56142 , n56140 , n56141 );
xnor ( n56143 , n56142 , n52213 );
xor ( n56144 , n56139 , n56143 );
and ( n56145 , n56105 , n56144 );
and ( n56146 , n56101 , n56144 );
or ( n56147 , n56106 , n56145 , n56146 );
and ( n56148 , n52829 , n53455 );
and ( n56149 , n52809 , n53453 );
nor ( n56150 , n56148 , n56149 );
xnor ( n56151 , n56150 , n53159 );
and ( n56152 , n56147 , n56151 );
xor ( n56153 , n55988 , n55992 );
xor ( n56154 , n56153 , n55995 );
and ( n56155 , n56151 , n56154 );
and ( n56156 , n56147 , n56154 );
or ( n56157 , n56152 , n56155 , n56156 );
and ( n56158 , n52565 , n53972 );
and ( n56159 , n52439 , n53970 );
nor ( n56160 , n56158 , n56159 );
xnor ( n56161 , n56160 , n53662 );
and ( n56162 , n56157 , n56161 );
and ( n56163 , n52809 , n53455 );
and ( n56164 , n52718 , n53453 );
nor ( n56165 , n56163 , n56164 );
xnor ( n56166 , n56165 , n53159 );
and ( n56167 , n56161 , n56166 );
and ( n56168 , n56157 , n56166 );
or ( n56169 , n56162 , n56167 , n56168 );
and ( n56170 , n52371 , n54285 );
and ( n56171 , n52307 , n54283 );
nor ( n56172 , n56170 , n56171 );
xnor ( n56173 , n56172 , n53794 );
and ( n56174 , n56169 , n56173 );
xor ( n56175 , n56010 , n56024 );
xor ( n56176 , n56175 , n56027 );
and ( n56177 , n56173 , n56176 );
and ( n56178 , n56169 , n56176 );
or ( n56179 , n56174 , n56177 , n56178 );
and ( n56180 , n52307 , n54693 );
and ( n56181 , n52271 , n54691 );
nor ( n56182 , n56180 , n56181 );
xnor ( n56183 , n56182 , n53892 );
and ( n56184 , n52664 , n53739 );
and ( n56185 , n52639 , n53737 );
nor ( n56186 , n56184 , n56185 );
xnor ( n56187 , n56186 , n53315 );
and ( n56188 , n56183 , n56187 );
and ( n56189 , n56134 , n56138 );
and ( n56190 , n56138 , n56143 );
and ( n56191 , n56134 , n56143 );
or ( n56192 , n56189 , n56190 , n56191 );
and ( n56193 , n53148 , n53021 );
and ( n56194 , n53150 , n53019 );
nor ( n56195 , n56193 , n56194 );
xnor ( n56196 , n56195 , n52839 );
and ( n56197 , n56192 , n56196 );
xor ( n56198 , n55786 , n55790 );
xor ( n56199 , n56198 , n55795 );
and ( n56200 , n56196 , n56199 );
and ( n56201 , n56192 , n56199 );
or ( n56202 , n56197 , n56200 , n56201 );
xor ( n56203 , n56014 , n56018 );
xor ( n56204 , n56203 , n56021 );
xor ( n56205 , n56202 , n56204 );
xor ( n56206 , n55798 , n55802 );
xor ( n56207 , n56206 , n55805 );
xor ( n56208 , n56205 , n56207 );
and ( n56209 , n56187 , n56208 );
and ( n56210 , n56183 , n56208 );
or ( n56211 , n56188 , n56209 , n56210 );
xor ( n56212 , n55942 , n55946 );
xor ( n56213 , n56212 , n55949 );
and ( n56214 , n56211 , n56213 );
and ( n56215 , n56202 , n56204 );
and ( n56216 , n56204 , n56207 );
and ( n56217 , n56202 , n56207 );
or ( n56218 , n56215 , n56216 , n56217 );
and ( n56219 , n52718 , n53455 );
and ( n56220 , n52664 , n53453 );
nor ( n56221 , n56219 , n56220 );
xnor ( n56222 , n56221 , n53159 );
xor ( n56223 , n56218 , n56222 );
xor ( n56224 , n55808 , n55812 );
xor ( n56225 , n56224 , n55815 );
xor ( n56226 , n56223 , n56225 );
and ( n56227 , n56213 , n56226 );
and ( n56228 , n56211 , n56226 );
or ( n56229 , n56214 , n56227 , n56228 );
and ( n56230 , n56179 , n56229 );
xor ( n56231 , n55952 , n55956 );
xor ( n56232 , n56231 , n55959 );
and ( n56233 , n56229 , n56232 );
and ( n56234 , n56179 , n56232 );
or ( n56235 , n56230 , n56233 , n56234 );
and ( n56236 , n53785 , n52617 );
and ( n56237 , n53652 , n52615 );
nor ( n56238 , n56236 , n56237 );
xnor ( n56239 , n56238 , n52558 );
and ( n56240 , n53895 , n52540 );
and ( n56241 , n53783 , n52538 );
nor ( n56242 , n56240 , n56241 );
xnor ( n56243 , n56242 , n52424 );
and ( n56244 , n56239 , n56243 );
xor ( n56245 , n55776 , n55780 );
xor ( n56246 , n56245 , n55783 );
and ( n56247 , n56243 , n56246 );
and ( n56248 , n56239 , n56246 );
or ( n56249 , n56244 , n56247 , n56248 );
and ( n56250 , n52952 , n53293 );
and ( n56251 , n52954 , n53291 );
nor ( n56252 , n56250 , n56251 );
xnor ( n56253 , n56252 , n52963 );
and ( n56254 , n56249 , n56253 );
and ( n56255 , n53499 , n52886 );
and ( n56256 , n53322 , n52884 );
nor ( n56257 , n56255 , n56256 );
xnor ( n56258 , n56257 , n52657 );
and ( n56259 , n56253 , n56258 );
and ( n56260 , n56249 , n56258 );
or ( n56261 , n56254 , n56259 , n56260 );
and ( n56262 , n52431 , n54285 );
and ( n56263 , n52371 , n54283 );
nor ( n56264 , n56262 , n56263 );
xnor ( n56265 , n56264 , n53794 );
and ( n56266 , n56261 , n56265 );
xor ( n56267 , n55998 , n56002 );
xor ( n56268 , n56267 , n56007 );
and ( n56269 , n56265 , n56268 );
and ( n56270 , n56261 , n56268 );
or ( n56271 , n56266 , n56269 , n56270 );
and ( n56272 , n52186 , n55033 );
and ( n56273 , n52159 , n55030 );
nor ( n56274 , n56272 , n56273 );
xnor ( n56275 , n56274 , n53885 );
and ( n56276 , n56271 , n56275 );
and ( n56277 , n52271 , n54693 );
and ( n56278 , n52220 , n54691 );
nor ( n56279 , n56277 , n56278 );
xnor ( n56280 , n56279 , n53892 );
and ( n56281 , n56275 , n56280 );
and ( n56282 , n56271 , n56280 );
or ( n56283 , n56276 , n56281 , n56282 );
and ( n56284 , n56218 , n56222 );
and ( n56285 , n56222 , n56225 );
and ( n56286 , n56218 , n56225 );
or ( n56287 , n56284 , n56285 , n56286 );
and ( n56288 , n56283 , n56287 );
xor ( n56289 , n55974 , n55978 );
xor ( n56290 , n56289 , n55981 );
and ( n56291 , n56287 , n56290 );
and ( n56292 , n56283 , n56290 );
or ( n56293 , n56288 , n56291 , n56292 );
and ( n56294 , n56235 , n56293 );
xor ( n56295 , n55984 , n56040 );
xor ( n56296 , n56295 , n56043 );
and ( n56297 , n56293 , n56296 );
and ( n56298 , n56235 , n56296 );
or ( n56299 , n56294 , n56297 , n56298 );
xor ( n56300 , n55867 , n55869 );
xor ( n56301 , n56300 , n55872 );
and ( n56302 , n56299 , n56301 );
xor ( n56303 , n55970 , n56046 );
xor ( n56304 , n56303 , n56049 );
and ( n56305 , n56301 , n56304 );
and ( n56306 , n56299 , n56304 );
or ( n56307 , n56302 , n56305 , n56306 );
xor ( n56308 , n56052 , n56054 );
xor ( n56309 , n56308 , n56057 );
and ( n56310 , n56307 , n56309 );
xor ( n56311 , n56299 , n56301 );
xor ( n56312 , n56311 , n56304 );
and ( n56313 , n53652 , n52886 );
and ( n56314 , n53644 , n52884 );
nor ( n56315 , n56313 , n56314 );
xnor ( n56316 , n56315 , n52657 );
and ( n56317 , n54078 , n52540 );
and ( n56318 , n53895 , n52538 );
nor ( n56319 , n56317 , n56318 );
xnor ( n56320 , n56319 , n52424 );
and ( n56321 , n56316 , n56320 );
xor ( n56322 , n56122 , n56126 );
xor ( n56323 , n56322 , n56131 );
and ( n56324 , n56320 , n56323 );
and ( n56325 , n56316 , n56323 );
or ( n56326 , n56321 , n56324 , n56325 );
and ( n56327 , n55769 , n52121 );
and ( n56328 , n55720 , n52119 );
nor ( n56329 , n56327 , n56328 );
xnor ( n56330 , n56329 , n52087 );
and ( n56331 , n56071 , n52092 );
and ( n56332 , n56073 , n52090 );
nor ( n56333 , n56331 , n56332 );
xnor ( n56334 , n56333 , n52072 );
and ( n56335 , n56330 , n56334 );
buf ( n56336 , n51717 );
and ( n56337 , n56336 , n52059 );
buf ( n56338 , n51716 );
and ( n56339 , n56338 , n52057 );
nor ( n56340 , n56337 , n56339 );
not ( n56341 , n56340 );
and ( n56342 , n56334 , n56341 );
and ( n56343 , n56330 , n56341 );
or ( n56344 , n56335 , n56342 , n56343 );
and ( n56345 , n56073 , n52092 );
and ( n56346 , n55769 , n52090 );
nor ( n56347 , n56345 , n56346 );
xnor ( n56348 , n56347 , n52072 );
and ( n56349 , n56344 , n56348 );
and ( n56350 , n56338 , n52059 );
and ( n56351 , n56071 , n52057 );
nor ( n56352 , n56350 , n56351 );
not ( n56353 , n56352 );
and ( n56354 , n56348 , n56353 );
and ( n56355 , n56344 , n56353 );
or ( n56356 , n56349 , n56354 , n56355 );
and ( n56357 , n55661 , n52121 );
and ( n56358 , n55406 , n52119 );
nor ( n56359 , n56357 , n56358 );
xnor ( n56360 , n56359 , n52087 );
and ( n56361 , n56356 , n56360 );
xor ( n56362 , n56065 , n56069 );
xor ( n56363 , n56362 , n56076 );
and ( n56364 , n56360 , n56363 );
and ( n56365 , n56356 , n56363 );
or ( n56366 , n56361 , n56364 , n56365 );
and ( n56367 , n54715 , n52346 );
and ( n56368 , n54466 , n52344 );
nor ( n56369 , n56367 , n56368 );
xnor ( n56370 , n56369 , n52300 );
and ( n56371 , n56366 , n56370 );
xor ( n56372 , n56110 , n56114 );
xor ( n56373 , n56372 , n56119 );
and ( n56374 , n56370 , n56373 );
and ( n56375 , n56366 , n56373 );
or ( n56376 , n56371 , n56374 , n56375 );
and ( n56377 , n53783 , n52617 );
and ( n56378 , n53785 , n52615 );
nor ( n56379 , n56377 , n56378 );
xnor ( n56380 , n56379 , n52558 );
and ( n56381 , n56376 , n56380 );
xor ( n56382 , n56091 , n56095 );
xor ( n56383 , n56382 , n56098 );
and ( n56384 , n56380 , n56383 );
and ( n56385 , n56376 , n56383 );
or ( n56386 , n56381 , n56384 , n56385 );
and ( n56387 , n56326 , n56386 );
and ( n56388 , n52954 , n53455 );
and ( n56389 , n52829 , n53453 );
nor ( n56390 , n56388 , n56389 );
xnor ( n56391 , n56390 , n53159 );
and ( n56392 , n56386 , n56391 );
and ( n56393 , n56326 , n56391 );
or ( n56394 , n56387 , n56392 , n56393 );
and ( n56395 , n53150 , n53293 );
and ( n56396 , n52952 , n53291 );
nor ( n56397 , n56395 , n56396 );
xnor ( n56398 , n56397 , n52963 );
and ( n56399 , n53322 , n53021 );
and ( n56400 , n53148 , n53019 );
nor ( n56401 , n56399 , n56400 );
xnor ( n56402 , n56401 , n52839 );
and ( n56403 , n56398 , n56402 );
xor ( n56404 , n56239 , n56243 );
xor ( n56405 , n56404 , n56246 );
and ( n56406 , n56402 , n56405 );
and ( n56407 , n56398 , n56405 );
or ( n56408 , n56403 , n56406 , n56407 );
and ( n56409 , n56394 , n56408 );
xor ( n56410 , n56192 , n56196 );
xor ( n56411 , n56410 , n56199 );
and ( n56412 , n56408 , n56411 );
and ( n56413 , n56394 , n56411 );
or ( n56414 , n56409 , n56412 , n56413 );
and ( n56415 , n52220 , n55033 );
and ( n56416 , n52186 , n55030 );
nor ( n56417 , n56415 , n56416 );
xnor ( n56418 , n56417 , n53885 );
and ( n56419 , n56414 , n56418 );
xor ( n56420 , n56261 , n56265 );
xor ( n56421 , n56420 , n56268 );
and ( n56422 , n56418 , n56421 );
and ( n56423 , n56414 , n56421 );
or ( n56424 , n56419 , n56422 , n56423 );
xor ( n56425 , n56271 , n56275 );
xor ( n56426 , n56425 , n56280 );
and ( n56427 , n56424 , n56426 );
xor ( n56428 , n56169 , n56173 );
xor ( n56429 , n56428 , n56176 );
and ( n56430 , n56426 , n56429 );
and ( n56431 , n56424 , n56429 );
or ( n56432 , n56427 , n56430 , n56431 );
xor ( n56433 , n56283 , n56287 );
xor ( n56434 , n56433 , n56290 );
and ( n56435 , n56432 , n56434 );
xor ( n56436 , n56030 , n56034 );
xor ( n56437 , n56436 , n56037 );
and ( n56438 , n56434 , n56437 );
and ( n56439 , n56432 , n56437 );
or ( n56440 , n56435 , n56438 , n56439 );
xor ( n56441 , n55962 , n55964 );
xor ( n56442 , n56441 , n55967 );
and ( n56443 , n56440 , n56442 );
xor ( n56444 , n56235 , n56293 );
xor ( n56445 , n56444 , n56296 );
and ( n56446 , n56442 , n56445 );
and ( n56447 , n56440 , n56445 );
or ( n56448 , n56443 , n56446 , n56447 );
and ( n56449 , n56312 , n56448 );
xor ( n56450 , n56440 , n56442 );
xor ( n56451 , n56450 , n56445 );
and ( n56452 , n52371 , n54693 );
and ( n56453 , n52307 , n54691 );
nor ( n56454 , n56452 , n56453 );
xnor ( n56455 , n56454 , n53892 );
and ( n56456 , n52639 , n53972 );
and ( n56457 , n52565 , n53970 );
nor ( n56458 , n56456 , n56457 );
xnor ( n56459 , n56458 , n53662 );
and ( n56460 , n56455 , n56459 );
and ( n56461 , n52718 , n53739 );
and ( n56462 , n52664 , n53737 );
nor ( n56463 , n56461 , n56462 );
xnor ( n56464 , n56463 , n53315 );
and ( n56465 , n56459 , n56464 );
and ( n56466 , n56455 , n56464 );
or ( n56467 , n56460 , n56465 , n56466 );
and ( n56468 , n52439 , n54285 );
and ( n56469 , n52431 , n54283 );
nor ( n56470 , n56468 , n56469 );
xnor ( n56471 , n56470 , n53794 );
xor ( n56472 , n56249 , n56253 );
xor ( n56473 , n56472 , n56258 );
and ( n56474 , n56471 , n56473 );
xor ( n56475 , n56147 , n56151 );
xor ( n56476 , n56475 , n56154 );
and ( n56477 , n56473 , n56476 );
and ( n56478 , n56471 , n56476 );
or ( n56479 , n56474 , n56477 , n56478 );
and ( n56480 , n56467 , n56479 );
xor ( n56481 , n56157 , n56161 );
xor ( n56482 , n56481 , n56166 );
and ( n56483 , n56479 , n56482 );
and ( n56484 , n56467 , n56482 );
or ( n56485 , n56480 , n56483 , n56484 );
and ( n56486 , n56073 , n52121 );
and ( n56487 , n55769 , n52119 );
nor ( n56488 , n56486 , n56487 );
xnor ( n56489 , n56488 , n52087 );
and ( n56490 , n56338 , n52092 );
and ( n56491 , n56071 , n52090 );
nor ( n56492 , n56490 , n56491 );
xnor ( n56493 , n56492 , n52072 );
and ( n56494 , n56489 , n56493 );
buf ( n56495 , n51718 );
and ( n56496 , n56495 , n52059 );
and ( n56497 , n56336 , n52057 );
nor ( n56498 , n56496 , n56497 );
not ( n56499 , n56498 );
and ( n56500 , n56493 , n56499 );
and ( n56501 , n56489 , n56499 );
or ( n56502 , n56494 , n56500 , n56501 );
and ( n56503 , n55365 , n52318 );
and ( n56504 , n55199 , n52316 );
nor ( n56505 , n56503 , n56504 );
xnor ( n56506 , n56505 , n52213 );
and ( n56507 , n56502 , n56506 );
and ( n56508 , n55661 , n52170 );
and ( n56509 , n55406 , n52168 );
nor ( n56510 , n56508 , n56509 );
xnor ( n56511 , n56510 , n52152 );
and ( n56512 , n56506 , n56511 );
and ( n56513 , n56502 , n56511 );
or ( n56514 , n56507 , n56512 , n56513 );
and ( n56515 , n54885 , n52346 );
and ( n56516 , n54767 , n52344 );
nor ( n56517 , n56515 , n56516 );
xnor ( n56518 , n56517 , n52300 );
and ( n56519 , n56514 , n56518 );
xor ( n56520 , n56344 , n56348 );
xor ( n56521 , n56520 , n56353 );
and ( n56522 , n56518 , n56521 );
and ( n56523 , n56514 , n56521 );
or ( n56524 , n56519 , n56522 , n56523 );
and ( n56525 , n54078 , n52617 );
and ( n56526 , n53895 , n52615 );
nor ( n56527 , n56525 , n56526 );
xnor ( n56528 , n56527 , n52558 );
and ( n56529 , n56524 , n56528 );
xor ( n56530 , n56356 , n56360 );
xor ( n56531 , n56530 , n56363 );
and ( n56532 , n56528 , n56531 );
and ( n56533 , n56524 , n56531 );
or ( n56534 , n56529 , n56532 , n56533 );
and ( n56535 , n53322 , n53293 );
and ( n56536 , n53148 , n53291 );
nor ( n56537 , n56535 , n56536 );
xnor ( n56538 , n56537 , n52963 );
and ( n56539 , n56534 , n56538 );
and ( n56540 , n55199 , n52318 );
and ( n56541 , n55055 , n52316 );
nor ( n56542 , n56540 , n56541 );
xnor ( n56543 , n56542 , n52213 );
and ( n56544 , n55406 , n52170 );
and ( n56545 , n55365 , n52168 );
nor ( n56546 , n56544 , n56545 );
xnor ( n56547 , n56546 , n52152 );
and ( n56548 , n56543 , n56547 );
and ( n56549 , n55720 , n52121 );
and ( n56550 , n55661 , n52119 );
nor ( n56551 , n56549 , n56550 );
xnor ( n56552 , n56551 , n52087 );
and ( n56553 , n56547 , n56552 );
and ( n56554 , n56543 , n56552 );
or ( n56555 , n56548 , n56553 , n56554 );
and ( n56556 , n54767 , n52346 );
and ( n56557 , n54715 , n52344 );
nor ( n56558 , n56556 , n56557 );
xnor ( n56559 , n56558 , n52300 );
and ( n56560 , n56555 , n56559 );
and ( n56561 , n55055 , n52318 );
and ( n56562 , n54885 , n52316 );
nor ( n56563 , n56561 , n56562 );
xnor ( n56564 , n56563 , n52213 );
and ( n56565 , n56559 , n56564 );
and ( n56566 , n56555 , n56564 );
or ( n56567 , n56560 , n56565 , n56566 );
and ( n56568 , n54364 , n52540 );
and ( n56569 , n54078 , n52538 );
nor ( n56570 , n56568 , n56569 );
xnor ( n56571 , n56570 , n52424 );
xor ( n56572 , n56567 , n56571 );
xor ( n56573 , n56079 , n56083 );
xor ( n56574 , n56573 , n56088 );
xor ( n56575 , n56572 , n56574 );
and ( n56576 , n56538 , n56575 );
and ( n56577 , n56534 , n56575 );
or ( n56578 , n56539 , n56576 , n56577 );
and ( n56579 , n52952 , n53455 );
and ( n56580 , n52954 , n53453 );
nor ( n56581 , n56579 , n56580 );
xnor ( n56582 , n56581 , n53159 );
and ( n56583 , n56578 , n56582 );
xor ( n56584 , n56376 , n56380 );
xor ( n56585 , n56584 , n56383 );
and ( n56586 , n56582 , n56585 );
and ( n56587 , n56578 , n56585 );
or ( n56588 , n56583 , n56586 , n56587 );
and ( n56589 , n52431 , n54693 );
and ( n56590 , n52371 , n54691 );
nor ( n56591 , n56589 , n56590 );
xnor ( n56592 , n56591 , n53892 );
and ( n56593 , n56588 , n56592 );
and ( n56594 , n52565 , n54285 );
and ( n56595 , n52439 , n54283 );
nor ( n56596 , n56594 , n56595 );
xnor ( n56597 , n56596 , n53794 );
and ( n56598 , n56592 , n56597 );
and ( n56599 , n56588 , n56597 );
or ( n56600 , n56593 , n56598 , n56599 );
and ( n56601 , n52664 , n53972 );
and ( n56602 , n52639 , n53970 );
nor ( n56603 , n56601 , n56602 );
xnor ( n56604 , n56603 , n53662 );
xor ( n56605 , n56326 , n56386 );
xor ( n56606 , n56605 , n56391 );
and ( n56607 , n56604 , n56606 );
xor ( n56608 , n56398 , n56402 );
xor ( n56609 , n56608 , n56405 );
and ( n56610 , n56606 , n56609 );
and ( n56611 , n56604 , n56609 );
or ( n56612 , n56607 , n56610 , n56611 );
and ( n56613 , n56600 , n56612 );
xor ( n56614 , n56455 , n56459 );
xor ( n56615 , n56614 , n56464 );
and ( n56616 , n56612 , n56615 );
and ( n56617 , n56600 , n56615 );
or ( n56618 , n56613 , n56616 , n56617 );
and ( n56619 , n56567 , n56571 );
and ( n56620 , n56571 , n56574 );
and ( n56621 , n56567 , n56574 );
or ( n56622 , n56619 , n56620 , n56621 );
and ( n56623 , n53148 , n53293 );
and ( n56624 , n53150 , n53291 );
nor ( n56625 , n56623 , n56624 );
xnor ( n56626 , n56625 , n52963 );
and ( n56627 , n56622 , n56626 );
and ( n56628 , n53499 , n53021 );
and ( n56629 , n53322 , n53019 );
nor ( n56630 , n56628 , n56629 );
xnor ( n56631 , n56630 , n52839 );
and ( n56632 , n56626 , n56631 );
and ( n56633 , n56622 , n56631 );
or ( n56634 , n56627 , n56632 , n56633 );
and ( n56635 , n53785 , n52886 );
and ( n56636 , n53652 , n52884 );
nor ( n56637 , n56635 , n56636 );
xnor ( n56638 , n56637 , n52657 );
and ( n56639 , n53895 , n52617 );
and ( n56640 , n53783 , n52615 );
nor ( n56641 , n56639 , n56640 );
xnor ( n56642 , n56641 , n52558 );
and ( n56643 , n56638 , n56642 );
xor ( n56644 , n56366 , n56370 );
xor ( n56645 , n56644 , n56373 );
and ( n56646 , n56642 , n56645 );
and ( n56647 , n56638 , n56645 );
or ( n56648 , n56643 , n56646 , n56647 );
and ( n56649 , n52829 , n53739 );
and ( n56650 , n52809 , n53737 );
nor ( n56651 , n56649 , n56650 );
xnor ( n56652 , n56651 , n53315 );
and ( n56653 , n56648 , n56652 );
xor ( n56654 , n56316 , n56320 );
xor ( n56655 , n56654 , n56323 );
and ( n56656 , n56652 , n56655 );
and ( n56657 , n56648 , n56655 );
or ( n56658 , n56653 , n56656 , n56657 );
and ( n56659 , n56634 , n56658 );
xor ( n56660 , n56101 , n56105 );
xor ( n56661 , n56660 , n56144 );
and ( n56662 , n56658 , n56661 );
and ( n56663 , n56634 , n56661 );
or ( n56664 , n56659 , n56662 , n56663 );
and ( n56665 , n52271 , n55033 );
and ( n56666 , n52220 , n55030 );
nor ( n56667 , n56665 , n56666 );
xnor ( n56668 , n56667 , n53885 );
and ( n56669 , n56664 , n56668 );
xor ( n56670 , n56394 , n56408 );
xor ( n56671 , n56670 , n56411 );
and ( n56672 , n56668 , n56671 );
and ( n56673 , n56664 , n56671 );
or ( n56674 , n56669 , n56672 , n56673 );
and ( n56675 , n56618 , n56674 );
xor ( n56676 , n56183 , n56187 );
xor ( n56677 , n56676 , n56208 );
and ( n56678 , n56674 , n56677 );
and ( n56679 , n56618 , n56677 );
or ( n56680 , n56675 , n56678 , n56679 );
and ( n56681 , n56485 , n56680 );
xor ( n56682 , n56211 , n56213 );
xor ( n56683 , n56682 , n56226 );
and ( n56684 , n56680 , n56683 );
and ( n56685 , n56485 , n56683 );
or ( n56686 , n56681 , n56684 , n56685 );
xor ( n56687 , n56179 , n56229 );
xor ( n56688 , n56687 , n56232 );
and ( n56689 , n56686 , n56688 );
xor ( n56690 , n56432 , n56434 );
xor ( n56691 , n56690 , n56437 );
and ( n56692 , n56688 , n56691 );
and ( n56693 , n56686 , n56691 );
or ( n56694 , n56689 , n56692 , n56693 );
and ( n56695 , n56451 , n56694 );
xor ( n56696 , n56686 , n56688 );
xor ( n56697 , n56696 , n56691 );
and ( n56698 , n52307 , n55033 );
and ( n56699 , n52271 , n55030 );
nor ( n56700 , n56698 , n56699 );
xnor ( n56701 , n56700 , n53885 );
and ( n56702 , n52809 , n53739 );
and ( n56703 , n52718 , n53737 );
nor ( n56704 , n56702 , n56703 );
xnor ( n56705 , n56704 , n53315 );
and ( n56706 , n56701 , n56705 );
xor ( n56707 , n56634 , n56658 );
xor ( n56708 , n56707 , n56661 );
and ( n56709 , n56705 , n56708 );
and ( n56710 , n56701 , n56708 );
or ( n56711 , n56706 , n56709 , n56710 );
xor ( n56712 , n56664 , n56668 );
xor ( n56713 , n56712 , n56671 );
and ( n56714 , n56711 , n56713 );
xor ( n56715 , n56471 , n56473 );
xor ( n56716 , n56715 , n56476 );
and ( n56717 , n56713 , n56716 );
and ( n56718 , n56711 , n56716 );
or ( n56719 , n56714 , n56717 , n56718 );
xor ( n56720 , n56467 , n56479 );
xor ( n56721 , n56720 , n56482 );
and ( n56722 , n56719 , n56721 );
xor ( n56723 , n56414 , n56418 );
xor ( n56724 , n56723 , n56421 );
and ( n56725 , n56721 , n56724 );
and ( n56726 , n56719 , n56724 );
or ( n56727 , n56722 , n56725 , n56726 );
xor ( n56728 , n56424 , n56426 );
xor ( n56729 , n56728 , n56429 );
and ( n56730 , n56727 , n56729 );
xor ( n56731 , n56485 , n56680 );
xor ( n56732 , n56731 , n56683 );
and ( n56733 , n56729 , n56732 );
and ( n56734 , n56727 , n56732 );
or ( n56735 , n56730 , n56733 , n56734 );
and ( n56736 , n56697 , n56735 );
xor ( n56737 , n56727 , n56729 );
xor ( n56738 , n56737 , n56732 );
and ( n56739 , n52371 , n55033 );
and ( n56740 , n52307 , n55030 );
nor ( n56741 , n56739 , n56740 );
xnor ( n56742 , n56741 , n53885 );
and ( n56743 , n52439 , n54693 );
and ( n56744 , n52431 , n54691 );
nor ( n56745 , n56743 , n56744 );
xnor ( n56746 , n56745 , n53892 );
and ( n56747 , n56742 , n56746 );
and ( n56748 , n52639 , n54285 );
and ( n56749 , n52565 , n54283 );
nor ( n56750 , n56748 , n56749 );
xnor ( n56751 , n56750 , n53794 );
and ( n56752 , n56746 , n56751 );
and ( n56753 , n56742 , n56751 );
or ( n56754 , n56747 , n56752 , n56753 );
xor ( n56755 , n56588 , n56592 );
xor ( n56756 , n56755 , n56597 );
and ( n56757 , n56754 , n56756 );
xor ( n56758 , n56701 , n56705 );
xor ( n56759 , n56758 , n56708 );
and ( n56760 , n56756 , n56759 );
and ( n56761 , n56754 , n56759 );
or ( n56762 , n56757 , n56760 , n56761 );
and ( n56763 , n53783 , n52886 );
and ( n56764 , n53785 , n52884 );
nor ( n56765 , n56763 , n56764 );
xnor ( n56766 , n56765 , n52657 );
and ( n56767 , n54466 , n52540 );
and ( n56768 , n54364 , n52538 );
nor ( n56769 , n56767 , n56768 );
xnor ( n56770 , n56769 , n52424 );
and ( n56771 , n56766 , n56770 );
xor ( n56772 , n56555 , n56559 );
xor ( n56773 , n56772 , n56564 );
and ( n56774 , n56770 , n56773 );
and ( n56775 , n56766 , n56773 );
or ( n56776 , n56771 , n56774 , n56775 );
and ( n56777 , n53150 , n53455 );
and ( n56778 , n52952 , n53453 );
nor ( n56779 , n56777 , n56778 );
xnor ( n56780 , n56779 , n53159 );
and ( n56781 , n56776 , n56780 );
and ( n56782 , n53644 , n53021 );
and ( n56783 , n53499 , n53019 );
nor ( n56784 , n56782 , n56783 );
xnor ( n56785 , n56784 , n52839 );
and ( n56786 , n56780 , n56785 );
and ( n56787 , n56776 , n56785 );
or ( n56788 , n56781 , n56786 , n56787 );
xor ( n56789 , n56622 , n56626 );
xor ( n56790 , n56789 , n56631 );
and ( n56791 , n56788 , n56790 );
xor ( n56792 , n56648 , n56652 );
xor ( n56793 , n56792 , n56655 );
and ( n56794 , n56790 , n56793 );
and ( n56795 , n56788 , n56793 );
or ( n56796 , n56791 , n56794 , n56795 );
and ( n56797 , n56071 , n52121 );
and ( n56798 , n56073 , n52119 );
nor ( n56799 , n56797 , n56798 );
xnor ( n56800 , n56799 , n52087 );
and ( n56801 , n56336 , n52092 );
and ( n56802 , n56338 , n52090 );
nor ( n56803 , n56801 , n56802 );
xnor ( n56804 , n56803 , n52072 );
and ( n56805 , n56800 , n56804 );
buf ( n56806 , n51719 );
and ( n56807 , n56806 , n52059 );
and ( n56808 , n56495 , n52057 );
nor ( n56809 , n56807 , n56808 );
not ( n56810 , n56809 );
and ( n56811 , n56804 , n56810 );
and ( n56812 , n56800 , n56810 );
or ( n56813 , n56805 , n56811 , n56812 );
and ( n56814 , n55406 , n52318 );
and ( n56815 , n55365 , n52316 );
nor ( n56816 , n56814 , n56815 );
xnor ( n56817 , n56816 , n52213 );
and ( n56818 , n56813 , n56817 );
and ( n56819 , n55720 , n52170 );
and ( n56820 , n55661 , n52168 );
nor ( n56821 , n56819 , n56820 );
xnor ( n56822 , n56821 , n52152 );
and ( n56823 , n56817 , n56822 );
and ( n56824 , n56813 , n56822 );
or ( n56825 , n56818 , n56823 , n56824 );
and ( n56826 , n55055 , n52346 );
and ( n56827 , n54885 , n52344 );
nor ( n56828 , n56826 , n56827 );
xnor ( n56829 , n56828 , n52300 );
and ( n56830 , n56825 , n56829 );
xor ( n56831 , n56330 , n56334 );
xor ( n56832 , n56831 , n56341 );
and ( n56833 , n56829 , n56832 );
and ( n56834 , n56825 , n56832 );
or ( n56835 , n56830 , n56833 , n56834 );
and ( n56836 , n54715 , n52540 );
and ( n56837 , n54466 , n52538 );
nor ( n56838 , n56836 , n56837 );
xnor ( n56839 , n56838 , n52424 );
and ( n56840 , n56835 , n56839 );
xor ( n56841 , n56543 , n56547 );
xor ( n56842 , n56841 , n56552 );
and ( n56843 , n56839 , n56842 );
and ( n56844 , n56835 , n56842 );
or ( n56845 , n56840 , n56843 , n56844 );
and ( n56846 , n56073 , n52170 );
and ( n56847 , n55769 , n52168 );
nor ( n56848 , n56846 , n56847 );
xnor ( n56849 , n56848 , n52152 );
and ( n56850 , n56495 , n52092 );
and ( n56851 , n56336 , n52090 );
nor ( n56852 , n56850 , n56851 );
xnor ( n56853 , n56852 , n52072 );
and ( n56854 , n56849 , n56853 );
buf ( n56855 , n51720 );
and ( n56856 , n56855 , n52059 );
and ( n56857 , n56806 , n52057 );
nor ( n56858 , n56856 , n56857 );
not ( n56859 , n56858 );
and ( n56860 , n56853 , n56859 );
and ( n56861 , n56849 , n56859 );
or ( n56862 , n56854 , n56860 , n56861 );
and ( n56863 , n55769 , n52170 );
and ( n56864 , n55720 , n52168 );
nor ( n56865 , n56863 , n56864 );
xnor ( n56866 , n56865 , n52152 );
and ( n56867 , n56862 , n56866 );
xor ( n56868 , n56800 , n56804 );
xor ( n56869 , n56868 , n56810 );
and ( n56870 , n56866 , n56869 );
and ( n56871 , n56862 , n56869 );
or ( n56872 , n56867 , n56870 , n56871 );
and ( n56873 , n55199 , n52346 );
and ( n56874 , n55055 , n52344 );
nor ( n56875 , n56873 , n56874 );
xnor ( n56876 , n56875 , n52300 );
and ( n56877 , n56872 , n56876 );
xor ( n56878 , n56489 , n56493 );
xor ( n56879 , n56878 , n56499 );
and ( n56880 , n56876 , n56879 );
and ( n56881 , n56872 , n56879 );
or ( n56882 , n56877 , n56880 , n56881 );
and ( n56883 , n54767 , n52540 );
and ( n56884 , n54715 , n52538 );
nor ( n56885 , n56883 , n56884 );
xnor ( n56886 , n56885 , n52424 );
and ( n56887 , n56882 , n56886 );
xor ( n56888 , n56502 , n56506 );
xor ( n56889 , n56888 , n56511 );
and ( n56890 , n56886 , n56889 );
and ( n56891 , n56882 , n56889 );
or ( n56892 , n56887 , n56890 , n56891 );
and ( n56893 , n54364 , n52617 );
and ( n56894 , n54078 , n52615 );
nor ( n56895 , n56893 , n56894 );
xnor ( n56896 , n56895 , n52558 );
and ( n56897 , n56892 , n56896 );
xor ( n56898 , n56514 , n56518 );
xor ( n56899 , n56898 , n56521 );
and ( n56900 , n56896 , n56899 );
and ( n56901 , n56892 , n56899 );
or ( n56902 , n56897 , n56900 , n56901 );
and ( n56903 , n56845 , n56902 );
and ( n56904 , n53652 , n53021 );
and ( n56905 , n53644 , n53019 );
nor ( n56906 , n56904 , n56905 );
xnor ( n56907 , n56906 , n52839 );
and ( n56908 , n56902 , n56907 );
and ( n56909 , n56845 , n56907 );
or ( n56910 , n56903 , n56908 , n56909 );
and ( n56911 , n52954 , n53739 );
and ( n56912 , n52829 , n53737 );
nor ( n56913 , n56911 , n56912 );
xnor ( n56914 , n56913 , n53315 );
and ( n56915 , n56910 , n56914 );
xor ( n56916 , n56638 , n56642 );
xor ( n56917 , n56916 , n56645 );
and ( n56918 , n56914 , n56917 );
and ( n56919 , n56910 , n56917 );
or ( n56920 , n56915 , n56918 , n56919 );
and ( n56921 , n52718 , n53972 );
and ( n56922 , n52664 , n53970 );
nor ( n56923 , n56921 , n56922 );
xnor ( n56924 , n56923 , n53662 );
and ( n56925 , n56920 , n56924 );
xor ( n56926 , n56578 , n56582 );
xor ( n56927 , n56926 , n56585 );
and ( n56928 , n56924 , n56927 );
and ( n56929 , n56920 , n56927 );
or ( n56930 , n56925 , n56928 , n56929 );
and ( n56931 , n56796 , n56930 );
xor ( n56932 , n56604 , n56606 );
xor ( n56933 , n56932 , n56609 );
and ( n56934 , n56930 , n56933 );
and ( n56935 , n56796 , n56933 );
or ( n56936 , n56931 , n56934 , n56935 );
and ( n56937 , n56762 , n56936 );
xor ( n56938 , n56600 , n56612 );
xor ( n56939 , n56938 , n56615 );
and ( n56940 , n56936 , n56939 );
and ( n56941 , n56762 , n56939 );
or ( n56942 , n56937 , n56940 , n56941 );
xor ( n56943 , n56719 , n56721 );
xor ( n56944 , n56943 , n56724 );
and ( n56945 , n56942 , n56944 );
xor ( n56946 , n56618 , n56674 );
xor ( n56947 , n56946 , n56677 );
and ( n56948 , n56944 , n56947 );
and ( n56949 , n56942 , n56947 );
or ( n56950 , n56945 , n56948 , n56949 );
and ( n56951 , n56738 , n56950 );
xor ( n56952 , n56942 , n56944 );
xor ( n56953 , n56952 , n56947 );
and ( n56954 , n53785 , n53021 );
and ( n56955 , n53652 , n53019 );
nor ( n56956 , n56954 , n56955 );
xnor ( n56957 , n56956 , n52839 );
and ( n56958 , n53895 , n52886 );
and ( n56959 , n53783 , n52884 );
nor ( n56960 , n56958 , n56959 );
xnor ( n56961 , n56960 , n52657 );
and ( n56962 , n56957 , n56961 );
xor ( n56963 , n56835 , n56839 );
xor ( n56964 , n56963 , n56842 );
and ( n56965 , n56961 , n56964 );
and ( n56966 , n56957 , n56964 );
or ( n56967 , n56962 , n56965 , n56966 );
and ( n56968 , n52952 , n53739 );
and ( n56969 , n52954 , n53737 );
nor ( n56970 , n56968 , n56969 );
xnor ( n56971 , n56970 , n53315 );
and ( n56972 , n56967 , n56971 );
xor ( n56973 , n56766 , n56770 );
xor ( n56974 , n56973 , n56773 );
and ( n56975 , n56971 , n56974 );
and ( n56976 , n56967 , n56974 );
or ( n56977 , n56972 , n56975 , n56976 );
and ( n56978 , n53148 , n53455 );
and ( n56979 , n53150 , n53453 );
nor ( n56980 , n56978 , n56979 );
xnor ( n56981 , n56980 , n53159 );
and ( n56982 , n53499 , n53293 );
and ( n56983 , n53322 , n53291 );
nor ( n56984 , n56982 , n56983 );
xnor ( n56985 , n56984 , n52963 );
and ( n56986 , n56981 , n56985 );
xor ( n56987 , n56524 , n56528 );
xor ( n56988 , n56987 , n56531 );
and ( n56989 , n56985 , n56988 );
and ( n56990 , n56981 , n56988 );
or ( n56991 , n56986 , n56989 , n56990 );
and ( n56992 , n56977 , n56991 );
xor ( n56993 , n56534 , n56538 );
xor ( n56994 , n56993 , n56575 );
and ( n56995 , n56991 , n56994 );
and ( n56996 , n56977 , n56994 );
or ( n56997 , n56992 , n56995 , n56996 );
and ( n56998 , n52664 , n54285 );
and ( n56999 , n52639 , n54283 );
nor ( n57000 , n56998 , n56999 );
xnor ( n57001 , n57000 , n53794 );
and ( n57002 , n52809 , n53972 );
and ( n57003 , n52718 , n53970 );
nor ( n57004 , n57002 , n57003 );
xnor ( n57005 , n57004 , n53662 );
and ( n57006 , n57001 , n57005 );
xor ( n57007 , n56910 , n56914 );
xor ( n57008 , n57007 , n56917 );
and ( n57009 , n57005 , n57008 );
and ( n57010 , n57001 , n57008 );
or ( n57011 , n57006 , n57009 , n57010 );
and ( n57012 , n56997 , n57011 );
xor ( n57013 , n56788 , n56790 );
xor ( n57014 , n57013 , n56793 );
and ( n57015 , n57011 , n57014 );
and ( n57016 , n56997 , n57014 );
or ( n57017 , n57012 , n57015 , n57016 );
and ( n57018 , n56336 , n52121 );
and ( n57019 , n56338 , n52119 );
nor ( n57020 , n57018 , n57019 );
xnor ( n57021 , n57020 , n52087 );
and ( n57022 , n56806 , n52092 );
and ( n57023 , n56495 , n52090 );
nor ( n57024 , n57022 , n57023 );
xnor ( n57025 , n57024 , n52072 );
and ( n57026 , n57021 , n57025 );
buf ( n57027 , n51721 );
and ( n57028 , n57027 , n52059 );
and ( n57029 , n56855 , n52057 );
nor ( n57030 , n57028 , n57029 );
not ( n57031 , n57030 );
and ( n57032 , n57025 , n57031 );
and ( n57033 , n57021 , n57031 );
or ( n57034 , n57026 , n57032 , n57033 );
and ( n57035 , n56338 , n52121 );
and ( n57036 , n56071 , n52119 );
nor ( n57037 , n57035 , n57036 );
xnor ( n57038 , n57037 , n52087 );
and ( n57039 , n57034 , n57038 );
xor ( n57040 , n56849 , n56853 );
xor ( n57041 , n57040 , n56859 );
and ( n57042 , n57038 , n57041 );
and ( n57043 , n57034 , n57041 );
or ( n57044 , n57039 , n57042 , n57043 );
and ( n57045 , n55365 , n52346 );
and ( n57046 , n55199 , n52344 );
nor ( n57047 , n57045 , n57046 );
xnor ( n57048 , n57047 , n52300 );
and ( n57049 , n57044 , n57048 );
and ( n57050 , n55661 , n52318 );
and ( n57051 , n55406 , n52316 );
nor ( n57052 , n57050 , n57051 );
xnor ( n57053 , n57052 , n52213 );
and ( n57054 , n57048 , n57053 );
and ( n57055 , n57044 , n57053 );
or ( n57056 , n57049 , n57054 , n57055 );
and ( n57057 , n54885 , n52540 );
and ( n57058 , n54767 , n52538 );
nor ( n57059 , n57057 , n57058 );
xnor ( n57060 , n57059 , n52424 );
and ( n57061 , n57056 , n57060 );
xor ( n57062 , n56813 , n56817 );
xor ( n57063 , n57062 , n56822 );
and ( n57064 , n57060 , n57063 );
and ( n57065 , n57056 , n57063 );
or ( n57066 , n57061 , n57064 , n57065 );
and ( n57067 , n54078 , n52886 );
and ( n57068 , n53895 , n52884 );
nor ( n57069 , n57067 , n57068 );
xnor ( n57070 , n57069 , n52657 );
and ( n57071 , n57066 , n57070 );
xor ( n57072 , n56825 , n56829 );
xor ( n57073 , n57072 , n56832 );
and ( n57074 , n57070 , n57073 );
and ( n57075 , n57066 , n57073 );
or ( n57076 , n57071 , n57074 , n57075 );
and ( n57077 , n53322 , n53455 );
and ( n57078 , n53148 , n53453 );
nor ( n57079 , n57077 , n57078 );
xnor ( n57080 , n57079 , n53159 );
and ( n57081 , n57076 , n57080 );
and ( n57082 , n53644 , n53293 );
and ( n57083 , n53499 , n53291 );
nor ( n57084 , n57082 , n57083 );
xnor ( n57085 , n57084 , n52963 );
and ( n57086 , n57080 , n57085 );
and ( n57087 , n57076 , n57085 );
or ( n57088 , n57081 , n57086 , n57087 );
and ( n57089 , n52829 , n53972 );
and ( n57090 , n52809 , n53970 );
nor ( n57091 , n57089 , n57090 );
xnor ( n57092 , n57091 , n53662 );
and ( n57093 , n57088 , n57092 );
xor ( n57094 , n56845 , n56902 );
xor ( n57095 , n57094 , n56907 );
and ( n57096 , n57092 , n57095 );
and ( n57097 , n57088 , n57095 );
or ( n57098 , n57093 , n57096 , n57097 );
and ( n57099 , n52431 , n55033 );
and ( n57100 , n52371 , n55030 );
nor ( n57101 , n57099 , n57100 );
xnor ( n57102 , n57101 , n53885 );
and ( n57103 , n57098 , n57102 );
xor ( n57104 , n56776 , n56780 );
xor ( n57105 , n57104 , n56785 );
and ( n57106 , n57102 , n57105 );
and ( n57107 , n57098 , n57105 );
or ( n57108 , n57103 , n57106 , n57107 );
xor ( n57109 , n56742 , n56746 );
xor ( n57110 , n57109 , n56751 );
and ( n57111 , n57108 , n57110 );
xor ( n57112 , n56920 , n56924 );
xor ( n57113 , n57112 , n56927 );
and ( n57114 , n57110 , n57113 );
and ( n57115 , n57108 , n57113 );
or ( n57116 , n57111 , n57114 , n57115 );
and ( n57117 , n57017 , n57116 );
xor ( n57118 , n56796 , n56930 );
xor ( n57119 , n57118 , n56933 );
and ( n57120 , n57116 , n57119 );
and ( n57121 , n57017 , n57119 );
or ( n57122 , n57117 , n57120 , n57121 );
xor ( n57123 , n56762 , n56936 );
xor ( n57124 , n57123 , n56939 );
and ( n57125 , n57122 , n57124 );
xor ( n57126 , n56711 , n56713 );
xor ( n57127 , n57126 , n56716 );
and ( n57128 , n57124 , n57127 );
and ( n57129 , n57122 , n57127 );
or ( n57130 , n57125 , n57128 , n57129 );
and ( n57131 , n56953 , n57130 );
xor ( n57132 , n57122 , n57124 );
xor ( n57133 , n57132 , n57127 );
and ( n57134 , n53652 , n53293 );
and ( n57135 , n53644 , n53291 );
nor ( n57136 , n57134 , n57135 );
xnor ( n57137 , n57136 , n52963 );
and ( n57138 , n54466 , n52617 );
and ( n57139 , n54364 , n52615 );
nor ( n57140 , n57138 , n57139 );
xnor ( n57141 , n57140 , n52558 );
and ( n57142 , n57137 , n57141 );
xor ( n57143 , n56882 , n56886 );
xor ( n57144 , n57143 , n56889 );
and ( n57145 , n57141 , n57144 );
and ( n57146 , n57137 , n57144 );
or ( n57147 , n57142 , n57145 , n57146 );
and ( n57148 , n53150 , n53739 );
and ( n57149 , n52952 , n53737 );
nor ( n57150 , n57148 , n57149 );
xnor ( n57151 , n57150 , n53315 );
and ( n57152 , n57147 , n57151 );
xor ( n57153 , n56892 , n56896 );
xor ( n57154 , n57153 , n56899 );
and ( n57155 , n57151 , n57154 );
and ( n57156 , n57147 , n57154 );
or ( n57157 , n57152 , n57155 , n57156 );
and ( n57158 , n52718 , n54285 );
and ( n57159 , n52664 , n54283 );
nor ( n57160 , n57158 , n57159 );
xnor ( n57161 , n57160 , n53794 );
and ( n57162 , n57157 , n57161 );
xor ( n57163 , n56981 , n56985 );
xor ( n57164 , n57163 , n56988 );
and ( n57165 , n57161 , n57164 );
and ( n57166 , n57157 , n57164 );
or ( n57167 , n57162 , n57165 , n57166 );
and ( n57168 , n52565 , n54693 );
and ( n57169 , n52439 , n54691 );
nor ( n57170 , n57168 , n57169 );
xnor ( n57171 , n57170 , n53892 );
and ( n57172 , n57167 , n57171 );
xor ( n57173 , n56977 , n56991 );
xor ( n57174 , n57173 , n56994 );
and ( n57175 , n57171 , n57174 );
and ( n57176 , n57167 , n57174 );
or ( n57177 , n57172 , n57175 , n57176 );
and ( n57178 , n53148 , n53739 );
and ( n57179 , n53150 , n53737 );
nor ( n57180 , n57178 , n57179 );
xnor ( n57181 , n57180 , n53315 );
and ( n57182 , n53499 , n53455 );
and ( n57183 , n53322 , n53453 );
nor ( n57184 , n57182 , n57183 );
xnor ( n57185 , n57184 , n53159 );
and ( n57186 , n57181 , n57185 );
xor ( n57187 , n57066 , n57070 );
xor ( n57188 , n57187 , n57073 );
and ( n57189 , n57185 , n57188 );
and ( n57190 , n57181 , n57188 );
or ( n57191 , n57186 , n57189 , n57190 );
and ( n57192 , n52954 , n53972 );
and ( n57193 , n52829 , n53970 );
nor ( n57194 , n57192 , n57193 );
xnor ( n57195 , n57194 , n53662 );
and ( n57196 , n57191 , n57195 );
xor ( n57197 , n56957 , n56961 );
xor ( n57198 , n57197 , n56964 );
and ( n57199 , n57195 , n57198 );
and ( n57200 , n57191 , n57198 );
or ( n57201 , n57196 , n57199 , n57200 );
xor ( n57202 , n57088 , n57092 );
xor ( n57203 , n57202 , n57095 );
and ( n57204 , n57201 , n57203 );
xor ( n57205 , n56967 , n56971 );
xor ( n57206 , n57205 , n56974 );
and ( n57207 , n57203 , n57206 );
and ( n57208 , n57201 , n57206 );
or ( n57209 , n57204 , n57207 , n57208 );
xor ( n57210 , n57098 , n57102 );
xor ( n57211 , n57210 , n57105 );
and ( n57212 , n57209 , n57211 );
xor ( n57213 , n57001 , n57005 );
xor ( n57214 , n57213 , n57008 );
and ( n57215 , n57211 , n57214 );
and ( n57216 , n57209 , n57214 );
or ( n57217 , n57212 , n57215 , n57216 );
and ( n57218 , n57177 , n57217 );
xor ( n57219 , n56997 , n57011 );
xor ( n57220 , n57219 , n57014 );
and ( n57221 , n57217 , n57220 );
and ( n57222 , n57177 , n57220 );
or ( n57223 , n57218 , n57221 , n57222 );
xor ( n57224 , n56754 , n56756 );
xor ( n57225 , n57224 , n56759 );
and ( n57226 , n57223 , n57225 );
xor ( n57227 , n57017 , n57116 );
xor ( n57228 , n57227 , n57119 );
and ( n57229 , n57225 , n57228 );
and ( n57230 , n57223 , n57228 );
or ( n57231 , n57226 , n57229 , n57230 );
and ( n57232 , n57133 , n57231 );
xor ( n57233 , n57223 , n57225 );
xor ( n57234 , n57233 , n57228 );
and ( n57235 , n56495 , n52121 );
and ( n57236 , n56336 , n52119 );
nor ( n57237 , n57235 , n57236 );
xnor ( n57238 , n57237 , n52087 );
and ( n57239 , n56855 , n52092 );
and ( n57240 , n56806 , n52090 );
nor ( n57241 , n57239 , n57240 );
xnor ( n57242 , n57241 , n52072 );
and ( n57243 , n57238 , n57242 );
buf ( n57244 , n51722 );
and ( n57245 , n57244 , n52059 );
and ( n57246 , n57027 , n52057 );
nor ( n57247 , n57245 , n57246 );
not ( n57248 , n57247 );
and ( n57249 , n57242 , n57248 );
and ( n57250 , n57238 , n57248 );
or ( n57251 , n57243 , n57249 , n57250 );
and ( n57252 , n55769 , n52318 );
and ( n57253 , n55720 , n52316 );
nor ( n57254 , n57252 , n57253 );
xnor ( n57255 , n57254 , n52213 );
and ( n57256 , n57251 , n57255 );
and ( n57257 , n56071 , n52170 );
and ( n57258 , n56073 , n52168 );
nor ( n57259 , n57257 , n57258 );
xnor ( n57260 , n57259 , n52152 );
and ( n57261 , n57255 , n57260 );
and ( n57262 , n57251 , n57260 );
or ( n57263 , n57256 , n57261 , n57262 );
and ( n57264 , n55406 , n52346 );
and ( n57265 , n55365 , n52344 );
nor ( n57266 , n57264 , n57265 );
xnor ( n57267 , n57266 , n52300 );
and ( n57268 , n57263 , n57267 );
and ( n57269 , n55720 , n52318 );
and ( n57270 , n55661 , n52316 );
nor ( n57271 , n57269 , n57270 );
xnor ( n57272 , n57271 , n52213 );
and ( n57273 , n57267 , n57272 );
and ( n57274 , n57263 , n57272 );
or ( n57275 , n57268 , n57273 , n57274 );
and ( n57276 , n54767 , n52617 );
and ( n57277 , n54715 , n52615 );
nor ( n57278 , n57276 , n57277 );
xnor ( n57279 , n57278 , n52558 );
and ( n57280 , n57275 , n57279 );
xor ( n57281 , n56862 , n56866 );
xor ( n57282 , n57281 , n56869 );
and ( n57283 , n57279 , n57282 );
and ( n57284 , n57275 , n57282 );
or ( n57285 , n57280 , n57283 , n57284 );
and ( n57286 , n54715 , n52617 );
and ( n57287 , n54466 , n52615 );
nor ( n57288 , n57286 , n57287 );
xnor ( n57289 , n57288 , n52558 );
and ( n57290 , n57285 , n57289 );
xor ( n57291 , n56872 , n56876 );
xor ( n57292 , n57291 , n56879 );
and ( n57293 , n57289 , n57292 );
and ( n57294 , n57285 , n57292 );
or ( n57295 , n57290 , n57293 , n57294 );
and ( n57296 , n55365 , n52540 );
and ( n57297 , n55199 , n52538 );
nor ( n57298 , n57296 , n57297 );
xnor ( n57299 , n57298 , n52424 );
and ( n57300 , n55661 , n52346 );
and ( n57301 , n55406 , n52344 );
nor ( n57302 , n57300 , n57301 );
xnor ( n57303 , n57302 , n52300 );
and ( n57304 , n57299 , n57303 );
xor ( n57305 , n57021 , n57025 );
xor ( n57306 , n57305 , n57031 );
and ( n57307 , n57303 , n57306 );
and ( n57308 , n57299 , n57306 );
or ( n57309 , n57304 , n57307 , n57308 );
and ( n57310 , n55199 , n52540 );
and ( n57311 , n55055 , n52538 );
nor ( n57312 , n57310 , n57311 );
xnor ( n57313 , n57312 , n52424 );
and ( n57314 , n57309 , n57313 );
xor ( n57315 , n57034 , n57038 );
xor ( n57316 , n57315 , n57041 );
and ( n57317 , n57313 , n57316 );
and ( n57318 , n57309 , n57316 );
or ( n57319 , n57314 , n57317 , n57318 );
and ( n57320 , n55055 , n52540 );
and ( n57321 , n54885 , n52538 );
nor ( n57322 , n57320 , n57321 );
xnor ( n57323 , n57322 , n52424 );
and ( n57324 , n57319 , n57323 );
xor ( n57325 , n57044 , n57048 );
xor ( n57326 , n57325 , n57053 );
and ( n57327 , n57323 , n57326 );
and ( n57328 , n57319 , n57326 );
or ( n57329 , n57324 , n57327 , n57328 );
and ( n57330 , n54364 , n52886 );
and ( n57331 , n54078 , n52884 );
nor ( n57332 , n57330 , n57331 );
xnor ( n57333 , n57332 , n52657 );
and ( n57334 , n57329 , n57333 );
xor ( n57335 , n57056 , n57060 );
xor ( n57336 , n57335 , n57063 );
and ( n57337 , n57333 , n57336 );
and ( n57338 , n57329 , n57336 );
or ( n57339 , n57334 , n57337 , n57338 );
and ( n57340 , n57295 , n57339 );
and ( n57341 , n53783 , n53021 );
and ( n57342 , n53785 , n53019 );
nor ( n57343 , n57341 , n57342 );
xnor ( n57344 , n57343 , n52839 );
and ( n57345 , n57339 , n57344 );
and ( n57346 , n57295 , n57344 );
or ( n57347 , n57340 , n57345 , n57346 );
xor ( n57348 , n57076 , n57080 );
xor ( n57349 , n57348 , n57085 );
and ( n57350 , n57347 , n57349 );
xor ( n57351 , n57147 , n57151 );
xor ( n57352 , n57351 , n57154 );
and ( n57353 , n57349 , n57352 );
and ( n57354 , n57347 , n57352 );
or ( n57355 , n57350 , n57353 , n57354 );
and ( n57356 , n52439 , n55033 );
and ( n57357 , n52431 , n55030 );
nor ( n57358 , n57356 , n57357 );
xnor ( n57359 , n57358 , n53885 );
and ( n57360 , n57355 , n57359 );
and ( n57361 , n52639 , n54693 );
and ( n57362 , n52565 , n54691 );
nor ( n57363 , n57361 , n57362 );
xnor ( n57364 , n57363 , n53892 );
and ( n57365 , n57359 , n57364 );
and ( n57366 , n57355 , n57364 );
or ( n57367 , n57360 , n57365 , n57366 );
and ( n57368 , n52565 , n55033 );
and ( n57369 , n52439 , n55030 );
nor ( n57370 , n57368 , n57369 );
xnor ( n57371 , n57370 , n53885 );
and ( n57372 , n52664 , n54693 );
and ( n57373 , n52639 , n54691 );
nor ( n57374 , n57372 , n57373 );
xnor ( n57375 , n57374 , n53892 );
and ( n57376 , n57371 , n57375 );
and ( n57377 , n52809 , n54285 );
and ( n57378 , n52718 , n54283 );
nor ( n57379 , n57377 , n57378 );
xnor ( n57380 , n57379 , n53794 );
and ( n57381 , n57375 , n57380 );
and ( n57382 , n57371 , n57380 );
or ( n57383 , n57376 , n57381 , n57382 );
and ( n57384 , n53322 , n53739 );
and ( n57385 , n53148 , n53737 );
nor ( n57386 , n57384 , n57385 );
xnor ( n57387 , n57386 , n53315 );
and ( n57388 , n53644 , n53455 );
and ( n57389 , n53499 , n53453 );
nor ( n57390 , n57388 , n57389 );
xnor ( n57391 , n57390 , n53159 );
and ( n57392 , n57387 , n57391 );
xor ( n57393 , n57285 , n57289 );
xor ( n57394 , n57393 , n57292 );
and ( n57395 , n57391 , n57394 );
and ( n57396 , n57387 , n57394 );
or ( n57397 , n57392 , n57395 , n57396 );
and ( n57398 , n52829 , n54285 );
and ( n57399 , n52809 , n54283 );
nor ( n57400 , n57398 , n57399 );
xnor ( n57401 , n57400 , n53794 );
and ( n57402 , n57397 , n57401 );
xor ( n57403 , n57295 , n57339 );
xor ( n57404 , n57403 , n57344 );
and ( n57405 , n57401 , n57404 );
and ( n57406 , n57397 , n57404 );
or ( n57407 , n57402 , n57405 , n57406 );
and ( n57408 , n54078 , n53021 );
and ( n57409 , n53895 , n53019 );
nor ( n57410 , n57408 , n57409 );
xnor ( n57411 , n57410 , n52839 );
and ( n57412 , n54466 , n52886 );
and ( n57413 , n54364 , n52884 );
nor ( n57414 , n57412 , n57413 );
xnor ( n57415 , n57414 , n52657 );
and ( n57416 , n57411 , n57415 );
xor ( n57417 , n57275 , n57279 );
xor ( n57418 , n57417 , n57282 );
and ( n57419 , n57415 , n57418 );
and ( n57420 , n57411 , n57418 );
or ( n57421 , n57416 , n57419 , n57420 );
and ( n57422 , n53785 , n53293 );
and ( n57423 , n53652 , n53291 );
nor ( n57424 , n57422 , n57423 );
xnor ( n57425 , n57424 , n52963 );
and ( n57426 , n57421 , n57425 );
and ( n57427 , n53895 , n53021 );
and ( n57428 , n53783 , n53019 );
nor ( n57429 , n57427 , n57428 );
xnor ( n57430 , n57429 , n52839 );
and ( n57431 , n57425 , n57430 );
and ( n57432 , n57421 , n57430 );
or ( n57433 , n57426 , n57431 , n57432 );
and ( n57434 , n52952 , n53972 );
and ( n57435 , n52954 , n53970 );
nor ( n57436 , n57434 , n57435 );
xnor ( n57437 , n57436 , n53662 );
and ( n57438 , n57433 , n57437 );
xor ( n57439 , n57137 , n57141 );
xor ( n57440 , n57439 , n57144 );
and ( n57441 , n57437 , n57440 );
and ( n57442 , n57433 , n57440 );
or ( n57443 , n57438 , n57441 , n57442 );
and ( n57444 , n57407 , n57443 );
xor ( n57445 , n57191 , n57195 );
xor ( n57446 , n57445 , n57198 );
and ( n57447 , n57443 , n57446 );
and ( n57448 , n57407 , n57446 );
or ( n57449 , n57444 , n57447 , n57448 );
and ( n57450 , n57383 , n57449 );
xor ( n57451 , n57157 , n57161 );
xor ( n57452 , n57451 , n57164 );
and ( n57453 , n57449 , n57452 );
and ( n57454 , n57383 , n57452 );
or ( n57455 , n57450 , n57453 , n57454 );
and ( n57456 , n57367 , n57455 );
xor ( n57457 , n57167 , n57171 );
xor ( n57458 , n57457 , n57174 );
and ( n57459 , n57455 , n57458 );
and ( n57460 , n57367 , n57458 );
or ( n57461 , n57456 , n57459 , n57460 );
xor ( n57462 , n57108 , n57110 );
xor ( n57463 , n57462 , n57113 );
and ( n57464 , n57461 , n57463 );
xor ( n57465 , n57177 , n57217 );
xor ( n57466 , n57465 , n57220 );
and ( n57467 , n57463 , n57466 );
and ( n57468 , n57461 , n57466 );
or ( n57469 , n57464 , n57467 , n57468 );
and ( n57470 , n57234 , n57469 );
xor ( n57471 , n57461 , n57463 );
xor ( n57472 , n57471 , n57466 );
and ( n57473 , n53148 , n53972 );
and ( n57474 , n53150 , n53970 );
nor ( n57475 , n57473 , n57474 );
xnor ( n57476 , n57475 , n53662 );
and ( n57477 , n53499 , n53739 );
and ( n57478 , n53322 , n53737 );
nor ( n57479 , n57477 , n57478 );
xnor ( n57480 , n57479 , n53315 );
and ( n57481 , n57476 , n57480 );
xor ( n57482 , n57411 , n57415 );
xor ( n57483 , n57482 , n57418 );
and ( n57484 , n57480 , n57483 );
and ( n57485 , n57476 , n57483 );
or ( n57486 , n57481 , n57484 , n57485 );
and ( n57487 , n52954 , n54285 );
and ( n57488 , n52829 , n54283 );
nor ( n57489 , n57487 , n57488 );
xnor ( n57490 , n57489 , n53794 );
and ( n57491 , n57486 , n57490 );
xor ( n57492 , n57421 , n57425 );
xor ( n57493 , n57492 , n57430 );
and ( n57494 , n57490 , n57493 );
and ( n57495 , n57486 , n57493 );
or ( n57496 , n57491 , n57494 , n57495 );
and ( n57497 , n52718 , n54693 );
and ( n57498 , n52664 , n54691 );
nor ( n57499 , n57497 , n57498 );
xnor ( n57500 , n57499 , n53892 );
and ( n57501 , n57496 , n57500 );
xor ( n57502 , n57433 , n57437 );
xor ( n57503 , n57502 , n57440 );
and ( n57504 , n57500 , n57503 );
and ( n57505 , n57496 , n57503 );
or ( n57506 , n57501 , n57504 , n57505 );
and ( n57507 , n57027 , n52121 );
and ( n57508 , n56855 , n52119 );
nor ( n57509 , n57507 , n57508 );
xnor ( n57510 , n57509 , n52087 );
buf ( n57511 , n51723 );
and ( n57512 , n57511 , n52092 );
and ( n57513 , n57244 , n52090 );
nor ( n57514 , n57512 , n57513 );
xnor ( n57515 , n57514 , n52072 );
and ( n57516 , n57510 , n57515 );
buf ( n57517 , n51725 );
and ( n57518 , n57517 , n52059 );
buf ( n57519 , n51724 );
and ( n57520 , n57519 , n52057 );
nor ( n57521 , n57518 , n57520 );
not ( n57522 , n57521 );
and ( n57523 , n57515 , n57522 );
and ( n57524 , n57510 , n57522 );
or ( n57525 , n57516 , n57523 , n57524 );
and ( n57526 , n57244 , n52092 );
and ( n57527 , n57027 , n52090 );
nor ( n57528 , n57526 , n57527 );
xnor ( n57529 , n57528 , n52072 );
and ( n57530 , n57525 , n57529 );
and ( n57531 , n57519 , n52059 );
and ( n57532 , n57511 , n52057 );
nor ( n57533 , n57531 , n57532 );
not ( n57534 , n57533 );
and ( n57535 , n57529 , n57534 );
and ( n57536 , n57525 , n57534 );
or ( n57537 , n57530 , n57535 , n57536 );
and ( n57538 , n57027 , n52092 );
and ( n57539 , n56855 , n52090 );
nor ( n57540 , n57538 , n57539 );
xnor ( n57541 , n57540 , n52072 );
and ( n57542 , n57537 , n57541 );
and ( n57543 , n57511 , n52059 );
and ( n57544 , n57244 , n52057 );
nor ( n57545 , n57543 , n57544 );
not ( n57546 , n57545 );
and ( n57547 , n57541 , n57546 );
and ( n57548 , n57537 , n57546 );
or ( n57549 , n57542 , n57547 , n57548 );
and ( n57550 , n56073 , n52318 );
and ( n57551 , n55769 , n52316 );
nor ( n57552 , n57550 , n57551 );
xnor ( n57553 , n57552 , n52213 );
and ( n57554 , n57549 , n57553 );
and ( n57555 , n56338 , n52170 );
and ( n57556 , n56071 , n52168 );
nor ( n57557 , n57555 , n57556 );
xnor ( n57558 , n57557 , n52152 );
and ( n57559 , n57553 , n57558 );
and ( n57560 , n57549 , n57558 );
or ( n57561 , n57554 , n57559 , n57560 );
and ( n57562 , n56071 , n52318 );
and ( n57563 , n56073 , n52316 );
nor ( n57564 , n57562 , n57563 );
xnor ( n57565 , n57564 , n52213 );
and ( n57566 , n56336 , n52170 );
and ( n57567 , n56338 , n52168 );
nor ( n57568 , n57566 , n57567 );
xnor ( n57569 , n57568 , n52152 );
and ( n57570 , n57565 , n57569 );
and ( n57571 , n56806 , n52121 );
and ( n57572 , n56495 , n52119 );
nor ( n57573 , n57571 , n57572 );
xnor ( n57574 , n57573 , n52087 );
and ( n57575 , n57569 , n57574 );
and ( n57576 , n57565 , n57574 );
or ( n57577 , n57570 , n57575 , n57576 );
and ( n57578 , n56495 , n52170 );
and ( n57579 , n56336 , n52168 );
nor ( n57580 , n57578 , n57579 );
xnor ( n57581 , n57580 , n52152 );
and ( n57582 , n56855 , n52121 );
and ( n57583 , n56806 , n52119 );
nor ( n57584 , n57582 , n57583 );
xnor ( n57585 , n57584 , n52087 );
and ( n57586 , n57581 , n57585 );
xor ( n57587 , n57525 , n57529 );
xor ( n57588 , n57587 , n57534 );
and ( n57589 , n57585 , n57588 );
and ( n57590 , n57581 , n57588 );
or ( n57591 , n57586 , n57589 , n57590 );
and ( n57592 , n55769 , n52346 );
and ( n57593 , n55720 , n52344 );
nor ( n57594 , n57592 , n57593 );
xnor ( n57595 , n57594 , n52300 );
and ( n57596 , n57591 , n57595 );
xor ( n57597 , n57537 , n57541 );
xor ( n57598 , n57597 , n57546 );
and ( n57599 , n57595 , n57598 );
and ( n57600 , n57591 , n57598 );
or ( n57601 , n57596 , n57599 , n57600 );
and ( n57602 , n57577 , n57601 );
xor ( n57603 , n57238 , n57242 );
xor ( n57604 , n57603 , n57248 );
and ( n57605 , n57601 , n57604 );
and ( n57606 , n57577 , n57604 );
or ( n57607 , n57602 , n57605 , n57606 );
and ( n57608 , n57561 , n57607 );
xor ( n57609 , n57251 , n57255 );
xor ( n57610 , n57609 , n57260 );
and ( n57611 , n57607 , n57610 );
and ( n57612 , n57561 , n57610 );
or ( n57613 , n57608 , n57611 , n57612 );
and ( n57614 , n54885 , n52617 );
and ( n57615 , n54767 , n52615 );
nor ( n57616 , n57614 , n57615 );
xnor ( n57617 , n57616 , n52558 );
and ( n57618 , n57613 , n57617 );
xor ( n57619 , n57263 , n57267 );
xor ( n57620 , n57619 , n57272 );
and ( n57621 , n57617 , n57620 );
and ( n57622 , n57613 , n57620 );
or ( n57623 , n57618 , n57621 , n57622 );
and ( n57624 , n53652 , n53455 );
and ( n57625 , n53644 , n53453 );
nor ( n57626 , n57624 , n57625 );
xnor ( n57627 , n57626 , n53159 );
and ( n57628 , n57623 , n57627 );
xor ( n57629 , n57319 , n57323 );
xor ( n57630 , n57629 , n57326 );
and ( n57631 , n57627 , n57630 );
and ( n57632 , n57623 , n57630 );
or ( n57633 , n57628 , n57631 , n57632 );
and ( n57634 , n53150 , n53972 );
and ( n57635 , n52952 , n53970 );
nor ( n57636 , n57634 , n57635 );
xnor ( n57637 , n57636 , n53662 );
and ( n57638 , n57633 , n57637 );
xor ( n57639 , n57329 , n57333 );
xor ( n57640 , n57639 , n57336 );
and ( n57641 , n57637 , n57640 );
and ( n57642 , n57633 , n57640 );
or ( n57643 , n57638 , n57641 , n57642 );
and ( n57644 , n52639 , n55033 );
and ( n57645 , n52565 , n55030 );
nor ( n57646 , n57644 , n57645 );
xnor ( n57647 , n57646 , n53885 );
and ( n57648 , n57643 , n57647 );
xor ( n57649 , n57181 , n57185 );
xor ( n57650 , n57649 , n57188 );
and ( n57651 , n57647 , n57650 );
and ( n57652 , n57643 , n57650 );
or ( n57653 , n57648 , n57651 , n57652 );
and ( n57654 , n57506 , n57653 );
xor ( n57655 , n57347 , n57349 );
xor ( n57656 , n57655 , n57352 );
and ( n57657 , n57653 , n57656 );
and ( n57658 , n57506 , n57656 );
or ( n57659 , n57654 , n57657 , n57658 );
xor ( n57660 , n57355 , n57359 );
xor ( n57661 , n57660 , n57364 );
and ( n57662 , n57659 , n57661 );
xor ( n57663 , n57201 , n57203 );
xor ( n57664 , n57663 , n57206 );
and ( n57665 , n57661 , n57664 );
and ( n57666 , n57659 , n57664 );
or ( n57667 , n57662 , n57665 , n57666 );
xor ( n57668 , n57209 , n57211 );
xor ( n57669 , n57668 , n57214 );
and ( n57670 , n57667 , n57669 );
xor ( n57671 , n57367 , n57455 );
xor ( n57672 , n57671 , n57458 );
and ( n57673 , n57669 , n57672 );
and ( n57674 , n57667 , n57672 );
or ( n57675 , n57670 , n57673 , n57674 );
and ( n57676 , n57472 , n57675 );
xor ( n57677 , n57667 , n57669 );
xor ( n57678 , n57677 , n57672 );
and ( n57679 , n57244 , n52121 );
and ( n57680 , n57027 , n52119 );
nor ( n57681 , n57679 , n57680 );
xnor ( n57682 , n57681 , n52087 );
and ( n57683 , n57519 , n52092 );
and ( n57684 , n57511 , n52090 );
nor ( n57685 , n57683 , n57684 );
xnor ( n57686 , n57685 , n52072 );
and ( n57687 , n57682 , n57686 );
buf ( n57688 , n51726 );
and ( n57689 , n57688 , n52059 );
and ( n57690 , n57517 , n52057 );
nor ( n57691 , n57689 , n57690 );
not ( n57692 , n57691 );
and ( n57693 , n57686 , n57692 );
and ( n57694 , n57682 , n57692 );
or ( n57695 , n57687 , n57693 , n57694 );
and ( n57696 , n56336 , n52318 );
and ( n57697 , n56338 , n52316 );
nor ( n57698 , n57696 , n57697 );
xnor ( n57699 , n57698 , n52213 );
and ( n57700 , n57695 , n57699 );
xor ( n57701 , n57510 , n57515 );
xor ( n57702 , n57701 , n57522 );
and ( n57703 , n57699 , n57702 );
and ( n57704 , n57695 , n57702 );
or ( n57705 , n57700 , n57703 , n57704 );
and ( n57706 , n56073 , n52346 );
and ( n57707 , n55769 , n52344 );
nor ( n57708 , n57706 , n57707 );
xnor ( n57709 , n57708 , n52300 );
and ( n57710 , n57705 , n57709 );
and ( n57711 , n56338 , n52318 );
and ( n57712 , n56071 , n52316 );
nor ( n57713 , n57711 , n57712 );
xnor ( n57714 , n57713 , n52213 );
and ( n57715 , n57709 , n57714 );
and ( n57716 , n57705 , n57714 );
or ( n57717 , n57710 , n57715 , n57716 );
and ( n57718 , n55365 , n52617 );
and ( n57719 , n55199 , n52615 );
nor ( n57720 , n57718 , n57719 );
xnor ( n57721 , n57720 , n52558 );
and ( n57722 , n57717 , n57721 );
xor ( n57723 , n57565 , n57569 );
xor ( n57724 , n57723 , n57574 );
and ( n57725 , n57721 , n57724 );
and ( n57726 , n57717 , n57724 );
or ( n57727 , n57722 , n57725 , n57726 );
and ( n57728 , n55199 , n52617 );
and ( n57729 , n55055 , n52615 );
nor ( n57730 , n57728 , n57729 );
xnor ( n57731 , n57730 , n52558 );
and ( n57732 , n57727 , n57731 );
xor ( n57733 , n57577 , n57601 );
xor ( n57734 , n57733 , n57604 );
and ( n57735 , n57731 , n57734 );
and ( n57736 , n57727 , n57734 );
or ( n57737 , n57732 , n57735 , n57736 );
and ( n57738 , n55055 , n52617 );
and ( n57739 , n54885 , n52615 );
nor ( n57740 , n57738 , n57739 );
xnor ( n57741 , n57740 , n52558 );
and ( n57742 , n57737 , n57741 );
xor ( n57743 , n57561 , n57607 );
xor ( n57744 , n57743 , n57610 );
and ( n57745 , n57741 , n57744 );
and ( n57746 , n57737 , n57744 );
or ( n57747 , n57742 , n57745 , n57746 );
and ( n57748 , n53895 , n53293 );
and ( n57749 , n53783 , n53291 );
nor ( n57750 , n57748 , n57749 );
xnor ( n57751 , n57750 , n52963 );
and ( n57752 , n57747 , n57751 );
and ( n57753 , n54364 , n53021 );
and ( n57754 , n54078 , n53019 );
nor ( n57755 , n57753 , n57754 );
xnor ( n57756 , n57755 , n52839 );
and ( n57757 , n57751 , n57756 );
and ( n57758 , n57747 , n57756 );
or ( n57759 , n57752 , n57757 , n57758 );
and ( n57760 , n55406 , n52540 );
and ( n57761 , n55365 , n52538 );
nor ( n57762 , n57760 , n57761 );
xnor ( n57763 , n57762 , n52424 );
and ( n57764 , n55720 , n52346 );
and ( n57765 , n55661 , n52344 );
nor ( n57766 , n57764 , n57765 );
xnor ( n57767 , n57766 , n52300 );
and ( n57768 , n57763 , n57767 );
xor ( n57769 , n57549 , n57553 );
xor ( n57770 , n57769 , n57558 );
and ( n57771 , n57767 , n57770 );
and ( n57772 , n57763 , n57770 );
or ( n57773 , n57768 , n57771 , n57772 );
and ( n57774 , n54767 , n52886 );
and ( n57775 , n54715 , n52884 );
nor ( n57776 , n57774 , n57775 );
xnor ( n57777 , n57776 , n52657 );
and ( n57778 , n57773 , n57777 );
xor ( n57779 , n57299 , n57303 );
xor ( n57780 , n57779 , n57306 );
and ( n57781 , n57777 , n57780 );
and ( n57782 , n57773 , n57780 );
or ( n57783 , n57778 , n57781 , n57782 );
and ( n57784 , n54715 , n52886 );
and ( n57785 , n54466 , n52884 );
nor ( n57786 , n57784 , n57785 );
xnor ( n57787 , n57786 , n52657 );
and ( n57788 , n57783 , n57787 );
xor ( n57789 , n57309 , n57313 );
xor ( n57790 , n57789 , n57316 );
and ( n57791 , n57787 , n57790 );
and ( n57792 , n57783 , n57790 );
or ( n57793 , n57788 , n57791 , n57792 );
and ( n57794 , n57759 , n57793 );
and ( n57795 , n53783 , n53293 );
and ( n57796 , n53785 , n53291 );
nor ( n57797 , n57795 , n57796 );
xnor ( n57798 , n57797 , n52963 );
and ( n57799 , n57793 , n57798 );
and ( n57800 , n57759 , n57798 );
or ( n57801 , n57794 , n57799 , n57800 );
and ( n57802 , n54078 , n53293 );
and ( n57803 , n53895 , n53291 );
nor ( n57804 , n57802 , n57803 );
xnor ( n57805 , n57804 , n52963 );
and ( n57806 , n54466 , n53021 );
and ( n57807 , n54364 , n53019 );
nor ( n57808 , n57806 , n57807 );
xnor ( n57809 , n57808 , n52839 );
and ( n57810 , n57805 , n57809 );
xor ( n57811 , n57773 , n57777 );
xor ( n57812 , n57811 , n57780 );
and ( n57813 , n57809 , n57812 );
and ( n57814 , n57805 , n57812 );
or ( n57815 , n57810 , n57813 , n57814 );
and ( n57816 , n53785 , n53455 );
and ( n57817 , n53652 , n53453 );
nor ( n57818 , n57816 , n57817 );
xnor ( n57819 , n57818 , n53159 );
and ( n57820 , n57815 , n57819 );
xor ( n57821 , n57613 , n57617 );
xor ( n57822 , n57821 , n57620 );
and ( n57823 , n57819 , n57822 );
and ( n57824 , n57815 , n57822 );
or ( n57825 , n57820 , n57823 , n57824 );
and ( n57826 , n52952 , n54285 );
and ( n57827 , n52954 , n54283 );
nor ( n57828 , n57826 , n57827 );
xnor ( n57829 , n57828 , n53794 );
and ( n57830 , n57825 , n57829 );
xor ( n57831 , n57623 , n57627 );
xor ( n57832 , n57831 , n57630 );
and ( n57833 , n57829 , n57832 );
and ( n57834 , n57825 , n57832 );
or ( n57835 , n57830 , n57833 , n57834 );
and ( n57836 , n57801 , n57835 );
xor ( n57837 , n57387 , n57391 );
xor ( n57838 , n57837 , n57394 );
and ( n57839 , n57835 , n57838 );
and ( n57840 , n57801 , n57838 );
or ( n57841 , n57836 , n57839 , n57840 );
and ( n57842 , n52809 , n54693 );
and ( n57843 , n52718 , n54691 );
nor ( n57844 , n57842 , n57843 );
xnor ( n57845 , n57844 , n53892 );
xor ( n57846 , n57486 , n57490 );
xor ( n57847 , n57846 , n57493 );
and ( n57848 , n57845 , n57847 );
xor ( n57849 , n57633 , n57637 );
xor ( n57850 , n57849 , n57640 );
and ( n57851 , n57847 , n57850 );
and ( n57852 , n57845 , n57850 );
or ( n57853 , n57848 , n57851 , n57852 );
and ( n57854 , n57841 , n57853 );
xor ( n57855 , n57397 , n57401 );
xor ( n57856 , n57855 , n57404 );
and ( n57857 , n57853 , n57856 );
and ( n57858 , n57841 , n57856 );
or ( n57859 , n57854 , n57857 , n57858 );
xor ( n57860 , n57371 , n57375 );
xor ( n57861 , n57860 , n57380 );
and ( n57862 , n57859 , n57861 );
xor ( n57863 , n57407 , n57443 );
xor ( n57864 , n57863 , n57446 );
and ( n57865 , n57861 , n57864 );
and ( n57866 , n57859 , n57864 );
or ( n57867 , n57862 , n57865 , n57866 );
xor ( n57868 , n57659 , n57661 );
xor ( n57869 , n57868 , n57664 );
and ( n57870 , n57867 , n57869 );
xor ( n57871 , n57383 , n57449 );
xor ( n57872 , n57871 , n57452 );
and ( n57873 , n57869 , n57872 );
and ( n57874 , n57867 , n57872 );
or ( n57875 , n57870 , n57873 , n57874 );
and ( n57876 , n57678 , n57875 );
xor ( n57877 , n57867 , n57869 );
xor ( n57878 , n57877 , n57872 );
and ( n57879 , n53322 , n53972 );
and ( n57880 , n53148 , n53970 );
nor ( n57881 , n57879 , n57880 );
xnor ( n57882 , n57881 , n53662 );
and ( n57883 , n53644 , n53739 );
and ( n57884 , n53499 , n53737 );
nor ( n57885 , n57883 , n57884 );
xnor ( n57886 , n57885 , n53315 );
and ( n57887 , n57882 , n57886 );
xor ( n57888 , n57783 , n57787 );
xor ( n57889 , n57888 , n57790 );
and ( n57890 , n57886 , n57889 );
and ( n57891 , n57882 , n57889 );
or ( n57892 , n57887 , n57890 , n57891 );
and ( n57893 , n52829 , n54693 );
and ( n57894 , n52809 , n54691 );
nor ( n57895 , n57893 , n57894 );
xnor ( n57896 , n57895 , n53892 );
and ( n57897 , n57892 , n57896 );
xor ( n57898 , n57759 , n57793 );
xor ( n57899 , n57898 , n57798 );
and ( n57900 , n57896 , n57899 );
and ( n57901 , n57892 , n57899 );
or ( n57902 , n57897 , n57900 , n57901 );
and ( n57903 , n52664 , n55033 );
and ( n57904 , n52639 , n55030 );
nor ( n57905 , n57903 , n57904 );
xnor ( n57906 , n57905 , n53885 );
and ( n57907 , n57902 , n57906 );
xor ( n57908 , n57801 , n57835 );
xor ( n57909 , n57908 , n57838 );
and ( n57910 , n57906 , n57909 );
and ( n57911 , n57902 , n57909 );
or ( n57912 , n57907 , n57910 , n57911 );
xor ( n57913 , n57496 , n57500 );
xor ( n57914 , n57913 , n57503 );
and ( n57915 , n57912 , n57914 );
xor ( n57916 , n57643 , n57647 );
xor ( n57917 , n57916 , n57650 );
and ( n57918 , n57914 , n57917 );
and ( n57919 , n57912 , n57917 );
or ( n57920 , n57915 , n57918 , n57919 );
xor ( n57921 , n57506 , n57653 );
xor ( n57922 , n57921 , n57656 );
and ( n57923 , n57920 , n57922 );
xor ( n57924 , n57859 , n57861 );
xor ( n57925 , n57924 , n57864 );
and ( n57926 , n57922 , n57925 );
and ( n57927 , n57920 , n57925 );
or ( n57928 , n57923 , n57926 , n57927 );
and ( n57929 , n57878 , n57928 );
xor ( n57930 , n57920 , n57922 );
xor ( n57931 , n57930 , n57925 );
and ( n57932 , n52718 , n55033 );
and ( n57933 , n52664 , n55030 );
nor ( n57934 , n57932 , n57933 );
xnor ( n57935 , n57934 , n53885 );
xor ( n57936 , n57892 , n57896 );
xor ( n57937 , n57936 , n57899 );
and ( n57938 , n57935 , n57937 );
xor ( n57939 , n57825 , n57829 );
xor ( n57940 , n57939 , n57832 );
and ( n57941 , n57937 , n57940 );
and ( n57942 , n57935 , n57940 );
or ( n57943 , n57938 , n57941 , n57942 );
and ( n57944 , n57511 , n52121 );
and ( n57945 , n57244 , n52119 );
nor ( n57946 , n57944 , n57945 );
xnor ( n57947 , n57946 , n52087 );
and ( n57948 , n57517 , n52092 );
and ( n57949 , n57519 , n52090 );
nor ( n57950 , n57948 , n57949 );
xnor ( n57951 , n57950 , n52072 );
and ( n57952 , n57947 , n57951 );
buf ( n57953 , n51727 );
and ( n57954 , n57953 , n52059 );
and ( n57955 , n57688 , n52057 );
nor ( n57956 , n57954 , n57955 );
not ( n57957 , n57956 );
and ( n57958 , n57951 , n57957 );
and ( n57959 , n57947 , n57957 );
or ( n57960 , n57952 , n57958 , n57959 );
and ( n57961 , n57519 , n52121 );
and ( n57962 , n57511 , n52119 );
nor ( n57963 , n57961 , n57962 );
xnor ( n57964 , n57963 , n52087 );
and ( n57965 , n57688 , n52092 );
and ( n57966 , n57517 , n52090 );
nor ( n57967 , n57965 , n57966 );
xnor ( n57968 , n57967 , n52072 );
and ( n57969 , n57964 , n57968 );
buf ( n57970 , n51728 );
and ( n57971 , n57970 , n52059 );
and ( n57972 , n57953 , n52057 );
nor ( n57973 , n57971 , n57972 );
not ( n57974 , n57973 );
and ( n57975 , n57968 , n57974 );
and ( n57976 , n57964 , n57974 );
or ( n57977 , n57969 , n57975 , n57976 );
and ( n57978 , n57027 , n52170 );
and ( n57979 , n56855 , n52168 );
nor ( n57980 , n57978 , n57979 );
xnor ( n57981 , n57980 , n52152 );
and ( n57982 , n57977 , n57981 );
xor ( n57983 , n57947 , n57951 );
xor ( n57984 , n57983 , n57957 );
and ( n57985 , n57981 , n57984 );
and ( n57986 , n57977 , n57984 );
or ( n57987 , n57982 , n57985 , n57986 );
and ( n57988 , n57960 , n57987 );
xor ( n57989 , n57682 , n57686 );
xor ( n57990 , n57989 , n57692 );
and ( n57991 , n57987 , n57990 );
and ( n57992 , n57960 , n57990 );
or ( n57993 , n57988 , n57991 , n57992 );
and ( n57994 , n56071 , n52346 );
and ( n57995 , n56073 , n52344 );
nor ( n57996 , n57994 , n57995 );
xnor ( n57997 , n57996 , n52300 );
and ( n57998 , n57993 , n57997 );
and ( n57999 , n56806 , n52170 );
and ( n58000 , n56495 , n52168 );
nor ( n58001 , n57999 , n58000 );
xnor ( n58002 , n58001 , n52152 );
and ( n58003 , n57997 , n58002 );
and ( n58004 , n57993 , n58002 );
or ( n58005 , n57998 , n58003 , n58004 );
and ( n58006 , n55406 , n52617 );
and ( n58007 , n55365 , n52615 );
nor ( n58008 , n58006 , n58007 );
xnor ( n58009 , n58008 , n52558 );
and ( n58010 , n58005 , n58009 );
xor ( n58011 , n57581 , n57585 );
xor ( n58012 , n58011 , n57588 );
and ( n58013 , n58009 , n58012 );
and ( n58014 , n58005 , n58012 );
or ( n58015 , n58010 , n58013 , n58014 );
and ( n58016 , n55661 , n52540 );
and ( n58017 , n55406 , n52538 );
nor ( n58018 , n58016 , n58017 );
xnor ( n58019 , n58018 , n52424 );
and ( n58020 , n58015 , n58019 );
xor ( n58021 , n57591 , n57595 );
xor ( n58022 , n58021 , n57598 );
and ( n58023 , n58019 , n58022 );
and ( n58024 , n58015 , n58022 );
or ( n58025 , n58020 , n58023 , n58024 );
and ( n58026 , n54885 , n52886 );
and ( n58027 , n54767 , n52884 );
nor ( n58028 , n58026 , n58027 );
xnor ( n58029 , n58028 , n52657 );
and ( n58030 , n58025 , n58029 );
xor ( n58031 , n57763 , n57767 );
xor ( n58032 , n58031 , n57770 );
and ( n58033 , n58029 , n58032 );
and ( n58034 , n58025 , n58032 );
or ( n58035 , n58030 , n58033 , n58034 );
and ( n58036 , n56495 , n52318 );
and ( n58037 , n56336 , n52316 );
nor ( n58038 , n58036 , n58037 );
xnor ( n58039 , n58038 , n52213 );
and ( n58040 , n56855 , n52170 );
and ( n58041 , n56806 , n52168 );
nor ( n58042 , n58040 , n58041 );
xnor ( n58043 , n58042 , n52152 );
and ( n58044 , n58039 , n58043 );
xor ( n58045 , n57960 , n57987 );
xor ( n58046 , n58045 , n57990 );
and ( n58047 , n58043 , n58046 );
and ( n58048 , n58039 , n58046 );
or ( n58049 , n58044 , n58047 , n58048 );
and ( n58050 , n55769 , n52540 );
and ( n58051 , n55720 , n52538 );
nor ( n58052 , n58050 , n58051 );
xnor ( n58053 , n58052 , n52424 );
and ( n58054 , n58049 , n58053 );
xor ( n58055 , n57695 , n57699 );
xor ( n58056 , n58055 , n57702 );
and ( n58057 , n58053 , n58056 );
and ( n58058 , n58049 , n58056 );
or ( n58059 , n58054 , n58057 , n58058 );
and ( n58060 , n55720 , n52540 );
and ( n58061 , n55661 , n52538 );
nor ( n58062 , n58060 , n58061 );
xnor ( n58063 , n58062 , n52424 );
and ( n58064 , n58059 , n58063 );
xor ( n58065 , n57705 , n57709 );
xor ( n58066 , n58065 , n57714 );
and ( n58067 , n58063 , n58066 );
and ( n58068 , n58059 , n58066 );
or ( n58069 , n58064 , n58067 , n58068 );
and ( n58070 , n55055 , n52886 );
and ( n58071 , n54885 , n52884 );
nor ( n58072 , n58070 , n58071 );
xnor ( n58073 , n58072 , n52657 );
and ( n58074 , n58069 , n58073 );
xor ( n58075 , n57717 , n57721 );
xor ( n58076 , n58075 , n57724 );
and ( n58077 , n58073 , n58076 );
and ( n58078 , n58069 , n58076 );
or ( n58079 , n58074 , n58077 , n58078 );
and ( n58080 , n54715 , n53021 );
and ( n58081 , n54466 , n53019 );
nor ( n58082 , n58080 , n58081 );
xnor ( n58083 , n58082 , n52839 );
and ( n58084 , n58079 , n58083 );
xor ( n58085 , n57727 , n57731 );
xor ( n58086 , n58085 , n57734 );
and ( n58087 , n58083 , n58086 );
and ( n58088 , n58079 , n58086 );
or ( n58089 , n58084 , n58087 , n58088 );
and ( n58090 , n58035 , n58089 );
and ( n58091 , n53652 , n53739 );
and ( n58092 , n53644 , n53737 );
nor ( n58093 , n58091 , n58092 );
xnor ( n58094 , n58093 , n53315 );
and ( n58095 , n58089 , n58094 );
and ( n58096 , n58035 , n58094 );
or ( n58097 , n58090 , n58095 , n58096 );
and ( n58098 , n53150 , n54285 );
and ( n58099 , n52952 , n54283 );
nor ( n58100 , n58098 , n58099 );
xnor ( n58101 , n58100 , n53794 );
and ( n58102 , n58097 , n58101 );
xor ( n58103 , n57747 , n57751 );
xor ( n58104 , n58103 , n57756 );
and ( n58105 , n58101 , n58104 );
and ( n58106 , n58097 , n58104 );
or ( n58107 , n58102 , n58105 , n58106 );
and ( n58108 , n57517 , n52121 );
and ( n58109 , n57519 , n52119 );
nor ( n58110 , n58108 , n58109 );
xnor ( n58111 , n58110 , n52087 );
and ( n58112 , n57953 , n52092 );
and ( n58113 , n57688 , n52090 );
nor ( n58114 , n58112 , n58113 );
xnor ( n58115 , n58114 , n52072 );
and ( n58116 , n58111 , n58115 );
buf ( n58117 , n51729 );
and ( n58118 , n58117 , n52059 );
and ( n58119 , n57970 , n52057 );
nor ( n58120 , n58118 , n58119 );
not ( n58121 , n58120 );
and ( n58122 , n58115 , n58121 );
and ( n58123 , n58111 , n58121 );
or ( n58124 , n58116 , n58122 , n58123 );
and ( n58125 , n57244 , n52170 );
and ( n58126 , n57027 , n52168 );
nor ( n58127 , n58125 , n58126 );
xnor ( n58128 , n58127 , n52152 );
and ( n58129 , n58124 , n58128 );
xor ( n58130 , n57964 , n57968 );
xor ( n58131 , n58130 , n57974 );
and ( n58132 , n58128 , n58131 );
and ( n58133 , n58124 , n58131 );
or ( n58134 , n58129 , n58132 , n58133 );
and ( n58135 , n57688 , n52121 );
and ( n58136 , n57517 , n52119 );
nor ( n58137 , n58135 , n58136 );
xnor ( n58138 , n58137 , n52087 );
and ( n58139 , n57970 , n52092 );
and ( n58140 , n57953 , n52090 );
nor ( n58141 , n58139 , n58140 );
xnor ( n58142 , n58141 , n52072 );
and ( n58143 , n58138 , n58142 );
buf ( n58144 , n51730 );
and ( n58145 , n58144 , n52059 );
and ( n58146 , n58117 , n52057 );
nor ( n58147 , n58145 , n58146 );
not ( n58148 , n58147 );
and ( n58149 , n58142 , n58148 );
and ( n58150 , n58138 , n58148 );
or ( n58151 , n58143 , n58149 , n58150 );
and ( n58152 , n57511 , n52170 );
and ( n58153 , n57244 , n52168 );
nor ( n58154 , n58152 , n58153 );
xnor ( n58155 , n58154 , n52152 );
and ( n58156 , n58151 , n58155 );
xor ( n58157 , n58111 , n58115 );
xor ( n58158 , n58157 , n58121 );
and ( n58159 , n58155 , n58158 );
and ( n58160 , n58151 , n58158 );
or ( n58161 , n58156 , n58159 , n58160 );
and ( n58162 , n57953 , n52121 );
and ( n58163 , n57688 , n52119 );
nor ( n58164 , n58162 , n58163 );
xnor ( n58165 , n58164 , n52087 );
and ( n58166 , n58117 , n52092 );
and ( n58167 , n57970 , n52090 );
nor ( n58168 , n58166 , n58167 );
xnor ( n58169 , n58168 , n52072 );
and ( n58170 , n58165 , n58169 );
buf ( n58171 , n51731 );
and ( n58172 , n58171 , n52059 );
and ( n58173 , n58144 , n52057 );
nor ( n58174 , n58172 , n58173 );
not ( n58175 , n58174 );
and ( n58176 , n58169 , n58175 );
and ( n58177 , n58165 , n58175 );
or ( n58178 , n58170 , n58176 , n58177 );
and ( n58179 , n57519 , n52170 );
and ( n58180 , n57511 , n52168 );
nor ( n58181 , n58179 , n58180 );
xnor ( n58182 , n58181 , n52152 );
and ( n58183 , n58178 , n58182 );
xor ( n58184 , n58138 , n58142 );
xor ( n58185 , n58184 , n58148 );
and ( n58186 , n58182 , n58185 );
and ( n58187 , n58178 , n58185 );
or ( n58188 , n58183 , n58186 , n58187 );
and ( n58189 , n57027 , n52318 );
and ( n58190 , n56855 , n52316 );
nor ( n58191 , n58189 , n58190 );
xnor ( n58192 , n58191 , n52213 );
and ( n58193 , n58188 , n58192 );
xor ( n58194 , n58151 , n58155 );
xor ( n58195 , n58194 , n58158 );
and ( n58196 , n58192 , n58195 );
and ( n58197 , n58188 , n58195 );
or ( n58198 , n58193 , n58196 , n58197 );
and ( n58199 , n58161 , n58198 );
xor ( n58200 , n58124 , n58128 );
xor ( n58201 , n58200 , n58131 );
and ( n58202 , n58198 , n58201 );
and ( n58203 , n58161 , n58201 );
or ( n58204 , n58199 , n58202 , n58203 );
and ( n58205 , n58134 , n58204 );
xor ( n58206 , n57977 , n57981 );
xor ( n58207 , n58206 , n57984 );
and ( n58208 , n58204 , n58207 );
and ( n58209 , n58134 , n58207 );
or ( n58210 , n58205 , n58208 , n58209 );
and ( n58211 , n56073 , n52540 );
and ( n58212 , n55769 , n52538 );
nor ( n58213 , n58211 , n58212 );
xnor ( n58214 , n58213 , n52424 );
and ( n58215 , n58210 , n58214 );
and ( n58216 , n56338 , n52346 );
and ( n58217 , n56071 , n52344 );
nor ( n58218 , n58216 , n58217 );
xnor ( n58219 , n58218 , n52300 );
and ( n58220 , n58214 , n58219 );
and ( n58221 , n58210 , n58219 );
or ( n58222 , n58215 , n58220 , n58221 );
and ( n58223 , n55365 , n52886 );
and ( n58224 , n55199 , n52884 );
nor ( n58225 , n58223 , n58224 );
xnor ( n58226 , n58225 , n52657 );
and ( n58227 , n58222 , n58226 );
xor ( n58228 , n57993 , n57997 );
xor ( n58229 , n58228 , n58002 );
and ( n58230 , n58226 , n58229 );
and ( n58231 , n58222 , n58229 );
or ( n58232 , n58227 , n58230 , n58231 );
and ( n58233 , n55199 , n52886 );
and ( n58234 , n55055 , n52884 );
nor ( n58235 , n58233 , n58234 );
xnor ( n58236 , n58235 , n52657 );
and ( n58237 , n58232 , n58236 );
xor ( n58238 , n58005 , n58009 );
xor ( n58239 , n58238 , n58012 );
and ( n58240 , n58236 , n58239 );
and ( n58241 , n58232 , n58239 );
or ( n58242 , n58237 , n58240 , n58241 );
and ( n58243 , n54767 , n53021 );
and ( n58244 , n54715 , n53019 );
nor ( n58245 , n58243 , n58244 );
xnor ( n58246 , n58245 , n52839 );
and ( n58247 , n58242 , n58246 );
xor ( n58248 , n58015 , n58019 );
xor ( n58249 , n58248 , n58022 );
and ( n58250 , n58246 , n58249 );
and ( n58251 , n58242 , n58249 );
or ( n58252 , n58247 , n58250 , n58251 );
and ( n58253 , n53895 , n53455 );
and ( n58254 , n53783 , n53453 );
nor ( n58255 , n58253 , n58254 );
xnor ( n58256 , n58255 , n53159 );
and ( n58257 , n58252 , n58256 );
and ( n58258 , n54364 , n53293 );
and ( n58259 , n54078 , n53291 );
nor ( n58260 , n58258 , n58259 );
xnor ( n58261 , n58260 , n52963 );
and ( n58262 , n58256 , n58261 );
and ( n58263 , n58252 , n58261 );
or ( n58264 , n58257 , n58262 , n58263 );
and ( n58265 , n53148 , n54285 );
and ( n58266 , n53150 , n54283 );
nor ( n58267 , n58265 , n58266 );
xnor ( n58268 , n58267 , n53794 );
and ( n58269 , n58264 , n58268 );
and ( n58270 , n53499 , n53972 );
and ( n58271 , n53322 , n53970 );
nor ( n58272 , n58270 , n58271 );
xnor ( n58273 , n58272 , n53662 );
and ( n58274 , n58268 , n58273 );
and ( n58275 , n58264 , n58273 );
or ( n58276 , n58269 , n58274 , n58275 );
and ( n58277 , n52954 , n54693 );
and ( n58278 , n52829 , n54691 );
nor ( n58279 , n58277 , n58278 );
xnor ( n58280 , n58279 , n53892 );
and ( n58281 , n58276 , n58280 );
xor ( n58282 , n57815 , n57819 );
xor ( n58283 , n58282 , n57822 );
and ( n58284 , n58280 , n58283 );
and ( n58285 , n58276 , n58283 );
or ( n58286 , n58281 , n58284 , n58285 );
and ( n58287 , n58107 , n58286 );
xor ( n58288 , n57476 , n57480 );
xor ( n58289 , n58288 , n57483 );
and ( n58290 , n58286 , n58289 );
and ( n58291 , n58107 , n58289 );
or ( n58292 , n58287 , n58290 , n58291 );
and ( n58293 , n57943 , n58292 );
xor ( n58294 , n57845 , n57847 );
xor ( n58295 , n58294 , n57850 );
and ( n58296 , n58292 , n58295 );
and ( n58297 , n57943 , n58295 );
or ( n58298 , n58293 , n58296 , n58297 );
xor ( n58299 , n57841 , n57853 );
xor ( n58300 , n58299 , n57856 );
and ( n58301 , n58298 , n58300 );
xor ( n58302 , n57912 , n57914 );
xor ( n58303 , n58302 , n57917 );
and ( n58304 , n58300 , n58303 );
and ( n58305 , n58298 , n58303 );
or ( n58306 , n58301 , n58304 , n58305 );
and ( n58307 , n57931 , n58306 );
xor ( n58308 , n58298 , n58300 );
xor ( n58309 , n58308 , n58303 );
and ( n58310 , n54078 , n53455 );
and ( n58311 , n53895 , n53453 );
nor ( n58312 , n58310 , n58311 );
xnor ( n58313 , n58312 , n53159 );
and ( n58314 , n54466 , n53293 );
and ( n58315 , n54364 , n53291 );
nor ( n58316 , n58314 , n58315 );
xnor ( n58317 , n58316 , n52963 );
and ( n58318 , n58313 , n58317 );
xor ( n58319 , n58069 , n58073 );
xor ( n58320 , n58319 , n58076 );
and ( n58321 , n58317 , n58320 );
and ( n58322 , n58313 , n58320 );
or ( n58323 , n58318 , n58321 , n58322 );
and ( n58324 , n53322 , n54285 );
and ( n58325 , n53148 , n54283 );
nor ( n58326 , n58324 , n58325 );
xnor ( n58327 , n58326 , n53794 );
and ( n58328 , n58323 , n58327 );
and ( n58329 , n53644 , n53972 );
and ( n58330 , n53499 , n53970 );
nor ( n58331 , n58329 , n58330 );
xnor ( n58332 , n58331 , n53662 );
and ( n58333 , n58327 , n58332 );
and ( n58334 , n58323 , n58332 );
or ( n58335 , n58328 , n58333 , n58334 );
and ( n58336 , n52952 , n54693 );
and ( n58337 , n52954 , n54691 );
nor ( n58338 , n58336 , n58337 );
xnor ( n58339 , n58338 , n53892 );
and ( n58340 , n58335 , n58339 );
and ( n58341 , n53783 , n53455 );
and ( n58342 , n53785 , n53453 );
nor ( n58343 , n58341 , n58342 );
xnor ( n58344 , n58343 , n53159 );
xor ( n58345 , n57737 , n57741 );
xor ( n58346 , n58345 , n57744 );
xor ( n58347 , n58344 , n58346 );
xor ( n58348 , n57805 , n57809 );
xor ( n58349 , n58348 , n57812 );
xor ( n58350 , n58347 , n58349 );
and ( n58351 , n58339 , n58350 );
and ( n58352 , n58335 , n58350 );
or ( n58353 , n58340 , n58351 , n58352 );
and ( n58354 , n52809 , n55033 );
and ( n58355 , n52718 , n55030 );
nor ( n58356 , n58354 , n58355 );
xnor ( n58357 , n58356 , n53885 );
and ( n58358 , n58353 , n58357 );
xor ( n58359 , n58097 , n58101 );
xor ( n58360 , n58359 , n58104 );
and ( n58361 , n58357 , n58360 );
and ( n58362 , n58353 , n58360 );
or ( n58363 , n58358 , n58361 , n58362 );
and ( n58364 , n53785 , n53739 );
and ( n58365 , n53652 , n53737 );
nor ( n58366 , n58364 , n58365 );
xnor ( n58367 , n58366 , n53315 );
xor ( n58368 , n58025 , n58029 );
xor ( n58369 , n58368 , n58032 );
and ( n58370 , n58367 , n58369 );
xor ( n58371 , n58079 , n58083 );
xor ( n58372 , n58371 , n58086 );
and ( n58373 , n58369 , n58372 );
and ( n58374 , n58367 , n58372 );
or ( n58375 , n58370 , n58373 , n58374 );
and ( n58376 , n52829 , n55033 );
and ( n58377 , n52809 , n55030 );
nor ( n58378 , n58376 , n58377 );
xnor ( n58379 , n58378 , n53885 );
and ( n58380 , n58375 , n58379 );
xor ( n58381 , n58035 , n58089 );
xor ( n58382 , n58381 , n58094 );
and ( n58383 , n58379 , n58382 );
and ( n58384 , n58375 , n58382 );
or ( n58385 , n58380 , n58383 , n58384 );
and ( n58386 , n58344 , n58346 );
and ( n58387 , n58346 , n58349 );
and ( n58388 , n58344 , n58349 );
or ( n58389 , n58386 , n58387 , n58388 );
and ( n58390 , n58385 , n58389 );
xor ( n58391 , n57882 , n57886 );
xor ( n58392 , n58391 , n57889 );
and ( n58393 , n58389 , n58392 );
and ( n58394 , n58385 , n58392 );
or ( n58395 , n58390 , n58393 , n58394 );
and ( n58396 , n58363 , n58395 );
xor ( n58397 , n58107 , n58286 );
xor ( n58398 , n58397 , n58289 );
and ( n58399 , n58395 , n58398 );
and ( n58400 , n58363 , n58398 );
or ( n58401 , n58396 , n58399 , n58400 );
xor ( n58402 , n57902 , n57906 );
xor ( n58403 , n58402 , n57909 );
and ( n58404 , n58401 , n58403 );
xor ( n58405 , n57943 , n58292 );
xor ( n58406 , n58405 , n58295 );
and ( n58407 , n58403 , n58406 );
and ( n58408 , n58401 , n58406 );
or ( n58409 , n58404 , n58407 , n58408 );
and ( n58410 , n58309 , n58409 );
xor ( n58411 , n58401 , n58403 );
xor ( n58412 , n58411 , n58406 );
and ( n58413 , n56071 , n52540 );
and ( n58414 , n56073 , n52538 );
nor ( n58415 , n58413 , n58414 );
xnor ( n58416 , n58415 , n52424 );
and ( n58417 , n56336 , n52346 );
and ( n58418 , n56338 , n52344 );
nor ( n58419 , n58417 , n58418 );
xnor ( n58420 , n58419 , n52300 );
and ( n58421 , n58416 , n58420 );
and ( n58422 , n56806 , n52318 );
and ( n58423 , n56495 , n52316 );
nor ( n58424 , n58422 , n58423 );
xnor ( n58425 , n58424 , n52213 );
and ( n58426 , n58420 , n58425 );
and ( n58427 , n58416 , n58425 );
or ( n58428 , n58421 , n58426 , n58427 );
and ( n58429 , n55406 , n52886 );
and ( n58430 , n55365 , n52884 );
nor ( n58431 , n58429 , n58430 );
xnor ( n58432 , n58431 , n52657 );
and ( n58433 , n58428 , n58432 );
xor ( n58434 , n58039 , n58043 );
xor ( n58435 , n58434 , n58046 );
and ( n58436 , n58432 , n58435 );
and ( n58437 , n58428 , n58435 );
or ( n58438 , n58433 , n58436 , n58437 );
and ( n58439 , n55661 , n52617 );
and ( n58440 , n55406 , n52615 );
nor ( n58441 , n58439 , n58440 );
xnor ( n58442 , n58441 , n52558 );
and ( n58443 , n58438 , n58442 );
xor ( n58444 , n58049 , n58053 );
xor ( n58445 , n58444 , n58056 );
and ( n58446 , n58442 , n58445 );
and ( n58447 , n58438 , n58445 );
or ( n58448 , n58443 , n58446 , n58447 );
and ( n58449 , n54885 , n53021 );
and ( n58450 , n54767 , n53019 );
nor ( n58451 , n58449 , n58450 );
xnor ( n58452 , n58451 , n52839 );
and ( n58453 , n58448 , n58452 );
xor ( n58454 , n58059 , n58063 );
xor ( n58455 , n58454 , n58066 );
and ( n58456 , n58452 , n58455 );
and ( n58457 , n58448 , n58455 );
or ( n58458 , n58453 , n58456 , n58457 );
and ( n58459 , n53783 , n53739 );
and ( n58460 , n53785 , n53737 );
nor ( n58461 , n58459 , n58460 );
xnor ( n58462 , n58461 , n53315 );
and ( n58463 , n58458 , n58462 );
xor ( n58464 , n58242 , n58246 );
xor ( n58465 , n58464 , n58249 );
and ( n58466 , n58462 , n58465 );
and ( n58467 , n58458 , n58465 );
or ( n58468 , n58463 , n58466 , n58467 );
and ( n58469 , n53150 , n54693 );
and ( n58470 , n52952 , n54691 );
nor ( n58471 , n58469 , n58470 );
xnor ( n58472 , n58471 , n53892 );
and ( n58473 , n58468 , n58472 );
xor ( n58474 , n58252 , n58256 );
xor ( n58475 , n58474 , n58261 );
and ( n58476 , n58472 , n58475 );
and ( n58477 , n58468 , n58475 );
or ( n58478 , n58473 , n58476 , n58477 );
xor ( n58479 , n58264 , n58268 );
xor ( n58480 , n58479 , n58273 );
and ( n58481 , n58478 , n58480 );
xor ( n58482 , n58375 , n58379 );
xor ( n58483 , n58482 , n58382 );
and ( n58484 , n58480 , n58483 );
and ( n58485 , n58478 , n58483 );
or ( n58486 , n58481 , n58484 , n58485 );
xor ( n58487 , n58276 , n58280 );
xor ( n58488 , n58487 , n58283 );
and ( n58489 , n58486 , n58488 );
xor ( n58490 , n58385 , n58389 );
xor ( n58491 , n58490 , n58392 );
and ( n58492 , n58488 , n58491 );
and ( n58493 , n58486 , n58491 );
or ( n58494 , n58489 , n58492 , n58493 );
xor ( n58495 , n57935 , n57937 );
xor ( n58496 , n58495 , n57940 );
and ( n58497 , n58494 , n58496 );
xor ( n58498 , n58363 , n58395 );
xor ( n58499 , n58498 , n58398 );
and ( n58500 , n58496 , n58499 );
and ( n58501 , n58494 , n58499 );
or ( n58502 , n58497 , n58500 , n58501 );
and ( n58503 , n58412 , n58502 );
and ( n58504 , n53895 , n53739 );
and ( n58505 , n53783 , n53737 );
nor ( n58506 , n58504 , n58505 );
xnor ( n58507 , n58506 , n53315 );
and ( n58508 , n54364 , n53455 );
and ( n58509 , n54078 , n53453 );
nor ( n58510 , n58508 , n58509 );
xnor ( n58511 , n58510 , n53159 );
and ( n58512 , n58507 , n58511 );
xor ( n58513 , n58448 , n58452 );
xor ( n58514 , n58513 , n58455 );
and ( n58515 , n58511 , n58514 );
and ( n58516 , n58507 , n58514 );
or ( n58517 , n58512 , n58515 , n58516 );
and ( n58518 , n53499 , n54285 );
and ( n58519 , n53322 , n54283 );
nor ( n58520 , n58518 , n58519 );
xnor ( n58521 , n58520 , n53794 );
and ( n58522 , n58517 , n58521 );
xor ( n58523 , n58313 , n58317 );
xor ( n58524 , n58523 , n58320 );
and ( n58525 , n58521 , n58524 );
and ( n58526 , n58517 , n58524 );
or ( n58527 , n58522 , n58525 , n58526 );
and ( n58528 , n56495 , n52346 );
and ( n58529 , n56336 , n52344 );
nor ( n58530 , n58528 , n58529 );
xnor ( n58531 , n58530 , n52300 );
and ( n58532 , n56855 , n52318 );
and ( n58533 , n56806 , n52316 );
nor ( n58534 , n58532 , n58533 );
xnor ( n58535 , n58534 , n52213 );
and ( n58536 , n58531 , n58535 );
xor ( n58537 , n58161 , n58198 );
xor ( n58538 , n58537 , n58201 );
and ( n58539 , n58535 , n58538 );
and ( n58540 , n58531 , n58538 );
or ( n58541 , n58536 , n58539 , n58540 );
and ( n58542 , n55769 , n52617 );
and ( n58543 , n55720 , n52615 );
nor ( n58544 , n58542 , n58543 );
xnor ( n58545 , n58544 , n52558 );
and ( n58546 , n58541 , n58545 );
xor ( n58547 , n58134 , n58204 );
xor ( n58548 , n58547 , n58207 );
and ( n58549 , n58545 , n58548 );
and ( n58550 , n58541 , n58548 );
or ( n58551 , n58546 , n58549 , n58550 );
and ( n58552 , n55720 , n52617 );
and ( n58553 , n55661 , n52615 );
nor ( n58554 , n58552 , n58553 );
xnor ( n58555 , n58554 , n52558 );
and ( n58556 , n58551 , n58555 );
xor ( n58557 , n58210 , n58214 );
xor ( n58558 , n58557 , n58219 );
and ( n58559 , n58555 , n58558 );
and ( n58560 , n58551 , n58558 );
or ( n58561 , n58556 , n58559 , n58560 );
and ( n58562 , n57970 , n52121 );
and ( n58563 , n57953 , n52119 );
nor ( n58564 , n58562 , n58563 );
xnor ( n58565 , n58564 , n52087 );
and ( n58566 , n58144 , n52092 );
and ( n58567 , n58117 , n52090 );
nor ( n58568 , n58566 , n58567 );
xnor ( n58569 , n58568 , n52072 );
and ( n58570 , n58565 , n58569 );
buf ( n58571 , n51732 );
and ( n58572 , n58571 , n52059 );
and ( n58573 , n58171 , n52057 );
nor ( n58574 , n58572 , n58573 );
not ( n58575 , n58574 );
and ( n58576 , n58569 , n58575 );
and ( n58577 , n58565 , n58575 );
or ( n58578 , n58570 , n58576 , n58577 );
and ( n58579 , n57517 , n52170 );
and ( n58580 , n57519 , n52168 );
nor ( n58581 , n58579 , n58580 );
xnor ( n58582 , n58581 , n52152 );
and ( n58583 , n58578 , n58582 );
xor ( n58584 , n58165 , n58169 );
xor ( n58585 , n58584 , n58175 );
and ( n58586 , n58582 , n58585 );
and ( n58587 , n58578 , n58585 );
or ( n58588 , n58583 , n58586 , n58587 );
and ( n58589 , n57244 , n52318 );
and ( n58590 , n57027 , n52316 );
nor ( n58591 , n58589 , n58590 );
xnor ( n58592 , n58591 , n52213 );
and ( n58593 , n58588 , n58592 );
xor ( n58594 , n58178 , n58182 );
xor ( n58595 , n58594 , n58185 );
and ( n58596 , n58592 , n58595 );
and ( n58597 , n58588 , n58595 );
or ( n58598 , n58593 , n58596 , n58597 );
and ( n58599 , n56806 , n52346 );
and ( n58600 , n56495 , n52344 );
nor ( n58601 , n58599 , n58600 );
xnor ( n58602 , n58601 , n52300 );
and ( n58603 , n58598 , n58602 );
xor ( n58604 , n58188 , n58192 );
xor ( n58605 , n58604 , n58195 );
and ( n58606 , n58602 , n58605 );
and ( n58607 , n58598 , n58605 );
or ( n58608 , n58603 , n58606 , n58607 );
and ( n58609 , n56073 , n52617 );
and ( n58610 , n55769 , n52615 );
nor ( n58611 , n58609 , n58610 );
xnor ( n58612 , n58611 , n52558 );
and ( n58613 , n58608 , n58612 );
and ( n58614 , n56338 , n52540 );
and ( n58615 , n56071 , n52538 );
nor ( n58616 , n58614 , n58615 );
xnor ( n58617 , n58616 , n52424 );
and ( n58618 , n58612 , n58617 );
and ( n58619 , n58608 , n58617 );
or ( n58620 , n58613 , n58618 , n58619 );
and ( n58621 , n55661 , n52886 );
and ( n58622 , n55406 , n52884 );
nor ( n58623 , n58621 , n58622 );
xnor ( n58624 , n58623 , n52657 );
and ( n58625 , n58620 , n58624 );
xor ( n58626 , n58416 , n58420 );
xor ( n58627 , n58626 , n58425 );
and ( n58628 , n58624 , n58627 );
and ( n58629 , n58620 , n58627 );
or ( n58630 , n58625 , n58628 , n58629 );
and ( n58631 , n55199 , n53021 );
and ( n58632 , n55055 , n53019 );
nor ( n58633 , n58631 , n58632 );
xnor ( n58634 , n58633 , n52839 );
and ( n58635 , n58630 , n58634 );
xor ( n58636 , n58428 , n58432 );
xor ( n58637 , n58636 , n58435 );
and ( n58638 , n58634 , n58637 );
and ( n58639 , n58630 , n58637 );
or ( n58640 , n58635 , n58638 , n58639 );
and ( n58641 , n58561 , n58640 );
xor ( n58642 , n58438 , n58442 );
xor ( n58643 , n58642 , n58445 );
and ( n58644 , n58640 , n58643 );
and ( n58645 , n58561 , n58643 );
or ( n58646 , n58641 , n58644 , n58645 );
and ( n58647 , n53785 , n53972 );
and ( n58648 , n53652 , n53970 );
nor ( n58649 , n58647 , n58648 );
xnor ( n58650 , n58649 , n53662 );
and ( n58651 , n58646 , n58650 );
and ( n58652 , n54767 , n53293 );
and ( n58653 , n54715 , n53291 );
nor ( n58654 , n58652 , n58653 );
xnor ( n58655 , n58654 , n52963 );
and ( n58656 , n55055 , n53021 );
and ( n58657 , n54885 , n53019 );
nor ( n58658 , n58656 , n58657 );
xnor ( n58659 , n58658 , n52839 );
and ( n58660 , n58655 , n58659 );
xor ( n58661 , n58222 , n58226 );
xor ( n58662 , n58661 , n58229 );
and ( n58663 , n58659 , n58662 );
and ( n58664 , n58655 , n58662 );
or ( n58665 , n58660 , n58663 , n58664 );
and ( n58666 , n54715 , n53293 );
and ( n58667 , n54466 , n53291 );
nor ( n58668 , n58666 , n58667 );
xnor ( n58669 , n58668 , n52963 );
xor ( n58670 , n58665 , n58669 );
xor ( n58671 , n58232 , n58236 );
xor ( n58672 , n58671 , n58239 );
xor ( n58673 , n58670 , n58672 );
and ( n58674 , n58650 , n58673 );
and ( n58675 , n58646 , n58673 );
or ( n58676 , n58651 , n58674 , n58675 );
and ( n58677 , n52952 , n55033 );
and ( n58678 , n52954 , n55030 );
nor ( n58679 , n58677 , n58678 );
xnor ( n58680 , n58679 , n53885 );
and ( n58681 , n58676 , n58680 );
xor ( n58682 , n58458 , n58462 );
xor ( n58683 , n58682 , n58465 );
and ( n58684 , n58680 , n58683 );
and ( n58685 , n58676 , n58683 );
or ( n58686 , n58681 , n58684 , n58685 );
and ( n58687 , n58527 , n58686 );
xor ( n58688 , n58323 , n58327 );
xor ( n58689 , n58688 , n58332 );
and ( n58690 , n58686 , n58689 );
and ( n58691 , n58527 , n58689 );
or ( n58692 , n58687 , n58690 , n58691 );
and ( n58693 , n58665 , n58669 );
and ( n58694 , n58669 , n58672 );
and ( n58695 , n58665 , n58672 );
or ( n58696 , n58693 , n58694 , n58695 );
and ( n58697 , n53148 , n54693 );
and ( n58698 , n53150 , n54691 );
nor ( n58699 , n58697 , n58698 );
xnor ( n58700 , n58699 , n53892 );
and ( n58701 , n58696 , n58700 );
and ( n58702 , n53652 , n53972 );
and ( n58703 , n53644 , n53970 );
nor ( n58704 , n58702 , n58703 );
xnor ( n58705 , n58704 , n53662 );
and ( n58706 , n58700 , n58705 );
and ( n58707 , n58696 , n58705 );
or ( n58708 , n58701 , n58706 , n58707 );
and ( n58709 , n52954 , n55033 );
and ( n58710 , n52829 , n55030 );
nor ( n58711 , n58709 , n58710 );
xnor ( n58712 , n58711 , n53885 );
and ( n58713 , n58708 , n58712 );
xor ( n58714 , n58367 , n58369 );
xor ( n58715 , n58714 , n58372 );
and ( n58716 , n58712 , n58715 );
and ( n58717 , n58708 , n58715 );
or ( n58718 , n58713 , n58716 , n58717 );
and ( n58719 , n58692 , n58718 );
xor ( n58720 , n58335 , n58339 );
xor ( n58721 , n58720 , n58350 );
and ( n58722 , n58718 , n58721 );
and ( n58723 , n58692 , n58721 );
or ( n58724 , n58719 , n58722 , n58723 );
xor ( n58725 , n58353 , n58357 );
xor ( n58726 , n58725 , n58360 );
and ( n58727 , n58724 , n58726 );
xor ( n58728 , n58486 , n58488 );
xor ( n58729 , n58728 , n58491 );
and ( n58730 , n58726 , n58729 );
and ( n58731 , n58724 , n58729 );
or ( n58732 , n58727 , n58730 , n58731 );
xor ( n58733 , n58494 , n58496 );
xor ( n58734 , n58733 , n58499 );
and ( n58735 , n58732 , n58734 );
xor ( n58736 , n58724 , n58726 );
xor ( n58737 , n58736 , n58729 );
and ( n58738 , n54078 , n53739 );
and ( n58739 , n53895 , n53737 );
nor ( n58740 , n58738 , n58739 );
xnor ( n58741 , n58740 , n53315 );
and ( n58742 , n54466 , n53455 );
and ( n58743 , n54364 , n53453 );
nor ( n58744 , n58742 , n58743 );
xnor ( n58745 , n58744 , n53159 );
and ( n58746 , n58741 , n58745 );
xor ( n58747 , n58655 , n58659 );
xor ( n58748 , n58747 , n58662 );
and ( n58749 , n58745 , n58748 );
and ( n58750 , n58741 , n58748 );
or ( n58751 , n58746 , n58749 , n58750 );
and ( n58752 , n53322 , n54693 );
and ( n58753 , n53148 , n54691 );
nor ( n58754 , n58752 , n58753 );
xnor ( n58755 , n58754 , n53892 );
and ( n58756 , n58751 , n58755 );
and ( n58757 , n53644 , n54285 );
and ( n58758 , n53499 , n54283 );
nor ( n58759 , n58757 , n58758 );
xnor ( n58760 , n58759 , n53794 );
and ( n58761 , n58755 , n58760 );
and ( n58762 , n58751 , n58760 );
or ( n58763 , n58756 , n58761 , n58762 );
xor ( n58764 , n58696 , n58700 );
xor ( n58765 , n58764 , n58705 );
and ( n58766 , n58763 , n58765 );
xor ( n58767 , n58517 , n58521 );
xor ( n58768 , n58767 , n58524 );
and ( n58769 , n58765 , n58768 );
and ( n58770 , n58763 , n58768 );
or ( n58771 , n58766 , n58769 , n58770 );
xor ( n58772 , n58468 , n58472 );
xor ( n58773 , n58772 , n58475 );
and ( n58774 , n58771 , n58773 );
xor ( n58775 , n58708 , n58712 );
xor ( n58776 , n58775 , n58715 );
and ( n58777 , n58773 , n58776 );
and ( n58778 , n58771 , n58776 );
or ( n58779 , n58774 , n58777 , n58778 );
xor ( n58780 , n58478 , n58480 );
xor ( n58781 , n58780 , n58483 );
and ( n58782 , n58779 , n58781 );
xor ( n58783 , n58692 , n58718 );
xor ( n58784 , n58783 , n58721 );
and ( n58785 , n58781 , n58784 );
and ( n58786 , n58779 , n58784 );
or ( n58787 , n58782 , n58785 , n58786 );
and ( n58788 , n58737 , n58787 );
xor ( n58789 , n58779 , n58781 );
xor ( n58790 , n58789 , n58784 );
and ( n58791 , n58117 , n52121 );
and ( n58792 , n57970 , n52119 );
nor ( n58793 , n58791 , n58792 );
xnor ( n58794 , n58793 , n52087 );
and ( n58795 , n58171 , n52092 );
and ( n58796 , n58144 , n52090 );
nor ( n58797 , n58795 , n58796 );
xnor ( n58798 , n58797 , n52072 );
and ( n58799 , n58794 , n58798 );
buf ( n58800 , n51733 );
and ( n58801 , n58800 , n52059 );
and ( n58802 , n58571 , n52057 );
nor ( n58803 , n58801 , n58802 );
not ( n58804 , n58803 );
and ( n58805 , n58798 , n58804 );
and ( n58806 , n58794 , n58804 );
or ( n58807 , n58799 , n58805 , n58806 );
and ( n58808 , n57688 , n52170 );
and ( n58809 , n57517 , n52168 );
nor ( n58810 , n58808 , n58809 );
xnor ( n58811 , n58810 , n52152 );
and ( n58812 , n58807 , n58811 );
xor ( n58813 , n58565 , n58569 );
xor ( n58814 , n58813 , n58575 );
and ( n58815 , n58811 , n58814 );
and ( n58816 , n58807 , n58814 );
or ( n58817 , n58812 , n58815 , n58816 );
and ( n58818 , n57511 , n52318 );
and ( n58819 , n57244 , n52316 );
nor ( n58820 , n58818 , n58819 );
xnor ( n58821 , n58820 , n52213 );
and ( n58822 , n58817 , n58821 );
xor ( n58823 , n58578 , n58582 );
xor ( n58824 , n58823 , n58585 );
and ( n58825 , n58821 , n58824 );
and ( n58826 , n58817 , n58824 );
or ( n58827 , n58822 , n58825 , n58826 );
and ( n58828 , n58144 , n52121 );
and ( n58829 , n58117 , n52119 );
nor ( n58830 , n58828 , n58829 );
xnor ( n58831 , n58830 , n52087 );
and ( n58832 , n58571 , n52092 );
and ( n58833 , n58171 , n52090 );
nor ( n58834 , n58832 , n58833 );
xnor ( n58835 , n58834 , n52072 );
and ( n58836 , n58831 , n58835 );
buf ( n58837 , n51734 );
and ( n58838 , n58837 , n52059 );
and ( n58839 , n58800 , n52057 );
nor ( n58840 , n58838 , n58839 );
not ( n58841 , n58840 );
and ( n58842 , n58835 , n58841 );
and ( n58843 , n58831 , n58841 );
or ( n58844 , n58836 , n58842 , n58843 );
and ( n58845 , n57953 , n52170 );
and ( n58846 , n57688 , n52168 );
nor ( n58847 , n58845 , n58846 );
xnor ( n58848 , n58847 , n52152 );
and ( n58849 , n58844 , n58848 );
xor ( n58850 , n58794 , n58798 );
xor ( n58851 , n58850 , n58804 );
and ( n58852 , n58848 , n58851 );
and ( n58853 , n58844 , n58851 );
or ( n58854 , n58849 , n58852 , n58853 );
and ( n58855 , n58171 , n52121 );
and ( n58856 , n58144 , n52119 );
nor ( n58857 , n58855 , n58856 );
xnor ( n58858 , n58857 , n52087 );
and ( n58859 , n58800 , n52092 );
and ( n58860 , n58571 , n52090 );
nor ( n58861 , n58859 , n58860 );
xnor ( n58862 , n58861 , n52072 );
and ( n58863 , n58858 , n58862 );
buf ( n58864 , n51735 );
and ( n58865 , n58864 , n52059 );
and ( n58866 , n58837 , n52057 );
nor ( n58867 , n58865 , n58866 );
not ( n58868 , n58867 );
and ( n58869 , n58862 , n58868 );
and ( n58870 , n58858 , n58868 );
or ( n58871 , n58863 , n58869 , n58870 );
and ( n58872 , n57970 , n52170 );
and ( n58873 , n57953 , n52168 );
nor ( n58874 , n58872 , n58873 );
xnor ( n58875 , n58874 , n52152 );
and ( n58876 , n58871 , n58875 );
xor ( n58877 , n58831 , n58835 );
xor ( n58878 , n58877 , n58841 );
and ( n58879 , n58875 , n58878 );
and ( n58880 , n58871 , n58878 );
or ( n58881 , n58876 , n58879 , n58880 );
and ( n58882 , n57517 , n52318 );
and ( n58883 , n57519 , n52316 );
nor ( n58884 , n58882 , n58883 );
xnor ( n58885 , n58884 , n52213 );
and ( n58886 , n58881 , n58885 );
xor ( n58887 , n58844 , n58848 );
xor ( n58888 , n58887 , n58851 );
and ( n58889 , n58885 , n58888 );
and ( n58890 , n58881 , n58888 );
or ( n58891 , n58886 , n58889 , n58890 );
and ( n58892 , n58854 , n58891 );
xor ( n58893 , n58807 , n58811 );
xor ( n58894 , n58893 , n58814 );
and ( n58895 , n58891 , n58894 );
and ( n58896 , n58854 , n58894 );
or ( n58897 , n58892 , n58895 , n58896 );
and ( n58898 , n57027 , n52346 );
and ( n58899 , n56855 , n52344 );
nor ( n58900 , n58898 , n58899 );
xnor ( n58901 , n58900 , n52300 );
and ( n58902 , n58897 , n58901 );
xor ( n58903 , n58817 , n58821 );
xor ( n58904 , n58903 , n58824 );
and ( n58905 , n58901 , n58904 );
and ( n58906 , n58897 , n58904 );
or ( n58907 , n58902 , n58905 , n58906 );
and ( n58908 , n58827 , n58907 );
xor ( n58909 , n58588 , n58592 );
xor ( n58910 , n58909 , n58595 );
and ( n58911 , n58907 , n58910 );
and ( n58912 , n58827 , n58910 );
or ( n58913 , n58908 , n58911 , n58912 );
and ( n58914 , n56071 , n52617 );
and ( n58915 , n56073 , n52615 );
nor ( n58916 , n58914 , n58915 );
xnor ( n58917 , n58916 , n52558 );
and ( n58918 , n58913 , n58917 );
and ( n58919 , n56336 , n52540 );
and ( n58920 , n56338 , n52538 );
nor ( n58921 , n58919 , n58920 );
xnor ( n58922 , n58921 , n52424 );
and ( n58923 , n58917 , n58922 );
and ( n58924 , n58913 , n58922 );
or ( n58925 , n58918 , n58923 , n58924 );
and ( n58926 , n55720 , n52886 );
and ( n58927 , n55661 , n52884 );
nor ( n58928 , n58926 , n58927 );
xnor ( n58929 , n58928 , n52657 );
and ( n58930 , n58925 , n58929 );
xor ( n58931 , n58531 , n58535 );
xor ( n58932 , n58931 , n58538 );
and ( n58933 , n58929 , n58932 );
and ( n58934 , n58925 , n58932 );
or ( n58935 , n58930 , n58933 , n58934 );
and ( n58936 , n55365 , n53021 );
and ( n58937 , n55199 , n53019 );
nor ( n58938 , n58936 , n58937 );
xnor ( n58939 , n58938 , n52839 );
and ( n58940 , n58935 , n58939 );
xor ( n58941 , n58541 , n58545 );
xor ( n58942 , n58941 , n58548 );
and ( n58943 , n58939 , n58942 );
and ( n58944 , n58935 , n58942 );
or ( n58945 , n58940 , n58943 , n58944 );
and ( n58946 , n54885 , n53293 );
and ( n58947 , n54767 , n53291 );
nor ( n58948 , n58946 , n58947 );
xnor ( n58949 , n58948 , n52963 );
and ( n58950 , n58945 , n58949 );
xor ( n58951 , n58551 , n58555 );
xor ( n58952 , n58951 , n58558 );
and ( n58953 , n58949 , n58952 );
and ( n58954 , n58945 , n58952 );
or ( n58955 , n58950 , n58953 , n58954 );
and ( n58956 , n53783 , n53972 );
and ( n58957 , n53785 , n53970 );
nor ( n58958 , n58956 , n58957 );
xnor ( n58959 , n58958 , n53662 );
and ( n58960 , n58955 , n58959 );
xor ( n58961 , n58561 , n58640 );
xor ( n58962 , n58961 , n58643 );
and ( n58963 , n58959 , n58962 );
and ( n58964 , n58955 , n58962 );
or ( n58965 , n58960 , n58963 , n58964 );
and ( n58966 , n53150 , n55033 );
and ( n58967 , n52952 , n55030 );
nor ( n58968 , n58966 , n58967 );
xnor ( n58969 , n58968 , n53885 );
and ( n58970 , n58965 , n58969 );
xor ( n58971 , n58507 , n58511 );
xor ( n58972 , n58971 , n58514 );
and ( n58973 , n58969 , n58972 );
and ( n58974 , n58965 , n58972 );
or ( n58975 , n58970 , n58973 , n58974 );
and ( n58976 , n56495 , n52540 );
and ( n58977 , n56336 , n52538 );
nor ( n58978 , n58976 , n58977 );
xnor ( n58979 , n58978 , n52424 );
and ( n58980 , n56855 , n52346 );
and ( n58981 , n56806 , n52344 );
nor ( n58982 , n58980 , n58981 );
xnor ( n58983 , n58982 , n52300 );
and ( n58984 , n58979 , n58983 );
xor ( n58985 , n58827 , n58907 );
xor ( n58986 , n58985 , n58910 );
and ( n58987 , n58983 , n58986 );
and ( n58988 , n58979 , n58986 );
or ( n58989 , n58984 , n58987 , n58988 );
and ( n58990 , n55769 , n52886 );
and ( n58991 , n55720 , n52884 );
nor ( n58992 , n58990 , n58991 );
xnor ( n58993 , n58992 , n52657 );
and ( n58994 , n58989 , n58993 );
xor ( n58995 , n58598 , n58602 );
xor ( n58996 , n58995 , n58605 );
and ( n58997 , n58993 , n58996 );
and ( n58998 , n58989 , n58996 );
or ( n58999 , n58994 , n58997 , n58998 );
and ( n59000 , n55406 , n53021 );
and ( n59001 , n55365 , n53019 );
nor ( n59002 , n59000 , n59001 );
xnor ( n59003 , n59002 , n52839 );
and ( n59004 , n58999 , n59003 );
xor ( n59005 , n58608 , n58612 );
xor ( n59006 , n59005 , n58617 );
and ( n59007 , n59003 , n59006 );
and ( n59008 , n58999 , n59006 );
or ( n59009 , n59004 , n59007 , n59008 );
and ( n59010 , n54767 , n53455 );
and ( n59011 , n54715 , n53453 );
nor ( n59012 , n59010 , n59011 );
xnor ( n59013 , n59012 , n53159 );
and ( n59014 , n59009 , n59013 );
and ( n59015 , n55055 , n53293 );
and ( n59016 , n54885 , n53291 );
nor ( n59017 , n59015 , n59016 );
xnor ( n59018 , n59017 , n52963 );
and ( n59019 , n59013 , n59018 );
and ( n59020 , n59009 , n59018 );
or ( n59021 , n59014 , n59019 , n59020 );
and ( n59022 , n54715 , n53455 );
and ( n59023 , n54466 , n53453 );
nor ( n59024 , n59022 , n59023 );
xnor ( n59025 , n59024 , n53159 );
and ( n59026 , n59021 , n59025 );
xor ( n59027 , n58630 , n58634 );
xor ( n59028 , n59027 , n58637 );
and ( n59029 , n59025 , n59028 );
and ( n59030 , n59021 , n59028 );
or ( n59031 , n59026 , n59029 , n59030 );
and ( n59032 , n53499 , n54693 );
and ( n59033 , n53322 , n54691 );
nor ( n59034 , n59032 , n59033 );
xnor ( n59035 , n59034 , n53892 );
and ( n59036 , n59031 , n59035 );
and ( n59037 , n53652 , n54285 );
and ( n59038 , n53644 , n54283 );
nor ( n59039 , n59037 , n59038 );
xnor ( n59040 , n59039 , n53794 );
and ( n59041 , n59035 , n59040 );
and ( n59042 , n59031 , n59040 );
or ( n59043 , n59036 , n59041 , n59042 );
and ( n59044 , n55365 , n53293 );
and ( n59045 , n55199 , n53291 );
nor ( n59046 , n59044 , n59045 );
xnor ( n59047 , n59046 , n52963 );
and ( n59048 , n55661 , n53021 );
and ( n59049 , n55406 , n53019 );
nor ( n59050 , n59048 , n59049 );
xnor ( n59051 , n59050 , n52839 );
and ( n59052 , n59047 , n59051 );
xor ( n59053 , n58913 , n58917 );
xor ( n59054 , n59053 , n58922 );
and ( n59055 , n59051 , n59054 );
and ( n59056 , n59047 , n59054 );
or ( n59057 , n59052 , n59055 , n59056 );
and ( n59058 , n55199 , n53293 );
and ( n59059 , n55055 , n53291 );
nor ( n59060 , n59058 , n59059 );
xnor ( n59061 , n59060 , n52963 );
and ( n59062 , n59057 , n59061 );
xor ( n59063 , n58925 , n58929 );
xor ( n59064 , n59063 , n58932 );
and ( n59065 , n59061 , n59064 );
and ( n59066 , n59057 , n59064 );
or ( n59067 , n59062 , n59065 , n59066 );
xor ( n59068 , n58620 , n58624 );
xor ( n59069 , n59068 , n58627 );
and ( n59070 , n59067 , n59069 );
xor ( n59071 , n58935 , n58939 );
xor ( n59072 , n59071 , n58942 );
and ( n59073 , n59069 , n59072 );
and ( n59074 , n59067 , n59072 );
or ( n59075 , n59070 , n59073 , n59074 );
and ( n59076 , n54364 , n53739 );
and ( n59077 , n54078 , n53737 );
nor ( n59078 , n59076 , n59077 );
xnor ( n59079 , n59078 , n53315 );
and ( n59080 , n59075 , n59079 );
xor ( n59081 , n58945 , n58949 );
xor ( n59082 , n59081 , n58952 );
and ( n59083 , n59079 , n59082 );
and ( n59084 , n59075 , n59082 );
or ( n59085 , n59080 , n59083 , n59084 );
and ( n59086 , n53148 , n55033 );
and ( n59087 , n53150 , n55030 );
nor ( n59088 , n59086 , n59087 );
xnor ( n59089 , n59088 , n53885 );
and ( n59090 , n59085 , n59089 );
xor ( n59091 , n58741 , n58745 );
xor ( n59092 , n59091 , n58748 );
and ( n59093 , n59089 , n59092 );
and ( n59094 , n59085 , n59092 );
or ( n59095 , n59090 , n59093 , n59094 );
and ( n59096 , n59043 , n59095 );
xor ( n59097 , n58646 , n58650 );
xor ( n59098 , n59097 , n58673 );
and ( n59099 , n59095 , n59098 );
and ( n59100 , n59043 , n59098 );
or ( n59101 , n59096 , n59099 , n59100 );
and ( n59102 , n58975 , n59101 );
xor ( n59103 , n58676 , n58680 );
xor ( n59104 , n59103 , n58683 );
and ( n59105 , n59101 , n59104 );
and ( n59106 , n58975 , n59104 );
or ( n59107 , n59102 , n59105 , n59106 );
xor ( n59108 , n58527 , n58686 );
xor ( n59109 , n59108 , n58689 );
and ( n59110 , n59107 , n59109 );
xor ( n59111 , n58771 , n58773 );
xor ( n59112 , n59111 , n58776 );
and ( n59113 , n59109 , n59112 );
and ( n59114 , n59107 , n59112 );
or ( n59115 , n59110 , n59113 , n59114 );
and ( n59116 , n58790 , n59115 );
xor ( n59117 , n59107 , n59109 );
xor ( n59118 , n59117 , n59112 );
and ( n59119 , n53785 , n54285 );
and ( n59120 , n53652 , n54283 );
nor ( n59121 , n59119 , n59120 );
xnor ( n59122 , n59121 , n53794 );
and ( n59123 , n53895 , n53972 );
and ( n59124 , n53783 , n53970 );
nor ( n59125 , n59123 , n59124 );
xnor ( n59126 , n59125 , n53662 );
and ( n59127 , n59122 , n59126 );
xor ( n59128 , n59021 , n59025 );
xor ( n59129 , n59128 , n59028 );
and ( n59130 , n59126 , n59129 );
and ( n59131 , n59122 , n59129 );
or ( n59132 , n59127 , n59130 , n59131 );
xor ( n59133 , n59031 , n59035 );
xor ( n59134 , n59133 , n59040 );
and ( n59135 , n59132 , n59134 );
xor ( n59136 , n58955 , n58959 );
xor ( n59137 , n59136 , n58962 );
and ( n59138 , n59134 , n59137 );
and ( n59139 , n59132 , n59137 );
or ( n59140 , n59135 , n59138 , n59139 );
xor ( n59141 , n58751 , n58755 );
xor ( n59142 , n59141 , n58760 );
and ( n59143 , n59140 , n59142 );
xor ( n59144 , n58965 , n58969 );
xor ( n59145 , n59144 , n58972 );
and ( n59146 , n59142 , n59145 );
and ( n59147 , n59140 , n59145 );
or ( n59148 , n59143 , n59146 , n59147 );
xor ( n59149 , n58763 , n58765 );
xor ( n59150 , n59149 , n58768 );
and ( n59151 , n59148 , n59150 );
xor ( n59152 , n58975 , n59101 );
xor ( n59153 , n59152 , n59104 );
and ( n59154 , n59150 , n59153 );
and ( n59155 , n59148 , n59153 );
or ( n59156 , n59151 , n59154 , n59155 );
and ( n59157 , n59118 , n59156 );
xor ( n59158 , n59148 , n59150 );
xor ( n59159 , n59158 , n59153 );
and ( n59160 , n54078 , n53972 );
and ( n59161 , n53895 , n53970 );
nor ( n59162 , n59160 , n59161 );
xnor ( n59163 , n59162 , n53662 );
and ( n59164 , n54466 , n53739 );
and ( n59165 , n54364 , n53737 );
nor ( n59166 , n59164 , n59165 );
xnor ( n59167 , n59166 , n53315 );
and ( n59168 , n59163 , n59167 );
xor ( n59169 , n59009 , n59013 );
xor ( n59170 , n59169 , n59018 );
and ( n59171 , n59167 , n59170 );
and ( n59172 , n59163 , n59170 );
or ( n59173 , n59168 , n59171 , n59172 );
and ( n59174 , n53322 , n55033 );
and ( n59175 , n53148 , n55030 );
nor ( n59176 , n59174 , n59175 );
xnor ( n59177 , n59176 , n53885 );
and ( n59178 , n59173 , n59177 );
and ( n59179 , n53644 , n54693 );
and ( n59180 , n53499 , n54691 );
nor ( n59181 , n59179 , n59180 );
xnor ( n59182 , n59181 , n53892 );
and ( n59183 , n59177 , n59182 );
and ( n59184 , n59173 , n59182 );
or ( n59185 , n59178 , n59183 , n59184 );
and ( n59186 , n57244 , n52346 );
and ( n59187 , n57027 , n52344 );
nor ( n59188 , n59186 , n59187 );
xnor ( n59189 , n59188 , n52300 );
and ( n59190 , n57519 , n52318 );
and ( n59191 , n57511 , n52316 );
nor ( n59192 , n59190 , n59191 );
xnor ( n59193 , n59192 , n52213 );
and ( n59194 , n59189 , n59193 );
xor ( n59195 , n58854 , n58891 );
xor ( n59196 , n59195 , n58894 );
and ( n59197 , n59193 , n59196 );
and ( n59198 , n59189 , n59196 );
or ( n59199 , n59194 , n59197 , n59198 );
and ( n59200 , n56336 , n52617 );
and ( n59201 , n56338 , n52615 );
nor ( n59202 , n59200 , n59201 );
xnor ( n59203 , n59202 , n52558 );
and ( n59204 , n59199 , n59203 );
xor ( n59205 , n58897 , n58901 );
xor ( n59206 , n59205 , n58904 );
and ( n59207 , n59203 , n59206 );
and ( n59208 , n59199 , n59206 );
or ( n59209 , n59204 , n59207 , n59208 );
and ( n59210 , n56073 , n52886 );
and ( n59211 , n55769 , n52884 );
nor ( n59212 , n59210 , n59211 );
xnor ( n59213 , n59212 , n52657 );
and ( n59214 , n59209 , n59213 );
and ( n59215 , n56338 , n52617 );
and ( n59216 , n56071 , n52615 );
nor ( n59217 , n59215 , n59216 );
xnor ( n59218 , n59217 , n52558 );
and ( n59219 , n59213 , n59218 );
and ( n59220 , n59209 , n59218 );
or ( n59221 , n59214 , n59219 , n59220 );
and ( n59222 , n58571 , n52121 );
and ( n59223 , n58171 , n52119 );
nor ( n59224 , n59222 , n59223 );
xnor ( n59225 , n59224 , n52087 );
and ( n59226 , n58837 , n52092 );
and ( n59227 , n58800 , n52090 );
nor ( n59228 , n59226 , n59227 );
xnor ( n59229 , n59228 , n52072 );
and ( n59230 , n59225 , n59229 );
and ( n59231 , n58864 , n52057 );
nor ( n59232 , n52059 , n59231 );
not ( n59233 , n59232 );
and ( n59234 , n59229 , n59233 );
and ( n59235 , n59225 , n59233 );
or ( n59236 , n59230 , n59234 , n59235 );
and ( n59237 , n58117 , n52170 );
and ( n59238 , n57970 , n52168 );
nor ( n59239 , n59237 , n59238 );
xnor ( n59240 , n59239 , n52152 );
and ( n59241 , n59236 , n59240 );
xor ( n59242 , n58858 , n58862 );
xor ( n59243 , n59242 , n58868 );
and ( n59244 , n59240 , n59243 );
and ( n59245 , n59236 , n59243 );
or ( n59246 , n59241 , n59244 , n59245 );
and ( n59247 , n57688 , n52318 );
and ( n59248 , n57517 , n52316 );
nor ( n59249 , n59247 , n59248 );
xnor ( n59250 , n59249 , n52213 );
and ( n59251 , n59246 , n59250 );
xor ( n59252 , n58871 , n58875 );
xor ( n59253 , n59252 , n58878 );
and ( n59254 , n59250 , n59253 );
and ( n59255 , n59246 , n59253 );
or ( n59256 , n59251 , n59254 , n59255 );
and ( n59257 , n57511 , n52346 );
and ( n59258 , n57244 , n52344 );
nor ( n59259 , n59257 , n59258 );
xnor ( n59260 , n59259 , n52300 );
and ( n59261 , n59256 , n59260 );
xor ( n59262 , n58881 , n58885 );
xor ( n59263 , n59262 , n58888 );
and ( n59264 , n59260 , n59263 );
and ( n59265 , n59256 , n59263 );
or ( n59266 , n59261 , n59264 , n59265 );
and ( n59267 , n58800 , n52121 );
and ( n59268 , n58571 , n52119 );
nor ( n59269 , n59267 , n59268 );
xnor ( n59270 , n59269 , n52087 );
and ( n59271 , n58864 , n52092 );
and ( n59272 , n58837 , n52090 );
nor ( n59273 , n59271 , n59272 );
xnor ( n59274 , n59273 , n52072 );
and ( n59275 , n59270 , n59274 );
nor ( n59276 , n52059 , n52057 );
not ( n59277 , n59276 );
and ( n59278 , n59274 , n59277 );
and ( n59279 , n59270 , n59277 );
or ( n59280 , n59275 , n59278 , n59279 );
and ( n59281 , n58144 , n52170 );
and ( n59282 , n58117 , n52168 );
nor ( n59283 , n59281 , n59282 );
xnor ( n59284 , n59283 , n52152 );
and ( n59285 , n59280 , n59284 );
xor ( n59286 , n59225 , n59229 );
xor ( n59287 , n59286 , n59233 );
and ( n59288 , n59284 , n59287 );
and ( n59289 , n59280 , n59287 );
or ( n59290 , n59285 , n59288 , n59289 );
and ( n59291 , n57953 , n52318 );
and ( n59292 , n57688 , n52316 );
nor ( n59293 , n59291 , n59292 );
xnor ( n59294 , n59293 , n52213 );
and ( n59295 , n59290 , n59294 );
xor ( n59296 , n59236 , n59240 );
xor ( n59297 , n59296 , n59243 );
and ( n59298 , n59294 , n59297 );
and ( n59299 , n59290 , n59297 );
or ( n59300 , n59295 , n59298 , n59299 );
and ( n59301 , n58837 , n52121 );
and ( n59302 , n58800 , n52119 );
nor ( n59303 , n59301 , n59302 );
xnor ( n59304 , n59303 , n52087 );
and ( n59305 , n58864 , n52090 );
nor ( n59306 , n52092 , n59305 );
xnor ( n59307 , n59306 , n52072 );
and ( n59308 , n59304 , n59307 );
nor ( n59309 , n52059 , n52057 );
not ( n59310 , n59309 );
and ( n59311 , n59307 , n59310 );
and ( n59312 , n59304 , n59310 );
or ( n59313 , n59308 , n59311 , n59312 );
and ( n59314 , n58171 , n52170 );
and ( n59315 , n58144 , n52168 );
nor ( n59316 , n59314 , n59315 );
xnor ( n59317 , n59316 , n52152 );
and ( n59318 , n59313 , n59317 );
xor ( n59319 , n59270 , n59274 );
xor ( n59320 , n59319 , n59277 );
and ( n59321 , n59317 , n59320 );
and ( n59322 , n59313 , n59320 );
or ( n59323 , n59318 , n59321 , n59322 );
and ( n59324 , n58864 , n52119 );
nor ( n59325 , n52121 , n59324 );
xnor ( n59326 , n59325 , n52087 );
nor ( n59327 , n52092 , n52090 );
xnor ( n59328 , n59327 , n52072 );
and ( n59329 , n59326 , n59328 );
nor ( n59330 , n52059 , n52057 );
not ( n59331 , n59330 );
and ( n59332 , n59328 , n59331 );
and ( n59333 , n59326 , n59331 );
or ( n59334 , n59329 , n59332 , n59333 );
nor ( n59335 , n52092 , n52090 );
xnor ( n59336 , n59335 , n52072 );
and ( n59337 , n59334 , n59336 );
nor ( n59338 , n52059 , n52057 );
not ( n59339 , n59338 );
and ( n59340 , n59336 , n59339 );
and ( n59341 , n59334 , n59339 );
or ( n59342 , n59337 , n59340 , n59341 );
and ( n59343 , n58571 , n52170 );
and ( n59344 , n58171 , n52168 );
nor ( n59345 , n59343 , n59344 );
xnor ( n59346 , n59345 , n52152 );
and ( n59347 , n59342 , n59346 );
xor ( n59348 , n59304 , n59307 );
xor ( n59349 , n59348 , n59310 );
and ( n59350 , n59346 , n59349 );
and ( n59351 , n59342 , n59349 );
or ( n59352 , n59347 , n59350 , n59351 );
and ( n59353 , n58117 , n52318 );
and ( n59354 , n57970 , n52316 );
nor ( n59355 , n59353 , n59354 );
xnor ( n59356 , n59355 , n52213 );
and ( n59357 , n59352 , n59356 );
xor ( n59358 , n59313 , n59317 );
xor ( n59359 , n59358 , n59320 );
and ( n59360 , n59356 , n59359 );
and ( n59361 , n59352 , n59359 );
or ( n59362 , n59357 , n59360 , n59361 );
and ( n59363 , n59323 , n59362 );
xor ( n59364 , n59280 , n59284 );
xor ( n59365 , n59364 , n59287 );
and ( n59366 , n59362 , n59365 );
and ( n59367 , n59323 , n59365 );
or ( n59368 , n59363 , n59366 , n59367 );
and ( n59369 , n57517 , n52346 );
and ( n59370 , n57519 , n52344 );
nor ( n59371 , n59369 , n59370 );
xnor ( n59372 , n59371 , n52300 );
and ( n59373 , n59368 , n59372 );
xor ( n59374 , n59290 , n59294 );
xor ( n59375 , n59374 , n59297 );
and ( n59376 , n59372 , n59375 );
and ( n59377 , n59368 , n59375 );
or ( n59378 , n59373 , n59376 , n59377 );
and ( n59379 , n59300 , n59378 );
xor ( n59380 , n59246 , n59250 );
xor ( n59381 , n59380 , n59253 );
and ( n59382 , n59378 , n59381 );
and ( n59383 , n59300 , n59381 );
or ( n59384 , n59379 , n59382 , n59383 );
and ( n59385 , n57027 , n52540 );
and ( n59386 , n56855 , n52538 );
nor ( n59387 , n59385 , n59386 );
xnor ( n59388 , n59387 , n52424 );
and ( n59389 , n59384 , n59388 );
xor ( n59390 , n59256 , n59260 );
xor ( n59391 , n59390 , n59263 );
and ( n59392 , n59388 , n59391 );
and ( n59393 , n59384 , n59391 );
or ( n59394 , n59389 , n59392 , n59393 );
and ( n59395 , n59266 , n59394 );
xor ( n59396 , n59189 , n59193 );
xor ( n59397 , n59396 , n59196 );
and ( n59398 , n59394 , n59397 );
and ( n59399 , n59266 , n59397 );
or ( n59400 , n59395 , n59398 , n59399 );
and ( n59401 , n56071 , n52886 );
and ( n59402 , n56073 , n52884 );
nor ( n59403 , n59401 , n59402 );
xnor ( n59404 , n59403 , n52657 );
and ( n59405 , n59400 , n59404 );
and ( n59406 , n56806 , n52540 );
and ( n59407 , n56495 , n52538 );
nor ( n59408 , n59406 , n59407 );
xnor ( n59409 , n59408 , n52424 );
and ( n59410 , n59404 , n59409 );
and ( n59411 , n59400 , n59409 );
or ( n59412 , n59405 , n59410 , n59411 );
and ( n59413 , n55720 , n53021 );
and ( n59414 , n55661 , n53019 );
nor ( n59415 , n59413 , n59414 );
xnor ( n59416 , n59415 , n52839 );
and ( n59417 , n59412 , n59416 );
xor ( n59418 , n58979 , n58983 );
xor ( n59419 , n59418 , n58986 );
and ( n59420 , n59416 , n59419 );
and ( n59421 , n59412 , n59419 );
or ( n59422 , n59417 , n59420 , n59421 );
and ( n59423 , n59221 , n59422 );
xor ( n59424 , n58989 , n58993 );
xor ( n59425 , n59424 , n58996 );
and ( n59426 , n59422 , n59425 );
and ( n59427 , n59221 , n59425 );
or ( n59428 , n59423 , n59426 , n59427 );
and ( n59429 , n54885 , n53455 );
and ( n59430 , n54767 , n53453 );
nor ( n59431 , n59429 , n59430 );
xnor ( n59432 , n59431 , n53159 );
and ( n59433 , n59428 , n59432 );
xor ( n59434 , n58999 , n59003 );
xor ( n59435 , n59434 , n59006 );
and ( n59436 , n59432 , n59435 );
and ( n59437 , n59428 , n59435 );
or ( n59438 , n59433 , n59436 , n59437 );
and ( n59439 , n53783 , n54285 );
and ( n59440 , n53785 , n54283 );
nor ( n59441 , n59439 , n59440 );
xnor ( n59442 , n59441 , n53794 );
and ( n59443 , n59438 , n59442 );
xor ( n59444 , n59067 , n59069 );
xor ( n59445 , n59444 , n59072 );
and ( n59446 , n59442 , n59445 );
and ( n59447 , n59438 , n59445 );
or ( n59448 , n59443 , n59446 , n59447 );
xor ( n59449 , n59075 , n59079 );
xor ( n59450 , n59449 , n59082 );
and ( n59451 , n59448 , n59450 );
xor ( n59452 , n59122 , n59126 );
xor ( n59453 , n59452 , n59129 );
and ( n59454 , n59450 , n59453 );
and ( n59455 , n59448 , n59453 );
or ( n59456 , n59451 , n59454 , n59455 );
and ( n59457 , n59185 , n59456 );
xor ( n59458 , n59085 , n59089 );
xor ( n59459 , n59458 , n59092 );
and ( n59460 , n59456 , n59459 );
and ( n59461 , n59185 , n59459 );
or ( n59462 , n59457 , n59460 , n59461 );
xor ( n59463 , n59140 , n59142 );
xor ( n59464 , n59463 , n59145 );
and ( n59465 , n59462 , n59464 );
xor ( n59466 , n59043 , n59095 );
xor ( n59467 , n59466 , n59098 );
and ( n59468 , n59464 , n59467 );
and ( n59469 , n59462 , n59467 );
or ( n59470 , n59465 , n59468 , n59469 );
and ( n59471 , n59159 , n59470 );
xor ( n59472 , n59462 , n59464 );
xor ( n59473 , n59472 , n59467 );
and ( n59474 , n56495 , n52617 );
and ( n59475 , n56336 , n52615 );
nor ( n59476 , n59474 , n59475 );
xnor ( n59477 , n59476 , n52558 );
and ( n59478 , n56855 , n52540 );
and ( n59479 , n56806 , n52538 );
nor ( n59480 , n59478 , n59479 );
xnor ( n59481 , n59480 , n52424 );
and ( n59482 , n59477 , n59481 );
xor ( n59483 , n59266 , n59394 );
xor ( n59484 , n59483 , n59397 );
and ( n59485 , n59481 , n59484 );
and ( n59486 , n59477 , n59484 );
or ( n59487 , n59482 , n59485 , n59486 );
and ( n59488 , n55769 , n53021 );
and ( n59489 , n55720 , n53019 );
nor ( n59490 , n59488 , n59489 );
xnor ( n59491 , n59490 , n52839 );
and ( n59492 , n59487 , n59491 );
xor ( n59493 , n59199 , n59203 );
xor ( n59494 , n59493 , n59206 );
and ( n59495 , n59491 , n59494 );
and ( n59496 , n59487 , n59494 );
or ( n59497 , n59492 , n59495 , n59496 );
and ( n59498 , n55406 , n53293 );
and ( n59499 , n55365 , n53291 );
nor ( n59500 , n59498 , n59499 );
xnor ( n59501 , n59500 , n52963 );
and ( n59502 , n59497 , n59501 );
xor ( n59503 , n59209 , n59213 );
xor ( n59504 , n59503 , n59218 );
and ( n59505 , n59501 , n59504 );
and ( n59506 , n59497 , n59504 );
or ( n59507 , n59502 , n59505 , n59506 );
and ( n59508 , n54767 , n53739 );
and ( n59509 , n54715 , n53737 );
nor ( n59510 , n59508 , n59509 );
xnor ( n59511 , n59510 , n53315 );
and ( n59512 , n59507 , n59511 );
xor ( n59513 , n59047 , n59051 );
xor ( n59514 , n59513 , n59054 );
and ( n59515 , n59511 , n59514 );
and ( n59516 , n59507 , n59514 );
or ( n59517 , n59512 , n59515 , n59516 );
and ( n59518 , n54715 , n53739 );
and ( n59519 , n54466 , n53737 );
nor ( n59520 , n59518 , n59519 );
xnor ( n59521 , n59520 , n53315 );
and ( n59522 , n59517 , n59521 );
xor ( n59523 , n59057 , n59061 );
xor ( n59524 , n59523 , n59064 );
and ( n59525 , n59521 , n59524 );
and ( n59526 , n59517 , n59524 );
or ( n59527 , n59522 , n59525 , n59526 );
and ( n59528 , n53499 , n55033 );
and ( n59529 , n53322 , n55030 );
nor ( n59530 , n59528 , n59529 );
xnor ( n59531 , n59530 , n53885 );
and ( n59532 , n59527 , n59531 );
and ( n59533 , n53652 , n54693 );
and ( n59534 , n53644 , n54691 );
nor ( n59535 , n59533 , n59534 );
xnor ( n59536 , n59535 , n53892 );
and ( n59537 , n59531 , n59536 );
and ( n59538 , n59527 , n59536 );
or ( n59539 , n59532 , n59537 , n59538 );
and ( n59540 , n55365 , n53455 );
and ( n59541 , n55199 , n53453 );
nor ( n59542 , n59540 , n59541 );
xnor ( n59543 , n59542 , n53159 );
and ( n59544 , n55661 , n53293 );
and ( n59545 , n55406 , n53291 );
nor ( n59546 , n59544 , n59545 );
xnor ( n59547 , n59546 , n52963 );
and ( n59548 , n59543 , n59547 );
xor ( n59549 , n59400 , n59404 );
xor ( n59550 , n59549 , n59409 );
and ( n59551 , n59547 , n59550 );
and ( n59552 , n59543 , n59550 );
or ( n59553 , n59548 , n59551 , n59552 );
and ( n59554 , n55199 , n53455 );
and ( n59555 , n55055 , n53453 );
nor ( n59556 , n59554 , n59555 );
xnor ( n59557 , n59556 , n53159 );
and ( n59558 , n59553 , n59557 );
xor ( n59559 , n59412 , n59416 );
xor ( n59560 , n59559 , n59419 );
and ( n59561 , n59557 , n59560 );
and ( n59562 , n59553 , n59560 );
or ( n59563 , n59558 , n59561 , n59562 );
and ( n59564 , n55055 , n53455 );
and ( n59565 , n54885 , n53453 );
nor ( n59566 , n59564 , n59565 );
xnor ( n59567 , n59566 , n53159 );
and ( n59568 , n59563 , n59567 );
xor ( n59569 , n59221 , n59422 );
xor ( n59570 , n59569 , n59425 );
and ( n59571 , n59567 , n59570 );
and ( n59572 , n59563 , n59570 );
or ( n59573 , n59568 , n59571 , n59572 );
and ( n59574 , n53895 , n54285 );
and ( n59575 , n53783 , n54283 );
nor ( n59576 , n59574 , n59575 );
xnor ( n59577 , n59576 , n53794 );
and ( n59578 , n59573 , n59577 );
and ( n59579 , n54364 , n53972 );
and ( n59580 , n54078 , n53970 );
nor ( n59581 , n59579 , n59580 );
xnor ( n59582 , n59581 , n53662 );
and ( n59583 , n59577 , n59582 );
and ( n59584 , n59573 , n59582 );
or ( n59585 , n59578 , n59583 , n59584 );
and ( n59586 , n53785 , n54693 );
and ( n59587 , n53652 , n54691 );
nor ( n59588 , n59586 , n59587 );
xnor ( n59589 , n59588 , n53892 );
xor ( n59590 , n59428 , n59432 );
xor ( n59591 , n59590 , n59435 );
and ( n59592 , n59589 , n59591 );
xor ( n59593 , n59517 , n59521 );
xor ( n59594 , n59593 , n59524 );
and ( n59595 , n59591 , n59594 );
and ( n59596 , n59589 , n59594 );
or ( n59597 , n59592 , n59595 , n59596 );
and ( n59598 , n59585 , n59597 );
xor ( n59599 , n59163 , n59167 );
xor ( n59600 , n59599 , n59170 );
and ( n59601 , n59597 , n59600 );
and ( n59602 , n59585 , n59600 );
or ( n59603 , n59598 , n59601 , n59602 );
and ( n59604 , n59539 , n59603 );
xor ( n59605 , n59173 , n59177 );
xor ( n59606 , n59605 , n59182 );
and ( n59607 , n59603 , n59606 );
and ( n59608 , n59539 , n59606 );
or ( n59609 , n59604 , n59607 , n59608 );
xor ( n59610 , n59185 , n59456 );
xor ( n59611 , n59610 , n59459 );
and ( n59612 , n59609 , n59611 );
xor ( n59613 , n59132 , n59134 );
xor ( n59614 , n59613 , n59137 );
and ( n59615 , n59611 , n59614 );
and ( n59616 , n59609 , n59614 );
or ( n59617 , n59612 , n59615 , n59616 );
and ( n59618 , n59473 , n59617 );
xor ( n59619 , n59609 , n59611 );
xor ( n59620 , n59619 , n59614 );
and ( n59621 , n57244 , n52540 );
and ( n59622 , n57027 , n52538 );
nor ( n59623 , n59621 , n59622 );
xnor ( n59624 , n59623 , n52424 );
and ( n59625 , n57519 , n52346 );
and ( n59626 , n57511 , n52344 );
nor ( n59627 , n59625 , n59626 );
xnor ( n59628 , n59627 , n52300 );
and ( n59629 , n59624 , n59628 );
xor ( n59630 , n59300 , n59378 );
xor ( n59631 , n59630 , n59381 );
and ( n59632 , n59628 , n59631 );
and ( n59633 , n59624 , n59631 );
or ( n59634 , n59629 , n59632 , n59633 );
and ( n59635 , n56336 , n52886 );
and ( n59636 , n56338 , n52884 );
nor ( n59637 , n59635 , n59636 );
xnor ( n59638 , n59637 , n52657 );
and ( n59639 , n59634 , n59638 );
xor ( n59640 , n59384 , n59388 );
xor ( n59641 , n59640 , n59391 );
and ( n59642 , n59638 , n59641 );
and ( n59643 , n59634 , n59641 );
or ( n59644 , n59639 , n59642 , n59643 );
and ( n59645 , n56073 , n53021 );
and ( n59646 , n55769 , n53019 );
nor ( n59647 , n59645 , n59646 );
xnor ( n59648 , n59647 , n52839 );
and ( n59649 , n59644 , n59648 );
and ( n59650 , n56338 , n52886 );
and ( n59651 , n56071 , n52884 );
nor ( n59652 , n59650 , n59651 );
xnor ( n59653 , n59652 , n52657 );
and ( n59654 , n59648 , n59653 );
and ( n59655 , n59644 , n59653 );
or ( n59656 , n59649 , n59654 , n59655 );
and ( n59657 , n57688 , n52346 );
and ( n59658 , n57517 , n52344 );
nor ( n59659 , n59657 , n59658 );
xnor ( n59660 , n59659 , n52300 );
and ( n59661 , n57970 , n52318 );
and ( n59662 , n57953 , n52316 );
nor ( n59663 , n59661 , n59662 );
xnor ( n59664 , n59663 , n52213 );
and ( n59665 , n59660 , n59664 );
xor ( n59666 , n59323 , n59362 );
xor ( n59667 , n59666 , n59365 );
and ( n59668 , n59664 , n59667 );
and ( n59669 , n59660 , n59667 );
or ( n59670 , n59665 , n59668 , n59669 );
and ( n59671 , n57511 , n52540 );
and ( n59672 , n57244 , n52538 );
nor ( n59673 , n59671 , n59672 );
xnor ( n59674 , n59673 , n52424 );
and ( n59675 , n59670 , n59674 );
xor ( n59676 , n59368 , n59372 );
xor ( n59677 , n59676 , n59375 );
and ( n59678 , n59674 , n59677 );
and ( n59679 , n59670 , n59677 );
or ( n59680 , n59675 , n59678 , n59679 );
and ( n59681 , n56855 , n52617 );
and ( n59682 , n56806 , n52615 );
nor ( n59683 , n59681 , n59682 );
xnor ( n59684 , n59683 , n52558 );
and ( n59685 , n59680 , n59684 );
xor ( n59686 , n59624 , n59628 );
xor ( n59687 , n59686 , n59631 );
and ( n59688 , n59684 , n59687 );
and ( n59689 , n59680 , n59687 );
or ( n59690 , n59685 , n59688 , n59689 );
and ( n59691 , n56071 , n53021 );
and ( n59692 , n56073 , n53019 );
nor ( n59693 , n59691 , n59692 );
xnor ( n59694 , n59693 , n52839 );
and ( n59695 , n59690 , n59694 );
and ( n59696 , n56806 , n52617 );
and ( n59697 , n56495 , n52615 );
nor ( n59698 , n59696 , n59697 );
xnor ( n59699 , n59698 , n52558 );
and ( n59700 , n59694 , n59699 );
and ( n59701 , n59690 , n59699 );
or ( n59702 , n59695 , n59700 , n59701 );
and ( n59703 , n55406 , n53455 );
and ( n59704 , n55365 , n53453 );
nor ( n59705 , n59703 , n59704 );
xnor ( n59706 , n59705 , n53159 );
and ( n59707 , n59702 , n59706 );
xor ( n59708 , n59477 , n59481 );
xor ( n59709 , n59708 , n59484 );
and ( n59710 , n59706 , n59709 );
and ( n59711 , n59702 , n59709 );
or ( n59712 , n59707 , n59710 , n59711 );
and ( n59713 , n59656 , n59712 );
xor ( n59714 , n59487 , n59491 );
xor ( n59715 , n59714 , n59494 );
and ( n59716 , n59712 , n59715 );
and ( n59717 , n59656 , n59715 );
or ( n59718 , n59713 , n59716 , n59717 );
and ( n59719 , n54885 , n53739 );
and ( n59720 , n54767 , n53737 );
nor ( n59721 , n59719 , n59720 );
xnor ( n59722 , n59721 , n53315 );
and ( n59723 , n59718 , n59722 );
xor ( n59724 , n59497 , n59501 );
xor ( n59725 , n59724 , n59504 );
and ( n59726 , n59722 , n59725 );
and ( n59727 , n59718 , n59725 );
or ( n59728 , n59723 , n59726 , n59727 );
and ( n59729 , n58800 , n52170 );
and ( n59730 , n58571 , n52168 );
nor ( n59731 , n59729 , n59730 );
xnor ( n59732 , n59731 , n52152 );
and ( n59733 , n58864 , n52121 );
and ( n59734 , n58837 , n52119 );
nor ( n59735 , n59733 , n59734 );
xnor ( n59736 , n59735 , n52087 );
and ( n59737 , n59732 , n59736 );
xor ( n59738 , n59334 , n59336 );
xor ( n59739 , n59738 , n59339 );
and ( n59740 , n59736 , n59739 );
and ( n59741 , n59732 , n59739 );
or ( n59742 , n59737 , n59740 , n59741 );
nor ( n59743 , n52121 , n52119 );
xnor ( n59744 , n59743 , n52087 );
nor ( n59745 , n52092 , n52090 );
xnor ( n59746 , n59745 , n52072 );
and ( n59747 , n59744 , n59746 );
nor ( n59748 , n52059 , n52057 );
not ( n59749 , n59748 );
and ( n59750 , n59746 , n59749 );
and ( n59751 , n59744 , n59749 );
or ( n59752 , n59747 , n59750 , n59751 );
and ( n59753 , n58837 , n52170 );
and ( n59754 , n58800 , n52168 );
nor ( n59755 , n59753 , n59754 );
xnor ( n59756 , n59755 , n52152 );
and ( n59757 , n59752 , n59756 );
xor ( n59758 , n59326 , n59328 );
xor ( n59759 , n59758 , n59331 );
and ( n59760 , n59756 , n59759 );
and ( n59761 , n59752 , n59759 );
or ( n59762 , n59757 , n59760 , n59761 );
and ( n59763 , n58864 , n52168 );
nor ( n59764 , n52170 , n59763 );
xnor ( n59765 , n59764 , n52152 );
nor ( n59766 , n52092 , n52090 );
xnor ( n59767 , n59766 , n52072 );
and ( n59768 , n59765 , n59767 );
nor ( n59769 , n52059 , n52057 );
not ( n59770 , n59769 );
and ( n59771 , n59767 , n59770 );
and ( n59772 , n59765 , n59770 );
or ( n59773 , n59768 , n59771 , n59772 );
and ( n59774 , n58864 , n52170 );
and ( n59775 , n58837 , n52168 );
nor ( n59776 , n59774 , n59775 );
xnor ( n59777 , n59776 , n52152 );
and ( n59778 , n59773 , n59777 );
xor ( n59779 , n59744 , n59746 );
xor ( n59780 , n59779 , n59749 );
and ( n59781 , n59777 , n59780 );
and ( n59782 , n59773 , n59780 );
or ( n59783 , n59778 , n59781 , n59782 );
and ( n59784 , n58571 , n52318 );
and ( n59785 , n58171 , n52316 );
nor ( n59786 , n59784 , n59785 );
xnor ( n59787 , n59786 , n52213 );
and ( n59788 , n59783 , n59787 );
xor ( n59789 , n59752 , n59756 );
xor ( n59790 , n59789 , n59759 );
and ( n59791 , n59787 , n59790 );
and ( n59792 , n59783 , n59790 );
or ( n59793 , n59788 , n59791 , n59792 );
and ( n59794 , n59762 , n59793 );
xor ( n59795 , n59732 , n59736 );
xor ( n59796 , n59795 , n59739 );
and ( n59797 , n59793 , n59796 );
and ( n59798 , n59762 , n59796 );
or ( n59799 , n59794 , n59797 , n59798 );
and ( n59800 , n59742 , n59799 );
xor ( n59801 , n59342 , n59346 );
xor ( n59802 , n59801 , n59349 );
and ( n59803 , n59799 , n59802 );
and ( n59804 , n59742 , n59802 );
or ( n59805 , n59800 , n59803 , n59804 );
and ( n59806 , n57953 , n52346 );
and ( n59807 , n57688 , n52344 );
nor ( n59808 , n59806 , n59807 );
xnor ( n59809 , n59808 , n52300 );
and ( n59810 , n59805 , n59809 );
xor ( n59811 , n59352 , n59356 );
xor ( n59812 , n59811 , n59359 );
and ( n59813 , n59809 , n59812 );
and ( n59814 , n59805 , n59812 );
or ( n59815 , n59810 , n59813 , n59814 );
and ( n59816 , n58117 , n52346 );
and ( n59817 , n57970 , n52344 );
nor ( n59818 , n59816 , n59817 );
xnor ( n59819 , n59818 , n52300 );
and ( n59820 , n58171 , n52318 );
and ( n59821 , n58144 , n52316 );
nor ( n59822 , n59820 , n59821 );
xnor ( n59823 , n59822 , n52213 );
and ( n59824 , n59819 , n59823 );
xor ( n59825 , n59762 , n59793 );
xor ( n59826 , n59825 , n59796 );
and ( n59827 , n59823 , n59826 );
and ( n59828 , n59819 , n59826 );
or ( n59829 , n59824 , n59827 , n59828 );
and ( n59830 , n58144 , n52318 );
and ( n59831 , n58117 , n52316 );
nor ( n59832 , n59830 , n59831 );
xnor ( n59833 , n59832 , n52213 );
and ( n59834 , n59829 , n59833 );
xor ( n59835 , n59742 , n59799 );
xor ( n59836 , n59835 , n59802 );
and ( n59837 , n59833 , n59836 );
and ( n59838 , n59829 , n59836 );
or ( n59839 , n59834 , n59837 , n59838 );
and ( n59840 , n57517 , n52540 );
and ( n59841 , n57519 , n52538 );
nor ( n59842 , n59840 , n59841 );
xnor ( n59843 , n59842 , n52424 );
and ( n59844 , n59839 , n59843 );
xor ( n59845 , n59805 , n59809 );
xor ( n59846 , n59845 , n59812 );
and ( n59847 , n59843 , n59846 );
and ( n59848 , n59839 , n59846 );
or ( n59849 , n59844 , n59847 , n59848 );
and ( n59850 , n59815 , n59849 );
xor ( n59851 , n59660 , n59664 );
xor ( n59852 , n59851 , n59667 );
and ( n59853 , n59849 , n59852 );
and ( n59854 , n59815 , n59852 );
or ( n59855 , n59850 , n59853 , n59854 );
and ( n59856 , n57027 , n52617 );
and ( n59857 , n56855 , n52615 );
nor ( n59858 , n59856 , n59857 );
xnor ( n59859 , n59858 , n52558 );
and ( n59860 , n59855 , n59859 );
xor ( n59861 , n59670 , n59674 );
xor ( n59862 , n59861 , n59677 );
and ( n59863 , n59859 , n59862 );
and ( n59864 , n59855 , n59862 );
or ( n59865 , n59860 , n59863 , n59864 );
and ( n59866 , n56495 , n52886 );
and ( n59867 , n56336 , n52884 );
nor ( n59868 , n59866 , n59867 );
xnor ( n59869 , n59868 , n52657 );
and ( n59870 , n59865 , n59869 );
xor ( n59871 , n59680 , n59684 );
xor ( n59872 , n59871 , n59687 );
and ( n59873 , n59869 , n59872 );
and ( n59874 , n59865 , n59872 );
or ( n59875 , n59870 , n59873 , n59874 );
and ( n59876 , n55769 , n53293 );
and ( n59877 , n55720 , n53291 );
nor ( n59878 , n59876 , n59877 );
xnor ( n59879 , n59878 , n52963 );
and ( n59880 , n59875 , n59879 );
xor ( n59881 , n59634 , n59638 );
xor ( n59882 , n59881 , n59641 );
and ( n59883 , n59879 , n59882 );
and ( n59884 , n59875 , n59882 );
or ( n59885 , n59880 , n59883 , n59884 );
and ( n59886 , n55720 , n53293 );
and ( n59887 , n55661 , n53291 );
nor ( n59888 , n59886 , n59887 );
xnor ( n59889 , n59888 , n52963 );
and ( n59890 , n59885 , n59889 );
xor ( n59891 , n59644 , n59648 );
xor ( n59892 , n59891 , n59653 );
and ( n59893 , n59889 , n59892 );
and ( n59894 , n59885 , n59892 );
or ( n59895 , n59890 , n59893 , n59894 );
and ( n59896 , n54767 , n53972 );
and ( n59897 , n54715 , n53970 );
nor ( n59898 , n59896 , n59897 );
xnor ( n59899 , n59898 , n53662 );
and ( n59900 , n59895 , n59899 );
xor ( n59901 , n59543 , n59547 );
xor ( n59902 , n59901 , n59550 );
and ( n59903 , n59899 , n59902 );
and ( n59904 , n59895 , n59902 );
or ( n59905 , n59900 , n59903 , n59904 );
and ( n59906 , n54715 , n53972 );
and ( n59907 , n54466 , n53970 );
nor ( n59908 , n59906 , n59907 );
xnor ( n59909 , n59908 , n53662 );
and ( n59910 , n59905 , n59909 );
xor ( n59911 , n59553 , n59557 );
xor ( n59912 , n59911 , n59560 );
and ( n59913 , n59909 , n59912 );
and ( n59914 , n59905 , n59912 );
or ( n59915 , n59910 , n59913 , n59914 );
and ( n59916 , n59728 , n59915 );
and ( n59917 , n53783 , n54693 );
and ( n59918 , n53785 , n54691 );
nor ( n59919 , n59917 , n59918 );
xnor ( n59920 , n59919 , n53892 );
and ( n59921 , n59915 , n59920 );
and ( n59922 , n59728 , n59920 );
or ( n59923 , n59916 , n59921 , n59922 );
and ( n59924 , n54078 , n54285 );
and ( n59925 , n53895 , n54283 );
nor ( n59926 , n59924 , n59925 );
xnor ( n59927 , n59926 , n53794 );
and ( n59928 , n54466 , n53972 );
and ( n59929 , n54364 , n53970 );
nor ( n59930 , n59928 , n59929 );
xnor ( n59931 , n59930 , n53662 );
and ( n59932 , n59927 , n59931 );
xor ( n59933 , n59507 , n59511 );
xor ( n59934 , n59933 , n59514 );
and ( n59935 , n59931 , n59934 );
and ( n59936 , n59927 , n59934 );
or ( n59937 , n59932 , n59935 , n59936 );
and ( n59938 , n59923 , n59937 );
and ( n59939 , n53644 , n55033 );
and ( n59940 , n53499 , n55030 );
nor ( n59941 , n59939 , n59940 );
xnor ( n59942 , n59941 , n53885 );
and ( n59943 , n59937 , n59942 );
and ( n59944 , n59923 , n59942 );
or ( n59945 , n59938 , n59943 , n59944 );
xor ( n59946 , n59527 , n59531 );
xor ( n59947 , n59946 , n59536 );
and ( n59948 , n59945 , n59947 );
xor ( n59949 , n59438 , n59442 );
xor ( n59950 , n59949 , n59445 );
and ( n59951 , n59947 , n59950 );
and ( n59952 , n59945 , n59950 );
or ( n59953 , n59948 , n59951 , n59952 );
xor ( n59954 , n59539 , n59603 );
xor ( n59955 , n59954 , n59606 );
and ( n59956 , n59953 , n59955 );
xor ( n59957 , n59448 , n59450 );
xor ( n59958 , n59957 , n59453 );
and ( n59959 , n59955 , n59958 );
and ( n59960 , n59953 , n59958 );
or ( n59961 , n59956 , n59959 , n59960 );
and ( n59962 , n59620 , n59961 );
xor ( n59963 , n59953 , n59955 );
xor ( n59964 , n59963 , n59958 );
and ( n59965 , n57244 , n52617 );
and ( n59966 , n57027 , n52615 );
nor ( n59967 , n59965 , n59966 );
xnor ( n59968 , n59967 , n52558 );
and ( n59969 , n57519 , n52540 );
and ( n59970 , n57511 , n52538 );
nor ( n59971 , n59969 , n59970 );
xnor ( n59972 , n59971 , n52424 );
and ( n59973 , n59968 , n59972 );
xor ( n59974 , n59815 , n59849 );
xor ( n59975 , n59974 , n59852 );
and ( n59976 , n59972 , n59975 );
and ( n59977 , n59968 , n59975 );
or ( n59978 , n59973 , n59976 , n59977 );
and ( n59979 , n56336 , n53021 );
and ( n59980 , n56338 , n53019 );
nor ( n59981 , n59979 , n59980 );
xnor ( n59982 , n59981 , n52839 );
and ( n59983 , n59978 , n59982 );
xor ( n59984 , n59855 , n59859 );
xor ( n59985 , n59984 , n59862 );
and ( n59986 , n59982 , n59985 );
and ( n59987 , n59978 , n59985 );
or ( n59988 , n59983 , n59986 , n59987 );
and ( n59989 , n56073 , n53293 );
and ( n59990 , n55769 , n53291 );
nor ( n59991 , n59989 , n59990 );
xnor ( n59992 , n59991 , n52963 );
and ( n59993 , n59988 , n59992 );
and ( n59994 , n56338 , n53021 );
and ( n59995 , n56071 , n53019 );
nor ( n59996 , n59994 , n59995 );
xnor ( n59997 , n59996 , n52839 );
and ( n59998 , n59992 , n59997 );
and ( n59999 , n59988 , n59997 );
or ( n60000 , n59993 , n59998 , n59999 );
and ( n60001 , n55661 , n53455 );
and ( n60002 , n55406 , n53453 );
nor ( n60003 , n60001 , n60002 );
xnor ( n60004 , n60003 , n53159 );
and ( n60005 , n60000 , n60004 );
xor ( n60006 , n59690 , n59694 );
xor ( n60007 , n60006 , n59699 );
and ( n60008 , n60004 , n60007 );
and ( n60009 , n60000 , n60007 );
or ( n60010 , n60005 , n60008 , n60009 );
and ( n60011 , n55199 , n53739 );
and ( n60012 , n55055 , n53737 );
nor ( n60013 , n60011 , n60012 );
xnor ( n60014 , n60013 , n53315 );
and ( n60015 , n60010 , n60014 );
xor ( n60016 , n59702 , n59706 );
xor ( n60017 , n60016 , n59709 );
and ( n60018 , n60014 , n60017 );
and ( n60019 , n60010 , n60017 );
or ( n60020 , n60015 , n60018 , n60019 );
and ( n60021 , n55055 , n53739 );
and ( n60022 , n54885 , n53737 );
nor ( n60023 , n60021 , n60022 );
xnor ( n60024 , n60023 , n53315 );
and ( n60025 , n60020 , n60024 );
xor ( n60026 , n59656 , n59712 );
xor ( n60027 , n60026 , n59715 );
and ( n60028 , n60024 , n60027 );
and ( n60029 , n60020 , n60027 );
or ( n60030 , n60025 , n60028 , n60029 );
and ( n60031 , n53895 , n54693 );
and ( n60032 , n53783 , n54691 );
nor ( n60033 , n60031 , n60032 );
xnor ( n60034 , n60033 , n53892 );
and ( n60035 , n60030 , n60034 );
and ( n60036 , n54364 , n54285 );
and ( n60037 , n54078 , n54283 );
nor ( n60038 , n60036 , n60037 );
xnor ( n60039 , n60038 , n53794 );
and ( n60040 , n60034 , n60039 );
and ( n60041 , n60030 , n60039 );
or ( n60042 , n60035 , n60040 , n60041 );
and ( n60043 , n53652 , n55033 );
and ( n60044 , n53644 , n55030 );
nor ( n60045 , n60043 , n60044 );
xnor ( n60046 , n60045 , n53885 );
and ( n60047 , n60042 , n60046 );
xor ( n60048 , n59563 , n59567 );
xor ( n60049 , n60048 , n59570 );
and ( n60050 , n60046 , n60049 );
and ( n60051 , n60042 , n60049 );
or ( n60052 , n60047 , n60050 , n60051 );
xor ( n60053 , n59573 , n59577 );
xor ( n60054 , n60053 , n59582 );
and ( n60055 , n60052 , n60054 );
xor ( n60056 , n59589 , n59591 );
xor ( n60057 , n60056 , n59594 );
and ( n60058 , n60054 , n60057 );
and ( n60059 , n60052 , n60057 );
or ( n60060 , n60055 , n60058 , n60059 );
xor ( n60061 , n59585 , n59597 );
xor ( n60062 , n60061 , n59600 );
and ( n60063 , n60060 , n60062 );
xor ( n60064 , n59945 , n59947 );
xor ( n60065 , n60064 , n59950 );
and ( n60066 , n60062 , n60065 );
and ( n60067 , n60060 , n60065 );
or ( n60068 , n60063 , n60066 , n60067 );
and ( n60069 , n59964 , n60068 );
xor ( n60070 , n60060 , n60062 );
xor ( n60071 , n60070 , n60065 );
and ( n60072 , n53785 , n55033 );
and ( n60073 , n53652 , n55030 );
nor ( n60074 , n60072 , n60073 );
xnor ( n60075 , n60074 , n53885 );
xor ( n60076 , n59718 , n59722 );
xor ( n60077 , n60076 , n59725 );
and ( n60078 , n60075 , n60077 );
xor ( n60079 , n59905 , n59909 );
xor ( n60080 , n60079 , n59912 );
and ( n60081 , n60077 , n60080 );
and ( n60082 , n60075 , n60080 );
or ( n60083 , n60078 , n60081 , n60082 );
xor ( n60084 , n59728 , n59915 );
xor ( n60085 , n60084 , n59920 );
and ( n60086 , n60083 , n60085 );
xor ( n60087 , n59927 , n59931 );
xor ( n60088 , n60087 , n59934 );
and ( n60089 , n60085 , n60088 );
and ( n60090 , n60083 , n60088 );
or ( n60091 , n60086 , n60089 , n60090 );
xor ( n60092 , n59923 , n59937 );
xor ( n60093 , n60092 , n59942 );
and ( n60094 , n60091 , n60093 );
xor ( n60095 , n60052 , n60054 );
xor ( n60096 , n60095 , n60057 );
and ( n60097 , n60093 , n60096 );
and ( n60098 , n60091 , n60096 );
or ( n60099 , n60094 , n60097 , n60098 );
and ( n60100 , n60071 , n60099 );
xor ( n60101 , n60091 , n60093 );
xor ( n60102 , n60101 , n60096 );
and ( n60103 , n57688 , n52540 );
and ( n60104 , n57517 , n52538 );
nor ( n60105 , n60103 , n60104 );
xnor ( n60106 , n60105 , n52424 );
and ( n60107 , n57970 , n52346 );
and ( n60108 , n57953 , n52344 );
nor ( n60109 , n60107 , n60108 );
xnor ( n60110 , n60109 , n52300 );
and ( n60111 , n60106 , n60110 );
xor ( n60112 , n59829 , n59833 );
xor ( n60113 , n60112 , n59836 );
and ( n60114 , n60110 , n60113 );
and ( n60115 , n60106 , n60113 );
or ( n60116 , n60111 , n60114 , n60115 );
and ( n60117 , n57511 , n52617 );
and ( n60118 , n57244 , n52615 );
nor ( n60119 , n60117 , n60118 );
xnor ( n60120 , n60119 , n52558 );
and ( n60121 , n60116 , n60120 );
xor ( n60122 , n59839 , n59843 );
xor ( n60123 , n60122 , n59846 );
and ( n60124 , n60120 , n60123 );
and ( n60125 , n60116 , n60123 );
or ( n60126 , n60121 , n60124 , n60125 );
nor ( n60127 , n52170 , n52168 );
xnor ( n60128 , n60127 , n52152 );
nor ( n60129 , n52092 , n52090 );
xnor ( n60130 , n60129 , n52072 );
and ( n60131 , n60128 , n60130 );
nor ( n60132 , n52059 , n52057 );
not ( n60133 , n60132 );
and ( n60134 , n60130 , n60133 );
and ( n60135 , n60128 , n60133 );
or ( n60136 , n60131 , n60134 , n60135 );
nor ( n60137 , n52121 , n52119 );
xnor ( n60138 , n60137 , n52087 );
and ( n60139 , n60136 , n60138 );
xor ( n60140 , n59765 , n59767 );
xor ( n60141 , n60140 , n59770 );
and ( n60142 , n60138 , n60141 );
and ( n60143 , n60136 , n60141 );
or ( n60144 , n60139 , n60142 , n60143 );
and ( n60145 , n58800 , n52318 );
and ( n60146 , n58571 , n52316 );
nor ( n60147 , n60145 , n60146 );
xnor ( n60148 , n60147 , n52213 );
and ( n60149 , n60144 , n60148 );
xor ( n60150 , n59773 , n59777 );
xor ( n60151 , n60150 , n59780 );
and ( n60152 , n60148 , n60151 );
and ( n60153 , n60144 , n60151 );
or ( n60154 , n60149 , n60152 , n60153 );
nor ( n60155 , n52170 , n52168 );
xnor ( n60156 , n60155 , n52152 );
nor ( n60157 , n52092 , n52090 );
xnor ( n60158 , n60157 , n52072 );
and ( n60159 , n60156 , n60158 );
and ( n60160 , n60158 , n52057 );
and ( n60161 , n60156 , n52057 );
or ( n60162 , n60159 , n60160 , n60161 );
and ( n60163 , n58864 , n52318 );
and ( n60164 , n58837 , n52316 );
nor ( n60165 , n60163 , n60164 );
xnor ( n60166 , n60165 , n52213 );
and ( n60167 , n60162 , n60166 );
nor ( n60168 , n52121 , n52119 );
xnor ( n60169 , n60168 , n52087 );
and ( n60170 , n60166 , n60169 );
and ( n60171 , n60162 , n60169 );
or ( n60172 , n60167 , n60170 , n60171 );
and ( n60173 , n58837 , n52318 );
and ( n60174 , n58800 , n52316 );
nor ( n60175 , n60173 , n60174 );
xnor ( n60176 , n60175 , n52213 );
and ( n60177 , n60172 , n60176 );
xor ( n60178 , n60136 , n60138 );
xor ( n60179 , n60178 , n60141 );
and ( n60180 , n60176 , n60179 );
and ( n60181 , n60172 , n60179 );
or ( n60182 , n60177 , n60180 , n60181 );
and ( n60183 , n58171 , n52346 );
and ( n60184 , n58144 , n52344 );
nor ( n60185 , n60183 , n60184 );
xnor ( n60186 , n60185 , n52300 );
and ( n60187 , n60182 , n60186 );
xor ( n60188 , n60144 , n60148 );
xor ( n60189 , n60188 , n60151 );
and ( n60190 , n60186 , n60189 );
and ( n60191 , n60182 , n60189 );
or ( n60192 , n60187 , n60190 , n60191 );
and ( n60193 , n60154 , n60192 );
xor ( n60194 , n59783 , n59787 );
xor ( n60195 , n60194 , n59790 );
and ( n60196 , n60192 , n60195 );
and ( n60197 , n60154 , n60195 );
or ( n60198 , n60193 , n60196 , n60197 );
and ( n60199 , n57953 , n52540 );
and ( n60200 , n57688 , n52538 );
nor ( n60201 , n60199 , n60200 );
xnor ( n60202 , n60201 , n52424 );
and ( n60203 , n60198 , n60202 );
xor ( n60204 , n59819 , n59823 );
xor ( n60205 , n60204 , n59826 );
and ( n60206 , n60202 , n60205 );
and ( n60207 , n60198 , n60205 );
or ( n60208 , n60203 , n60206 , n60207 );
and ( n60209 , n57519 , n52617 );
and ( n60210 , n57511 , n52615 );
nor ( n60211 , n60209 , n60210 );
xnor ( n60212 , n60211 , n52558 );
and ( n60213 , n60208 , n60212 );
xor ( n60214 , n60106 , n60110 );
xor ( n60215 , n60214 , n60113 );
and ( n60216 , n60212 , n60215 );
and ( n60217 , n60208 , n60215 );
or ( n60218 , n60213 , n60216 , n60217 );
and ( n60219 , n57027 , n52886 );
and ( n60220 , n56855 , n52884 );
nor ( n60221 , n60219 , n60220 );
xnor ( n60222 , n60221 , n52657 );
and ( n60223 , n60218 , n60222 );
xor ( n60224 , n60116 , n60120 );
xor ( n60225 , n60224 , n60123 );
and ( n60226 , n60222 , n60225 );
and ( n60227 , n60218 , n60225 );
or ( n60228 , n60223 , n60226 , n60227 );
and ( n60229 , n60126 , n60228 );
xor ( n60230 , n59968 , n59972 );
xor ( n60231 , n60230 , n59975 );
and ( n60232 , n60228 , n60231 );
and ( n60233 , n60126 , n60231 );
or ( n60234 , n60229 , n60232 , n60233 );
and ( n60235 , n56071 , n53293 );
and ( n60236 , n56073 , n53291 );
nor ( n60237 , n60235 , n60236 );
xnor ( n60238 , n60237 , n52963 );
and ( n60239 , n60234 , n60238 );
and ( n60240 , n56806 , n52886 );
and ( n60241 , n56495 , n52884 );
nor ( n60242 , n60240 , n60241 );
xnor ( n60243 , n60242 , n52657 );
and ( n60244 , n60238 , n60243 );
and ( n60245 , n60234 , n60243 );
or ( n60246 , n60239 , n60244 , n60245 );
xor ( n60247 , n59988 , n59992 );
xor ( n60248 , n60247 , n59997 );
and ( n60249 , n60246 , n60248 );
xor ( n60250 , n59865 , n59869 );
xor ( n60251 , n60250 , n59872 );
and ( n60252 , n60248 , n60251 );
and ( n60253 , n60246 , n60251 );
or ( n60254 , n60249 , n60252 , n60253 );
and ( n60255 , n55365 , n53739 );
and ( n60256 , n55199 , n53737 );
nor ( n60257 , n60255 , n60256 );
xnor ( n60258 , n60257 , n53315 );
and ( n60259 , n60254 , n60258 );
xor ( n60260 , n59875 , n59879 );
xor ( n60261 , n60260 , n59882 );
and ( n60262 , n60258 , n60261 );
and ( n60263 , n60254 , n60261 );
or ( n60264 , n60259 , n60262 , n60263 );
and ( n60265 , n54885 , n53972 );
and ( n60266 , n54767 , n53970 );
nor ( n60267 , n60265 , n60266 );
xnor ( n60268 , n60267 , n53662 );
and ( n60269 , n60264 , n60268 );
xor ( n60270 , n59885 , n59889 );
xor ( n60271 , n60270 , n59892 );
and ( n60272 , n60268 , n60271 );
and ( n60273 , n60264 , n60271 );
or ( n60274 , n60269 , n60272 , n60273 );
and ( n60275 , n56495 , n53021 );
and ( n60276 , n56336 , n53019 );
nor ( n60277 , n60275 , n60276 );
xnor ( n60278 , n60277 , n52839 );
and ( n60279 , n56855 , n52886 );
and ( n60280 , n56806 , n52884 );
nor ( n60281 , n60279 , n60280 );
xnor ( n60282 , n60281 , n52657 );
and ( n60283 , n60278 , n60282 );
xor ( n60284 , n60126 , n60228 );
xor ( n60285 , n60284 , n60231 );
and ( n60286 , n60282 , n60285 );
and ( n60287 , n60278 , n60285 );
or ( n60288 , n60283 , n60286 , n60287 );
and ( n60289 , n55769 , n53455 );
and ( n60290 , n55720 , n53453 );
nor ( n60291 , n60289 , n60290 );
xnor ( n60292 , n60291 , n53159 );
and ( n60293 , n60288 , n60292 );
xor ( n60294 , n59978 , n59982 );
xor ( n60295 , n60294 , n59985 );
and ( n60296 , n60292 , n60295 );
and ( n60297 , n60288 , n60295 );
or ( n60298 , n60293 , n60296 , n60297 );
and ( n60299 , n55406 , n53739 );
and ( n60300 , n55365 , n53737 );
nor ( n60301 , n60299 , n60300 );
xnor ( n60302 , n60301 , n53315 );
and ( n60303 , n60298 , n60302 );
and ( n60304 , n55720 , n53455 );
and ( n60305 , n55661 , n53453 );
nor ( n60306 , n60304 , n60305 );
xnor ( n60307 , n60306 , n53159 );
and ( n60308 , n60302 , n60307 );
and ( n60309 , n60298 , n60307 );
or ( n60310 , n60303 , n60308 , n60309 );
and ( n60311 , n54767 , n54285 );
and ( n60312 , n54715 , n54283 );
nor ( n60313 , n60311 , n60312 );
xnor ( n60314 , n60313 , n53794 );
and ( n60315 , n60310 , n60314 );
and ( n60316 , n55055 , n53972 );
and ( n60317 , n54885 , n53970 );
nor ( n60318 , n60316 , n60317 );
xnor ( n60319 , n60318 , n53662 );
and ( n60320 , n60314 , n60319 );
and ( n60321 , n60310 , n60319 );
or ( n60322 , n60315 , n60320 , n60321 );
and ( n60323 , n54715 , n54285 );
and ( n60324 , n54466 , n54283 );
nor ( n60325 , n60323 , n60324 );
xnor ( n60326 , n60325 , n53794 );
and ( n60327 , n60322 , n60326 );
xor ( n60328 , n60010 , n60014 );
xor ( n60329 , n60328 , n60017 );
and ( n60330 , n60326 , n60329 );
and ( n60331 , n60322 , n60329 );
or ( n60332 , n60327 , n60330 , n60331 );
and ( n60333 , n60274 , n60332 );
and ( n60334 , n53783 , n55033 );
and ( n60335 , n53785 , n55030 );
nor ( n60336 , n60334 , n60335 );
xnor ( n60337 , n60336 , n53885 );
and ( n60338 , n60332 , n60337 );
and ( n60339 , n60274 , n60337 );
or ( n60340 , n60333 , n60338 , n60339 );
and ( n60341 , n54078 , n54693 );
and ( n60342 , n53895 , n54691 );
nor ( n60343 , n60341 , n60342 );
xnor ( n60344 , n60343 , n53892 );
and ( n60345 , n54466 , n54285 );
and ( n60346 , n54364 , n54283 );
nor ( n60347 , n60345 , n60346 );
xnor ( n60348 , n60347 , n53794 );
and ( n60349 , n60344 , n60348 );
xor ( n60350 , n59895 , n59899 );
xor ( n60351 , n60350 , n59902 );
and ( n60352 , n60348 , n60351 );
and ( n60353 , n60344 , n60351 );
or ( n60354 , n60349 , n60352 , n60353 );
and ( n60355 , n60340 , n60354 );
xor ( n60356 , n60030 , n60034 );
xor ( n60357 , n60356 , n60039 );
and ( n60358 , n60354 , n60357 );
and ( n60359 , n60340 , n60357 );
or ( n60360 , n60355 , n60358 , n60359 );
xor ( n60361 , n60083 , n60085 );
xor ( n60362 , n60361 , n60088 );
and ( n60363 , n60360 , n60362 );
xor ( n60364 , n60042 , n60046 );
xor ( n60365 , n60364 , n60049 );
and ( n60366 , n60362 , n60365 );
and ( n60367 , n60360 , n60365 );
or ( n60368 , n60363 , n60366 , n60367 );
and ( n60369 , n60102 , n60368 );
xor ( n60370 , n60360 , n60362 );
xor ( n60371 , n60370 , n60365 );
and ( n60372 , n53895 , n55033 );
and ( n60373 , n53783 , n55030 );
nor ( n60374 , n60372 , n60373 );
xnor ( n60375 , n60374 , n53885 );
and ( n60376 , n54364 , n54693 );
and ( n60377 , n54078 , n54691 );
nor ( n60378 , n60376 , n60377 );
xnor ( n60379 , n60378 , n53892 );
and ( n60380 , n60375 , n60379 );
xor ( n60381 , n60264 , n60268 );
xor ( n60382 , n60381 , n60271 );
and ( n60383 , n60379 , n60382 );
and ( n60384 , n60375 , n60382 );
or ( n60385 , n60380 , n60383 , n60384 );
xor ( n60386 , n60344 , n60348 );
xor ( n60387 , n60386 , n60351 );
and ( n60388 , n60385 , n60387 );
xor ( n60389 , n60020 , n60024 );
xor ( n60390 , n60389 , n60027 );
and ( n60391 , n60387 , n60390 );
and ( n60392 , n60385 , n60390 );
or ( n60393 , n60388 , n60391 , n60392 );
xor ( n60394 , n60340 , n60354 );
xor ( n60395 , n60394 , n60357 );
and ( n60396 , n60393 , n60395 );
xor ( n60397 , n60075 , n60077 );
xor ( n60398 , n60397 , n60080 );
and ( n60399 , n60395 , n60398 );
and ( n60400 , n60393 , n60398 );
or ( n60401 , n60396 , n60399 , n60400 );
and ( n60402 , n60371 , n60401 );
and ( n60403 , n54078 , n55033 );
and ( n60404 , n53895 , n55030 );
nor ( n60405 , n60403 , n60404 );
xnor ( n60406 , n60405 , n53885 );
and ( n60407 , n54466 , n54693 );
and ( n60408 , n54364 , n54691 );
nor ( n60409 , n60407 , n60408 );
xnor ( n60410 , n60409 , n53892 );
and ( n60411 , n60406 , n60410 );
xor ( n60412 , n60310 , n60314 );
xor ( n60413 , n60412 , n60319 );
and ( n60414 , n60410 , n60413 );
and ( n60415 , n60406 , n60413 );
or ( n60416 , n60411 , n60414 , n60415 );
nor ( n60417 , n52170 , n52168 );
xnor ( n60418 , n60417 , n52152 );
and ( n60419 , n52091 , n52072 );
and ( n60420 , n60418 , n60419 );
and ( n60421 , n58864 , n52316 );
nor ( n60422 , n52318 , n60421 );
xnor ( n60423 , n60422 , n52213 );
and ( n60424 , n60420 , n60423 );
nor ( n60425 , n52121 , n52119 );
xnor ( n60426 , n60425 , n52087 );
and ( n60427 , n60423 , n60426 );
and ( n60428 , n60420 , n60426 );
or ( n60429 , n60424 , n60427 , n60428 );
xor ( n60430 , n60128 , n60130 );
xor ( n60431 , n60430 , n60133 );
and ( n60432 , n60429 , n60431 );
xor ( n60433 , n60162 , n60166 );
xor ( n60434 , n60433 , n60169 );
and ( n60435 , n60431 , n60434 );
and ( n60436 , n60429 , n60434 );
or ( n60437 , n60432 , n60435 , n60436 );
and ( n60438 , n58571 , n52346 );
and ( n60439 , n58171 , n52344 );
nor ( n60440 , n60438 , n60439 );
xnor ( n60441 , n60440 , n52300 );
and ( n60442 , n60437 , n60441 );
xor ( n60443 , n60172 , n60176 );
xor ( n60444 , n60443 , n60179 );
and ( n60445 , n60441 , n60444 );
and ( n60446 , n60437 , n60444 );
or ( n60447 , n60442 , n60445 , n60446 );
and ( n60448 , n58117 , n52540 );
and ( n60449 , n57970 , n52538 );
nor ( n60450 , n60448 , n60449 );
xnor ( n60451 , n60450 , n52424 );
and ( n60452 , n60447 , n60451 );
xor ( n60453 , n60182 , n60186 );
xor ( n60454 , n60453 , n60189 );
and ( n60455 , n60451 , n60454 );
and ( n60456 , n60447 , n60454 );
or ( n60457 , n60452 , n60455 , n60456 );
and ( n60458 , n58144 , n52346 );
and ( n60459 , n58117 , n52344 );
nor ( n60460 , n60458 , n60459 );
xnor ( n60461 , n60460 , n52300 );
and ( n60462 , n60457 , n60461 );
xor ( n60463 , n60154 , n60192 );
xor ( n60464 , n60463 , n60195 );
and ( n60465 , n60461 , n60464 );
and ( n60466 , n60457 , n60464 );
or ( n60467 , n60462 , n60465 , n60466 );
and ( n60468 , n57517 , n52617 );
and ( n60469 , n57519 , n52615 );
nor ( n60470 , n60468 , n60469 );
xnor ( n60471 , n60470 , n52558 );
and ( n60472 , n60467 , n60471 );
xor ( n60473 , n60198 , n60202 );
xor ( n60474 , n60473 , n60205 );
and ( n60475 , n60471 , n60474 );
and ( n60476 , n60467 , n60474 );
or ( n60477 , n60472 , n60475 , n60476 );
and ( n60478 , n57244 , n52886 );
and ( n60479 , n57027 , n52884 );
nor ( n60480 , n60478 , n60479 );
xnor ( n60481 , n60480 , n52657 );
and ( n60482 , n60477 , n60481 );
xor ( n60483 , n60208 , n60212 );
xor ( n60484 , n60483 , n60215 );
and ( n60485 , n60481 , n60484 );
and ( n60486 , n60477 , n60484 );
or ( n60487 , n60482 , n60485 , n60486 );
and ( n60488 , n56806 , n53021 );
and ( n60489 , n56495 , n53019 );
nor ( n60490 , n60488 , n60489 );
xnor ( n60491 , n60490 , n52839 );
and ( n60492 , n60487 , n60491 );
xor ( n60493 , n60218 , n60222 );
xor ( n60494 , n60493 , n60225 );
and ( n60495 , n60491 , n60494 );
and ( n60496 , n60487 , n60494 );
or ( n60497 , n60492 , n60495 , n60496 );
and ( n60498 , n56073 , n53455 );
and ( n60499 , n55769 , n53453 );
nor ( n60500 , n60498 , n60499 );
xnor ( n60501 , n60500 , n53159 );
and ( n60502 , n60497 , n60501 );
and ( n60503 , n56338 , n53293 );
and ( n60504 , n56071 , n53291 );
nor ( n60505 , n60503 , n60504 );
xnor ( n60506 , n60505 , n52963 );
and ( n60507 , n60501 , n60506 );
and ( n60508 , n60497 , n60506 );
or ( n60509 , n60502 , n60507 , n60508 );
and ( n60510 , n55365 , n53972 );
and ( n60511 , n55199 , n53970 );
nor ( n60512 , n60510 , n60511 );
xnor ( n60513 , n60512 , n53662 );
and ( n60514 , n60509 , n60513 );
xor ( n60515 , n60234 , n60238 );
xor ( n60516 , n60515 , n60243 );
and ( n60517 , n60513 , n60516 );
and ( n60518 , n60509 , n60516 );
or ( n60519 , n60514 , n60517 , n60518 );
and ( n60520 , n55199 , n53972 );
and ( n60521 , n55055 , n53970 );
nor ( n60522 , n60520 , n60521 );
xnor ( n60523 , n60522 , n53662 );
and ( n60524 , n60519 , n60523 );
xor ( n60525 , n60246 , n60248 );
xor ( n60526 , n60525 , n60251 );
and ( n60527 , n60523 , n60526 );
and ( n60528 , n60519 , n60526 );
or ( n60529 , n60524 , n60527 , n60528 );
xor ( n60530 , n60000 , n60004 );
xor ( n60531 , n60530 , n60007 );
and ( n60532 , n60529 , n60531 );
xor ( n60533 , n60254 , n60258 );
xor ( n60534 , n60533 , n60261 );
and ( n60535 , n60531 , n60534 );
and ( n60536 , n60529 , n60534 );
or ( n60537 , n60532 , n60535 , n60536 );
and ( n60538 , n60416 , n60537 );
xor ( n60539 , n60322 , n60326 );
xor ( n60540 , n60539 , n60329 );
and ( n60541 , n60537 , n60540 );
and ( n60542 , n60416 , n60540 );
or ( n60543 , n60538 , n60541 , n60542 );
xor ( n60544 , n60274 , n60332 );
xor ( n60545 , n60544 , n60337 );
and ( n60546 , n60543 , n60545 );
xor ( n60547 , n60385 , n60387 );
xor ( n60548 , n60547 , n60390 );
and ( n60549 , n60545 , n60548 );
and ( n60550 , n60543 , n60548 );
or ( n60551 , n60546 , n60549 , n60550 );
xor ( n60552 , n60393 , n60395 );
xor ( n60553 , n60552 , n60398 );
and ( n60554 , n60551 , n60553 );
xor ( n60555 , n60543 , n60545 );
xor ( n60556 , n60555 , n60548 );
and ( n60557 , n57688 , n52617 );
and ( n60558 , n57517 , n52615 );
nor ( n60559 , n60557 , n60558 );
xnor ( n60560 , n60559 , n52558 );
and ( n60561 , n57970 , n52540 );
and ( n60562 , n57953 , n52538 );
nor ( n60563 , n60561 , n60562 );
xnor ( n60564 , n60563 , n52424 );
and ( n60565 , n60560 , n60564 );
xor ( n60566 , n60457 , n60461 );
xor ( n60567 , n60566 , n60464 );
and ( n60568 , n60564 , n60567 );
and ( n60569 , n60560 , n60567 );
or ( n60570 , n60565 , n60568 , n60569 );
and ( n60571 , n57511 , n52886 );
and ( n60572 , n57244 , n52884 );
nor ( n60573 , n60571 , n60572 );
xnor ( n60574 , n60573 , n52657 );
and ( n60575 , n60570 , n60574 );
xor ( n60576 , n60467 , n60471 );
xor ( n60577 , n60576 , n60474 );
and ( n60578 , n60574 , n60577 );
and ( n60579 , n60570 , n60577 );
or ( n60580 , n60575 , n60578 , n60579 );
and ( n60581 , n56855 , n53021 );
and ( n60582 , n56806 , n53019 );
nor ( n60583 , n60581 , n60582 );
xnor ( n60584 , n60583 , n52839 );
and ( n60585 , n60580 , n60584 );
xor ( n60586 , n60477 , n60481 );
xor ( n60587 , n60586 , n60484 );
and ( n60588 , n60584 , n60587 );
and ( n60589 , n60580 , n60587 );
or ( n60590 , n60585 , n60588 , n60589 );
and ( n60591 , n56071 , n53455 );
and ( n60592 , n56073 , n53453 );
nor ( n60593 , n60591 , n60592 );
xnor ( n60594 , n60593 , n53159 );
and ( n60595 , n60590 , n60594 );
and ( n60596 , n56336 , n53293 );
and ( n60597 , n56338 , n53291 );
nor ( n60598 , n60596 , n60597 );
xnor ( n60599 , n60598 , n52963 );
and ( n60600 , n60594 , n60599 );
and ( n60601 , n60590 , n60599 );
or ( n60602 , n60595 , n60600 , n60601 );
and ( n60603 , n55406 , n53972 );
and ( n60604 , n55365 , n53970 );
nor ( n60605 , n60603 , n60604 );
xnor ( n60606 , n60605 , n53662 );
and ( n60607 , n60602 , n60606 );
xor ( n60608 , n60278 , n60282 );
xor ( n60609 , n60608 , n60285 );
and ( n60610 , n60606 , n60609 );
and ( n60611 , n60602 , n60609 );
or ( n60612 , n60607 , n60610 , n60611 );
and ( n60613 , n55661 , n53739 );
and ( n60614 , n55406 , n53737 );
nor ( n60615 , n60613 , n60614 );
xnor ( n60616 , n60615 , n53315 );
and ( n60617 , n60612 , n60616 );
xor ( n60618 , n60288 , n60292 );
xor ( n60619 , n60618 , n60295 );
and ( n60620 , n60616 , n60619 );
and ( n60621 , n60612 , n60619 );
or ( n60622 , n60617 , n60620 , n60621 );
and ( n60623 , n54885 , n54285 );
and ( n60624 , n54767 , n54283 );
nor ( n60625 , n60623 , n60624 );
xnor ( n60626 , n60625 , n53794 );
and ( n60627 , n60622 , n60626 );
xor ( n60628 , n60298 , n60302 );
xor ( n60629 , n60628 , n60307 );
and ( n60630 , n60626 , n60629 );
and ( n60631 , n60622 , n60629 );
or ( n60632 , n60627 , n60630 , n60631 );
and ( n60633 , n54767 , n54693 );
and ( n60634 , n54715 , n54691 );
nor ( n60635 , n60633 , n60634 );
xnor ( n60636 , n60635 , n53892 );
and ( n60637 , n55055 , n54285 );
and ( n60638 , n54885 , n54283 );
nor ( n60639 , n60637 , n60638 );
xnor ( n60640 , n60639 , n53794 );
and ( n60641 , n60636 , n60640 );
xor ( n60642 , n60509 , n60513 );
xor ( n60643 , n60642 , n60516 );
and ( n60644 , n60640 , n60643 );
and ( n60645 , n60636 , n60643 );
or ( n60646 , n60641 , n60644 , n60645 );
and ( n60647 , n54715 , n54693 );
and ( n60648 , n54466 , n54691 );
nor ( n60649 , n60647 , n60648 );
xnor ( n60650 , n60649 , n53892 );
and ( n60651 , n60646 , n60650 );
xor ( n60652 , n60519 , n60523 );
xor ( n60653 , n60652 , n60526 );
and ( n60654 , n60650 , n60653 );
and ( n60655 , n60646 , n60653 );
or ( n60656 , n60651 , n60654 , n60655 );
and ( n60657 , n60632 , n60656 );
xor ( n60658 , n60529 , n60531 );
xor ( n60659 , n60658 , n60534 );
and ( n60660 , n60656 , n60659 );
and ( n60661 , n60632 , n60659 );
or ( n60662 , n60657 , n60660 , n60661 );
xor ( n60663 , n60375 , n60379 );
xor ( n60664 , n60663 , n60382 );
and ( n60665 , n60662 , n60664 );
xor ( n60666 , n60416 , n60537 );
xor ( n60667 , n60666 , n60540 );
and ( n60668 , n60664 , n60667 );
and ( n60669 , n60662 , n60667 );
or ( n60670 , n60665 , n60668 , n60669 );
and ( n60671 , n60556 , n60670 );
xor ( n60672 , n60662 , n60664 );
xor ( n60673 , n60672 , n60667 );
nor ( n60674 , n52318 , n52316 );
xnor ( n60675 , n60674 , n52213 );
nor ( n60676 , n52121 , n52119 );
xnor ( n60677 , n60676 , n52087 );
and ( n60678 , n60675 , n60677 );
nor ( n60679 , n52092 , n52090 );
xnor ( n60680 , n60679 , n52072 );
and ( n60681 , n60677 , n60680 );
and ( n60682 , n60675 , n60680 );
or ( n60683 , n60678 , n60681 , n60682 );
xor ( n60684 , n60156 , n60158 );
xor ( n60685 , n60684 , n52057 );
and ( n60686 , n60683 , n60685 );
xor ( n60687 , n60420 , n60423 );
xor ( n60688 , n60687 , n60426 );
and ( n60689 , n60685 , n60688 );
and ( n60690 , n60683 , n60688 );
or ( n60691 , n60686 , n60689 , n60690 );
and ( n60692 , n58800 , n52346 );
and ( n60693 , n58571 , n52344 );
nor ( n60694 , n60692 , n60693 );
xnor ( n60695 , n60694 , n52300 );
and ( n60696 , n60691 , n60695 );
xor ( n60697 , n60429 , n60431 );
xor ( n60698 , n60697 , n60434 );
and ( n60699 , n60695 , n60698 );
and ( n60700 , n60691 , n60698 );
or ( n60701 , n60696 , n60699 , n60700 );
xor ( n60702 , n60418 , n60419 );
nor ( n60703 , n52170 , n52168 );
xnor ( n60704 , n60703 , n52152 );
nor ( n60705 , n52121 , n52119 );
xnor ( n60706 , n60705 , n52087 );
and ( n60707 , n60704 , n60706 );
and ( n60708 , n60706 , n52090 );
and ( n60709 , n60704 , n52090 );
or ( n60710 , n60707 , n60708 , n60709 );
and ( n60711 , n60702 , n60710 );
and ( n60712 , n58864 , n52346 );
and ( n60713 , n58837 , n52344 );
nor ( n60714 , n60712 , n60713 );
xnor ( n60715 , n60714 , n52300 );
and ( n60716 , n60710 , n60715 );
and ( n60717 , n60702 , n60715 );
or ( n60718 , n60711 , n60716 , n60717 );
and ( n60719 , n58837 , n52346 );
and ( n60720 , n58800 , n52344 );
nor ( n60721 , n60719 , n60720 );
xnor ( n60722 , n60721 , n52300 );
and ( n60723 , n60718 , n60722 );
xor ( n60724 , n60683 , n60685 );
xor ( n60725 , n60724 , n60688 );
and ( n60726 , n60722 , n60725 );
and ( n60727 , n60718 , n60725 );
or ( n60728 , n60723 , n60726 , n60727 );
and ( n60729 , n58171 , n52540 );
and ( n60730 , n58144 , n52538 );
nor ( n60731 , n60729 , n60730 );
xnor ( n60732 , n60731 , n52424 );
and ( n60733 , n60728 , n60732 );
xor ( n60734 , n60691 , n60695 );
xor ( n60735 , n60734 , n60698 );
and ( n60736 , n60732 , n60735 );
and ( n60737 , n60728 , n60735 );
or ( n60738 , n60733 , n60736 , n60737 );
and ( n60739 , n60701 , n60738 );
xor ( n60740 , n60437 , n60441 );
xor ( n60741 , n60740 , n60444 );
and ( n60742 , n60738 , n60741 );
and ( n60743 , n60701 , n60741 );
or ( n60744 , n60739 , n60742 , n60743 );
and ( n60745 , n57953 , n52617 );
and ( n60746 , n57688 , n52615 );
nor ( n60747 , n60745 , n60746 );
xnor ( n60748 , n60747 , n52558 );
and ( n60749 , n60744 , n60748 );
xor ( n60750 , n60447 , n60451 );
xor ( n60751 , n60750 , n60454 );
and ( n60752 , n60748 , n60751 );
and ( n60753 , n60744 , n60751 );
or ( n60754 , n60749 , n60752 , n60753 );
and ( n60755 , n57970 , n52617 );
and ( n60756 , n57953 , n52615 );
nor ( n60757 , n60755 , n60756 );
xnor ( n60758 , n60757 , n52558 );
and ( n60759 , n58144 , n52540 );
and ( n60760 , n58117 , n52538 );
nor ( n60761 , n60759 , n60760 );
xnor ( n60762 , n60761 , n52424 );
and ( n60763 , n60758 , n60762 );
xor ( n60764 , n60701 , n60738 );
xor ( n60765 , n60764 , n60741 );
and ( n60766 , n60762 , n60765 );
and ( n60767 , n60758 , n60765 );
or ( n60768 , n60763 , n60766 , n60767 );
and ( n60769 , n57517 , n52886 );
and ( n60770 , n57519 , n52884 );
nor ( n60771 , n60769 , n60770 );
xnor ( n60772 , n60771 , n52657 );
and ( n60773 , n60768 , n60772 );
xor ( n60774 , n60744 , n60748 );
xor ( n60775 , n60774 , n60751 );
and ( n60776 , n60772 , n60775 );
and ( n60777 , n60768 , n60775 );
or ( n60778 , n60773 , n60776 , n60777 );
and ( n60779 , n60754 , n60778 );
xor ( n60780 , n60560 , n60564 );
xor ( n60781 , n60780 , n60567 );
and ( n60782 , n60778 , n60781 );
and ( n60783 , n60754 , n60781 );
or ( n60784 , n60779 , n60782 , n60783 );
and ( n60785 , n57027 , n53021 );
and ( n60786 , n56855 , n53019 );
nor ( n60787 , n60785 , n60786 );
xnor ( n60788 , n60787 , n52839 );
and ( n60789 , n60784 , n60788 );
xor ( n60790 , n60570 , n60574 );
xor ( n60791 , n60790 , n60577 );
and ( n60792 , n60788 , n60791 );
and ( n60793 , n60784 , n60791 );
or ( n60794 , n60789 , n60792 , n60793 );
and ( n60795 , n56495 , n53293 );
and ( n60796 , n56336 , n53291 );
nor ( n60797 , n60795 , n60796 );
xnor ( n60798 , n60797 , n52963 );
and ( n60799 , n60794 , n60798 );
xor ( n60800 , n60580 , n60584 );
xor ( n60801 , n60800 , n60587 );
and ( n60802 , n60798 , n60801 );
and ( n60803 , n60794 , n60801 );
or ( n60804 , n60799 , n60802 , n60803 );
and ( n60805 , n55769 , n53739 );
and ( n60806 , n55720 , n53737 );
nor ( n60807 , n60805 , n60806 );
xnor ( n60808 , n60807 , n53315 );
and ( n60809 , n60804 , n60808 );
xor ( n60810 , n60487 , n60491 );
xor ( n60811 , n60810 , n60494 );
and ( n60812 , n60808 , n60811 );
and ( n60813 , n60804 , n60811 );
or ( n60814 , n60809 , n60812 , n60813 );
and ( n60815 , n55720 , n53739 );
and ( n60816 , n55661 , n53737 );
nor ( n60817 , n60815 , n60816 );
xnor ( n60818 , n60817 , n53315 );
and ( n60819 , n60814 , n60818 );
xor ( n60820 , n60497 , n60501 );
xor ( n60821 , n60820 , n60506 );
and ( n60822 , n60818 , n60821 );
and ( n60823 , n60814 , n60821 );
or ( n60824 , n60819 , n60822 , n60823 );
and ( n60825 , n57244 , n53021 );
and ( n60826 , n57027 , n53019 );
nor ( n60827 , n60825 , n60826 );
xnor ( n60828 , n60827 , n52839 );
and ( n60829 , n57519 , n52886 );
and ( n60830 , n57511 , n52884 );
nor ( n60831 , n60829 , n60830 );
xnor ( n60832 , n60831 , n52657 );
and ( n60833 , n60828 , n60832 );
xor ( n60834 , n60754 , n60778 );
xor ( n60835 , n60834 , n60781 );
and ( n60836 , n60832 , n60835 );
and ( n60837 , n60828 , n60835 );
or ( n60838 , n60833 , n60836 , n60837 );
and ( n60839 , n56806 , n53293 );
and ( n60840 , n56495 , n53291 );
nor ( n60841 , n60839 , n60840 );
xnor ( n60842 , n60841 , n52963 );
and ( n60843 , n60838 , n60842 );
xor ( n60844 , n60784 , n60788 );
xor ( n60845 , n60844 , n60791 );
and ( n60846 , n60842 , n60845 );
and ( n60847 , n60838 , n60845 );
or ( n60848 , n60843 , n60846 , n60847 );
and ( n60849 , n56073 , n53739 );
and ( n60850 , n55769 , n53737 );
nor ( n60851 , n60849 , n60850 );
xnor ( n60852 , n60851 , n53315 );
and ( n60853 , n60848 , n60852 );
and ( n60854 , n56338 , n53455 );
and ( n60855 , n56071 , n53453 );
nor ( n60856 , n60854 , n60855 );
xnor ( n60857 , n60856 , n53159 );
and ( n60858 , n60852 , n60857 );
and ( n60859 , n60848 , n60857 );
or ( n60860 , n60853 , n60858 , n60859 );
and ( n60861 , n55661 , n53972 );
and ( n60862 , n55406 , n53970 );
nor ( n60863 , n60861 , n60862 );
xnor ( n60864 , n60863 , n53662 );
and ( n60865 , n60860 , n60864 );
xor ( n60866 , n60590 , n60594 );
xor ( n60867 , n60866 , n60599 );
and ( n60868 , n60864 , n60867 );
and ( n60869 , n60860 , n60867 );
or ( n60870 , n60865 , n60868 , n60869 );
and ( n60871 , n55199 , n54285 );
and ( n60872 , n55055 , n54283 );
nor ( n60873 , n60871 , n60872 );
xnor ( n60874 , n60873 , n53794 );
and ( n60875 , n60870 , n60874 );
xor ( n60876 , n60602 , n60606 );
xor ( n60877 , n60876 , n60609 );
and ( n60878 , n60874 , n60877 );
and ( n60879 , n60870 , n60877 );
or ( n60880 , n60875 , n60878 , n60879 );
and ( n60881 , n60824 , n60880 );
xor ( n60882 , n60612 , n60616 );
xor ( n60883 , n60882 , n60619 );
and ( n60884 , n60880 , n60883 );
and ( n60885 , n60824 , n60883 );
or ( n60886 , n60881 , n60884 , n60885 );
and ( n60887 , n54364 , n55033 );
and ( n60888 , n54078 , n55030 );
nor ( n60889 , n60887 , n60888 );
xnor ( n60890 , n60889 , n53885 );
and ( n60891 , n60886 , n60890 );
xor ( n60892 , n60622 , n60626 );
xor ( n60893 , n60892 , n60629 );
and ( n60894 , n60890 , n60893 );
and ( n60895 , n60886 , n60893 );
or ( n60896 , n60891 , n60894 , n60895 );
xor ( n60897 , n60406 , n60410 );
xor ( n60898 , n60897 , n60413 );
and ( n60899 , n60896 , n60898 );
xor ( n60900 , n60632 , n60656 );
xor ( n60901 , n60900 , n60659 );
and ( n60902 , n60898 , n60901 );
and ( n60903 , n60896 , n60901 );
or ( n60904 , n60899 , n60902 , n60903 );
and ( n60905 , n60673 , n60904 );
xor ( n60906 , n60896 , n60898 );
xor ( n60907 , n60906 , n60901 );
nor ( n60908 , n52170 , n52168 );
xnor ( n60909 , n60908 , n52152 );
and ( n60910 , n52120 , n52087 );
and ( n60911 , n60909 , n60910 );
and ( n60912 , n58864 , n52344 );
nor ( n60913 , n52346 , n60912 );
xnor ( n60914 , n60913 , n52300 );
and ( n60915 , n60911 , n60914 );
nor ( n60916 , n52318 , n52316 );
xnor ( n60917 , n60916 , n52213 );
and ( n60918 , n60914 , n60917 );
and ( n60919 , n60911 , n60917 );
or ( n60920 , n60915 , n60918 , n60919 );
xor ( n60921 , n60675 , n60677 );
xor ( n60922 , n60921 , n60680 );
and ( n60923 , n60920 , n60922 );
xor ( n60924 , n60702 , n60710 );
xor ( n60925 , n60924 , n60715 );
and ( n60926 , n60922 , n60925 );
and ( n60927 , n60920 , n60925 );
or ( n60928 , n60923 , n60926 , n60927 );
and ( n60929 , n58571 , n52540 );
and ( n60930 , n58171 , n52538 );
nor ( n60931 , n60929 , n60930 );
xnor ( n60932 , n60931 , n52424 );
and ( n60933 , n60928 , n60932 );
xor ( n60934 , n60718 , n60722 );
xor ( n60935 , n60934 , n60725 );
and ( n60936 , n60932 , n60935 );
and ( n60937 , n60928 , n60935 );
or ( n60938 , n60933 , n60936 , n60937 );
and ( n60939 , n58117 , n52617 );
and ( n60940 , n57970 , n52615 );
nor ( n60941 , n60939 , n60940 );
xnor ( n60942 , n60941 , n52558 );
and ( n60943 , n60938 , n60942 );
xor ( n60944 , n60728 , n60732 );
xor ( n60945 , n60944 , n60735 );
and ( n60946 , n60942 , n60945 );
and ( n60947 , n60938 , n60945 );
or ( n60948 , n60943 , n60946 , n60947 );
and ( n60949 , n57688 , n52886 );
and ( n60950 , n57517 , n52884 );
nor ( n60951 , n60949 , n60950 );
xnor ( n60952 , n60951 , n52657 );
and ( n60953 , n60948 , n60952 );
xor ( n60954 , n60758 , n60762 );
xor ( n60955 , n60954 , n60765 );
and ( n60956 , n60952 , n60955 );
and ( n60957 , n60948 , n60955 );
or ( n60958 , n60953 , n60956 , n60957 );
and ( n60959 , n57511 , n53021 );
and ( n60960 , n57244 , n53019 );
nor ( n60961 , n60959 , n60960 );
xnor ( n60962 , n60961 , n52839 );
and ( n60963 , n60958 , n60962 );
xor ( n60964 , n60768 , n60772 );
xor ( n60965 , n60964 , n60775 );
and ( n60966 , n60962 , n60965 );
and ( n60967 , n60958 , n60965 );
or ( n60968 , n60963 , n60966 , n60967 );
and ( n60969 , n56855 , n53293 );
and ( n60970 , n56806 , n53291 );
nor ( n60971 , n60969 , n60970 );
xnor ( n60972 , n60971 , n52963 );
and ( n60973 , n60968 , n60972 );
xor ( n60974 , n60828 , n60832 );
xor ( n60975 , n60974 , n60835 );
and ( n60976 , n60972 , n60975 );
and ( n60977 , n60968 , n60975 );
or ( n60978 , n60973 , n60976 , n60977 );
and ( n60979 , n56071 , n53739 );
and ( n60980 , n56073 , n53737 );
nor ( n60981 , n60979 , n60980 );
xnor ( n60982 , n60981 , n53315 );
and ( n60983 , n60978 , n60982 );
and ( n60984 , n56336 , n53455 );
and ( n60985 , n56338 , n53453 );
nor ( n60986 , n60984 , n60985 );
xnor ( n60987 , n60986 , n53159 );
and ( n60988 , n60982 , n60987 );
and ( n60989 , n60978 , n60987 );
or ( n60990 , n60983 , n60988 , n60989 );
and ( n60991 , n55406 , n54285 );
and ( n60992 , n55365 , n54283 );
nor ( n60993 , n60991 , n60992 );
xnor ( n60994 , n60993 , n53794 );
and ( n60995 , n60990 , n60994 );
xor ( n60996 , n60794 , n60798 );
xor ( n60997 , n60996 , n60801 );
and ( n60998 , n60994 , n60997 );
and ( n60999 , n60990 , n60997 );
or ( n61000 , n60995 , n60998 , n60999 );
and ( n61001 , n55365 , n54285 );
and ( n61002 , n55199 , n54283 );
nor ( n61003 , n61001 , n61002 );
xnor ( n61004 , n61003 , n53794 );
and ( n61005 , n61000 , n61004 );
xor ( n61006 , n60804 , n60808 );
xor ( n61007 , n61006 , n60811 );
and ( n61008 , n61004 , n61007 );
and ( n61009 , n61000 , n61007 );
or ( n61010 , n61005 , n61008 , n61009 );
and ( n61011 , n54885 , n54693 );
and ( n61012 , n54767 , n54691 );
nor ( n61013 , n61011 , n61012 );
xnor ( n61014 , n61013 , n53892 );
and ( n61015 , n61010 , n61014 );
xor ( n61016 , n60814 , n60818 );
xor ( n61017 , n61016 , n60821 );
and ( n61018 , n61014 , n61017 );
and ( n61019 , n61010 , n61017 );
or ( n61020 , n61015 , n61018 , n61019 );
and ( n61021 , n54466 , n55033 );
and ( n61022 , n54364 , n55030 );
nor ( n61023 , n61021 , n61022 );
xnor ( n61024 , n61023 , n53885 );
and ( n61025 , n61020 , n61024 );
xor ( n61026 , n60636 , n60640 );
xor ( n61027 , n61026 , n60643 );
and ( n61028 , n61024 , n61027 );
and ( n61029 , n61020 , n61027 );
or ( n61030 , n61025 , n61028 , n61029 );
xor ( n61031 , n60886 , n60890 );
xor ( n61032 , n61031 , n60893 );
and ( n61033 , n61030 , n61032 );
xor ( n61034 , n60646 , n60650 );
xor ( n61035 , n61034 , n60653 );
and ( n61036 , n61032 , n61035 );
and ( n61037 , n61030 , n61035 );
or ( n61038 , n61033 , n61036 , n61037 );
and ( n61039 , n60907 , n61038 );
xor ( n61040 , n61030 , n61032 );
xor ( n61041 , n61040 , n61035 );
nor ( n61042 , n52346 , n52344 );
xnor ( n61043 , n61042 , n52300 );
nor ( n61044 , n52318 , n52316 );
xnor ( n61045 , n61044 , n52213 );
and ( n61046 , n61043 , n61045 );
nor ( n61047 , n52121 , n52119 );
xnor ( n61048 , n61047 , n52087 );
and ( n61049 , n61045 , n61048 );
and ( n61050 , n61043 , n61048 );
or ( n61051 , n61046 , n61049 , n61050 );
xor ( n61052 , n60704 , n60706 );
xor ( n61053 , n61052 , n52090 );
and ( n61054 , n61051 , n61053 );
xor ( n61055 , n60911 , n60914 );
xor ( n61056 , n61055 , n60917 );
and ( n61057 , n61053 , n61056 );
and ( n61058 , n61051 , n61056 );
or ( n61059 , n61054 , n61057 , n61058 );
and ( n61060 , n58800 , n52540 );
and ( n61061 , n58571 , n52538 );
nor ( n61062 , n61060 , n61061 );
xnor ( n61063 , n61062 , n52424 );
and ( n61064 , n61059 , n61063 );
xor ( n61065 , n60920 , n60922 );
xor ( n61066 , n61065 , n60925 );
and ( n61067 , n61063 , n61066 );
and ( n61068 , n61059 , n61066 );
or ( n61069 , n61064 , n61067 , n61068 );
and ( n61070 , n58144 , n52617 );
and ( n61071 , n58117 , n52615 );
nor ( n61072 , n61070 , n61071 );
xnor ( n61073 , n61072 , n52558 );
and ( n61074 , n61069 , n61073 );
xor ( n61075 , n60928 , n60932 );
xor ( n61076 , n61075 , n60935 );
and ( n61077 , n61073 , n61076 );
and ( n61078 , n61069 , n61076 );
or ( n61079 , n61074 , n61077 , n61078 );
and ( n61080 , n57953 , n52886 );
and ( n61081 , n57688 , n52884 );
nor ( n61082 , n61080 , n61081 );
xnor ( n61083 , n61082 , n52657 );
and ( n61084 , n61079 , n61083 );
xor ( n61085 , n60938 , n60942 );
xor ( n61086 , n61085 , n60945 );
and ( n61087 , n61083 , n61086 );
and ( n61088 , n61079 , n61086 );
or ( n61089 , n61084 , n61087 , n61088 );
and ( n61090 , n57519 , n53021 );
and ( n61091 , n57511 , n53019 );
nor ( n61092 , n61090 , n61091 );
xnor ( n61093 , n61092 , n52839 );
and ( n61094 , n61089 , n61093 );
xor ( n61095 , n60948 , n60952 );
xor ( n61096 , n61095 , n60955 );
and ( n61097 , n61093 , n61096 );
and ( n61098 , n61089 , n61096 );
or ( n61099 , n61094 , n61097 , n61098 );
and ( n61100 , n57027 , n53293 );
and ( n61101 , n56855 , n53291 );
nor ( n61102 , n61100 , n61101 );
xnor ( n61103 , n61102 , n52963 );
and ( n61104 , n61099 , n61103 );
xor ( n61105 , n60958 , n60962 );
xor ( n61106 , n61105 , n60965 );
and ( n61107 , n61103 , n61106 );
and ( n61108 , n61099 , n61106 );
or ( n61109 , n61104 , n61107 , n61108 );
and ( n61110 , n56495 , n53455 );
and ( n61111 , n56336 , n53453 );
nor ( n61112 , n61110 , n61111 );
xnor ( n61113 , n61112 , n53159 );
and ( n61114 , n61109 , n61113 );
xor ( n61115 , n60968 , n60972 );
xor ( n61116 , n61115 , n60975 );
and ( n61117 , n61113 , n61116 );
and ( n61118 , n61109 , n61116 );
or ( n61119 , n61114 , n61117 , n61118 );
and ( n61120 , n55769 , n53972 );
and ( n61121 , n55720 , n53970 );
nor ( n61122 , n61120 , n61121 );
xnor ( n61123 , n61122 , n53662 );
and ( n61124 , n61119 , n61123 );
xor ( n61125 , n60838 , n60842 );
xor ( n61126 , n61125 , n60845 );
and ( n61127 , n61123 , n61126 );
and ( n61128 , n61119 , n61126 );
or ( n61129 , n61124 , n61127 , n61128 );
and ( n61130 , n55720 , n53972 );
and ( n61131 , n55661 , n53970 );
nor ( n61132 , n61130 , n61131 );
xnor ( n61133 , n61132 , n53662 );
and ( n61134 , n61129 , n61133 );
xor ( n61135 , n60848 , n60852 );
xor ( n61136 , n61135 , n60857 );
and ( n61137 , n61133 , n61136 );
and ( n61138 , n61129 , n61136 );
or ( n61139 , n61134 , n61137 , n61138 );
and ( n61140 , n54767 , n55033 );
and ( n61141 , n54715 , n55030 );
nor ( n61142 , n61140 , n61141 );
xnor ( n61143 , n61142 , n53885 );
and ( n61144 , n61139 , n61143 );
xor ( n61145 , n60860 , n60864 );
xor ( n61146 , n61145 , n60867 );
and ( n61147 , n61143 , n61146 );
and ( n61148 , n61139 , n61146 );
or ( n61149 , n61144 , n61147 , n61148 );
and ( n61150 , n54715 , n55033 );
and ( n61151 , n54466 , n55030 );
nor ( n61152 , n61150 , n61151 );
xnor ( n61153 , n61152 , n53885 );
and ( n61154 , n61149 , n61153 );
xor ( n61155 , n60870 , n60874 );
xor ( n61156 , n61155 , n60877 );
and ( n61157 , n61153 , n61156 );
and ( n61158 , n61149 , n61156 );
or ( n61159 , n61154 , n61157 , n61158 );
xor ( n61160 , n61020 , n61024 );
xor ( n61161 , n61160 , n61027 );
and ( n61162 , n61159 , n61161 );
xor ( n61163 , n60824 , n60880 );
xor ( n61164 , n61163 , n60883 );
and ( n61165 , n61161 , n61164 );
and ( n61166 , n61159 , n61164 );
or ( n61167 , n61162 , n61165 , n61166 );
and ( n61168 , n61041 , n61167 );
xor ( n61169 , n61159 , n61161 );
xor ( n61170 , n61169 , n61164 );
xor ( n61171 , n60909 , n60910 );
and ( n61172 , n58864 , n52538 );
nor ( n61173 , n52540 , n61172 );
xnor ( n61174 , n61173 , n52424 );
nor ( n61175 , n52170 , n52168 );
xnor ( n61176 , n61175 , n52152 );
and ( n61177 , n61174 , n61176 );
and ( n61178 , n61176 , n52119 );
and ( n61179 , n61174 , n52119 );
or ( n61180 , n61177 , n61178 , n61179 );
and ( n61181 , n61171 , n61180 );
and ( n61182 , n58864 , n52540 );
and ( n61183 , n58837 , n52538 );
nor ( n61184 , n61182 , n61183 );
xnor ( n61185 , n61184 , n52424 );
and ( n61186 , n61180 , n61185 );
and ( n61187 , n61171 , n61185 );
or ( n61188 , n61181 , n61186 , n61187 );
and ( n61189 , n58837 , n52540 );
and ( n61190 , n58800 , n52538 );
nor ( n61191 , n61189 , n61190 );
xnor ( n61192 , n61191 , n52424 );
and ( n61193 , n61188 , n61192 );
xor ( n61194 , n61051 , n61053 );
xor ( n61195 , n61194 , n61056 );
and ( n61196 , n61192 , n61195 );
and ( n61197 , n61188 , n61195 );
or ( n61198 , n61193 , n61196 , n61197 );
and ( n61199 , n58171 , n52617 );
and ( n61200 , n58144 , n52615 );
nor ( n61201 , n61199 , n61200 );
xnor ( n61202 , n61201 , n52558 );
and ( n61203 , n61198 , n61202 );
xor ( n61204 , n61059 , n61063 );
xor ( n61205 , n61204 , n61066 );
and ( n61206 , n61202 , n61205 );
and ( n61207 , n61198 , n61205 );
or ( n61208 , n61203 , n61206 , n61207 );
and ( n61209 , n57970 , n52886 );
and ( n61210 , n57953 , n52884 );
nor ( n61211 , n61209 , n61210 );
xnor ( n61212 , n61211 , n52657 );
and ( n61213 , n61208 , n61212 );
xor ( n61214 , n61069 , n61073 );
xor ( n61215 , n61214 , n61076 );
and ( n61216 , n61212 , n61215 );
and ( n61217 , n61208 , n61215 );
or ( n61218 , n61213 , n61216 , n61217 );
and ( n61219 , n57517 , n53021 );
and ( n61220 , n57519 , n53019 );
nor ( n61221 , n61219 , n61220 );
xnor ( n61222 , n61221 , n52839 );
and ( n61223 , n61218 , n61222 );
xor ( n61224 , n61079 , n61083 );
xor ( n61225 , n61224 , n61086 );
and ( n61226 , n61222 , n61225 );
and ( n61227 , n61218 , n61225 );
or ( n61228 , n61223 , n61226 , n61227 );
and ( n61229 , n57244 , n53293 );
and ( n61230 , n57027 , n53291 );
nor ( n61231 , n61229 , n61230 );
xnor ( n61232 , n61231 , n52963 );
and ( n61233 , n61228 , n61232 );
xor ( n61234 , n61089 , n61093 );
xor ( n61235 , n61234 , n61096 );
and ( n61236 , n61232 , n61235 );
and ( n61237 , n61228 , n61235 );
or ( n61238 , n61233 , n61236 , n61237 );
and ( n61239 , n56806 , n53455 );
and ( n61240 , n56495 , n53453 );
nor ( n61241 , n61239 , n61240 );
xnor ( n61242 , n61241 , n53159 );
and ( n61243 , n61238 , n61242 );
xor ( n61244 , n61099 , n61103 );
xor ( n61245 , n61244 , n61106 );
and ( n61246 , n61242 , n61245 );
and ( n61247 , n61238 , n61245 );
or ( n61248 , n61243 , n61246 , n61247 );
and ( n61249 , n56073 , n53972 );
and ( n61250 , n55769 , n53970 );
nor ( n61251 , n61249 , n61250 );
xnor ( n61252 , n61251 , n53662 );
and ( n61253 , n61248 , n61252 );
and ( n61254 , n56338 , n53739 );
and ( n61255 , n56071 , n53737 );
nor ( n61256 , n61254 , n61255 );
xnor ( n61257 , n61256 , n53315 );
and ( n61258 , n61252 , n61257 );
and ( n61259 , n61248 , n61257 );
or ( n61260 , n61253 , n61258 , n61259 );
and ( n61261 , n55365 , n54693 );
and ( n61262 , n55199 , n54691 );
nor ( n61263 , n61261 , n61262 );
xnor ( n61264 , n61263 , n53892 );
and ( n61265 , n61260 , n61264 );
xor ( n61266 , n60978 , n60982 );
xor ( n61267 , n61266 , n60987 );
and ( n61268 , n61264 , n61267 );
and ( n61269 , n61260 , n61267 );
or ( n61270 , n61265 , n61268 , n61269 );
and ( n61271 , n55199 , n54693 );
and ( n61272 , n55055 , n54691 );
nor ( n61273 , n61271 , n61272 );
xnor ( n61274 , n61273 , n53892 );
and ( n61275 , n61270 , n61274 );
xor ( n61276 , n60990 , n60994 );
xor ( n61277 , n61276 , n60997 );
and ( n61278 , n61274 , n61277 );
and ( n61279 , n61270 , n61277 );
or ( n61280 , n61275 , n61278 , n61279 );
and ( n61281 , n55055 , n54693 );
and ( n61282 , n54885 , n54691 );
nor ( n61283 , n61281 , n61282 );
xnor ( n61284 , n61283 , n53892 );
and ( n61285 , n61280 , n61284 );
xor ( n61286 , n61000 , n61004 );
xor ( n61287 , n61286 , n61007 );
and ( n61288 , n61284 , n61287 );
and ( n61289 , n61280 , n61287 );
or ( n61290 , n61285 , n61288 , n61289 );
xor ( n61291 , n61010 , n61014 );
xor ( n61292 , n61291 , n61017 );
and ( n61293 , n61290 , n61292 );
xor ( n61294 , n61149 , n61153 );
xor ( n61295 , n61294 , n61156 );
and ( n61296 , n61292 , n61295 );
and ( n61297 , n61290 , n61295 );
or ( n61298 , n61293 , n61296 , n61297 );
and ( n61299 , n61170 , n61298 );
xor ( n61300 , n61139 , n61143 );
xor ( n61301 , n61300 , n61146 );
xor ( n61302 , n61280 , n61284 );
xor ( n61303 , n61302 , n61287 );
and ( n61304 , n61301 , n61303 );
and ( n61305 , n54885 , n55033 );
and ( n61306 , n54767 , n55030 );
nor ( n61307 , n61305 , n61306 );
xnor ( n61308 , n61307 , n53885 );
xor ( n61309 , n61129 , n61133 );
xor ( n61310 , n61309 , n61136 );
and ( n61311 , n61308 , n61310 );
and ( n61312 , n61303 , n61311 );
and ( n61313 , n61301 , n61311 );
or ( n61314 , n61304 , n61312 , n61313 );
xor ( n61315 , n61290 , n61292 );
xor ( n61316 , n61315 , n61295 );
and ( n61317 , n61314 , n61316 );
and ( n61318 , n55055 , n55033 );
and ( n61319 , n54885 , n55030 );
nor ( n61320 , n61318 , n61319 );
xnor ( n61321 , n61320 , n53885 );
and ( n61322 , n55199 , n55033 );
and ( n61323 , n55055 , n55030 );
nor ( n61324 , n61322 , n61323 );
xnor ( n61325 , n61324 , n53885 );
and ( n61326 , n55720 , n54285 );
and ( n61327 , n55661 , n54283 );
nor ( n61328 , n61326 , n61327 );
xnor ( n61329 , n61328 , n53794 );
and ( n61330 , n61325 , n61329 );
and ( n61331 , n55365 , n55033 );
and ( n61332 , n55199 , n55030 );
nor ( n61333 , n61331 , n61332 );
xnor ( n61334 , n61333 , n53885 );
and ( n61335 , n55661 , n54693 );
and ( n61336 , n55406 , n54691 );
nor ( n61337 , n61335 , n61336 );
xnor ( n61338 , n61337 , n53892 );
and ( n61339 , n61334 , n61338 );
and ( n61340 , n56071 , n53972 );
and ( n61341 , n56073 , n53970 );
nor ( n61342 , n61340 , n61341 );
xnor ( n61343 , n61342 , n53662 );
and ( n61344 , n61338 , n61343 );
and ( n61345 , n61334 , n61343 );
or ( n61346 , n61339 , n61344 , n61345 );
and ( n61347 , n61329 , n61346 );
and ( n61348 , n61325 , n61346 );
or ( n61349 , n61330 , n61347 , n61348 );
and ( n61350 , n61321 , n61349 );
and ( n61351 , n56336 , n53739 );
and ( n61352 , n56338 , n53737 );
nor ( n61353 , n61351 , n61352 );
xnor ( n61354 , n61353 , n53315 );
and ( n61355 , n56495 , n53739 );
and ( n61356 , n56336 , n53737 );
nor ( n61357 , n61355 , n61356 );
xnor ( n61358 , n61357 , n53315 );
and ( n61359 , n56855 , n53455 );
and ( n61360 , n56806 , n53453 );
nor ( n61361 , n61359 , n61360 );
xnor ( n61362 , n61361 , n53159 );
and ( n61363 , n61358 , n61362 );
and ( n61364 , n61354 , n61363 );
and ( n61365 , n56073 , n54285 );
and ( n61366 , n55769 , n54283 );
nor ( n61367 , n61365 , n61366 );
xnor ( n61368 , n61367 , n53794 );
and ( n61369 , n56338 , n53972 );
and ( n61370 , n56071 , n53970 );
nor ( n61371 , n61369 , n61370 );
xnor ( n61372 , n61371 , n53662 );
and ( n61373 , n61368 , n61372 );
and ( n61374 , n61363 , n61373 );
and ( n61375 , n61354 , n61373 );
or ( n61376 , n61364 , n61374 , n61375 );
xor ( n61377 , n61325 , n61329 );
xor ( n61378 , n61377 , n61346 );
and ( n61379 , n61376 , n61378 );
and ( n61380 , n55406 , n55033 );
and ( n61381 , n55365 , n55030 );
nor ( n61382 , n61380 , n61381 );
xnor ( n61383 , n61382 , n53885 );
and ( n61384 , n55720 , n54693 );
and ( n61385 , n55661 , n54691 );
nor ( n61386 , n61384 , n61385 );
xnor ( n61387 , n61386 , n53892 );
and ( n61388 , n61383 , n61387 );
xor ( n61389 , n61334 , n61338 );
xor ( n61390 , n61389 , n61343 );
and ( n61391 , n61388 , n61390 );
xor ( n61392 , n61358 , n61362 );
xor ( n61393 , n61368 , n61372 );
and ( n61394 , n61392 , n61393 );
xor ( n61395 , n61383 , n61387 );
and ( n61396 , n61393 , n61395 );
and ( n61397 , n61392 , n61395 );
or ( n61398 , n61394 , n61396 , n61397 );
and ( n61399 , n61390 , n61398 );
and ( n61400 , n61388 , n61398 );
or ( n61401 , n61391 , n61399 , n61400 );
and ( n61402 , n61378 , n61401 );
and ( n61403 , n61376 , n61401 );
or ( n61404 , n61379 , n61402 , n61403 );
and ( n61405 , n61349 , n61404 );
and ( n61406 , n61321 , n61404 );
or ( n61407 , n61350 , n61405 , n61406 );
xor ( n61408 , n61270 , n61274 );
xor ( n61409 , n61408 , n61277 );
and ( n61410 , n61407 , n61409 );
and ( n61411 , n55661 , n54285 );
and ( n61412 , n55406 , n54283 );
nor ( n61413 , n61411 , n61412 );
xnor ( n61414 , n61413 , n53794 );
xor ( n61415 , n61119 , n61123 );
xor ( n61416 , n61415 , n61126 );
and ( n61417 , n61414 , n61416 );
and ( n61418 , n61409 , n61417 );
and ( n61419 , n61407 , n61417 );
or ( n61420 , n61410 , n61418 , n61419 );
xor ( n61421 , n61321 , n61349 );
xor ( n61422 , n61421 , n61404 );
xor ( n61423 , n61354 , n61363 );
xor ( n61424 , n61423 , n61373 );
and ( n61425 , n55661 , n55033 );
and ( n61426 , n55406 , n55030 );
nor ( n61427 , n61425 , n61426 );
xnor ( n61428 , n61427 , n53885 );
and ( n61429 , n55769 , n54693 );
and ( n61430 , n55720 , n54691 );
nor ( n61431 , n61429 , n61430 );
xnor ( n61432 , n61431 , n53892 );
and ( n61433 , n61428 , n61432 );
and ( n61434 , n56071 , n54285 );
and ( n61435 , n56073 , n54283 );
nor ( n61436 , n61434 , n61435 );
xnor ( n61437 , n61436 , n53794 );
and ( n61438 , n61432 , n61437 );
and ( n61439 , n61428 , n61437 );
or ( n61440 , n61433 , n61438 , n61439 );
and ( n61441 , n56336 , n53972 );
and ( n61442 , n56338 , n53970 );
nor ( n61443 , n61441 , n61442 );
xnor ( n61444 , n61443 , n53662 );
and ( n61445 , n56806 , n53739 );
and ( n61446 , n56495 , n53737 );
nor ( n61447 , n61445 , n61446 );
xnor ( n61448 , n61447 , n53315 );
and ( n61449 , n61444 , n61448 );
and ( n61450 , n57027 , n53455 );
and ( n61451 , n56855 , n53453 );
nor ( n61452 , n61450 , n61451 );
xnor ( n61453 , n61452 , n53159 );
and ( n61454 , n61448 , n61453 );
and ( n61455 , n61444 , n61453 );
or ( n61456 , n61449 , n61454 , n61455 );
and ( n61457 , n61440 , n61456 );
and ( n61458 , n56073 , n54693 );
and ( n61459 , n55769 , n54691 );
nor ( n61460 , n61458 , n61459 );
xnor ( n61461 , n61460 , n53892 );
and ( n61462 , n56338 , n54285 );
and ( n61463 , n56071 , n54283 );
nor ( n61464 , n61462 , n61463 );
xnor ( n61465 , n61464 , n53794 );
and ( n61466 , n61461 , n61465 );
and ( n61467 , n55720 , n55033 );
and ( n61468 , n55661 , n55030 );
nor ( n61469 , n61467 , n61468 );
xnor ( n61470 , n61469 , n53885 );
and ( n61471 , n56495 , n53972 );
and ( n61472 , n56336 , n53970 );
nor ( n61473 , n61471 , n61472 );
xnor ( n61474 , n61473 , n53662 );
and ( n61475 , n61470 , n61474 );
and ( n61476 , n56855 , n53739 );
and ( n61477 , n56806 , n53737 );
nor ( n61478 , n61476 , n61477 );
xnor ( n61479 , n61478 , n53315 );
and ( n61480 , n61474 , n61479 );
and ( n61481 , n61470 , n61479 );
or ( n61482 , n61475 , n61480 , n61481 );
and ( n61483 , n61466 , n61482 );
xor ( n61484 , n61428 , n61432 );
xor ( n61485 , n61484 , n61437 );
and ( n61486 , n61482 , n61485 );
and ( n61487 , n61466 , n61485 );
or ( n61488 , n61483 , n61486 , n61487 );
and ( n61489 , n61456 , n61488 );
and ( n61490 , n61440 , n61488 );
or ( n61491 , n61457 , n61489 , n61490 );
and ( n61492 , n61424 , n61491 );
xor ( n61493 , n61388 , n61390 );
xor ( n61494 , n61493 , n61398 );
and ( n61495 , n61491 , n61494 );
and ( n61496 , n61424 , n61494 );
or ( n61497 , n61492 , n61495 , n61496 );
xor ( n61498 , n61376 , n61378 );
xor ( n61499 , n61498 , n61401 );
and ( n61500 , n61497 , n61499 );
xor ( n61501 , n61392 , n61393 );
xor ( n61502 , n61501 , n61395 );
xor ( n61503 , n61444 , n61448 );
xor ( n61504 , n61503 , n61453 );
and ( n61505 , n57244 , n53455 );
and ( n61506 , n57027 , n53453 );
nor ( n61507 , n61505 , n61506 );
xnor ( n61508 , n61507 , n53159 );
and ( n61509 , n57519 , n53293 );
and ( n61510 , n57511 , n53291 );
nor ( n61511 , n61509 , n61510 );
xnor ( n61512 , n61511 , n52963 );
and ( n61513 , n61508 , n61512 );
xor ( n61514 , n61461 , n61465 );
and ( n61515 , n61512 , n61514 );
and ( n61516 , n61508 , n61514 );
or ( n61517 , n61513 , n61515 , n61516 );
and ( n61518 , n61504 , n61517 );
and ( n61519 , n55769 , n55033 );
and ( n61520 , n55720 , n55030 );
nor ( n61521 , n61519 , n61520 );
xnor ( n61522 , n61521 , n53885 );
and ( n61523 , n56071 , n54693 );
and ( n61524 , n56073 , n54691 );
nor ( n61525 , n61523 , n61524 );
xnor ( n61526 , n61525 , n53892 );
and ( n61527 , n61522 , n61526 );
and ( n61528 , n56336 , n54285 );
and ( n61529 , n56338 , n54283 );
nor ( n61530 , n61528 , n61529 );
xnor ( n61531 , n61530 , n53794 );
and ( n61532 , n61526 , n61531 );
and ( n61533 , n61522 , n61531 );
or ( n61534 , n61527 , n61532 , n61533 );
and ( n61535 , n56806 , n53972 );
and ( n61536 , n56495 , n53970 );
nor ( n61537 , n61535 , n61536 );
xnor ( n61538 , n61537 , n53662 );
and ( n61539 , n57027 , n53739 );
and ( n61540 , n56855 , n53737 );
nor ( n61541 , n61539 , n61540 );
xnor ( n61542 , n61541 , n53315 );
and ( n61543 , n61538 , n61542 );
and ( n61544 , n57511 , n53455 );
and ( n61545 , n57244 , n53453 );
nor ( n61546 , n61544 , n61545 );
xnor ( n61547 , n61546 , n53159 );
and ( n61548 , n61542 , n61547 );
and ( n61549 , n61538 , n61547 );
or ( n61550 , n61543 , n61548 , n61549 );
and ( n61551 , n61534 , n61550 );
xor ( n61552 , n61470 , n61474 );
xor ( n61553 , n61552 , n61479 );
and ( n61554 , n61550 , n61553 );
and ( n61555 , n61534 , n61553 );
or ( n61556 , n61551 , n61554 , n61555 );
and ( n61557 , n61517 , n61556 );
and ( n61558 , n61504 , n61556 );
or ( n61559 , n61518 , n61557 , n61558 );
and ( n61560 , n61502 , n61559 );
xor ( n61561 , n61440 , n61456 );
xor ( n61562 , n61561 , n61488 );
and ( n61563 , n61559 , n61562 );
and ( n61564 , n61502 , n61562 );
or ( n61565 , n61560 , n61563 , n61564 );
xor ( n61566 , n61424 , n61491 );
xor ( n61567 , n61566 , n61494 );
and ( n61568 , n61565 , n61567 );
xor ( n61569 , n61466 , n61482 );
xor ( n61570 , n61569 , n61485 );
and ( n61571 , n57517 , n53293 );
and ( n61572 , n57519 , n53291 );
nor ( n61573 , n61571 , n61572 );
xnor ( n61574 , n61573 , n52963 );
and ( n61575 , n57953 , n53021 );
and ( n61576 , n57688 , n53019 );
nor ( n61577 , n61575 , n61576 );
xnor ( n61578 , n61577 , n52839 );
and ( n61579 , n61574 , n61578 );
and ( n61580 , n57244 , n53739 );
and ( n61581 , n57027 , n53737 );
nor ( n61582 , n61580 , n61581 );
xnor ( n61583 , n61582 , n53315 );
and ( n61584 , n57519 , n53455 );
and ( n61585 , n57511 , n53453 );
nor ( n61586 , n61584 , n61585 );
xnor ( n61587 , n61586 , n53159 );
and ( n61588 , n61583 , n61587 );
and ( n61589 , n61578 , n61588 );
and ( n61590 , n61574 , n61588 );
or ( n61591 , n61579 , n61589 , n61590 );
and ( n61592 , n56495 , n54285 );
and ( n61593 , n56336 , n54283 );
nor ( n61594 , n61592 , n61593 );
xnor ( n61595 , n61594 , n53794 );
and ( n61596 , n56855 , n53972 );
and ( n61597 , n56806 , n53970 );
nor ( n61598 , n61596 , n61597 );
xnor ( n61599 , n61598 , n53662 );
and ( n61600 , n61595 , n61599 );
and ( n61601 , n56073 , n55033 );
and ( n61602 , n55769 , n55030 );
nor ( n61603 , n61601 , n61602 );
xnor ( n61604 , n61603 , n53885 );
and ( n61605 , n56338 , n54693 );
and ( n61606 , n56071 , n54691 );
nor ( n61607 , n61605 , n61606 );
xnor ( n61608 , n61607 , n53892 );
and ( n61609 , n61604 , n61608 );
and ( n61610 , n61600 , n61609 );
and ( n61611 , n57688 , n53293 );
and ( n61612 , n57517 , n53291 );
nor ( n61613 , n61611 , n61612 );
xnor ( n61614 , n61613 , n52963 );
and ( n61615 , n57970 , n53021 );
and ( n61616 , n57953 , n53019 );
nor ( n61617 , n61615 , n61616 );
xnor ( n61618 , n61617 , n52839 );
and ( n61619 , n61614 , n61618 );
and ( n61620 , n58144 , n52886 );
and ( n61621 , n58117 , n52884 );
nor ( n61622 , n61620 , n61621 );
xnor ( n61623 , n61622 , n52657 );
and ( n61624 , n61618 , n61623 );
and ( n61625 , n61614 , n61623 );
or ( n61626 , n61619 , n61624 , n61625 );
and ( n61627 , n61609 , n61626 );
and ( n61628 , n61600 , n61626 );
or ( n61629 , n61610 , n61627 , n61628 );
and ( n61630 , n61591 , n61629 );
xor ( n61631 , n61508 , n61512 );
xor ( n61632 , n61631 , n61514 );
and ( n61633 , n61629 , n61632 );
and ( n61634 , n61591 , n61632 );
or ( n61635 , n61630 , n61633 , n61634 );
and ( n61636 , n61570 , n61635 );
xor ( n61637 , n61504 , n61517 );
xor ( n61638 , n61637 , n61556 );
and ( n61639 , n61635 , n61638 );
and ( n61640 , n61570 , n61638 );
or ( n61641 , n61636 , n61639 , n61640 );
xor ( n61642 , n61502 , n61559 );
xor ( n61643 , n61642 , n61562 );
and ( n61644 , n61641 , n61643 );
xor ( n61645 , n61534 , n61550 );
xor ( n61646 , n61645 , n61553 );
xor ( n61647 , n61522 , n61526 );
xor ( n61648 , n61647 , n61531 );
xor ( n61649 , n61538 , n61542 );
xor ( n61650 , n61649 , n61547 );
and ( n61651 , n61648 , n61650 );
xor ( n61652 , n61583 , n61587 );
xor ( n61653 , n61595 , n61599 );
and ( n61654 , n61652 , n61653 );
xor ( n61655 , n61604 , n61608 );
and ( n61656 , n61653 , n61655 );
and ( n61657 , n61652 , n61655 );
or ( n61658 , n61654 , n61656 , n61657 );
and ( n61659 , n61650 , n61658 );
and ( n61660 , n61648 , n61658 );
or ( n61661 , n61651 , n61659 , n61660 );
and ( n61662 , n61646 , n61661 );
and ( n61663 , n56071 , n55033 );
and ( n61664 , n56073 , n55030 );
nor ( n61665 , n61663 , n61664 );
xnor ( n61666 , n61665 , n53885 );
and ( n61667 , n56336 , n54693 );
and ( n61668 , n56338 , n54691 );
nor ( n61669 , n61667 , n61668 );
xnor ( n61670 , n61669 , n53892 );
and ( n61671 , n61666 , n61670 );
and ( n61672 , n56806 , n54285 );
and ( n61673 , n56495 , n54283 );
nor ( n61674 , n61672 , n61673 );
xnor ( n61675 , n61674 , n53794 );
and ( n61676 , n61670 , n61675 );
and ( n61677 , n61666 , n61675 );
or ( n61678 , n61671 , n61676 , n61677 );
and ( n61679 , n57027 , n53972 );
and ( n61680 , n56855 , n53970 );
nor ( n61681 , n61679 , n61680 );
xnor ( n61682 , n61681 , n53662 );
and ( n61683 , n57511 , n53739 );
and ( n61684 , n57244 , n53737 );
nor ( n61685 , n61683 , n61684 );
xnor ( n61686 , n61685 , n53315 );
and ( n61687 , n61682 , n61686 );
and ( n61688 , n57517 , n53455 );
and ( n61689 , n57519 , n53453 );
nor ( n61690 , n61688 , n61689 );
xnor ( n61691 , n61690 , n53159 );
and ( n61692 , n61686 , n61691 );
and ( n61693 , n61682 , n61691 );
or ( n61694 , n61687 , n61692 , n61693 );
and ( n61695 , n61678 , n61694 );
xor ( n61696 , n61614 , n61618 );
xor ( n61697 , n61696 , n61623 );
and ( n61698 , n61694 , n61697 );
and ( n61699 , n61678 , n61697 );
or ( n61700 , n61695 , n61698 , n61699 );
xor ( n61701 , n61574 , n61578 );
xor ( n61702 , n61701 , n61588 );
and ( n61703 , n61700 , n61702 );
xor ( n61704 , n61600 , n61609 );
xor ( n61705 , n61704 , n61626 );
and ( n61706 , n61702 , n61705 );
and ( n61707 , n61700 , n61705 );
or ( n61708 , n61703 , n61706 , n61707 );
and ( n61709 , n61661 , n61708 );
and ( n61710 , n61646 , n61708 );
or ( n61711 , n61662 , n61709 , n61710 );
xor ( n61712 , n61570 , n61635 );
xor ( n61713 , n61712 , n61638 );
and ( n61714 , n61711 , n61713 );
xor ( n61715 , n61591 , n61629 );
xor ( n61716 , n61715 , n61632 );
and ( n61717 , n57953 , n53293 );
and ( n61718 , n57688 , n53291 );
nor ( n61719 , n61717 , n61718 );
xnor ( n61720 , n61719 , n52963 );
and ( n61721 , n58117 , n53021 );
and ( n61722 , n57970 , n53019 );
nor ( n61723 , n61721 , n61722 );
xnor ( n61724 , n61723 , n52839 );
and ( n61725 , n61720 , n61724 );
and ( n61726 , n57244 , n53972 );
and ( n61727 , n57027 , n53970 );
nor ( n61728 , n61726 , n61727 );
xnor ( n61729 , n61728 , n53662 );
and ( n61730 , n57519 , n53739 );
and ( n61731 , n57511 , n53737 );
nor ( n61732 , n61730 , n61731 );
xnor ( n61733 , n61732 , n53315 );
and ( n61734 , n61729 , n61733 );
and ( n61735 , n61724 , n61734 );
and ( n61736 , n61720 , n61734 );
or ( n61737 , n61725 , n61735 , n61736 );
and ( n61738 , n56495 , n54693 );
and ( n61739 , n56336 , n54691 );
nor ( n61740 , n61738 , n61739 );
xnor ( n61741 , n61740 , n53892 );
and ( n61742 , n56855 , n54285 );
and ( n61743 , n56806 , n54283 );
nor ( n61744 , n61742 , n61743 );
xnor ( n61745 , n61744 , n53794 );
and ( n61746 , n61741 , n61745 );
and ( n61747 , n56338 , n55033 );
and ( n61748 , n56071 , n55030 );
nor ( n61749 , n61747 , n61748 );
xnor ( n61750 , n61749 , n53885 );
and ( n61751 , n57688 , n53455 );
and ( n61752 , n57517 , n53453 );
nor ( n61753 , n61751 , n61752 );
xnor ( n61754 , n61753 , n53159 );
and ( n61755 , n61750 , n61754 );
and ( n61756 , n57970 , n53293 );
and ( n61757 , n57953 , n53291 );
nor ( n61758 , n61756 , n61757 );
xnor ( n61759 , n61758 , n52963 );
and ( n61760 , n61754 , n61759 );
and ( n61761 , n61750 , n61759 );
or ( n61762 , n61755 , n61760 , n61761 );
and ( n61763 , n61746 , n61762 );
and ( n61764 , n58144 , n53021 );
and ( n61765 , n58117 , n53019 );
nor ( n61766 , n61764 , n61765 );
xnor ( n61767 , n61766 , n52839 );
and ( n61768 , n58571 , n52886 );
and ( n61769 , n58171 , n52884 );
nor ( n61770 , n61768 , n61769 );
xnor ( n61771 , n61770 , n52657 );
and ( n61772 , n61767 , n61771 );
and ( n61773 , n58837 , n52617 );
and ( n61774 , n58800 , n52615 );
nor ( n61775 , n61773 , n61774 );
xnor ( n61776 , n61775 , n52558 );
and ( n61777 , n61771 , n61776 );
and ( n61778 , n61767 , n61776 );
or ( n61779 , n61772 , n61777 , n61778 );
and ( n61780 , n61762 , n61779 );
and ( n61781 , n61746 , n61779 );
or ( n61782 , n61763 , n61780 , n61781 );
and ( n61783 , n61737 , n61782 );
xor ( n61784 , n61652 , n61653 );
xor ( n61785 , n61784 , n61655 );
and ( n61786 , n61782 , n61785 );
and ( n61787 , n61737 , n61785 );
or ( n61788 , n61783 , n61786 , n61787 );
xor ( n61789 , n61648 , n61650 );
xor ( n61790 , n61789 , n61658 );
and ( n61791 , n61788 , n61790 );
xor ( n61792 , n61700 , n61702 );
xor ( n61793 , n61792 , n61705 );
and ( n61794 , n61790 , n61793 );
and ( n61795 , n61788 , n61793 );
or ( n61796 , n61791 , n61794 , n61795 );
and ( n61797 , n61716 , n61796 );
xor ( n61798 , n61646 , n61661 );
xor ( n61799 , n61798 , n61708 );
and ( n61800 , n61796 , n61799 );
and ( n61801 , n61716 , n61799 );
or ( n61802 , n61797 , n61800 , n61801 );
and ( n61803 , n61713 , n61802 );
and ( n61804 , n61711 , n61802 );
or ( n61805 , n61714 , n61803 , n61804 );
and ( n61806 , n61643 , n61805 );
and ( n61807 , n61641 , n61805 );
or ( n61808 , n61644 , n61806 , n61807 );
and ( n61809 , n61567 , n61808 );
and ( n61810 , n61565 , n61808 );
or ( n61811 , n61568 , n61809 , n61810 );
and ( n61812 , n61499 , n61811 );
and ( n61813 , n61497 , n61811 );
or ( n61814 , n61500 , n61812 , n61813 );
and ( n61815 , n61422 , n61814 );
xor ( n61816 , n61260 , n61264 );
xor ( n61817 , n61816 , n61267 );
and ( n61818 , n61814 , n61817 );
and ( n61819 , n61422 , n61817 );
or ( n61820 , n61815 , n61818 , n61819 );
xor ( n61821 , n61308 , n61310 );
and ( n61822 , n61820 , n61821 );
and ( n61823 , n55406 , n54693 );
and ( n61824 , n55365 , n54691 );
nor ( n61825 , n61823 , n61824 );
xnor ( n61826 , n61825 , n53892 );
xor ( n61827 , n61248 , n61252 );
xor ( n61828 , n61827 , n61257 );
and ( n61829 , n61826 , n61828 );
xor ( n61830 , n61497 , n61499 );
xor ( n61831 , n61830 , n61811 );
xor ( n61832 , n61109 , n61113 );
xor ( n61833 , n61832 , n61116 );
and ( n61834 , n61831 , n61833 );
and ( n61835 , n55769 , n54285 );
and ( n61836 , n55720 , n54283 );
nor ( n61837 , n61835 , n61836 );
xnor ( n61838 , n61837 , n53794 );
xor ( n61839 , n61238 , n61242 );
xor ( n61840 , n61839 , n61245 );
and ( n61841 , n61838 , n61840 );
and ( n61842 , n61833 , n61841 );
and ( n61843 , n61831 , n61841 );
or ( n61844 , n61834 , n61842 , n61843 );
and ( n61845 , n61829 , n61844 );
xor ( n61846 , n61414 , n61416 );
and ( n61847 , n61844 , n61846 );
and ( n61848 , n61829 , n61846 );
or ( n61849 , n61845 , n61847 , n61848 );
and ( n61850 , n61821 , n61849 );
and ( n61851 , n61820 , n61849 );
or ( n61852 , n61822 , n61850 , n61851 );
and ( n61853 , n61420 , n61852 );
xor ( n61854 , n61301 , n61303 );
xor ( n61855 , n61854 , n61311 );
and ( n61856 , n61852 , n61855 );
and ( n61857 , n61420 , n61855 );
or ( n61858 , n61853 , n61856 , n61857 );
and ( n61859 , n61316 , n61858 );
and ( n61860 , n61314 , n61858 );
or ( n61861 , n61317 , n61859 , n61860 );
and ( n61862 , n61298 , n61861 );
and ( n61863 , n61170 , n61861 );
or ( n61864 , n61299 , n61862 , n61863 );
and ( n61865 , n61167 , n61864 );
and ( n61866 , n61041 , n61864 );
or ( n61867 , n61168 , n61865 , n61866 );
and ( n61868 , n61038 , n61867 );
and ( n61869 , n60907 , n61867 );
or ( n61870 , n61039 , n61868 , n61869 );
and ( n61871 , n60904 , n61870 );
and ( n61872 , n60673 , n61870 );
or ( n61873 , n60905 , n61871 , n61872 );
and ( n61874 , n60670 , n61873 );
and ( n61875 , n60556 , n61873 );
or ( n61876 , n60671 , n61874 , n61875 );
and ( n61877 , n60553 , n61876 );
and ( n61878 , n60551 , n61876 );
or ( n61879 , n60554 , n61877 , n61878 );
and ( n61880 , n60401 , n61879 );
and ( n61881 , n60371 , n61879 );
or ( n61882 , n60402 , n61880 , n61881 );
and ( n61883 , n60368 , n61882 );
and ( n61884 , n60102 , n61882 );
or ( n61885 , n60369 , n61883 , n61884 );
and ( n61886 , n60099 , n61885 );
and ( n61887 , n60071 , n61885 );
or ( n61888 , n60100 , n61886 , n61887 );
and ( n61889 , n60068 , n61888 );
and ( n61890 , n59964 , n61888 );
or ( n61891 , n60069 , n61889 , n61890 );
and ( n61892 , n59961 , n61891 );
and ( n61893 , n59620 , n61891 );
or ( n61894 , n59962 , n61892 , n61893 );
and ( n61895 , n59617 , n61894 );
and ( n61896 , n59473 , n61894 );
or ( n61897 , n59618 , n61895 , n61896 );
and ( n61898 , n59470 , n61897 );
and ( n61899 , n59159 , n61897 );
or ( n61900 , n59471 , n61898 , n61899 );
and ( n61901 , n59156 , n61900 );
and ( n61902 , n59118 , n61900 );
or ( n61903 , n59157 , n61901 , n61902 );
and ( n61904 , n59115 , n61903 );
and ( n61905 , n58790 , n61903 );
or ( n61906 , n59116 , n61904 , n61905 );
and ( n61907 , n58787 , n61906 );
and ( n61908 , n58737 , n61906 );
or ( n61909 , n58788 , n61907 , n61908 );
and ( n61910 , n58734 , n61909 );
and ( n61911 , n58732 , n61909 );
or ( n61912 , n58735 , n61910 , n61911 );
and ( n61913 , n58502 , n61912 );
and ( n61914 , n58412 , n61912 );
or ( n61915 , n58503 , n61913 , n61914 );
and ( n61916 , n58409 , n61915 );
and ( n61917 , n58309 , n61915 );
or ( n61918 , n58410 , n61916 , n61917 );
and ( n61919 , n58306 , n61918 );
and ( n61920 , n57931 , n61918 );
or ( n61921 , n58307 , n61919 , n61920 );
and ( n61922 , n57928 , n61921 );
and ( n61923 , n57878 , n61921 );
or ( n61924 , n57929 , n61922 , n61923 );
and ( n61925 , n57875 , n61924 );
and ( n61926 , n57678 , n61924 );
or ( n61927 , n57876 , n61925 , n61926 );
and ( n61928 , n57675 , n61927 );
and ( n61929 , n57472 , n61927 );
or ( n61930 , n57676 , n61928 , n61929 );
and ( n61931 , n57469 , n61930 );
and ( n61932 , n57234 , n61930 );
or ( n61933 , n57470 , n61931 , n61932 );
and ( n61934 , n57231 , n61933 );
and ( n61935 , n57133 , n61933 );
or ( n61936 , n57232 , n61934 , n61935 );
and ( n61937 , n57130 , n61936 );
and ( n61938 , n56953 , n61936 );
or ( n61939 , n57131 , n61937 , n61938 );
and ( n61940 , n56950 , n61939 );
and ( n61941 , n56738 , n61939 );
or ( n61942 , n56951 , n61940 , n61941 );
and ( n61943 , n56735 , n61942 );
and ( n61944 , n56697 , n61942 );
or ( n61945 , n56736 , n61943 , n61944 );
and ( n61946 , n56694 , n61945 );
and ( n61947 , n56451 , n61945 );
or ( n61948 , n56695 , n61946 , n61947 );
and ( n61949 , n56448 , n61948 );
and ( n61950 , n56312 , n61948 );
or ( n61951 , n56449 , n61949 , n61950 );
and ( n61952 , n56309 , n61951 );
and ( n61953 , n56307 , n61951 );
or ( n61954 , n56310 , n61952 , n61953 );
and ( n61955 , n56060 , n61954 );
and ( n61956 , n55938 , n61954 );
or ( n61957 , n56061 , n61955 , n61956 );
and ( n61958 , n55935 , n61957 );
and ( n61959 , n55865 , n61957 );
or ( n61960 , n55936 , n61958 , n61959 );
and ( n61961 , n55862 , n61960 );
and ( n61962 , n55565 , n61960 );
or ( n61963 , n55863 , n61961 , n61962 );
and ( n61964 , n55562 , n61963 );
and ( n61965 , n55320 , n61963 );
or ( n61966 , n55563 , n61964 , n61965 );
and ( n61967 , n55317 , n61966 );
and ( n61968 , n55299 , n61966 );
or ( n61969 , n55318 , n61967 , n61968 );
and ( n61970 , n55296 , n61969 );
and ( n61971 , n55294 , n61969 );
or ( n61972 , n55297 , n61970 , n61971 );
and ( n61973 , n54996 , n61972 );
and ( n61974 , n54859 , n61972 );
or ( n61975 , n54997 , n61973 , n61974 );
and ( n61976 , n54856 , n61975 );
and ( n61977 , n54637 , n61975 );
or ( n61978 , n54857 , n61976 , n61977 );
and ( n61979 , n54634 , n61978 );
and ( n61980 , n54586 , n61978 );
or ( n61981 , n54635 , n61979 , n61980 );
and ( n61982 , n54583 , n61981 );
and ( n61983 , n54440 , n61981 );
or ( n61984 , n54584 , n61982 , n61983 );
and ( n61985 , n54437 , n61984 );
and ( n61986 , n54435 , n61984 );
or ( n61987 , n54438 , n61985 , n61986 );
and ( n61988 , n54264 , n61987 );
and ( n61989 , n54196 , n61987 );
or ( n61990 , n54265 , n61988 , n61989 );
and ( n61991 , n54193 , n61990 );
and ( n61992 , n53884 , n61990 );
or ( n61993 , n54194 , n61991 , n61992 );
and ( n61994 , n53881 , n61993 );
and ( n61995 , n53715 , n61993 );
or ( n61996 , n53882 , n61994 , n61995 );
and ( n61997 , n53712 , n61996 );
and ( n61998 , n53563 , n61996 );
or ( n61999 , n53713 , n61997 , n61998 );
and ( n62000 , n53560 , n61999 );
and ( n62001 , n53451 , n61999 );
or ( n62002 , n53561 , n62000 , n62001 );
and ( n62003 , n53448 , n62002 );
and ( n62004 , n53396 , n62002 );
or ( n62005 , n53449 , n62003 , n62004 );
and ( n62006 , n53393 , n62005 );
and ( n62007 , n53257 , n62005 );
or ( n62008 , n53394 , n62006 , n62007 );
and ( n62009 , n53254 , n62008 );
and ( n62010 , n53089 , n62008 );
or ( n62011 , n53255 , n62009 , n62010 );
and ( n62012 , n53086 , n62011 );
and ( n62013 , n53017 , n62011 );
or ( n62014 , n53087 , n62012 , n62013 );
and ( n62015 , n53014 , n62014 );
and ( n62016 , n52882 , n62014 );
or ( n62017 , n53015 , n62015 , n62016 );
and ( n62018 , n52879 , n62017 );
and ( n62019 , n52799 , n62017 );
or ( n62020 , n52880 , n62018 , n62019 );
and ( n62021 , n52796 , n62020 );
and ( n62022 , n52708 , n62020 );
or ( n62023 , n52797 , n62021 , n62022 );
and ( n62024 , n52705 , n62023 );
and ( n62025 , n52613 , n62023 );
or ( n62026 , n52706 , n62024 , n62025 );
and ( n62027 , n52610 , n62026 );
and ( n62028 , n52493 , n62026 );
or ( n62029 , n52611 , n62027 , n62028 );
and ( n62030 , n52490 , n62029 );
and ( n62031 , n52419 , n62029 );
or ( n62032 , n52491 , n62030 , n62031 );
and ( n62033 , n52416 , n62032 );
and ( n62034 , n52414 , n62032 );
or ( n62035 , n52417 , n62033 , n62034 );
and ( n62036 , n52395 , n62035 );
and ( n62037 , n52295 , n62035 );
or ( n62038 , n52396 , n62036 , n62037 );
and ( n62039 , n52292 , n62038 );
and ( n62040 , n52244 , n62038 );
or ( n62041 , n52293 , n62039 , n62040 );
and ( n62042 , n52241 , n62041 );
and ( n62043 , n52208 , n62041 );
or ( n62044 , n52242 , n62042 , n62043 );
and ( n62045 , n52205 , n62044 );
and ( n62046 , n52147 , n62044 );
or ( n62047 , n52206 , n62045 , n62046 );
and ( n62048 , n52144 , n62047 );
and ( n62049 , n52117 , n62047 );
or ( n62050 , n52145 , n62048 , n62049 );
and ( n62051 , n52114 , n62050 );
and ( n62052 , n52112 , n62050 );
or ( n62053 , n52115 , n62051 , n62052 );
xor ( n62054 , n52082 , n62053 );
not ( n62055 , n62054 );
xor ( n62056 , n52112 , n52114 );
xor ( n62057 , n62056 , n62050 );
xor ( n62058 , n52117 , n52144 );
xor ( n62059 , n62058 , n62047 );
xor ( n62060 , n52147 , n52205 );
xor ( n62061 , n62060 , n62044 );
xor ( n62062 , n52208 , n52241 );
xor ( n62063 , n62062 , n62041 );
xor ( n62064 , n52244 , n52292 );
xor ( n62065 , n62064 , n62038 );
xor ( n62066 , n52295 , n52395 );
xor ( n62067 , n62066 , n62035 );
xor ( n62068 , n52414 , n52416 );
xor ( n62069 , n62068 , n62032 );
xor ( n62070 , n52419 , n52490 );
xor ( n62071 , n62070 , n62029 );
xor ( n62072 , n52493 , n52610 );
xor ( n62073 , n62072 , n62026 );
xor ( n62074 , n52613 , n52705 );
xor ( n62075 , n62074 , n62023 );
xor ( n62076 , n52708 , n52796 );
xor ( n62077 , n62076 , n62020 );
xor ( n62078 , n52799 , n52879 );
xor ( n62079 , n62078 , n62017 );
xor ( n62080 , n52882 , n53014 );
xor ( n62081 , n62080 , n62014 );
xor ( n62082 , n53017 , n53086 );
xor ( n62083 , n62082 , n62011 );
xor ( n62084 , n53089 , n53254 );
xor ( n62085 , n62084 , n62008 );
xor ( n62086 , n53257 , n53393 );
xor ( n62087 , n62086 , n62005 );
xor ( n62088 , n53396 , n53448 );
xor ( n62089 , n62088 , n62002 );
xor ( n62090 , n53451 , n53560 );
xor ( n62091 , n62090 , n61999 );
xor ( n62092 , n53563 , n53712 );
xor ( n62093 , n62092 , n61996 );
xor ( n62094 , n53715 , n53881 );
xor ( n62095 , n62094 , n61993 );
xor ( n62096 , n53884 , n54193 );
xor ( n62097 , n62096 , n61990 );
xor ( n62098 , n54196 , n54264 );
xor ( n62099 , n62098 , n61987 );
xor ( n62100 , n54435 , n54437 );
xor ( n62101 , n62100 , n61984 );
xor ( n62102 , n54440 , n54583 );
xor ( n62103 , n62102 , n61981 );
xor ( n62104 , n54586 , n54634 );
xor ( n62105 , n62104 , n61978 );
xor ( n62106 , n54637 , n54856 );
xor ( n62107 , n62106 , n61975 );
xor ( n62108 , n54859 , n54996 );
xor ( n62109 , n62108 , n61972 );
xor ( n62110 , n55294 , n55296 );
xor ( n62111 , n62110 , n61969 );
xor ( n62112 , n55299 , n55317 );
xor ( n62113 , n62112 , n61966 );
xor ( n62114 , n55320 , n55562 );
xor ( n62115 , n62114 , n61963 );
xor ( n62116 , n55565 , n55862 );
xor ( n62117 , n62116 , n61960 );
xor ( n62118 , n55865 , n55935 );
xor ( n62119 , n62118 , n61957 );
xor ( n62120 , n55938 , n56060 );
xor ( n62121 , n62120 , n61954 );
xor ( n62122 , n56307 , n56309 );
xor ( n62123 , n62122 , n61951 );
xor ( n62124 , n56312 , n56448 );
xor ( n62125 , n62124 , n61948 );
xor ( n62126 , n56451 , n56694 );
xor ( n62127 , n62126 , n61945 );
xor ( n62128 , n56697 , n56735 );
xor ( n62129 , n62128 , n61942 );
xor ( n62130 , n56738 , n56950 );
xor ( n62131 , n62130 , n61939 );
xor ( n62132 , n56953 , n57130 );
xor ( n62133 , n62132 , n61936 );
xor ( n62134 , n57133 , n57231 );
xor ( n62135 , n62134 , n61933 );
xor ( n62136 , n57234 , n57469 );
xor ( n62137 , n62136 , n61930 );
xor ( n62138 , n57472 , n57675 );
xor ( n62139 , n62138 , n61927 );
xor ( n62140 , n57678 , n57875 );
xor ( n62141 , n62140 , n61924 );
xor ( n62142 , n57878 , n57928 );
xor ( n62143 , n62142 , n61921 );
xor ( n62144 , n57931 , n58306 );
xor ( n62145 , n62144 , n61918 );
xor ( n62146 , n58309 , n58409 );
xor ( n62147 , n62146 , n61915 );
xor ( n62148 , n58412 , n58502 );
xor ( n62149 , n62148 , n61912 );
xor ( n62150 , n58732 , n58734 );
xor ( n62151 , n62150 , n61909 );
xor ( n62152 , n58737 , n58787 );
xor ( n62153 , n62152 , n61906 );
xor ( n62154 , n58790 , n59115 );
xor ( n62155 , n62154 , n61903 );
xor ( n62156 , n59118 , n59156 );
xor ( n62157 , n62156 , n61900 );
xor ( n62158 , n59159 , n59470 );
xor ( n62159 , n62158 , n61897 );
xor ( n62160 , n59473 , n59617 );
xor ( n62161 , n62160 , n61894 );
xor ( n62162 , n59620 , n59961 );
xor ( n62163 , n62162 , n61891 );
xor ( n62164 , n59964 , n60068 );
xor ( n62165 , n62164 , n61888 );
xor ( n62166 , n60071 , n60099 );
xor ( n62167 , n62166 , n61885 );
xor ( n62168 , n60102 , n60368 );
xor ( n62169 , n62168 , n61882 );
xor ( n62170 , n60371 , n60401 );
xor ( n62171 , n62170 , n61879 );
xor ( n62172 , n60551 , n60553 );
xor ( n62173 , n62172 , n61876 );
xor ( n62174 , n60556 , n60670 );
xor ( n62175 , n62174 , n61873 );
xor ( n62176 , n60673 , n60904 );
xor ( n62177 , n62176 , n61870 );
xor ( n62178 , n60907 , n61038 );
xor ( n62179 , n62178 , n61867 );
xor ( n62180 , n61041 , n61167 );
xor ( n62181 , n62180 , n61864 );
xor ( n62182 , n61170 , n61298 );
xor ( n62183 , n62182 , n61861 );
xor ( n62184 , n61314 , n61316 );
xor ( n62185 , n62184 , n61858 );
xor ( n62186 , n61407 , n61409 );
xor ( n62187 , n62186 , n61417 );
xor ( n62188 , n61826 , n61828 );
xor ( n62189 , n61565 , n61567 );
xor ( n62190 , n62189 , n61808 );
nor ( n62191 , n52346 , n52344 );
xnor ( n62192 , n62191 , n52300 );
nor ( n62193 , n52318 , n52316 );
xnor ( n62194 , n62193 , n52213 );
and ( n62195 , n62192 , n62194 );
xor ( n62196 , n62192 , n62194 );
nor ( n62197 , n52540 , n52538 );
xnor ( n62198 , n62197 , n52424 );
nor ( n62199 , n52346 , n52344 );
xnor ( n62200 , n62199 , n52300 );
and ( n62201 , n62198 , n62200 );
nor ( n62202 , n52318 , n52316 );
xnor ( n62203 , n62202 , n52213 );
and ( n62204 , n62200 , n62203 );
and ( n62205 , n62198 , n62203 );
or ( n62206 , n62201 , n62204 , n62205 );
and ( n62207 , n62196 , n62206 );
xor ( n62208 , n61174 , n61176 );
xor ( n62209 , n62208 , n52119 );
and ( n62210 , n62206 , n62209 );
and ( n62211 , n62196 , n62209 );
or ( n62212 , n62207 , n62210 , n62211 );
and ( n62213 , n62195 , n62212 );
xor ( n62214 , n61043 , n61045 );
xor ( n62215 , n62214 , n61048 );
and ( n62216 , n62212 , n62215 );
and ( n62217 , n62195 , n62215 );
or ( n62218 , n62213 , n62216 , n62217 );
and ( n62219 , n58571 , n52617 );
and ( n62220 , n58171 , n52615 );
nor ( n62221 , n62219 , n62220 );
xnor ( n62222 , n62221 , n52558 );
and ( n62223 , n62218 , n62222 );
xor ( n62224 , n61188 , n61192 );
xor ( n62225 , n62224 , n61195 );
and ( n62226 , n62222 , n62225 );
and ( n62227 , n62218 , n62225 );
or ( n62228 , n62223 , n62226 , n62227 );
and ( n62229 , n58117 , n52886 );
and ( n62230 , n57970 , n52884 );
nor ( n62231 , n62229 , n62230 );
xnor ( n62232 , n62231 , n52657 );
and ( n62233 , n62228 , n62232 );
xor ( n62234 , n61198 , n61202 );
xor ( n62235 , n62234 , n61205 );
and ( n62236 , n62232 , n62235 );
and ( n62237 , n62228 , n62235 );
or ( n62238 , n62233 , n62236 , n62237 );
and ( n62239 , n57688 , n53021 );
and ( n62240 , n57517 , n53019 );
nor ( n62241 , n62239 , n62240 );
xnor ( n62242 , n62241 , n52839 );
and ( n62243 , n62238 , n62242 );
xor ( n62244 , n61208 , n61212 );
xor ( n62245 , n62244 , n61215 );
and ( n62246 , n62242 , n62245 );
and ( n62247 , n62238 , n62245 );
or ( n62248 , n62243 , n62246 , n62247 );
and ( n62249 , n57511 , n53293 );
and ( n62250 , n57244 , n53291 );
nor ( n62251 , n62249 , n62250 );
xnor ( n62252 , n62251 , n52963 );
and ( n62253 , n62248 , n62252 );
xor ( n62254 , n61218 , n61222 );
xor ( n62255 , n62254 , n61225 );
and ( n62256 , n62252 , n62255 );
and ( n62257 , n62248 , n62255 );
or ( n62258 , n62253 , n62256 , n62257 );
xor ( n62259 , n61228 , n61232 );
xor ( n62260 , n62259 , n61235 );
and ( n62261 , n62258 , n62260 );
and ( n62262 , n62190 , n62261 );
xor ( n62263 , n61838 , n61840 );
and ( n62264 , n62261 , n62263 );
and ( n62265 , n62190 , n62263 );
or ( n62266 , n62262 , n62264 , n62265 );
and ( n62267 , n62188 , n62266 );
xor ( n62268 , n61831 , n61833 );
xor ( n62269 , n62268 , n61841 );
and ( n62270 , n62266 , n62269 );
and ( n62271 , n62188 , n62269 );
or ( n62272 , n62267 , n62270 , n62271 );
xor ( n62273 , n61422 , n61814 );
xor ( n62274 , n62273 , n61817 );
and ( n62275 , n62272 , n62274 );
xor ( n62276 , n61829 , n61844 );
xor ( n62277 , n62276 , n61846 );
and ( n62278 , n62274 , n62277 );
and ( n62279 , n62272 , n62277 );
or ( n62280 , n62275 , n62278 , n62279 );
and ( n62281 , n62187 , n62280 );
xor ( n62282 , n61820 , n61821 );
xor ( n62283 , n62282 , n61849 );
and ( n62284 , n62280 , n62283 );
and ( n62285 , n62187 , n62283 );
or ( n62286 , n62281 , n62284 , n62285 );
xor ( n62287 , n61420 , n61852 );
xor ( n62288 , n62287 , n61855 );
and ( n62289 , n62286 , n62288 );
xor ( n62290 , n62286 , n62288 );
xor ( n62291 , n62187 , n62280 );
xor ( n62292 , n62291 , n62283 );
xor ( n62293 , n62272 , n62274 );
xor ( n62294 , n62293 , n62277 );
xor ( n62295 , n62188 , n62266 );
xor ( n62296 , n62295 , n62269 );
xor ( n62297 , n61641 , n61643 );
xor ( n62298 , n62297 , n61805 );
xor ( n62299 , n61711 , n61713 );
xor ( n62300 , n62299 , n61802 );
xor ( n62301 , n61716 , n61796 );
xor ( n62302 , n62301 , n61799 );
xor ( n62303 , n61678 , n61694 );
xor ( n62304 , n62303 , n61697 );
and ( n62305 , n58800 , n52617 );
and ( n62306 , n58571 , n52615 );
nor ( n62307 , n62305 , n62306 );
xnor ( n62308 , n62307 , n52558 );
xor ( n62309 , n61171 , n61180 );
xor ( n62310 , n62309 , n61185 );
and ( n62311 , n62308 , n62310 );
and ( n62312 , n62304 , n62311 );
xor ( n62313 , n61666 , n61670 );
xor ( n62314 , n62313 , n61675 );
xor ( n62315 , n61682 , n61686 );
xor ( n62316 , n62315 , n61691 );
and ( n62317 , n62314 , n62316 );
xor ( n62318 , n61729 , n61733 );
xor ( n62319 , n61741 , n61745 );
and ( n62320 , n62318 , n62319 );
and ( n62321 , n56336 , n55033 );
and ( n62322 , n56338 , n55030 );
nor ( n62323 , n62321 , n62322 );
xnor ( n62324 , n62323 , n53885 );
and ( n62325 , n56806 , n54693 );
and ( n62326 , n56495 , n54691 );
nor ( n62327 , n62325 , n62326 );
xnor ( n62328 , n62327 , n53892 );
and ( n62329 , n62324 , n62328 );
and ( n62330 , n57027 , n54285 );
and ( n62331 , n56855 , n54283 );
nor ( n62332 , n62330 , n62331 );
xnor ( n62333 , n62332 , n53794 );
and ( n62334 , n62328 , n62333 );
and ( n62335 , n62324 , n62333 );
or ( n62336 , n62329 , n62334 , n62335 );
and ( n62337 , n62319 , n62336 );
and ( n62338 , n62318 , n62336 );
or ( n62339 , n62320 , n62337 , n62338 );
and ( n62340 , n62316 , n62339 );
and ( n62341 , n62314 , n62339 );
or ( n62342 , n62317 , n62340 , n62341 );
and ( n62343 , n62311 , n62342 );
and ( n62344 , n62304 , n62342 );
or ( n62345 , n62312 , n62343 , n62344 );
xor ( n62346 , n61788 , n61790 );
xor ( n62347 , n62346 , n61793 );
and ( n62348 , n62345 , n62347 );
and ( n62349 , n57511 , n53972 );
and ( n62350 , n57244 , n53970 );
nor ( n62351 , n62349 , n62350 );
xnor ( n62352 , n62351 , n53662 );
and ( n62353 , n57517 , n53739 );
and ( n62354 , n57519 , n53737 );
nor ( n62355 , n62353 , n62354 );
xnor ( n62356 , n62355 , n53315 );
and ( n62357 , n62352 , n62356 );
and ( n62358 , n57953 , n53455 );
and ( n62359 , n57688 , n53453 );
nor ( n62360 , n62358 , n62359 );
xnor ( n62361 , n62360 , n53159 );
and ( n62362 , n62356 , n62361 );
and ( n62363 , n62352 , n62361 );
or ( n62364 , n62357 , n62362 , n62363 );
and ( n62365 , n58117 , n53293 );
and ( n62366 , n57970 , n53291 );
nor ( n62367 , n62365 , n62366 );
xnor ( n62368 , n62367 , n52963 );
and ( n62369 , n58171 , n53021 );
and ( n62370 , n58144 , n53019 );
nor ( n62371 , n62369 , n62370 );
xnor ( n62372 , n62371 , n52839 );
and ( n62373 , n62368 , n62372 );
and ( n62374 , n58800 , n52886 );
and ( n62375 , n58571 , n52884 );
nor ( n62376 , n62374 , n62375 );
xnor ( n62377 , n62376 , n52657 );
and ( n62378 , n62372 , n62377 );
and ( n62379 , n62368 , n62377 );
or ( n62380 , n62373 , n62378 , n62379 );
and ( n62381 , n62364 , n62380 );
and ( n62382 , n58864 , n52617 );
and ( n62383 , n58837 , n52615 );
nor ( n62384 , n62382 , n62383 );
xnor ( n62385 , n62384 , n52558 );
nor ( n62386 , n52170 , n52168 );
xnor ( n62387 , n62386 , n52152 );
and ( n62388 , n62385 , n62387 );
and ( n62389 , n52169 , n52152 );
and ( n62390 , n62387 , n62389 );
and ( n62391 , n62385 , n62389 );
or ( n62392 , n62388 , n62390 , n62391 );
and ( n62393 , n62380 , n62392 );
and ( n62394 , n62364 , n62392 );
or ( n62395 , n62381 , n62393 , n62394 );
xor ( n62396 , n61720 , n61724 );
xor ( n62397 , n62396 , n61734 );
and ( n62398 , n62395 , n62397 );
xor ( n62399 , n61746 , n61762 );
xor ( n62400 , n62399 , n61779 );
and ( n62401 , n62397 , n62400 );
and ( n62402 , n62395 , n62400 );
or ( n62403 , n62398 , n62401 , n62402 );
xor ( n62404 , n61737 , n61782 );
xor ( n62405 , n62404 , n61785 );
and ( n62406 , n62403 , n62405 );
and ( n62407 , n58171 , n52886 );
and ( n62408 , n58144 , n52884 );
nor ( n62409 , n62407 , n62408 );
xnor ( n62410 , n62409 , n52657 );
xor ( n62411 , n62195 , n62212 );
xor ( n62412 , n62411 , n62215 );
and ( n62413 , n62410 , n62412 );
and ( n62414 , n62405 , n62413 );
and ( n62415 , n62403 , n62413 );
or ( n62416 , n62406 , n62414 , n62415 );
and ( n62417 , n62347 , n62416 );
and ( n62418 , n62345 , n62416 );
or ( n62419 , n62348 , n62417 , n62418 );
and ( n62420 , n62302 , n62419 );
xor ( n62421 , n62228 , n62232 );
xor ( n62422 , n62421 , n62235 );
xor ( n62423 , n62308 , n62310 );
xor ( n62424 , n61750 , n61754 );
xor ( n62425 , n62424 , n61759 );
xor ( n62426 , n61767 , n61771 );
xor ( n62427 , n62426 , n61776 );
and ( n62428 , n62425 , n62427 );
xor ( n62429 , n62196 , n62206 );
xor ( n62430 , n62429 , n62209 );
and ( n62431 , n62427 , n62430 );
and ( n62432 , n62425 , n62430 );
or ( n62433 , n62428 , n62431 , n62432 );
and ( n62434 , n62423 , n62433 );
xor ( n62435 , n62198 , n62200 );
xor ( n62436 , n62435 , n62203 );
nor ( n62437 , n52540 , n52538 );
xnor ( n62438 , n62437 , n52424 );
nor ( n62439 , n52346 , n52344 );
xnor ( n62440 , n62439 , n52300 );
and ( n62441 , n62438 , n62440 );
and ( n62442 , n62440 , n52168 );
and ( n62443 , n62438 , n52168 );
or ( n62444 , n62441 , n62442 , n62443 );
and ( n62445 , n62436 , n62444 );
and ( n62446 , n58864 , n52615 );
nor ( n62447 , n52617 , n62446 );
xnor ( n62448 , n62447 , n52558 );
nor ( n62449 , n52318 , n52316 );
xnor ( n62450 , n62449 , n52213 );
and ( n62451 , n62448 , n62450 );
and ( n62452 , n62444 , n62451 );
and ( n62453 , n62436 , n62451 );
or ( n62454 , n62445 , n62452 , n62453 );
and ( n62455 , n56495 , n55033 );
and ( n62456 , n56336 , n55030 );
nor ( n62457 , n62455 , n62456 );
xnor ( n62458 , n62457 , n53885 );
and ( n62459 , n56855 , n54693 );
and ( n62460 , n56806 , n54691 );
nor ( n62461 , n62459 , n62460 );
xnor ( n62462 , n62461 , n53892 );
and ( n62463 , n62458 , n62462 );
and ( n62464 , n57244 , n54285 );
and ( n62465 , n57027 , n54283 );
nor ( n62466 , n62464 , n62465 );
xnor ( n62467 , n62466 , n53794 );
and ( n62468 , n62462 , n62467 );
and ( n62469 , n62458 , n62467 );
or ( n62470 , n62463 , n62468 , n62469 );
and ( n62471 , n57519 , n53972 );
and ( n62472 , n57511 , n53970 );
nor ( n62473 , n62471 , n62472 );
xnor ( n62474 , n62473 , n53662 );
and ( n62475 , n57688 , n53739 );
and ( n62476 , n57517 , n53737 );
nor ( n62477 , n62475 , n62476 );
xnor ( n62478 , n62477 , n53315 );
and ( n62479 , n62474 , n62478 );
and ( n62480 , n57970 , n53455 );
and ( n62481 , n57953 , n53453 );
nor ( n62482 , n62480 , n62481 );
xnor ( n62483 , n62482 , n53159 );
and ( n62484 , n62478 , n62483 );
and ( n62485 , n62474 , n62483 );
or ( n62486 , n62479 , n62484 , n62485 );
and ( n62487 , n62470 , n62486 );
and ( n62488 , n58144 , n53293 );
and ( n62489 , n58117 , n53291 );
nor ( n62490 , n62488 , n62489 );
xnor ( n62491 , n62490 , n52963 );
and ( n62492 , n58571 , n53021 );
and ( n62493 , n58171 , n53019 );
nor ( n62494 , n62492 , n62493 );
xnor ( n62495 , n62494 , n52839 );
and ( n62496 , n62491 , n62495 );
and ( n62497 , n58837 , n52886 );
and ( n62498 , n58800 , n52884 );
nor ( n62499 , n62497 , n62498 );
xnor ( n62500 , n62499 , n52657 );
and ( n62501 , n62495 , n62500 );
and ( n62502 , n62491 , n62500 );
or ( n62503 , n62496 , n62501 , n62502 );
and ( n62504 , n62486 , n62503 );
and ( n62505 , n62470 , n62503 );
or ( n62506 , n62487 , n62504 , n62505 );
and ( n62507 , n62454 , n62506 );
xor ( n62508 , n62324 , n62328 );
xor ( n62509 , n62508 , n62333 );
xor ( n62510 , n62352 , n62356 );
xor ( n62511 , n62510 , n62361 );
and ( n62512 , n62509 , n62511 );
xor ( n62513 , n62368 , n62372 );
xor ( n62514 , n62513 , n62377 );
and ( n62515 , n62511 , n62514 );
and ( n62516 , n62509 , n62514 );
or ( n62517 , n62512 , n62515 , n62516 );
and ( n62518 , n62506 , n62517 );
and ( n62519 , n62454 , n62517 );
or ( n62520 , n62507 , n62518 , n62519 );
and ( n62521 , n62433 , n62520 );
and ( n62522 , n62423 , n62520 );
or ( n62523 , n62434 , n62521 , n62522 );
xor ( n62524 , n62304 , n62311 );
xor ( n62525 , n62524 , n62342 );
and ( n62526 , n62523 , n62525 );
xor ( n62527 , n62218 , n62222 );
xor ( n62528 , n62527 , n62225 );
and ( n62529 , n62525 , n62528 );
and ( n62530 , n62523 , n62528 );
or ( n62531 , n62526 , n62529 , n62530 );
and ( n62532 , n62422 , n62531 );
xor ( n62533 , n62314 , n62316 );
xor ( n62534 , n62533 , n62339 );
xor ( n62535 , n62395 , n62397 );
xor ( n62536 , n62535 , n62400 );
and ( n62537 , n62534 , n62536 );
xor ( n62538 , n62410 , n62412 );
and ( n62539 , n62536 , n62538 );
and ( n62540 , n62534 , n62538 );
or ( n62541 , n62537 , n62539 , n62540 );
xor ( n62542 , n62318 , n62319 );
xor ( n62543 , n62542 , n62336 );
xor ( n62544 , n62364 , n62380 );
xor ( n62545 , n62544 , n62392 );
and ( n62546 , n62543 , n62545 );
xor ( n62547 , n62385 , n62387 );
xor ( n62548 , n62547 , n62389 );
xor ( n62549 , n62438 , n62440 );
xor ( n62550 , n62549 , n52168 );
xor ( n62551 , n62448 , n62450 );
and ( n62552 , n62550 , n62551 );
nor ( n62553 , n52617 , n52615 );
xnor ( n62554 , n62553 , n52558 );
nor ( n62555 , n52540 , n52538 );
xnor ( n62556 , n62555 , n52424 );
and ( n62557 , n62554 , n62556 );
nor ( n62558 , n52346 , n52344 );
xnor ( n62559 , n62558 , n52300 );
and ( n62560 , n62556 , n62559 );
and ( n62561 , n62554 , n62559 );
or ( n62562 , n62557 , n62560 , n62561 );
and ( n62563 , n62551 , n62562 );
and ( n62564 , n62550 , n62562 );
or ( n62565 , n62552 , n62563 , n62564 );
and ( n62566 , n62548 , n62565 );
and ( n62567 , n56806 , n55033 );
and ( n62568 , n56495 , n55030 );
nor ( n62569 , n62567 , n62568 );
xnor ( n62570 , n62569 , n53885 );
and ( n62571 , n57027 , n54693 );
and ( n62572 , n56855 , n54691 );
nor ( n62573 , n62571 , n62572 );
xnor ( n62574 , n62573 , n53892 );
and ( n62575 , n62570 , n62574 );
and ( n62576 , n57511 , n54285 );
and ( n62577 , n57244 , n54283 );
nor ( n62578 , n62576 , n62577 );
xnor ( n62579 , n62578 , n53794 );
and ( n62580 , n62574 , n62579 );
and ( n62581 , n62570 , n62579 );
or ( n62582 , n62575 , n62580 , n62581 );
and ( n62583 , n57517 , n53972 );
and ( n62584 , n57519 , n53970 );
nor ( n62585 , n62583 , n62584 );
xnor ( n62586 , n62585 , n53662 );
and ( n62587 , n57953 , n53739 );
and ( n62588 , n57688 , n53737 );
nor ( n62589 , n62587 , n62588 );
xnor ( n62590 , n62589 , n53315 );
and ( n62591 , n62586 , n62590 );
and ( n62592 , n58117 , n53455 );
and ( n62593 , n57970 , n53453 );
nor ( n62594 , n62592 , n62593 );
xnor ( n62595 , n62594 , n53159 );
and ( n62596 , n62590 , n62595 );
and ( n62597 , n62586 , n62595 );
or ( n62598 , n62591 , n62596 , n62597 );
and ( n62599 , n62582 , n62598 );
and ( n62600 , n58171 , n53293 );
and ( n62601 , n58144 , n53291 );
nor ( n62602 , n62600 , n62601 );
xnor ( n62603 , n62602 , n52963 );
and ( n62604 , n58800 , n53021 );
and ( n62605 , n58571 , n53019 );
nor ( n62606 , n62604 , n62605 );
xnor ( n62607 , n62606 , n52839 );
and ( n62608 , n62603 , n62607 );
and ( n62609 , n58864 , n52886 );
and ( n62610 , n58837 , n52884 );
nor ( n62611 , n62609 , n62610 );
xnor ( n62612 , n62611 , n52657 );
and ( n62613 , n62607 , n62612 );
and ( n62614 , n62603 , n62612 );
or ( n62615 , n62608 , n62613 , n62614 );
and ( n62616 , n62598 , n62615 );
and ( n62617 , n62582 , n62615 );
or ( n62618 , n62599 , n62616 , n62617 );
and ( n62619 , n62565 , n62618 );
and ( n62620 , n62548 , n62618 );
or ( n62621 , n62566 , n62619 , n62620 );
and ( n62622 , n62545 , n62621 );
and ( n62623 , n62543 , n62621 );
or ( n62624 , n62546 , n62622 , n62623 );
xor ( n62625 , n62458 , n62462 );
xor ( n62626 , n62625 , n62467 );
xor ( n62627 , n62474 , n62478 );
xor ( n62628 , n62627 , n62483 );
and ( n62629 , n62626 , n62628 );
xor ( n62630 , n62491 , n62495 );
xor ( n62631 , n62630 , n62500 );
and ( n62632 , n62628 , n62631 );
and ( n62633 , n62626 , n62631 );
or ( n62634 , n62629 , n62632 , n62633 );
xor ( n62635 , n62436 , n62444 );
xor ( n62636 , n62635 , n62451 );
and ( n62637 , n62634 , n62636 );
xor ( n62638 , n62470 , n62486 );
xor ( n62639 , n62638 , n62503 );
and ( n62640 , n62636 , n62639 );
and ( n62641 , n62634 , n62639 );
or ( n62642 , n62637 , n62640 , n62641 );
xor ( n62643 , n62425 , n62427 );
xor ( n62644 , n62643 , n62430 );
and ( n62645 , n62642 , n62644 );
xor ( n62646 , n62454 , n62506 );
xor ( n62647 , n62646 , n62517 );
and ( n62648 , n62644 , n62647 );
and ( n62649 , n62642 , n62647 );
or ( n62650 , n62645 , n62648 , n62649 );
and ( n62651 , n62624 , n62650 );
xor ( n62652 , n62423 , n62433 );
xor ( n62653 , n62652 , n62520 );
and ( n62654 , n62650 , n62653 );
and ( n62655 , n62624 , n62653 );
or ( n62656 , n62651 , n62654 , n62655 );
and ( n62657 , n62541 , n62656 );
xor ( n62658 , n62403 , n62405 );
xor ( n62659 , n62658 , n62413 );
and ( n62660 , n62656 , n62659 );
and ( n62661 , n62541 , n62659 );
or ( n62662 , n62657 , n62660 , n62661 );
and ( n62663 , n62531 , n62662 );
and ( n62664 , n62422 , n62662 );
or ( n62665 , n62532 , n62663 , n62664 );
and ( n62666 , n62419 , n62665 );
and ( n62667 , n62302 , n62665 );
or ( n62668 , n62420 , n62666 , n62667 );
and ( n62669 , n62300 , n62668 );
xor ( n62670 , n62248 , n62252 );
xor ( n62671 , n62670 , n62255 );
and ( n62672 , n62668 , n62671 );
and ( n62673 , n62300 , n62671 );
or ( n62674 , n62669 , n62672 , n62673 );
and ( n62675 , n62298 , n62674 );
xor ( n62676 , n62258 , n62260 );
and ( n62677 , n62674 , n62676 );
and ( n62678 , n62298 , n62676 );
or ( n62679 , n62675 , n62677 , n62678 );
xor ( n62680 , n62190 , n62261 );
xor ( n62681 , n62680 , n62263 );
and ( n62682 , n62679 , n62681 );
xor ( n62683 , n62679 , n62681 );
xor ( n62684 , n62298 , n62674 );
xor ( n62685 , n62684 , n62676 );
xor ( n62686 , n62238 , n62242 );
xor ( n62687 , n62686 , n62245 );
xor ( n62688 , n62345 , n62347 );
xor ( n62689 , n62688 , n62416 );
xor ( n62690 , n62509 , n62511 );
xor ( n62691 , n62690 , n62514 );
nor ( n62692 , n52318 , n52316 );
xnor ( n62693 , n62692 , n52213 );
and ( n62694 , n52317 , n52213 );
and ( n62695 , n62693 , n62694 );
xor ( n62696 , n62554 , n62556 );
xor ( n62697 , n62696 , n62559 );
and ( n62698 , n62694 , n62697 );
and ( n62699 , n62693 , n62697 );
or ( n62700 , n62695 , n62698 , n62699 );
nor ( n62701 , n52617 , n52615 );
xnor ( n62702 , n62701 , n52558 );
nor ( n62703 , n52540 , n52538 );
xnor ( n62704 , n62703 , n52424 );
and ( n62705 , n62702 , n62704 );
nor ( n62706 , n52346 , n52344 );
xnor ( n62707 , n62706 , n52300 );
and ( n62708 , n62704 , n62707 );
and ( n62709 , n62702 , n62707 );
or ( n62710 , n62705 , n62708 , n62709 );
and ( n62711 , n58864 , n52884 );
nor ( n62712 , n52886 , n62711 );
xnor ( n62713 , n62712 , n52657 );
and ( n62714 , n62713 , n52316 );
and ( n62715 , n62710 , n62714 );
and ( n62716 , n56855 , n55033 );
and ( n62717 , n56806 , n55030 );
nor ( n62718 , n62716 , n62717 );
xnor ( n62719 , n62718 , n53885 );
and ( n62720 , n57244 , n54693 );
and ( n62721 , n57027 , n54691 );
nor ( n62722 , n62720 , n62721 );
xnor ( n62723 , n62722 , n53892 );
and ( n62724 , n62719 , n62723 );
and ( n62725 , n57519 , n54285 );
and ( n62726 , n57511 , n54283 );
nor ( n62727 , n62725 , n62726 );
xnor ( n62728 , n62727 , n53794 );
and ( n62729 , n62723 , n62728 );
and ( n62730 , n62719 , n62728 );
or ( n62731 , n62724 , n62729 , n62730 );
and ( n62732 , n62714 , n62731 );
and ( n62733 , n62710 , n62731 );
or ( n62734 , n62715 , n62732 , n62733 );
and ( n62735 , n62700 , n62734 );
and ( n62736 , n57688 , n53972 );
and ( n62737 , n57517 , n53970 );
nor ( n62738 , n62736 , n62737 );
xnor ( n62739 , n62738 , n53662 );
and ( n62740 , n57970 , n53739 );
and ( n62741 , n57953 , n53737 );
nor ( n62742 , n62740 , n62741 );
xnor ( n62743 , n62742 , n53315 );
and ( n62744 , n62739 , n62743 );
and ( n62745 , n58144 , n53455 );
and ( n62746 , n58117 , n53453 );
nor ( n62747 , n62745 , n62746 );
xnor ( n62748 , n62747 , n53159 );
and ( n62749 , n62743 , n62748 );
and ( n62750 , n62739 , n62748 );
or ( n62751 , n62744 , n62749 , n62750 );
xor ( n62752 , n62570 , n62574 );
xor ( n62753 , n62752 , n62579 );
and ( n62754 , n62751 , n62753 );
xor ( n62755 , n62586 , n62590 );
xor ( n62756 , n62755 , n62595 );
and ( n62757 , n62753 , n62756 );
and ( n62758 , n62751 , n62756 );
or ( n62759 , n62754 , n62757 , n62758 );
and ( n62760 , n62734 , n62759 );
and ( n62761 , n62700 , n62759 );
or ( n62762 , n62735 , n62760 , n62761 );
and ( n62763 , n62691 , n62762 );
xor ( n62764 , n62550 , n62551 );
xor ( n62765 , n62764 , n62562 );
xor ( n62766 , n62582 , n62598 );
xor ( n62767 , n62766 , n62615 );
and ( n62768 , n62765 , n62767 );
xor ( n62769 , n62626 , n62628 );
xor ( n62770 , n62769 , n62631 );
and ( n62771 , n62767 , n62770 );
and ( n62772 , n62765 , n62770 );
or ( n62773 , n62768 , n62771 , n62772 );
and ( n62774 , n62762 , n62773 );
and ( n62775 , n62691 , n62773 );
or ( n62776 , n62763 , n62774 , n62775 );
xor ( n62777 , n62543 , n62545 );
xor ( n62778 , n62777 , n62621 );
and ( n62779 , n62776 , n62778 );
xor ( n62780 , n62642 , n62644 );
xor ( n62781 , n62780 , n62647 );
and ( n62782 , n62778 , n62781 );
and ( n62783 , n62776 , n62781 );
or ( n62784 , n62779 , n62782 , n62783 );
xor ( n62785 , n62534 , n62536 );
xor ( n62786 , n62785 , n62538 );
and ( n62787 , n62784 , n62786 );
xor ( n62788 , n62624 , n62650 );
xor ( n62789 , n62788 , n62653 );
and ( n62790 , n62786 , n62789 );
and ( n62791 , n62784 , n62789 );
or ( n62792 , n62787 , n62790 , n62791 );
xor ( n62793 , n62523 , n62525 );
xor ( n62794 , n62793 , n62528 );
and ( n62795 , n62792 , n62794 );
xor ( n62796 , n62541 , n62656 );
xor ( n62797 , n62796 , n62659 );
and ( n62798 , n62794 , n62797 );
and ( n62799 , n62792 , n62797 );
or ( n62800 , n62795 , n62798 , n62799 );
and ( n62801 , n62689 , n62800 );
xor ( n62802 , n62422 , n62531 );
xor ( n62803 , n62802 , n62662 );
and ( n62804 , n62800 , n62803 );
and ( n62805 , n62689 , n62803 );
or ( n62806 , n62801 , n62804 , n62805 );
and ( n62807 , n62687 , n62806 );
xor ( n62808 , n62302 , n62419 );
xor ( n62809 , n62808 , n62665 );
and ( n62810 , n62806 , n62809 );
and ( n62811 , n62687 , n62809 );
or ( n62812 , n62807 , n62810 , n62811 );
xor ( n62813 , n62300 , n62668 );
xor ( n62814 , n62813 , n62671 );
and ( n62815 , n62812 , n62814 );
xor ( n62816 , n62812 , n62814 );
xor ( n62817 , n62687 , n62806 );
xor ( n62818 , n62817 , n62809 );
xor ( n62819 , n62689 , n62800 );
xor ( n62820 , n62819 , n62803 );
xor ( n62821 , n62792 , n62794 );
xor ( n62822 , n62821 , n62797 );
xor ( n62823 , n62784 , n62786 );
xor ( n62824 , n62823 , n62789 );
xor ( n62825 , n62548 , n62565 );
xor ( n62826 , n62825 , n62618 );
xor ( n62827 , n62634 , n62636 );
xor ( n62828 , n62827 , n62639 );
and ( n62829 , n62826 , n62828 );
xor ( n62830 , n62603 , n62607 );
xor ( n62831 , n62830 , n62612 );
and ( n62832 , n58571 , n53293 );
and ( n62833 , n58171 , n53291 );
nor ( n62834 , n62832 , n62833 );
xnor ( n62835 , n62834 , n52963 );
and ( n62836 , n58837 , n53021 );
and ( n62837 , n58800 , n53019 );
nor ( n62838 , n62836 , n62837 );
xnor ( n62839 , n62838 , n52839 );
and ( n62840 , n62835 , n62839 );
xor ( n62841 , n62702 , n62704 );
xor ( n62842 , n62841 , n62707 );
and ( n62843 , n62839 , n62842 );
and ( n62844 , n62835 , n62842 );
or ( n62845 , n62840 , n62843 , n62844 );
and ( n62846 , n62831 , n62845 );
xor ( n62847 , n62713 , n52316 );
nor ( n62848 , n52886 , n52884 );
xnor ( n62849 , n62848 , n52657 );
nor ( n62850 , n52617 , n52615 );
xnor ( n62851 , n62850 , n52558 );
and ( n62852 , n62849 , n62851 );
nor ( n62853 , n52540 , n52538 );
xnor ( n62854 , n62853 , n52424 );
and ( n62855 , n62851 , n62854 );
and ( n62856 , n62849 , n62854 );
or ( n62857 , n62852 , n62855 , n62856 );
and ( n62858 , n62847 , n62857 );
and ( n62859 , n57027 , n55033 );
and ( n62860 , n56855 , n55030 );
nor ( n62861 , n62859 , n62860 );
xnor ( n62862 , n62861 , n53885 );
and ( n62863 , n57511 , n54693 );
and ( n62864 , n57244 , n54691 );
nor ( n62865 , n62863 , n62864 );
xnor ( n62866 , n62865 , n53892 );
and ( n62867 , n62862 , n62866 );
and ( n62868 , n57517 , n54285 );
and ( n62869 , n57519 , n54283 );
nor ( n62870 , n62868 , n62869 );
xnor ( n62871 , n62870 , n53794 );
and ( n62872 , n62866 , n62871 );
and ( n62873 , n62862 , n62871 );
or ( n62874 , n62867 , n62872 , n62873 );
and ( n62875 , n62857 , n62874 );
and ( n62876 , n62847 , n62874 );
or ( n62877 , n62858 , n62875 , n62876 );
and ( n62878 , n62845 , n62877 );
and ( n62879 , n62831 , n62877 );
or ( n62880 , n62846 , n62878 , n62879 );
and ( n62881 , n57953 , n53972 );
and ( n62882 , n57688 , n53970 );
nor ( n62883 , n62881 , n62882 );
xnor ( n62884 , n62883 , n53662 );
and ( n62885 , n58117 , n53739 );
and ( n62886 , n57970 , n53737 );
nor ( n62887 , n62885 , n62886 );
xnor ( n62888 , n62887 , n53315 );
and ( n62889 , n62884 , n62888 );
and ( n62890 , n58171 , n53455 );
and ( n62891 , n58144 , n53453 );
nor ( n62892 , n62890 , n62891 );
xnor ( n62893 , n62892 , n53159 );
and ( n62894 , n62888 , n62893 );
and ( n62895 , n62884 , n62893 );
or ( n62896 , n62889 , n62894 , n62895 );
and ( n62897 , n58800 , n53293 );
and ( n62898 , n58571 , n53291 );
nor ( n62899 , n62897 , n62898 );
xnor ( n62900 , n62899 , n52963 );
and ( n62901 , n58864 , n53021 );
and ( n62902 , n58837 , n53019 );
nor ( n62903 , n62901 , n62902 );
xnor ( n62904 , n62903 , n52839 );
and ( n62905 , n62900 , n62904 );
nor ( n62906 , n52346 , n52344 );
xnor ( n62907 , n62906 , n52300 );
and ( n62908 , n62904 , n62907 );
and ( n62909 , n62900 , n62907 );
or ( n62910 , n62905 , n62908 , n62909 );
and ( n62911 , n62896 , n62910 );
xor ( n62912 , n62719 , n62723 );
xor ( n62913 , n62912 , n62728 );
and ( n62914 , n62910 , n62913 );
and ( n62915 , n62896 , n62913 );
or ( n62916 , n62911 , n62914 , n62915 );
xor ( n62917 , n62693 , n62694 );
xor ( n62918 , n62917 , n62697 );
and ( n62919 , n62916 , n62918 );
xor ( n62920 , n62710 , n62714 );
xor ( n62921 , n62920 , n62731 );
and ( n62922 , n62918 , n62921 );
and ( n62923 , n62916 , n62921 );
or ( n62924 , n62919 , n62922 , n62923 );
and ( n62925 , n62880 , n62924 );
xor ( n62926 , n62700 , n62734 );
xor ( n62927 , n62926 , n62759 );
and ( n62928 , n62924 , n62927 );
and ( n62929 , n62880 , n62927 );
or ( n62930 , n62925 , n62928 , n62929 );
and ( n62931 , n62828 , n62930 );
and ( n62932 , n62826 , n62930 );
or ( n62933 , n62829 , n62931 , n62932 );
xor ( n62934 , n62776 , n62778 );
xor ( n62935 , n62934 , n62781 );
and ( n62936 , n62933 , n62935 );
xor ( n62937 , n62691 , n62762 );
xor ( n62938 , n62937 , n62773 );
xor ( n62939 , n62765 , n62767 );
xor ( n62940 , n62939 , n62770 );
xor ( n62941 , n62751 , n62753 );
xor ( n62942 , n62941 , n62756 );
xor ( n62943 , n62739 , n62743 );
xor ( n62944 , n62943 , n62748 );
and ( n62945 , n52345 , n52300 );
xor ( n62946 , n62849 , n62851 );
xor ( n62947 , n62946 , n62854 );
and ( n62948 , n62945 , n62947 );
nor ( n62949 , n52886 , n52884 );
xnor ( n62950 , n62949 , n52657 );
nor ( n62951 , n52617 , n52615 );
xnor ( n62952 , n62951 , n52558 );
and ( n62953 , n62950 , n62952 );
nor ( n62954 , n52540 , n52538 );
xnor ( n62955 , n62954 , n52424 );
and ( n62956 , n62952 , n62955 );
and ( n62957 , n62950 , n62955 );
or ( n62958 , n62953 , n62956 , n62957 );
and ( n62959 , n62947 , n62958 );
and ( n62960 , n62945 , n62958 );
or ( n62961 , n62948 , n62959 , n62960 );
and ( n62962 , n62944 , n62961 );
and ( n62963 , n58864 , n53019 );
nor ( n62964 , n53021 , n62963 );
xnor ( n62965 , n62964 , n52839 );
and ( n62966 , n62965 , n52344 );
and ( n62967 , n57244 , n55033 );
and ( n62968 , n57027 , n55030 );
nor ( n62969 , n62967 , n62968 );
xnor ( n62970 , n62969 , n53885 );
and ( n62971 , n57519 , n54693 );
and ( n62972 , n57511 , n54691 );
nor ( n62973 , n62971 , n62972 );
xnor ( n62974 , n62973 , n53892 );
and ( n62975 , n62970 , n62974 );
and ( n62976 , n57688 , n54285 );
and ( n62977 , n57517 , n54283 );
nor ( n62978 , n62976 , n62977 );
xnor ( n62979 , n62978 , n53794 );
and ( n62980 , n62974 , n62979 );
and ( n62981 , n62970 , n62979 );
or ( n62982 , n62975 , n62980 , n62981 );
and ( n62983 , n62966 , n62982 );
and ( n62984 , n57970 , n53972 );
and ( n62985 , n57953 , n53970 );
nor ( n62986 , n62984 , n62985 );
xnor ( n62987 , n62986 , n53662 );
and ( n62988 , n58144 , n53739 );
and ( n62989 , n58117 , n53737 );
nor ( n62990 , n62988 , n62989 );
xnor ( n62991 , n62990 , n53315 );
and ( n62992 , n62987 , n62991 );
and ( n62993 , n58571 , n53455 );
and ( n62994 , n58171 , n53453 );
nor ( n62995 , n62993 , n62994 );
xnor ( n62996 , n62995 , n53159 );
and ( n62997 , n62991 , n62996 );
and ( n62998 , n62987 , n62996 );
or ( n62999 , n62992 , n62997 , n62998 );
and ( n63000 , n62982 , n62999 );
and ( n63001 , n62966 , n62999 );
or ( n63002 , n62983 , n63000 , n63001 );
and ( n63003 , n62961 , n63002 );
and ( n63004 , n62944 , n63002 );
or ( n63005 , n62962 , n63003 , n63004 );
and ( n63006 , n62942 , n63005 );
xor ( n63007 , n62862 , n62866 );
xor ( n63008 , n63007 , n62871 );
xor ( n63009 , n62884 , n62888 );
xor ( n63010 , n63009 , n62893 );
and ( n63011 , n63008 , n63010 );
xor ( n63012 , n62900 , n62904 );
xor ( n63013 , n63012 , n62907 );
and ( n63014 , n63010 , n63013 );
and ( n63015 , n63008 , n63013 );
or ( n63016 , n63011 , n63014 , n63015 );
xor ( n63017 , n62835 , n62839 );
xor ( n63018 , n63017 , n62842 );
and ( n63019 , n63016 , n63018 );
xor ( n63020 , n62847 , n62857 );
xor ( n63021 , n63020 , n62874 );
and ( n63022 , n63018 , n63021 );
and ( n63023 , n63016 , n63021 );
or ( n63024 , n63019 , n63022 , n63023 );
and ( n63025 , n63005 , n63024 );
and ( n63026 , n62942 , n63024 );
or ( n63027 , n63006 , n63025 , n63026 );
and ( n63028 , n62940 , n63027 );
xor ( n63029 , n62880 , n62924 );
xor ( n63030 , n63029 , n62927 );
and ( n63031 , n63027 , n63030 );
and ( n63032 , n62940 , n63030 );
or ( n63033 , n63028 , n63031 , n63032 );
and ( n63034 , n62938 , n63033 );
xor ( n63035 , n62826 , n62828 );
xor ( n63036 , n63035 , n62930 );
and ( n63037 , n63033 , n63036 );
and ( n63038 , n62938 , n63036 );
or ( n63039 , n63034 , n63037 , n63038 );
and ( n63040 , n62935 , n63039 );
and ( n63041 , n62933 , n63039 );
or ( n63042 , n62936 , n63040 , n63041 );
and ( n63043 , n62824 , n63042 );
xor ( n63044 , n62824 , n63042 );
xor ( n63045 , n62933 , n62935 );
xor ( n63046 , n63045 , n63039 );
xor ( n63047 , n62938 , n63033 );
xor ( n63048 , n63047 , n63036 );
xor ( n63049 , n62831 , n62845 );
xor ( n63050 , n63049 , n62877 );
xor ( n63051 , n62916 , n62918 );
xor ( n63052 , n63051 , n62921 );
and ( n63053 , n63050 , n63052 );
xor ( n63054 , n62896 , n62910 );
xor ( n63055 , n63054 , n62913 );
and ( n63056 , n58837 , n53293 );
and ( n63057 , n58800 , n53291 );
nor ( n63058 , n63056 , n63057 );
xnor ( n63059 , n63058 , n52963 );
xor ( n63060 , n62950 , n62952 );
xor ( n63061 , n63060 , n62955 );
and ( n63062 , n63059 , n63061 );
xor ( n63063 , n62965 , n52344 );
and ( n63064 , n63061 , n63063 );
and ( n63065 , n63059 , n63063 );
or ( n63066 , n63062 , n63064 , n63065 );
nor ( n63067 , n52886 , n52884 );
xnor ( n63068 , n63067 , n52657 );
nor ( n63069 , n52617 , n52615 );
xnor ( n63070 , n63069 , n52558 );
and ( n63071 , n63068 , n63070 );
nor ( n63072 , n52540 , n52538 );
xnor ( n63073 , n63072 , n52424 );
and ( n63074 , n63070 , n63073 );
and ( n63075 , n63068 , n63073 );
or ( n63076 , n63071 , n63074 , n63075 );
nor ( n63077 , n53021 , n53019 );
xnor ( n63078 , n63077 , n52839 );
and ( n63079 , n52539 , n52424 );
and ( n63080 , n63078 , n63079 );
and ( n63081 , n63076 , n63080 );
and ( n63082 , n57511 , n55033 );
and ( n63083 , n57244 , n55030 );
nor ( n63084 , n63082 , n63083 );
xnor ( n63085 , n63084 , n53885 );
and ( n63086 , n57517 , n54693 );
and ( n63087 , n57519 , n54691 );
nor ( n63088 , n63086 , n63087 );
xnor ( n63089 , n63088 , n53892 );
and ( n63090 , n63085 , n63089 );
and ( n63091 , n57953 , n54285 );
and ( n63092 , n57688 , n54283 );
nor ( n63093 , n63091 , n63092 );
xnor ( n63094 , n63093 , n53794 );
and ( n63095 , n63089 , n63094 );
and ( n63096 , n63085 , n63094 );
or ( n63097 , n63090 , n63095 , n63096 );
and ( n63098 , n63080 , n63097 );
and ( n63099 , n63076 , n63097 );
or ( n63100 , n63081 , n63098 , n63099 );
and ( n63101 , n63066 , n63100 );
and ( n63102 , n58117 , n53972 );
and ( n63103 , n57970 , n53970 );
nor ( n63104 , n63102 , n63103 );
xnor ( n63105 , n63104 , n53662 );
and ( n63106 , n58171 , n53739 );
and ( n63107 , n58144 , n53737 );
nor ( n63108 , n63106 , n63107 );
xnor ( n63109 , n63108 , n53315 );
and ( n63110 , n63105 , n63109 );
and ( n63111 , n58800 , n53455 );
and ( n63112 , n58571 , n53453 );
nor ( n63113 , n63111 , n63112 );
xnor ( n63114 , n63113 , n53159 );
and ( n63115 , n63109 , n63114 );
and ( n63116 , n63105 , n63114 );
or ( n63117 , n63110 , n63115 , n63116 );
xor ( n63118 , n62970 , n62974 );
xor ( n63119 , n63118 , n62979 );
and ( n63120 , n63117 , n63119 );
xor ( n63121 , n62987 , n62991 );
xor ( n63122 , n63121 , n62996 );
and ( n63123 , n63119 , n63122 );
and ( n63124 , n63117 , n63122 );
or ( n63125 , n63120 , n63123 , n63124 );
and ( n63126 , n63100 , n63125 );
and ( n63127 , n63066 , n63125 );
or ( n63128 , n63101 , n63126 , n63127 );
and ( n63129 , n63055 , n63128 );
xor ( n63130 , n62945 , n62947 );
xor ( n63131 , n63130 , n62958 );
xor ( n63132 , n62966 , n62982 );
xor ( n63133 , n63132 , n62999 );
and ( n63134 , n63131 , n63133 );
xor ( n63135 , n63008 , n63010 );
xor ( n63136 , n63135 , n63013 );
and ( n63137 , n63133 , n63136 );
and ( n63138 , n63131 , n63136 );
or ( n63139 , n63134 , n63137 , n63138 );
and ( n63140 , n63128 , n63139 );
and ( n63141 , n63055 , n63139 );
or ( n63142 , n63129 , n63140 , n63141 );
and ( n63143 , n63052 , n63142 );
and ( n63144 , n63050 , n63142 );
or ( n63145 , n63053 , n63143 , n63144 );
xor ( n63146 , n62940 , n63027 );
xor ( n63147 , n63146 , n63030 );
and ( n63148 , n63145 , n63147 );
xor ( n63149 , n62942 , n63005 );
xor ( n63150 , n63149 , n63024 );
xor ( n63151 , n62944 , n62961 );
xor ( n63152 , n63151 , n63002 );
xor ( n63153 , n63016 , n63018 );
xor ( n63154 , n63153 , n63021 );
and ( n63155 , n63152 , n63154 );
and ( n63156 , n58864 , n53291 );
nor ( n63157 , n53293 , n63156 );
xnor ( n63158 , n63157 , n52963 );
nor ( n63159 , n53021 , n53019 );
xnor ( n63160 , n63159 , n52839 );
and ( n63161 , n63158 , n63160 );
and ( n63162 , n63160 , n52538 );
and ( n63163 , n63158 , n52538 );
or ( n63164 , n63161 , n63162 , n63163 );
xor ( n63165 , n63078 , n63079 );
and ( n63166 , n63164 , n63165 );
and ( n63167 , n58864 , n53293 );
and ( n63168 , n58837 , n53291 );
nor ( n63169 , n63167 , n63168 );
xnor ( n63170 , n63169 , n52963 );
xor ( n63171 , n63068 , n63070 );
xor ( n63172 , n63171 , n63073 );
and ( n63173 , n63170 , n63172 );
and ( n63174 , n63166 , n63173 );
and ( n63175 , n57519 , n55033 );
and ( n63176 , n57511 , n55030 );
nor ( n63177 , n63175 , n63176 );
xnor ( n63178 , n63177 , n53885 );
and ( n63179 , n57688 , n54693 );
and ( n63180 , n57517 , n54691 );
nor ( n63181 , n63179 , n63180 );
xnor ( n63182 , n63181 , n53892 );
and ( n63183 , n63178 , n63182 );
and ( n63184 , n57970 , n54285 );
and ( n63185 , n57953 , n54283 );
nor ( n63186 , n63184 , n63185 );
xnor ( n63187 , n63186 , n53794 );
and ( n63188 , n63182 , n63187 );
and ( n63189 , n63178 , n63187 );
or ( n63190 , n63183 , n63188 , n63189 );
and ( n63191 , n58144 , n53972 );
and ( n63192 , n58117 , n53970 );
nor ( n63193 , n63191 , n63192 );
xnor ( n63194 , n63193 , n53662 );
and ( n63195 , n58571 , n53739 );
and ( n63196 , n58171 , n53737 );
nor ( n63197 , n63195 , n63196 );
xnor ( n63198 , n63197 , n53315 );
and ( n63199 , n63194 , n63198 );
and ( n63200 , n58837 , n53455 );
and ( n63201 , n58800 , n53453 );
nor ( n63202 , n63200 , n63201 );
xnor ( n63203 , n63202 , n53159 );
and ( n63204 , n63198 , n63203 );
and ( n63205 , n63194 , n63203 );
or ( n63206 , n63199 , n63204 , n63205 );
and ( n63207 , n63190 , n63206 );
xor ( n63208 , n63085 , n63089 );
xor ( n63209 , n63208 , n63094 );
and ( n63210 , n63206 , n63209 );
and ( n63211 , n63190 , n63209 );
or ( n63212 , n63207 , n63210 , n63211 );
and ( n63213 , n63173 , n63212 );
and ( n63214 , n63166 , n63212 );
or ( n63215 , n63174 , n63213 , n63214 );
xor ( n63216 , n63059 , n63061 );
xor ( n63217 , n63216 , n63063 );
xor ( n63218 , n63076 , n63080 );
xor ( n63219 , n63218 , n63097 );
and ( n63220 , n63217 , n63219 );
xor ( n63221 , n63117 , n63119 );
xor ( n63222 , n63221 , n63122 );
and ( n63223 , n63219 , n63222 );
and ( n63224 , n63217 , n63222 );
or ( n63225 , n63220 , n63223 , n63224 );
and ( n63226 , n63215 , n63225 );
xor ( n63227 , n63066 , n63100 );
xor ( n63228 , n63227 , n63125 );
and ( n63229 , n63225 , n63228 );
and ( n63230 , n63215 , n63228 );
or ( n63231 , n63226 , n63229 , n63230 );
and ( n63232 , n63154 , n63231 );
and ( n63233 , n63152 , n63231 );
or ( n63234 , n63155 , n63232 , n63233 );
and ( n63235 , n63150 , n63234 );
xor ( n63236 , n63050 , n63052 );
xor ( n63237 , n63236 , n63142 );
and ( n63238 , n63234 , n63237 );
and ( n63239 , n63150 , n63237 );
or ( n63240 , n63235 , n63238 , n63239 );
and ( n63241 , n63147 , n63240 );
and ( n63242 , n63145 , n63240 );
or ( n63243 , n63148 , n63241 , n63242 );
and ( n63244 , n63048 , n63243 );
xor ( n63245 , n63048 , n63243 );
xor ( n63246 , n63145 , n63147 );
xor ( n63247 , n63246 , n63240 );
xor ( n63248 , n63055 , n63128 );
xor ( n63249 , n63248 , n63139 );
xor ( n63250 , n63131 , n63133 );
xor ( n63251 , n63250 , n63136 );
xor ( n63252 , n63105 , n63109 );
xor ( n63253 , n63252 , n63114 );
xor ( n63254 , n63164 , n63165 );
and ( n63255 , n63253 , n63254 );
xor ( n63256 , n63170 , n63172 );
and ( n63257 , n63254 , n63256 );
and ( n63258 , n63253 , n63256 );
or ( n63259 , n63255 , n63257 , n63258 );
nor ( n63260 , n52886 , n52884 );
xnor ( n63261 , n63260 , n52657 );
nor ( n63262 , n52617 , n52615 );
xnor ( n63263 , n63262 , n52558 );
and ( n63264 , n63261 , n63263 );
xor ( n63265 , n63158 , n63160 );
xor ( n63266 , n63265 , n52538 );
and ( n63267 , n63263 , n63266 );
and ( n63268 , n63261 , n63266 );
or ( n63269 , n63264 , n63267 , n63268 );
nor ( n63270 , n53293 , n53291 );
xnor ( n63271 , n63270 , n52963 );
nor ( n63272 , n53021 , n53019 );
xnor ( n63273 , n63272 , n52839 );
and ( n63274 , n63271 , n63273 );
nor ( n63275 , n52886 , n52884 );
xnor ( n63276 , n63275 , n52657 );
and ( n63277 , n63273 , n63276 );
and ( n63278 , n63271 , n63276 );
or ( n63279 , n63274 , n63277 , n63278 );
and ( n63280 , n57517 , n55033 );
and ( n63281 , n57519 , n55030 );
nor ( n63282 , n63280 , n63281 );
xnor ( n63283 , n63282 , n53885 );
and ( n63284 , n57953 , n54693 );
and ( n63285 , n57688 , n54691 );
nor ( n63286 , n63284 , n63285 );
xnor ( n63287 , n63286 , n53892 );
and ( n63288 , n63283 , n63287 );
and ( n63289 , n58117 , n54285 );
and ( n63290 , n57970 , n54283 );
nor ( n63291 , n63289 , n63290 );
xnor ( n63292 , n63291 , n53794 );
and ( n63293 , n63287 , n63292 );
and ( n63294 , n63283 , n63292 );
or ( n63295 , n63288 , n63293 , n63294 );
and ( n63296 , n63279 , n63295 );
and ( n63297 , n58171 , n53972 );
and ( n63298 , n58144 , n53970 );
nor ( n63299 , n63297 , n63298 );
xnor ( n63300 , n63299 , n53662 );
and ( n63301 , n58800 , n53739 );
and ( n63302 , n58571 , n53737 );
nor ( n63303 , n63301 , n63302 );
xnor ( n63304 , n63303 , n53315 );
and ( n63305 , n63300 , n63304 );
and ( n63306 , n58864 , n53455 );
and ( n63307 , n58837 , n53453 );
nor ( n63308 , n63306 , n63307 );
xnor ( n63309 , n63308 , n53159 );
and ( n63310 , n63304 , n63309 );
and ( n63311 , n63300 , n63309 );
or ( n63312 , n63305 , n63310 , n63311 );
and ( n63313 , n63295 , n63312 );
and ( n63314 , n63279 , n63312 );
or ( n63315 , n63296 , n63313 , n63314 );
and ( n63316 , n63269 , n63315 );
xor ( n63317 , n63190 , n63206 );
xor ( n63318 , n63317 , n63209 );
and ( n63319 , n63315 , n63318 );
and ( n63320 , n63269 , n63318 );
or ( n63321 , n63316 , n63319 , n63320 );
and ( n63322 , n63259 , n63321 );
xor ( n63323 , n63166 , n63173 );
xor ( n63324 , n63323 , n63212 );
and ( n63325 , n63321 , n63324 );
and ( n63326 , n63259 , n63324 );
or ( n63327 , n63322 , n63325 , n63326 );
and ( n63328 , n63251 , n63327 );
xor ( n63329 , n63215 , n63225 );
xor ( n63330 , n63329 , n63228 );
and ( n63331 , n63327 , n63330 );
and ( n63332 , n63251 , n63330 );
or ( n63333 , n63328 , n63331 , n63332 );
and ( n63334 , n63249 , n63333 );
xor ( n63335 , n63152 , n63154 );
xor ( n63336 , n63335 , n63231 );
and ( n63337 , n63333 , n63336 );
and ( n63338 , n63249 , n63336 );
or ( n63339 , n63334 , n63337 , n63338 );
xor ( n63340 , n63150 , n63234 );
xor ( n63341 , n63340 , n63237 );
and ( n63342 , n63339 , n63341 );
xor ( n63343 , n63339 , n63341 );
xor ( n63344 , n63249 , n63333 );
xor ( n63345 , n63344 , n63336 );
xor ( n63346 , n63217 , n63219 );
xor ( n63347 , n63346 , n63222 );
xor ( n63348 , n63178 , n63182 );
xor ( n63349 , n63348 , n63187 );
xor ( n63350 , n63194 , n63198 );
xor ( n63351 , n63350 , n63203 );
and ( n63352 , n63349 , n63351 );
nor ( n63353 , n52617 , n52615 );
xnor ( n63354 , n63353 , n52558 );
and ( n63355 , n52616 , n52558 );
and ( n63356 , n63354 , n63355 );
xor ( n63357 , n63271 , n63273 );
xor ( n63358 , n63357 , n63276 );
and ( n63359 , n63355 , n63358 );
and ( n63360 , n63354 , n63358 );
or ( n63361 , n63356 , n63359 , n63360 );
and ( n63362 , n63351 , n63361 );
and ( n63363 , n63349 , n63361 );
or ( n63364 , n63352 , n63362 , n63363 );
nor ( n63365 , n53293 , n53291 );
xnor ( n63366 , n63365 , n52963 );
nor ( n63367 , n53021 , n53019 );
xnor ( n63368 , n63367 , n52839 );
and ( n63369 , n63366 , n63368 );
nor ( n63370 , n52886 , n52884 );
xnor ( n63371 , n63370 , n52657 );
and ( n63372 , n63368 , n63371 );
and ( n63373 , n63366 , n63371 );
or ( n63374 , n63369 , n63372 , n63373 );
and ( n63375 , n57688 , n55033 );
and ( n63376 , n57517 , n55030 );
nor ( n63377 , n63375 , n63376 );
xnor ( n63378 , n63377 , n53885 );
and ( n63379 , n57970 , n54693 );
and ( n63380 , n57953 , n54691 );
nor ( n63381 , n63379 , n63380 );
xnor ( n63382 , n63381 , n53892 );
and ( n63383 , n63378 , n63382 );
and ( n63384 , n58144 , n54285 );
and ( n63385 , n58117 , n54283 );
nor ( n63386 , n63384 , n63385 );
xnor ( n63387 , n63386 , n53794 );
and ( n63388 , n63382 , n63387 );
and ( n63389 , n63378 , n63387 );
or ( n63390 , n63383 , n63388 , n63389 );
and ( n63391 , n63374 , n63390 );
and ( n63392 , n58571 , n53972 );
and ( n63393 , n58171 , n53970 );
nor ( n63394 , n63392 , n63393 );
xnor ( n63395 , n63394 , n53662 );
and ( n63396 , n58837 , n53739 );
and ( n63397 , n58800 , n53737 );
nor ( n63398 , n63396 , n63397 );
xnor ( n63399 , n63398 , n53315 );
and ( n63400 , n63395 , n63399 );
and ( n63401 , n58864 , n53453 );
nor ( n63402 , n53455 , n63401 );
xnor ( n63403 , n63402 , n53159 );
and ( n63404 , n63399 , n63403 );
and ( n63405 , n63395 , n63403 );
or ( n63406 , n63400 , n63404 , n63405 );
and ( n63407 , n63390 , n63406 );
and ( n63408 , n63374 , n63406 );
or ( n63409 , n63391 , n63407 , n63408 );
xor ( n63410 , n63261 , n63263 );
xor ( n63411 , n63410 , n63266 );
and ( n63412 , n63409 , n63411 );
xor ( n63413 , n63279 , n63295 );
xor ( n63414 , n63413 , n63312 );
and ( n63415 , n63411 , n63414 );
and ( n63416 , n63409 , n63414 );
or ( n63417 , n63412 , n63415 , n63416 );
and ( n63418 , n63364 , n63417 );
xor ( n63419 , n63253 , n63254 );
xor ( n63420 , n63419 , n63256 );
and ( n63421 , n63417 , n63420 );
and ( n63422 , n63364 , n63420 );
or ( n63423 , n63418 , n63421 , n63422 );
and ( n63424 , n63347 , n63423 );
xor ( n63425 , n63259 , n63321 );
xor ( n63426 , n63425 , n63324 );
and ( n63427 , n63423 , n63426 );
and ( n63428 , n63347 , n63426 );
or ( n63429 , n63424 , n63427 , n63428 );
xor ( n63430 , n63251 , n63327 );
xor ( n63431 , n63430 , n63330 );
and ( n63432 , n63429 , n63431 );
xor ( n63433 , n63429 , n63431 );
xor ( n63434 , n63269 , n63315 );
xor ( n63435 , n63434 , n63318 );
xor ( n63436 , n63283 , n63287 );
xor ( n63437 , n63436 , n63292 );
xor ( n63438 , n63300 , n63304 );
xor ( n63439 , n63438 , n63309 );
and ( n63440 , n63437 , n63439 );
xor ( n63441 , n63366 , n63368 );
xor ( n63442 , n63441 , n63371 );
and ( n63443 , n52615 , n63442 );
nor ( n63444 , n53455 , n53453 );
xnor ( n63445 , n63444 , n53159 );
nor ( n63446 , n53293 , n53291 );
xnor ( n63447 , n63446 , n52963 );
and ( n63448 , n63445 , n63447 );
nor ( n63449 , n53021 , n53019 );
xnor ( n63450 , n63449 , n52839 );
and ( n63451 , n63447 , n63450 );
and ( n63452 , n63445 , n63450 );
or ( n63453 , n63448 , n63451 , n63452 );
and ( n63454 , n63442 , n63453 );
and ( n63455 , n52615 , n63453 );
or ( n63456 , n63443 , n63454 , n63455 );
and ( n63457 , n63439 , n63456 );
and ( n63458 , n63437 , n63456 );
or ( n63459 , n63440 , n63457 , n63458 );
and ( n63460 , n57953 , n55033 );
and ( n63461 , n57688 , n55030 );
nor ( n63462 , n63460 , n63461 );
xnor ( n63463 , n63462 , n53885 );
and ( n63464 , n58117 , n54693 );
and ( n63465 , n57970 , n54691 );
nor ( n63466 , n63464 , n63465 );
xnor ( n63467 , n63466 , n53892 );
and ( n63468 , n63463 , n63467 );
and ( n63469 , n58171 , n54285 );
and ( n63470 , n58144 , n54283 );
nor ( n63471 , n63469 , n63470 );
xnor ( n63472 , n63471 , n53794 );
and ( n63473 , n63467 , n63472 );
and ( n63474 , n63463 , n63472 );
or ( n63475 , n63468 , n63473 , n63474 );
and ( n63476 , n58800 , n53972 );
and ( n63477 , n58571 , n53970 );
nor ( n63478 , n63476 , n63477 );
xnor ( n63479 , n63478 , n53662 );
and ( n63480 , n58864 , n53739 );
and ( n63481 , n58837 , n53737 );
nor ( n63482 , n63480 , n63481 );
xnor ( n63483 , n63482 , n53315 );
and ( n63484 , n63479 , n63483 );
nor ( n63485 , n52886 , n52884 );
xnor ( n63486 , n63485 , n52657 );
and ( n63487 , n63483 , n63486 );
and ( n63488 , n63479 , n63486 );
or ( n63489 , n63484 , n63487 , n63488 );
and ( n63490 , n63475 , n63489 );
xor ( n63491 , n63378 , n63382 );
xor ( n63492 , n63491 , n63387 );
and ( n63493 , n63489 , n63492 );
and ( n63494 , n63475 , n63492 );
or ( n63495 , n63490 , n63493 , n63494 );
xor ( n63496 , n63354 , n63355 );
xor ( n63497 , n63496 , n63358 );
and ( n63498 , n63495 , n63497 );
xor ( n63499 , n63374 , n63390 );
xor ( n63500 , n63499 , n63406 );
and ( n63501 , n63497 , n63500 );
and ( n63502 , n63495 , n63500 );
or ( n63503 , n63498 , n63501 , n63502 );
and ( n63504 , n63459 , n63503 );
xor ( n63505 , n63349 , n63351 );
xor ( n63506 , n63505 , n63361 );
and ( n63507 , n63503 , n63506 );
and ( n63508 , n63459 , n63506 );
or ( n63509 , n63504 , n63507 , n63508 );
and ( n63510 , n63435 , n63509 );
xor ( n63511 , n63364 , n63417 );
xor ( n63512 , n63511 , n63420 );
and ( n63513 , n63509 , n63512 );
and ( n63514 , n63435 , n63512 );
or ( n63515 , n63510 , n63513 , n63514 );
xor ( n63516 , n63347 , n63423 );
xor ( n63517 , n63516 , n63426 );
and ( n63518 , n63515 , n63517 );
xor ( n63519 , n63515 , n63517 );
xor ( n63520 , n63409 , n63411 );
xor ( n63521 , n63520 , n63414 );
xor ( n63522 , n63395 , n63399 );
xor ( n63523 , n63522 , n63403 );
and ( n63524 , n52885 , n52657 );
xor ( n63525 , n63445 , n63447 );
xor ( n63526 , n63525 , n63450 );
and ( n63527 , n63524 , n63526 );
nor ( n63528 , n53455 , n53453 );
xnor ( n63529 , n63528 , n53159 );
nor ( n63530 , n53293 , n53291 );
xnor ( n63531 , n63530 , n52963 );
and ( n63532 , n63529 , n63531 );
nor ( n63533 , n53021 , n53019 );
xnor ( n63534 , n63533 , n52839 );
and ( n63535 , n63531 , n63534 );
and ( n63536 , n63529 , n63534 );
or ( n63537 , n63532 , n63535 , n63536 );
and ( n63538 , n63526 , n63537 );
and ( n63539 , n63524 , n63537 );
or ( n63540 , n63527 , n63538 , n63539 );
and ( n63541 , n63523 , n63540 );
and ( n63542 , n58864 , n53737 );
nor ( n63543 , n53739 , n63542 );
xnor ( n63544 , n63543 , n53315 );
and ( n63545 , n63544 , n52884 );
and ( n63546 , n57970 , n55033 );
and ( n63547 , n57953 , n55030 );
nor ( n63548 , n63546 , n63547 );
xnor ( n63549 , n63548 , n53885 );
and ( n63550 , n58144 , n54693 );
and ( n63551 , n58117 , n54691 );
nor ( n63552 , n63550 , n63551 );
xnor ( n63553 , n63552 , n53892 );
and ( n63554 , n63549 , n63553 );
and ( n63555 , n58571 , n54285 );
and ( n63556 , n58171 , n54283 );
nor ( n63557 , n63555 , n63556 );
xnor ( n63558 , n63557 , n53794 );
and ( n63559 , n63553 , n63558 );
and ( n63560 , n63549 , n63558 );
or ( n63561 , n63554 , n63559 , n63560 );
and ( n63562 , n63545 , n63561 );
xor ( n63563 , n63463 , n63467 );
xor ( n63564 , n63563 , n63472 );
and ( n63565 , n63561 , n63564 );
and ( n63566 , n63545 , n63564 );
or ( n63567 , n63562 , n63565 , n63566 );
and ( n63568 , n63540 , n63567 );
and ( n63569 , n63523 , n63567 );
or ( n63570 , n63541 , n63568 , n63569 );
xor ( n63571 , n63437 , n63439 );
xor ( n63572 , n63571 , n63456 );
and ( n63573 , n63570 , n63572 );
xor ( n63574 , n63495 , n63497 );
xor ( n63575 , n63574 , n63500 );
and ( n63576 , n63572 , n63575 );
and ( n63577 , n63570 , n63575 );
or ( n63578 , n63573 , n63576 , n63577 );
and ( n63579 , n63521 , n63578 );
xor ( n63580 , n63459 , n63503 );
xor ( n63581 , n63580 , n63506 );
and ( n63582 , n63578 , n63581 );
and ( n63583 , n63521 , n63581 );
or ( n63584 , n63579 , n63582 , n63583 );
xor ( n63585 , n63435 , n63509 );
xor ( n63586 , n63585 , n63512 );
and ( n63587 , n63584 , n63586 );
xor ( n63588 , n63584 , n63586 );
xor ( n63589 , n63521 , n63578 );
xor ( n63590 , n63589 , n63581 );
xor ( n63591 , n52615 , n63442 );
xor ( n63592 , n63591 , n63453 );
xor ( n63593 , n63475 , n63489 );
xor ( n63594 , n63593 , n63492 );
and ( n63595 , n63592 , n63594 );
xor ( n63596 , n63479 , n63483 );
xor ( n63597 , n63596 , n63486 );
and ( n63598 , n58837 , n53972 );
and ( n63599 , n58800 , n53970 );
nor ( n63600 , n63598 , n63599 );
xnor ( n63601 , n63600 , n53662 );
xor ( n63602 , n63529 , n63531 );
xor ( n63603 , n63602 , n63534 );
and ( n63604 , n63601 , n63603 );
xor ( n63605 , n63544 , n52884 );
and ( n63606 , n63603 , n63605 );
and ( n63607 , n63601 , n63605 );
or ( n63608 , n63604 , n63606 , n63607 );
and ( n63609 , n63597 , n63608 );
nor ( n63610 , n53739 , n53737 );
xnor ( n63611 , n63610 , n53315 );
nor ( n63612 , n53455 , n53453 );
xnor ( n63613 , n63612 , n53159 );
and ( n63614 , n63611 , n63613 );
nor ( n63615 , n53293 , n53291 );
xnor ( n63616 , n63615 , n52963 );
and ( n63617 , n63613 , n63616 );
and ( n63618 , n63611 , n63616 );
or ( n63619 , n63614 , n63617 , n63618 );
and ( n63620 , n58117 , n55033 );
and ( n63621 , n57970 , n55030 );
nor ( n63622 , n63620 , n63621 );
xnor ( n63623 , n63622 , n53885 );
and ( n63624 , n58171 , n54693 );
and ( n63625 , n58144 , n54691 );
nor ( n63626 , n63624 , n63625 );
xnor ( n63627 , n63626 , n53892 );
and ( n63628 , n63623 , n63627 );
and ( n63629 , n58800 , n54285 );
and ( n63630 , n58571 , n54283 );
nor ( n63631 , n63629 , n63630 );
xnor ( n63632 , n63631 , n53794 );
and ( n63633 , n63627 , n63632 );
and ( n63634 , n63623 , n63632 );
or ( n63635 , n63628 , n63633 , n63634 );
and ( n63636 , n63619 , n63635 );
and ( n63637 , n58864 , n53972 );
and ( n63638 , n58837 , n53970 );
nor ( n63639 , n63637 , n63638 );
xnor ( n63640 , n63639 , n53662 );
nor ( n63641 , n53021 , n53019 );
xnor ( n63642 , n63641 , n52839 );
and ( n63643 , n63640 , n63642 );
and ( n63644 , n53020 , n52839 );
and ( n63645 , n63642 , n63644 );
and ( n63646 , n63640 , n63644 );
or ( n63647 , n63643 , n63645 , n63646 );
and ( n63648 , n63635 , n63647 );
and ( n63649 , n63619 , n63647 );
or ( n63650 , n63636 , n63648 , n63649 );
and ( n63651 , n63608 , n63650 );
and ( n63652 , n63597 , n63650 );
or ( n63653 , n63609 , n63651 , n63652 );
and ( n63654 , n63594 , n63653 );
and ( n63655 , n63592 , n63653 );
or ( n63656 , n63595 , n63654 , n63655 );
xor ( n63657 , n63570 , n63572 );
xor ( n63658 , n63657 , n63575 );
and ( n63659 , n63656 , n63658 );
xor ( n63660 , n63523 , n63540 );
xor ( n63661 , n63660 , n63567 );
xor ( n63662 , n63524 , n63526 );
xor ( n63663 , n63662 , n63537 );
xor ( n63664 , n63545 , n63561 );
xor ( n63665 , n63664 , n63564 );
and ( n63666 , n63663 , n63665 );
xor ( n63667 , n63549 , n63553 );
xor ( n63668 , n63667 , n63558 );
xor ( n63669 , n63611 , n63613 );
xor ( n63670 , n63669 , n63616 );
nor ( n63671 , n53739 , n53737 );
xnor ( n63672 , n63671 , n53315 );
nor ( n63673 , n53455 , n53453 );
xnor ( n63674 , n63673 , n53159 );
and ( n63675 , n63672 , n63674 );
nor ( n63676 , n53293 , n53291 );
xnor ( n63677 , n63676 , n52963 );
and ( n63678 , n63674 , n63677 );
and ( n63679 , n63672 , n63677 );
or ( n63680 , n63675 , n63678 , n63679 );
and ( n63681 , n63670 , n63680 );
xor ( n63682 , n63623 , n63627 );
xor ( n63683 , n63682 , n63632 );
and ( n63684 , n63680 , n63683 );
and ( n63685 , n63670 , n63683 );
or ( n63686 , n63681 , n63684 , n63685 );
and ( n63687 , n63668 , n63686 );
xor ( n63688 , n63601 , n63603 );
xor ( n63689 , n63688 , n63605 );
and ( n63690 , n63686 , n63689 );
and ( n63691 , n63668 , n63689 );
or ( n63692 , n63687 , n63690 , n63691 );
and ( n63693 , n63665 , n63692 );
and ( n63694 , n63663 , n63692 );
or ( n63695 , n63666 , n63693 , n63694 );
and ( n63696 , n63661 , n63695 );
xor ( n63697 , n63592 , n63594 );
xor ( n63698 , n63697 , n63653 );
and ( n63699 , n63695 , n63698 );
and ( n63700 , n63661 , n63698 );
or ( n63701 , n63696 , n63699 , n63700 );
and ( n63702 , n63658 , n63701 );
and ( n63703 , n63656 , n63701 );
or ( n63704 , n63659 , n63702 , n63703 );
and ( n63705 , n63590 , n63704 );
xor ( n63706 , n63590 , n63704 );
xor ( n63707 , n63656 , n63658 );
xor ( n63708 , n63707 , n63701 );
xor ( n63709 , n63597 , n63608 );
xor ( n63710 , n63709 , n63650 );
xor ( n63711 , n63619 , n63635 );
xor ( n63712 , n63711 , n63647 );
xor ( n63713 , n63640 , n63642 );
xor ( n63714 , n63713 , n63644 );
nor ( n63715 , n53972 , n53970 );
xnor ( n63716 , n63715 , n53662 );
and ( n63717 , n53292 , n52963 );
and ( n63718 , n63716 , n63717 );
and ( n63719 , n58864 , n53970 );
nor ( n63720 , n53972 , n63719 );
xnor ( n63721 , n63720 , n53662 );
and ( n63722 , n63718 , n63721 );
and ( n63723 , n63721 , n53019 );
and ( n63724 , n63718 , n53019 );
or ( n63725 , n63722 , n63723 , n63724 );
and ( n63726 , n63714 , n63725 );
xor ( n63727 , n63670 , n63680 );
xor ( n63728 , n63727 , n63683 );
and ( n63729 , n63725 , n63728 );
and ( n63730 , n63714 , n63728 );
or ( n63731 , n63726 , n63729 , n63730 );
and ( n63732 , n63712 , n63731 );
xor ( n63733 , n63668 , n63686 );
xor ( n63734 , n63733 , n63689 );
and ( n63735 , n63731 , n63734 );
and ( n63736 , n63712 , n63734 );
or ( n63737 , n63732 , n63735 , n63736 );
and ( n63738 , n63710 , n63737 );
xor ( n63739 , n63663 , n63665 );
xor ( n63740 , n63739 , n63692 );
and ( n63741 , n63737 , n63740 );
and ( n63742 , n63710 , n63740 );
or ( n63743 , n63738 , n63741 , n63742 );
xor ( n63744 , n63661 , n63695 );
xor ( n63745 , n63744 , n63698 );
and ( n63746 , n63743 , n63745 );
xor ( n63747 , n63743 , n63745 );
xor ( n63748 , n63710 , n63737 );
xor ( n63749 , n63748 , n63740 );
xor ( n63750 , n63712 , n63731 );
xor ( n63751 , n63750 , n63734 );
nor ( n63752 , n53739 , n53737 );
xnor ( n63753 , n63752 , n53315 );
nor ( n63754 , n53455 , n53453 );
xnor ( n63755 , n63754 , n53159 );
and ( n63756 , n63753 , n63755 );
nor ( n63757 , n53293 , n53291 );
xnor ( n63758 , n63757 , n52963 );
and ( n63759 , n63755 , n63758 );
and ( n63760 , n63753 , n63758 );
or ( n63761 , n63756 , n63759 , n63760 );
xor ( n63762 , n63672 , n63674 );
xor ( n63763 , n63762 , n63677 );
and ( n63764 , n63761 , n63763 );
xor ( n63765 , n63718 , n63721 );
xor ( n63766 , n63765 , n53019 );
and ( n63767 , n63763 , n63766 );
and ( n63768 , n63761 , n63766 );
or ( n63769 , n63764 , n63767 , n63768 );
xor ( n63770 , n63714 , n63725 );
xor ( n63771 , n63770 , n63728 );
and ( n63772 , n63769 , n63771 );
xor ( n63773 , n63716 , n63717 );
and ( n63774 , n58864 , n54283 );
nor ( n63775 , n54285 , n63774 );
xnor ( n63776 , n63775 , n53794 );
nor ( n63777 , n53972 , n53970 );
xnor ( n63778 , n63777 , n53662 );
and ( n63779 , n63776 , n63778 );
and ( n63780 , n63778 , n53291 );
and ( n63781 , n63776 , n53291 );
or ( n63782 , n63779 , n63780 , n63781 );
and ( n63783 , n63773 , n63782 );
nor ( n63784 , n54285 , n54283 );
xnor ( n63785 , n63784 , n53794 );
nor ( n63786 , n53972 , n53970 );
xnor ( n63787 , n63786 , n53662 );
and ( n63788 , n63785 , n63787 );
nor ( n63789 , n53739 , n53737 );
xnor ( n63790 , n63789 , n53315 );
and ( n63791 , n63788 , n63790 );
nor ( n63792 , n53455 , n53453 );
xnor ( n63793 , n63792 , n53159 );
and ( n63794 , n63790 , n63793 );
and ( n63795 , n63788 , n63793 );
or ( n63796 , n63791 , n63794 , n63795 );
and ( n63797 , n63782 , n63796 );
and ( n63798 , n63773 , n63796 );
or ( n63799 , n63783 , n63797 , n63798 );
and ( n63800 , n58837 , n54285 );
and ( n63801 , n58800 , n54283 );
nor ( n63802 , n63800 , n63801 );
xnor ( n63803 , n63802 , n53794 );
and ( n63804 , n63799 , n63803 );
xor ( n63805 , n63761 , n63763 );
xor ( n63806 , n63805 , n63766 );
and ( n63807 , n63803 , n63806 );
and ( n63808 , n63799 , n63806 );
or ( n63809 , n63804 , n63807 , n63808 );
and ( n63810 , n63771 , n63809 );
and ( n63811 , n63769 , n63809 );
or ( n63812 , n63772 , n63810 , n63811 );
and ( n63813 , n63751 , n63812 );
and ( n63814 , n58864 , n54285 );
and ( n63815 , n58837 , n54283 );
nor ( n63816 , n63814 , n63815 );
xnor ( n63817 , n63816 , n53794 );
xor ( n63818 , n63753 , n63755 );
xor ( n63819 , n63818 , n63758 );
and ( n63820 , n63817 , n63819 );
xor ( n63821 , n63773 , n63782 );
xor ( n63822 , n63821 , n63796 );
and ( n63823 , n63819 , n63822 );
and ( n63824 , n63817 , n63822 );
or ( n63825 , n63820 , n63823 , n63824 );
and ( n63826 , n58571 , n54693 );
and ( n63827 , n58171 , n54691 );
nor ( n63828 , n63826 , n63827 );
xnor ( n63829 , n63828 , n53892 );
and ( n63830 , n63825 , n63829 );
xor ( n63831 , n63799 , n63803 );
xor ( n63832 , n63831 , n63806 );
and ( n63833 , n63829 , n63832 );
and ( n63834 , n63825 , n63832 );
or ( n63835 , n63830 , n63833 , n63834 );
xor ( n63836 , n63769 , n63771 );
xor ( n63837 , n63836 , n63809 );
and ( n63838 , n63835 , n63837 );
xor ( n63839 , n63785 , n63787 );
nor ( n63840 , n53739 , n53737 );
xnor ( n63841 , n63840 , n53315 );
and ( n63842 , n63839 , n63841 );
and ( n63843 , n53454 , n53159 );
and ( n63844 , n63841 , n63843 );
and ( n63845 , n63839 , n63843 );
or ( n63846 , n63842 , n63844 , n63845 );
xor ( n63847 , n63776 , n63778 );
xor ( n63848 , n63847 , n53291 );
and ( n63849 , n63846 , n63848 );
xor ( n63850 , n63788 , n63790 );
xor ( n63851 , n63850 , n63793 );
and ( n63852 , n63848 , n63851 );
and ( n63853 , n63846 , n63851 );
or ( n63854 , n63849 , n63852 , n63853 );
and ( n63855 , n58800 , n54693 );
and ( n63856 , n58571 , n54691 );
nor ( n63857 , n63855 , n63856 );
xnor ( n63858 , n63857 , n53892 );
and ( n63859 , n63854 , n63858 );
xor ( n63860 , n63817 , n63819 );
xor ( n63861 , n63860 , n63822 );
and ( n63862 , n63858 , n63861 );
and ( n63863 , n63854 , n63861 );
or ( n63864 , n63859 , n63862 , n63863 );
xor ( n63865 , n63825 , n63829 );
xor ( n63866 , n63865 , n63832 );
and ( n63867 , n63864 , n63866 );
and ( n63868 , n63837 , n63867 );
and ( n63869 , n63835 , n63867 );
or ( n63870 , n63838 , n63868 , n63869 );
and ( n63871 , n63812 , n63870 );
and ( n63872 , n63751 , n63870 );
or ( n63873 , n63813 , n63871 , n63872 );
and ( n63874 , n63749 , n63873 );
xor ( n63875 , n63749 , n63873 );
xor ( n63876 , n63751 , n63812 );
xor ( n63877 , n63876 , n63870 );
and ( n63878 , n58144 , n55033 );
and ( n63879 , n58117 , n55030 );
nor ( n63880 , n63878 , n63879 );
xnor ( n63881 , n63880 , n53885 );
and ( n63882 , n58171 , n55033 );
and ( n63883 , n58144 , n55030 );
nor ( n63884 , n63882 , n63883 );
xnor ( n63885 , n63884 , n53885 );
and ( n63886 , n58571 , n55033 );
and ( n63887 , n58171 , n55030 );
nor ( n63888 , n63886 , n63887 );
xnor ( n63889 , n63888 , n53885 );
and ( n63890 , n58837 , n54693 );
and ( n63891 , n58800 , n54691 );
nor ( n63892 , n63890 , n63891 );
xnor ( n63893 , n63892 , n53892 );
and ( n63894 , n63889 , n63893 );
and ( n63895 , n58864 , n54691 );
nor ( n63896 , n54693 , n63895 );
xnor ( n63897 , n63896 , n53892 );
nor ( n63898 , n53972 , n53970 );
xnor ( n63899 , n63898 , n53662 );
and ( n63900 , n63897 , n63899 );
and ( n63901 , n63899 , n53453 );
and ( n63902 , n63897 , n53453 );
or ( n63903 , n63900 , n63901 , n63902 );
nor ( n63904 , n53455 , n53453 );
xnor ( n63905 , n63904 , n53159 );
and ( n63906 , n63903 , n63905 );
and ( n63907 , n63893 , n63906 );
and ( n63908 , n63889 , n63906 );
or ( n63909 , n63894 , n63907 , n63908 );
and ( n63910 , n63885 , n63909 );
xor ( n63911 , n63846 , n63848 );
xor ( n63912 , n63911 , n63851 );
and ( n63913 , n58864 , n54693 );
and ( n63914 , n58837 , n54691 );
nor ( n63915 , n63913 , n63914 );
xnor ( n63916 , n63915 , n53892 );
xor ( n63917 , n63839 , n63841 );
xor ( n63918 , n63917 , n63843 );
and ( n63919 , n63916 , n63918 );
and ( n63920 , n63912 , n63919 );
and ( n63921 , n58800 , n55033 );
and ( n63922 , n58571 , n55030 );
nor ( n63923 , n63921 , n63922 );
xnor ( n63924 , n63923 , n53885 );
and ( n63925 , n58837 , n55033 );
and ( n63926 , n58800 , n55030 );
nor ( n63927 , n63925 , n63926 );
xnor ( n63928 , n63927 , n53885 );
nor ( n63929 , n54285 , n54283 );
xnor ( n63930 , n63929 , n53794 );
and ( n63931 , n63928 , n63930 );
nor ( n63932 , n53739 , n53737 );
xnor ( n63933 , n63932 , n53315 );
and ( n63934 , n63930 , n63933 );
and ( n63935 , n63928 , n63933 );
or ( n63936 , n63931 , n63934 , n63935 );
and ( n63937 , n63924 , n63936 );
xor ( n63938 , n63903 , n63905 );
and ( n63939 , n63936 , n63938 );
and ( n63940 , n63924 , n63938 );
or ( n63941 , n63937 , n63939 , n63940 );
and ( n63942 , n63919 , n63941 );
and ( n63943 , n63912 , n63941 );
or ( n63944 , n63920 , n63942 , n63943 );
and ( n63945 , n63909 , n63944 );
and ( n63946 , n63885 , n63944 );
or ( n63947 , n63910 , n63945 , n63946 );
and ( n63948 , n63881 , n63947 );
xor ( n63949 , n63864 , n63866 );
and ( n63950 , n63947 , n63949 );
and ( n63951 , n63881 , n63949 );
or ( n63952 , n63948 , n63950 , n63951 );
xor ( n63953 , n63835 , n63837 );
xor ( n63954 , n63953 , n63867 );
and ( n63955 , n63952 , n63954 );
xor ( n63956 , n63952 , n63954 );
xor ( n63957 , n63854 , n63858 );
xor ( n63958 , n63957 , n63861 );
xor ( n63959 , n63889 , n63893 );
xor ( n63960 , n63959 , n63906 );
xor ( n63961 , n63897 , n63899 );
xor ( n63962 , n63961 , n53453 );
nor ( n63963 , n54693 , n54691 );
xnor ( n63964 , n63963 , n53892 );
nor ( n63965 , n54285 , n54283 );
xnor ( n63966 , n63965 , n53794 );
and ( n63967 , n63964 , n63966 );
nor ( n63968 , n53972 , n53970 );
xnor ( n63969 , n63968 , n53662 );
and ( n63970 , n63966 , n63969 );
and ( n63971 , n63964 , n63969 );
or ( n63972 , n63967 , n63970 , n63971 );
and ( n63973 , n63962 , n63972 );
and ( n63974 , n58864 , n55033 );
and ( n63975 , n58837 , n55030 );
nor ( n63976 , n63974 , n63975 );
xnor ( n63977 , n63976 , n53885 );
nor ( n63978 , n53739 , n53737 );
xnor ( n63979 , n63978 , n53315 );
and ( n63980 , n63977 , n63979 );
and ( n63981 , n53738 , n53315 );
and ( n63982 , n63979 , n63981 );
and ( n63983 , n63977 , n63981 );
or ( n63984 , n63980 , n63982 , n63983 );
and ( n63985 , n63972 , n63984 );
and ( n63986 , n63962 , n63984 );
or ( n63987 , n63973 , n63985 , n63986 );
xor ( n63988 , n63916 , n63918 );
and ( n63989 , n63987 , n63988 );
xor ( n63990 , n63928 , n63930 );
xor ( n63991 , n63990 , n63933 );
xor ( n63992 , n63964 , n63966 );
xor ( n63993 , n63992 , n63969 );
nor ( n63994 , n54693 , n54691 );
xnor ( n63995 , n63994 , n53892 );
nor ( n63996 , n54285 , n54283 );
xnor ( n63997 , n63996 , n53794 );
and ( n63998 , n63995 , n63997 );
nor ( n63999 , n53972 , n53970 );
xnor ( n64000 , n63999 , n53662 );
and ( n64001 , n63997 , n64000 );
and ( n64002 , n63995 , n64000 );
or ( n64003 , n63998 , n64001 , n64002 );
and ( n64004 , n63993 , n64003 );
and ( n64005 , n58864 , n55030 );
nor ( n64006 , n55033 , n64005 );
xnor ( n64007 , n64006 , n53885 );
and ( n64008 , n64007 , n53737 );
and ( n64009 , n64003 , n64008 );
and ( n64010 , n63993 , n64008 );
or ( n64011 , n64004 , n64009 , n64010 );
and ( n64012 , n63991 , n64011 );
xor ( n64013 , n63962 , n63972 );
xor ( n64014 , n64013 , n63984 );
and ( n64015 , n64011 , n64014 );
and ( n64016 , n63991 , n64014 );
or ( n64017 , n64012 , n64015 , n64016 );
and ( n64018 , n63988 , n64017 );
and ( n64019 , n63987 , n64017 );
or ( n64020 , n63989 , n64018 , n64019 );
and ( n64021 , n63960 , n64020 );
xor ( n64022 , n63912 , n63919 );
xor ( n64023 , n64022 , n63941 );
and ( n64024 , n64020 , n64023 );
and ( n64025 , n63960 , n64023 );
or ( n64026 , n64021 , n64024 , n64025 );
and ( n64027 , n63958 , n64026 );
xor ( n64028 , n63885 , n63909 );
xor ( n64029 , n64028 , n63944 );
and ( n64030 , n64026 , n64029 );
and ( n64031 , n63958 , n64029 );
or ( n64032 , n64027 , n64030 , n64031 );
xor ( n64033 , n63881 , n63947 );
xor ( n64034 , n64033 , n63949 );
and ( n64035 , n64032 , n64034 );
xor ( n64036 , n64032 , n64034 );
xor ( n64037 , n63958 , n64026 );
xor ( n64038 , n64037 , n64029 );
xor ( n64039 , n63960 , n64020 );
xor ( n64040 , n64039 , n64023 );
xor ( n64041 , n63924 , n63936 );
xor ( n64042 , n64041 , n63938 );
xor ( n64043 , n63987 , n63988 );
xor ( n64044 , n64043 , n64017 );
and ( n64045 , n64042 , n64044 );
xor ( n64046 , n64042 , n64044 );
xor ( n64047 , n63977 , n63979 );
xor ( n64048 , n64047 , n63981 );
xor ( n64049 , n63995 , n63997 );
xor ( n64050 , n64049 , n64000 );
xor ( n64051 , n64007 , n53737 );
and ( n64052 , n64050 , n64051 );
nor ( n64053 , n54693 , n54691 );
xnor ( n64054 , n64053 , n53892 );
nor ( n64055 , n54285 , n54283 );
xnor ( n64056 , n64055 , n53794 );
and ( n64057 , n64054 , n64056 );
nor ( n64058 , n53972 , n53970 );
xnor ( n64059 , n64058 , n53662 );
and ( n64060 , n64056 , n64059 );
and ( n64061 , n64054 , n64059 );
or ( n64062 , n64057 , n64060 , n64061 );
and ( n64063 , n64051 , n64062 );
and ( n64064 , n64050 , n64062 );
or ( n64065 , n64052 , n64063 , n64064 );
and ( n64066 , n64048 , n64065 );
xor ( n64067 , n63993 , n64003 );
xor ( n64068 , n64067 , n64008 );
and ( n64069 , n64065 , n64068 );
and ( n64070 , n64048 , n64068 );
or ( n64071 , n64066 , n64069 , n64070 );
xor ( n64072 , n63991 , n64011 );
xor ( n64073 , n64072 , n64014 );
and ( n64074 , n64071 , n64073 );
xor ( n64075 , n64071 , n64073 );
nor ( n64076 , n55033 , n55030 );
xnor ( n64077 , n64076 , n53885 );
and ( n64078 , n53971 , n53662 );
and ( n64079 , n64077 , n64078 );
xor ( n64080 , n64077 , n64078 );
nor ( n64081 , n55033 , n55030 );
xnor ( n64082 , n64081 , n53885 );
nor ( n64083 , n54693 , n54691 );
xnor ( n64084 , n64083 , n53892 );
and ( n64085 , n64082 , n64084 );
and ( n64086 , n64084 , n53970 );
and ( n64087 , n64082 , n53970 );
or ( n64088 , n64085 , n64086 , n64087 );
and ( n64089 , n64080 , n64088 );
xor ( n64090 , n64054 , n64056 );
xor ( n64091 , n64090 , n64059 );
and ( n64092 , n64088 , n64091 );
and ( n64093 , n64080 , n64091 );
or ( n64094 , n64089 , n64092 , n64093 );
and ( n64095 , n64079 , n64094 );
xor ( n64096 , n64050 , n64051 );
xor ( n64097 , n64096 , n64062 );
and ( n64098 , n64094 , n64097 );
and ( n64099 , n64079 , n64097 );
or ( n64100 , n64095 , n64098 , n64099 );
xor ( n64101 , n64048 , n64065 );
xor ( n64102 , n64101 , n64068 );
and ( n64103 , n64100 , n64102 );
xor ( n64104 , n64100 , n64102 );
xor ( n64105 , n64079 , n64094 );
xor ( n64106 , n64105 , n64097 );
xor ( n64107 , n64080 , n64088 );
xor ( n64108 , n64107 , n64091 );
nor ( n64109 , n55033 , n55030 );
xnor ( n64110 , n64109 , n53885 );
and ( n64111 , n54284 , n53794 );
and ( n64112 , n64110 , n64111 );
nor ( n64113 , n54285 , n54283 );
xnor ( n64114 , n64113 , n53794 );
and ( n64115 , n64112 , n64114 );
xor ( n64116 , n64082 , n64084 );
xor ( n64117 , n64116 , n53970 );
and ( n64118 , n64114 , n64117 );
and ( n64119 , n64112 , n64117 );
or ( n64120 , n64115 , n64118 , n64119 );
and ( n64121 , n64108 , n64120 );
xor ( n64122 , n64108 , n64120 );
xor ( n64123 , n64112 , n64114 );
xor ( n64124 , n64123 , n64117 );
xor ( n64125 , n64110 , n64111 );
nor ( n64126 , n54693 , n54691 );
xnor ( n64127 , n64126 , n53892 );
and ( n64128 , n64125 , n64127 );
nor ( n64129 , n54285 , n54283 );
xnor ( n64130 , n64129 , n53794 );
and ( n64131 , n64127 , n64130 );
and ( n64132 , n64125 , n64130 );
or ( n64133 , n64128 , n64131 , n64132 );
and ( n64134 , n64124 , n64133 );
xor ( n64135 , n64124 , n64133 );
nor ( n64136 , n55033 , n55030 );
xnor ( n64137 , n64136 , n53885 );
nor ( n64138 , n54693 , n54691 );
xnor ( n64139 , n64138 , n53892 );
and ( n64140 , n64137 , n64139 );
and ( n64141 , n64139 , n54283 );
and ( n64142 , n64137 , n54283 );
or ( n64143 , n64140 , n64141 , n64142 );
xor ( n64144 , n64125 , n64127 );
xor ( n64145 , n64144 , n64130 );
and ( n64146 , n64143 , n64145 );
xor ( n64147 , n64143 , n64145 );
xor ( n64148 , n64137 , n64139 );
xor ( n64149 , n64148 , n54283 );
nor ( n64150 , n55033 , n55030 );
xnor ( n64151 , n64150 , n53885 );
and ( n64152 , n54692 , n53892 );
and ( n64153 , n64151 , n64152 );
and ( n64154 , n64149 , n64153 );
xor ( n64155 , n64149 , n64153 );
nor ( n64156 , n54693 , n54691 );
xnor ( n64157 , n64156 , n53892 );
xor ( n64158 , n64151 , n64152 );
and ( n64159 , n64157 , n64158 );
xor ( n64160 , n64157 , n64158 );
nor ( n64161 , n55033 , n55030 );
xnor ( n64162 , n64161 , n53885 );
and ( n64163 , n64162 , n54691 );
xor ( n64164 , n64162 , n54691 );
nor ( n64165 , n55033 , n55030 );
xnor ( n64166 , n64165 , n53885 );
and ( n64167 , n55032 , n53885 );
and ( n64168 , n64166 , n64167 );
and ( n64169 , n64164 , n64168 );
or ( n64170 , n64163 , n64169 );
and ( n64171 , n64160 , n64170 );
or ( n64172 , n64159 , n64171 );
and ( n64173 , n64155 , n64172 );
or ( n64174 , n64154 , n64173 );
and ( n64175 , n64147 , n64174 );
or ( n64176 , n64146 , n64175 );
and ( n64177 , n64135 , n64176 );
or ( n64178 , n64134 , n64177 );
and ( n64179 , n64122 , n64178 );
or ( n64180 , n64121 , n64179 );
and ( n64181 , n64106 , n64180 );
and ( n64182 , n64104 , n64181 );
or ( n64183 , n64103 , n64182 );
and ( n64184 , n64075 , n64183 );
or ( n64185 , n64074 , n64184 );
and ( n64186 , n64046 , n64185 );
or ( n64187 , n64045 , n64186 );
and ( n64188 , n64040 , n64187 );
and ( n64189 , n64038 , n64188 );
and ( n64190 , n64036 , n64189 );
or ( n64191 , n64035 , n64190 );
and ( n64192 , n63956 , n64191 );
or ( n64193 , n63955 , n64192 );
and ( n64194 , n63877 , n64193 );
and ( n64195 , n63875 , n64194 );
or ( n64196 , n63874 , n64195 );
and ( n64197 , n63747 , n64196 );
or ( n64198 , n63746 , n64197 );
and ( n64199 , n63708 , n64198 );
and ( n64200 , n63706 , n64199 );
or ( n64201 , n63705 , n64200 );
and ( n64202 , n63588 , n64201 );
or ( n64203 , n63587 , n64202 );
and ( n64204 , n63519 , n64203 );
or ( n64205 , n63518 , n64204 );
and ( n64206 , n63433 , n64205 );
or ( n64207 , n63432 , n64206 );
and ( n64208 , n63345 , n64207 );
and ( n64209 , n63343 , n64208 );
or ( n64210 , n63342 , n64209 );
and ( n64211 , n63247 , n64210 );
and ( n64212 , n63245 , n64211 );
or ( n64213 , n63244 , n64212 );
and ( n64214 , n63046 , n64213 );
and ( n64215 , n63044 , n64214 );
or ( n64216 , n63043 , n64215 );
and ( n64217 , n62822 , n64216 );
and ( n64218 , n62820 , n64217 );
and ( n64219 , n62818 , n64218 );
and ( n64220 , n62816 , n64219 );
or ( n64221 , n62815 , n64220 );
and ( n64222 , n62685 , n64221 );
and ( n64223 , n62683 , n64222 );
or ( n64224 , n62682 , n64223 );
and ( n64225 , n62296 , n64224 );
and ( n64226 , n62294 , n64225 );
and ( n64227 , n62292 , n64226 );
and ( n64228 , n62290 , n64227 );
or ( n64229 , n62289 , n64228 );
and ( n64230 , n62185 , n64229 );
and ( n64231 , n62183 , n64230 );
and ( n64232 , n62181 , n64231 );
and ( n64233 , n62179 , n64232 );
and ( n64234 , n62177 , n64233 );
and ( n64235 , n62175 , n64234 );
and ( n64236 , n62173 , n64235 );
and ( n64237 , n62171 , n64236 );
and ( n64238 , n62169 , n64237 );
and ( n64239 , n62167 , n64238 );
and ( n64240 , n62165 , n64239 );
and ( n64241 , n62163 , n64240 );
and ( n64242 , n62161 , n64241 );
and ( n64243 , n62159 , n64242 );
and ( n64244 , n62157 , n64243 );
and ( n64245 , n62155 , n64244 );
and ( n64246 , n62153 , n64245 );
and ( n64247 , n62151 , n64246 );
and ( n64248 , n62149 , n64247 );
and ( n64249 , n62147 , n64248 );
and ( n64250 , n62145 , n64249 );
and ( n64251 , n62143 , n64250 );
and ( n64252 , n62141 , n64251 );
and ( n64253 , n62139 , n64252 );
and ( n64254 , n62137 , n64253 );
and ( n64255 , n62135 , n64254 );
and ( n64256 , n62133 , n64255 );
and ( n64257 , n62131 , n64256 );
and ( n64258 , n62129 , n64257 );
and ( n64259 , n62127 , n64258 );
and ( n64260 , n62125 , n64259 );
and ( n64261 , n62123 , n64260 );
and ( n64262 , n62121 , n64261 );
and ( n64263 , n62119 , n64262 );
and ( n64264 , n62117 , n64263 );
and ( n64265 , n62115 , n64264 );
and ( n64266 , n62113 , n64265 );
and ( n64267 , n62111 , n64266 );
and ( n64268 , n62109 , n64267 );
and ( n64269 , n62107 , n64268 );
and ( n64270 , n62105 , n64269 );
and ( n64271 , n62103 , n64270 );
and ( n64272 , n62101 , n64271 );
and ( n64273 , n62099 , n64272 );
and ( n64274 , n62097 , n64273 );
and ( n64275 , n62095 , n64274 );
and ( n64276 , n62093 , n64275 );
and ( n64277 , n62091 , n64276 );
and ( n64278 , n62089 , n64277 );
and ( n64279 , n62087 , n64278 );
and ( n64280 , n62085 , n64279 );
and ( n64281 , n62083 , n64280 );
and ( n64282 , n62081 , n64281 );
and ( n64283 , n62079 , n64282 );
and ( n64284 , n62077 , n64283 );
and ( n64285 , n62075 , n64284 );
and ( n64286 , n62073 , n64285 );
and ( n64287 , n62071 , n64286 );
and ( n64288 , n62069 , n64287 );
and ( n64289 , n62067 , n64288 );
and ( n64290 , n62065 , n64289 );
and ( n64291 , n62063 , n64290 );
and ( n64292 , n62061 , n64291 );
and ( n64293 , n62059 , n64292 );
and ( n64294 , n62057 , n64293 );
xor ( n64295 , n62055 , n64294 );
buf ( n64296 , n64295 );
xor ( n64297 , n62057 , n64293 );
buf ( n64298 , n64297 );
xor ( n64299 , n62059 , n64292 );
buf ( n64300 , n64299 );
xor ( n64301 , n62061 , n64291 );
buf ( n64302 , n64301 );
xor ( n64303 , n62063 , n64290 );
buf ( n64304 , n64303 );
xor ( n64305 , n62065 , n64289 );
buf ( n64306 , n64305 );
xor ( n64307 , n62067 , n64288 );
buf ( n64308 , n64307 );
xor ( n64309 , n62069 , n64287 );
buf ( n64310 , n64309 );
xor ( n64311 , n62071 , n64286 );
buf ( n64312 , n64311 );
xor ( n64313 , n62073 , n64285 );
buf ( n64314 , n64313 );
xor ( n64315 , n62075 , n64284 );
buf ( n64316 , n64315 );
xor ( n64317 , n62077 , n64283 );
buf ( n64318 , n64317 );
xor ( n64319 , n62079 , n64282 );
buf ( n64320 , n64319 );
xor ( n64321 , n62081 , n64281 );
buf ( n64322 , n64321 );
xor ( n64323 , n62083 , n64280 );
buf ( n64324 , n64323 );
xor ( n64325 , n62085 , n64279 );
buf ( n64326 , n64325 );
xor ( n64327 , n62087 , n64278 );
buf ( n64328 , n64327 );
xor ( n64329 , n62089 , n64277 );
buf ( n64330 , n64329 );
xor ( n64331 , n62091 , n64276 );
buf ( n64332 , n64331 );
xor ( n64333 , n62093 , n64275 );
buf ( n64334 , n64333 );
xor ( n64335 , n62095 , n64274 );
buf ( n64336 , n64335 );
xor ( n64337 , n62097 , n64273 );
buf ( n64338 , n64337 );
xor ( n64339 , n62099 , n64272 );
buf ( n64340 , n64339 );
xor ( n64341 , n62101 , n64271 );
buf ( n64342 , n64341 );
xor ( n64343 , n62103 , n64270 );
buf ( n64344 , n64343 );
xor ( n64345 , n62105 , n64269 );
buf ( n64346 , n64345 );
xor ( n64347 , n62107 , n64268 );
buf ( n64348 , n64347 );
xor ( n64349 , n62109 , n64267 );
buf ( n64350 , n64349 );
xor ( n64351 , n62111 , n64266 );
buf ( n64352 , n64351 );
xor ( n64353 , n62113 , n64265 );
buf ( n64354 , n64353 );
xor ( n64355 , n62115 , n64264 );
buf ( n64356 , n64355 );
xor ( n64357 , n62117 , n64263 );
buf ( n64358 , n64357 );
xor ( n64359 , n62119 , n64262 );
buf ( n64360 , n64359 );
xor ( n64361 , n62121 , n64261 );
buf ( n64362 , n64361 );
xor ( n64363 , n62123 , n64260 );
buf ( n64364 , n64363 );
xor ( n64365 , n62125 , n64259 );
buf ( n64366 , n64365 );
xor ( n64367 , n62127 , n64258 );
buf ( n64368 , n64367 );
xor ( n64369 , n62129 , n64257 );
buf ( n64370 , n64369 );
xor ( n64371 , n62131 , n64256 );
buf ( n64372 , n64371 );
xor ( n64373 , n62133 , n64255 );
buf ( n64374 , n64373 );
xor ( n64375 , n62135 , n64254 );
buf ( n64376 , n64375 );
xor ( n64377 , n62137 , n64253 );
buf ( n64378 , n64377 );
xor ( n64379 , n62139 , n64252 );
buf ( n64380 , n64379 );
xor ( n64381 , n62141 , n64251 );
buf ( n64382 , n64381 );
xor ( n64383 , n62143 , n64250 );
buf ( n64384 , n64383 );
xor ( n64385 , n62145 , n64249 );
buf ( n64386 , n64385 );
xor ( n64387 , n62147 , n64248 );
buf ( n64388 , n64387 );
xor ( n64389 , n62149 , n64247 );
buf ( n64390 , n64389 );
xor ( n64391 , n62151 , n64246 );
buf ( n64392 , n64391 );
xor ( n64393 , n62153 , n64245 );
buf ( n64394 , n64393 );
xor ( n64395 , n62155 , n64244 );
buf ( n64396 , n64395 );
xor ( n64397 , n62157 , n64243 );
buf ( n64398 , n64397 );
xor ( n64399 , n62159 , n64242 );
buf ( n64400 , n64399 );
xor ( n64401 , n62161 , n64241 );
buf ( n64402 , n64401 );
xor ( n64403 , n62163 , n64240 );
buf ( n64404 , n64403 );
xor ( n64405 , n62165 , n64239 );
buf ( n64406 , n64405 );
xor ( n64407 , n62167 , n64238 );
buf ( n64408 , n64407 );
xor ( n64409 , n62169 , n64237 );
buf ( n64410 , n64409 );
xor ( n64411 , n62171 , n64236 );
buf ( n64412 , n64411 );
xor ( n64413 , n62173 , n64235 );
buf ( n64414 , n64413 );
xor ( n64415 , n62175 , n64234 );
buf ( n64416 , n64415 );
xor ( n64417 , n62177 , n64233 );
buf ( n64418 , n64417 );
xor ( n64419 , n62179 , n64232 );
buf ( n64420 , n64419 );
xor ( n64421 , n62181 , n64231 );
buf ( n64422 , n64421 );
xor ( n64423 , n62183 , n64230 );
buf ( n64424 , n64423 );
xor ( n64425 , n62185 , n64229 );
buf ( n64426 , n64425 );
xor ( n64427 , n62290 , n64227 );
buf ( n64428 , n64427 );
xor ( n64429 , n62292 , n64226 );
buf ( n64430 , n64429 );
xor ( n64431 , n62294 , n64225 );
buf ( n64432 , n64431 );
xor ( n64433 , n62296 , n64224 );
buf ( n64434 , n64433 );
xor ( n64435 , n62683 , n64222 );
buf ( n64436 , n64435 );
xor ( n64437 , n62685 , n64221 );
buf ( n64438 , n64437 );
xor ( n64439 , n62816 , n64219 );
buf ( n64440 , n64439 );
xor ( n64441 , n62818 , n64218 );
buf ( n64442 , n64441 );
xor ( n64443 , n62820 , n64217 );
buf ( n64444 , n64443 );
xor ( n64445 , n62822 , n64216 );
buf ( n64446 , n64445 );
xor ( n64447 , n63044 , n64214 );
buf ( n64448 , n64447 );
xor ( n64449 , n63046 , n64213 );
buf ( n64450 , n64449 );
xor ( n64451 , n63245 , n64211 );
buf ( n64452 , n64451 );
xor ( n64453 , n63247 , n64210 );
buf ( n64454 , n64453 );
xor ( n64455 , n63343 , n64208 );
buf ( n64456 , n64455 );
xor ( n64457 , n63345 , n64207 );
buf ( n64458 , n64457 );
xor ( n64459 , n63433 , n64205 );
buf ( n64460 , n64459 );
xor ( n64461 , n63519 , n64203 );
buf ( n64462 , n64461 );
xor ( n64463 , n63588 , n64201 );
buf ( n64464 , n64463 );
xor ( n64465 , n63706 , n64199 );
buf ( n64466 , n64465 );
xor ( n64467 , n63708 , n64198 );
buf ( n64468 , n64467 );
xor ( n64469 , n63747 , n64196 );
buf ( n64470 , n64469 );
xor ( n64471 , n63875 , n64194 );
buf ( n64472 , n64471 );
xor ( n64473 , n63877 , n64193 );
buf ( n64474 , n64473 );
xor ( n64475 , n63956 , n64191 );
buf ( n64476 , n64475 );
xor ( n64477 , n64036 , n64189 );
buf ( n64478 , n64477 );
xor ( n64479 , n64038 , n64188 );
buf ( n64480 , n64479 );
xor ( n64481 , n64040 , n64187 );
buf ( n64482 , n64481 );
xor ( n64483 , n64046 , n64185 );
buf ( n64484 , n64483 );
xor ( n64485 , n64075 , n64183 );
buf ( n64486 , n64485 );
xor ( n64487 , n64104 , n64181 );
buf ( n64488 , n64487 );
xor ( n64489 , n64106 , n64180 );
buf ( n64490 , n64489 );
xor ( n64491 , n64122 , n64178 );
buf ( n64492 , n64491 );
xor ( n64493 , n64135 , n64176 );
buf ( n64494 , n64493 );
xor ( n64495 , n64147 , n64174 );
buf ( n64496 , n64495 );
xor ( n64497 , n64155 , n64172 );
buf ( n64498 , n64497 );
xor ( n64499 , n64160 , n64170 );
buf ( n64500 , n64499 );
xor ( n64501 , n64164 , n64168 );
buf ( n64502 , n64501 );
xor ( n64503 , n64166 , n64167 );
buf ( n64504 , n64503 );
buf ( n64505 , n55030 );
buf ( n64506 , n64505 );
buf ( n64507 , n30153 );
buf ( n64508 , n30156 );
buf ( n64509 , n30159 );
buf ( n64510 , n30162 );
buf ( n64511 , n30165 );
buf ( n64512 , n30168 );
buf ( n64513 , n30171 );
buf ( n64514 , n30174 );
buf ( n64515 , n30177 );
buf ( n64516 , n30180 );
buf ( n64517 , n30183 );
buf ( n64518 , n30186 );
buf ( n64519 , n30189 );
buf ( n64520 , n30192 );
buf ( n64521 , n30195 );
buf ( n64522 , n30198 );
buf ( n64523 , n30201 );
buf ( n64524 , n30204 );
buf ( n64525 , n30207 );
buf ( n64526 , n30210 );
buf ( n64527 , n30213 );
buf ( n64528 , n30216 );
buf ( n64529 , n30219 );
buf ( n64530 , n30222 );
buf ( n64531 , n30225 );
buf ( n64532 , n30228 );
buf ( n64533 , n30231 );
buf ( n64534 , n30234 );
buf ( n64535 , n30237 );
buf ( n64536 , n30240 );
buf ( n64537 , n30243 );
buf ( n64538 , n30246 );
buf ( n64539 , n30249 );
buf ( n64540 , n30252 );
buf ( n64541 , n30255 );
buf ( n64542 , n30258 );
buf ( n64543 , n30261 );
buf ( n64544 , n30264 );
buf ( n64545 , n30267 );
buf ( n64546 , n30270 );
buf ( n64547 , n30273 );
buf ( n64548 , n30276 );
buf ( n64549 , n30279 );
buf ( n64550 , n30282 );
buf ( n64551 , n30285 );
buf ( n64552 , n30288 );
buf ( n64553 , n30291 );
buf ( n64554 , n30294 );
buf ( n64555 , n30297 );
buf ( n64556 , n30300 );
buf ( n64557 , n30303 );
buf ( n64558 , n30306 );
buf ( n64559 , n30309 );
buf ( n64560 , n30312 );
buf ( n64561 , n30315 );
buf ( n64562 , n30318 );
buf ( n64563 , n30321 );
buf ( n64564 , n30324 );
buf ( n64565 , n30327 );
buf ( n64566 , n30330 );
buf ( n64567 , n30333 );
buf ( n64568 , n30336 );
buf ( n64569 , n30339 );
buf ( n64570 , n30342 );
buf ( n64571 , n30344 );
buf ( n64572 , n1186 );
buf ( n64573 , n1187 );
buf ( n64574 , n1188 );
buf ( n64575 , n1189 );
buf ( n64576 , n1190 );
buf ( n64577 , n1191 );
buf ( n64578 , n1192 );
buf ( n64579 , n1193 );
buf ( n64580 , n1194 );
buf ( n64581 , n1195 );
buf ( n64582 , n1196 );
buf ( n64583 , n1197 );
buf ( n64584 , n1198 );
buf ( n64585 , n1199 );
buf ( n64586 , n1200 );
buf ( n64587 , n1201 );
buf ( n64588 , n1202 );
buf ( n64589 , n1203 );
buf ( n64590 , n1204 );
buf ( n64591 , n1205 );
buf ( n64592 , n1206 );
buf ( n64593 , n1207 );
buf ( n64594 , n1208 );
buf ( n64595 , n1209 );
buf ( n64596 , n1210 );
buf ( n64597 , n1211 );
buf ( n64598 , n1212 );
buf ( n64599 , n1213 );
buf ( n64600 , n1214 );
buf ( n64601 , n1215 );
buf ( n64602 , n1216 );
buf ( n64603 , n1217 );
buf ( n64604 , n64574 );
buf ( n64605 , n64575 );
buf ( n64606 , n64576 );
and ( n64607 , n64605 , n64606 );
not ( n64608 , n64607 );
and ( n64609 , n64604 , n64608 );
not ( n64610 , n64609 );
buf ( n64611 , n64508 );
buf ( n64612 , n64572 );
buf ( n64613 , n64573 );
xor ( n64614 , n64612 , n64613 );
xor ( n64615 , n64613 , n64604 );
not ( n64616 , n64615 );
and ( n64617 , n64614 , n64616 );
and ( n64618 , n64611 , n64617 );
buf ( n64619 , n64507 );
and ( n64620 , n64619 , n64615 );
nor ( n64621 , n64618 , n64620 );
and ( n64622 , n64613 , n64604 );
not ( n64623 , n64622 );
and ( n64624 , n64612 , n64623 );
xnor ( n64625 , n64621 , n64624 );
and ( n64626 , n64610 , n64625 );
buf ( n64627 , n64509 );
and ( n64628 , n64627 , n64612 );
and ( n64629 , n64625 , n64628 );
and ( n64630 , n64610 , n64628 );
or ( n64631 , n64626 , n64629 , n64630 );
and ( n64632 , n64619 , n64617 );
not ( n64633 , n64632 );
xnor ( n64634 , n64633 , n64624 );
and ( n64635 , n64631 , n64634 );
and ( n64636 , n64611 , n64612 );
not ( n64637 , n64636 );
and ( n64638 , n64634 , n64637 );
and ( n64639 , n64631 , n64637 );
or ( n64640 , n64635 , n64638 , n64639 );
buf ( n64641 , n64636 );
not ( n64642 , n64624 );
xor ( n64643 , n64641 , n64642 );
and ( n64644 , n64619 , n64612 );
xor ( n64645 , n64643 , n64644 );
xor ( n64646 , n64640 , n64645 );
xor ( n64647 , n64631 , n64634 );
xor ( n64648 , n64647 , n64637 );
xor ( n64649 , n64604 , n64605 );
xor ( n64650 , n64605 , n64606 );
not ( n64651 , n64650 );
and ( n64652 , n64649 , n64651 );
and ( n64653 , n64619 , n64652 );
not ( n64654 , n64653 );
xnor ( n64655 , n64654 , n64609 );
not ( n64656 , n64655 );
and ( n64657 , n64627 , n64617 );
and ( n64658 , n64611 , n64615 );
nor ( n64659 , n64657 , n64658 );
xnor ( n64660 , n64659 , n64624 );
and ( n64661 , n64656 , n64660 );
buf ( n64662 , n64510 );
and ( n64663 , n64662 , n64612 );
and ( n64664 , n64660 , n64663 );
and ( n64665 , n64656 , n64663 );
or ( n64666 , n64661 , n64664 , n64665 );
buf ( n64667 , n64655 );
and ( n64668 , n64666 , n64667 );
xor ( n64669 , n64610 , n64625 );
xor ( n64670 , n64669 , n64628 );
and ( n64671 , n64667 , n64670 );
and ( n64672 , n64666 , n64670 );
or ( n64673 , n64668 , n64671 , n64672 );
and ( n64674 , n64648 , n64673 );
xor ( n64675 , n64648 , n64673 );
xor ( n64676 , n64666 , n64667 );
xor ( n64677 , n64676 , n64670 );
buf ( n64678 , n64577 );
buf ( n64679 , n64578 );
and ( n64680 , n64678 , n64679 );
not ( n64681 , n64680 );
and ( n64682 , n64606 , n64681 );
not ( n64683 , n64682 );
and ( n64684 , n64611 , n64652 );
and ( n64685 , n64619 , n64650 );
nor ( n64686 , n64684 , n64685 );
xnor ( n64687 , n64686 , n64609 );
and ( n64688 , n64683 , n64687 );
buf ( n64689 , n64511 );
and ( n64690 , n64689 , n64612 );
and ( n64691 , n64687 , n64690 );
and ( n64692 , n64683 , n64690 );
or ( n64693 , n64688 , n64691 , n64692 );
and ( n64694 , n64627 , n64652 );
and ( n64695 , n64611 , n64650 );
nor ( n64696 , n64694 , n64695 );
xnor ( n64697 , n64696 , n64609 );
and ( n64698 , n64689 , n64617 );
and ( n64699 , n64662 , n64615 );
nor ( n64700 , n64698 , n64699 );
xnor ( n64701 , n64700 , n64624 );
and ( n64702 , n64697 , n64701 );
buf ( n64703 , n64512 );
and ( n64704 , n64703 , n64612 );
and ( n64705 , n64701 , n64704 );
and ( n64706 , n64697 , n64704 );
or ( n64707 , n64702 , n64705 , n64706 );
xor ( n64708 , n64606 , n64678 );
xor ( n64709 , n64678 , n64679 );
not ( n64710 , n64709 );
and ( n64711 , n64708 , n64710 );
and ( n64712 , n64619 , n64711 );
not ( n64713 , n64712 );
xnor ( n64714 , n64713 , n64682 );
buf ( n64715 , n64714 );
and ( n64716 , n64707 , n64715 );
and ( n64717 , n64662 , n64617 );
and ( n64718 , n64627 , n64615 );
nor ( n64719 , n64717 , n64718 );
xnor ( n64720 , n64719 , n64624 );
and ( n64721 , n64715 , n64720 );
and ( n64722 , n64707 , n64720 );
or ( n64723 , n64716 , n64721 , n64722 );
and ( n64724 , n64693 , n64723 );
xor ( n64725 , n64656 , n64660 );
xor ( n64726 , n64725 , n64663 );
and ( n64727 , n64723 , n64726 );
and ( n64728 , n64693 , n64726 );
or ( n64729 , n64724 , n64727 , n64728 );
and ( n64730 , n64677 , n64729 );
xor ( n64731 , n64677 , n64729 );
xor ( n64732 , n64693 , n64723 );
xor ( n64733 , n64732 , n64726 );
buf ( n64734 , n64579 );
buf ( n64735 , n64580 );
and ( n64736 , n64734 , n64735 );
not ( n64737 , n64736 );
and ( n64738 , n64679 , n64737 );
not ( n64739 , n64738 );
and ( n64740 , n64611 , n64711 );
and ( n64741 , n64619 , n64709 );
nor ( n64742 , n64740 , n64741 );
xnor ( n64743 , n64742 , n64682 );
and ( n64744 , n64739 , n64743 );
and ( n64745 , n64703 , n64617 );
and ( n64746 , n64689 , n64615 );
nor ( n64747 , n64745 , n64746 );
xnor ( n64748 , n64747 , n64624 );
and ( n64749 , n64743 , n64748 );
and ( n64750 , n64739 , n64748 );
or ( n64751 , n64744 , n64749 , n64750 );
not ( n64752 , n64714 );
and ( n64753 , n64751 , n64752 );
xor ( n64754 , n64697 , n64701 );
xor ( n64755 , n64754 , n64704 );
and ( n64756 , n64752 , n64755 );
and ( n64757 , n64751 , n64755 );
or ( n64758 , n64753 , n64756 , n64757 );
xor ( n64759 , n64683 , n64687 );
xor ( n64760 , n64759 , n64690 );
and ( n64761 , n64758 , n64760 );
xor ( n64762 , n64707 , n64715 );
xor ( n64763 , n64762 , n64720 );
and ( n64764 , n64760 , n64763 );
and ( n64765 , n64758 , n64763 );
or ( n64766 , n64761 , n64764 , n64765 );
and ( n64767 , n64733 , n64766 );
xor ( n64768 , n64733 , n64766 );
xor ( n64769 , n64758 , n64760 );
xor ( n64770 , n64769 , n64763 );
and ( n64771 , n64627 , n64711 );
and ( n64772 , n64611 , n64709 );
nor ( n64773 , n64771 , n64772 );
xnor ( n64774 , n64773 , n64682 );
buf ( n64775 , n64774 );
and ( n64776 , n64662 , n64652 );
and ( n64777 , n64627 , n64650 );
nor ( n64778 , n64776 , n64777 );
xnor ( n64779 , n64778 , n64609 );
and ( n64780 , n64775 , n64779 );
buf ( n64781 , n64513 );
and ( n64782 , n64781 , n64612 );
and ( n64783 , n64779 , n64782 );
and ( n64784 , n64775 , n64782 );
or ( n64785 , n64780 , n64783 , n64784 );
xor ( n64786 , n64679 , n64734 );
xor ( n64787 , n64734 , n64735 );
not ( n64788 , n64787 );
and ( n64789 , n64786 , n64788 );
and ( n64790 , n64619 , n64789 );
not ( n64791 , n64790 );
xnor ( n64792 , n64791 , n64738 );
and ( n64793 , n64781 , n64617 );
and ( n64794 , n64703 , n64615 );
nor ( n64795 , n64793 , n64794 );
xnor ( n64796 , n64795 , n64624 );
and ( n64797 , n64792 , n64796 );
buf ( n64798 , n64514 );
and ( n64799 , n64798 , n64612 );
and ( n64800 , n64796 , n64799 );
and ( n64801 , n64792 , n64799 );
or ( n64802 , n64797 , n64800 , n64801 );
xor ( n64803 , n64739 , n64743 );
xor ( n64804 , n64803 , n64748 );
and ( n64805 , n64802 , n64804 );
xor ( n64806 , n64775 , n64779 );
xor ( n64807 , n64806 , n64782 );
and ( n64808 , n64804 , n64807 );
and ( n64809 , n64802 , n64807 );
or ( n64810 , n64805 , n64808 , n64809 );
and ( n64811 , n64785 , n64810 );
xor ( n64812 , n64751 , n64752 );
xor ( n64813 , n64812 , n64755 );
and ( n64814 , n64810 , n64813 );
and ( n64815 , n64785 , n64813 );
or ( n64816 , n64811 , n64814 , n64815 );
and ( n64817 , n64770 , n64816 );
xor ( n64818 , n64770 , n64816 );
xor ( n64819 , n64785 , n64810 );
xor ( n64820 , n64819 , n64813 );
and ( n64821 , n64662 , n64711 );
and ( n64822 , n64627 , n64709 );
nor ( n64823 , n64821 , n64822 );
xnor ( n64824 , n64823 , n64682 );
and ( n64825 , n64703 , n64652 );
and ( n64826 , n64689 , n64650 );
nor ( n64827 , n64825 , n64826 );
xnor ( n64828 , n64827 , n64609 );
and ( n64829 , n64824 , n64828 );
and ( n64830 , n64798 , n64617 );
and ( n64831 , n64781 , n64615 );
nor ( n64832 , n64830 , n64831 );
xnor ( n64833 , n64832 , n64624 );
and ( n64834 , n64828 , n64833 );
and ( n64835 , n64824 , n64833 );
or ( n64836 , n64829 , n64834 , n64835 );
not ( n64837 , n64774 );
and ( n64838 , n64836 , n64837 );
and ( n64839 , n64689 , n64652 );
and ( n64840 , n64662 , n64650 );
nor ( n64841 , n64839 , n64840 );
xnor ( n64842 , n64841 , n64609 );
and ( n64843 , n64837 , n64842 );
and ( n64844 , n64836 , n64842 );
or ( n64845 , n64838 , n64843 , n64844 );
buf ( n64846 , n64581 );
buf ( n64847 , n64582 );
and ( n64848 , n64846 , n64847 );
not ( n64849 , n64848 );
and ( n64850 , n64735 , n64849 );
not ( n64851 , n64850 );
and ( n64852 , n64611 , n64789 );
and ( n64853 , n64619 , n64787 );
nor ( n64854 , n64852 , n64853 );
xnor ( n64855 , n64854 , n64738 );
and ( n64856 , n64851 , n64855 );
buf ( n64857 , n64515 );
and ( n64858 , n64857 , n64612 );
and ( n64859 , n64855 , n64858 );
and ( n64860 , n64851 , n64858 );
or ( n64861 , n64856 , n64859 , n64860 );
xor ( n64862 , n64792 , n64796 );
xor ( n64863 , n64862 , n64799 );
and ( n64864 , n64861 , n64863 );
xor ( n64865 , n64836 , n64837 );
xor ( n64866 , n64865 , n64842 );
and ( n64867 , n64863 , n64866 );
and ( n64868 , n64861 , n64866 );
or ( n64869 , n64864 , n64867 , n64868 );
and ( n64870 , n64845 , n64869 );
xor ( n64871 , n64802 , n64804 );
xor ( n64872 , n64871 , n64807 );
and ( n64873 , n64869 , n64872 );
and ( n64874 , n64845 , n64872 );
or ( n64875 , n64870 , n64873 , n64874 );
and ( n64876 , n64820 , n64875 );
xor ( n64877 , n64820 , n64875 );
and ( n64878 , n64627 , n64789 );
and ( n64879 , n64611 , n64787 );
nor ( n64880 , n64878 , n64879 );
xnor ( n64881 , n64880 , n64738 );
and ( n64882 , n64781 , n64652 );
and ( n64883 , n64703 , n64650 );
nor ( n64884 , n64882 , n64883 );
xnor ( n64885 , n64884 , n64609 );
and ( n64886 , n64881 , n64885 );
and ( n64887 , n64857 , n64617 );
and ( n64888 , n64798 , n64615 );
nor ( n64889 , n64887 , n64888 );
xnor ( n64890 , n64889 , n64624 );
and ( n64891 , n64885 , n64890 );
and ( n64892 , n64881 , n64890 );
or ( n64893 , n64886 , n64891 , n64892 );
xor ( n64894 , n64735 , n64846 );
xor ( n64895 , n64846 , n64847 );
not ( n64896 , n64895 );
and ( n64897 , n64894 , n64896 );
and ( n64898 , n64619 , n64897 );
not ( n64899 , n64898 );
xnor ( n64900 , n64899 , n64850 );
and ( n64901 , n64689 , n64711 );
and ( n64902 , n64662 , n64709 );
nor ( n64903 , n64901 , n64902 );
xnor ( n64904 , n64903 , n64682 );
and ( n64905 , n64900 , n64904 );
buf ( n64906 , n64516 );
and ( n64907 , n64906 , n64612 );
not ( n64908 , n64907 );
and ( n64909 , n64904 , n64908 );
and ( n64910 , n64900 , n64908 );
or ( n64911 , n64905 , n64909 , n64910 );
and ( n64912 , n64893 , n64911 );
buf ( n64913 , n64907 );
and ( n64914 , n64911 , n64913 );
and ( n64915 , n64893 , n64913 );
or ( n64916 , n64912 , n64914 , n64915 );
xor ( n64917 , n64851 , n64855 );
xor ( n64918 , n64917 , n64858 );
xor ( n64919 , n64824 , n64828 );
xor ( n64920 , n64919 , n64833 );
and ( n64921 , n64918 , n64920 );
xor ( n64922 , n64893 , n64911 );
xor ( n64923 , n64922 , n64913 );
and ( n64924 , n64920 , n64923 );
and ( n64925 , n64918 , n64923 );
or ( n64926 , n64921 , n64924 , n64925 );
and ( n64927 , n64916 , n64926 );
xor ( n64928 , n64861 , n64863 );
xor ( n64929 , n64928 , n64866 );
and ( n64930 , n64926 , n64929 );
and ( n64931 , n64916 , n64929 );
or ( n64932 , n64927 , n64930 , n64931 );
xor ( n64933 , n64845 , n64869 );
xor ( n64934 , n64933 , n64872 );
and ( n64935 , n64932 , n64934 );
xor ( n64936 , n64932 , n64934 );
xor ( n64937 , n64916 , n64926 );
xor ( n64938 , n64937 , n64929 );
buf ( n64939 , n64583 );
buf ( n64940 , n64584 );
and ( n64941 , n64939 , n64940 );
not ( n64942 , n64941 );
and ( n64943 , n64847 , n64942 );
not ( n64944 , n64943 );
and ( n64945 , n64906 , n64617 );
and ( n64946 , n64857 , n64615 );
nor ( n64947 , n64945 , n64946 );
xnor ( n64948 , n64947 , n64624 );
and ( n64949 , n64944 , n64948 );
buf ( n64950 , n64517 );
and ( n64951 , n64950 , n64612 );
and ( n64952 , n64948 , n64951 );
and ( n64953 , n64944 , n64951 );
or ( n64954 , n64949 , n64952 , n64953 );
buf ( n64955 , n64518 );
and ( n64956 , n64955 , n64612 );
buf ( n64957 , n64956 );
and ( n64958 , n64611 , n64897 );
and ( n64959 , n64619 , n64895 );
nor ( n64960 , n64958 , n64959 );
xnor ( n64961 , n64960 , n64850 );
and ( n64962 , n64957 , n64961 );
and ( n64963 , n64703 , n64711 );
and ( n64964 , n64689 , n64709 );
nor ( n64965 , n64963 , n64964 );
xnor ( n64966 , n64965 , n64682 );
and ( n64967 , n64961 , n64966 );
and ( n64968 , n64957 , n64966 );
or ( n64969 , n64962 , n64967 , n64968 );
and ( n64970 , n64954 , n64969 );
xor ( n64971 , n64900 , n64904 );
xor ( n64972 , n64971 , n64908 );
and ( n64973 , n64969 , n64972 );
and ( n64974 , n64954 , n64972 );
or ( n64975 , n64970 , n64973 , n64974 );
and ( n64976 , n64662 , n64789 );
and ( n64977 , n64627 , n64787 );
nor ( n64978 , n64976 , n64977 );
xnor ( n64979 , n64978 , n64738 );
and ( n64980 , n64798 , n64652 );
and ( n64981 , n64781 , n64650 );
nor ( n64982 , n64980 , n64981 );
xnor ( n64983 , n64982 , n64609 );
and ( n64984 , n64979 , n64983 );
xor ( n64985 , n64944 , n64948 );
xor ( n64986 , n64985 , n64951 );
and ( n64987 , n64983 , n64986 );
and ( n64988 , n64979 , n64986 );
or ( n64989 , n64984 , n64987 , n64988 );
buf ( n64990 , n64585 );
buf ( n64991 , n64586 );
and ( n64992 , n64990 , n64991 );
not ( n64993 , n64992 );
and ( n64994 , n64940 , n64993 );
not ( n64995 , n64994 );
and ( n64996 , n64955 , n64617 );
and ( n64997 , n64950 , n64615 );
nor ( n64998 , n64996 , n64997 );
xnor ( n64999 , n64998 , n64624 );
and ( n65000 , n64995 , n64999 );
buf ( n65001 , n64519 );
and ( n65002 , n65001 , n64612 );
and ( n65003 , n64999 , n65002 );
and ( n65004 , n64995 , n65002 );
or ( n65005 , n65000 , n65003 , n65004 );
and ( n65006 , n64781 , n64711 );
and ( n65007 , n64703 , n64709 );
nor ( n65008 , n65006 , n65007 );
xnor ( n65009 , n65008 , n64682 );
and ( n65010 , n65005 , n65009 );
and ( n65011 , n64857 , n64652 );
and ( n65012 , n64798 , n64650 );
nor ( n65013 , n65011 , n65012 );
xnor ( n65014 , n65013 , n64609 );
and ( n65015 , n65009 , n65014 );
and ( n65016 , n65005 , n65014 );
or ( n65017 , n65010 , n65015 , n65016 );
and ( n65018 , n64627 , n64897 );
and ( n65019 , n64611 , n64895 );
nor ( n65020 , n65018 , n65019 );
xnor ( n65021 , n65020 , n64850 );
and ( n65022 , n64950 , n64617 );
and ( n65023 , n64906 , n64615 );
nor ( n65024 , n65022 , n65023 );
xnor ( n65025 , n65024 , n64624 );
and ( n65026 , n65021 , n65025 );
not ( n65027 , n64956 );
and ( n65028 , n65025 , n65027 );
and ( n65029 , n65021 , n65027 );
or ( n65030 , n65026 , n65028 , n65029 );
and ( n65031 , n65017 , n65030 );
xor ( n65032 , n64979 , n64983 );
xor ( n65033 , n65032 , n64986 );
and ( n65034 , n65030 , n65033 );
and ( n65035 , n65017 , n65033 );
or ( n65036 , n65031 , n65034 , n65035 );
and ( n65037 , n64989 , n65036 );
xor ( n65038 , n64881 , n64885 );
xor ( n65039 , n65038 , n64890 );
and ( n65040 , n65036 , n65039 );
and ( n65041 , n64989 , n65039 );
or ( n65042 , n65037 , n65040 , n65041 );
and ( n65043 , n64975 , n65042 );
xor ( n65044 , n64918 , n64920 );
xor ( n65045 , n65044 , n64923 );
and ( n65046 , n65042 , n65045 );
and ( n65047 , n64975 , n65045 );
or ( n65048 , n65043 , n65046 , n65047 );
and ( n65049 , n64938 , n65048 );
xor ( n65050 , n64938 , n65048 );
xor ( n65051 , n64975 , n65042 );
xor ( n65052 , n65051 , n65045 );
xor ( n65053 , n64847 , n64939 );
xor ( n65054 , n64939 , n64940 );
not ( n65055 , n65054 );
and ( n65056 , n65053 , n65055 );
and ( n65057 , n64611 , n65056 );
and ( n65058 , n64619 , n65054 );
nor ( n65059 , n65057 , n65058 );
xnor ( n65060 , n65059 , n64943 );
and ( n65061 , n64662 , n64897 );
and ( n65062 , n64627 , n64895 );
nor ( n65063 , n65061 , n65062 );
xnor ( n65064 , n65063 , n64850 );
and ( n65065 , n65060 , n65064 );
and ( n65066 , n64798 , n64711 );
and ( n65067 , n64781 , n64709 );
nor ( n65068 , n65066 , n65067 );
xnor ( n65069 , n65068 , n64682 );
and ( n65070 , n65064 , n65069 );
and ( n65071 , n65060 , n65069 );
or ( n65072 , n65065 , n65070 , n65071 );
and ( n65073 , n64619 , n65056 );
not ( n65074 , n65073 );
xnor ( n65075 , n65074 , n64943 );
and ( n65076 , n65072 , n65075 );
and ( n65077 , n64689 , n64789 );
and ( n65078 , n64662 , n64787 );
nor ( n65079 , n65077 , n65078 );
xnor ( n65080 , n65079 , n64738 );
and ( n65081 , n65075 , n65080 );
and ( n65082 , n65072 , n65080 );
or ( n65083 , n65076 , n65081 , n65082 );
xor ( n65084 , n64957 , n64961 );
xor ( n65085 , n65084 , n64966 );
and ( n65086 , n65083 , n65085 );
xor ( n65087 , n65017 , n65030 );
xor ( n65088 , n65087 , n65033 );
and ( n65089 , n65085 , n65088 );
and ( n65090 , n65083 , n65088 );
or ( n65091 , n65086 , n65089 , n65090 );
xor ( n65092 , n64954 , n64969 );
xor ( n65093 , n65092 , n64972 );
and ( n65094 , n65091 , n65093 );
xor ( n65095 , n64989 , n65036 );
xor ( n65096 , n65095 , n65039 );
and ( n65097 , n65093 , n65096 );
and ( n65098 , n65091 , n65096 );
or ( n65099 , n65094 , n65097 , n65098 );
and ( n65100 , n65052 , n65099 );
xor ( n65101 , n65052 , n65099 );
xor ( n65102 , n65091 , n65093 );
xor ( n65103 , n65102 , n65096 );
and ( n65104 , n65001 , n64617 );
and ( n65105 , n64955 , n64615 );
nor ( n65106 , n65104 , n65105 );
xnor ( n65107 , n65106 , n64624 );
buf ( n65108 , n65107 );
and ( n65109 , n64703 , n64789 );
and ( n65110 , n64689 , n64787 );
nor ( n65111 , n65109 , n65110 );
xnor ( n65112 , n65111 , n64738 );
and ( n65113 , n65108 , n65112 );
and ( n65114 , n64906 , n64652 );
and ( n65115 , n64857 , n64650 );
nor ( n65116 , n65114 , n65115 );
xnor ( n65117 , n65116 , n64609 );
and ( n65118 , n65112 , n65117 );
and ( n65119 , n65108 , n65117 );
or ( n65120 , n65113 , n65118 , n65119 );
xor ( n65121 , n65005 , n65009 );
xor ( n65122 , n65121 , n65014 );
and ( n65123 , n65120 , n65122 );
xor ( n65124 , n65021 , n65025 );
xor ( n65125 , n65124 , n65027 );
and ( n65126 , n65122 , n65125 );
and ( n65127 , n65120 , n65125 );
or ( n65128 , n65123 , n65126 , n65127 );
and ( n65129 , n64950 , n64652 );
and ( n65130 , n64906 , n64650 );
nor ( n65131 , n65129 , n65130 );
xnor ( n65132 , n65131 , n64609 );
not ( n65133 , n65107 );
and ( n65134 , n65132 , n65133 );
buf ( n65135 , n64520 );
and ( n65136 , n65135 , n64612 );
and ( n65137 , n65133 , n65136 );
and ( n65138 , n65132 , n65136 );
or ( n65139 , n65134 , n65137 , n65138 );
xor ( n65140 , n64995 , n64999 );
xor ( n65141 , n65140 , n65002 );
and ( n65142 , n65139 , n65141 );
xor ( n65143 , n65108 , n65112 );
xor ( n65144 , n65143 , n65117 );
and ( n65145 , n65141 , n65144 );
and ( n65146 , n65139 , n65144 );
or ( n65147 , n65142 , n65145 , n65146 );
and ( n65148 , n64627 , n65056 );
and ( n65149 , n64611 , n65054 );
nor ( n65150 , n65148 , n65149 );
xnor ( n65151 , n65150 , n64943 );
and ( n65152 , n64781 , n64789 );
and ( n65153 , n64703 , n64787 );
nor ( n65154 , n65152 , n65153 );
xnor ( n65155 , n65154 , n64738 );
and ( n65156 , n65151 , n65155 );
and ( n65157 , n64857 , n64711 );
and ( n65158 , n64798 , n64709 );
nor ( n65159 , n65157 , n65158 );
xnor ( n65160 , n65159 , n64682 );
and ( n65161 , n65155 , n65160 );
and ( n65162 , n65151 , n65160 );
or ( n65163 , n65156 , n65161 , n65162 );
buf ( n65164 , n64587 );
buf ( n65165 , n64588 );
and ( n65166 , n65164 , n65165 );
not ( n65167 , n65166 );
and ( n65168 , n64991 , n65167 );
not ( n65169 , n65168 );
and ( n65170 , n65135 , n64617 );
and ( n65171 , n65001 , n64615 );
nor ( n65172 , n65170 , n65171 );
xnor ( n65173 , n65172 , n64624 );
and ( n65174 , n65169 , n65173 );
buf ( n65175 , n64521 );
and ( n65176 , n65175 , n64612 );
and ( n65177 , n65173 , n65176 );
and ( n65178 , n65169 , n65176 );
or ( n65179 , n65174 , n65177 , n65178 );
xor ( n65180 , n64940 , n64990 );
xor ( n65181 , n64990 , n64991 );
not ( n65182 , n65181 );
and ( n65183 , n65180 , n65182 );
and ( n65184 , n64619 , n65183 );
not ( n65185 , n65184 );
xnor ( n65186 , n65185 , n64994 );
and ( n65187 , n65179 , n65186 );
and ( n65188 , n64689 , n64897 );
and ( n65189 , n64662 , n64895 );
nor ( n65190 , n65188 , n65189 );
xnor ( n65191 , n65190 , n64850 );
and ( n65192 , n65186 , n65191 );
and ( n65193 , n65179 , n65191 );
or ( n65194 , n65187 , n65192 , n65193 );
and ( n65195 , n65163 , n65194 );
xor ( n65196 , n65060 , n65064 );
xor ( n65197 , n65196 , n65069 );
and ( n65198 , n65194 , n65197 );
and ( n65199 , n65163 , n65197 );
or ( n65200 , n65195 , n65198 , n65199 );
and ( n65201 , n65147 , n65200 );
xor ( n65202 , n65072 , n65075 );
xor ( n65203 , n65202 , n65080 );
and ( n65204 , n65200 , n65203 );
and ( n65205 , n65147 , n65203 );
or ( n65206 , n65201 , n65204 , n65205 );
and ( n65207 , n65128 , n65206 );
xor ( n65208 , n65083 , n65085 );
xor ( n65209 , n65208 , n65088 );
and ( n65210 , n65206 , n65209 );
and ( n65211 , n65128 , n65209 );
or ( n65212 , n65207 , n65210 , n65211 );
and ( n65213 , n65103 , n65212 );
xor ( n65214 , n65103 , n65212 );
xor ( n65215 , n65128 , n65206 );
xor ( n65216 , n65215 , n65209 );
and ( n65217 , n64611 , n65183 );
and ( n65218 , n64619 , n65181 );
nor ( n65219 , n65217 , n65218 );
xnor ( n65220 , n65219 , n64994 );
and ( n65221 , n64703 , n64897 );
and ( n65222 , n64689 , n64895 );
nor ( n65223 , n65221 , n65222 );
xnor ( n65224 , n65223 , n64850 );
and ( n65225 , n65220 , n65224 );
and ( n65226 , n64798 , n64789 );
and ( n65227 , n64781 , n64787 );
nor ( n65228 , n65226 , n65227 );
xnor ( n65229 , n65228 , n64738 );
and ( n65230 , n65224 , n65229 );
and ( n65231 , n65220 , n65229 );
or ( n65232 , n65225 , n65230 , n65231 );
and ( n65233 , n65001 , n64652 );
and ( n65234 , n64955 , n64650 );
nor ( n65235 , n65233 , n65234 );
xnor ( n65236 , n65235 , n64609 );
buf ( n65237 , n65236 );
and ( n65238 , n64906 , n64711 );
and ( n65239 , n64857 , n64709 );
nor ( n65240 , n65238 , n65239 );
xnor ( n65241 , n65240 , n64682 );
and ( n65242 , n65237 , n65241 );
and ( n65243 , n64955 , n64652 );
and ( n65244 , n64950 , n64650 );
nor ( n65245 , n65243 , n65244 );
xnor ( n65246 , n65245 , n64609 );
and ( n65247 , n65241 , n65246 );
and ( n65248 , n65237 , n65246 );
or ( n65249 , n65242 , n65247 , n65248 );
and ( n65250 , n65232 , n65249 );
xor ( n65251 , n65132 , n65133 );
xor ( n65252 , n65251 , n65136 );
and ( n65253 , n65249 , n65252 );
and ( n65254 , n65232 , n65252 );
or ( n65255 , n65250 , n65253 , n65254 );
and ( n65256 , n64950 , n64711 );
and ( n65257 , n64906 , n64709 );
nor ( n65258 , n65256 , n65257 );
xnor ( n65259 , n65258 , n64682 );
and ( n65260 , n65175 , n64617 );
and ( n65261 , n65135 , n64615 );
nor ( n65262 , n65260 , n65261 );
xnor ( n65263 , n65262 , n64624 );
and ( n65264 , n65259 , n65263 );
buf ( n65265 , n64522 );
and ( n65266 , n65265 , n64612 );
and ( n65267 , n65263 , n65266 );
and ( n65268 , n65259 , n65266 );
or ( n65269 , n65264 , n65267 , n65268 );
and ( n65270 , n64662 , n65056 );
and ( n65271 , n64627 , n65054 );
nor ( n65272 , n65270 , n65271 );
xnor ( n65273 , n65272 , n64943 );
and ( n65274 , n65269 , n65273 );
xor ( n65275 , n65169 , n65173 );
xor ( n65276 , n65275 , n65176 );
and ( n65277 , n65273 , n65276 );
and ( n65278 , n65269 , n65276 );
or ( n65279 , n65274 , n65277 , n65278 );
xor ( n65280 , n65151 , n65155 );
xor ( n65281 , n65280 , n65160 );
and ( n65282 , n65279 , n65281 );
xor ( n65283 , n65179 , n65186 );
xor ( n65284 , n65283 , n65191 );
and ( n65285 , n65281 , n65284 );
and ( n65286 , n65279 , n65284 );
or ( n65287 , n65282 , n65285 , n65286 );
and ( n65288 , n65255 , n65287 );
xor ( n65289 , n65139 , n65141 );
xor ( n65290 , n65289 , n65144 );
and ( n65291 , n65287 , n65290 );
and ( n65292 , n65255 , n65290 );
or ( n65293 , n65288 , n65291 , n65292 );
xor ( n65294 , n65120 , n65122 );
xor ( n65295 , n65294 , n65125 );
and ( n65296 , n65293 , n65295 );
xor ( n65297 , n65147 , n65200 );
xor ( n65298 , n65297 , n65203 );
and ( n65299 , n65295 , n65298 );
and ( n65300 , n65293 , n65298 );
or ( n65301 , n65296 , n65299 , n65300 );
and ( n65302 , n65216 , n65301 );
xor ( n65303 , n65216 , n65301 );
xor ( n65304 , n65293 , n65295 );
xor ( n65305 , n65304 , n65298 );
buf ( n65306 , n64524 );
and ( n65307 , n65306 , n64612 );
buf ( n65308 , n65307 );
buf ( n65309 , n64589 );
buf ( n65310 , n64590 );
and ( n65311 , n65309 , n65310 );
not ( n65312 , n65311 );
and ( n65313 , n65165 , n65312 );
not ( n65314 , n65313 );
and ( n65315 , n65308 , n65314 );
and ( n65316 , n65265 , n64617 );
and ( n65317 , n65175 , n64615 );
nor ( n65318 , n65316 , n65317 );
xnor ( n65319 , n65318 , n64624 );
and ( n65320 , n65314 , n65319 );
and ( n65321 , n65308 , n65319 );
or ( n65322 , n65315 , n65320 , n65321 );
and ( n65323 , n64689 , n65056 );
and ( n65324 , n64662 , n65054 );
nor ( n65325 , n65323 , n65324 );
xnor ( n65326 , n65325 , n64943 );
and ( n65327 , n65322 , n65326 );
and ( n65328 , n64857 , n64789 );
and ( n65329 , n64798 , n64787 );
nor ( n65330 , n65328 , n65329 );
xnor ( n65331 , n65330 , n64738 );
and ( n65332 , n65326 , n65331 );
and ( n65333 , n65322 , n65331 );
or ( n65334 , n65327 , n65332 , n65333 );
and ( n65335 , n64627 , n65183 );
and ( n65336 , n64611 , n65181 );
nor ( n65337 , n65335 , n65336 );
xnor ( n65338 , n65337 , n64994 );
and ( n65339 , n64781 , n64897 );
and ( n65340 , n64703 , n64895 );
nor ( n65341 , n65339 , n65340 );
xnor ( n65342 , n65341 , n64850 );
and ( n65343 , n65338 , n65342 );
not ( n65344 , n65236 );
and ( n65345 , n65342 , n65344 );
and ( n65346 , n65338 , n65344 );
or ( n65347 , n65343 , n65345 , n65346 );
and ( n65348 , n65334 , n65347 );
xor ( n65349 , n65237 , n65241 );
xor ( n65350 , n65349 , n65246 );
and ( n65351 , n65347 , n65350 );
and ( n65352 , n65334 , n65350 );
or ( n65353 , n65348 , n65351 , n65352 );
and ( n65354 , n64955 , n64711 );
and ( n65355 , n64950 , n64709 );
nor ( n65356 , n65354 , n65355 );
xnor ( n65357 , n65356 , n64682 );
and ( n65358 , n65135 , n64652 );
and ( n65359 , n65001 , n64650 );
nor ( n65360 , n65358 , n65359 );
xnor ( n65361 , n65360 , n64609 );
and ( n65362 , n65357 , n65361 );
buf ( n65363 , n64523 );
and ( n65364 , n65363 , n64612 );
and ( n65365 , n65361 , n65364 );
and ( n65366 , n65357 , n65364 );
or ( n65367 , n65362 , n65365 , n65366 );
xor ( n65368 , n64991 , n65164 );
xor ( n65369 , n65164 , n65165 );
not ( n65370 , n65369 );
and ( n65371 , n65368 , n65370 );
and ( n65372 , n64619 , n65371 );
not ( n65373 , n65372 );
xnor ( n65374 , n65373 , n65168 );
and ( n65375 , n65367 , n65374 );
xor ( n65376 , n65259 , n65263 );
xor ( n65377 , n65376 , n65266 );
and ( n65378 , n65374 , n65377 );
and ( n65379 , n65367 , n65377 );
or ( n65380 , n65375 , n65378 , n65379 );
xor ( n65381 , n65220 , n65224 );
xor ( n65382 , n65381 , n65229 );
and ( n65383 , n65380 , n65382 );
xor ( n65384 , n65269 , n65273 );
xor ( n65385 , n65384 , n65276 );
and ( n65386 , n65382 , n65385 );
and ( n65387 , n65380 , n65385 );
or ( n65388 , n65383 , n65386 , n65387 );
and ( n65389 , n65353 , n65388 );
xor ( n65390 , n65232 , n65249 );
xor ( n65391 , n65390 , n65252 );
and ( n65392 , n65388 , n65391 );
and ( n65393 , n65353 , n65391 );
or ( n65394 , n65389 , n65392 , n65393 );
xor ( n65395 , n65163 , n65194 );
xor ( n65396 , n65395 , n65197 );
and ( n65397 , n65394 , n65396 );
xor ( n65398 , n65255 , n65287 );
xor ( n65399 , n65398 , n65290 );
and ( n65400 , n65396 , n65399 );
and ( n65401 , n65394 , n65399 );
or ( n65402 , n65397 , n65400 , n65401 );
and ( n65403 , n65305 , n65402 );
xor ( n65404 , n65305 , n65402 );
xor ( n65405 , n65394 , n65396 );
xor ( n65406 , n65405 , n65399 );
and ( n65407 , n64611 , n65371 );
and ( n65408 , n64619 , n65369 );
nor ( n65409 , n65407 , n65408 );
xnor ( n65410 , n65409 , n65168 );
and ( n65411 , n64662 , n65183 );
and ( n65412 , n64627 , n65181 );
nor ( n65413 , n65411 , n65412 );
xnor ( n65414 , n65413 , n64994 );
and ( n65415 , n65410 , n65414 );
and ( n65416 , n64798 , n64897 );
and ( n65417 , n64781 , n64895 );
nor ( n65418 , n65416 , n65417 );
xnor ( n65419 , n65418 , n64850 );
and ( n65420 , n65414 , n65419 );
and ( n65421 , n65410 , n65419 );
or ( n65422 , n65415 , n65420 , n65421 );
and ( n65423 , n64703 , n65056 );
and ( n65424 , n64689 , n65054 );
nor ( n65425 , n65423 , n65424 );
xnor ( n65426 , n65425 , n64943 );
and ( n65427 , n64906 , n64789 );
and ( n65428 , n64857 , n64787 );
nor ( n65429 , n65427 , n65428 );
xnor ( n65430 , n65429 , n64738 );
and ( n65431 , n65426 , n65430 );
xor ( n65432 , n65308 , n65314 );
xor ( n65433 , n65432 , n65319 );
and ( n65434 , n65430 , n65433 );
and ( n65435 , n65426 , n65433 );
or ( n65436 , n65431 , n65434 , n65435 );
and ( n65437 , n65422 , n65436 );
xor ( n65438 , n65338 , n65342 );
xor ( n65439 , n65438 , n65344 );
and ( n65440 , n65436 , n65439 );
and ( n65441 , n65422 , n65439 );
or ( n65442 , n65437 , n65440 , n65441 );
buf ( n65443 , n64526 );
and ( n65444 , n65443 , n64612 );
buf ( n65445 , n65444 );
buf ( n65446 , n64591 );
buf ( n65447 , n64592 );
and ( n65448 , n65446 , n65447 );
not ( n65449 , n65448 );
and ( n65450 , n65310 , n65449 );
not ( n65451 , n65450 );
and ( n65452 , n65445 , n65451 );
buf ( n65453 , n64525 );
and ( n65454 , n65453 , n64612 );
and ( n65455 , n65451 , n65454 );
and ( n65456 , n65445 , n65454 );
or ( n65457 , n65452 , n65455 , n65456 );
and ( n65458 , n64950 , n64789 );
and ( n65459 , n64906 , n64787 );
nor ( n65460 , n65458 , n65459 );
xnor ( n65461 , n65460 , n64738 );
and ( n65462 , n65457 , n65461 );
and ( n65463 , n65175 , n64652 );
and ( n65464 , n65135 , n64650 );
nor ( n65465 , n65463 , n65464 );
xnor ( n65466 , n65465 , n64609 );
and ( n65467 , n65461 , n65466 );
and ( n65468 , n65457 , n65466 );
or ( n65469 , n65462 , n65467 , n65468 );
and ( n65470 , n65001 , n64711 );
and ( n65471 , n64955 , n64709 );
nor ( n65472 , n65470 , n65471 );
xnor ( n65473 , n65472 , n64682 );
and ( n65474 , n65363 , n64617 );
and ( n65475 , n65265 , n64615 );
nor ( n65476 , n65474 , n65475 );
xnor ( n65477 , n65476 , n64624 );
and ( n65478 , n65473 , n65477 );
not ( n65479 , n65307 );
and ( n65480 , n65477 , n65479 );
and ( n65481 , n65473 , n65479 );
or ( n65482 , n65478 , n65480 , n65481 );
and ( n65483 , n65469 , n65482 );
xor ( n65484 , n65357 , n65361 );
xor ( n65485 , n65484 , n65364 );
and ( n65486 , n65482 , n65485 );
and ( n65487 , n65469 , n65485 );
or ( n65488 , n65483 , n65486 , n65487 );
xor ( n65489 , n65322 , n65326 );
xor ( n65490 , n65489 , n65331 );
and ( n65491 , n65488 , n65490 );
xor ( n65492 , n65367 , n65374 );
xor ( n65493 , n65492 , n65377 );
and ( n65494 , n65490 , n65493 );
and ( n65495 , n65488 , n65493 );
or ( n65496 , n65491 , n65494 , n65495 );
and ( n65497 , n65442 , n65496 );
xor ( n65498 , n65334 , n65347 );
xor ( n65499 , n65498 , n65350 );
and ( n65500 , n65496 , n65499 );
and ( n65501 , n65442 , n65499 );
or ( n65502 , n65497 , n65500 , n65501 );
xor ( n65503 , n65279 , n65281 );
xor ( n65504 , n65503 , n65284 );
and ( n65505 , n65502 , n65504 );
xor ( n65506 , n65353 , n65388 );
xor ( n65507 , n65506 , n65391 );
and ( n65508 , n65504 , n65507 );
and ( n65509 , n65502 , n65507 );
or ( n65510 , n65505 , n65508 , n65509 );
and ( n65511 , n65406 , n65510 );
xor ( n65512 , n65406 , n65510 );
xor ( n65513 , n65502 , n65504 );
xor ( n65514 , n65513 , n65507 );
and ( n65515 , n64627 , n65371 );
and ( n65516 , n64611 , n65369 );
nor ( n65517 , n65515 , n65516 );
xnor ( n65518 , n65517 , n65168 );
and ( n65519 , n64781 , n65056 );
and ( n65520 , n64703 , n65054 );
nor ( n65521 , n65519 , n65520 );
xnor ( n65522 , n65521 , n64943 );
and ( n65523 , n65518 , n65522 );
and ( n65524 , n64857 , n64897 );
and ( n65525 , n64798 , n64895 );
nor ( n65526 , n65524 , n65525 );
xnor ( n65527 , n65526 , n64850 );
and ( n65528 , n65522 , n65527 );
and ( n65529 , n65518 , n65527 );
or ( n65530 , n65523 , n65528 , n65529 );
and ( n65531 , n65135 , n64711 );
and ( n65532 , n65001 , n64709 );
nor ( n65533 , n65531 , n65532 );
xnor ( n65534 , n65533 , n64682 );
and ( n65535 , n65265 , n64652 );
and ( n65536 , n65175 , n64650 );
nor ( n65537 , n65535 , n65536 );
xnor ( n65538 , n65537 , n64609 );
and ( n65539 , n65534 , n65538 );
and ( n65540 , n65306 , n64617 );
and ( n65541 , n65363 , n64615 );
nor ( n65542 , n65540 , n65541 );
xnor ( n65543 , n65542 , n64624 );
and ( n65544 , n65538 , n65543 );
and ( n65545 , n65534 , n65543 );
or ( n65546 , n65539 , n65544 , n65545 );
xor ( n65547 , n65165 , n65309 );
xor ( n65548 , n65309 , n65310 );
not ( n65549 , n65548 );
and ( n65550 , n65547 , n65549 );
and ( n65551 , n64619 , n65550 );
not ( n65552 , n65551 );
xnor ( n65553 , n65552 , n65313 );
and ( n65554 , n65546 , n65553 );
and ( n65555 , n64689 , n65183 );
and ( n65556 , n64662 , n65181 );
nor ( n65557 , n65555 , n65556 );
xnor ( n65558 , n65557 , n64994 );
and ( n65559 , n65553 , n65558 );
and ( n65560 , n65546 , n65558 );
or ( n65561 , n65554 , n65559 , n65560 );
and ( n65562 , n65530 , n65561 );
xor ( n65563 , n65426 , n65430 );
xor ( n65564 , n65563 , n65433 );
and ( n65565 , n65561 , n65564 );
and ( n65566 , n65530 , n65564 );
or ( n65567 , n65562 , n65565 , n65566 );
xor ( n65568 , n65422 , n65436 );
xor ( n65569 , n65568 , n65439 );
and ( n65570 , n65567 , n65569 );
xor ( n65571 , n65488 , n65490 );
xor ( n65572 , n65571 , n65493 );
and ( n65573 , n65569 , n65572 );
and ( n65574 , n65567 , n65572 );
or ( n65575 , n65570 , n65573 , n65574 );
xor ( n65576 , n65380 , n65382 );
xor ( n65577 , n65576 , n65385 );
and ( n65578 , n65575 , n65577 );
xor ( n65579 , n65442 , n65496 );
xor ( n65580 , n65579 , n65499 );
and ( n65581 , n65577 , n65580 );
and ( n65582 , n65575 , n65580 );
or ( n65583 , n65578 , n65581 , n65582 );
and ( n65584 , n65514 , n65583 );
xor ( n65585 , n65514 , n65583 );
xor ( n65586 , n65575 , n65577 );
xor ( n65587 , n65586 , n65580 );
and ( n65588 , n64906 , n64897 );
and ( n65589 , n64857 , n64895 );
nor ( n65590 , n65588 , n65589 );
xnor ( n65591 , n65590 , n64850 );
and ( n65592 , n64955 , n64789 );
and ( n65593 , n64950 , n64787 );
nor ( n65594 , n65592 , n65593 );
xnor ( n65595 , n65594 , n64738 );
and ( n65596 , n65591 , n65595 );
xor ( n65597 , n65445 , n65451 );
xor ( n65598 , n65597 , n65454 );
and ( n65599 , n65595 , n65598 );
and ( n65600 , n65591 , n65598 );
or ( n65601 , n65596 , n65599 , n65600 );
xor ( n65602 , n65457 , n65461 );
xor ( n65603 , n65602 , n65466 );
and ( n65604 , n65601 , n65603 );
xor ( n65605 , n65473 , n65477 );
xor ( n65606 , n65605 , n65479 );
and ( n65607 , n65603 , n65606 );
and ( n65608 , n65601 , n65606 );
or ( n65609 , n65604 , n65607 , n65608 );
xor ( n65610 , n65410 , n65414 );
xor ( n65611 , n65610 , n65419 );
and ( n65612 , n65609 , n65611 );
xor ( n65613 , n65469 , n65482 );
xor ( n65614 , n65613 , n65485 );
and ( n65615 , n65611 , n65614 );
and ( n65616 , n65609 , n65614 );
or ( n65617 , n65612 , n65615 , n65616 );
and ( n65618 , n65001 , n64789 );
and ( n65619 , n64955 , n64787 );
nor ( n65620 , n65618 , n65619 );
xnor ( n65621 , n65620 , n64738 );
and ( n65622 , n65175 , n64711 );
and ( n65623 , n65135 , n64709 );
nor ( n65624 , n65622 , n65623 );
xnor ( n65625 , n65624 , n64682 );
and ( n65626 , n65621 , n65625 );
and ( n65627 , n65363 , n64652 );
and ( n65628 , n65265 , n64650 );
nor ( n65629 , n65627 , n65628 );
xnor ( n65630 , n65629 , n64609 );
and ( n65631 , n65625 , n65630 );
and ( n65632 , n65621 , n65630 );
or ( n65633 , n65626 , n65631 , n65632 );
and ( n65634 , n64662 , n65371 );
and ( n65635 , n64627 , n65369 );
nor ( n65636 , n65634 , n65635 );
xnor ( n65637 , n65636 , n65168 );
and ( n65638 , n65633 , n65637 );
and ( n65639 , n64798 , n65056 );
and ( n65640 , n64781 , n65054 );
nor ( n65641 , n65639 , n65640 );
xnor ( n65642 , n65641 , n64943 );
and ( n65643 , n65637 , n65642 );
and ( n65644 , n65633 , n65642 );
or ( n65645 , n65638 , n65643 , n65644 );
buf ( n65646 , n64593 );
buf ( n65647 , n64594 );
and ( n65648 , n65646 , n65647 );
not ( n65649 , n65648 );
and ( n65650 , n65447 , n65649 );
not ( n65651 , n65650 );
and ( n65652 , n65443 , n64617 );
and ( n65653 , n65453 , n64615 );
nor ( n65654 , n65652 , n65653 );
xnor ( n65655 , n65654 , n64624 );
and ( n65656 , n65651 , n65655 );
buf ( n65657 , n64527 );
and ( n65658 , n65657 , n64612 );
and ( n65659 , n65655 , n65658 );
and ( n65660 , n65651 , n65658 );
or ( n65661 , n65656 , n65659 , n65660 );
and ( n65662 , n65453 , n64617 );
and ( n65663 , n65306 , n64615 );
nor ( n65664 , n65662 , n65663 );
xnor ( n65665 , n65664 , n64624 );
and ( n65666 , n65661 , n65665 );
not ( n65667 , n65444 );
and ( n65668 , n65665 , n65667 );
and ( n65669 , n65661 , n65667 );
or ( n65670 , n65666 , n65668 , n65669 );
and ( n65671 , n64611 , n65550 );
and ( n65672 , n64619 , n65548 );
nor ( n65673 , n65671 , n65672 );
xnor ( n65674 , n65673 , n65313 );
and ( n65675 , n65670 , n65674 );
and ( n65676 , n64703 , n65183 );
and ( n65677 , n64689 , n65181 );
nor ( n65678 , n65676 , n65677 );
xnor ( n65679 , n65678 , n64994 );
and ( n65680 , n65674 , n65679 );
and ( n65681 , n65670 , n65679 );
or ( n65682 , n65675 , n65680 , n65681 );
and ( n65683 , n65645 , n65682 );
xor ( n65684 , n65546 , n65553 );
xor ( n65685 , n65684 , n65558 );
and ( n65686 , n65682 , n65685 );
and ( n65687 , n65645 , n65685 );
or ( n65688 , n65683 , n65686 , n65687 );
and ( n65689 , n65453 , n64652 );
and ( n65690 , n65306 , n64650 );
nor ( n65691 , n65689 , n65690 );
xnor ( n65692 , n65691 , n64609 );
and ( n65693 , n65657 , n64617 );
and ( n65694 , n65443 , n64615 );
nor ( n65695 , n65693 , n65694 );
xnor ( n65696 , n65695 , n64624 );
and ( n65697 , n65692 , n65696 );
buf ( n65698 , n64528 );
and ( n65699 , n65698 , n64612 );
not ( n65700 , n65699 );
and ( n65701 , n65696 , n65700 );
and ( n65702 , n65692 , n65700 );
or ( n65703 , n65697 , n65701 , n65702 );
buf ( n65704 , n65699 );
and ( n65705 , n65703 , n65704 );
xor ( n65706 , n65651 , n65655 );
xor ( n65707 , n65706 , n65658 );
and ( n65708 , n65704 , n65707 );
and ( n65709 , n65703 , n65707 );
or ( n65710 , n65705 , n65708 , n65709 );
and ( n65711 , n64950 , n64897 );
and ( n65712 , n64906 , n64895 );
nor ( n65713 , n65711 , n65712 );
xnor ( n65714 , n65713 , n64850 );
and ( n65715 , n65710 , n65714 );
xor ( n65716 , n65661 , n65665 );
xor ( n65717 , n65716 , n65667 );
and ( n65718 , n65714 , n65717 );
and ( n65719 , n65710 , n65717 );
or ( n65720 , n65715 , n65718 , n65719 );
xor ( n65721 , n65534 , n65538 );
xor ( n65722 , n65721 , n65543 );
and ( n65723 , n65720 , n65722 );
xor ( n65724 , n65591 , n65595 );
xor ( n65725 , n65724 , n65598 );
and ( n65726 , n65722 , n65725 );
and ( n65727 , n65720 , n65725 );
or ( n65728 , n65723 , n65726 , n65727 );
xor ( n65729 , n65518 , n65522 );
xor ( n65730 , n65729 , n65527 );
and ( n65731 , n65728 , n65730 );
xor ( n65732 , n65601 , n65603 );
xor ( n65733 , n65732 , n65606 );
and ( n65734 , n65730 , n65733 );
and ( n65735 , n65728 , n65733 );
or ( n65736 , n65731 , n65734 , n65735 );
and ( n65737 , n65688 , n65736 );
xor ( n65738 , n65530 , n65561 );
xor ( n65739 , n65738 , n65564 );
and ( n65740 , n65736 , n65739 );
and ( n65741 , n65688 , n65739 );
or ( n65742 , n65737 , n65740 , n65741 );
and ( n65743 , n65617 , n65742 );
xor ( n65744 , n65567 , n65569 );
xor ( n65745 , n65744 , n65572 );
and ( n65746 , n65742 , n65745 );
and ( n65747 , n65617 , n65745 );
or ( n65748 , n65743 , n65746 , n65747 );
and ( n65749 , n65587 , n65748 );
xor ( n65750 , n65587 , n65748 );
xor ( n65751 , n65617 , n65742 );
xor ( n65752 , n65751 , n65745 );
xor ( n65753 , n65310 , n65446 );
xor ( n65754 , n65446 , n65447 );
not ( n65755 , n65754 );
and ( n65756 , n65753 , n65755 );
and ( n65757 , n64619 , n65756 );
not ( n65758 , n65757 );
xnor ( n65759 , n65758 , n65450 );
and ( n65760 , n64689 , n65371 );
and ( n65761 , n64662 , n65369 );
nor ( n65762 , n65760 , n65761 );
xnor ( n65763 , n65762 , n65168 );
and ( n65764 , n65759 , n65763 );
and ( n65765 , n64857 , n65056 );
and ( n65766 , n64798 , n65054 );
nor ( n65767 , n65765 , n65766 );
xnor ( n65768 , n65767 , n64943 );
and ( n65769 , n65763 , n65768 );
and ( n65770 , n65759 , n65768 );
or ( n65771 , n65764 , n65769 , n65770 );
and ( n65772 , n65135 , n64789 );
and ( n65773 , n65001 , n64787 );
nor ( n65774 , n65772 , n65773 );
xnor ( n65775 , n65774 , n64738 );
and ( n65776 , n65265 , n64711 );
and ( n65777 , n65175 , n64709 );
nor ( n65778 , n65776 , n65777 );
xnor ( n65779 , n65778 , n64682 );
and ( n65780 , n65775 , n65779 );
and ( n65781 , n65306 , n64652 );
and ( n65782 , n65363 , n64650 );
nor ( n65783 , n65781 , n65782 );
xnor ( n65784 , n65783 , n64609 );
and ( n65785 , n65779 , n65784 );
and ( n65786 , n65775 , n65784 );
or ( n65787 , n65780 , n65785 , n65786 );
and ( n65788 , n64627 , n65550 );
and ( n65789 , n64611 , n65548 );
nor ( n65790 , n65788 , n65789 );
xnor ( n65791 , n65790 , n65313 );
and ( n65792 , n65787 , n65791 );
and ( n65793 , n64781 , n65183 );
and ( n65794 , n64703 , n65181 );
nor ( n65795 , n65793 , n65794 );
xnor ( n65796 , n65795 , n64994 );
and ( n65797 , n65791 , n65796 );
and ( n65798 , n65787 , n65796 );
or ( n65799 , n65792 , n65797 , n65798 );
and ( n65800 , n65771 , n65799 );
xor ( n65801 , n65633 , n65637 );
xor ( n65802 , n65801 , n65642 );
and ( n65803 , n65799 , n65802 );
and ( n65804 , n65771 , n65802 );
or ( n65805 , n65800 , n65803 , n65804 );
and ( n65806 , n64703 , n65371 );
and ( n65807 , n64689 , n65369 );
nor ( n65808 , n65806 , n65807 );
xnor ( n65809 , n65808 , n65168 );
and ( n65810 , n64906 , n65056 );
and ( n65811 , n64857 , n65054 );
nor ( n65812 , n65810 , n65811 );
xnor ( n65813 , n65812 , n64943 );
and ( n65814 , n65809 , n65813 );
and ( n65815 , n64955 , n64897 );
and ( n65816 , n64950 , n64895 );
nor ( n65817 , n65815 , n65816 );
xnor ( n65818 , n65817 , n64850 );
and ( n65819 , n65813 , n65818 );
and ( n65820 , n65809 , n65818 );
or ( n65821 , n65814 , n65819 , n65820 );
xor ( n65822 , n65621 , n65625 );
xor ( n65823 , n65822 , n65630 );
and ( n65824 , n65821 , n65823 );
xor ( n65825 , n65710 , n65714 );
xor ( n65826 , n65825 , n65717 );
and ( n65827 , n65823 , n65826 );
and ( n65828 , n65821 , n65826 );
or ( n65829 , n65824 , n65827 , n65828 );
xor ( n65830 , n65670 , n65674 );
xor ( n65831 , n65830 , n65679 );
and ( n65832 , n65829 , n65831 );
xor ( n65833 , n65720 , n65722 );
xor ( n65834 , n65833 , n65725 );
and ( n65835 , n65831 , n65834 );
and ( n65836 , n65829 , n65834 );
or ( n65837 , n65832 , n65835 , n65836 );
and ( n65838 , n65805 , n65837 );
xor ( n65839 , n65645 , n65682 );
xor ( n65840 , n65839 , n65685 );
and ( n65841 , n65837 , n65840 );
and ( n65842 , n65805 , n65840 );
or ( n65843 , n65838 , n65841 , n65842 );
xor ( n65844 , n65609 , n65611 );
xor ( n65845 , n65844 , n65614 );
and ( n65846 , n65843 , n65845 );
xor ( n65847 , n65688 , n65736 );
xor ( n65848 , n65847 , n65739 );
and ( n65849 , n65845 , n65848 );
and ( n65850 , n65843 , n65848 );
or ( n65851 , n65846 , n65849 , n65850 );
and ( n65852 , n65752 , n65851 );
xor ( n65853 , n65752 , n65851 );
xor ( n65854 , n65843 , n65845 );
xor ( n65855 , n65854 , n65848 );
and ( n65856 , n64950 , n65056 );
and ( n65857 , n64906 , n65054 );
nor ( n65858 , n65856 , n65857 );
xnor ( n65859 , n65858 , n64943 );
and ( n65860 , n65001 , n64897 );
and ( n65861 , n64955 , n64895 );
nor ( n65862 , n65860 , n65861 );
xnor ( n65863 , n65862 , n64850 );
and ( n65864 , n65859 , n65863 );
and ( n65865 , n65175 , n64789 );
and ( n65866 , n65135 , n64787 );
nor ( n65867 , n65865 , n65866 );
xnor ( n65868 , n65867 , n64738 );
and ( n65869 , n65863 , n65868 );
and ( n65870 , n65859 , n65868 );
or ( n65871 , n65864 , n65869 , n65870 );
buf ( n65872 , n64595 );
buf ( n65873 , n64596 );
and ( n65874 , n65872 , n65873 );
not ( n65875 , n65874 );
and ( n65876 , n65647 , n65875 );
not ( n65877 , n65876 );
and ( n65878 , n65698 , n64617 );
and ( n65879 , n65657 , n64615 );
nor ( n65880 , n65878 , n65879 );
xnor ( n65881 , n65880 , n64624 );
and ( n65882 , n65877 , n65881 );
buf ( n65883 , n64529 );
and ( n65884 , n65883 , n64612 );
and ( n65885 , n65881 , n65884 );
and ( n65886 , n65877 , n65884 );
or ( n65887 , n65882 , n65885 , n65886 );
and ( n65888 , n65363 , n64711 );
and ( n65889 , n65265 , n64709 );
nor ( n65890 , n65888 , n65889 );
xnor ( n65891 , n65890 , n64682 );
and ( n65892 , n65887 , n65891 );
xor ( n65893 , n65692 , n65696 );
xor ( n65894 , n65893 , n65700 );
and ( n65895 , n65891 , n65894 );
and ( n65896 , n65887 , n65894 );
or ( n65897 , n65892 , n65895 , n65896 );
and ( n65898 , n65871 , n65897 );
and ( n65899 , n64662 , n65550 );
and ( n65900 , n64627 , n65548 );
nor ( n65901 , n65899 , n65900 );
xnor ( n65902 , n65901 , n65313 );
and ( n65903 , n65897 , n65902 );
and ( n65904 , n65871 , n65902 );
or ( n65905 , n65898 , n65903 , n65904 );
and ( n65906 , n64611 , n65756 );
and ( n65907 , n64619 , n65754 );
nor ( n65908 , n65906 , n65907 );
xnor ( n65909 , n65908 , n65450 );
and ( n65910 , n64798 , n65183 );
and ( n65911 , n64781 , n65181 );
nor ( n65912 , n65910 , n65911 );
xnor ( n65913 , n65912 , n64994 );
and ( n65914 , n65909 , n65913 );
xor ( n65915 , n65703 , n65704 );
xor ( n65916 , n65915 , n65707 );
and ( n65917 , n65913 , n65916 );
and ( n65918 , n65909 , n65916 );
or ( n65919 , n65914 , n65917 , n65918 );
and ( n65920 , n65905 , n65919 );
xor ( n65921 , n65759 , n65763 );
xor ( n65922 , n65921 , n65768 );
and ( n65923 , n65919 , n65922 );
and ( n65924 , n65905 , n65922 );
or ( n65925 , n65920 , n65923 , n65924 );
and ( n65926 , n65453 , n64711 );
and ( n65927 , n65306 , n64709 );
nor ( n65928 , n65926 , n65927 );
xnor ( n65929 , n65928 , n64682 );
and ( n65930 , n65657 , n64652 );
and ( n65931 , n65443 , n64650 );
nor ( n65932 , n65930 , n65931 );
xnor ( n65933 , n65932 , n64609 );
and ( n65934 , n65929 , n65933 );
buf ( n65935 , n64530 );
and ( n65936 , n65935 , n64612 );
and ( n65937 , n65933 , n65936 );
and ( n65938 , n65929 , n65936 );
or ( n65939 , n65934 , n65937 , n65938 );
and ( n65940 , n65135 , n64897 );
and ( n65941 , n65001 , n64895 );
nor ( n65942 , n65940 , n65941 );
xnor ( n65943 , n65942 , n64850 );
and ( n65944 , n65939 , n65943 );
and ( n65945 , n65265 , n64789 );
and ( n65946 , n65175 , n64787 );
nor ( n65947 , n65945 , n65946 );
xnor ( n65948 , n65947 , n64738 );
and ( n65949 , n65943 , n65948 );
and ( n65950 , n65939 , n65948 );
or ( n65951 , n65944 , n65949 , n65950 );
and ( n65952 , n65883 , n64617 );
and ( n65953 , n65698 , n64615 );
nor ( n65954 , n65952 , n65953 );
xnor ( n65955 , n65954 , n64624 );
buf ( n65956 , n65955 );
and ( n65957 , n65443 , n64652 );
and ( n65958 , n65453 , n64650 );
nor ( n65959 , n65957 , n65958 );
xnor ( n65960 , n65959 , n64609 );
and ( n65961 , n65956 , n65960 );
xor ( n65962 , n65877 , n65881 );
xor ( n65963 , n65962 , n65884 );
and ( n65964 , n65960 , n65963 );
and ( n65965 , n65956 , n65963 );
or ( n65966 , n65961 , n65964 , n65965 );
and ( n65967 , n65951 , n65966 );
and ( n65968 , n64781 , n65371 );
and ( n65969 , n64703 , n65369 );
nor ( n65970 , n65968 , n65969 );
xnor ( n65971 , n65970 , n65168 );
and ( n65972 , n65966 , n65971 );
and ( n65973 , n65951 , n65971 );
or ( n65974 , n65967 , n65972 , n65973 );
xor ( n65975 , n65775 , n65779 );
xor ( n65976 , n65975 , n65784 );
and ( n65977 , n65974 , n65976 );
xor ( n65978 , n65809 , n65813 );
xor ( n65979 , n65978 , n65818 );
and ( n65980 , n65976 , n65979 );
and ( n65981 , n65974 , n65979 );
or ( n65982 , n65977 , n65980 , n65981 );
and ( n65983 , n64627 , n65756 );
and ( n65984 , n64611 , n65754 );
nor ( n65985 , n65983 , n65984 );
xnor ( n65986 , n65985 , n65450 );
and ( n65987 , n64689 , n65550 );
and ( n65988 , n64662 , n65548 );
nor ( n65989 , n65987 , n65988 );
xnor ( n65990 , n65989 , n65313 );
and ( n65991 , n65986 , n65990 );
and ( n65992 , n64857 , n65183 );
and ( n65993 , n64798 , n65181 );
nor ( n65994 , n65992 , n65993 );
xnor ( n65995 , n65994 , n64994 );
and ( n65996 , n65990 , n65995 );
and ( n65997 , n65986 , n65995 );
or ( n65998 , n65991 , n65996 , n65997 );
and ( n65999 , n64955 , n65056 );
and ( n66000 , n64950 , n65054 );
nor ( n66001 , n65999 , n66000 );
xnor ( n66002 , n66001 , n64943 );
and ( n66003 , n65306 , n64711 );
and ( n66004 , n65363 , n64709 );
nor ( n66005 , n66003 , n66004 );
xnor ( n66006 , n66005 , n64682 );
and ( n66007 , n66002 , n66006 );
xor ( n66008 , n65956 , n65960 );
xor ( n66009 , n66008 , n65963 );
and ( n66010 , n66006 , n66009 );
and ( n66011 , n66002 , n66009 );
or ( n66012 , n66007 , n66010 , n66011 );
xor ( n66013 , n65447 , n65646 );
xor ( n66014 , n65646 , n65647 );
not ( n66015 , n66014 );
and ( n66016 , n66013 , n66015 );
and ( n66017 , n64619 , n66016 );
not ( n66018 , n66017 );
xnor ( n66019 , n66018 , n65650 );
and ( n66020 , n66012 , n66019 );
xor ( n66021 , n65859 , n65863 );
xor ( n66022 , n66021 , n65868 );
and ( n66023 , n66019 , n66022 );
and ( n66024 , n66012 , n66022 );
or ( n66025 , n66020 , n66023 , n66024 );
and ( n66026 , n65998 , n66025 );
xor ( n66027 , n65871 , n65897 );
xor ( n66028 , n66027 , n65902 );
and ( n66029 , n66025 , n66028 );
and ( n66030 , n65998 , n66028 );
or ( n66031 , n66026 , n66029 , n66030 );
and ( n66032 , n65982 , n66031 );
xor ( n66033 , n65787 , n65791 );
xor ( n66034 , n66033 , n65796 );
and ( n66035 , n66031 , n66034 );
and ( n66036 , n65982 , n66034 );
or ( n66037 , n66032 , n66035 , n66036 );
and ( n66038 , n65925 , n66037 );
xor ( n66039 , n65771 , n65799 );
xor ( n66040 , n66039 , n65802 );
and ( n66041 , n66037 , n66040 );
and ( n66042 , n65925 , n66040 );
or ( n66043 , n66038 , n66041 , n66042 );
xor ( n66044 , n65728 , n65730 );
xor ( n66045 , n66044 , n65733 );
and ( n66046 , n66043 , n66045 );
xor ( n66047 , n65805 , n65837 );
xor ( n66048 , n66047 , n65840 );
and ( n66049 , n66045 , n66048 );
and ( n66050 , n66043 , n66048 );
or ( n66051 , n66046 , n66049 , n66050 );
and ( n66052 , n65855 , n66051 );
xor ( n66053 , n65855 , n66051 );
xor ( n66054 , n66043 , n66045 );
xor ( n66055 , n66054 , n66048 );
xor ( n66056 , n65905 , n65919 );
xor ( n66057 , n66056 , n65922 );
xor ( n66058 , n65982 , n66031 );
xor ( n66059 , n66058 , n66034 );
and ( n66060 , n66057 , n66059 );
xor ( n66061 , n65821 , n65823 );
xor ( n66062 , n66061 , n65826 );
and ( n66063 , n66059 , n66062 );
and ( n66064 , n66057 , n66062 );
or ( n66065 , n66060 , n66063 , n66064 );
xor ( n66066 , n65925 , n66037 );
xor ( n66067 , n66066 , n66040 );
and ( n66068 , n66065 , n66067 );
xor ( n66069 , n65829 , n65831 );
xor ( n66070 , n66069 , n65834 );
and ( n66071 , n66067 , n66070 );
and ( n66072 , n66065 , n66070 );
or ( n66073 , n66068 , n66071 , n66072 );
and ( n66074 , n66055 , n66073 );
xor ( n66075 , n66055 , n66073 );
xor ( n66076 , n66065 , n66067 );
xor ( n66077 , n66076 , n66070 );
and ( n66078 , n64662 , n65756 );
and ( n66079 , n64627 , n65754 );
nor ( n66080 , n66078 , n66079 );
xnor ( n66081 , n66080 , n65450 );
xor ( n66082 , n65939 , n65943 );
xor ( n66083 , n66082 , n65948 );
and ( n66084 , n66081 , n66083 );
xor ( n66085 , n66002 , n66006 );
xor ( n66086 , n66085 , n66009 );
and ( n66087 , n66083 , n66086 );
and ( n66088 , n66081 , n66086 );
or ( n66089 , n66084 , n66087 , n66088 );
xor ( n66090 , n65986 , n65990 );
xor ( n66091 , n66090 , n65995 );
and ( n66092 , n66089 , n66091 );
xor ( n66093 , n65951 , n65966 );
xor ( n66094 , n66093 , n65971 );
and ( n66095 , n66091 , n66094 );
and ( n66096 , n66089 , n66094 );
or ( n66097 , n66092 , n66095 , n66096 );
and ( n66098 , n65001 , n65056 );
and ( n66099 , n64955 , n65054 );
nor ( n66100 , n66098 , n66099 );
xnor ( n66101 , n66100 , n64943 );
and ( n66102 , n65175 , n64897 );
and ( n66103 , n65135 , n64895 );
nor ( n66104 , n66102 , n66103 );
xnor ( n66105 , n66104 , n64850 );
and ( n66106 , n66101 , n66105 );
and ( n66107 , n65363 , n64789 );
and ( n66108 , n65265 , n64787 );
nor ( n66109 , n66107 , n66108 );
xnor ( n66110 , n66109 , n64738 );
and ( n66111 , n66105 , n66110 );
and ( n66112 , n66101 , n66110 );
or ( n66113 , n66106 , n66111 , n66112 );
and ( n66114 , n64611 , n66016 );
and ( n66115 , n64619 , n66014 );
nor ( n66116 , n66114 , n66115 );
xnor ( n66117 , n66116 , n65650 );
and ( n66118 , n66113 , n66117 );
and ( n66119 , n64798 , n65371 );
and ( n66120 , n64781 , n65369 );
nor ( n66121 , n66119 , n66120 );
xnor ( n66122 , n66121 , n65168 );
and ( n66123 , n66117 , n66122 );
and ( n66124 , n66113 , n66122 );
or ( n66125 , n66118 , n66123 , n66124 );
buf ( n66126 , n64597 );
buf ( n66127 , n64598 );
and ( n66128 , n66126 , n66127 );
not ( n66129 , n66128 );
and ( n66130 , n65873 , n66129 );
not ( n66131 , n66130 );
and ( n66132 , n65935 , n64617 );
and ( n66133 , n65883 , n64615 );
nor ( n66134 , n66132 , n66133 );
xnor ( n66135 , n66134 , n64624 );
and ( n66136 , n66131 , n66135 );
buf ( n66137 , n64531 );
and ( n66138 , n66137 , n64612 );
and ( n66139 , n66135 , n66138 );
and ( n66140 , n66131 , n66138 );
or ( n66141 , n66136 , n66139 , n66140 );
buf ( n66142 , n64532 );
and ( n66143 , n66142 , n64612 );
buf ( n66144 , n66143 );
and ( n66145 , n65443 , n64711 );
and ( n66146 , n65453 , n64709 );
nor ( n66147 , n66145 , n66146 );
xnor ( n66148 , n66147 , n64682 );
and ( n66149 , n66144 , n66148 );
and ( n66150 , n65698 , n64652 );
and ( n66151 , n65657 , n64650 );
nor ( n66152 , n66150 , n66151 );
xnor ( n66153 , n66152 , n64609 );
and ( n66154 , n66148 , n66153 );
and ( n66155 , n66144 , n66153 );
or ( n66156 , n66149 , n66154 , n66155 );
and ( n66157 , n66141 , n66156 );
not ( n66158 , n65955 );
and ( n66159 , n66156 , n66158 );
and ( n66160 , n66141 , n66158 );
or ( n66161 , n66157 , n66159 , n66160 );
and ( n66162 , n64703 , n65550 );
and ( n66163 , n64689 , n65548 );
nor ( n66164 , n66162 , n66163 );
xnor ( n66165 , n66164 , n65313 );
and ( n66166 , n66161 , n66165 );
and ( n66167 , n64906 , n65183 );
and ( n66168 , n64857 , n65181 );
nor ( n66169 , n66167 , n66168 );
xnor ( n66170 , n66169 , n64994 );
and ( n66171 , n66165 , n66170 );
and ( n66172 , n66161 , n66170 );
or ( n66173 , n66166 , n66171 , n66172 );
and ( n66174 , n66125 , n66173 );
xor ( n66175 , n65887 , n65891 );
xor ( n66176 , n66175 , n65894 );
and ( n66177 , n66173 , n66176 );
and ( n66178 , n66125 , n66176 );
or ( n66179 , n66174 , n66177 , n66178 );
and ( n66180 , n66097 , n66179 );
xor ( n66181 , n65909 , n65913 );
xor ( n66182 , n66181 , n65916 );
and ( n66183 , n66179 , n66182 );
and ( n66184 , n66097 , n66182 );
or ( n66185 , n66180 , n66183 , n66184 );
xor ( n66186 , n65974 , n65976 );
xor ( n66187 , n66186 , n65979 );
xor ( n66188 , n65998 , n66025 );
xor ( n66189 , n66188 , n66028 );
and ( n66190 , n66187 , n66189 );
xor ( n66191 , n66097 , n66179 );
xor ( n66192 , n66191 , n66182 );
and ( n66193 , n66189 , n66192 );
and ( n66194 , n66187 , n66192 );
or ( n66195 , n66190 , n66193 , n66194 );
and ( n66196 , n66185 , n66195 );
xor ( n66197 , n66057 , n66059 );
xor ( n66198 , n66197 , n66062 );
and ( n66199 , n66195 , n66198 );
and ( n66200 , n66185 , n66198 );
or ( n66201 , n66196 , n66199 , n66200 );
and ( n66202 , n66077 , n66201 );
xor ( n66203 , n66077 , n66201 );
xor ( n66204 , n66185 , n66195 );
xor ( n66205 , n66204 , n66198 );
and ( n66206 , n64627 , n66016 );
and ( n66207 , n64611 , n66014 );
nor ( n66208 , n66206 , n66207 );
xnor ( n66209 , n66208 , n65650 );
and ( n66210 , n64689 , n65756 );
and ( n66211 , n64662 , n65754 );
nor ( n66212 , n66210 , n66211 );
xnor ( n66213 , n66212 , n65450 );
and ( n66214 , n66209 , n66213 );
and ( n66215 , n64857 , n65371 );
and ( n66216 , n64798 , n65369 );
nor ( n66217 , n66215 , n66216 );
xnor ( n66218 , n66217 , n65168 );
and ( n66219 , n66213 , n66218 );
and ( n66220 , n66209 , n66218 );
or ( n66221 , n66214 , n66219 , n66220 );
and ( n66222 , n64906 , n65371 );
and ( n66223 , n64857 , n65369 );
nor ( n66224 , n66222 , n66223 );
xnor ( n66225 , n66224 , n65168 );
and ( n66226 , n64955 , n65183 );
and ( n66227 , n64950 , n65181 );
nor ( n66228 , n66226 , n66227 );
xnor ( n66229 , n66228 , n64994 );
and ( n66230 , n66225 , n66229 );
and ( n66231 , n65306 , n64789 );
and ( n66232 , n65363 , n64787 );
nor ( n66233 , n66231 , n66232 );
xnor ( n66234 , n66233 , n64738 );
and ( n66235 , n66229 , n66234 );
and ( n66236 , n66225 , n66234 );
or ( n66237 , n66230 , n66235 , n66236 );
xor ( n66238 , n65647 , n65872 );
xor ( n66239 , n65872 , n65873 );
not ( n66240 , n66239 );
and ( n66241 , n66238 , n66240 );
and ( n66242 , n64619 , n66241 );
not ( n66243 , n66242 );
xnor ( n66244 , n66243 , n65876 );
and ( n66245 , n66237 , n66244 );
xor ( n66246 , n66101 , n66105 );
xor ( n66247 , n66246 , n66110 );
and ( n66248 , n66244 , n66247 );
and ( n66249 , n66237 , n66247 );
or ( n66250 , n66245 , n66248 , n66249 );
and ( n66251 , n66221 , n66250 );
xor ( n66252 , n66113 , n66117 );
xor ( n66253 , n66252 , n66122 );
and ( n66254 , n66250 , n66253 );
and ( n66255 , n66221 , n66253 );
or ( n66256 , n66251 , n66254 , n66255 );
and ( n66257 , n65883 , n64711 );
and ( n66258 , n65698 , n64709 );
nor ( n66259 , n66257 , n66258 );
xnor ( n66260 , n66259 , n64682 );
and ( n66261 , n66137 , n64652 );
and ( n66262 , n65935 , n64650 );
nor ( n66263 , n66261 , n66262 );
xnor ( n66264 , n66263 , n64609 );
and ( n66265 , n66260 , n66264 );
buf ( n66266 , n64534 );
and ( n66267 , n66266 , n64612 );
and ( n66268 , n66264 , n66267 );
and ( n66269 , n66260 , n66267 );
or ( n66270 , n66265 , n66268 , n66269 );
and ( n66271 , n65443 , n64789 );
and ( n66272 , n65453 , n64787 );
nor ( n66273 , n66271 , n66272 );
xnor ( n66274 , n66273 , n64738 );
and ( n66275 , n66270 , n66274 );
buf ( n66276 , n64533 );
and ( n66277 , n66276 , n64617 );
and ( n66278 , n66142 , n64615 );
nor ( n66279 , n66277 , n66278 );
xnor ( n66280 , n66279 , n64624 );
buf ( n66281 , n66280 );
buf ( n66282 , n64599 );
buf ( n66283 , n64600 );
and ( n66284 , n66282 , n66283 );
not ( n66285 , n66284 );
and ( n66286 , n66127 , n66285 );
not ( n66287 , n66286 );
xor ( n66288 , n66281 , n66287 );
and ( n66289 , n66276 , n64612 );
xor ( n66290 , n66288 , n66289 );
and ( n66291 , n66274 , n66290 );
and ( n66292 , n66270 , n66290 );
or ( n66293 , n66275 , n66291 , n66292 );
and ( n66294 , n65001 , n65183 );
and ( n66295 , n64955 , n65181 );
nor ( n66296 , n66294 , n66295 );
xnor ( n66297 , n66296 , n64994 );
and ( n66298 , n66293 , n66297 );
and ( n66299 , n65175 , n65056 );
and ( n66300 , n65135 , n65054 );
nor ( n66301 , n66299 , n66300 );
xnor ( n66302 , n66301 , n64943 );
and ( n66303 , n66297 , n66302 );
and ( n66304 , n66293 , n66302 );
or ( n66305 , n66298 , n66303 , n66304 );
and ( n66306 , n64611 , n66241 );
and ( n66307 , n64619 , n66239 );
nor ( n66308 , n66306 , n66307 );
xnor ( n66309 , n66308 , n65876 );
and ( n66310 , n66305 , n66309 );
and ( n66311 , n64798 , n65550 );
and ( n66312 , n64781 , n65548 );
nor ( n66313 , n66311 , n66312 );
xnor ( n66314 , n66313 , n65313 );
and ( n66315 , n66309 , n66314 );
and ( n66316 , n66305 , n66314 );
or ( n66317 , n66310 , n66315 , n66316 );
and ( n66318 , n65698 , n64711 );
and ( n66319 , n65657 , n64709 );
nor ( n66320 , n66318 , n66319 );
xnor ( n66321 , n66320 , n64682 );
and ( n66322 , n65935 , n64652 );
and ( n66323 , n65883 , n64650 );
nor ( n66324 , n66322 , n66323 );
xnor ( n66325 , n66324 , n64609 );
and ( n66326 , n66321 , n66325 );
and ( n66327 , n66142 , n64617 );
and ( n66328 , n66137 , n64615 );
nor ( n66329 , n66327 , n66328 );
xnor ( n66330 , n66329 , n64624 );
and ( n66331 , n66325 , n66330 );
and ( n66332 , n66321 , n66330 );
or ( n66333 , n66326 , n66331 , n66332 );
and ( n66334 , n65363 , n64897 );
and ( n66335 , n65265 , n64895 );
nor ( n66336 , n66334 , n66335 );
xnor ( n66337 , n66336 , n64850 );
and ( n66338 , n66333 , n66337 );
and ( n66339 , n65883 , n64652 );
and ( n66340 , n65698 , n64650 );
nor ( n66341 , n66339 , n66340 );
xnor ( n66342 , n66341 , n64609 );
and ( n66343 , n66137 , n64617 );
and ( n66344 , n65935 , n64615 );
nor ( n66345 , n66343 , n66344 );
xnor ( n66346 , n66345 , n64624 );
xor ( n66347 , n66342 , n66346 );
not ( n66348 , n66143 );
xor ( n66349 , n66347 , n66348 );
and ( n66350 , n66337 , n66349 );
and ( n66351 , n66333 , n66349 );
or ( n66352 , n66338 , n66350 , n66351 );
and ( n66353 , n64703 , n65756 );
and ( n66354 , n64689 , n65754 );
nor ( n66355 , n66353 , n66354 );
xnor ( n66356 , n66355 , n65450 );
and ( n66357 , n66352 , n66356 );
and ( n66358 , n66342 , n66346 );
and ( n66359 , n66346 , n66348 );
and ( n66360 , n66342 , n66348 );
or ( n66361 , n66358 , n66359 , n66360 );
xor ( n66362 , n66131 , n66135 );
xor ( n66363 , n66362 , n66138 );
xor ( n66364 , n66361 , n66363 );
xor ( n66365 , n66144 , n66148 );
xor ( n66366 , n66365 , n66153 );
xor ( n66367 , n66364 , n66366 );
and ( n66368 , n66356 , n66367 );
and ( n66369 , n66352 , n66367 );
or ( n66370 , n66357 , n66368 , n66369 );
and ( n66371 , n66317 , n66370 );
and ( n66372 , n66361 , n66363 );
and ( n66373 , n66363 , n66366 );
and ( n66374 , n66361 , n66366 );
or ( n66375 , n66372 , n66373 , n66374 );
and ( n66376 , n64950 , n65183 );
and ( n66377 , n64906 , n65181 );
nor ( n66378 , n66376 , n66377 );
xnor ( n66379 , n66378 , n64994 );
xor ( n66380 , n66375 , n66379 );
xor ( n66381 , n65929 , n65933 );
xor ( n66382 , n66381 , n65936 );
xor ( n66383 , n66380 , n66382 );
and ( n66384 , n66370 , n66383 );
and ( n66385 , n66317 , n66383 );
or ( n66386 , n66371 , n66384 , n66385 );
and ( n66387 , n66375 , n66379 );
and ( n66388 , n66379 , n66382 );
and ( n66389 , n66375 , n66382 );
or ( n66390 , n66387 , n66388 , n66389 );
and ( n66391 , n66281 , n66287 );
and ( n66392 , n66287 , n66289 );
and ( n66393 , n66281 , n66289 );
or ( n66394 , n66391 , n66392 , n66393 );
and ( n66395 , n65453 , n64789 );
and ( n66396 , n65306 , n64787 );
nor ( n66397 , n66395 , n66396 );
xnor ( n66398 , n66397 , n64738 );
and ( n66399 , n66394 , n66398 );
and ( n66400 , n65657 , n64711 );
and ( n66401 , n65443 , n64709 );
nor ( n66402 , n66400 , n66401 );
xnor ( n66403 , n66402 , n64682 );
and ( n66404 , n66398 , n66403 );
and ( n66405 , n66394 , n66403 );
or ( n66406 , n66399 , n66404 , n66405 );
and ( n66407 , n65135 , n65056 );
and ( n66408 , n65001 , n65054 );
nor ( n66409 , n66407 , n66408 );
xnor ( n66410 , n66409 , n64943 );
and ( n66411 , n66406 , n66410 );
and ( n66412 , n65265 , n64897 );
and ( n66413 , n65175 , n64895 );
nor ( n66414 , n66412 , n66413 );
xnor ( n66415 , n66414 , n64850 );
and ( n66416 , n66410 , n66415 );
and ( n66417 , n66406 , n66415 );
or ( n66418 , n66411 , n66416 , n66417 );
and ( n66419 , n64781 , n65550 );
and ( n66420 , n64703 , n65548 );
nor ( n66421 , n66419 , n66420 );
xnor ( n66422 , n66421 , n65313 );
and ( n66423 , n66418 , n66422 );
xor ( n66424 , n66141 , n66156 );
xor ( n66425 , n66424 , n66158 );
and ( n66426 , n66422 , n66425 );
and ( n66427 , n66418 , n66425 );
or ( n66428 , n66423 , n66426 , n66427 );
xor ( n66429 , n66390 , n66428 );
xor ( n66430 , n66161 , n66165 );
xor ( n66431 , n66430 , n66170 );
xor ( n66432 , n66429 , n66431 );
and ( n66433 , n66386 , n66432 );
xor ( n66434 , n66081 , n66083 );
xor ( n66435 , n66434 , n66086 );
and ( n66436 , n66432 , n66435 );
and ( n66437 , n66386 , n66435 );
or ( n66438 , n66433 , n66436 , n66437 );
and ( n66439 , n66256 , n66438 );
xor ( n66440 , n66089 , n66091 );
xor ( n66441 , n66440 , n66094 );
and ( n66442 , n66438 , n66441 );
and ( n66443 , n66256 , n66441 );
or ( n66444 , n66439 , n66442 , n66443 );
and ( n66445 , n66390 , n66428 );
and ( n66446 , n66428 , n66431 );
and ( n66447 , n66390 , n66431 );
or ( n66448 , n66445 , n66446 , n66447 );
xor ( n66449 , n66012 , n66019 );
xor ( n66450 , n66449 , n66022 );
and ( n66451 , n66448 , n66450 );
xor ( n66452 , n66125 , n66173 );
xor ( n66453 , n66452 , n66176 );
and ( n66454 , n66450 , n66453 );
and ( n66455 , n66448 , n66453 );
or ( n66456 , n66451 , n66454 , n66455 );
and ( n66457 , n66444 , n66456 );
xor ( n66458 , n66187 , n66189 );
xor ( n66459 , n66458 , n66192 );
and ( n66460 , n66456 , n66459 );
and ( n66461 , n66444 , n66459 );
or ( n66462 , n66457 , n66460 , n66461 );
and ( n66463 , n66205 , n66462 );
xor ( n66464 , n66205 , n66462 );
xor ( n66465 , n66444 , n66456 );
xor ( n66466 , n66465 , n66459 );
and ( n66467 , n64662 , n66016 );
and ( n66468 , n64627 , n66014 );
nor ( n66469 , n66467 , n66468 );
xnor ( n66470 , n66469 , n65650 );
xor ( n66471 , n66225 , n66229 );
xor ( n66472 , n66471 , n66234 );
and ( n66473 , n66470 , n66472 );
xor ( n66474 , n66406 , n66410 );
xor ( n66475 , n66474 , n66415 );
and ( n66476 , n66472 , n66475 );
and ( n66477 , n66470 , n66475 );
or ( n66478 , n66473 , n66476 , n66477 );
xor ( n66479 , n66209 , n66213 );
xor ( n66480 , n66479 , n66218 );
and ( n66481 , n66478 , n66480 );
xor ( n66482 , n66418 , n66422 );
xor ( n66483 , n66482 , n66425 );
and ( n66484 , n66480 , n66483 );
and ( n66485 , n66478 , n66483 );
or ( n66486 , n66481 , n66484 , n66485 );
xor ( n66487 , n66221 , n66250 );
xor ( n66488 , n66487 , n66253 );
and ( n66489 , n66486 , n66488 );
xor ( n66490 , n66386 , n66432 );
xor ( n66491 , n66490 , n66435 );
and ( n66492 , n66488 , n66491 );
and ( n66493 , n66486 , n66491 );
or ( n66494 , n66489 , n66492 , n66493 );
xor ( n66495 , n66256 , n66438 );
xor ( n66496 , n66495 , n66441 );
and ( n66497 , n66494 , n66496 );
xor ( n66498 , n66448 , n66450 );
xor ( n66499 , n66498 , n66453 );
and ( n66500 , n66496 , n66499 );
and ( n66501 , n66494 , n66499 );
or ( n66502 , n66497 , n66500 , n66501 );
and ( n66503 , n66466 , n66502 );
xor ( n66504 , n66466 , n66502 );
xor ( n66505 , n66494 , n66496 );
xor ( n66506 , n66505 , n66499 );
buf ( n66507 , n64536 );
and ( n66508 , n66507 , n64612 );
buf ( n66509 , n66508 );
buf ( n66510 , n64601 );
buf ( n66511 , n64602 );
and ( n66512 , n66510 , n66511 );
not ( n66513 , n66512 );
and ( n66514 , n66283 , n66513 );
not ( n66515 , n66514 );
and ( n66516 , n66509 , n66515 );
buf ( n66517 , n64535 );
and ( n66518 , n66517 , n64612 );
and ( n66519 , n66515 , n66518 );
and ( n66520 , n66509 , n66518 );
or ( n66521 , n66516 , n66519 , n66520 );
and ( n66522 , n65657 , n64789 );
and ( n66523 , n65443 , n64787 );
nor ( n66524 , n66522 , n66523 );
xnor ( n66525 , n66524 , n64738 );
and ( n66526 , n66521 , n66525 );
not ( n66527 , n66280 );
and ( n66528 , n66525 , n66527 );
and ( n66529 , n66521 , n66527 );
or ( n66530 , n66526 , n66528 , n66529 );
and ( n66531 , n65265 , n65056 );
and ( n66532 , n65175 , n65054 );
nor ( n66533 , n66531 , n66532 );
xnor ( n66534 , n66533 , n64943 );
and ( n66535 , n66530 , n66534 );
xor ( n66536 , n66321 , n66325 );
xor ( n66537 , n66536 , n66330 );
and ( n66538 , n66534 , n66537 );
and ( n66539 , n66530 , n66537 );
or ( n66540 , n66535 , n66538 , n66539 );
and ( n66541 , n64627 , n66241 );
and ( n66542 , n64611 , n66239 );
nor ( n66543 , n66541 , n66542 );
xnor ( n66544 , n66543 , n65876 );
and ( n66545 , n66540 , n66544 );
and ( n66546 , n64857 , n65550 );
and ( n66547 , n64798 , n65548 );
nor ( n66548 , n66546 , n66547 );
xnor ( n66549 , n66548 , n65313 );
and ( n66550 , n66544 , n66549 );
and ( n66551 , n66540 , n66549 );
or ( n66552 , n66545 , n66550 , n66551 );
and ( n66553 , n64781 , n65756 );
and ( n66554 , n64703 , n65754 );
nor ( n66555 , n66553 , n66554 );
xnor ( n66556 , n66555 , n65450 );
and ( n66557 , n64950 , n65371 );
and ( n66558 , n64906 , n65369 );
nor ( n66559 , n66557 , n66558 );
xnor ( n66560 , n66559 , n65168 );
and ( n66561 , n66556 , n66560 );
xor ( n66562 , n66394 , n66398 );
xor ( n66563 , n66562 , n66403 );
and ( n66564 , n66560 , n66563 );
and ( n66565 , n66556 , n66563 );
or ( n66566 , n66561 , n66564 , n66565 );
and ( n66567 , n66552 , n66566 );
and ( n66568 , n64955 , n65371 );
and ( n66569 , n64950 , n65369 );
nor ( n66570 , n66568 , n66569 );
xnor ( n66571 , n66570 , n65168 );
and ( n66572 , n65135 , n65183 );
and ( n66573 , n65001 , n65181 );
nor ( n66574 , n66572 , n66573 );
xnor ( n66575 , n66574 , n64994 );
and ( n66576 , n66571 , n66575 );
and ( n66577 , n65306 , n64897 );
and ( n66578 , n65363 , n64895 );
nor ( n66579 , n66577 , n66578 );
xnor ( n66580 , n66579 , n64850 );
and ( n66581 , n66575 , n66580 );
and ( n66582 , n66571 , n66580 );
or ( n66583 , n66576 , n66581 , n66582 );
and ( n66584 , n64689 , n66016 );
and ( n66585 , n64662 , n66014 );
nor ( n66586 , n66584 , n66585 );
xnor ( n66587 , n66586 , n65650 );
and ( n66588 , n66583 , n66587 );
xor ( n66589 , n66333 , n66337 );
xor ( n66590 , n66589 , n66349 );
and ( n66591 , n66587 , n66590 );
and ( n66592 , n66583 , n66590 );
or ( n66593 , n66588 , n66591 , n66592 );
and ( n66594 , n66566 , n66593 );
and ( n66595 , n66552 , n66593 );
or ( n66596 , n66567 , n66594 , n66595 );
and ( n66597 , n65935 , n64711 );
and ( n66598 , n65883 , n64709 );
nor ( n66599 , n66597 , n66598 );
xnor ( n66600 , n66599 , n64682 );
and ( n66601 , n66142 , n64652 );
and ( n66602 , n66137 , n64650 );
nor ( n66603 , n66601 , n66602 );
xnor ( n66604 , n66603 , n64609 );
and ( n66605 , n66600 , n66604 );
and ( n66606 , n66266 , n64617 );
and ( n66607 , n66276 , n64615 );
nor ( n66608 , n66606 , n66607 );
xnor ( n66609 , n66608 , n64624 );
and ( n66610 , n66604 , n66609 );
and ( n66611 , n66600 , n66609 );
or ( n66612 , n66605 , n66610 , n66611 );
and ( n66613 , n66276 , n64652 );
and ( n66614 , n66142 , n64650 );
nor ( n66615 , n66613 , n66614 );
xnor ( n66616 , n66615 , n64609 );
and ( n66617 , n66517 , n64617 );
and ( n66618 , n66266 , n64615 );
nor ( n66619 , n66617 , n66618 );
xnor ( n66620 , n66619 , n64624 );
and ( n66621 , n66616 , n66620 );
not ( n66622 , n66508 );
and ( n66623 , n66620 , n66622 );
and ( n66624 , n66616 , n66622 );
or ( n66625 , n66621 , n66623 , n66624 );
and ( n66626 , n65698 , n64789 );
and ( n66627 , n65657 , n64787 );
nor ( n66628 , n66626 , n66627 );
xnor ( n66629 , n66628 , n64738 );
and ( n66630 , n66625 , n66629 );
xor ( n66631 , n66509 , n66515 );
xor ( n66632 , n66631 , n66518 );
and ( n66633 , n66629 , n66632 );
and ( n66634 , n66625 , n66632 );
or ( n66635 , n66630 , n66633 , n66634 );
and ( n66636 , n66612 , n66635 );
and ( n66637 , n65453 , n64897 );
and ( n66638 , n65306 , n64895 );
nor ( n66639 , n66637 , n66638 );
xnor ( n66640 , n66639 , n64850 );
and ( n66641 , n66635 , n66640 );
and ( n66642 , n66612 , n66640 );
or ( n66643 , n66636 , n66641 , n66642 );
and ( n66644 , n64906 , n65550 );
and ( n66645 , n64857 , n65548 );
nor ( n66646 , n66644 , n66645 );
xnor ( n66647 , n66646 , n65313 );
and ( n66648 , n66643 , n66647 );
xor ( n66649 , n66270 , n66274 );
xor ( n66650 , n66649 , n66290 );
and ( n66651 , n66647 , n66650 );
and ( n66652 , n66643 , n66650 );
or ( n66653 , n66648 , n66651 , n66652 );
xor ( n66654 , n65873 , n66126 );
xor ( n66655 , n66126 , n66127 );
not ( n66656 , n66655 );
and ( n66657 , n66654 , n66656 );
and ( n66658 , n64619 , n66657 );
not ( n66659 , n66658 );
xnor ( n66660 , n66659 , n66130 );
and ( n66661 , n66653 , n66660 );
xor ( n66662 , n66293 , n66297 );
xor ( n66663 , n66662 , n66302 );
and ( n66664 , n66660 , n66663 );
and ( n66665 , n66653 , n66663 );
or ( n66666 , n66661 , n66664 , n66665 );
xor ( n66667 , n66305 , n66309 );
xor ( n66668 , n66667 , n66314 );
and ( n66669 , n66666 , n66668 );
xor ( n66670 , n66352 , n66356 );
xor ( n66671 , n66670 , n66367 );
and ( n66672 , n66668 , n66671 );
and ( n66673 , n66666 , n66671 );
or ( n66674 , n66669 , n66672 , n66673 );
and ( n66675 , n66596 , n66674 );
xor ( n66676 , n66237 , n66244 );
xor ( n66677 , n66676 , n66247 );
and ( n66678 , n66674 , n66677 );
and ( n66679 , n66596 , n66677 );
or ( n66680 , n66675 , n66678 , n66679 );
xor ( n66681 , n66317 , n66370 );
xor ( n66682 , n66681 , n66383 );
xor ( n66683 , n66478 , n66480 );
xor ( n66684 , n66683 , n66483 );
and ( n66685 , n66682 , n66684 );
xor ( n66686 , n66596 , n66674 );
xor ( n66687 , n66686 , n66677 );
and ( n66688 , n66684 , n66687 );
and ( n66689 , n66682 , n66687 );
or ( n66690 , n66685 , n66688 , n66689 );
and ( n66691 , n66680 , n66690 );
xor ( n66692 , n66486 , n66488 );
xor ( n66693 , n66692 , n66491 );
and ( n66694 , n66690 , n66693 );
and ( n66695 , n66680 , n66693 );
or ( n66696 , n66691 , n66694 , n66695 );
and ( n66697 , n66506 , n66696 );
xor ( n66698 , n66506 , n66696 );
xor ( n66699 , n66680 , n66690 );
xor ( n66700 , n66699 , n66693 );
and ( n66701 , n64611 , n66657 );
and ( n66702 , n64619 , n66655 );
nor ( n66703 , n66701 , n66702 );
xnor ( n66704 , n66703 , n66130 );
and ( n66705 , n64703 , n66016 );
and ( n66706 , n64689 , n66014 );
nor ( n66707 , n66705 , n66706 );
xnor ( n66708 , n66707 , n65650 );
and ( n66709 , n66704 , n66708 );
and ( n66710 , n64798 , n65756 );
and ( n66711 , n64781 , n65754 );
nor ( n66712 , n66710 , n66711 );
xnor ( n66713 , n66712 , n65450 );
and ( n66714 , n66708 , n66713 );
and ( n66715 , n66704 , n66713 );
or ( n66716 , n66709 , n66714 , n66715 );
and ( n66717 , n65363 , n65056 );
and ( n66718 , n65265 , n65054 );
nor ( n66719 , n66717 , n66718 );
xnor ( n66720 , n66719 , n64943 );
xor ( n66721 , n66260 , n66264 );
xor ( n66722 , n66721 , n66267 );
and ( n66723 , n66720 , n66722 );
xor ( n66724 , n66521 , n66525 );
xor ( n66725 , n66724 , n66527 );
and ( n66726 , n66722 , n66725 );
and ( n66727 , n66720 , n66725 );
or ( n66728 , n66723 , n66726 , n66727 );
and ( n66729 , n64662 , n66241 );
and ( n66730 , n64627 , n66239 );
nor ( n66731 , n66729 , n66730 );
xnor ( n66732 , n66731 , n65876 );
and ( n66733 , n66728 , n66732 );
xor ( n66734 , n66530 , n66534 );
xor ( n66735 , n66734 , n66537 );
and ( n66736 , n66732 , n66735 );
and ( n66737 , n66728 , n66735 );
or ( n66738 , n66733 , n66736 , n66737 );
and ( n66739 , n66716 , n66738 );
xor ( n66740 , n66556 , n66560 );
xor ( n66741 , n66740 , n66563 );
and ( n66742 , n66738 , n66741 );
and ( n66743 , n66716 , n66741 );
or ( n66744 , n66739 , n66742 , n66743 );
xor ( n66745 , n66552 , n66566 );
xor ( n66746 , n66745 , n66593 );
and ( n66747 , n66744 , n66746 );
xor ( n66748 , n66470 , n66472 );
xor ( n66749 , n66748 , n66475 );
and ( n66750 , n66746 , n66749 );
and ( n66751 , n66744 , n66749 );
or ( n66752 , n66747 , n66750 , n66751 );
and ( n66753 , n64955 , n65550 );
and ( n66754 , n64950 , n65548 );
nor ( n66755 , n66753 , n66754 );
xnor ( n66756 , n66755 , n65313 );
and ( n66757 , n65135 , n65371 );
and ( n66758 , n65001 , n65369 );
nor ( n66759 , n66757 , n66758 );
xnor ( n66760 , n66759 , n65168 );
and ( n66761 , n66756 , n66760 );
and ( n66762 , n65306 , n65056 );
and ( n66763 , n65363 , n65054 );
nor ( n66764 , n66762 , n66763 );
xnor ( n66765 , n66764 , n64943 );
and ( n66766 , n66760 , n66765 );
and ( n66767 , n66756 , n66765 );
or ( n66768 , n66761 , n66766 , n66767 );
and ( n66769 , n64689 , n66241 );
and ( n66770 , n64662 , n66239 );
nor ( n66771 , n66769 , n66770 );
xnor ( n66772 , n66771 , n65876 );
and ( n66773 , n66768 , n66772 );
and ( n66774 , n64857 , n65756 );
and ( n66775 , n64798 , n65754 );
nor ( n66776 , n66774 , n66775 );
xnor ( n66777 , n66776 , n65450 );
and ( n66778 , n66772 , n66777 );
and ( n66779 , n66768 , n66777 );
or ( n66780 , n66773 , n66778 , n66779 );
buf ( n66781 , n64537 );
and ( n66782 , n66781 , n64617 );
and ( n66783 , n66507 , n64615 );
nor ( n66784 , n66782 , n66783 );
xnor ( n66785 , n66784 , n64624 );
buf ( n66786 , n64538 );
and ( n66787 , n66786 , n64612 );
and ( n66788 , n66785 , n66787 );
and ( n66789 , n66266 , n64652 );
and ( n66790 , n66276 , n64650 );
nor ( n66791 , n66789 , n66790 );
xnor ( n66792 , n66791 , n64609 );
and ( n66793 , n66788 , n66792 );
and ( n66794 , n66507 , n64617 );
and ( n66795 , n66517 , n64615 );
nor ( n66796 , n66794 , n66795 );
xnor ( n66797 , n66796 , n64624 );
and ( n66798 , n66792 , n66797 );
and ( n66799 , n66788 , n66797 );
or ( n66800 , n66793 , n66798 , n66799 );
and ( n66801 , n65453 , n65056 );
and ( n66802 , n65306 , n65054 );
nor ( n66803 , n66801 , n66802 );
xnor ( n66804 , n66803 , n64943 );
and ( n66805 , n66800 , n66804 );
and ( n66806 , n65657 , n64897 );
and ( n66807 , n65443 , n64895 );
nor ( n66808 , n66806 , n66807 );
xnor ( n66809 , n66808 , n64850 );
and ( n66810 , n66804 , n66809 );
and ( n66811 , n66800 , n66809 );
or ( n66812 , n66805 , n66810 , n66811 );
and ( n66813 , n65265 , n65183 );
and ( n66814 , n65175 , n65181 );
nor ( n66815 , n66813 , n66814 );
xnor ( n66816 , n66815 , n64994 );
and ( n66817 , n66812 , n66816 );
xor ( n66818 , n66625 , n66629 );
xor ( n66819 , n66818 , n66632 );
and ( n66820 , n66816 , n66819 );
and ( n66821 , n66812 , n66819 );
or ( n66822 , n66817 , n66820 , n66821 );
and ( n66823 , n64950 , n65550 );
and ( n66824 , n64906 , n65548 );
nor ( n66825 , n66823 , n66824 );
xnor ( n66826 , n66825 , n65313 );
and ( n66827 , n66822 , n66826 );
xor ( n66828 , n66612 , n66635 );
xor ( n66829 , n66828 , n66640 );
and ( n66830 , n66826 , n66829 );
and ( n66831 , n66822 , n66829 );
or ( n66832 , n66827 , n66830 , n66831 );
and ( n66833 , n66780 , n66832 );
and ( n66834 , n64627 , n66657 );
and ( n66835 , n64611 , n66655 );
nor ( n66836 , n66834 , n66835 );
xnor ( n66837 , n66836 , n66130 );
and ( n66838 , n64781 , n66016 );
and ( n66839 , n64703 , n66014 );
nor ( n66840 , n66838 , n66839 );
xnor ( n66841 , n66840 , n65650 );
and ( n66842 , n66837 , n66841 );
xor ( n66843 , n66720 , n66722 );
xor ( n66844 , n66843 , n66725 );
and ( n66845 , n66841 , n66844 );
and ( n66846 , n66837 , n66844 );
or ( n66847 , n66842 , n66845 , n66846 );
and ( n66848 , n66832 , n66847 );
and ( n66849 , n66780 , n66847 );
or ( n66850 , n66833 , n66848 , n66849 );
not ( n66851 , n66511 );
and ( n66852 , n66781 , n64612 );
xnor ( n66853 , n66851 , n66852 );
and ( n66854 , n65935 , n64789 );
and ( n66855 , n65883 , n64787 );
nor ( n66856 , n66854 , n66855 );
xnor ( n66857 , n66856 , n64738 );
and ( n66858 , n66853 , n66857 );
and ( n66859 , n66142 , n64711 );
and ( n66860 , n66137 , n64709 );
nor ( n66861 , n66859 , n66860 );
xnor ( n66862 , n66861 , n64682 );
and ( n66863 , n66857 , n66862 );
and ( n66864 , n66853 , n66862 );
or ( n66865 , n66858 , n66863 , n66864 );
or ( n66866 , n66851 , n66852 );
and ( n66867 , n65883 , n64789 );
and ( n66868 , n65698 , n64787 );
nor ( n66869 , n66867 , n66868 );
xnor ( n66870 , n66869 , n64738 );
xor ( n66871 , n66866 , n66870 );
and ( n66872 , n66137 , n64711 );
and ( n66873 , n65935 , n64709 );
nor ( n66874 , n66872 , n66873 );
xnor ( n66875 , n66874 , n64682 );
xor ( n66876 , n66871 , n66875 );
and ( n66877 , n66865 , n66876 );
xor ( n66878 , n66616 , n66620 );
xor ( n66879 , n66878 , n66622 );
and ( n66880 , n66876 , n66879 );
and ( n66881 , n66865 , n66879 );
or ( n66882 , n66877 , n66880 , n66881 );
and ( n66883 , n64906 , n65756 );
and ( n66884 , n64857 , n65754 );
nor ( n66885 , n66883 , n66884 );
xnor ( n66886 , n66885 , n65450 );
and ( n66887 , n66882 , n66886 );
and ( n66888 , n66866 , n66870 );
and ( n66889 , n66870 , n66875 );
and ( n66890 , n66866 , n66875 );
or ( n66891 , n66888 , n66889 , n66890 );
and ( n66892 , n65443 , n64897 );
and ( n66893 , n65453 , n64895 );
nor ( n66894 , n66892 , n66893 );
xnor ( n66895 , n66894 , n64850 );
xor ( n66896 , n66891 , n66895 );
xor ( n66897 , n66600 , n66604 );
xor ( n66898 , n66897 , n66609 );
xor ( n66899 , n66896 , n66898 );
and ( n66900 , n66886 , n66899 );
and ( n66901 , n66882 , n66899 );
or ( n66902 , n66887 , n66900 , n66901 );
xor ( n66903 , n66127 , n66282 );
xor ( n66904 , n66282 , n66283 );
not ( n66905 , n66904 );
and ( n66906 , n66903 , n66905 );
and ( n66907 , n64619 , n66906 );
not ( n66908 , n66907 );
xnor ( n66909 , n66908 , n66286 );
and ( n66910 , n66902 , n66909 );
and ( n66911 , n66891 , n66895 );
and ( n66912 , n66895 , n66898 );
and ( n66913 , n66891 , n66898 );
or ( n66914 , n66911 , n66912 , n66913 );
and ( n66915 , n65001 , n65371 );
and ( n66916 , n64955 , n65369 );
nor ( n66917 , n66915 , n66916 );
xnor ( n66918 , n66917 , n65168 );
xor ( n66919 , n66914 , n66918 );
and ( n66920 , n65175 , n65183 );
and ( n66921 , n65135 , n65181 );
nor ( n66922 , n66920 , n66921 );
xnor ( n66923 , n66922 , n64994 );
xor ( n66924 , n66919 , n66923 );
and ( n66925 , n66909 , n66924 );
and ( n66926 , n66902 , n66924 );
or ( n66927 , n66910 , n66925 , n66926 );
xor ( n66928 , n66704 , n66708 );
xor ( n66929 , n66928 , n66713 );
and ( n66930 , n66927 , n66929 );
xor ( n66931 , n66728 , n66732 );
xor ( n66932 , n66931 , n66735 );
and ( n66933 , n66929 , n66932 );
and ( n66934 , n66927 , n66932 );
or ( n66935 , n66930 , n66933 , n66934 );
and ( n66936 , n66850 , n66935 );
xor ( n66937 , n66653 , n66660 );
xor ( n66938 , n66937 , n66663 );
and ( n66939 , n66935 , n66938 );
and ( n66940 , n66850 , n66938 );
or ( n66941 , n66936 , n66939 , n66940 );
and ( n66942 , n66914 , n66918 );
and ( n66943 , n66918 , n66923 );
and ( n66944 , n66914 , n66923 );
or ( n66945 , n66942 , n66943 , n66944 );
xor ( n66946 , n66571 , n66575 );
xor ( n66947 , n66946 , n66580 );
and ( n66948 , n66945 , n66947 );
xor ( n66949 , n66643 , n66647 );
xor ( n66950 , n66949 , n66650 );
and ( n66951 , n66947 , n66950 );
and ( n66952 , n66945 , n66950 );
or ( n66953 , n66948 , n66951 , n66952 );
xor ( n66954 , n66540 , n66544 );
xor ( n66955 , n66954 , n66549 );
and ( n66956 , n66953 , n66955 );
xor ( n66957 , n66583 , n66587 );
xor ( n66958 , n66957 , n66590 );
and ( n66959 , n66955 , n66958 );
and ( n66960 , n66953 , n66958 );
or ( n66961 , n66956 , n66959 , n66960 );
and ( n66962 , n66941 , n66961 );
xor ( n66963 , n66666 , n66668 );
xor ( n66964 , n66963 , n66671 );
and ( n66965 , n66961 , n66964 );
and ( n66966 , n66941 , n66964 );
or ( n66967 , n66962 , n66965 , n66966 );
and ( n66968 , n66752 , n66967 );
xor ( n66969 , n66682 , n66684 );
xor ( n66970 , n66969 , n66687 );
and ( n66971 , n66967 , n66970 );
and ( n66972 , n66752 , n66970 );
or ( n66973 , n66968 , n66971 , n66972 );
and ( n66974 , n66700 , n66973 );
xor ( n66975 , n66700 , n66973 );
xor ( n66976 , n66785 , n66787 );
and ( n66977 , n66786 , n64617 );
and ( n66978 , n66781 , n64615 );
nor ( n66979 , n66977 , n66978 );
xnor ( n66980 , n66979 , n64624 );
buf ( n66981 , n64539 );
and ( n66982 , n66981 , n64612 );
and ( n66983 , n66980 , n66982 );
and ( n66984 , n66976 , n66983 );
and ( n66985 , n66276 , n64711 );
and ( n66986 , n66142 , n64709 );
nor ( n66987 , n66985 , n66986 );
xnor ( n66988 , n66987 , n64682 );
and ( n66989 , n66983 , n66988 );
and ( n66990 , n66976 , n66988 );
or ( n66991 , n66984 , n66989 , n66990 );
and ( n66992 , n65443 , n65056 );
and ( n66993 , n65453 , n65054 );
nor ( n66994 , n66992 , n66993 );
xnor ( n66995 , n66994 , n64943 );
and ( n66996 , n66991 , n66995 );
and ( n66997 , n65698 , n64897 );
and ( n66998 , n65657 , n64895 );
nor ( n66999 , n66997 , n66998 );
xnor ( n67000 , n66999 , n64850 );
and ( n67001 , n66995 , n67000 );
and ( n67002 , n66991 , n67000 );
or ( n67003 , n66996 , n67001 , n67002 );
and ( n67004 , n65001 , n65550 );
and ( n67005 , n64955 , n65548 );
nor ( n67006 , n67004 , n67005 );
xnor ( n67007 , n67006 , n65313 );
and ( n67008 , n67003 , n67007 );
and ( n67009 , n65363 , n65183 );
and ( n67010 , n65265 , n65181 );
nor ( n67011 , n67009 , n67010 );
xnor ( n67012 , n67011 , n64994 );
and ( n67013 , n67007 , n67012 );
and ( n67014 , n67003 , n67012 );
or ( n67015 , n67008 , n67013 , n67014 );
and ( n67016 , n64662 , n66657 );
and ( n67017 , n64627 , n66655 );
nor ( n67018 , n67016 , n67017 );
xnor ( n67019 , n67018 , n66130 );
and ( n67020 , n67015 , n67019 );
and ( n67021 , n64798 , n66016 );
and ( n67022 , n64781 , n66014 );
nor ( n67023 , n67021 , n67022 );
xnor ( n67024 , n67023 , n65650 );
and ( n67025 , n67019 , n67024 );
and ( n67026 , n67015 , n67024 );
or ( n67027 , n67020 , n67025 , n67026 );
and ( n67028 , n64611 , n66906 );
and ( n67029 , n64619 , n66904 );
nor ( n67030 , n67028 , n67029 );
xnor ( n67031 , n67030 , n66286 );
and ( n67032 , n64703 , n66241 );
and ( n67033 , n64689 , n66239 );
nor ( n67034 , n67032 , n67033 );
xnor ( n67035 , n67034 , n65876 );
and ( n67036 , n67031 , n67035 );
xor ( n67037 , n66812 , n66816 );
xor ( n67038 , n67037 , n66819 );
and ( n67039 , n67035 , n67038 );
and ( n67040 , n67031 , n67038 );
or ( n67041 , n67036 , n67039 , n67040 );
and ( n67042 , n67027 , n67041 );
xor ( n67043 , n66822 , n66826 );
xor ( n67044 , n67043 , n66829 );
and ( n67045 , n67041 , n67044 );
and ( n67046 , n67027 , n67044 );
or ( n67047 , n67042 , n67045 , n67046 );
xor ( n67048 , n66780 , n66832 );
xor ( n67049 , n67048 , n66847 );
and ( n67050 , n67047 , n67049 );
xor ( n67051 , n66945 , n66947 );
xor ( n67052 , n67051 , n66950 );
and ( n67053 , n67049 , n67052 );
and ( n67054 , n67047 , n67052 );
or ( n67055 , n67050 , n67053 , n67054 );
xor ( n67056 , n66716 , n66738 );
xor ( n67057 , n67056 , n66741 );
and ( n67058 , n67055 , n67057 );
xor ( n67059 , n66953 , n66955 );
xor ( n67060 , n67059 , n66958 );
and ( n67061 , n67057 , n67060 );
and ( n67062 , n67055 , n67060 );
or ( n67063 , n67058 , n67061 , n67062 );
xor ( n67064 , n66744 , n66746 );
xor ( n67065 , n67064 , n66749 );
and ( n67066 , n67063 , n67065 );
xor ( n67067 , n66941 , n66961 );
xor ( n67068 , n67067 , n66964 );
and ( n67069 , n67065 , n67068 );
and ( n67070 , n67063 , n67068 );
or ( n67071 , n67066 , n67069 , n67070 );
xor ( n67072 , n66752 , n66967 );
xor ( n67073 , n67072 , n66970 );
and ( n67074 , n67071 , n67073 );
xor ( n67075 , n67071 , n67073 );
xor ( n67076 , n67063 , n67065 );
xor ( n67077 , n67076 , n67068 );
and ( n67078 , n64955 , n65756 );
and ( n67079 , n64950 , n65754 );
nor ( n67080 , n67078 , n67079 );
xnor ( n67081 , n67080 , n65450 );
and ( n67082 , n65135 , n65550 );
and ( n67083 , n65001 , n65548 );
nor ( n67084 , n67082 , n67083 );
xnor ( n67085 , n67084 , n65313 );
and ( n67086 , n67081 , n67085 );
and ( n67087 , n65306 , n65183 );
and ( n67088 , n65363 , n65181 );
nor ( n67089 , n67087 , n67088 );
xnor ( n67090 , n67089 , n64994 );
and ( n67091 , n67085 , n67090 );
and ( n67092 , n67081 , n67090 );
or ( n67093 , n67086 , n67091 , n67092 );
and ( n67094 , n64627 , n66906 );
and ( n67095 , n64611 , n66904 );
nor ( n67096 , n67094 , n67095 );
xnor ( n67097 , n67096 , n66286 );
and ( n67098 , n67093 , n67097 );
and ( n67099 , n64781 , n66241 );
and ( n67100 , n64703 , n66239 );
nor ( n67101 , n67099 , n67100 );
xnor ( n67102 , n67101 , n65876 );
and ( n67103 , n67097 , n67102 );
and ( n67104 , n67093 , n67102 );
or ( n67105 , n67098 , n67103 , n67104 );
xor ( n67106 , n66980 , n66982 );
and ( n67107 , n66781 , n64652 );
and ( n67108 , n66507 , n64650 );
nor ( n67109 , n67107 , n67108 );
xnor ( n67110 , n67109 , n64609 );
buf ( n67111 , n64540 );
and ( n67112 , n67111 , n64612 );
and ( n67113 , n67110 , n67112 );
and ( n67114 , n67106 , n67113 );
and ( n67115 , n66507 , n64652 );
and ( n67116 , n66517 , n64650 );
nor ( n67117 , n67115 , n67116 );
xnor ( n67118 , n67117 , n64609 );
and ( n67119 , n67113 , n67118 );
and ( n67120 , n67106 , n67118 );
or ( n67121 , n67114 , n67119 , n67120 );
and ( n67122 , n65453 , n65183 );
and ( n67123 , n65306 , n65181 );
nor ( n67124 , n67122 , n67123 );
xnor ( n67125 , n67124 , n64994 );
and ( n67126 , n67121 , n67125 );
and ( n67127 , n65657 , n65056 );
and ( n67128 , n65443 , n65054 );
nor ( n67129 , n67127 , n67128 );
xnor ( n67130 , n67129 , n64943 );
and ( n67131 , n67125 , n67130 );
and ( n67132 , n67121 , n67130 );
or ( n67133 , n67126 , n67131 , n67132 );
and ( n67134 , n65265 , n65371 );
and ( n67135 , n65175 , n65369 );
nor ( n67136 , n67134 , n67135 );
xnor ( n67137 , n67136 , n65168 );
and ( n67138 , n67133 , n67137 );
xor ( n67139 , n66991 , n66995 );
xor ( n67140 , n67139 , n67000 );
and ( n67141 , n67137 , n67140 );
and ( n67142 , n67133 , n67140 );
or ( n67143 , n67138 , n67141 , n67142 );
and ( n67144 , n64689 , n66657 );
and ( n67145 , n64662 , n66655 );
nor ( n67146 , n67144 , n67145 );
xnor ( n67147 , n67146 , n66130 );
and ( n67148 , n67143 , n67147 );
and ( n67149 , n64857 , n66016 );
and ( n67150 , n64798 , n66014 );
nor ( n67151 , n67149 , n67150 );
xnor ( n67152 , n67151 , n65650 );
and ( n67153 , n67147 , n67152 );
and ( n67154 , n67143 , n67152 );
or ( n67155 , n67148 , n67153 , n67154 );
and ( n67156 , n67105 , n67155 );
xor ( n67157 , n66283 , n66510 );
xor ( n67158 , n66510 , n66511 );
not ( n67159 , n67158 );
and ( n67160 , n67157 , n67159 );
and ( n67161 , n64619 , n67160 );
not ( n67162 , n67161 );
xnor ( n67163 , n67162 , n66514 );
and ( n67164 , n64950 , n65756 );
and ( n67165 , n64906 , n65754 );
nor ( n67166 , n67164 , n67165 );
xnor ( n67167 , n67166 , n65450 );
and ( n67168 , n67163 , n67167 );
xor ( n67169 , n66865 , n66876 );
xor ( n67170 , n67169 , n66879 );
and ( n67171 , n67167 , n67170 );
and ( n67172 , n67163 , n67170 );
or ( n67173 , n67168 , n67171 , n67172 );
and ( n67174 , n67155 , n67173 );
and ( n67175 , n67105 , n67173 );
or ( n67176 , n67156 , n67174 , n67175 );
and ( n67177 , n65935 , n64897 );
and ( n67178 , n65883 , n64895 );
nor ( n67179 , n67177 , n67178 );
xnor ( n67180 , n67179 , n64850 );
and ( n67181 , n66142 , n64789 );
and ( n67182 , n66137 , n64787 );
nor ( n67183 , n67181 , n67182 );
xnor ( n67184 , n67183 , n64738 );
and ( n67185 , n67180 , n67184 );
and ( n67186 , n66266 , n64711 );
and ( n67187 , n66276 , n64709 );
nor ( n67188 , n67186 , n67187 );
xnor ( n67189 , n67188 , n64682 );
and ( n67190 , n67184 , n67189 );
and ( n67191 , n67180 , n67189 );
or ( n67192 , n67185 , n67190 , n67191 );
and ( n67193 , n65883 , n64897 );
and ( n67194 , n65698 , n64895 );
nor ( n67195 , n67193 , n67194 );
xnor ( n67196 , n67195 , n64850 );
and ( n67197 , n66137 , n64789 );
and ( n67198 , n65935 , n64787 );
nor ( n67199 , n67197 , n67198 );
xnor ( n67200 , n67199 , n64738 );
xor ( n67201 , n67196 , n67200 );
and ( n67202 , n66517 , n64652 );
and ( n67203 , n66266 , n64650 );
nor ( n67204 , n67202 , n67203 );
xnor ( n67205 , n67204 , n64609 );
xor ( n67206 , n67201 , n67205 );
and ( n67207 , n67192 , n67206 );
xor ( n67208 , n66976 , n66983 );
xor ( n67209 , n67208 , n66988 );
and ( n67210 , n67206 , n67209 );
and ( n67211 , n67192 , n67209 );
or ( n67212 , n67207 , n67210 , n67211 );
and ( n67213 , n64906 , n66016 );
and ( n67214 , n64857 , n66014 );
nor ( n67215 , n67213 , n67214 );
xnor ( n67216 , n67215 , n65650 );
and ( n67217 , n67212 , n67216 );
and ( n67218 , n67196 , n67200 );
and ( n67219 , n67200 , n67205 );
and ( n67220 , n67196 , n67205 );
or ( n67221 , n67218 , n67219 , n67220 );
xor ( n67222 , n66788 , n66792 );
xor ( n67223 , n67222 , n66797 );
xor ( n67224 , n67221 , n67223 );
xor ( n67225 , n66853 , n66857 );
xor ( n67226 , n67225 , n66862 );
xor ( n67227 , n67224 , n67226 );
and ( n67228 , n67216 , n67227 );
and ( n67229 , n67212 , n67227 );
or ( n67230 , n67217 , n67228 , n67229 );
xor ( n67231 , n67003 , n67007 );
xor ( n67232 , n67231 , n67012 );
and ( n67233 , n67230 , n67232 );
and ( n67234 , n67221 , n67223 );
and ( n67235 , n67223 , n67226 );
and ( n67236 , n67221 , n67226 );
or ( n67237 , n67234 , n67235 , n67236 );
and ( n67238 , n65175 , n65371 );
and ( n67239 , n65135 , n65369 );
nor ( n67240 , n67238 , n67239 );
xnor ( n67241 , n67240 , n65168 );
xor ( n67242 , n67237 , n67241 );
xor ( n67243 , n66800 , n66804 );
xor ( n67244 , n67243 , n66809 );
xor ( n67245 , n67242 , n67244 );
and ( n67246 , n67232 , n67245 );
and ( n67247 , n67230 , n67245 );
or ( n67248 , n67233 , n67246 , n67247 );
xor ( n67249 , n67015 , n67019 );
xor ( n67250 , n67249 , n67024 );
and ( n67251 , n67248 , n67250 );
xor ( n67252 , n67031 , n67035 );
xor ( n67253 , n67252 , n67038 );
and ( n67254 , n67250 , n67253 );
and ( n67255 , n67248 , n67253 );
or ( n67256 , n67251 , n67254 , n67255 );
and ( n67257 , n67176 , n67256 );
xor ( n67258 , n66902 , n66909 );
xor ( n67259 , n67258 , n66924 );
and ( n67260 , n67256 , n67259 );
and ( n67261 , n67176 , n67259 );
or ( n67262 , n67257 , n67260 , n67261 );
and ( n67263 , n67237 , n67241 );
and ( n67264 , n67241 , n67244 );
and ( n67265 , n67237 , n67244 );
or ( n67266 , n67263 , n67264 , n67265 );
xor ( n67267 , n66756 , n66760 );
xor ( n67268 , n67267 , n66765 );
and ( n67269 , n67266 , n67268 );
xor ( n67270 , n66882 , n66886 );
xor ( n67271 , n67270 , n66899 );
and ( n67272 , n67268 , n67271 );
and ( n67273 , n67266 , n67271 );
or ( n67274 , n67269 , n67272 , n67273 );
xor ( n67275 , n66768 , n66772 );
xor ( n67276 , n67275 , n66777 );
and ( n67277 , n67274 , n67276 );
xor ( n67278 , n66837 , n66841 );
xor ( n67279 , n67278 , n66844 );
and ( n67280 , n67276 , n67279 );
and ( n67281 , n67274 , n67279 );
or ( n67282 , n67277 , n67280 , n67281 );
and ( n67283 , n67262 , n67282 );
xor ( n67284 , n66927 , n66929 );
xor ( n67285 , n67284 , n66932 );
and ( n67286 , n67282 , n67285 );
and ( n67287 , n67262 , n67285 );
or ( n67288 , n67283 , n67286 , n67287 );
xor ( n67289 , n66850 , n66935 );
xor ( n67290 , n67289 , n66938 );
and ( n67291 , n67288 , n67290 );
xor ( n67292 , n67055 , n67057 );
xor ( n67293 , n67292 , n67060 );
and ( n67294 , n67290 , n67293 );
and ( n67295 , n67288 , n67293 );
or ( n67296 , n67291 , n67294 , n67295 );
and ( n67297 , n67077 , n67296 );
xor ( n67298 , n67077 , n67296 );
xor ( n67299 , n67288 , n67290 );
xor ( n67300 , n67299 , n67293 );
xor ( n67301 , n67110 , n67112 );
buf ( n67302 , n64541 );
and ( n67303 , n67302 , n64617 );
and ( n67304 , n67111 , n64615 );
nor ( n67305 , n67303 , n67304 );
xnor ( n67306 , n67305 , n64624 );
buf ( n67307 , n64542 );
and ( n67308 , n67307 , n64612 );
and ( n67309 , n67306 , n67308 );
and ( n67310 , n67302 , n64612 );
and ( n67311 , n67309 , n67310 );
and ( n67312 , n67301 , n67311 );
and ( n67313 , n66981 , n64617 );
and ( n67314 , n66786 , n64615 );
nor ( n67315 , n67313 , n67314 );
xnor ( n67316 , n67315 , n64624 );
and ( n67317 , n67311 , n67316 );
and ( n67318 , n67301 , n67316 );
or ( n67319 , n67312 , n67317 , n67318 );
and ( n67320 , n65443 , n65183 );
and ( n67321 , n65453 , n65181 );
nor ( n67322 , n67320 , n67321 );
xnor ( n67323 , n67322 , n64994 );
and ( n67324 , n67319 , n67323 );
and ( n67325 , n65698 , n65056 );
and ( n67326 , n65657 , n65054 );
nor ( n67327 , n67325 , n67326 );
xnor ( n67328 , n67327 , n64943 );
and ( n67329 , n67323 , n67328 );
and ( n67330 , n67319 , n67328 );
or ( n67331 , n67324 , n67329 , n67330 );
and ( n67332 , n65001 , n65756 );
and ( n67333 , n64955 , n65754 );
nor ( n67334 , n67332 , n67333 );
xnor ( n67335 , n67334 , n65450 );
and ( n67336 , n67331 , n67335 );
and ( n67337 , n65363 , n65371 );
and ( n67338 , n65265 , n65369 );
nor ( n67339 , n67337 , n67338 );
xnor ( n67340 , n67339 , n65168 );
and ( n67341 , n67335 , n67340 );
and ( n67342 , n67331 , n67340 );
or ( n67343 , n67336 , n67341 , n67342 );
and ( n67344 , n64611 , n67160 );
and ( n67345 , n64619 , n67158 );
nor ( n67346 , n67344 , n67345 );
xnor ( n67347 , n67346 , n66514 );
and ( n67348 , n67343 , n67347 );
and ( n67349 , n64703 , n66657 );
and ( n67350 , n64689 , n66655 );
nor ( n67351 , n67349 , n67350 );
xnor ( n67352 , n67351 , n66130 );
and ( n67353 , n67347 , n67352 );
and ( n67354 , n67343 , n67352 );
or ( n67355 , n67348 , n67353 , n67354 );
and ( n67356 , n64662 , n66906 );
and ( n67357 , n64627 , n66904 );
nor ( n67358 , n67356 , n67357 );
xnor ( n67359 , n67358 , n66286 );
and ( n67360 , n64798 , n66241 );
and ( n67361 , n64781 , n66239 );
nor ( n67362 , n67360 , n67361 );
xnor ( n67363 , n67362 , n65876 );
and ( n67364 , n67359 , n67363 );
xor ( n67365 , n67133 , n67137 );
xor ( n67366 , n67365 , n67140 );
and ( n67367 , n67363 , n67366 );
and ( n67368 , n67359 , n67366 );
or ( n67369 , n67364 , n67367 , n67368 );
and ( n67370 , n67355 , n67369 );
xor ( n67371 , n67163 , n67167 );
xor ( n67372 , n67371 , n67170 );
and ( n67373 , n67369 , n67372 );
and ( n67374 , n67355 , n67372 );
or ( n67375 , n67370 , n67373 , n67374 );
xor ( n67376 , n67105 , n67155 );
xor ( n67377 , n67376 , n67173 );
and ( n67378 , n67375 , n67377 );
xor ( n67379 , n67266 , n67268 );
xor ( n67380 , n67379 , n67271 );
and ( n67381 , n67377 , n67380 );
and ( n67382 , n67375 , n67380 );
or ( n67383 , n67378 , n67381 , n67382 );
xor ( n67384 , n67027 , n67041 );
xor ( n67385 , n67384 , n67044 );
and ( n67386 , n67383 , n67385 );
xor ( n67387 , n67274 , n67276 );
xor ( n67388 , n67387 , n67279 );
and ( n67389 , n67385 , n67388 );
and ( n67390 , n67383 , n67388 );
or ( n67391 , n67386 , n67389 , n67390 );
xor ( n67392 , n67047 , n67049 );
xor ( n67393 , n67392 , n67052 );
and ( n67394 , n67391 , n67393 );
xor ( n67395 , n67262 , n67282 );
xor ( n67396 , n67395 , n67285 );
and ( n67397 , n67393 , n67396 );
and ( n67398 , n67391 , n67396 );
or ( n67399 , n67394 , n67397 , n67398 );
and ( n67400 , n67300 , n67399 );
xor ( n67401 , n67300 , n67399 );
xor ( n67402 , n67391 , n67393 );
xor ( n67403 , n67402 , n67396 );
xor ( n67404 , n67309 , n67310 );
and ( n67405 , n66786 , n64652 );
and ( n67406 , n66781 , n64650 );
nor ( n67407 , n67405 , n67406 );
xnor ( n67408 , n67407 , n64609 );
and ( n67409 , n67404 , n67408 );
and ( n67410 , n67111 , n64617 );
and ( n67411 , n66981 , n64615 );
nor ( n67412 , n67410 , n67411 );
xnor ( n67413 , n67412 , n64624 );
and ( n67414 , n67408 , n67413 );
and ( n67415 , n67404 , n67413 );
or ( n67416 , n67409 , n67414 , n67415 );
and ( n67417 , n66276 , n64789 );
and ( n67418 , n66142 , n64787 );
nor ( n67419 , n67417 , n67418 );
xnor ( n67420 , n67419 , n64738 );
and ( n67421 , n67416 , n67420 );
and ( n67422 , n66517 , n64711 );
and ( n67423 , n66266 , n64709 );
nor ( n67424 , n67422 , n67423 );
xnor ( n67425 , n67424 , n64682 );
and ( n67426 , n67420 , n67425 );
and ( n67427 , n67416 , n67425 );
or ( n67428 , n67421 , n67426 , n67427 );
and ( n67429 , n65883 , n65056 );
and ( n67430 , n65698 , n65054 );
nor ( n67431 , n67429 , n67430 );
xnor ( n67432 , n67431 , n64943 );
and ( n67433 , n66137 , n64897 );
and ( n67434 , n65935 , n64895 );
nor ( n67435 , n67433 , n67434 );
xnor ( n67436 , n67435 , n64850 );
and ( n67437 , n67432 , n67436 );
xor ( n67438 , n67301 , n67311 );
xor ( n67439 , n67438 , n67316 );
and ( n67440 , n67436 , n67439 );
and ( n67441 , n67432 , n67439 );
or ( n67442 , n67437 , n67440 , n67441 );
and ( n67443 , n67428 , n67442 );
xor ( n67444 , n67106 , n67113 );
xor ( n67445 , n67444 , n67118 );
and ( n67446 , n67442 , n67445 );
and ( n67447 , n67428 , n67445 );
or ( n67448 , n67443 , n67446 , n67447 );
and ( n67449 , n65175 , n65550 );
and ( n67450 , n65135 , n65548 );
nor ( n67451 , n67449 , n67450 );
xnor ( n67452 , n67451 , n65313 );
and ( n67453 , n67448 , n67452 );
xor ( n67454 , n67121 , n67125 );
xor ( n67455 , n67454 , n67130 );
and ( n67456 , n67452 , n67455 );
and ( n67457 , n67448 , n67455 );
or ( n67458 , n67453 , n67456 , n67457 );
xor ( n67459 , n67081 , n67085 );
xor ( n67460 , n67459 , n67090 );
and ( n67461 , n67458 , n67460 );
xor ( n67462 , n67212 , n67216 );
xor ( n67463 , n67462 , n67227 );
and ( n67464 , n67460 , n67463 );
and ( n67465 , n67458 , n67463 );
or ( n67466 , n67461 , n67464 , n67465 );
xor ( n67467 , n67093 , n67097 );
xor ( n67468 , n67467 , n67102 );
and ( n67469 , n67466 , n67468 );
xor ( n67470 , n67143 , n67147 );
xor ( n67471 , n67470 , n67152 );
and ( n67472 , n67468 , n67471 );
and ( n67473 , n67466 , n67471 );
or ( n67474 , n67469 , n67472 , n67473 );
xor ( n67475 , n67248 , n67250 );
xor ( n67476 , n67475 , n67253 );
and ( n67477 , n67474 , n67476 );
xor ( n67478 , n67375 , n67377 );
xor ( n67479 , n67478 , n67380 );
and ( n67480 , n67476 , n67479 );
and ( n67481 , n67474 , n67479 );
or ( n67482 , n67477 , n67480 , n67481 );
xor ( n67483 , n67176 , n67256 );
xor ( n67484 , n67483 , n67259 );
and ( n67485 , n67482 , n67484 );
xor ( n67486 , n67383 , n67385 );
xor ( n67487 , n67486 , n67388 );
and ( n67488 , n67484 , n67487 );
and ( n67489 , n67482 , n67487 );
or ( n67490 , n67485 , n67488 , n67489 );
and ( n67491 , n67403 , n67490 );
xor ( n67492 , n67403 , n67490 );
xor ( n67493 , n67482 , n67484 );
xor ( n67494 , n67493 , n67487 );
buf ( n67495 , n64603 );
xor ( n67496 , n66511 , n67495 );
not ( n67497 , n67495 );
and ( n67498 , n67496 , n67497 );
and ( n67499 , n64619 , n67498 );
not ( n67500 , n67499 );
xnor ( n67501 , n67500 , n66511 );
and ( n67502 , n64689 , n66906 );
and ( n67503 , n64662 , n66904 );
nor ( n67504 , n67502 , n67503 );
xnor ( n67505 , n67504 , n66286 );
and ( n67506 , n67501 , n67505 );
and ( n67507 , n64857 , n66241 );
and ( n67508 , n64798 , n66239 );
nor ( n67509 , n67507 , n67508 );
xnor ( n67510 , n67509 , n65876 );
and ( n67511 , n67505 , n67510 );
and ( n67512 , n67501 , n67510 );
or ( n67513 , n67506 , n67511 , n67512 );
and ( n67514 , n64955 , n66016 );
and ( n67515 , n64950 , n66014 );
nor ( n67516 , n67514 , n67515 );
xnor ( n67517 , n67516 , n65650 );
and ( n67518 , n65265 , n65550 );
and ( n67519 , n65175 , n65548 );
nor ( n67520 , n67518 , n67519 );
xnor ( n67521 , n67520 , n65313 );
and ( n67522 , n67517 , n67521 );
and ( n67523 , n65306 , n65371 );
and ( n67524 , n65363 , n65369 );
nor ( n67525 , n67523 , n67524 );
xnor ( n67526 , n67525 , n65168 );
and ( n67527 , n67521 , n67526 );
and ( n67528 , n67517 , n67526 );
or ( n67529 , n67522 , n67527 , n67528 );
and ( n67530 , n64627 , n67160 );
and ( n67531 , n64611 , n67158 );
nor ( n67532 , n67530 , n67531 );
xnor ( n67533 , n67532 , n66514 );
and ( n67534 , n67529 , n67533 );
and ( n67535 , n64781 , n66657 );
and ( n67536 , n64703 , n66655 );
nor ( n67537 , n67535 , n67536 );
xnor ( n67538 , n67537 , n66130 );
and ( n67539 , n67533 , n67538 );
and ( n67540 , n67529 , n67538 );
or ( n67541 , n67534 , n67539 , n67540 );
and ( n67542 , n67513 , n67541 );
xor ( n67543 , n67306 , n67308 );
and ( n67544 , n67307 , n64617 );
and ( n67545 , n67302 , n64615 );
nor ( n67546 , n67544 , n67545 );
xnor ( n67547 , n67546 , n64624 );
buf ( n67548 , n64543 );
and ( n67549 , n67548 , n64612 );
and ( n67550 , n67547 , n67549 );
and ( n67551 , n67543 , n67550 );
and ( n67552 , n66781 , n64711 );
and ( n67553 , n66507 , n64709 );
nor ( n67554 , n67552 , n67553 );
xnor ( n67555 , n67554 , n64682 );
and ( n67556 , n67550 , n67555 );
and ( n67557 , n67543 , n67555 );
or ( n67558 , n67551 , n67556 , n67557 );
and ( n67559 , n66266 , n64789 );
and ( n67560 , n66276 , n64787 );
nor ( n67561 , n67559 , n67560 );
xnor ( n67562 , n67561 , n64738 );
and ( n67563 , n67558 , n67562 );
and ( n67564 , n66507 , n64711 );
and ( n67565 , n66517 , n64709 );
nor ( n67566 , n67564 , n67565 );
xnor ( n67567 , n67566 , n64682 );
and ( n67568 , n67562 , n67567 );
and ( n67569 , n67558 , n67567 );
or ( n67570 , n67563 , n67568 , n67569 );
and ( n67571 , n65453 , n65371 );
and ( n67572 , n65306 , n65369 );
nor ( n67573 , n67571 , n67572 );
xnor ( n67574 , n67573 , n65168 );
and ( n67575 , n67570 , n67574 );
and ( n67576 , n65657 , n65183 );
and ( n67577 , n65443 , n65181 );
nor ( n67578 , n67576 , n67577 );
xnor ( n67579 , n67578 , n64994 );
and ( n67580 , n67574 , n67579 );
and ( n67581 , n67570 , n67579 );
or ( n67582 , n67575 , n67580 , n67581 );
xor ( n67583 , n67180 , n67184 );
xor ( n67584 , n67583 , n67189 );
and ( n67585 , n67582 , n67584 );
xor ( n67586 , n67319 , n67323 );
xor ( n67587 , n67586 , n67328 );
and ( n67588 , n67584 , n67587 );
and ( n67589 , n67582 , n67587 );
or ( n67590 , n67585 , n67588 , n67589 );
and ( n67591 , n64950 , n66016 );
and ( n67592 , n64906 , n66014 );
nor ( n67593 , n67591 , n67592 );
xnor ( n67594 , n67593 , n65650 );
and ( n67595 , n67590 , n67594 );
xor ( n67596 , n67192 , n67206 );
xor ( n67597 , n67596 , n67209 );
and ( n67598 , n67594 , n67597 );
and ( n67599 , n67590 , n67597 );
or ( n67600 , n67595 , n67598 , n67599 );
and ( n67601 , n67541 , n67600 );
and ( n67602 , n67513 , n67600 );
or ( n67603 , n67542 , n67601 , n67602 );
and ( n67604 , n65935 , n65056 );
and ( n67605 , n65883 , n65054 );
nor ( n67606 , n67604 , n67605 );
xnor ( n67607 , n67606 , n64943 );
and ( n67608 , n66142 , n64897 );
and ( n67609 , n66137 , n64895 );
nor ( n67610 , n67608 , n67609 );
xnor ( n67611 , n67610 , n64850 );
and ( n67612 , n67607 , n67611 );
xor ( n67613 , n67404 , n67408 );
xor ( n67614 , n67613 , n67413 );
and ( n67615 , n67611 , n67614 );
and ( n67616 , n67607 , n67614 );
or ( n67617 , n67612 , n67615 , n67616 );
xor ( n67618 , n67416 , n67420 );
xor ( n67619 , n67618 , n67425 );
and ( n67620 , n67617 , n67619 );
xor ( n67621 , n67432 , n67436 );
xor ( n67622 , n67621 , n67439 );
and ( n67623 , n67619 , n67622 );
and ( n67624 , n67617 , n67622 );
or ( n67625 , n67620 , n67623 , n67624 );
and ( n67626 , n65135 , n65756 );
and ( n67627 , n65001 , n65754 );
nor ( n67628 , n67626 , n67627 );
xnor ( n67629 , n67628 , n65450 );
and ( n67630 , n67625 , n67629 );
xor ( n67631 , n67428 , n67442 );
xor ( n67632 , n67631 , n67445 );
and ( n67633 , n67629 , n67632 );
and ( n67634 , n67625 , n67632 );
or ( n67635 , n67630 , n67633 , n67634 );
xor ( n67636 , n67331 , n67335 );
xor ( n67637 , n67636 , n67340 );
and ( n67638 , n67635 , n67637 );
xor ( n67639 , n67448 , n67452 );
xor ( n67640 , n67639 , n67455 );
and ( n67641 , n67637 , n67640 );
and ( n67642 , n67635 , n67640 );
or ( n67643 , n67638 , n67641 , n67642 );
xor ( n67644 , n67343 , n67347 );
xor ( n67645 , n67644 , n67352 );
and ( n67646 , n67643 , n67645 );
xor ( n67647 , n67359 , n67363 );
xor ( n67648 , n67647 , n67366 );
and ( n67649 , n67645 , n67648 );
and ( n67650 , n67643 , n67648 );
or ( n67651 , n67646 , n67649 , n67650 );
and ( n67652 , n67603 , n67651 );
xor ( n67653 , n67230 , n67232 );
xor ( n67654 , n67653 , n67245 );
and ( n67655 , n67651 , n67654 );
and ( n67656 , n67603 , n67654 );
or ( n67657 , n67652 , n67655 , n67656 );
xor ( n67658 , n67466 , n67468 );
xor ( n67659 , n67658 , n67471 );
xor ( n67660 , n67355 , n67369 );
xor ( n67661 , n67660 , n67372 );
and ( n67662 , n67659 , n67661 );
xor ( n67663 , n67603 , n67651 );
xor ( n67664 , n67663 , n67654 );
and ( n67665 , n67661 , n67664 );
and ( n67666 , n67659 , n67664 );
or ( n67667 , n67662 , n67665 , n67666 );
and ( n67668 , n67657 , n67667 );
xor ( n67669 , n67474 , n67476 );
xor ( n67670 , n67669 , n67479 );
and ( n67671 , n67667 , n67670 );
and ( n67672 , n67657 , n67670 );
or ( n67673 , n67668 , n67671 , n67672 );
and ( n67674 , n67494 , n67673 );
xor ( n67675 , n67494 , n67673 );
xor ( n67676 , n67657 , n67667 );
xor ( n67677 , n67676 , n67670 );
and ( n67678 , n64703 , n66906 );
and ( n67679 , n64689 , n66904 );
nor ( n67680 , n67678 , n67679 );
xnor ( n67681 , n67680 , n66286 );
and ( n67682 , n64798 , n66657 );
and ( n67683 , n64781 , n66655 );
nor ( n67684 , n67682 , n67683 );
xnor ( n67685 , n67684 , n66130 );
and ( n67686 , n67681 , n67685 );
and ( n67687 , n64906 , n66241 );
and ( n67688 , n64857 , n66239 );
nor ( n67689 , n67687 , n67688 );
xnor ( n67690 , n67689 , n65876 );
and ( n67691 , n67685 , n67690 );
and ( n67692 , n67681 , n67690 );
or ( n67693 , n67686 , n67691 , n67692 );
and ( n67694 , n64611 , n67498 );
and ( n67695 , n64619 , n67495 );
nor ( n67696 , n67694 , n67695 );
xnor ( n67697 , n67696 , n66511 );
and ( n67698 , n64662 , n67160 );
and ( n67699 , n64627 , n67158 );
nor ( n67700 , n67698 , n67699 );
xnor ( n67701 , n67700 , n66514 );
and ( n67702 , n67697 , n67701 );
xor ( n67703 , n67582 , n67584 );
xor ( n67704 , n67703 , n67587 );
and ( n67705 , n67701 , n67704 );
and ( n67706 , n67697 , n67704 );
or ( n67707 , n67702 , n67705 , n67706 );
and ( n67708 , n67693 , n67707 );
xor ( n67709 , n67590 , n67594 );
xor ( n67710 , n67709 , n67597 );
and ( n67711 , n67707 , n67710 );
and ( n67712 , n67693 , n67710 );
or ( n67713 , n67708 , n67711 , n67712 );
xor ( n67714 , n67513 , n67541 );
xor ( n67715 , n67714 , n67600 );
and ( n67716 , n67713 , n67715 );
xor ( n67717 , n67458 , n67460 );
xor ( n67718 , n67717 , n67463 );
and ( n67719 , n67715 , n67718 );
and ( n67720 , n67713 , n67718 );
or ( n67721 , n67716 , n67719 , n67720 );
xor ( n67722 , n67547 , n67549 );
and ( n67723 , n67302 , n64652 );
and ( n67724 , n67111 , n64650 );
nor ( n67725 , n67723 , n67724 );
xnor ( n67726 , n67725 , n64609 );
buf ( n67727 , n64544 );
and ( n67728 , n67727 , n64612 );
and ( n67729 , n67726 , n67728 );
and ( n67730 , n67722 , n67729 );
and ( n67731 , n67111 , n64652 );
and ( n67732 , n66981 , n64650 );
nor ( n67733 , n67731 , n67732 );
xnor ( n67734 , n67733 , n64609 );
and ( n67735 , n67729 , n67734 );
and ( n67736 , n67722 , n67734 );
or ( n67737 , n67730 , n67735 , n67736 );
and ( n67738 , n66276 , n64897 );
and ( n67739 , n66142 , n64895 );
nor ( n67740 , n67738 , n67739 );
xnor ( n67741 , n67740 , n64850 );
and ( n67742 , n67737 , n67741 );
and ( n67743 , n66981 , n64652 );
and ( n67744 , n66786 , n64650 );
nor ( n67745 , n67743 , n67744 );
xnor ( n67746 , n67745 , n64609 );
and ( n67747 , n67741 , n67746 );
and ( n67748 , n67737 , n67746 );
or ( n67749 , n67742 , n67747 , n67748 );
and ( n67750 , n65443 , n65371 );
and ( n67751 , n65453 , n65369 );
nor ( n67752 , n67750 , n67751 );
xnor ( n67753 , n67752 , n65168 );
and ( n67754 , n67749 , n67753 );
and ( n67755 , n65698 , n65183 );
and ( n67756 , n65657 , n65181 );
nor ( n67757 , n67755 , n67756 );
xnor ( n67758 , n67757 , n64994 );
and ( n67759 , n67753 , n67758 );
and ( n67760 , n67749 , n67758 );
or ( n67761 , n67754 , n67759 , n67760 );
and ( n67762 , n65001 , n66016 );
and ( n67763 , n64955 , n66014 );
nor ( n67764 , n67762 , n67763 );
xnor ( n67765 , n67764 , n65650 );
and ( n67766 , n67761 , n67765 );
and ( n67767 , n65363 , n65550 );
and ( n67768 , n65265 , n65548 );
nor ( n67769 , n67767 , n67768 );
xnor ( n67770 , n67769 , n65313 );
and ( n67771 , n67765 , n67770 );
and ( n67772 , n67761 , n67770 );
or ( n67773 , n67766 , n67771 , n67772 );
and ( n67774 , n65175 , n65756 );
and ( n67775 , n65135 , n65754 );
nor ( n67776 , n67774 , n67775 );
xnor ( n67777 , n67776 , n65450 );
xor ( n67778 , n67570 , n67574 );
xor ( n67779 , n67778 , n67579 );
and ( n67780 , n67777 , n67779 );
xor ( n67781 , n67617 , n67619 );
xor ( n67782 , n67781 , n67622 );
and ( n67783 , n67779 , n67782 );
and ( n67784 , n67777 , n67782 );
or ( n67785 , n67780 , n67783 , n67784 );
and ( n67786 , n67773 , n67785 );
xor ( n67787 , n67517 , n67521 );
xor ( n67788 , n67787 , n67526 );
and ( n67789 , n67785 , n67788 );
and ( n67790 , n67773 , n67788 );
or ( n67791 , n67786 , n67789 , n67790 );
xor ( n67792 , n67501 , n67505 );
xor ( n67793 , n67792 , n67510 );
and ( n67794 , n67791 , n67793 );
xor ( n67795 , n67529 , n67533 );
xor ( n67796 , n67795 , n67538 );
and ( n67797 , n67793 , n67796 );
and ( n67798 , n67791 , n67796 );
or ( n67799 , n67794 , n67797 , n67798 );
and ( n67800 , n64955 , n66241 );
and ( n67801 , n64950 , n66239 );
nor ( n67802 , n67800 , n67801 );
xnor ( n67803 , n67802 , n65876 );
and ( n67804 , n65135 , n66016 );
and ( n67805 , n65001 , n66014 );
nor ( n67806 , n67804 , n67805 );
xnor ( n67807 , n67806 , n65650 );
and ( n67808 , n67803 , n67807 );
and ( n67809 , n65306 , n65550 );
and ( n67810 , n65363 , n65548 );
nor ( n67811 , n67809 , n67810 );
xnor ( n67812 , n67811 , n65313 );
and ( n67813 , n67807 , n67812 );
and ( n67814 , n67803 , n67812 );
or ( n67815 , n67808 , n67813 , n67814 );
and ( n67816 , n64627 , n67498 );
and ( n67817 , n64611 , n67495 );
nor ( n67818 , n67816 , n67817 );
xnor ( n67819 , n67818 , n66511 );
and ( n67820 , n67815 , n67819 );
and ( n67821 , n64857 , n66657 );
and ( n67822 , n64798 , n66655 );
nor ( n67823 , n67821 , n67822 );
xnor ( n67824 , n67823 , n66130 );
and ( n67825 , n67819 , n67824 );
and ( n67826 , n67815 , n67824 );
or ( n67827 , n67820 , n67825 , n67826 );
xor ( n67828 , n67726 , n67728 );
and ( n67829 , n67727 , n64617 );
and ( n67830 , n67548 , n64615 );
nor ( n67831 , n67829 , n67830 );
xnor ( n67832 , n67831 , n64624 );
buf ( n67833 , n64545 );
and ( n67834 , n67833 , n64612 );
and ( n67835 , n67832 , n67834 );
and ( n67836 , n67828 , n67835 );
and ( n67837 , n67548 , n64617 );
and ( n67838 , n67307 , n64615 );
nor ( n67839 , n67837 , n67838 );
xnor ( n67840 , n67839 , n64624 );
and ( n67841 , n67835 , n67840 );
and ( n67842 , n67828 , n67840 );
or ( n67843 , n67836 , n67841 , n67842 );
and ( n67844 , n66507 , n64789 );
and ( n67845 , n66517 , n64787 );
nor ( n67846 , n67844 , n67845 );
xnor ( n67847 , n67846 , n64738 );
and ( n67848 , n67843 , n67847 );
and ( n67849 , n66786 , n64711 );
and ( n67850 , n66781 , n64709 );
nor ( n67851 , n67849 , n67850 );
xnor ( n67852 , n67851 , n64682 );
and ( n67853 , n67847 , n67852 );
and ( n67854 , n67843 , n67852 );
or ( n67855 , n67848 , n67853 , n67854 );
and ( n67856 , n65453 , n65550 );
and ( n67857 , n65306 , n65548 );
nor ( n67858 , n67856 , n67857 );
xnor ( n67859 , n67858 , n65313 );
and ( n67860 , n67855 , n67859 );
and ( n67861 , n65883 , n65183 );
and ( n67862 , n65698 , n65181 );
nor ( n67863 , n67861 , n67862 );
xnor ( n67864 , n67863 , n64994 );
and ( n67865 , n67859 , n67864 );
and ( n67866 , n67855 , n67864 );
or ( n67867 , n67860 , n67865 , n67866 );
xor ( n67868 , n67832 , n67834 );
and ( n67869 , n67833 , n64617 );
and ( n67870 , n67727 , n64615 );
nor ( n67871 , n67869 , n67870 );
xnor ( n67872 , n67871 , n64624 );
buf ( n67873 , n64546 );
and ( n67874 , n67873 , n64612 );
and ( n67875 , n67872 , n67874 );
and ( n67876 , n67868 , n67875 );
and ( n67877 , n67307 , n64652 );
and ( n67878 , n67302 , n64650 );
nor ( n67879 , n67877 , n67878 );
xnor ( n67880 , n67879 , n64609 );
and ( n67881 , n67875 , n67880 );
and ( n67882 , n67868 , n67880 );
or ( n67883 , n67876 , n67881 , n67882 );
and ( n67884 , n66781 , n64789 );
and ( n67885 , n66507 , n64787 );
nor ( n67886 , n67884 , n67885 );
xnor ( n67887 , n67886 , n64738 );
and ( n67888 , n67883 , n67887 );
and ( n67889 , n66981 , n64711 );
and ( n67890 , n66786 , n64709 );
nor ( n67891 , n67889 , n67890 );
xnor ( n67892 , n67891 , n64682 );
and ( n67893 , n67887 , n67892 );
and ( n67894 , n67883 , n67892 );
or ( n67895 , n67888 , n67893 , n67894 );
and ( n67896 , n66266 , n64897 );
and ( n67897 , n66276 , n64895 );
nor ( n67898 , n67896 , n67897 );
xnor ( n67899 , n67898 , n64850 );
and ( n67900 , n67895 , n67899 );
xor ( n67901 , n67722 , n67729 );
xor ( n67902 , n67901 , n67734 );
and ( n67903 , n67899 , n67902 );
and ( n67904 , n67895 , n67902 );
or ( n67905 , n67900 , n67903 , n67904 );
and ( n67906 , n65657 , n65371 );
and ( n67907 , n65443 , n65369 );
nor ( n67908 , n67906 , n67907 );
xnor ( n67909 , n67908 , n65168 );
and ( n67910 , n67905 , n67909 );
xor ( n67911 , n67737 , n67741 );
xor ( n67912 , n67911 , n67746 );
and ( n67913 , n67909 , n67912 );
and ( n67914 , n67905 , n67912 );
or ( n67915 , n67910 , n67913 , n67914 );
and ( n67916 , n67867 , n67915 );
xor ( n67917 , n67749 , n67753 );
xor ( n67918 , n67917 , n67758 );
and ( n67919 , n67915 , n67918 );
and ( n67920 , n67867 , n67918 );
or ( n67921 , n67916 , n67919 , n67920 );
and ( n67922 , n66137 , n65056 );
and ( n67923 , n65935 , n65054 );
nor ( n67924 , n67922 , n67923 );
xnor ( n67925 , n67924 , n64943 );
and ( n67926 , n66517 , n64789 );
and ( n67927 , n66266 , n64787 );
nor ( n67928 , n67926 , n67927 );
xnor ( n67929 , n67928 , n64738 );
and ( n67930 , n67925 , n67929 );
xor ( n67931 , n67543 , n67550 );
xor ( n67932 , n67931 , n67555 );
and ( n67933 , n67929 , n67932 );
and ( n67934 , n67925 , n67932 );
or ( n67935 , n67930 , n67933 , n67934 );
xor ( n67936 , n67558 , n67562 );
xor ( n67937 , n67936 , n67567 );
and ( n67938 , n67935 , n67937 );
xor ( n67939 , n67607 , n67611 );
xor ( n67940 , n67939 , n67614 );
and ( n67941 , n67937 , n67940 );
and ( n67942 , n67935 , n67940 );
or ( n67943 , n67938 , n67941 , n67942 );
and ( n67944 , n67921 , n67943 );
and ( n67945 , n64950 , n66241 );
and ( n67946 , n64906 , n66239 );
nor ( n67947 , n67945 , n67946 );
xnor ( n67948 , n67947 , n65876 );
and ( n67949 , n67943 , n67948 );
and ( n67950 , n67921 , n67948 );
or ( n67951 , n67944 , n67949 , n67950 );
and ( n67952 , n67827 , n67951 );
xor ( n67953 , n67625 , n67629 );
xor ( n67954 , n67953 , n67632 );
and ( n67955 , n67951 , n67954 );
and ( n67956 , n67827 , n67954 );
or ( n67957 , n67952 , n67955 , n67956 );
and ( n67958 , n64906 , n66657 );
and ( n67959 , n64857 , n66655 );
nor ( n67960 , n67958 , n67959 );
xnor ( n67961 , n67960 , n66130 );
and ( n67962 , n65265 , n65756 );
and ( n67963 , n65175 , n65754 );
nor ( n67964 , n67962 , n67963 );
xnor ( n67965 , n67964 , n65450 );
and ( n67966 , n67961 , n67965 );
xor ( n67967 , n67935 , n67937 );
xor ( n67968 , n67967 , n67940 );
and ( n67969 , n67965 , n67968 );
and ( n67970 , n67961 , n67968 );
or ( n67971 , n67966 , n67969 , n67970 );
and ( n67972 , n64689 , n67160 );
and ( n67973 , n64662 , n67158 );
nor ( n67974 , n67972 , n67973 );
xnor ( n67975 , n67974 , n66514 );
and ( n67976 , n67971 , n67975 );
and ( n67977 , n64781 , n66906 );
and ( n67978 , n64703 , n66904 );
nor ( n67979 , n67977 , n67978 );
xnor ( n67980 , n67979 , n66286 );
and ( n67981 , n67975 , n67980 );
and ( n67982 , n67971 , n67980 );
or ( n67983 , n67976 , n67981 , n67982 );
xor ( n67984 , n67681 , n67685 );
xor ( n67985 , n67984 , n67690 );
and ( n67986 , n67983 , n67985 );
xor ( n67987 , n67697 , n67701 );
xor ( n67988 , n67987 , n67704 );
and ( n67989 , n67985 , n67988 );
and ( n67990 , n67983 , n67988 );
or ( n67991 , n67986 , n67989 , n67990 );
and ( n67992 , n67957 , n67991 );
xor ( n67993 , n67635 , n67637 );
xor ( n67994 , n67993 , n67640 );
and ( n67995 , n67991 , n67994 );
and ( n67996 , n67957 , n67994 );
or ( n67997 , n67992 , n67995 , n67996 );
and ( n67998 , n67799 , n67997 );
xor ( n67999 , n67643 , n67645 );
xor ( n68000 , n67999 , n67648 );
and ( n68001 , n67997 , n68000 );
and ( n68002 , n67799 , n68000 );
or ( n68003 , n67998 , n68001 , n68002 );
and ( n68004 , n67721 , n68003 );
xor ( n68005 , n67659 , n67661 );
xor ( n68006 , n68005 , n67664 );
and ( n68007 , n68003 , n68006 );
and ( n68008 , n67721 , n68006 );
or ( n68009 , n68004 , n68007 , n68008 );
and ( n68010 , n67677 , n68009 );
xor ( n68011 , n67677 , n68009 );
xor ( n68012 , n67721 , n68003 );
xor ( n68013 , n68012 , n68006 );
xor ( n68014 , n67761 , n67765 );
xor ( n68015 , n68014 , n67770 );
xor ( n68016 , n67921 , n67943 );
xor ( n68017 , n68016 , n67948 );
and ( n68018 , n68015 , n68017 );
xor ( n68019 , n67777 , n67779 );
xor ( n68020 , n68019 , n67782 );
and ( n68021 , n68017 , n68020 );
and ( n68022 , n68015 , n68020 );
or ( n68023 , n68018 , n68021 , n68022 );
xor ( n68024 , n67773 , n67785 );
xor ( n68025 , n68024 , n67788 );
and ( n68026 , n68023 , n68025 );
xor ( n68027 , n67827 , n67951 );
xor ( n68028 , n68027 , n67954 );
and ( n68029 , n68025 , n68028 );
and ( n68030 , n68023 , n68028 );
or ( n68031 , n68026 , n68029 , n68030 );
xor ( n68032 , n67791 , n67793 );
xor ( n68033 , n68032 , n67796 );
and ( n68034 , n68031 , n68033 );
xor ( n68035 , n67693 , n67707 );
xor ( n68036 , n68035 , n67710 );
and ( n68037 , n68033 , n68036 );
and ( n68038 , n68031 , n68036 );
or ( n68039 , n68034 , n68037 , n68038 );
xor ( n68040 , n67713 , n67715 );
xor ( n68041 , n68040 , n67718 );
and ( n68042 , n68039 , n68041 );
xor ( n68043 , n67799 , n67997 );
xor ( n68044 , n68043 , n68000 );
and ( n68045 , n68041 , n68044 );
and ( n68046 , n68039 , n68044 );
or ( n68047 , n68042 , n68045 , n68046 );
and ( n68048 , n68013 , n68047 );
xor ( n68049 , n68013 , n68047 );
xor ( n68050 , n68039 , n68041 );
xor ( n68051 , n68050 , n68044 );
and ( n68052 , n65001 , n66241 );
and ( n68053 , n64955 , n66239 );
nor ( n68054 , n68052 , n68053 );
xnor ( n68055 , n68054 , n65876 );
xor ( n68056 , n67855 , n67859 );
xor ( n68057 , n68056 , n67864 );
and ( n68058 , n68055 , n68057 );
xor ( n68059 , n67905 , n67909 );
xor ( n68060 , n68059 , n67912 );
and ( n68061 , n68057 , n68060 );
and ( n68062 , n68055 , n68060 );
or ( n68063 , n68058 , n68061 , n68062 );
and ( n68064 , n64662 , n67498 );
and ( n68065 , n64627 , n67495 );
nor ( n68066 , n68064 , n68065 );
xnor ( n68067 , n68066 , n66511 );
and ( n68068 , n68063 , n68067 );
and ( n68069 , n64798 , n66906 );
and ( n68070 , n64781 , n66904 );
nor ( n68071 , n68069 , n68070 );
xnor ( n68072 , n68071 , n66286 );
and ( n68073 , n68067 , n68072 );
and ( n68074 , n68063 , n68072 );
or ( n68075 , n68068 , n68073 , n68074 );
and ( n68076 , n65698 , n65371 );
and ( n68077 , n65657 , n65369 );
nor ( n68078 , n68076 , n68077 );
xnor ( n68079 , n68078 , n65168 );
and ( n68080 , n65935 , n65183 );
and ( n68081 , n65883 , n65181 );
nor ( n68082 , n68080 , n68081 );
xnor ( n68083 , n68082 , n64994 );
and ( n68084 , n68079 , n68083 );
and ( n68085 , n66142 , n65056 );
and ( n68086 , n66137 , n65054 );
nor ( n68087 , n68085 , n68086 );
xnor ( n68088 , n68087 , n64943 );
and ( n68089 , n68083 , n68088 );
and ( n68090 , n68079 , n68088 );
or ( n68091 , n68084 , n68089 , n68090 );
and ( n68092 , n66276 , n65056 );
and ( n68093 , n66142 , n65054 );
nor ( n68094 , n68092 , n68093 );
xnor ( n68095 , n68094 , n64943 );
and ( n68096 , n66517 , n64897 );
and ( n68097 , n66266 , n64895 );
nor ( n68098 , n68096 , n68097 );
xnor ( n68099 , n68098 , n64850 );
and ( n68100 , n68095 , n68099 );
xor ( n68101 , n67828 , n67835 );
xor ( n68102 , n68101 , n67840 );
and ( n68103 , n68099 , n68102 );
and ( n68104 , n68095 , n68102 );
or ( n68105 , n68100 , n68103 , n68104 );
and ( n68106 , n65443 , n65550 );
and ( n68107 , n65453 , n65548 );
nor ( n68108 , n68106 , n68107 );
xnor ( n68109 , n68108 , n65313 );
and ( n68110 , n68105 , n68109 );
xor ( n68111 , n67843 , n67847 );
xor ( n68112 , n68111 , n67852 );
and ( n68113 , n68109 , n68112 );
and ( n68114 , n68105 , n68112 );
or ( n68115 , n68110 , n68113 , n68114 );
and ( n68116 , n68091 , n68115 );
xor ( n68117 , n67925 , n67929 );
xor ( n68118 , n68117 , n67932 );
and ( n68119 , n68115 , n68118 );
and ( n68120 , n68091 , n68118 );
or ( n68121 , n68116 , n68119 , n68120 );
and ( n68122 , n64703 , n67160 );
and ( n68123 , n64689 , n67158 );
nor ( n68124 , n68122 , n68123 );
xnor ( n68125 , n68124 , n66514 );
and ( n68126 , n68121 , n68125 );
xor ( n68127 , n67867 , n67915 );
xor ( n68128 , n68127 , n67918 );
and ( n68129 , n68125 , n68128 );
and ( n68130 , n68121 , n68128 );
or ( n68131 , n68126 , n68129 , n68130 );
and ( n68132 , n68075 , n68131 );
xor ( n68133 , n67971 , n67975 );
xor ( n68134 , n68133 , n67980 );
and ( n68135 , n68131 , n68134 );
and ( n68136 , n68075 , n68134 );
or ( n68137 , n68132 , n68135 , n68136 );
and ( n68138 , n64950 , n66657 );
and ( n68139 , n64906 , n66655 );
nor ( n68140 , n68138 , n68139 );
xnor ( n68141 , n68140 , n66130 );
and ( n68142 , n65175 , n66016 );
and ( n68143 , n65135 , n66014 );
nor ( n68144 , n68142 , n68143 );
xnor ( n68145 , n68144 , n65650 );
and ( n68146 , n68141 , n68145 );
and ( n68147 , n65363 , n65756 );
and ( n68148 , n65265 , n65754 );
nor ( n68149 , n68147 , n68148 );
xnor ( n68150 , n68149 , n65450 );
and ( n68151 , n68145 , n68150 );
and ( n68152 , n68141 , n68150 );
or ( n68153 , n68146 , n68151 , n68152 );
xor ( n68154 , n67803 , n67807 );
xor ( n68155 , n68154 , n67812 );
and ( n68156 , n68153 , n68155 );
xor ( n68157 , n67961 , n67965 );
xor ( n68158 , n68157 , n67968 );
and ( n68159 , n68155 , n68158 );
and ( n68160 , n68153 , n68158 );
or ( n68161 , n68156 , n68159 , n68160 );
xor ( n68162 , n67815 , n67819 );
xor ( n68163 , n68162 , n67824 );
and ( n68164 , n68161 , n68163 );
xor ( n68165 , n68015 , n68017 );
xor ( n68166 , n68165 , n68020 );
and ( n68167 , n68163 , n68166 );
and ( n68168 , n68161 , n68166 );
or ( n68169 , n68164 , n68167 , n68168 );
and ( n68170 , n68137 , n68169 );
xor ( n68171 , n67983 , n67985 );
xor ( n68172 , n68171 , n67988 );
and ( n68173 , n68169 , n68172 );
and ( n68174 , n68137 , n68172 );
or ( n68175 , n68170 , n68173 , n68174 );
xor ( n68176 , n67957 , n67991 );
xor ( n68177 , n68176 , n67994 );
and ( n68178 , n68175 , n68177 );
xor ( n68179 , n68031 , n68033 );
xor ( n68180 , n68179 , n68036 );
and ( n68181 , n68177 , n68180 );
and ( n68182 , n68175 , n68180 );
or ( n68183 , n68178 , n68181 , n68182 );
and ( n68184 , n68051 , n68183 );
xor ( n68185 , n68051 , n68183 );
xor ( n68186 , n68175 , n68177 );
xor ( n68187 , n68186 , n68180 );
and ( n68188 , n67873 , n64617 );
and ( n68189 , n67833 , n64615 );
nor ( n68190 , n68188 , n68189 );
xnor ( n68191 , n68190 , n64624 );
buf ( n68192 , n64547 );
and ( n68193 , n68192 , n64612 );
xor ( n68194 , n68191 , n68193 );
and ( n68195 , n67833 , n64652 );
and ( n68196 , n67727 , n64650 );
nor ( n68197 , n68195 , n68196 );
xnor ( n68198 , n68197 , n64609 );
buf ( n68199 , n64548 );
and ( n68200 , n68199 , n64612 );
and ( n68201 , n68198 , n68200 );
and ( n68202 , n68194 , n68201 );
and ( n68203 , n67727 , n64652 );
and ( n68204 , n67548 , n64650 );
nor ( n68205 , n68203 , n68204 );
xnor ( n68206 , n68205 , n64609 );
and ( n68207 , n68201 , n68206 );
and ( n68208 , n68194 , n68206 );
or ( n68209 , n68202 , n68207 , n68208 );
and ( n68210 , n67548 , n64652 );
and ( n68211 , n67307 , n64650 );
nor ( n68212 , n68210 , n68211 );
xnor ( n68213 , n68212 , n64609 );
and ( n68214 , n68209 , n68213 );
xor ( n68215 , n67872 , n67874 );
and ( n68216 , n68191 , n68193 );
xor ( n68217 , n68215 , n68216 );
and ( n68218 , n67302 , n64711 );
and ( n68219 , n67111 , n64709 );
nor ( n68220 , n68218 , n68219 );
xnor ( n68221 , n68220 , n64682 );
xor ( n68222 , n68217 , n68221 );
and ( n68223 , n68213 , n68222 );
and ( n68224 , n68209 , n68222 );
or ( n68225 , n68214 , n68223 , n68224 );
and ( n68226 , n66507 , n64897 );
and ( n68227 , n66517 , n64895 );
nor ( n68228 , n68226 , n68227 );
xnor ( n68229 , n68228 , n64850 );
and ( n68230 , n68225 , n68229 );
xor ( n68231 , n67868 , n67875 );
xor ( n68232 , n68231 , n67880 );
and ( n68233 , n68229 , n68232 );
and ( n68234 , n68225 , n68232 );
or ( n68235 , n68230 , n68233 , n68234 );
and ( n68236 , n65657 , n65550 );
and ( n68237 , n65443 , n65548 );
nor ( n68238 , n68236 , n68237 );
xnor ( n68239 , n68238 , n65313 );
and ( n68240 , n68235 , n68239 );
xor ( n68241 , n67883 , n67887 );
xor ( n68242 , n68241 , n67892 );
and ( n68243 , n68239 , n68242 );
and ( n68244 , n68235 , n68242 );
or ( n68245 , n68240 , n68243 , n68244 );
and ( n68246 , n64955 , n66657 );
and ( n68247 , n64950 , n66655 );
nor ( n68248 , n68246 , n68247 );
xnor ( n68249 , n68248 , n66130 );
and ( n68250 , n68245 , n68249 );
xor ( n68251 , n68105 , n68109 );
xor ( n68252 , n68251 , n68112 );
and ( n68253 , n68249 , n68252 );
and ( n68254 , n68245 , n68252 );
or ( n68255 , n68250 , n68253 , n68254 );
and ( n68256 , n64689 , n67498 );
and ( n68257 , n64662 , n67495 );
nor ( n68258 , n68256 , n68257 );
xnor ( n68259 , n68258 , n66511 );
and ( n68260 , n68255 , n68259 );
and ( n68261 , n64857 , n66906 );
and ( n68262 , n64798 , n66904 );
nor ( n68263 , n68261 , n68262 );
xnor ( n68264 , n68263 , n66286 );
and ( n68265 , n68259 , n68264 );
and ( n68266 , n68255 , n68264 );
or ( n68267 , n68260 , n68265 , n68266 );
and ( n68268 , n68215 , n68216 );
and ( n68269 , n68216 , n68221 );
and ( n68270 , n68215 , n68221 );
or ( n68271 , n68268 , n68269 , n68270 );
and ( n68272 , n66786 , n64789 );
and ( n68273 , n66781 , n64787 );
nor ( n68274 , n68272 , n68273 );
xnor ( n68275 , n68274 , n64738 );
and ( n68276 , n68271 , n68275 );
and ( n68277 , n67111 , n64711 );
and ( n68278 , n66981 , n64709 );
nor ( n68279 , n68277 , n68278 );
xnor ( n68280 , n68279 , n64682 );
and ( n68281 , n68275 , n68280 );
and ( n68282 , n68271 , n68280 );
or ( n68283 , n68276 , n68281 , n68282 );
and ( n68284 , n65883 , n65371 );
and ( n68285 , n65698 , n65369 );
nor ( n68286 , n68284 , n68285 );
xnor ( n68287 , n68286 , n65168 );
and ( n68288 , n68283 , n68287 );
and ( n68289 , n66137 , n65183 );
and ( n68290 , n65935 , n65181 );
nor ( n68291 , n68289 , n68290 );
xnor ( n68292 , n68291 , n64994 );
and ( n68293 , n68287 , n68292 );
and ( n68294 , n68283 , n68292 );
or ( n68295 , n68288 , n68293 , n68294 );
xor ( n68296 , n68079 , n68083 );
xor ( n68297 , n68296 , n68088 );
and ( n68298 , n68295 , n68297 );
xor ( n68299 , n67895 , n67899 );
xor ( n68300 , n68299 , n67902 );
and ( n68301 , n68297 , n68300 );
and ( n68302 , n68295 , n68300 );
or ( n68303 , n68298 , n68301 , n68302 );
and ( n68304 , n64781 , n67160 );
and ( n68305 , n64703 , n67158 );
nor ( n68306 , n68304 , n68305 );
xnor ( n68307 , n68306 , n66514 );
and ( n68308 , n68303 , n68307 );
xor ( n68309 , n68091 , n68115 );
xor ( n68310 , n68309 , n68118 );
and ( n68311 , n68307 , n68310 );
and ( n68312 , n68303 , n68310 );
or ( n68313 , n68308 , n68311 , n68312 );
and ( n68314 , n68267 , n68313 );
xor ( n68315 , n68063 , n68067 );
xor ( n68316 , n68315 , n68072 );
and ( n68317 , n68313 , n68316 );
and ( n68318 , n68267 , n68316 );
or ( n68319 , n68314 , n68317 , n68318 );
and ( n68320 , n65935 , n65371 );
and ( n68321 , n65883 , n65369 );
nor ( n68322 , n68320 , n68321 );
xnor ( n68323 , n68322 , n65168 );
and ( n68324 , n66266 , n65056 );
and ( n68325 , n66276 , n65054 );
nor ( n68326 , n68324 , n68325 );
xnor ( n68327 , n68326 , n64943 );
and ( n68328 , n68323 , n68327 );
xor ( n68329 , n68271 , n68275 );
xor ( n68330 , n68329 , n68280 );
and ( n68331 , n68327 , n68330 );
and ( n68332 , n68323 , n68330 );
or ( n68333 , n68328 , n68331 , n68332 );
and ( n68334 , n65453 , n65756 );
and ( n68335 , n65306 , n65754 );
nor ( n68336 , n68334 , n68335 );
xnor ( n68337 , n68336 , n65450 );
and ( n68338 , n68333 , n68337 );
xor ( n68339 , n68095 , n68099 );
xor ( n68340 , n68339 , n68102 );
and ( n68341 , n68337 , n68340 );
and ( n68342 , n68333 , n68340 );
or ( n68343 , n68338 , n68341 , n68342 );
and ( n68344 , n65135 , n66241 );
and ( n68345 , n65001 , n66239 );
nor ( n68346 , n68344 , n68345 );
xnor ( n68347 , n68346 , n65876 );
and ( n68348 , n68343 , n68347 );
and ( n68349 , n65265 , n66016 );
and ( n68350 , n65175 , n66014 );
nor ( n68351 , n68349 , n68350 );
xnor ( n68352 , n68351 , n65650 );
and ( n68353 , n68347 , n68352 );
and ( n68354 , n68343 , n68352 );
or ( n68355 , n68348 , n68353 , n68354 );
and ( n68356 , n64906 , n66906 );
and ( n68357 , n64857 , n66904 );
nor ( n68358 , n68356 , n68357 );
xnor ( n68359 , n68358 , n66286 );
and ( n68360 , n65306 , n65756 );
and ( n68361 , n65363 , n65754 );
nor ( n68362 , n68360 , n68361 );
xnor ( n68363 , n68362 , n65450 );
and ( n68364 , n68359 , n68363 );
xor ( n68365 , n68295 , n68297 );
xor ( n68366 , n68365 , n68300 );
and ( n68367 , n68363 , n68366 );
and ( n68368 , n68359 , n68366 );
or ( n68369 , n68364 , n68367 , n68368 );
and ( n68370 , n68355 , n68369 );
xor ( n68371 , n68141 , n68145 );
xor ( n68372 , n68371 , n68150 );
and ( n68373 , n68369 , n68372 );
and ( n68374 , n68355 , n68372 );
or ( n68375 , n68370 , n68373 , n68374 );
xor ( n68376 , n68121 , n68125 );
xor ( n68377 , n68376 , n68128 );
and ( n68378 , n68375 , n68377 );
xor ( n68379 , n68153 , n68155 );
xor ( n68380 , n68379 , n68158 );
and ( n68381 , n68377 , n68380 );
and ( n68382 , n68375 , n68380 );
or ( n68383 , n68378 , n68381 , n68382 );
and ( n68384 , n68319 , n68383 );
xor ( n68385 , n68075 , n68131 );
xor ( n68386 , n68385 , n68134 );
and ( n68387 , n68383 , n68386 );
and ( n68388 , n68319 , n68386 );
or ( n68389 , n68384 , n68387 , n68388 );
xor ( n68390 , n68023 , n68025 );
xor ( n68391 , n68390 , n68028 );
and ( n68392 , n68389 , n68391 );
xor ( n68393 , n68137 , n68169 );
xor ( n68394 , n68393 , n68172 );
and ( n68395 , n68391 , n68394 );
and ( n68396 , n68389 , n68394 );
or ( n68397 , n68392 , n68395 , n68396 );
and ( n68398 , n68187 , n68397 );
xor ( n68399 , n68187 , n68397 );
xor ( n68400 , n68389 , n68391 );
xor ( n68401 , n68400 , n68394 );
and ( n68402 , n66276 , n65183 );
and ( n68403 , n66142 , n65181 );
nor ( n68404 , n68402 , n68403 );
xnor ( n68405 , n68404 , n64994 );
and ( n68406 , n66517 , n65056 );
and ( n68407 , n66266 , n65054 );
nor ( n68408 , n68406 , n68407 );
xnor ( n68409 , n68408 , n64943 );
and ( n68410 , n68405 , n68409 );
xor ( n68411 , n68209 , n68213 );
xor ( n68412 , n68411 , n68222 );
and ( n68413 , n68409 , n68412 );
and ( n68414 , n68405 , n68412 );
or ( n68415 , n68410 , n68413 , n68414 );
and ( n68416 , n65443 , n65756 );
and ( n68417 , n65453 , n65754 );
nor ( n68418 , n68416 , n68417 );
xnor ( n68419 , n68418 , n65450 );
and ( n68420 , n68415 , n68419 );
xor ( n68421 , n68225 , n68229 );
xor ( n68422 , n68421 , n68232 );
and ( n68423 , n68419 , n68422 );
and ( n68424 , n68415 , n68422 );
or ( n68425 , n68420 , n68423 , n68424 );
and ( n68426 , n65001 , n66657 );
and ( n68427 , n64955 , n66655 );
nor ( n68428 , n68426 , n68427 );
xnor ( n68429 , n68428 , n66130 );
and ( n68430 , n68425 , n68429 );
and ( n68431 , n65175 , n66241 );
and ( n68432 , n65135 , n66239 );
nor ( n68433 , n68431 , n68432 );
xnor ( n68434 , n68433 , n65876 );
and ( n68435 , n68429 , n68434 );
and ( n68436 , n68425 , n68434 );
or ( n68437 , n68430 , n68435 , n68436 );
xor ( n68438 , n68198 , n68200 );
buf ( n68439 , n64549 );
and ( n68440 , n68439 , n64617 );
and ( n68441 , n68199 , n64615 );
nor ( n68442 , n68440 , n68441 );
xnor ( n68443 , n68442 , n64624 );
buf ( n68444 , n64550 );
and ( n68445 , n68444 , n64612 );
and ( n68446 , n68443 , n68445 );
and ( n68447 , n68439 , n64612 );
and ( n68448 , n68446 , n68447 );
and ( n68449 , n68438 , n68448 );
and ( n68450 , n68192 , n64617 );
and ( n68451 , n67873 , n64615 );
nor ( n68452 , n68450 , n68451 );
xnor ( n68453 , n68452 , n64624 );
and ( n68454 , n68448 , n68453 );
and ( n68455 , n68438 , n68453 );
or ( n68456 , n68449 , n68454 , n68455 );
and ( n68457 , n67307 , n64711 );
and ( n68458 , n67302 , n64709 );
nor ( n68459 , n68457 , n68458 );
xnor ( n68460 , n68459 , n64682 );
and ( n68461 , n68456 , n68460 );
xor ( n68462 , n68194 , n68201 );
xor ( n68463 , n68462 , n68206 );
and ( n68464 , n68460 , n68463 );
and ( n68465 , n68456 , n68463 );
or ( n68466 , n68461 , n68464 , n68465 );
and ( n68467 , n66781 , n64897 );
and ( n68468 , n66507 , n64895 );
nor ( n68469 , n68467 , n68468 );
xnor ( n68470 , n68469 , n64850 );
and ( n68471 , n68466 , n68470 );
and ( n68472 , n66981 , n64789 );
and ( n68473 , n66786 , n64787 );
nor ( n68474 , n68472 , n68473 );
xnor ( n68475 , n68474 , n64738 );
and ( n68476 , n68470 , n68475 );
and ( n68477 , n68466 , n68475 );
or ( n68478 , n68471 , n68476 , n68477 );
and ( n68479 , n65698 , n65550 );
and ( n68480 , n65657 , n65548 );
nor ( n68481 , n68479 , n68480 );
xnor ( n68482 , n68481 , n65313 );
and ( n68483 , n68478 , n68482 );
and ( n68484 , n66142 , n65183 );
and ( n68485 , n66137 , n65181 );
nor ( n68486 , n68484 , n68485 );
xnor ( n68487 , n68486 , n64994 );
and ( n68488 , n68482 , n68487 );
and ( n68489 , n68478 , n68487 );
or ( n68490 , n68483 , n68488 , n68489 );
xor ( n68491 , n68283 , n68287 );
xor ( n68492 , n68491 , n68292 );
and ( n68493 , n68490 , n68492 );
xor ( n68494 , n68235 , n68239 );
xor ( n68495 , n68494 , n68242 );
and ( n68496 , n68492 , n68495 );
and ( n68497 , n68490 , n68495 );
or ( n68498 , n68493 , n68496 , n68497 );
and ( n68499 , n68437 , n68498 );
and ( n68500 , n64798 , n67160 );
and ( n68501 , n64781 , n67158 );
nor ( n68502 , n68500 , n68501 );
xnor ( n68503 , n68502 , n66514 );
and ( n68504 , n68498 , n68503 );
and ( n68505 , n68437 , n68503 );
or ( n68506 , n68499 , n68504 , n68505 );
xor ( n68507 , n68055 , n68057 );
xor ( n68508 , n68507 , n68060 );
and ( n68509 , n68506 , n68508 );
xor ( n68510 , n68303 , n68307 );
xor ( n68511 , n68510 , n68310 );
and ( n68512 , n68508 , n68511 );
and ( n68513 , n68506 , n68511 );
or ( n68514 , n68509 , n68512 , n68513 );
xor ( n68515 , n68267 , n68313 );
xor ( n68516 , n68515 , n68316 );
and ( n68517 , n68514 , n68516 );
xor ( n68518 , n68375 , n68377 );
xor ( n68519 , n68518 , n68380 );
and ( n68520 , n68516 , n68519 );
and ( n68521 , n68514 , n68519 );
or ( n68522 , n68517 , n68520 , n68521 );
xor ( n68523 , n68319 , n68383 );
xor ( n68524 , n68523 , n68386 );
and ( n68525 , n68522 , n68524 );
xor ( n68526 , n68161 , n68163 );
xor ( n68527 , n68526 , n68166 );
and ( n68528 , n68524 , n68527 );
and ( n68529 , n68522 , n68527 );
or ( n68530 , n68525 , n68528 , n68529 );
and ( n68531 , n68401 , n68530 );
xor ( n68532 , n68401 , n68530 );
xor ( n68533 , n68522 , n68524 );
xor ( n68534 , n68533 , n68527 );
xor ( n68535 , n68446 , n68447 );
and ( n68536 , n67873 , n64652 );
and ( n68537 , n67833 , n64650 );
nor ( n68538 , n68536 , n68537 );
xnor ( n68539 , n68538 , n64609 );
and ( n68540 , n68535 , n68539 );
and ( n68541 , n68199 , n64617 );
and ( n68542 , n68192 , n64615 );
nor ( n68543 , n68541 , n68542 );
xnor ( n68544 , n68543 , n64624 );
and ( n68545 , n68539 , n68544 );
and ( n68546 , n68535 , n68544 );
or ( n68547 , n68540 , n68545 , n68546 );
and ( n68548 , n67302 , n64789 );
and ( n68549 , n67111 , n64787 );
nor ( n68550 , n68548 , n68549 );
xnor ( n68551 , n68550 , n64738 );
and ( n68552 , n68547 , n68551 );
and ( n68553 , n67548 , n64711 );
and ( n68554 , n67307 , n64709 );
nor ( n68555 , n68553 , n68554 );
xnor ( n68556 , n68555 , n64682 );
and ( n68557 , n68551 , n68556 );
and ( n68558 , n68547 , n68556 );
or ( n68559 , n68552 , n68557 , n68558 );
and ( n68560 , n66786 , n64897 );
and ( n68561 , n66781 , n64895 );
nor ( n68562 , n68560 , n68561 );
xnor ( n68563 , n68562 , n64850 );
and ( n68564 , n68559 , n68563 );
and ( n68565 , n67111 , n64789 );
and ( n68566 , n66981 , n64787 );
nor ( n68567 , n68565 , n68566 );
xnor ( n68568 , n68567 , n64738 );
and ( n68569 , n68563 , n68568 );
and ( n68570 , n68559 , n68568 );
or ( n68571 , n68564 , n68569 , n68570 );
and ( n68572 , n65883 , n65550 );
and ( n68573 , n65698 , n65548 );
nor ( n68574 , n68572 , n68573 );
xnor ( n68575 , n68574 , n65313 );
and ( n68576 , n68571 , n68575 );
and ( n68577 , n66137 , n65371 );
and ( n68578 , n65935 , n65369 );
nor ( n68579 , n68577 , n68578 );
xnor ( n68580 , n68579 , n65168 );
and ( n68581 , n68575 , n68580 );
and ( n68582 , n68571 , n68580 );
or ( n68583 , n68576 , n68581 , n68582 );
xor ( n68584 , n68478 , n68482 );
xor ( n68585 , n68584 , n68487 );
and ( n68586 , n68583 , n68585 );
xor ( n68587 , n68323 , n68327 );
xor ( n68588 , n68587 , n68330 );
and ( n68589 , n68585 , n68588 );
and ( n68590 , n68583 , n68588 );
or ( n68591 , n68586 , n68589 , n68590 );
and ( n68592 , n65363 , n66016 );
and ( n68593 , n65265 , n66014 );
nor ( n68594 , n68592 , n68593 );
xnor ( n68595 , n68594 , n65650 );
and ( n68596 , n68591 , n68595 );
xor ( n68597 , n68333 , n68337 );
xor ( n68598 , n68597 , n68340 );
and ( n68599 , n68595 , n68598 );
and ( n68600 , n68591 , n68598 );
or ( n68601 , n68596 , n68599 , n68600 );
and ( n68602 , n64703 , n67498 );
and ( n68603 , n64689 , n67495 );
nor ( n68604 , n68602 , n68603 );
xnor ( n68605 , n68604 , n66511 );
and ( n68606 , n68601 , n68605 );
xor ( n68607 , n68245 , n68249 );
xor ( n68608 , n68607 , n68252 );
and ( n68609 , n68605 , n68608 );
and ( n68610 , n68601 , n68608 );
or ( n68611 , n68606 , n68609 , n68610 );
xor ( n68612 , n68255 , n68259 );
xor ( n68613 , n68612 , n68264 );
and ( n68614 , n68611 , n68613 );
xor ( n68615 , n68355 , n68369 );
xor ( n68616 , n68615 , n68372 );
and ( n68617 , n68613 , n68616 );
and ( n68618 , n68611 , n68616 );
or ( n68619 , n68614 , n68617 , n68618 );
xor ( n68620 , n68443 , n68445 );
and ( n68621 , n68444 , n64617 );
and ( n68622 , n68439 , n64615 );
nor ( n68623 , n68621 , n68622 );
xnor ( n68624 , n68623 , n64624 );
buf ( n68625 , n64551 );
and ( n68626 , n68625 , n64612 );
and ( n68627 , n68624 , n68626 );
and ( n68628 , n68620 , n68627 );
and ( n68629 , n67833 , n64711 );
and ( n68630 , n67727 , n64709 );
nor ( n68631 , n68629 , n68630 );
xnor ( n68632 , n68631 , n64682 );
and ( n68633 , n68627 , n68632 );
and ( n68634 , n68620 , n68632 );
or ( n68635 , n68628 , n68633 , n68634 );
and ( n68636 , n67307 , n64789 );
and ( n68637 , n67302 , n64787 );
nor ( n68638 , n68636 , n68637 );
xnor ( n68639 , n68638 , n64738 );
and ( n68640 , n68635 , n68639 );
and ( n68641 , n67727 , n64711 );
and ( n68642 , n67548 , n64709 );
nor ( n68643 , n68641 , n68642 );
xnor ( n68644 , n68643 , n64682 );
and ( n68645 , n68639 , n68644 );
and ( n68646 , n68635 , n68644 );
or ( n68647 , n68640 , n68645 , n68646 );
and ( n68648 , n66981 , n64897 );
and ( n68649 , n66786 , n64895 );
nor ( n68650 , n68648 , n68649 );
xnor ( n68651 , n68650 , n64850 );
and ( n68652 , n68647 , n68651 );
xor ( n68653 , n68438 , n68448 );
xor ( n68654 , n68653 , n68453 );
and ( n68655 , n68651 , n68654 );
and ( n68656 , n68647 , n68654 );
or ( n68657 , n68652 , n68655 , n68656 );
and ( n68658 , n65935 , n65550 );
and ( n68659 , n65883 , n65548 );
nor ( n68660 , n68658 , n68659 );
xnor ( n68661 , n68660 , n65313 );
and ( n68662 , n68657 , n68661 );
xor ( n68663 , n68559 , n68563 );
xor ( n68664 , n68663 , n68568 );
and ( n68665 , n68661 , n68664 );
and ( n68666 , n68657 , n68664 );
or ( n68667 , n68662 , n68665 , n68666 );
and ( n68668 , n65657 , n65756 );
and ( n68669 , n65443 , n65754 );
nor ( n68670 , n68668 , n68669 );
xnor ( n68671 , n68670 , n65450 );
and ( n68672 , n68667 , n68671 );
xor ( n68673 , n68405 , n68409 );
xor ( n68674 , n68673 , n68412 );
and ( n68675 , n68671 , n68674 );
and ( n68676 , n68667 , n68674 );
or ( n68677 , n68672 , n68675 , n68676 );
and ( n68678 , n64955 , n66906 );
and ( n68679 , n64950 , n66904 );
nor ( n68680 , n68678 , n68679 );
xnor ( n68681 , n68680 , n66286 );
and ( n68682 , n68677 , n68681 );
and ( n68683 , n65265 , n66241 );
and ( n68684 , n65175 , n66239 );
nor ( n68685 , n68683 , n68684 );
xnor ( n68686 , n68685 , n65876 );
and ( n68687 , n68681 , n68686 );
and ( n68688 , n68677 , n68686 );
or ( n68689 , n68682 , n68687 , n68688 );
and ( n68690 , n64781 , n67498 );
and ( n68691 , n64703 , n67495 );
nor ( n68692 , n68690 , n68691 );
xnor ( n68693 , n68692 , n66511 );
and ( n68694 , n68689 , n68693 );
and ( n68695 , n64857 , n67160 );
and ( n68696 , n64798 , n67158 );
nor ( n68697 , n68695 , n68696 );
xnor ( n68698 , n68697 , n66514 );
and ( n68699 , n68693 , n68698 );
and ( n68700 , n68689 , n68698 );
or ( n68701 , n68694 , n68699 , n68700 );
xor ( n68702 , n68343 , n68347 );
xor ( n68703 , n68702 , n68352 );
and ( n68704 , n68701 , n68703 );
xor ( n68705 , n68359 , n68363 );
xor ( n68706 , n68705 , n68366 );
and ( n68707 , n68703 , n68706 );
and ( n68708 , n68701 , n68706 );
or ( n68709 , n68704 , n68707 , n68708 );
and ( n68710 , n66266 , n65183 );
and ( n68711 , n66276 , n65181 );
nor ( n68712 , n68710 , n68711 );
xnor ( n68713 , n68712 , n64994 );
and ( n68714 , n66507 , n65056 );
and ( n68715 , n66517 , n65054 );
nor ( n68716 , n68714 , n68715 );
xnor ( n68717 , n68716 , n64943 );
and ( n68718 , n68713 , n68717 );
xor ( n68719 , n68456 , n68460 );
xor ( n68720 , n68719 , n68463 );
and ( n68721 , n68717 , n68720 );
and ( n68722 , n68713 , n68720 );
or ( n68723 , n68718 , n68721 , n68722 );
and ( n68724 , n65453 , n66016 );
and ( n68725 , n65306 , n66014 );
nor ( n68726 , n68724 , n68725 );
xnor ( n68727 , n68726 , n65650 );
and ( n68728 , n68723 , n68727 );
xor ( n68729 , n68466 , n68470 );
xor ( n68730 , n68729 , n68475 );
and ( n68731 , n68727 , n68730 );
and ( n68732 , n68723 , n68730 );
or ( n68733 , n68728 , n68731 , n68732 );
and ( n68734 , n65135 , n66657 );
and ( n68735 , n65001 , n66655 );
nor ( n68736 , n68734 , n68735 );
xnor ( n68737 , n68736 , n66130 );
and ( n68738 , n68733 , n68737 );
xor ( n68739 , n68415 , n68419 );
xor ( n68740 , n68739 , n68422 );
and ( n68741 , n68737 , n68740 );
and ( n68742 , n68733 , n68740 );
or ( n68743 , n68738 , n68741 , n68742 );
and ( n68744 , n64950 , n66906 );
and ( n68745 , n64906 , n66904 );
nor ( n68746 , n68744 , n68745 );
xnor ( n68747 , n68746 , n66286 );
and ( n68748 , n68743 , n68747 );
xor ( n68749 , n68490 , n68492 );
xor ( n68750 , n68749 , n68495 );
and ( n68751 , n68747 , n68750 );
and ( n68752 , n68743 , n68750 );
or ( n68753 , n68748 , n68751 , n68752 );
and ( n68754 , n64906 , n67160 );
and ( n68755 , n64857 , n67158 );
nor ( n68756 , n68754 , n68755 );
xnor ( n68757 , n68756 , n66514 );
and ( n68758 , n65306 , n66016 );
and ( n68759 , n65363 , n66014 );
nor ( n68760 , n68758 , n68759 );
xnor ( n68761 , n68760 , n65650 );
and ( n68762 , n68757 , n68761 );
xor ( n68763 , n68583 , n68585 );
xor ( n68764 , n68763 , n68588 );
and ( n68765 , n68761 , n68764 );
and ( n68766 , n68757 , n68764 );
or ( n68767 , n68762 , n68765 , n68766 );
xor ( n68768 , n68425 , n68429 );
xor ( n68769 , n68768 , n68434 );
and ( n68770 , n68767 , n68769 );
xor ( n68771 , n68591 , n68595 );
xor ( n68772 , n68771 , n68598 );
and ( n68773 , n68769 , n68772 );
and ( n68774 , n68767 , n68772 );
or ( n68775 , n68770 , n68773 , n68774 );
and ( n68776 , n68753 , n68775 );
xor ( n68777 , n68601 , n68605 );
xor ( n68778 , n68777 , n68608 );
and ( n68779 , n68775 , n68778 );
and ( n68780 , n68753 , n68778 );
or ( n68781 , n68776 , n68779 , n68780 );
and ( n68782 , n68709 , n68781 );
xor ( n68783 , n68506 , n68508 );
xor ( n68784 , n68783 , n68511 );
and ( n68785 , n68781 , n68784 );
and ( n68786 , n68709 , n68784 );
or ( n68787 , n68782 , n68785 , n68786 );
and ( n68788 , n68619 , n68787 );
xor ( n68789 , n68514 , n68516 );
xor ( n68790 , n68789 , n68519 );
and ( n68791 , n68787 , n68790 );
and ( n68792 , n68619 , n68790 );
or ( n68793 , n68788 , n68791 , n68792 );
and ( n68794 , n68534 , n68793 );
xor ( n68795 , n68534 , n68793 );
xor ( n68796 , n68619 , n68787 );
xor ( n68797 , n68796 , n68790 );
and ( n68798 , n66276 , n65371 );
and ( n68799 , n66142 , n65369 );
nor ( n68800 , n68798 , n68799 );
xnor ( n68801 , n68800 , n65168 );
and ( n68802 , n66781 , n65056 );
and ( n68803 , n66507 , n65054 );
nor ( n68804 , n68802 , n68803 );
xnor ( n68805 , n68804 , n64943 );
and ( n68806 , n68801 , n68805 );
xor ( n68807 , n68547 , n68551 );
xor ( n68808 , n68807 , n68556 );
and ( n68809 , n68805 , n68808 );
and ( n68810 , n68801 , n68808 );
or ( n68811 , n68806 , n68809 , n68810 );
and ( n68812 , n65698 , n65756 );
and ( n68813 , n65657 , n65754 );
nor ( n68814 , n68812 , n68813 );
xnor ( n68815 , n68814 , n65450 );
and ( n68816 , n68811 , n68815 );
and ( n68817 , n66142 , n65371 );
and ( n68818 , n66137 , n65369 );
nor ( n68819 , n68817 , n68818 );
xnor ( n68820 , n68819 , n65168 );
and ( n68821 , n68815 , n68820 );
and ( n68822 , n68811 , n68820 );
or ( n68823 , n68816 , n68821 , n68822 );
xor ( n68824 , n68571 , n68575 );
xor ( n68825 , n68824 , n68580 );
and ( n68826 , n68823 , n68825 );
xor ( n68827 , n68723 , n68727 );
xor ( n68828 , n68827 , n68730 );
and ( n68829 , n68825 , n68828 );
and ( n68830 , n68823 , n68828 );
or ( n68831 , n68826 , n68829 , n68830 );
xor ( n68832 , n68624 , n68626 );
and ( n68833 , n68625 , n64617 );
and ( n68834 , n68444 , n64615 );
nor ( n68835 , n68833 , n68834 );
xnor ( n68836 , n68835 , n64624 );
buf ( n68837 , n64552 );
and ( n68838 , n68837 , n64612 );
and ( n68839 , n68836 , n68838 );
and ( n68840 , n68832 , n68839 );
and ( n68841 , n67873 , n64711 );
and ( n68842 , n67833 , n64709 );
nor ( n68843 , n68841 , n68842 );
xnor ( n68844 , n68843 , n64682 );
and ( n68845 , n68839 , n68844 );
and ( n68846 , n68832 , n68844 );
or ( n68847 , n68840 , n68845 , n68846 );
and ( n68848 , n68192 , n64652 );
and ( n68849 , n67873 , n64650 );
nor ( n68850 , n68848 , n68849 );
xnor ( n68851 , n68850 , n64609 );
and ( n68852 , n68847 , n68851 );
xor ( n68853 , n68620 , n68627 );
xor ( n68854 , n68853 , n68632 );
and ( n68855 , n68851 , n68854 );
and ( n68856 , n68847 , n68854 );
or ( n68857 , n68852 , n68855 , n68856 );
and ( n68858 , n67111 , n64897 );
and ( n68859 , n66981 , n64895 );
nor ( n68860 , n68858 , n68859 );
xnor ( n68861 , n68860 , n64850 );
and ( n68862 , n68857 , n68861 );
xor ( n68863 , n68535 , n68539 );
xor ( n68864 , n68863 , n68544 );
and ( n68865 , n68861 , n68864 );
and ( n68866 , n68857 , n68864 );
or ( n68867 , n68862 , n68865 , n68866 );
xor ( n68868 , n68836 , n68838 );
and ( n68869 , n68444 , n64652 );
and ( n68870 , n68439 , n64650 );
nor ( n68871 , n68869 , n68870 );
xnor ( n68872 , n68871 , n64609 );
buf ( n68873 , n64553 );
and ( n68874 , n68873 , n64612 );
and ( n68875 , n68872 , n68874 );
and ( n68876 , n68868 , n68875 );
and ( n68877 , n68439 , n64652 );
and ( n68878 , n68199 , n64650 );
nor ( n68879 , n68877 , n68878 );
xnor ( n68880 , n68879 , n64609 );
and ( n68881 , n68875 , n68880 );
and ( n68882 , n68868 , n68880 );
or ( n68883 , n68876 , n68881 , n68882 );
and ( n68884 , n67727 , n64789 );
and ( n68885 , n67548 , n64787 );
nor ( n68886 , n68884 , n68885 );
xnor ( n68887 , n68886 , n64738 );
and ( n68888 , n68883 , n68887 );
and ( n68889 , n68199 , n64652 );
and ( n68890 , n68192 , n64650 );
nor ( n68891 , n68889 , n68890 );
xnor ( n68892 , n68891 , n64609 );
and ( n68893 , n68887 , n68892 );
and ( n68894 , n68883 , n68892 );
or ( n68895 , n68888 , n68893 , n68894 );
and ( n68896 , n67302 , n64897 );
and ( n68897 , n67111 , n64895 );
nor ( n68898 , n68896 , n68897 );
xnor ( n68899 , n68898 , n64850 );
and ( n68900 , n68895 , n68899 );
and ( n68901 , n67548 , n64789 );
and ( n68902 , n67307 , n64787 );
nor ( n68903 , n68901 , n68902 );
xnor ( n68904 , n68903 , n64738 );
and ( n68905 , n68899 , n68904 );
and ( n68906 , n68895 , n68904 );
or ( n68907 , n68900 , n68905 , n68906 );
and ( n68908 , n66786 , n65056 );
and ( n68909 , n66781 , n65054 );
nor ( n68910 , n68908 , n68909 );
xnor ( n68911 , n68910 , n64943 );
and ( n68912 , n68907 , n68911 );
xor ( n68913 , n68635 , n68639 );
xor ( n68914 , n68913 , n68644 );
and ( n68915 , n68911 , n68914 );
and ( n68916 , n68907 , n68914 );
or ( n68917 , n68912 , n68915 , n68916 );
and ( n68918 , n68867 , n68917 );
and ( n68919 , n66517 , n65183 );
and ( n68920 , n66266 , n65181 );
nor ( n68921 , n68919 , n68920 );
xnor ( n68922 , n68921 , n64994 );
and ( n68923 , n68917 , n68922 );
and ( n68924 , n68867 , n68922 );
or ( n68925 , n68918 , n68923 , n68924 );
and ( n68926 , n65443 , n66016 );
and ( n68927 , n65453 , n66014 );
nor ( n68928 , n68926 , n68927 );
xnor ( n68929 , n68928 , n65650 );
and ( n68930 , n68925 , n68929 );
xor ( n68931 , n68713 , n68717 );
xor ( n68932 , n68931 , n68720 );
and ( n68933 , n68929 , n68932 );
and ( n68934 , n68925 , n68932 );
or ( n68935 , n68930 , n68933 , n68934 );
and ( n68936 , n65175 , n66657 );
and ( n68937 , n65135 , n66655 );
nor ( n68938 , n68936 , n68937 );
xnor ( n68939 , n68938 , n66130 );
and ( n68940 , n68935 , n68939 );
xor ( n68941 , n68667 , n68671 );
xor ( n68942 , n68941 , n68674 );
and ( n68943 , n68939 , n68942 );
and ( n68944 , n68935 , n68942 );
or ( n68945 , n68940 , n68943 , n68944 );
and ( n68946 , n68831 , n68945 );
and ( n68947 , n64798 , n67498 );
and ( n68948 , n64781 , n67495 );
nor ( n68949 , n68947 , n68948 );
xnor ( n68950 , n68949 , n66511 );
and ( n68951 , n68945 , n68950 );
and ( n68952 , n68831 , n68950 );
or ( n68953 , n68946 , n68951 , n68952 );
xor ( n68954 , n68689 , n68693 );
xor ( n68955 , n68954 , n68698 );
and ( n68956 , n68953 , n68955 );
xor ( n68957 , n68743 , n68747 );
xor ( n68958 , n68957 , n68750 );
and ( n68959 , n68955 , n68958 );
and ( n68960 , n68953 , n68958 );
or ( n68961 , n68956 , n68959 , n68960 );
xor ( n68962 , n68437 , n68498 );
xor ( n68963 , n68962 , n68503 );
and ( n68964 , n68961 , n68963 );
xor ( n68965 , n68701 , n68703 );
xor ( n68966 , n68965 , n68706 );
and ( n68967 , n68963 , n68966 );
and ( n68968 , n68961 , n68966 );
or ( n68969 , n68964 , n68967 , n68968 );
xor ( n68970 , n68611 , n68613 );
xor ( n68971 , n68970 , n68616 );
and ( n68972 , n68969 , n68971 );
xor ( n68973 , n68709 , n68781 );
xor ( n68974 , n68973 , n68784 );
and ( n68975 , n68971 , n68974 );
and ( n68976 , n68969 , n68974 );
or ( n68977 , n68972 , n68975 , n68976 );
and ( n68978 , n68797 , n68977 );
xor ( n68979 , n68797 , n68977 );
xor ( n68980 , n68969 , n68971 );
xor ( n68981 , n68980 , n68974 );
and ( n68982 , n64950 , n67160 );
and ( n68983 , n64906 , n67158 );
nor ( n68984 , n68982 , n68983 );
xnor ( n68985 , n68984 , n66514 );
and ( n68986 , n65001 , n66906 );
and ( n68987 , n64955 , n66904 );
nor ( n68988 , n68986 , n68987 );
xnor ( n68989 , n68988 , n66286 );
and ( n68990 , n68985 , n68989 );
and ( n68991 , n65363 , n66241 );
and ( n68992 , n65265 , n66239 );
nor ( n68993 , n68991 , n68992 );
xnor ( n68994 , n68993 , n65876 );
and ( n68995 , n68989 , n68994 );
and ( n68996 , n68985 , n68994 );
or ( n68997 , n68990 , n68995 , n68996 );
xor ( n68998 , n68677 , n68681 );
xor ( n68999 , n68998 , n68686 );
and ( n69000 , n68997 , n68999 );
xor ( n69001 , n68733 , n68737 );
xor ( n69002 , n69001 , n68740 );
and ( n69003 , n68999 , n69002 );
and ( n69004 , n68997 , n69002 );
or ( n69005 , n69000 , n69003 , n69004 );
xor ( n69006 , n68767 , n68769 );
xor ( n69007 , n69006 , n68772 );
and ( n69008 , n69005 , n69007 );
xor ( n69009 , n68953 , n68955 );
xor ( n69010 , n69009 , n68958 );
and ( n69011 , n69007 , n69010 );
and ( n69012 , n69005 , n69010 );
or ( n69013 , n69008 , n69011 , n69012 );
xor ( n69014 , n68753 , n68775 );
xor ( n69015 , n69014 , n68778 );
and ( n69016 , n69013 , n69015 );
xor ( n69017 , n68961 , n68963 );
xor ( n69018 , n69017 , n68966 );
and ( n69019 , n69015 , n69018 );
and ( n69020 , n69013 , n69018 );
or ( n69021 , n69016 , n69019 , n69020 );
and ( n69022 , n68981 , n69021 );
xor ( n69023 , n68981 , n69021 );
xor ( n69024 , n69013 , n69015 );
xor ( n69025 , n69024 , n69018 );
and ( n69026 , n66266 , n65371 );
and ( n69027 , n66276 , n65369 );
nor ( n69028 , n69026 , n69027 );
xnor ( n69029 , n69028 , n65168 );
and ( n69030 , n66507 , n65183 );
and ( n69031 , n66517 , n65181 );
nor ( n69032 , n69030 , n69031 );
xnor ( n69033 , n69032 , n64994 );
and ( n69034 , n69029 , n69033 );
xor ( n69035 , n68857 , n68861 );
xor ( n69036 , n69035 , n68864 );
and ( n69037 , n69033 , n69036 );
and ( n69038 , n69029 , n69036 );
or ( n69039 , n69034 , n69037 , n69038 );
and ( n69040 , n65657 , n66016 );
and ( n69041 , n65443 , n66014 );
nor ( n69042 , n69040 , n69041 );
xnor ( n69043 , n69042 , n65650 );
and ( n69044 , n69039 , n69043 );
xor ( n69045 , n68801 , n68805 );
xor ( n69046 , n69045 , n68808 );
and ( n69047 , n69043 , n69046 );
and ( n69048 , n69039 , n69046 );
or ( n69049 , n69044 , n69047 , n69048 );
and ( n69050 , n65135 , n66906 );
and ( n69051 , n65001 , n66904 );
nor ( n69052 , n69050 , n69051 );
xnor ( n69053 , n69052 , n66286 );
and ( n69054 , n69049 , n69053 );
and ( n69055 , n65265 , n66657 );
and ( n69056 , n65175 , n66655 );
nor ( n69057 , n69055 , n69056 );
xnor ( n69058 , n69057 , n66130 );
and ( n69059 , n69053 , n69058 );
and ( n69060 , n69049 , n69058 );
or ( n69061 , n69054 , n69059 , n69060 );
and ( n69062 , n65883 , n65756 );
and ( n69063 , n65698 , n65754 );
nor ( n69064 , n69062 , n69063 );
xnor ( n69065 , n69064 , n65450 );
and ( n69066 , n66137 , n65550 );
and ( n69067 , n65935 , n65548 );
nor ( n69068 , n69066 , n69067 );
xnor ( n69069 , n69068 , n65313 );
and ( n69070 , n69065 , n69069 );
xor ( n69071 , n68647 , n68651 );
xor ( n69072 , n69071 , n68654 );
and ( n69073 , n69069 , n69072 );
and ( n69074 , n69065 , n69072 );
or ( n69075 , n69070 , n69073 , n69074 );
xor ( n69076 , n68811 , n68815 );
xor ( n69077 , n69076 , n68820 );
and ( n69078 , n69075 , n69077 );
xor ( n69079 , n68657 , n68661 );
xor ( n69080 , n69079 , n68664 );
and ( n69081 , n69077 , n69080 );
and ( n69082 , n69075 , n69080 );
or ( n69083 , n69078 , n69081 , n69082 );
and ( n69084 , n69061 , n69083 );
xor ( n69085 , n68823 , n68825 );
xor ( n69086 , n69085 , n68828 );
and ( n69087 , n69083 , n69086 );
and ( n69088 , n69061 , n69086 );
or ( n69089 , n69084 , n69087 , n69088 );
xor ( n69090 , n68872 , n68874 );
and ( n69091 , n68873 , n64617 );
and ( n69092 , n68837 , n64615 );
nor ( n69093 , n69091 , n69092 );
xnor ( n69094 , n69093 , n64624 );
buf ( n69095 , n64554 );
and ( n69096 , n69095 , n64612 );
and ( n69097 , n69094 , n69096 );
and ( n69098 , n69090 , n69097 );
and ( n69099 , n68837 , n64617 );
and ( n69100 , n68625 , n64615 );
nor ( n69101 , n69099 , n69100 );
xnor ( n69102 , n69101 , n64624 );
and ( n69103 , n69097 , n69102 );
and ( n69104 , n69090 , n69102 );
or ( n69105 , n69098 , n69103 , n69104 );
and ( n69106 , n67833 , n64789 );
and ( n69107 , n67727 , n64787 );
nor ( n69108 , n69106 , n69107 );
xnor ( n69109 , n69108 , n64738 );
and ( n69110 , n69105 , n69109 );
and ( n69111 , n68192 , n64711 );
and ( n69112 , n67873 , n64709 );
nor ( n69113 , n69111 , n69112 );
xnor ( n69114 , n69113 , n64682 );
and ( n69115 , n69109 , n69114 );
and ( n69116 , n69105 , n69114 );
or ( n69117 , n69110 , n69115 , n69116 );
and ( n69118 , n67307 , n64897 );
and ( n69119 , n67302 , n64895 );
nor ( n69120 , n69118 , n69119 );
xnor ( n69121 , n69120 , n64850 );
and ( n69122 , n69117 , n69121 );
xor ( n69123 , n68832 , n68839 );
xor ( n69124 , n69123 , n68844 );
and ( n69125 , n69121 , n69124 );
and ( n69126 , n69117 , n69124 );
or ( n69127 , n69122 , n69125 , n69126 );
and ( n69128 , n66981 , n65056 );
and ( n69129 , n66786 , n65054 );
nor ( n69130 , n69128 , n69129 );
xnor ( n69131 , n69130 , n64943 );
and ( n69132 , n69127 , n69131 );
xor ( n69133 , n68847 , n68851 );
xor ( n69134 , n69133 , n68854 );
and ( n69135 , n69131 , n69134 );
and ( n69136 , n69127 , n69134 );
or ( n69137 , n69132 , n69135 , n69136 );
and ( n69138 , n65935 , n65756 );
and ( n69139 , n65883 , n65754 );
nor ( n69140 , n69138 , n69139 );
xnor ( n69141 , n69140 , n65450 );
and ( n69142 , n69137 , n69141 );
and ( n69143 , n66142 , n65550 );
and ( n69144 , n66137 , n65548 );
nor ( n69145 , n69143 , n69144 );
xnor ( n69146 , n69145 , n65313 );
and ( n69147 , n69141 , n69146 );
and ( n69148 , n69137 , n69146 );
or ( n69149 , n69142 , n69147 , n69148 );
and ( n69150 , n65453 , n66241 );
and ( n69151 , n65306 , n66239 );
nor ( n69152 , n69150 , n69151 );
xnor ( n69153 , n69152 , n65876 );
and ( n69154 , n69149 , n69153 );
xor ( n69155 , n68867 , n68917 );
xor ( n69156 , n69155 , n68922 );
and ( n69157 , n69153 , n69156 );
and ( n69158 , n69149 , n69156 );
or ( n69159 , n69154 , n69157 , n69158 );
and ( n69160 , n65306 , n66241 );
and ( n69161 , n65363 , n66239 );
nor ( n69162 , n69160 , n69161 );
xnor ( n69163 , n69162 , n65876 );
and ( n69164 , n69159 , n69163 );
xor ( n69165 , n68925 , n68929 );
xor ( n69166 , n69165 , n68932 );
and ( n69167 , n69163 , n69166 );
and ( n69168 , n69159 , n69166 );
or ( n69169 , n69164 , n69167 , n69168 );
and ( n69170 , n64857 , n67498 );
and ( n69171 , n64798 , n67495 );
nor ( n69172 , n69170 , n69171 );
xnor ( n69173 , n69172 , n66511 );
and ( n69174 , n69169 , n69173 );
xor ( n69175 , n68935 , n68939 );
xor ( n69176 , n69175 , n68942 );
and ( n69177 , n69173 , n69176 );
and ( n69178 , n69169 , n69176 );
or ( n69179 , n69174 , n69177 , n69178 );
and ( n69180 , n69089 , n69179 );
xor ( n69181 , n68757 , n68761 );
xor ( n69182 , n69181 , n68764 );
and ( n69183 , n69179 , n69182 );
and ( n69184 , n69089 , n69182 );
or ( n69185 , n69180 , n69183 , n69184 );
and ( n69186 , n64906 , n67498 );
and ( n69187 , n64857 , n67495 );
nor ( n69188 , n69186 , n69187 );
xnor ( n69189 , n69188 , n66511 );
and ( n69190 , n64955 , n67160 );
and ( n69191 , n64950 , n67158 );
nor ( n69192 , n69190 , n69191 );
xnor ( n69193 , n69192 , n66514 );
and ( n69194 , n69189 , n69193 );
xor ( n69195 , n69075 , n69077 );
xor ( n69196 , n69195 , n69080 );
and ( n69197 , n69193 , n69196 );
and ( n69198 , n69189 , n69196 );
or ( n69199 , n69194 , n69197 , n69198 );
xor ( n69200 , n68985 , n68989 );
xor ( n69201 , n69200 , n68994 );
and ( n69202 , n69199 , n69201 );
xor ( n69203 , n69061 , n69083 );
xor ( n69204 , n69203 , n69086 );
and ( n69205 , n69201 , n69204 );
and ( n69206 , n69199 , n69204 );
or ( n69207 , n69202 , n69205 , n69206 );
xor ( n69208 , n68831 , n68945 );
xor ( n69209 , n69208 , n68950 );
and ( n69210 , n69207 , n69209 );
xor ( n69211 , n68997 , n68999 );
xor ( n69212 , n69211 , n69002 );
and ( n69213 , n69209 , n69212 );
and ( n69214 , n69207 , n69212 );
or ( n69215 , n69210 , n69213 , n69214 );
and ( n69216 , n69185 , n69215 );
xor ( n69217 , n69005 , n69007 );
xor ( n69218 , n69217 , n69010 );
and ( n69219 , n69215 , n69218 );
and ( n69220 , n69185 , n69218 );
or ( n69221 , n69216 , n69219 , n69220 );
and ( n69222 , n69025 , n69221 );
xor ( n69223 , n69025 , n69221 );
and ( n69224 , n64950 , n67498 );
and ( n69225 , n64906 , n67495 );
nor ( n69226 , n69224 , n69225 );
xnor ( n69227 , n69226 , n66511 );
and ( n69228 , n65001 , n67160 );
and ( n69229 , n64955 , n67158 );
nor ( n69230 , n69228 , n69229 );
xnor ( n69231 , n69230 , n66514 );
and ( n69232 , n69227 , n69231 );
and ( n69233 , n65175 , n66906 );
and ( n69234 , n65135 , n66904 );
nor ( n69235 , n69233 , n69234 );
xnor ( n69236 , n69235 , n66286 );
and ( n69237 , n69231 , n69236 );
and ( n69238 , n69227 , n69236 );
or ( n69239 , n69232 , n69237 , n69238 );
and ( n69240 , n68625 , n64652 );
and ( n69241 , n68444 , n64650 );
nor ( n69242 , n69240 , n69241 );
xnor ( n69243 , n69242 , n64609 );
xor ( n69244 , n69094 , n69096 );
and ( n69245 , n69243 , n69244 );
and ( n69246 , n67873 , n64789 );
and ( n69247 , n67833 , n64787 );
nor ( n69248 , n69246 , n69247 );
xnor ( n69249 , n69248 , n64738 );
and ( n69250 , n69245 , n69249 );
and ( n69251 , n68199 , n64711 );
and ( n69252 , n68192 , n64709 );
nor ( n69253 , n69251 , n69252 );
xnor ( n69254 , n69253 , n64682 );
and ( n69255 , n69249 , n69254 );
and ( n69256 , n69245 , n69254 );
or ( n69257 , n69250 , n69255 , n69256 );
and ( n69258 , n67548 , n64897 );
and ( n69259 , n67307 , n64895 );
nor ( n69260 , n69258 , n69259 );
xnor ( n69261 , n69260 , n64850 );
and ( n69262 , n69257 , n69261 );
xor ( n69263 , n68868 , n68875 );
xor ( n69264 , n69263 , n68880 );
and ( n69265 , n69261 , n69264 );
and ( n69266 , n69257 , n69264 );
or ( n69267 , n69262 , n69265 , n69266 );
and ( n69268 , n67111 , n65056 );
and ( n69269 , n66981 , n65054 );
nor ( n69270 , n69268 , n69269 );
xnor ( n69271 , n69270 , n64943 );
and ( n69272 , n69267 , n69271 );
xor ( n69273 , n68883 , n68887 );
xor ( n69274 , n69273 , n68892 );
and ( n69275 , n69271 , n69274 );
and ( n69276 , n69267 , n69274 );
or ( n69277 , n69272 , n69275 , n69276 );
and ( n69278 , n66517 , n65371 );
and ( n69279 , n66266 , n65369 );
nor ( n69280 , n69278 , n69279 );
xnor ( n69281 , n69280 , n65168 );
and ( n69282 , n69277 , n69281 );
xor ( n69283 , n69127 , n69131 );
xor ( n69284 , n69283 , n69134 );
and ( n69285 , n69281 , n69284 );
and ( n69286 , n69277 , n69284 );
or ( n69287 , n69282 , n69285 , n69286 );
and ( n69288 , n65443 , n66241 );
and ( n69289 , n65453 , n66239 );
nor ( n69290 , n69288 , n69289 );
xnor ( n69291 , n69290 , n65876 );
and ( n69292 , n69287 , n69291 );
xor ( n69293 , n69029 , n69033 );
xor ( n69294 , n69293 , n69036 );
and ( n69295 , n69291 , n69294 );
and ( n69296 , n69287 , n69294 );
or ( n69297 , n69292 , n69295 , n69296 );
and ( n69298 , n65363 , n66657 );
and ( n69299 , n65265 , n66655 );
nor ( n69300 , n69298 , n69299 );
xnor ( n69301 , n69300 , n66130 );
and ( n69302 , n69297 , n69301 );
xor ( n69303 , n69149 , n69153 );
xor ( n69304 , n69303 , n69156 );
and ( n69305 , n69301 , n69304 );
and ( n69306 , n69297 , n69304 );
or ( n69307 , n69302 , n69305 , n69306 );
and ( n69308 , n69239 , n69307 );
and ( n69309 , n66276 , n65550 );
and ( n69310 , n66142 , n65548 );
nor ( n69311 , n69309 , n69310 );
xnor ( n69312 , n69311 , n65313 );
and ( n69313 , n66781 , n65183 );
and ( n69314 , n66507 , n65181 );
nor ( n69315 , n69313 , n69314 );
xnor ( n69316 , n69315 , n64994 );
and ( n69317 , n69312 , n69316 );
xor ( n69318 , n68895 , n68899 );
xor ( n69319 , n69318 , n68904 );
and ( n69320 , n69316 , n69319 );
and ( n69321 , n69312 , n69319 );
or ( n69322 , n69317 , n69320 , n69321 );
and ( n69323 , n65698 , n66016 );
and ( n69324 , n65657 , n66014 );
nor ( n69325 , n69323 , n69324 );
xnor ( n69326 , n69325 , n65650 );
and ( n69327 , n69322 , n69326 );
xor ( n69328 , n68907 , n68911 );
xor ( n69329 , n69328 , n68914 );
and ( n69330 , n69326 , n69329 );
and ( n69331 , n69322 , n69329 );
or ( n69332 , n69327 , n69330 , n69331 );
xor ( n69333 , n69065 , n69069 );
xor ( n69334 , n69333 , n69072 );
and ( n69335 , n69332 , n69334 );
xor ( n69336 , n69039 , n69043 );
xor ( n69337 , n69336 , n69046 );
and ( n69338 , n69334 , n69337 );
and ( n69339 , n69332 , n69337 );
or ( n69340 , n69335 , n69338 , n69339 );
and ( n69341 , n69307 , n69340 );
and ( n69342 , n69239 , n69340 );
or ( n69343 , n69308 , n69341 , n69342 );
xor ( n69344 , n69049 , n69053 );
xor ( n69345 , n69344 , n69058 );
xor ( n69346 , n69189 , n69193 );
xor ( n69347 , n69346 , n69196 );
and ( n69348 , n69345 , n69347 );
xor ( n69349 , n69159 , n69163 );
xor ( n69350 , n69349 , n69166 );
and ( n69351 , n69347 , n69350 );
and ( n69352 , n69345 , n69350 );
or ( n69353 , n69348 , n69351 , n69352 );
and ( n69354 , n69343 , n69353 );
xor ( n69355 , n69169 , n69173 );
xor ( n69356 , n69355 , n69176 );
and ( n69357 , n69353 , n69356 );
and ( n69358 , n69343 , n69356 );
or ( n69359 , n69354 , n69357 , n69358 );
xor ( n69360 , n69089 , n69179 );
xor ( n69361 , n69360 , n69182 );
and ( n69362 , n69359 , n69361 );
xor ( n69363 , n69207 , n69209 );
xor ( n69364 , n69363 , n69212 );
and ( n69365 , n69361 , n69364 );
and ( n69366 , n69359 , n69364 );
or ( n69367 , n69362 , n69365 , n69366 );
xor ( n69368 , n69185 , n69215 );
xor ( n69369 , n69368 , n69218 );
and ( n69370 , n69367 , n69369 );
xor ( n69371 , n69367 , n69369 );
xor ( n69372 , n69359 , n69361 );
xor ( n69373 , n69372 , n69364 );
and ( n69374 , n65135 , n67160 );
and ( n69375 , n65001 , n67158 );
nor ( n69376 , n69374 , n69375 );
xnor ( n69377 , n69376 , n66514 );
and ( n69378 , n65306 , n66657 );
and ( n69379 , n65363 , n66655 );
nor ( n69380 , n69378 , n69379 );
xnor ( n69381 , n69380 , n66130 );
and ( n69382 , n69377 , n69381 );
xor ( n69383 , n69287 , n69291 );
xor ( n69384 , n69383 , n69294 );
and ( n69385 , n69381 , n69384 );
and ( n69386 , n69377 , n69384 );
or ( n69387 , n69382 , n69385 , n69386 );
xor ( n69388 , n69227 , n69231 );
xor ( n69389 , n69388 , n69236 );
and ( n69390 , n69387 , n69389 );
xor ( n69391 , n69297 , n69301 );
xor ( n69392 , n69391 , n69304 );
and ( n69393 , n69389 , n69392 );
and ( n69394 , n69387 , n69392 );
or ( n69395 , n69390 , n69393 , n69394 );
and ( n69396 , n66507 , n65371 );
and ( n69397 , n66517 , n65369 );
nor ( n69398 , n69396 , n69397 );
xnor ( n69399 , n69398 , n65168 );
and ( n69400 , n66786 , n65183 );
and ( n69401 , n66781 , n65181 );
nor ( n69402 , n69400 , n69401 );
xnor ( n69403 , n69402 , n64994 );
and ( n69404 , n69399 , n69403 );
xor ( n69405 , n69117 , n69121 );
xor ( n69406 , n69405 , n69124 );
and ( n69407 , n69403 , n69406 );
and ( n69408 , n69399 , n69406 );
or ( n69409 , n69404 , n69407 , n69408 );
and ( n69410 , n65883 , n66016 );
and ( n69411 , n65698 , n66014 );
nor ( n69412 , n69410 , n69411 );
xnor ( n69413 , n69412 , n65650 );
and ( n69414 , n69409 , n69413 );
and ( n69415 , n66137 , n65756 );
and ( n69416 , n65935 , n65754 );
nor ( n69417 , n69415 , n69416 );
xnor ( n69418 , n69417 , n65450 );
and ( n69419 , n69413 , n69418 );
and ( n69420 , n69409 , n69418 );
or ( n69421 , n69414 , n69419 , n69420 );
and ( n69422 , n65657 , n66241 );
and ( n69423 , n65443 , n66239 );
nor ( n69424 , n69422 , n69423 );
xnor ( n69425 , n69424 , n65876 );
xor ( n69426 , n69312 , n69316 );
xor ( n69427 , n69426 , n69319 );
and ( n69428 , n69425 , n69427 );
xor ( n69429 , n69277 , n69281 );
xor ( n69430 , n69429 , n69284 );
and ( n69431 , n69427 , n69430 );
and ( n69432 , n69425 , n69430 );
or ( n69433 , n69428 , n69431 , n69432 );
and ( n69434 , n69421 , n69433 );
xor ( n69435 , n69137 , n69141 );
xor ( n69436 , n69435 , n69146 );
and ( n69437 , n69433 , n69436 );
and ( n69438 , n69421 , n69436 );
or ( n69439 , n69434 , n69437 , n69438 );
and ( n69440 , n68444 , n64711 );
and ( n69441 , n68439 , n64709 );
nor ( n69442 , n69440 , n69441 );
xnor ( n69443 , n69442 , n64682 );
and ( n69444 , n69095 , n64617 );
and ( n69445 , n68873 , n64615 );
nor ( n69446 , n69444 , n69445 );
xnor ( n69447 , n69446 , n64624 );
and ( n69448 , n69443 , n69447 );
buf ( n69449 , n64555 );
and ( n69450 , n69449 , n64612 );
and ( n69451 , n69447 , n69450 );
and ( n69452 , n69443 , n69450 );
or ( n69453 , n69448 , n69451 , n69452 );
and ( n69454 , n67833 , n64897 );
and ( n69455 , n67727 , n64895 );
nor ( n69456 , n69454 , n69455 );
xnor ( n69457 , n69456 , n64850 );
and ( n69458 , n69453 , n69457 );
and ( n69459 , n68439 , n64711 );
and ( n69460 , n68199 , n64709 );
nor ( n69461 , n69459 , n69460 );
xnor ( n69462 , n69461 , n64682 );
and ( n69463 , n69457 , n69462 );
and ( n69464 , n69453 , n69462 );
or ( n69465 , n69458 , n69463 , n69464 );
and ( n69466 , n67727 , n64897 );
and ( n69467 , n67548 , n64895 );
nor ( n69468 , n69466 , n69467 );
xnor ( n69469 , n69468 , n64850 );
and ( n69470 , n69465 , n69469 );
xor ( n69471 , n69090 , n69097 );
xor ( n69472 , n69471 , n69102 );
and ( n69473 , n69469 , n69472 );
and ( n69474 , n69465 , n69472 );
or ( n69475 , n69470 , n69473 , n69474 );
and ( n69476 , n67302 , n65056 );
and ( n69477 , n67111 , n65054 );
nor ( n69478 , n69476 , n69477 );
xnor ( n69479 , n69478 , n64943 );
and ( n69480 , n69475 , n69479 );
xor ( n69481 , n69105 , n69109 );
xor ( n69482 , n69481 , n69114 );
and ( n69483 , n69479 , n69482 );
and ( n69484 , n69475 , n69482 );
or ( n69485 , n69480 , n69483 , n69484 );
and ( n69486 , n66781 , n65371 );
and ( n69487 , n66507 , n65369 );
nor ( n69488 , n69486 , n69487 );
xnor ( n69489 , n69488 , n65168 );
and ( n69490 , n66981 , n65183 );
and ( n69491 , n66786 , n65181 );
nor ( n69492 , n69490 , n69491 );
xnor ( n69493 , n69492 , n64994 );
and ( n69494 , n69489 , n69493 );
xor ( n69495 , n69257 , n69261 );
xor ( n69496 , n69495 , n69264 );
and ( n69497 , n69493 , n69496 );
and ( n69498 , n69489 , n69496 );
or ( n69499 , n69494 , n69497 , n69498 );
and ( n69500 , n69485 , n69499 );
and ( n69501 , n66266 , n65550 );
and ( n69502 , n66276 , n65548 );
nor ( n69503 , n69501 , n69502 );
xnor ( n69504 , n69503 , n65313 );
and ( n69505 , n69499 , n69504 );
and ( n69506 , n69485 , n69504 );
or ( n69507 , n69500 , n69505 , n69506 );
and ( n69508 , n65935 , n66016 );
and ( n69509 , n65883 , n66014 );
nor ( n69510 , n69508 , n69509 );
xnor ( n69511 , n69510 , n65650 );
xor ( n69512 , n69267 , n69271 );
xor ( n69513 , n69512 , n69274 );
and ( n69514 , n69511 , n69513 );
xor ( n69515 , n69399 , n69403 );
xor ( n69516 , n69515 , n69406 );
and ( n69517 , n69513 , n69516 );
and ( n69518 , n69511 , n69516 );
or ( n69519 , n69514 , n69517 , n69518 );
and ( n69520 , n69507 , n69519 );
and ( n69521 , n65453 , n66657 );
and ( n69522 , n65306 , n66655 );
nor ( n69523 , n69521 , n69522 );
xnor ( n69524 , n69523 , n66130 );
and ( n69525 , n69519 , n69524 );
and ( n69526 , n69507 , n69524 );
or ( n69527 , n69520 , n69525 , n69526 );
and ( n69528 , n65265 , n66906 );
and ( n69529 , n65175 , n66904 );
nor ( n69530 , n69528 , n69529 );
xnor ( n69531 , n69530 , n66286 );
and ( n69532 , n69527 , n69531 );
xor ( n69533 , n69322 , n69326 );
xor ( n69534 , n69533 , n69329 );
and ( n69535 , n69531 , n69534 );
and ( n69536 , n69527 , n69534 );
or ( n69537 , n69532 , n69535 , n69536 );
and ( n69538 , n69439 , n69537 );
xor ( n69539 , n69332 , n69334 );
xor ( n69540 , n69539 , n69337 );
and ( n69541 , n69537 , n69540 );
and ( n69542 , n69439 , n69540 );
or ( n69543 , n69538 , n69541 , n69542 );
and ( n69544 , n69395 , n69543 );
xor ( n69545 , n69239 , n69307 );
xor ( n69546 , n69545 , n69340 );
and ( n69547 , n69543 , n69546 );
and ( n69548 , n69395 , n69546 );
or ( n69549 , n69544 , n69547 , n69548 );
xor ( n69550 , n69199 , n69201 );
xor ( n69551 , n69550 , n69204 );
and ( n69552 , n69549 , n69551 );
xor ( n69553 , n69343 , n69353 );
xor ( n69554 , n69553 , n69356 );
and ( n69555 , n69551 , n69554 );
and ( n69556 , n69549 , n69554 );
or ( n69557 , n69552 , n69555 , n69556 );
and ( n69558 , n69373 , n69557 );
xor ( n69559 , n69373 , n69557 );
xor ( n69560 , n69549 , n69551 );
xor ( n69561 , n69560 , n69554 );
and ( n69562 , n68873 , n64711 );
and ( n69563 , n68837 , n64709 );
nor ( n69564 , n69562 , n69563 );
xnor ( n69565 , n69564 , n64682 );
buf ( n69566 , n64557 );
and ( n69567 , n69566 , n64617 );
buf ( n69568 , n64556 );
and ( n69569 , n69568 , n64615 );
nor ( n69570 , n69567 , n69569 );
xnor ( n69571 , n69570 , n64624 );
and ( n69572 , n69565 , n69571 );
buf ( n69573 , n64558 );
and ( n69574 , n69573 , n64612 );
and ( n69575 , n69571 , n69574 );
and ( n69576 , n69565 , n69574 );
or ( n69577 , n69572 , n69575 , n69576 );
and ( n69578 , n68444 , n64789 );
and ( n69579 , n68439 , n64787 );
nor ( n69580 , n69578 , n69579 );
xnor ( n69581 , n69580 , n64738 );
and ( n69582 , n69577 , n69581 );
and ( n69583 , n68837 , n64711 );
and ( n69584 , n68625 , n64709 );
nor ( n69585 , n69583 , n69584 );
xnor ( n69586 , n69585 , n64682 );
and ( n69587 , n69581 , n69586 );
and ( n69588 , n69577 , n69586 );
or ( n69589 , n69582 , n69587 , n69588 );
and ( n69590 , n68192 , n64897 );
and ( n69591 , n67873 , n64895 );
nor ( n69592 , n69590 , n69591 );
xnor ( n69593 , n69592 , n64850 );
and ( n69594 , n69589 , n69593 );
and ( n69595 , n68873 , n64652 );
and ( n69596 , n68837 , n64650 );
nor ( n69597 , n69595 , n69596 );
xnor ( n69598 , n69597 , n64609 );
and ( n69599 , n69449 , n64617 );
and ( n69600 , n69095 , n64615 );
nor ( n69601 , n69599 , n69600 );
xnor ( n69602 , n69601 , n64624 );
xor ( n69603 , n69598 , n69602 );
and ( n69604 , n69568 , n64612 );
xor ( n69605 , n69603 , n69604 );
and ( n69606 , n69593 , n69605 );
and ( n69607 , n69589 , n69605 );
or ( n69608 , n69594 , n69606 , n69607 );
and ( n69609 , n67727 , n65056 );
and ( n69610 , n67548 , n65054 );
nor ( n69611 , n69609 , n69610 );
xnor ( n69612 , n69611 , n64943 );
and ( n69613 , n69608 , n69612 );
and ( n69614 , n69598 , n69602 );
and ( n69615 , n69602 , n69604 );
and ( n69616 , n69598 , n69604 );
or ( n69617 , n69614 , n69615 , n69616 );
and ( n69618 , n68837 , n64652 );
and ( n69619 , n68625 , n64650 );
nor ( n69620 , n69618 , n69619 );
xnor ( n69621 , n69620 , n64609 );
xor ( n69622 , n69617 , n69621 );
xor ( n69623 , n69443 , n69447 );
xor ( n69624 , n69623 , n69450 );
xor ( n69625 , n69622 , n69624 );
and ( n69626 , n69612 , n69625 );
and ( n69627 , n69608 , n69625 );
or ( n69628 , n69613 , n69626 , n69627 );
and ( n69629 , n67302 , n65183 );
and ( n69630 , n67111 , n65181 );
nor ( n69631 , n69629 , n69630 );
xnor ( n69632 , n69631 , n64994 );
and ( n69633 , n69628 , n69632 );
xor ( n69634 , n69243 , n69244 );
and ( n69635 , n69617 , n69621 );
and ( n69636 , n69621 , n69624 );
and ( n69637 , n69617 , n69624 );
or ( n69638 , n69635 , n69636 , n69637 );
xor ( n69639 , n69634 , n69638 );
and ( n69640 , n68192 , n64789 );
and ( n69641 , n67873 , n64787 );
nor ( n69642 , n69640 , n69641 );
xnor ( n69643 , n69642 , n64738 );
xor ( n69644 , n69639 , n69643 );
and ( n69645 , n69632 , n69644 );
and ( n69646 , n69628 , n69644 );
or ( n69647 , n69633 , n69645 , n69646 );
and ( n69648 , n66786 , n65371 );
and ( n69649 , n66781 , n65369 );
nor ( n69650 , n69648 , n69649 );
xnor ( n69651 , n69650 , n65168 );
and ( n69652 , n69647 , n69651 );
and ( n69653 , n69634 , n69638 );
and ( n69654 , n69638 , n69643 );
and ( n69655 , n69634 , n69643 );
or ( n69656 , n69653 , n69654 , n69655 );
and ( n69657 , n67307 , n65056 );
and ( n69658 , n67302 , n65054 );
nor ( n69659 , n69657 , n69658 );
xnor ( n69660 , n69659 , n64943 );
xor ( n69661 , n69656 , n69660 );
xor ( n69662 , n69245 , n69249 );
xor ( n69663 , n69662 , n69254 );
xor ( n69664 , n69661 , n69663 );
and ( n69665 , n69651 , n69664 );
and ( n69666 , n69647 , n69664 );
or ( n69667 , n69652 , n69665 , n69666 );
and ( n69668 , n65883 , n66241 );
and ( n69669 , n65698 , n66239 );
nor ( n69670 , n69668 , n69669 );
xnor ( n69671 , n69670 , n65876 );
and ( n69672 , n69667 , n69671 );
xor ( n69673 , n69489 , n69493 );
xor ( n69674 , n69673 , n69496 );
and ( n69675 , n69671 , n69674 );
and ( n69676 , n69667 , n69674 );
or ( n69677 , n69672 , n69675 , n69676 );
and ( n69678 , n65443 , n66657 );
and ( n69679 , n65453 , n66655 );
nor ( n69680 , n69678 , n69679 );
xnor ( n69681 , n69680 , n66130 );
and ( n69682 , n69677 , n69681 );
xor ( n69683 , n69485 , n69499 );
xor ( n69684 , n69683 , n69504 );
and ( n69685 , n69681 , n69684 );
and ( n69686 , n69677 , n69684 );
or ( n69687 , n69682 , n69685 , n69686 );
and ( n69688 , n65001 , n67498 );
and ( n69689 , n64955 , n67495 );
nor ( n69690 , n69688 , n69689 );
xnor ( n69691 , n69690 , n66511 );
and ( n69692 , n69687 , n69691 );
xor ( n69693 , n69425 , n69427 );
xor ( n69694 , n69693 , n69430 );
and ( n69695 , n69691 , n69694 );
and ( n69696 , n69687 , n69694 );
or ( n69697 , n69692 , n69695 , n69696 );
and ( n69698 , n64955 , n67498 );
and ( n69699 , n64950 , n67495 );
nor ( n69700 , n69698 , n69699 );
xnor ( n69701 , n69700 , n66511 );
and ( n69702 , n69697 , n69701 );
xor ( n69703 , n69421 , n69433 );
xor ( n69704 , n69703 , n69436 );
and ( n69705 , n69701 , n69704 );
and ( n69706 , n69697 , n69704 );
or ( n69707 , n69702 , n69705 , n69706 );
and ( n69708 , n69656 , n69660 );
and ( n69709 , n69660 , n69663 );
and ( n69710 , n69656 , n69663 );
or ( n69711 , n69708 , n69709 , n69710 );
and ( n69712 , n66517 , n65550 );
and ( n69713 , n66266 , n65548 );
nor ( n69714 , n69712 , n69713 );
xnor ( n69715 , n69714 , n65313 );
and ( n69716 , n69711 , n69715 );
xor ( n69717 , n69475 , n69479 );
xor ( n69718 , n69717 , n69482 );
and ( n69719 , n69715 , n69718 );
and ( n69720 , n69711 , n69718 );
or ( n69721 , n69716 , n69719 , n69720 );
and ( n69722 , n65698 , n66241 );
and ( n69723 , n65657 , n66239 );
nor ( n69724 , n69722 , n69723 );
xnor ( n69725 , n69724 , n65876 );
and ( n69726 , n69721 , n69725 );
and ( n69727 , n66142 , n65756 );
and ( n69728 , n66137 , n65754 );
nor ( n69729 , n69727 , n69728 );
xnor ( n69730 , n69729 , n65450 );
and ( n69731 , n69725 , n69730 );
and ( n69732 , n69721 , n69730 );
or ( n69733 , n69726 , n69731 , n69732 );
and ( n69734 , n65175 , n67160 );
and ( n69735 , n65135 , n67158 );
nor ( n69736 , n69734 , n69735 );
xnor ( n69737 , n69736 , n66514 );
and ( n69738 , n69733 , n69737 );
xor ( n69739 , n69409 , n69413 );
xor ( n69740 , n69739 , n69418 );
and ( n69741 , n69737 , n69740 );
and ( n69742 , n69733 , n69740 );
or ( n69743 , n69738 , n69741 , n69742 );
xor ( n69744 , n69527 , n69531 );
xor ( n69745 , n69744 , n69534 );
and ( n69746 , n69743 , n69745 );
xor ( n69747 , n69377 , n69381 );
xor ( n69748 , n69747 , n69384 );
and ( n69749 , n69745 , n69748 );
and ( n69750 , n69743 , n69748 );
or ( n69751 , n69746 , n69749 , n69750 );
and ( n69752 , n69707 , n69751 );
xor ( n69753 , n69439 , n69537 );
xor ( n69754 , n69753 , n69540 );
and ( n69755 , n69751 , n69754 );
and ( n69756 , n69707 , n69754 );
or ( n69757 , n69752 , n69755 , n69756 );
xor ( n69758 , n69395 , n69543 );
xor ( n69759 , n69758 , n69546 );
and ( n69760 , n69757 , n69759 );
xor ( n69761 , n69345 , n69347 );
xor ( n69762 , n69761 , n69350 );
and ( n69763 , n69759 , n69762 );
and ( n69764 , n69757 , n69762 );
or ( n69765 , n69760 , n69763 , n69764 );
and ( n69766 , n69561 , n69765 );
xor ( n69767 , n69561 , n69765 );
xor ( n69768 , n69757 , n69759 );
xor ( n69769 , n69768 , n69762 );
and ( n69770 , n69095 , n64652 );
and ( n69771 , n68873 , n64650 );
nor ( n69772 , n69770 , n69771 );
xnor ( n69773 , n69772 , n64609 );
and ( n69774 , n69568 , n64617 );
and ( n69775 , n69449 , n64615 );
nor ( n69776 , n69774 , n69775 );
xnor ( n69777 , n69776 , n64624 );
and ( n69778 , n69773 , n69777 );
and ( n69779 , n69566 , n64612 );
and ( n69780 , n69777 , n69779 );
and ( n69781 , n69773 , n69779 );
or ( n69782 , n69778 , n69780 , n69781 );
and ( n69783 , n68439 , n64789 );
and ( n69784 , n68199 , n64787 );
nor ( n69785 , n69783 , n69784 );
xnor ( n69786 , n69785 , n64738 );
and ( n69787 , n69782 , n69786 );
and ( n69788 , n68625 , n64711 );
and ( n69789 , n68444 , n64709 );
nor ( n69790 , n69788 , n69789 );
xnor ( n69791 , n69790 , n64682 );
and ( n69792 , n69786 , n69791 );
and ( n69793 , n69782 , n69791 );
or ( n69794 , n69787 , n69792 , n69793 );
and ( n69795 , n67873 , n64897 );
and ( n69796 , n67833 , n64895 );
nor ( n69797 , n69795 , n69796 );
xnor ( n69798 , n69797 , n64850 );
and ( n69799 , n69794 , n69798 );
and ( n69800 , n68199 , n64789 );
and ( n69801 , n68192 , n64787 );
nor ( n69802 , n69800 , n69801 );
xnor ( n69803 , n69802 , n64738 );
and ( n69804 , n69798 , n69803 );
and ( n69805 , n69794 , n69803 );
or ( n69806 , n69799 , n69804 , n69805 );
and ( n69807 , n67548 , n65056 );
and ( n69808 , n67307 , n65054 );
nor ( n69809 , n69807 , n69808 );
xnor ( n69810 , n69809 , n64943 );
and ( n69811 , n69806 , n69810 );
xor ( n69812 , n69453 , n69457 );
xor ( n69813 , n69812 , n69462 );
and ( n69814 , n69810 , n69813 );
and ( n69815 , n69806 , n69813 );
or ( n69816 , n69811 , n69814 , n69815 );
and ( n69817 , n67111 , n65183 );
and ( n69818 , n66981 , n65181 );
nor ( n69819 , n69817 , n69818 );
xnor ( n69820 , n69819 , n64994 );
and ( n69821 , n69816 , n69820 );
xor ( n69822 , n69465 , n69469 );
xor ( n69823 , n69822 , n69472 );
and ( n69824 , n69820 , n69823 );
and ( n69825 , n69816 , n69823 );
or ( n69826 , n69821 , n69824 , n69825 );
and ( n69827 , n66137 , n66016 );
and ( n69828 , n65935 , n66014 );
nor ( n69829 , n69827 , n69828 );
xnor ( n69830 , n69829 , n65650 );
and ( n69831 , n69826 , n69830 );
and ( n69832 , n66276 , n65756 );
and ( n69833 , n66142 , n65754 );
nor ( n69834 , n69832 , n69833 );
xnor ( n69835 , n69834 , n65450 );
and ( n69836 , n69830 , n69835 );
and ( n69837 , n69826 , n69835 );
or ( n69838 , n69831 , n69836 , n69837 );
xor ( n69839 , n69721 , n69725 );
xor ( n69840 , n69839 , n69730 );
and ( n69841 , n69838 , n69840 );
xor ( n69842 , n69511 , n69513 );
xor ( n69843 , n69842 , n69516 );
and ( n69844 , n69840 , n69843 );
and ( n69845 , n69838 , n69843 );
or ( n69846 , n69841 , n69844 , n69845 );
and ( n69847 , n65363 , n66906 );
and ( n69848 , n65265 , n66904 );
nor ( n69849 , n69847 , n69848 );
xnor ( n69850 , n69849 , n66286 );
and ( n69851 , n69846 , n69850 );
xor ( n69852 , n69507 , n69519 );
xor ( n69853 , n69852 , n69524 );
and ( n69854 , n69850 , n69853 );
and ( n69855 , n69846 , n69853 );
or ( n69856 , n69851 , n69854 , n69855 );
and ( n69857 , n66781 , n65550 );
and ( n69858 , n66507 , n65548 );
nor ( n69859 , n69857 , n69858 );
xnor ( n69860 , n69859 , n65313 );
and ( n69861 , n66981 , n65371 );
and ( n69862 , n66786 , n65369 );
nor ( n69863 , n69861 , n69862 );
xnor ( n69864 , n69863 , n65168 );
and ( n69865 , n69860 , n69864 );
xor ( n69866 , n69806 , n69810 );
xor ( n69867 , n69866 , n69813 );
and ( n69868 , n69864 , n69867 );
and ( n69869 , n69860 , n69867 );
or ( n69870 , n69865 , n69868 , n69869 );
and ( n69871 , n65935 , n66241 );
and ( n69872 , n65883 , n66239 );
nor ( n69873 , n69871 , n69872 );
xnor ( n69874 , n69873 , n65876 );
and ( n69875 , n69870 , n69874 );
xor ( n69876 , n69647 , n69651 );
xor ( n69877 , n69876 , n69664 );
and ( n69878 , n69874 , n69877 );
and ( n69879 , n69870 , n69877 );
or ( n69880 , n69875 , n69878 , n69879 );
and ( n69881 , n65657 , n66657 );
and ( n69882 , n65443 , n66655 );
nor ( n69883 , n69881 , n69882 );
xnor ( n69884 , n69883 , n66130 );
and ( n69885 , n69880 , n69884 );
xor ( n69886 , n69826 , n69830 );
xor ( n69887 , n69886 , n69835 );
and ( n69888 , n69884 , n69887 );
and ( n69889 , n69880 , n69887 );
or ( n69890 , n69885 , n69888 , n69889 );
and ( n69891 , n66266 , n65756 );
and ( n69892 , n66276 , n65754 );
nor ( n69893 , n69891 , n69892 );
xnor ( n69894 , n69893 , n65450 );
and ( n69895 , n66507 , n65550 );
and ( n69896 , n66517 , n65548 );
nor ( n69897 , n69895 , n69896 );
xnor ( n69898 , n69897 , n65313 );
and ( n69899 , n69894 , n69898 );
xor ( n69900 , n69816 , n69820 );
xor ( n69901 , n69900 , n69823 );
and ( n69902 , n69898 , n69901 );
and ( n69903 , n69894 , n69901 );
or ( n69904 , n69899 , n69902 , n69903 );
and ( n69905 , n65453 , n66906 );
and ( n69906 , n65306 , n66904 );
nor ( n69907 , n69905 , n69906 );
xnor ( n69908 , n69907 , n66286 );
and ( n69909 , n69904 , n69908 );
xor ( n69910 , n69711 , n69715 );
xor ( n69911 , n69910 , n69718 );
and ( n69912 , n69908 , n69911 );
and ( n69913 , n69904 , n69911 );
or ( n69914 , n69909 , n69912 , n69913 );
and ( n69915 , n69890 , n69914 );
and ( n69916 , n65265 , n67160 );
and ( n69917 , n65175 , n67158 );
nor ( n69918 , n69916 , n69917 );
xnor ( n69919 , n69918 , n66514 );
and ( n69920 , n69914 , n69919 );
and ( n69921 , n69890 , n69919 );
or ( n69922 , n69915 , n69920 , n69921 );
and ( n69923 , n65135 , n67498 );
and ( n69924 , n65001 , n67495 );
nor ( n69925 , n69923 , n69924 );
xnor ( n69926 , n69925 , n66511 );
and ( n69927 , n65306 , n66906 );
and ( n69928 , n65363 , n66904 );
nor ( n69929 , n69927 , n69928 );
xnor ( n69930 , n69929 , n66286 );
and ( n69931 , n69926 , n69930 );
xor ( n69932 , n69677 , n69681 );
xor ( n69933 , n69932 , n69684 );
and ( n69934 , n69930 , n69933 );
and ( n69935 , n69926 , n69933 );
or ( n69936 , n69931 , n69934 , n69935 );
and ( n69937 , n69922 , n69936 );
xor ( n69938 , n69733 , n69737 );
xor ( n69939 , n69938 , n69740 );
and ( n69940 , n69936 , n69939 );
and ( n69941 , n69922 , n69939 );
or ( n69942 , n69937 , n69940 , n69941 );
and ( n69943 , n69856 , n69942 );
xor ( n69944 , n69697 , n69701 );
xor ( n69945 , n69944 , n69704 );
and ( n69946 , n69942 , n69945 );
and ( n69947 , n69856 , n69945 );
or ( n69948 , n69943 , n69946 , n69947 );
xor ( n69949 , n69387 , n69389 );
xor ( n69950 , n69949 , n69392 );
and ( n69951 , n69948 , n69950 );
xor ( n69952 , n69707 , n69751 );
xor ( n69953 , n69952 , n69754 );
and ( n69954 , n69950 , n69953 );
and ( n69955 , n69948 , n69953 );
or ( n69956 , n69951 , n69954 , n69955 );
and ( n69957 , n69769 , n69956 );
xor ( n69958 , n69769 , n69956 );
xor ( n69959 , n69948 , n69950 );
xor ( n69960 , n69959 , n69953 );
and ( n69961 , n65175 , n67498 );
and ( n69962 , n65135 , n67495 );
nor ( n69963 , n69961 , n69962 );
xnor ( n69964 , n69963 , n66511 );
and ( n69965 , n65363 , n67160 );
and ( n69966 , n65265 , n67158 );
nor ( n69967 , n69965 , n69966 );
xnor ( n69968 , n69967 , n66514 );
and ( n69969 , n69964 , n69968 );
xor ( n69970 , n69904 , n69908 );
xor ( n69971 , n69970 , n69911 );
and ( n69972 , n69968 , n69971 );
and ( n69973 , n69964 , n69971 );
or ( n69974 , n69969 , n69972 , n69973 );
and ( n69975 , n69566 , n64652 );
and ( n69976 , n69568 , n64650 );
nor ( n69977 , n69975 , n69976 );
xnor ( n69978 , n69977 , n64609 );
buf ( n69979 , n64559 );
and ( n69980 , n69979 , n64617 );
and ( n69981 , n69573 , n64615 );
nor ( n69982 , n69980 , n69981 );
xnor ( n69983 , n69982 , n64624 );
and ( n69984 , n69978 , n69983 );
buf ( n69985 , n64560 );
and ( n69986 , n69985 , n64612 );
and ( n69987 , n69983 , n69986 );
and ( n69988 , n69978 , n69986 );
or ( n69989 , n69984 , n69987 , n69988 );
and ( n69990 , n69573 , n64617 );
and ( n69991 , n69566 , n64615 );
nor ( n69992 , n69990 , n69991 );
xnor ( n69993 , n69992 , n64624 );
and ( n69994 , n69989 , n69993 );
and ( n69995 , n69979 , n64612 );
and ( n69996 , n69993 , n69995 );
and ( n69997 , n69989 , n69995 );
or ( n69998 , n69994 , n69996 , n69997 );
and ( n69999 , n68625 , n64789 );
and ( n70000 , n68444 , n64787 );
nor ( n70001 , n69999 , n70000 );
xnor ( n70002 , n70001 , n64738 );
and ( n70003 , n69998 , n70002 );
and ( n70004 , n69449 , n64652 );
and ( n70005 , n69095 , n64650 );
nor ( n70006 , n70004 , n70005 );
xnor ( n70007 , n70006 , n64609 );
and ( n70008 , n70002 , n70007 );
and ( n70009 , n69998 , n70007 );
or ( n70010 , n70003 , n70008 , n70009 );
and ( n70011 , n69095 , n64711 );
and ( n70012 , n68873 , n64709 );
nor ( n70013 , n70011 , n70012 );
xnor ( n70014 , n70013 , n64682 );
and ( n70015 , n69568 , n64652 );
and ( n70016 , n69449 , n64650 );
nor ( n70017 , n70015 , n70016 );
xnor ( n70018 , n70017 , n64609 );
and ( n70019 , n70014 , n70018 );
xor ( n70020 , n69989 , n69993 );
xor ( n70021 , n70020 , n69995 );
and ( n70022 , n70018 , n70021 );
and ( n70023 , n70014 , n70021 );
or ( n70024 , n70019 , n70022 , n70023 );
and ( n70025 , n68439 , n64897 );
and ( n70026 , n68199 , n64895 );
nor ( n70027 , n70025 , n70026 );
xnor ( n70028 , n70027 , n64850 );
and ( n70029 , n70024 , n70028 );
xor ( n70030 , n69565 , n69571 );
xor ( n70031 , n70030 , n69574 );
and ( n70032 , n70028 , n70031 );
and ( n70033 , n70024 , n70031 );
or ( n70034 , n70029 , n70032 , n70033 );
and ( n70035 , n70010 , n70034 );
xor ( n70036 , n69773 , n69777 );
xor ( n70037 , n70036 , n69779 );
and ( n70038 , n70034 , n70037 );
and ( n70039 , n70010 , n70037 );
or ( n70040 , n70035 , n70038 , n70039 );
and ( n70041 , n67833 , n65056 );
and ( n70042 , n67727 , n65054 );
nor ( n70043 , n70041 , n70042 );
xnor ( n70044 , n70043 , n64943 );
and ( n70045 , n70040 , n70044 );
xor ( n70046 , n69782 , n69786 );
xor ( n70047 , n70046 , n69791 );
and ( n70048 , n70044 , n70047 );
and ( n70049 , n70040 , n70047 );
or ( n70050 , n70045 , n70048 , n70049 );
and ( n70051 , n67307 , n65183 );
and ( n70052 , n67302 , n65181 );
nor ( n70053 , n70051 , n70052 );
xnor ( n70054 , n70053 , n64994 );
and ( n70055 , n70050 , n70054 );
xor ( n70056 , n69794 , n69798 );
xor ( n70057 , n70056 , n69803 );
and ( n70058 , n70054 , n70057 );
and ( n70059 , n70050 , n70057 );
or ( n70060 , n70055 , n70058 , n70059 );
and ( n70061 , n66276 , n66016 );
and ( n70062 , n66142 , n66014 );
nor ( n70063 , n70061 , n70062 );
xnor ( n70064 , n70063 , n65650 );
and ( n70065 , n70060 , n70064 );
xor ( n70066 , n69628 , n69632 );
xor ( n70067 , n70066 , n69644 );
and ( n70068 , n70064 , n70067 );
and ( n70069 , n70060 , n70067 );
or ( n70070 , n70065 , n70068 , n70069 );
and ( n70071 , n65698 , n66657 );
and ( n70072 , n65657 , n66655 );
nor ( n70073 , n70071 , n70072 );
xnor ( n70074 , n70073 , n66130 );
and ( n70075 , n70070 , n70074 );
and ( n70076 , n66142 , n66016 );
and ( n70077 , n66137 , n66014 );
nor ( n70078 , n70076 , n70077 );
xnor ( n70079 , n70078 , n65650 );
and ( n70080 , n70074 , n70079 );
and ( n70081 , n70070 , n70079 );
or ( n70082 , n70075 , n70080 , n70081 );
and ( n70083 , n66507 , n65756 );
and ( n70084 , n66517 , n65754 );
nor ( n70085 , n70083 , n70084 );
xnor ( n70086 , n70085 , n65450 );
and ( n70087 , n66786 , n65550 );
and ( n70088 , n66781 , n65548 );
nor ( n70089 , n70087 , n70088 );
xnor ( n70090 , n70089 , n65313 );
and ( n70091 , n70086 , n70090 );
xor ( n70092 , n70050 , n70054 );
xor ( n70093 , n70092 , n70057 );
and ( n70094 , n70090 , n70093 );
and ( n70095 , n70086 , n70093 );
or ( n70096 , n70091 , n70094 , n70095 );
and ( n70097 , n65883 , n66657 );
and ( n70098 , n65698 , n66655 );
nor ( n70099 , n70097 , n70098 );
xnor ( n70100 , n70099 , n66130 );
and ( n70101 , n70096 , n70100 );
xor ( n70102 , n69860 , n69864 );
xor ( n70103 , n70102 , n69867 );
and ( n70104 , n70100 , n70103 );
and ( n70105 , n70096 , n70103 );
or ( n70106 , n70101 , n70104 , n70105 );
and ( n70107 , n65443 , n66906 );
and ( n70108 , n65453 , n66904 );
nor ( n70109 , n70107 , n70108 );
xnor ( n70110 , n70109 , n66286 );
and ( n70111 , n70106 , n70110 );
xor ( n70112 , n69894 , n69898 );
xor ( n70113 , n70112 , n69901 );
and ( n70114 , n70110 , n70113 );
and ( n70115 , n70106 , n70113 );
or ( n70116 , n70111 , n70114 , n70115 );
and ( n70117 , n70082 , n70116 );
xor ( n70118 , n69667 , n69671 );
xor ( n70119 , n70118 , n69674 );
and ( n70120 , n70116 , n70119 );
and ( n70121 , n70082 , n70119 );
or ( n70122 , n70117 , n70120 , n70121 );
and ( n70123 , n69974 , n70122 );
xor ( n70124 , n69838 , n69840 );
xor ( n70125 , n70124 , n69843 );
and ( n70126 , n70122 , n70125 );
and ( n70127 , n69974 , n70125 );
or ( n70128 , n70123 , n70126 , n70127 );
xor ( n70129 , n69846 , n69850 );
xor ( n70130 , n70129 , n69853 );
and ( n70131 , n70128 , n70130 );
xor ( n70132 , n69687 , n69691 );
xor ( n70133 , n70132 , n69694 );
and ( n70134 , n70130 , n70133 );
and ( n70135 , n70128 , n70133 );
or ( n70136 , n70131 , n70134 , n70135 );
xor ( n70137 , n69856 , n69942 );
xor ( n70138 , n70137 , n69945 );
and ( n70139 , n70136 , n70138 );
xor ( n70140 , n69743 , n69745 );
xor ( n70141 , n70140 , n69748 );
and ( n70142 , n70138 , n70141 );
and ( n70143 , n70136 , n70141 );
or ( n70144 , n70139 , n70142 , n70143 );
and ( n70145 , n69960 , n70144 );
xor ( n70146 , n69960 , n70144 );
xor ( n70147 , n70136 , n70138 );
xor ( n70148 , n70147 , n70141 );
and ( n70149 , n66781 , n65756 );
and ( n70150 , n66507 , n65754 );
nor ( n70151 , n70149 , n70150 );
xnor ( n70152 , n70151 , n65450 );
and ( n70153 , n66981 , n65550 );
and ( n70154 , n66786 , n65548 );
nor ( n70155 , n70153 , n70154 );
xnor ( n70156 , n70155 , n65313 );
and ( n70157 , n70152 , n70156 );
and ( n70158 , n67873 , n65056 );
and ( n70159 , n67833 , n65054 );
nor ( n70160 , n70158 , n70159 );
xnor ( n70161 , n70160 , n64943 );
and ( n70162 , n68199 , n64897 );
and ( n70163 , n68192 , n64895 );
nor ( n70164 , n70162 , n70163 );
xnor ( n70165 , n70164 , n64850 );
and ( n70166 , n70161 , n70165 );
xor ( n70167 , n69577 , n69581 );
xor ( n70168 , n70167 , n69586 );
and ( n70169 , n70165 , n70168 );
and ( n70170 , n70161 , n70168 );
or ( n70171 , n70166 , n70169 , n70170 );
and ( n70172 , n67302 , n65371 );
and ( n70173 , n67111 , n65369 );
nor ( n70174 , n70172 , n70173 );
xnor ( n70175 , n70174 , n65168 );
xor ( n70176 , n70171 , n70175 );
and ( n70177 , n67548 , n65183 );
and ( n70178 , n67307 , n65181 );
nor ( n70179 , n70177 , n70178 );
xnor ( n70180 , n70179 , n64994 );
xor ( n70181 , n70176 , n70180 );
and ( n70182 , n70156 , n70181 );
and ( n70183 , n70152 , n70181 );
or ( n70184 , n70157 , n70182 , n70183 );
and ( n70185 , n65935 , n66657 );
and ( n70186 , n65883 , n66655 );
nor ( n70187 , n70185 , n70186 );
xnor ( n70188 , n70187 , n66130 );
and ( n70189 , n70184 , n70188 );
and ( n70190 , n66142 , n66241 );
and ( n70191 , n66137 , n66239 );
nor ( n70192 , n70190 , n70191 );
xnor ( n70193 , n70192 , n65876 );
and ( n70194 , n70188 , n70193 );
and ( n70195 , n70184 , n70193 );
or ( n70196 , n70189 , n70194 , n70195 );
and ( n70197 , n65453 , n67160 );
and ( n70198 , n65306 , n67158 );
nor ( n70199 , n70197 , n70198 );
xnor ( n70200 , n70199 , n66514 );
and ( n70201 , n70196 , n70200 );
and ( n70202 , n70171 , n70175 );
and ( n70203 , n70175 , n70180 );
and ( n70204 , n70171 , n70180 );
or ( n70205 , n70202 , n70203 , n70204 );
and ( n70206 , n67111 , n65371 );
and ( n70207 , n66981 , n65369 );
nor ( n70208 , n70206 , n70207 );
xnor ( n70209 , n70208 , n65168 );
and ( n70210 , n70205 , n70209 );
xor ( n70211 , n69608 , n69612 );
xor ( n70212 , n70211 , n69625 );
and ( n70213 , n70209 , n70212 );
and ( n70214 , n70205 , n70212 );
or ( n70215 , n70210 , n70213 , n70214 );
and ( n70216 , n66137 , n66241 );
and ( n70217 , n65935 , n66239 );
nor ( n70218 , n70216 , n70217 );
xnor ( n70219 , n70218 , n65876 );
xor ( n70220 , n70215 , n70219 );
and ( n70221 , n66517 , n65756 );
and ( n70222 , n66266 , n65754 );
nor ( n70223 , n70221 , n70222 );
xnor ( n70224 , n70223 , n65450 );
xor ( n70225 , n70220 , n70224 );
and ( n70226 , n70200 , n70225 );
and ( n70227 , n70196 , n70225 );
or ( n70228 , n70201 , n70226 , n70227 );
and ( n70229 , n69573 , n64652 );
and ( n70230 , n69566 , n64650 );
nor ( n70231 , n70229 , n70230 );
xnor ( n70232 , n70231 , n64609 );
and ( n70233 , n69985 , n64617 );
and ( n70234 , n69979 , n64615 );
nor ( n70235 , n70233 , n70234 );
xnor ( n70236 , n70235 , n64624 );
and ( n70237 , n70232 , n70236 );
buf ( n70238 , n64561 );
and ( n70239 , n70238 , n64612 );
and ( n70240 , n70236 , n70239 );
and ( n70241 , n70232 , n70239 );
or ( n70242 , n70237 , n70240 , n70241 );
and ( n70243 , n69979 , n64652 );
and ( n70244 , n69573 , n64650 );
nor ( n70245 , n70243 , n70244 );
xnor ( n70246 , n70245 , n64609 );
and ( n70247 , n70238 , n64617 );
and ( n70248 , n69985 , n64615 );
nor ( n70249 , n70247 , n70248 );
xnor ( n70250 , n70249 , n64624 );
and ( n70251 , n70246 , n70250 );
buf ( n70252 , n64562 );
and ( n70253 , n70252 , n64612 );
and ( n70254 , n70250 , n70253 );
and ( n70255 , n70246 , n70253 );
or ( n70256 , n70251 , n70254 , n70255 );
and ( n70257 , n69985 , n64652 );
and ( n70258 , n69979 , n64650 );
nor ( n70259 , n70257 , n70258 );
xnor ( n70260 , n70259 , n64609 );
and ( n70261 , n70252 , n64617 );
and ( n70262 , n70238 , n64615 );
nor ( n70263 , n70261 , n70262 );
xnor ( n70264 , n70263 , n64624 );
and ( n70265 , n70260 , n70264 );
buf ( n70266 , n64563 );
and ( n70267 , n70266 , n64612 );
and ( n70268 , n70264 , n70267 );
and ( n70269 , n70260 , n70267 );
or ( n70270 , n70265 , n70268 , n70269 );
and ( n70271 , n69566 , n64711 );
and ( n70272 , n69568 , n64709 );
nor ( n70273 , n70271 , n70272 );
xnor ( n70274 , n70273 , n64682 );
and ( n70275 , n70270 , n70274 );
xor ( n70276 , n70246 , n70250 );
xor ( n70277 , n70276 , n70253 );
and ( n70278 , n70274 , n70277 );
and ( n70279 , n70270 , n70277 );
or ( n70280 , n70275 , n70278 , n70279 );
and ( n70281 , n70256 , n70280 );
xor ( n70282 , n70232 , n70236 );
xor ( n70283 , n70282 , n70239 );
and ( n70284 , n70280 , n70283 );
and ( n70285 , n70256 , n70283 );
or ( n70286 , n70281 , n70284 , n70285 );
and ( n70287 , n70242 , n70286 );
xor ( n70288 , n69978 , n69983 );
xor ( n70289 , n70288 , n69986 );
and ( n70290 , n70286 , n70289 );
and ( n70291 , n70242 , n70289 );
or ( n70292 , n70287 , n70290 , n70291 );
and ( n70293 , n68444 , n64897 );
and ( n70294 , n68439 , n64895 );
nor ( n70295 , n70293 , n70294 );
xnor ( n70296 , n70295 , n64850 );
and ( n70297 , n70292 , n70296 );
and ( n70298 , n68837 , n64789 );
and ( n70299 , n68625 , n64787 );
nor ( n70300 , n70298 , n70299 );
xnor ( n70301 , n70300 , n64738 );
and ( n70302 , n70296 , n70301 );
and ( n70303 , n70292 , n70301 );
or ( n70304 , n70297 , n70302 , n70303 );
and ( n70305 , n68192 , n65056 );
and ( n70306 , n67873 , n65054 );
nor ( n70307 , n70305 , n70306 );
xnor ( n70308 , n70307 , n64943 );
and ( n70309 , n70304 , n70308 );
xor ( n70310 , n69998 , n70002 );
xor ( n70311 , n70310 , n70007 );
and ( n70312 , n70308 , n70311 );
and ( n70313 , n70304 , n70311 );
or ( n70314 , n70309 , n70312 , n70313 );
and ( n70315 , n67727 , n65183 );
and ( n70316 , n67548 , n65181 );
nor ( n70317 , n70315 , n70316 );
xnor ( n70318 , n70317 , n64994 );
and ( n70319 , n70314 , n70318 );
xor ( n70320 , n70010 , n70034 );
xor ( n70321 , n70320 , n70037 );
and ( n70322 , n70318 , n70321 );
and ( n70323 , n70314 , n70321 );
or ( n70324 , n70319 , n70322 , n70323 );
xor ( n70325 , n69589 , n69593 );
xor ( n70326 , n70325 , n69605 );
and ( n70327 , n70324 , n70326 );
xor ( n70328 , n70040 , n70044 );
xor ( n70329 , n70328 , n70047 );
and ( n70330 , n70326 , n70329 );
and ( n70331 , n70324 , n70329 );
or ( n70332 , n70327 , n70330 , n70331 );
and ( n70333 , n66266 , n66016 );
and ( n70334 , n66276 , n66014 );
nor ( n70335 , n70333 , n70334 );
xnor ( n70336 , n70335 , n65650 );
and ( n70337 , n70332 , n70336 );
xor ( n70338 , n70205 , n70209 );
xor ( n70339 , n70338 , n70212 );
and ( n70340 , n70336 , n70339 );
and ( n70341 , n70332 , n70339 );
or ( n70342 , n70337 , n70340 , n70341 );
and ( n70343 , n65657 , n66906 );
and ( n70344 , n65443 , n66904 );
nor ( n70345 , n70343 , n70344 );
xnor ( n70346 , n70345 , n66286 );
and ( n70347 , n70342 , n70346 );
xor ( n70348 , n70060 , n70064 );
xor ( n70349 , n70348 , n70067 );
and ( n70350 , n70346 , n70349 );
and ( n70351 , n70342 , n70349 );
or ( n70352 , n70347 , n70350 , n70351 );
and ( n70353 , n70228 , n70352 );
and ( n70354 , n65306 , n67160 );
and ( n70355 , n65363 , n67158 );
nor ( n70356 , n70354 , n70355 );
xnor ( n70357 , n70356 , n66514 );
and ( n70358 , n70352 , n70357 );
and ( n70359 , n70228 , n70357 );
or ( n70360 , n70353 , n70358 , n70359 );
and ( n70361 , n70215 , n70219 );
and ( n70362 , n70219 , n70224 );
and ( n70363 , n70215 , n70224 );
or ( n70364 , n70361 , n70362 , n70363 );
xor ( n70365 , n70070 , n70074 );
xor ( n70366 , n70365 , n70079 );
and ( n70367 , n70364 , n70366 );
xor ( n70368 , n69870 , n69874 );
xor ( n70369 , n70368 , n69877 );
and ( n70370 , n70366 , n70369 );
and ( n70371 , n70364 , n70369 );
or ( n70372 , n70367 , n70370 , n70371 );
and ( n70373 , n70360 , n70372 );
xor ( n70374 , n69880 , n69884 );
xor ( n70375 , n70374 , n69887 );
and ( n70376 , n70372 , n70375 );
and ( n70377 , n70360 , n70375 );
or ( n70378 , n70373 , n70376 , n70377 );
xor ( n70379 , n69890 , n69914 );
xor ( n70380 , n70379 , n69919 );
and ( n70381 , n70378 , n70380 );
xor ( n70382 , n69926 , n69930 );
xor ( n70383 , n70382 , n69933 );
and ( n70384 , n70380 , n70383 );
and ( n70385 , n70378 , n70383 );
or ( n70386 , n70381 , n70384 , n70385 );
xor ( n70387 , n69922 , n69936 );
xor ( n70388 , n70387 , n69939 );
and ( n70389 , n70386 , n70388 );
xor ( n70390 , n70128 , n70130 );
xor ( n70391 , n70390 , n70133 );
and ( n70392 , n70388 , n70391 );
and ( n70393 , n70386 , n70391 );
or ( n70394 , n70389 , n70392 , n70393 );
and ( n70395 , n70148 , n70394 );
xor ( n70396 , n70148 , n70394 );
xor ( n70397 , n70386 , n70388 );
xor ( n70398 , n70397 , n70391 );
and ( n70399 , n65265 , n67498 );
and ( n70400 , n65175 , n67495 );
nor ( n70401 , n70399 , n70400 );
xnor ( n70402 , n70401 , n66511 );
xor ( n70403 , n70364 , n70366 );
xor ( n70404 , n70403 , n70369 );
and ( n70405 , n70402 , n70404 );
xor ( n70406 , n70106 , n70110 );
xor ( n70407 , n70406 , n70113 );
and ( n70408 , n70404 , n70407 );
and ( n70409 , n70402 , n70407 );
or ( n70410 , n70405 , n70408 , n70409 );
xor ( n70411 , n69964 , n69968 );
xor ( n70412 , n70411 , n69971 );
and ( n70413 , n70410 , n70412 );
xor ( n70414 , n70082 , n70116 );
xor ( n70415 , n70414 , n70119 );
and ( n70416 , n70412 , n70415 );
and ( n70417 , n70410 , n70415 );
or ( n70418 , n70413 , n70416 , n70417 );
xor ( n70419 , n70378 , n70380 );
xor ( n70420 , n70419 , n70383 );
and ( n70421 , n70418 , n70420 );
xor ( n70422 , n69974 , n70122 );
xor ( n70423 , n70422 , n70125 );
and ( n70424 , n70420 , n70423 );
and ( n70425 , n70418 , n70423 );
or ( n70426 , n70421 , n70424 , n70425 );
and ( n70427 , n70398 , n70426 );
xor ( n70428 , n70398 , n70426 );
and ( n70429 , n68625 , n64897 );
and ( n70430 , n68444 , n64895 );
nor ( n70431 , n70429 , n70430 );
xnor ( n70432 , n70431 , n64850 );
and ( n70433 , n68873 , n64789 );
and ( n70434 , n68837 , n64787 );
nor ( n70435 , n70433 , n70434 );
xnor ( n70436 , n70435 , n64738 );
and ( n70437 , n70432 , n70436 );
and ( n70438 , n69449 , n64711 );
and ( n70439 , n69095 , n64709 );
nor ( n70440 , n70438 , n70439 );
xnor ( n70441 , n70440 , n64682 );
and ( n70442 , n70436 , n70441 );
and ( n70443 , n70432 , n70441 );
or ( n70444 , n70437 , n70442 , n70443 );
and ( n70445 , n68199 , n65056 );
and ( n70446 , n68192 , n65054 );
nor ( n70447 , n70445 , n70446 );
xnor ( n70448 , n70447 , n64943 );
and ( n70449 , n70444 , n70448 );
xor ( n70450 , n70014 , n70018 );
xor ( n70451 , n70450 , n70021 );
and ( n70452 , n70448 , n70451 );
and ( n70453 , n70444 , n70451 );
or ( n70454 , n70449 , n70452 , n70453 );
and ( n70455 , n67833 , n65183 );
and ( n70456 , n67727 , n65181 );
nor ( n70457 , n70455 , n70456 );
xnor ( n70458 , n70457 , n64994 );
and ( n70459 , n70454 , n70458 );
xor ( n70460 , n70024 , n70028 );
xor ( n70461 , n70460 , n70031 );
and ( n70462 , n70458 , n70461 );
and ( n70463 , n70454 , n70461 );
or ( n70464 , n70459 , n70462 , n70463 );
and ( n70465 , n67307 , n65371 );
and ( n70466 , n67302 , n65369 );
nor ( n70467 , n70465 , n70466 );
xnor ( n70468 , n70467 , n65168 );
and ( n70469 , n70464 , n70468 );
xor ( n70470 , n70161 , n70165 );
xor ( n70471 , n70470 , n70168 );
and ( n70472 , n70468 , n70471 );
and ( n70473 , n70464 , n70471 );
or ( n70474 , n70469 , n70472 , n70473 );
and ( n70475 , n66517 , n66016 );
and ( n70476 , n66266 , n66014 );
nor ( n70477 , n70475 , n70476 );
xnor ( n70478 , n70477 , n65650 );
and ( n70479 , n70474 , n70478 );
xor ( n70480 , n70324 , n70326 );
xor ( n70481 , n70480 , n70329 );
and ( n70482 , n70478 , n70481 );
and ( n70483 , n70474 , n70481 );
or ( n70484 , n70479 , n70482 , n70483 );
and ( n70485 , n65698 , n66906 );
and ( n70486 , n65657 , n66904 );
nor ( n70487 , n70485 , n70486 );
xnor ( n70488 , n70487 , n66286 );
and ( n70489 , n70484 , n70488 );
xor ( n70490 , n70086 , n70090 );
xor ( n70491 , n70490 , n70093 );
and ( n70492 , n70488 , n70491 );
and ( n70493 , n70484 , n70491 );
or ( n70494 , n70489 , n70492 , n70493 );
and ( n70495 , n65363 , n67498 );
and ( n70496 , n65265 , n67495 );
nor ( n70497 , n70495 , n70496 );
xnor ( n70498 , n70497 , n66511 );
and ( n70499 , n70494 , n70498 );
xor ( n70500 , n70096 , n70100 );
xor ( n70501 , n70500 , n70103 );
and ( n70502 , n70498 , n70501 );
and ( n70503 , n70494 , n70501 );
or ( n70504 , n70499 , n70502 , n70503 );
and ( n70505 , n69095 , n64789 );
and ( n70506 , n68873 , n64787 );
nor ( n70507 , n70505 , n70506 );
xnor ( n70508 , n70507 , n64738 );
and ( n70509 , n69568 , n64711 );
and ( n70510 , n69449 , n64709 );
nor ( n70511 , n70509 , n70510 );
xnor ( n70512 , n70511 , n64682 );
and ( n70513 , n70508 , n70512 );
xor ( n70514 , n70256 , n70280 );
xor ( n70515 , n70514 , n70283 );
and ( n70516 , n70512 , n70515 );
and ( n70517 , n70508 , n70515 );
or ( n70518 , n70513 , n70516 , n70517 );
and ( n70519 , n68439 , n65056 );
and ( n70520 , n68199 , n65054 );
nor ( n70521 , n70519 , n70520 );
xnor ( n70522 , n70521 , n64943 );
and ( n70523 , n70518 , n70522 );
xor ( n70524 , n70242 , n70286 );
xor ( n70525 , n70524 , n70289 );
and ( n70526 , n70522 , n70525 );
and ( n70527 , n70518 , n70525 );
or ( n70528 , n70523 , n70526 , n70527 );
and ( n70529 , n67873 , n65183 );
and ( n70530 , n67833 , n65181 );
nor ( n70531 , n70529 , n70530 );
xnor ( n70532 , n70531 , n64994 );
and ( n70533 , n70528 , n70532 );
xor ( n70534 , n70292 , n70296 );
xor ( n70535 , n70534 , n70301 );
and ( n70536 , n70532 , n70535 );
and ( n70537 , n70528 , n70535 );
or ( n70538 , n70533 , n70536 , n70537 );
and ( n70539 , n67302 , n65550 );
and ( n70540 , n67111 , n65548 );
nor ( n70541 , n70539 , n70540 );
xnor ( n70542 , n70541 , n65313 );
and ( n70543 , n70538 , n70542 );
and ( n70544 , n67548 , n65371 );
and ( n70545 , n67307 , n65369 );
nor ( n70546 , n70544 , n70545 );
xnor ( n70547 , n70546 , n65168 );
and ( n70548 , n70542 , n70547 );
and ( n70549 , n70538 , n70547 );
or ( n70550 , n70543 , n70548 , n70549 );
and ( n70551 , n67111 , n65550 );
and ( n70552 , n66981 , n65548 );
nor ( n70553 , n70551 , n70552 );
xnor ( n70554 , n70553 , n65313 );
and ( n70555 , n70550 , n70554 );
xor ( n70556 , n70314 , n70318 );
xor ( n70557 , n70556 , n70321 );
and ( n70558 , n70554 , n70557 );
and ( n70559 , n70550 , n70557 );
or ( n70560 , n70555 , n70558 , n70559 );
and ( n70561 , n65883 , n66906 );
and ( n70562 , n65698 , n66904 );
nor ( n70563 , n70561 , n70562 );
xnor ( n70564 , n70563 , n66286 );
and ( n70565 , n70560 , n70564 );
and ( n70566 , n66276 , n66241 );
and ( n70567 , n66142 , n66239 );
nor ( n70568 , n70566 , n70567 );
xnor ( n70569 , n70568 , n65876 );
and ( n70570 , n70564 , n70569 );
and ( n70571 , n70560 , n70569 );
or ( n70572 , n70565 , n70570 , n70571 );
and ( n70573 , n65443 , n67160 );
and ( n70574 , n65453 , n67158 );
nor ( n70575 , n70573 , n70574 );
xnor ( n70576 , n70575 , n66514 );
and ( n70577 , n70572 , n70576 );
xor ( n70578 , n70332 , n70336 );
xor ( n70579 , n70578 , n70339 );
and ( n70580 , n70576 , n70579 );
and ( n70581 , n70572 , n70579 );
or ( n70582 , n70577 , n70580 , n70581 );
xor ( n70583 , n70196 , n70200 );
xor ( n70584 , n70583 , n70225 );
and ( n70585 , n70582 , n70584 );
xor ( n70586 , n70342 , n70346 );
xor ( n70587 , n70586 , n70349 );
and ( n70588 , n70584 , n70587 );
and ( n70589 , n70582 , n70587 );
or ( n70590 , n70585 , n70588 , n70589 );
and ( n70591 , n70504 , n70590 );
xor ( n70592 , n70228 , n70352 );
xor ( n70593 , n70592 , n70357 );
and ( n70594 , n70590 , n70593 );
and ( n70595 , n70504 , n70593 );
or ( n70596 , n70591 , n70594 , n70595 );
xor ( n70597 , n70360 , n70372 );
xor ( n70598 , n70597 , n70375 );
and ( n70599 , n70596 , n70598 );
xor ( n70600 , n70410 , n70412 );
xor ( n70601 , n70600 , n70415 );
and ( n70602 , n70598 , n70601 );
and ( n70603 , n70596 , n70601 );
or ( n70604 , n70599 , n70602 , n70603 );
xor ( n70605 , n70418 , n70420 );
xor ( n70606 , n70605 , n70423 );
and ( n70607 , n70604 , n70606 );
xor ( n70608 , n70604 , n70606 );
xor ( n70609 , n70596 , n70598 );
xor ( n70610 , n70609 , n70601 );
and ( n70611 , n66266 , n66241 );
and ( n70612 , n66276 , n66239 );
nor ( n70613 , n70611 , n70612 );
xnor ( n70614 , n70613 , n65876 );
and ( n70615 , n66507 , n66016 );
and ( n70616 , n66517 , n66014 );
nor ( n70617 , n70615 , n70616 );
xnor ( n70618 , n70617 , n65650 );
and ( n70619 , n70614 , n70618 );
xor ( n70620 , n70550 , n70554 );
xor ( n70621 , n70620 , n70557 );
and ( n70622 , n70618 , n70621 );
and ( n70623 , n70614 , n70621 );
or ( n70624 , n70619 , n70622 , n70623 );
and ( n70625 , n65453 , n67498 );
and ( n70626 , n65306 , n67495 );
nor ( n70627 , n70625 , n70626 );
xnor ( n70628 , n70627 , n66511 );
and ( n70629 , n70624 , n70628 );
and ( n70630 , n65657 , n67160 );
and ( n70631 , n65443 , n67158 );
nor ( n70632 , n70630 , n70631 );
xnor ( n70633 , n70632 , n66514 );
and ( n70634 , n70628 , n70633 );
and ( n70635 , n70624 , n70633 );
or ( n70636 , n70629 , n70634 , n70635 );
and ( n70637 , n67833 , n65371 );
and ( n70638 , n67727 , n65369 );
nor ( n70639 , n70637 , n70638 );
xnor ( n70640 , n70639 , n65168 );
and ( n70641 , n68192 , n65183 );
and ( n70642 , n67873 , n65181 );
nor ( n70643 , n70641 , n70642 );
xnor ( n70644 , n70643 , n64994 );
and ( n70645 , n70640 , n70644 );
xor ( n70646 , n70432 , n70436 );
xor ( n70647 , n70646 , n70441 );
and ( n70648 , n70644 , n70647 );
and ( n70649 , n70640 , n70647 );
or ( n70650 , n70645 , n70648 , n70649 );
and ( n70651 , n67727 , n65371 );
and ( n70652 , n67548 , n65369 );
nor ( n70653 , n70651 , n70652 );
xnor ( n70654 , n70653 , n65168 );
and ( n70655 , n70650 , n70654 );
xor ( n70656 , n70444 , n70448 );
xor ( n70657 , n70656 , n70451 );
and ( n70658 , n70654 , n70657 );
and ( n70659 , n70650 , n70657 );
or ( n70660 , n70655 , n70658 , n70659 );
xor ( n70661 , n70304 , n70308 );
xor ( n70662 , n70661 , n70311 );
and ( n70663 , n70660 , n70662 );
xor ( n70664 , n70454 , n70458 );
xor ( n70665 , n70664 , n70461 );
and ( n70666 , n70662 , n70665 );
and ( n70667 , n70660 , n70665 );
or ( n70668 , n70663 , n70666 , n70667 );
and ( n70669 , n66786 , n65756 );
and ( n70670 , n66781 , n65754 );
nor ( n70671 , n70669 , n70670 );
xnor ( n70672 , n70671 , n65450 );
and ( n70673 , n70668 , n70672 );
xor ( n70674 , n70464 , n70468 );
xor ( n70675 , n70674 , n70471 );
and ( n70676 , n70672 , n70675 );
and ( n70677 , n70668 , n70675 );
or ( n70678 , n70673 , n70676 , n70677 );
and ( n70679 , n66137 , n66657 );
and ( n70680 , n65935 , n66655 );
nor ( n70681 , n70679 , n70680 );
xnor ( n70682 , n70681 , n66130 );
and ( n70683 , n70678 , n70682 );
xor ( n70684 , n70152 , n70156 );
xor ( n70685 , n70684 , n70181 );
and ( n70686 , n70682 , n70685 );
and ( n70687 , n70678 , n70685 );
or ( n70688 , n70683 , n70686 , n70687 );
and ( n70689 , n70636 , n70688 );
xor ( n70690 , n70184 , n70188 );
xor ( n70691 , n70690 , n70193 );
and ( n70692 , n70688 , n70691 );
and ( n70693 , n70636 , n70691 );
or ( n70694 , n70689 , n70692 , n70693 );
and ( n70695 , n66781 , n66016 );
and ( n70696 , n66507 , n66014 );
nor ( n70697 , n70695 , n70696 );
xnor ( n70698 , n70697 , n65650 );
and ( n70699 , n66981 , n65756 );
and ( n70700 , n66786 , n65754 );
nor ( n70701 , n70699 , n70700 );
xnor ( n70702 , n70701 , n65450 );
and ( n70703 , n70698 , n70702 );
xor ( n70704 , n70538 , n70542 );
xor ( n70705 , n70704 , n70547 );
and ( n70706 , n70702 , n70705 );
and ( n70707 , n70698 , n70705 );
or ( n70708 , n70703 , n70706 , n70707 );
and ( n70709 , n65935 , n66906 );
and ( n70710 , n65883 , n66904 );
nor ( n70711 , n70709 , n70710 );
xnor ( n70712 , n70711 , n66286 );
and ( n70713 , n70708 , n70712 );
and ( n70714 , n66142 , n66657 );
and ( n70715 , n66137 , n66655 );
nor ( n70716 , n70714 , n70715 );
xnor ( n70717 , n70716 , n66130 );
and ( n70718 , n70712 , n70717 );
and ( n70719 , n70708 , n70717 );
or ( n70720 , n70713 , n70718 , n70719 );
xor ( n70721 , n70560 , n70564 );
xor ( n70722 , n70721 , n70569 );
and ( n70723 , n70720 , n70722 );
xor ( n70724 , n70474 , n70478 );
xor ( n70725 , n70724 , n70481 );
and ( n70726 , n70722 , n70725 );
and ( n70727 , n70720 , n70725 );
or ( n70728 , n70723 , n70726 , n70727 );
and ( n70729 , n65306 , n67498 );
and ( n70730 , n65363 , n67495 );
nor ( n70731 , n70729 , n70730 );
xnor ( n70732 , n70731 , n66511 );
and ( n70733 , n70728 , n70732 );
xor ( n70734 , n70484 , n70488 );
xor ( n70735 , n70734 , n70491 );
and ( n70736 , n70732 , n70735 );
and ( n70737 , n70728 , n70735 );
or ( n70738 , n70733 , n70736 , n70737 );
and ( n70739 , n70694 , n70738 );
xor ( n70740 , n70494 , n70498 );
xor ( n70741 , n70740 , n70501 );
and ( n70742 , n70738 , n70741 );
and ( n70743 , n70694 , n70741 );
or ( n70744 , n70739 , n70742 , n70743 );
xor ( n70745 , n70504 , n70590 );
xor ( n70746 , n70745 , n70593 );
and ( n70747 , n70744 , n70746 );
xor ( n70748 , n70402 , n70404 );
xor ( n70749 , n70748 , n70407 );
and ( n70750 , n70746 , n70749 );
and ( n70751 , n70744 , n70749 );
or ( n70752 , n70747 , n70750 , n70751 );
and ( n70753 , n70610 , n70752 );
xor ( n70754 , n70610 , n70752 );
xor ( n70755 , n70744 , n70746 );
xor ( n70756 , n70755 , n70749 );
and ( n70757 , n70238 , n64652 );
and ( n70758 , n69985 , n64650 );
nor ( n70759 , n70757 , n70758 );
xnor ( n70760 , n70759 , n64609 );
and ( n70761 , n70266 , n64617 );
and ( n70762 , n70252 , n64615 );
nor ( n70763 , n70761 , n70762 );
xnor ( n70764 , n70763 , n64624 );
and ( n70765 , n70760 , n70764 );
buf ( n70766 , n64564 );
and ( n70767 , n70766 , n64612 );
and ( n70768 , n70764 , n70767 );
and ( n70769 , n70760 , n70767 );
or ( n70770 , n70765 , n70768 , n70769 );
and ( n70771 , n69573 , n64711 );
and ( n70772 , n69566 , n64709 );
nor ( n70773 , n70771 , n70772 );
xnor ( n70774 , n70773 , n64682 );
and ( n70775 , n70770 , n70774 );
xor ( n70776 , n70260 , n70264 );
xor ( n70777 , n70776 , n70267 );
and ( n70778 , n70774 , n70777 );
and ( n70779 , n70770 , n70777 );
or ( n70780 , n70775 , n70778 , n70779 );
buf ( n70781 , n64571 );
and ( n70782 , n70781 , n64615 );
not ( n70783 , n70782 );
and ( n70784 , n70783 , n64624 );
and ( n70785 , n70781 , n64617 );
buf ( n70786 , n64570 );
and ( n70787 , n70786 , n64615 );
nor ( n70788 , n70785 , n70787 );
xnor ( n70789 , n70788 , n64624 );
and ( n70790 , n70784 , n70789 );
and ( n70791 , n70786 , n64617 );
buf ( n70792 , n64569 );
and ( n70793 , n70792 , n64615 );
nor ( n70794 , n70791 , n70793 );
xnor ( n70795 , n70794 , n64624 );
and ( n70796 , n70790 , n70795 );
and ( n70797 , n70781 , n64612 );
and ( n70798 , n70795 , n70797 );
and ( n70799 , n70790 , n70797 );
or ( n70800 , n70796 , n70798 , n70799 );
and ( n70801 , n70792 , n64617 );
buf ( n70802 , n64568 );
and ( n70803 , n70802 , n64615 );
nor ( n70804 , n70801 , n70803 );
xnor ( n70805 , n70804 , n64624 );
and ( n70806 , n70800 , n70805 );
and ( n70807 , n70786 , n64612 );
and ( n70808 , n70805 , n70807 );
and ( n70809 , n70800 , n70807 );
or ( n70810 , n70806 , n70808 , n70809 );
and ( n70811 , n70802 , n64617 );
buf ( n70812 , n64567 );
and ( n70813 , n70812 , n64615 );
nor ( n70814 , n70811 , n70813 );
xnor ( n70815 , n70814 , n64624 );
and ( n70816 , n70810 , n70815 );
and ( n70817 , n70792 , n64612 );
and ( n70818 , n70815 , n70817 );
and ( n70819 , n70810 , n70817 );
or ( n70820 , n70816 , n70818 , n70819 );
and ( n70821 , n70812 , n64617 );
buf ( n70822 , n64566 );
and ( n70823 , n70822 , n64615 );
nor ( n70824 , n70821 , n70823 );
xnor ( n70825 , n70824 , n64624 );
and ( n70826 , n70820 , n70825 );
and ( n70827 , n70802 , n64612 );
and ( n70828 , n70825 , n70827 );
and ( n70829 , n70820 , n70827 );
or ( n70830 , n70826 , n70828 , n70829 );
and ( n70831 , n70822 , n64617 );
buf ( n70832 , n64565 );
and ( n70833 , n70832 , n64615 );
nor ( n70834 , n70831 , n70833 );
xnor ( n70835 , n70834 , n64624 );
and ( n70836 , n70830 , n70835 );
and ( n70837 , n70812 , n64612 );
and ( n70838 , n70835 , n70837 );
and ( n70839 , n70830 , n70837 );
or ( n70840 , n70836 , n70838 , n70839 );
and ( n70841 , n70832 , n64617 );
and ( n70842 , n70766 , n64615 );
nor ( n70843 , n70841 , n70842 );
xnor ( n70844 , n70843 , n64624 );
and ( n70845 , n70840 , n70844 );
and ( n70846 , n70822 , n64612 );
and ( n70847 , n70844 , n70846 );
and ( n70848 , n70840 , n70846 );
or ( n70849 , n70845 , n70847 , n70848 );
and ( n70850 , n70766 , n64617 );
and ( n70851 , n70266 , n64615 );
nor ( n70852 , n70850 , n70851 );
xnor ( n70853 , n70852 , n64624 );
and ( n70854 , n70849 , n70853 );
and ( n70855 , n70832 , n64612 );
and ( n70856 , n70853 , n70855 );
and ( n70857 , n70849 , n70855 );
or ( n70858 , n70854 , n70856 , n70857 );
and ( n70859 , n69979 , n64711 );
and ( n70860 , n69573 , n64709 );
nor ( n70861 , n70859 , n70860 );
xnor ( n70862 , n70861 , n64682 );
and ( n70863 , n70858 , n70862 );
xor ( n70864 , n70760 , n70764 );
xor ( n70865 , n70864 , n70767 );
and ( n70866 , n70862 , n70865 );
and ( n70867 , n70858 , n70865 );
or ( n70868 , n70863 , n70866 , n70867 );
and ( n70869 , n70238 , n64711 );
and ( n70870 , n69985 , n64709 );
nor ( n70871 , n70869 , n70870 );
xnor ( n70872 , n70871 , n64682 );
and ( n70873 , n70266 , n64652 );
and ( n70874 , n70252 , n64650 );
nor ( n70875 , n70873 , n70874 );
xnor ( n70876 , n70875 , n64609 );
and ( n70877 , n70872 , n70876 );
xor ( n70878 , n70840 , n70844 );
xor ( n70879 , n70878 , n70846 );
and ( n70880 , n70876 , n70879 );
and ( n70881 , n70872 , n70879 );
or ( n70882 , n70877 , n70880 , n70881 );
and ( n70883 , n70252 , n64652 );
and ( n70884 , n70238 , n64650 );
nor ( n70885 , n70883 , n70884 );
xnor ( n70886 , n70885 , n64609 );
and ( n70887 , n70882 , n70886 );
xor ( n70888 , n70849 , n70853 );
xor ( n70889 , n70888 , n70855 );
and ( n70890 , n70886 , n70889 );
and ( n70891 , n70882 , n70889 );
or ( n70892 , n70887 , n70890 , n70891 );
and ( n70893 , n69566 , n64789 );
and ( n70894 , n69568 , n64787 );
nor ( n70895 , n70893 , n70894 );
xnor ( n70896 , n70895 , n64738 );
and ( n70897 , n70892 , n70896 );
xor ( n70898 , n70858 , n70862 );
xor ( n70899 , n70898 , n70865 );
and ( n70900 , n70896 , n70899 );
and ( n70901 , n70892 , n70899 );
or ( n70902 , n70897 , n70900 , n70901 );
and ( n70903 , n70868 , n70902 );
xor ( n70904 , n70770 , n70774 );
xor ( n70905 , n70904 , n70777 );
and ( n70906 , n70902 , n70905 );
and ( n70907 , n70868 , n70905 );
or ( n70908 , n70903 , n70906 , n70907 );
and ( n70909 , n70780 , n70908 );
xor ( n70910 , n70270 , n70274 );
xor ( n70911 , n70910 , n70277 );
and ( n70912 , n70908 , n70911 );
and ( n70913 , n70780 , n70911 );
or ( n70914 , n70909 , n70912 , n70913 );
and ( n70915 , n68444 , n65056 );
and ( n70916 , n68439 , n65054 );
nor ( n70917 , n70915 , n70916 );
xnor ( n70918 , n70917 , n64943 );
and ( n70919 , n70914 , n70918 );
and ( n70920 , n68837 , n64897 );
and ( n70921 , n68625 , n64895 );
nor ( n70922 , n70920 , n70921 );
xnor ( n70923 , n70922 , n64850 );
and ( n70924 , n70918 , n70923 );
and ( n70925 , n70914 , n70923 );
or ( n70926 , n70919 , n70924 , n70925 );
and ( n70927 , n68625 , n65056 );
and ( n70928 , n68444 , n65054 );
nor ( n70929 , n70927 , n70928 );
xnor ( n70930 , n70929 , n64943 );
and ( n70931 , n68873 , n64897 );
and ( n70932 , n68837 , n64895 );
nor ( n70933 , n70931 , n70932 );
xnor ( n70934 , n70933 , n64850 );
and ( n70935 , n70930 , n70934 );
and ( n70936 , n69449 , n64789 );
and ( n70937 , n69095 , n64787 );
nor ( n70938 , n70936 , n70937 );
xnor ( n70939 , n70938 , n64738 );
and ( n70940 , n70934 , n70939 );
and ( n70941 , n70930 , n70939 );
or ( n70942 , n70935 , n70940 , n70941 );
and ( n70943 , n67873 , n65371 );
and ( n70944 , n67833 , n65369 );
nor ( n70945 , n70943 , n70944 );
xnor ( n70946 , n70945 , n65168 );
and ( n70947 , n70942 , n70946 );
xor ( n70948 , n70508 , n70512 );
xor ( n70949 , n70948 , n70515 );
and ( n70950 , n70946 , n70949 );
and ( n70951 , n70942 , n70949 );
or ( n70952 , n70947 , n70950 , n70951 );
and ( n70953 , n70926 , n70952 );
xor ( n70954 , n70518 , n70522 );
xor ( n70955 , n70954 , n70525 );
and ( n70956 , n70952 , n70955 );
and ( n70957 , n70926 , n70955 );
or ( n70958 , n70953 , n70956 , n70957 );
and ( n70959 , n67307 , n65550 );
and ( n70960 , n67302 , n65548 );
nor ( n70961 , n70959 , n70960 );
xnor ( n70962 , n70961 , n65313 );
and ( n70963 , n70958 , n70962 );
xor ( n70964 , n70528 , n70532 );
xor ( n70965 , n70964 , n70535 );
and ( n70966 , n70962 , n70965 );
and ( n70967 , n70958 , n70965 );
or ( n70968 , n70963 , n70966 , n70967 );
and ( n70969 , n66517 , n66241 );
and ( n70970 , n66266 , n66239 );
nor ( n70971 , n70969 , n70970 );
xnor ( n70972 , n70971 , n65876 );
and ( n70973 , n70968 , n70972 );
xor ( n70974 , n70660 , n70662 );
xor ( n70975 , n70974 , n70665 );
and ( n70976 , n70972 , n70975 );
and ( n70977 , n70968 , n70975 );
or ( n70978 , n70973 , n70976 , n70977 );
and ( n70979 , n65698 , n67160 );
and ( n70980 , n65657 , n67158 );
nor ( n70981 , n70979 , n70980 );
xnor ( n70982 , n70981 , n66514 );
and ( n70983 , n70978 , n70982 );
xor ( n70984 , n70668 , n70672 );
xor ( n70985 , n70984 , n70675 );
and ( n70986 , n70982 , n70985 );
and ( n70987 , n70978 , n70985 );
or ( n70988 , n70983 , n70986 , n70987 );
and ( n70989 , n67302 , n65756 );
and ( n70990 , n67111 , n65754 );
nor ( n70991 , n70989 , n70990 );
xnor ( n70992 , n70991 , n65450 );
and ( n70993 , n67548 , n65550 );
and ( n70994 , n67307 , n65548 );
nor ( n70995 , n70993 , n70994 );
xnor ( n70996 , n70995 , n65313 );
and ( n70997 , n70992 , n70996 );
xor ( n70998 , n70640 , n70644 );
xor ( n70999 , n70998 , n70647 );
and ( n71000 , n70996 , n70999 );
and ( n71001 , n70992 , n70999 );
or ( n71002 , n70997 , n71000 , n71001 );
and ( n71003 , n67111 , n65756 );
and ( n71004 , n66981 , n65754 );
nor ( n71005 , n71003 , n71004 );
xnor ( n71006 , n71005 , n65450 );
and ( n71007 , n71002 , n71006 );
xor ( n71008 , n70650 , n70654 );
xor ( n71009 , n71008 , n70657 );
and ( n71010 , n71006 , n71009 );
and ( n71011 , n71002 , n71009 );
or ( n71012 , n71007 , n71010 , n71011 );
and ( n71013 , n66276 , n66657 );
and ( n71014 , n66142 , n66655 );
nor ( n71015 , n71013 , n71014 );
xnor ( n71016 , n71015 , n66130 );
and ( n71017 , n71012 , n71016 );
xor ( n71018 , n70698 , n70702 );
xor ( n71019 , n71018 , n70705 );
and ( n71020 , n71016 , n71019 );
and ( n71021 , n71012 , n71019 );
or ( n71022 , n71017 , n71020 , n71021 );
and ( n71023 , n65443 , n67498 );
and ( n71024 , n65453 , n67495 );
nor ( n71025 , n71023 , n71024 );
xnor ( n71026 , n71025 , n66511 );
and ( n71027 , n71022 , n71026 );
xor ( n71028 , n70614 , n70618 );
xor ( n71029 , n71028 , n70621 );
and ( n71030 , n71026 , n71029 );
and ( n71031 , n71022 , n71029 );
or ( n71032 , n71027 , n71030 , n71031 );
and ( n71033 , n70988 , n71032 );
xor ( n71034 , n70678 , n70682 );
xor ( n71035 , n71034 , n70685 );
and ( n71036 , n71032 , n71035 );
and ( n71037 , n70988 , n71035 );
or ( n71038 , n71033 , n71036 , n71037 );
xor ( n71039 , n70636 , n70688 );
xor ( n71040 , n71039 , n70691 );
and ( n71041 , n71038 , n71040 );
xor ( n71042 , n70572 , n70576 );
xor ( n71043 , n71042 , n70579 );
and ( n71044 , n71040 , n71043 );
and ( n71045 , n71038 , n71043 );
or ( n71046 , n71041 , n71044 , n71045 );
xor ( n71047 , n70694 , n70738 );
xor ( n71048 , n71047 , n70741 );
and ( n71049 , n71046 , n71048 );
xor ( n71050 , n70582 , n70584 );
xor ( n71051 , n71050 , n70587 );
and ( n71052 , n71048 , n71051 );
and ( n71053 , n71046 , n71051 );
or ( n71054 , n71049 , n71052 , n71053 );
and ( n71055 , n70756 , n71054 );
xor ( n71056 , n70756 , n71054 );
xor ( n71057 , n71046 , n71048 );
xor ( n71058 , n71057 , n71051 );
and ( n71059 , n69095 , n64897 );
and ( n71060 , n68873 , n64895 );
nor ( n71061 , n71059 , n71060 );
xnor ( n71062 , n71061 , n64850 );
and ( n71063 , n69568 , n64789 );
and ( n71064 , n69449 , n64787 );
nor ( n71065 , n71063 , n71064 );
xnor ( n71066 , n71065 , n64738 );
and ( n71067 , n71062 , n71066 );
xor ( n71068 , n70868 , n70902 );
xor ( n71069 , n71068 , n70905 );
and ( n71070 , n71066 , n71069 );
and ( n71071 , n71062 , n71069 );
or ( n71072 , n71067 , n71070 , n71071 );
and ( n71073 , n68439 , n65183 );
and ( n71074 , n68199 , n65181 );
nor ( n71075 , n71073 , n71074 );
xnor ( n71076 , n71075 , n64994 );
and ( n71077 , n71072 , n71076 );
xor ( n71078 , n70780 , n70908 );
xor ( n71079 , n71078 , n70911 );
and ( n71080 , n71076 , n71079 );
and ( n71081 , n71072 , n71079 );
or ( n71082 , n71077 , n71080 , n71081 );
and ( n71083 , n68199 , n65183 );
and ( n71084 , n68192 , n65181 );
nor ( n71085 , n71083 , n71084 );
xnor ( n71086 , n71085 , n64994 );
and ( n71087 , n71082 , n71086 );
xor ( n71088 , n70914 , n70918 );
xor ( n71089 , n71088 , n70923 );
and ( n71090 , n71086 , n71089 );
and ( n71091 , n71082 , n71089 );
or ( n71092 , n71087 , n71090 , n71091 );
and ( n71093 , n69573 , n64789 );
and ( n71094 , n69566 , n64787 );
nor ( n71095 , n71093 , n71094 );
xnor ( n71096 , n71095 , n64738 );
and ( n71097 , n69985 , n64711 );
and ( n71098 , n69979 , n64709 );
nor ( n71099 , n71097 , n71098 );
xnor ( n71100 , n71099 , n64682 );
and ( n71101 , n71096 , n71100 );
xor ( n71102 , n70882 , n70886 );
xor ( n71103 , n71102 , n70889 );
and ( n71104 , n71100 , n71103 );
and ( n71105 , n71096 , n71103 );
or ( n71106 , n71101 , n71104 , n71105 );
xor ( n71107 , n70784 , n70789 );
and ( n71108 , n70781 , n64650 );
not ( n71109 , n71108 );
and ( n71110 , n71109 , n64609 );
and ( n71111 , n70781 , n64652 );
and ( n71112 , n70786 , n64650 );
nor ( n71113 , n71111 , n71112 );
xnor ( n71114 , n71113 , n64609 );
and ( n71115 , n71110 , n71114 );
and ( n71116 , n70786 , n64652 );
and ( n71117 , n70792 , n64650 );
nor ( n71118 , n71116 , n71117 );
xnor ( n71119 , n71118 , n64609 );
and ( n71120 , n71115 , n71119 );
and ( n71121 , n71119 , n70782 );
and ( n71122 , n71115 , n70782 );
or ( n71123 , n71120 , n71121 , n71122 );
and ( n71124 , n71107 , n71123 );
and ( n71125 , n70792 , n64652 );
and ( n71126 , n70802 , n64650 );
nor ( n71127 , n71125 , n71126 );
xnor ( n71128 , n71127 , n64609 );
and ( n71129 , n71123 , n71128 );
and ( n71130 , n71107 , n71128 );
or ( n71131 , n71124 , n71129 , n71130 );
and ( n71132 , n70802 , n64652 );
and ( n71133 , n70812 , n64650 );
nor ( n71134 , n71132 , n71133 );
xnor ( n71135 , n71134 , n64609 );
and ( n71136 , n71131 , n71135 );
xor ( n71137 , n70790 , n70795 );
xor ( n71138 , n71137 , n70797 );
and ( n71139 , n71135 , n71138 );
and ( n71140 , n71131 , n71138 );
or ( n71141 , n71136 , n71139 , n71140 );
and ( n71142 , n70812 , n64652 );
and ( n71143 , n70822 , n64650 );
nor ( n71144 , n71142 , n71143 );
xnor ( n71145 , n71144 , n64609 );
and ( n71146 , n71141 , n71145 );
xor ( n71147 , n70800 , n70805 );
xor ( n71148 , n71147 , n70807 );
and ( n71149 , n71145 , n71148 );
and ( n71150 , n71141 , n71148 );
or ( n71151 , n71146 , n71149 , n71150 );
and ( n71152 , n70822 , n64652 );
and ( n71153 , n70832 , n64650 );
nor ( n71154 , n71152 , n71153 );
xnor ( n71155 , n71154 , n64609 );
and ( n71156 , n71151 , n71155 );
xor ( n71157 , n70810 , n70815 );
xor ( n71158 , n71157 , n70817 );
and ( n71159 , n71155 , n71158 );
and ( n71160 , n71151 , n71158 );
or ( n71161 , n71156 , n71159 , n71160 );
and ( n71162 , n70832 , n64652 );
and ( n71163 , n70766 , n64650 );
nor ( n71164 , n71162 , n71163 );
xnor ( n71165 , n71164 , n64609 );
and ( n71166 , n71161 , n71165 );
xor ( n71167 , n70820 , n70825 );
xor ( n71168 , n71167 , n70827 );
and ( n71169 , n71165 , n71168 );
and ( n71170 , n71161 , n71168 );
or ( n71171 , n71166 , n71169 , n71170 );
and ( n71172 , n70766 , n64652 );
and ( n71173 , n70266 , n64650 );
nor ( n71174 , n71172 , n71173 );
xnor ( n71175 , n71174 , n64609 );
and ( n71176 , n71171 , n71175 );
xor ( n71177 , n70830 , n70835 );
xor ( n71178 , n71177 , n70837 );
and ( n71179 , n71175 , n71178 );
and ( n71180 , n71171 , n71178 );
or ( n71181 , n71176 , n71179 , n71180 );
and ( n71182 , n69979 , n64789 );
and ( n71183 , n69573 , n64787 );
nor ( n71184 , n71182 , n71183 );
xnor ( n71185 , n71184 , n64738 );
and ( n71186 , n71181 , n71185 );
xor ( n71187 , n70872 , n70876 );
xor ( n71188 , n71187 , n70879 );
and ( n71189 , n71185 , n71188 );
and ( n71190 , n71181 , n71188 );
or ( n71191 , n71186 , n71189 , n71190 );
and ( n71192 , n70238 , n64789 );
and ( n71193 , n69985 , n64787 );
nor ( n71194 , n71192 , n71193 );
xnor ( n71195 , n71194 , n64738 );
and ( n71196 , n70266 , n64711 );
and ( n71197 , n70252 , n64709 );
nor ( n71198 , n71196 , n71197 );
xnor ( n71199 , n71198 , n64682 );
and ( n71200 , n71195 , n71199 );
xor ( n71201 , n71161 , n71165 );
xor ( n71202 , n71201 , n71168 );
and ( n71203 , n71199 , n71202 );
and ( n71204 , n71195 , n71202 );
or ( n71205 , n71200 , n71203 , n71204 );
and ( n71206 , n70252 , n64711 );
and ( n71207 , n70238 , n64709 );
nor ( n71208 , n71206 , n71207 );
xnor ( n71209 , n71208 , n64682 );
and ( n71210 , n71205 , n71209 );
xor ( n71211 , n71171 , n71175 );
xor ( n71212 , n71211 , n71178 );
and ( n71213 , n71209 , n71212 );
and ( n71214 , n71205 , n71212 );
or ( n71215 , n71210 , n71213 , n71214 );
and ( n71216 , n69566 , n64897 );
and ( n71217 , n69568 , n64895 );
nor ( n71218 , n71216 , n71217 );
xnor ( n71219 , n71218 , n64850 );
and ( n71220 , n71215 , n71219 );
xor ( n71221 , n71181 , n71185 );
xor ( n71222 , n71221 , n71188 );
and ( n71223 , n71219 , n71222 );
and ( n71224 , n71215 , n71222 );
or ( n71225 , n71220 , n71223 , n71224 );
and ( n71226 , n71191 , n71225 );
xor ( n71227 , n71096 , n71100 );
xor ( n71228 , n71227 , n71103 );
and ( n71229 , n71225 , n71228 );
and ( n71230 , n71191 , n71228 );
or ( n71231 , n71226 , n71229 , n71230 );
and ( n71232 , n71106 , n71231 );
xor ( n71233 , n70892 , n70896 );
xor ( n71234 , n71233 , n70899 );
and ( n71235 , n71231 , n71234 );
and ( n71236 , n71106 , n71234 );
or ( n71237 , n71232 , n71235 , n71236 );
and ( n71238 , n68444 , n65183 );
and ( n71239 , n68439 , n65181 );
nor ( n71240 , n71238 , n71239 );
xnor ( n71241 , n71240 , n64994 );
and ( n71242 , n71237 , n71241 );
and ( n71243 , n68837 , n65056 );
and ( n71244 , n68625 , n65054 );
nor ( n71245 , n71243 , n71244 );
xnor ( n71246 , n71245 , n64943 );
and ( n71247 , n71241 , n71246 );
and ( n71248 , n71237 , n71246 );
or ( n71249 , n71242 , n71247 , n71248 );
and ( n71250 , n67833 , n65550 );
and ( n71251 , n67727 , n65548 );
nor ( n71252 , n71250 , n71251 );
xnor ( n71253 , n71252 , n65313 );
and ( n71254 , n71249 , n71253 );
xor ( n71255 , n70930 , n70934 );
xor ( n71256 , n71255 , n70939 );
and ( n71257 , n71253 , n71256 );
and ( n71258 , n71249 , n71256 );
or ( n71259 , n71254 , n71257 , n71258 );
and ( n71260 , n67727 , n65550 );
and ( n71261 , n67548 , n65548 );
nor ( n71262 , n71260 , n71261 );
xnor ( n71263 , n71262 , n65313 );
and ( n71264 , n71259 , n71263 );
xor ( n71265 , n70942 , n70946 );
xor ( n71266 , n71265 , n70949 );
and ( n71267 , n71263 , n71266 );
and ( n71268 , n71259 , n71266 );
or ( n71269 , n71264 , n71267 , n71268 );
and ( n71270 , n71092 , n71269 );
xor ( n71271 , n70926 , n70952 );
xor ( n71272 , n71271 , n70955 );
and ( n71273 , n71269 , n71272 );
and ( n71274 , n71092 , n71272 );
or ( n71275 , n71270 , n71273 , n71274 );
and ( n71276 , n66786 , n66016 );
and ( n71277 , n66781 , n66014 );
nor ( n71278 , n71276 , n71277 );
xnor ( n71279 , n71278 , n65650 );
and ( n71280 , n71275 , n71279 );
xor ( n71281 , n70958 , n70962 );
xor ( n71282 , n71281 , n70965 );
and ( n71283 , n71279 , n71282 );
and ( n71284 , n71275 , n71282 );
or ( n71285 , n71280 , n71283 , n71284 );
and ( n71286 , n65883 , n67160 );
and ( n71287 , n65698 , n67158 );
nor ( n71288 , n71286 , n71287 );
xnor ( n71289 , n71288 , n66514 );
and ( n71290 , n71285 , n71289 );
and ( n71291 , n66137 , n66906 );
and ( n71292 , n65935 , n66904 );
nor ( n71293 , n71291 , n71292 );
xnor ( n71294 , n71293 , n66286 );
and ( n71295 , n71289 , n71294 );
and ( n71296 , n71285 , n71294 );
or ( n71297 , n71290 , n71295 , n71296 );
and ( n71298 , n66266 , n66657 );
and ( n71299 , n66276 , n66655 );
nor ( n71300 , n71298 , n71299 );
xnor ( n71301 , n71300 , n66130 );
and ( n71302 , n66507 , n66241 );
and ( n71303 , n66517 , n66239 );
nor ( n71304 , n71302 , n71303 );
xnor ( n71305 , n71304 , n65876 );
and ( n71306 , n71301 , n71305 );
xor ( n71307 , n71002 , n71006 );
xor ( n71308 , n71307 , n71009 );
and ( n71309 , n71305 , n71308 );
and ( n71310 , n71301 , n71308 );
or ( n71311 , n71306 , n71309 , n71310 );
and ( n71312 , n65657 , n67498 );
and ( n71313 , n65443 , n67495 );
nor ( n71314 , n71312 , n71313 );
xnor ( n71315 , n71314 , n66511 );
and ( n71316 , n71311 , n71315 );
xor ( n71317 , n70968 , n70972 );
xor ( n71318 , n71317 , n70975 );
and ( n71319 , n71315 , n71318 );
and ( n71320 , n71311 , n71318 );
or ( n71321 , n71316 , n71319 , n71320 );
and ( n71322 , n71297 , n71321 );
xor ( n71323 , n70708 , n70712 );
xor ( n71324 , n71323 , n70717 );
and ( n71325 , n71321 , n71324 );
and ( n71326 , n71297 , n71324 );
or ( n71327 , n71322 , n71325 , n71326 );
xor ( n71328 , n70624 , n70628 );
xor ( n71329 , n71328 , n70633 );
and ( n71330 , n71327 , n71329 );
xor ( n71331 , n70720 , n70722 );
xor ( n71332 , n71331 , n70725 );
and ( n71333 , n71329 , n71332 );
and ( n71334 , n71327 , n71332 );
or ( n71335 , n71330 , n71333 , n71334 );
xor ( n71336 , n70728 , n70732 );
xor ( n71337 , n71336 , n70735 );
and ( n71338 , n71335 , n71337 );
xor ( n71339 , n71038 , n71040 );
xor ( n71340 , n71339 , n71043 );
and ( n71341 , n71337 , n71340 );
and ( n71342 , n71335 , n71340 );
or ( n71343 , n71338 , n71341 , n71342 );
and ( n71344 , n71058 , n71343 );
xor ( n71345 , n71058 , n71343 );
xor ( n71346 , n71335 , n71337 );
xor ( n71347 , n71346 , n71340 );
and ( n71348 , n66781 , n66241 );
and ( n71349 , n66507 , n66239 );
nor ( n71350 , n71348 , n71349 );
xnor ( n71351 , n71350 , n65876 );
and ( n71352 , n66981 , n66016 );
and ( n71353 , n66786 , n66014 );
nor ( n71354 , n71352 , n71353 );
xnor ( n71355 , n71354 , n65650 );
and ( n71356 , n71351 , n71355 );
xor ( n71357 , n70992 , n70996 );
xor ( n71358 , n71357 , n70999 );
and ( n71359 , n71355 , n71358 );
and ( n71360 , n71351 , n71358 );
or ( n71361 , n71356 , n71359 , n71360 );
and ( n71362 , n65935 , n67160 );
and ( n71363 , n65883 , n67158 );
nor ( n71364 , n71362 , n71363 );
xnor ( n71365 , n71364 , n66514 );
and ( n71366 , n71361 , n71365 );
and ( n71367 , n66142 , n66906 );
and ( n71368 , n66137 , n66904 );
nor ( n71369 , n71367 , n71368 );
xnor ( n71370 , n71369 , n66286 );
and ( n71371 , n71365 , n71370 );
and ( n71372 , n71361 , n71370 );
or ( n71373 , n71366 , n71371 , n71372 );
and ( n71374 , n68625 , n65183 );
and ( n71375 , n68444 , n65181 );
nor ( n71376 , n71374 , n71375 );
xnor ( n71377 , n71376 , n64994 );
and ( n71378 , n68873 , n65056 );
and ( n71379 , n68837 , n65054 );
nor ( n71380 , n71378 , n71379 );
xnor ( n71381 , n71380 , n64943 );
and ( n71382 , n71377 , n71381 );
and ( n71383 , n69449 , n64897 );
and ( n71384 , n69095 , n64895 );
nor ( n71385 , n71383 , n71384 );
xnor ( n71386 , n71385 , n64850 );
and ( n71387 , n71381 , n71386 );
and ( n71388 , n71377 , n71386 );
or ( n71389 , n71382 , n71387 , n71388 );
xor ( n71390 , n71237 , n71241 );
xor ( n71391 , n71390 , n71246 );
and ( n71392 , n71389 , n71391 );
xor ( n71393 , n71062 , n71066 );
xor ( n71394 , n71393 , n71069 );
and ( n71395 , n71391 , n71394 );
and ( n71396 , n71389 , n71394 );
or ( n71397 , n71392 , n71395 , n71396 );
and ( n71398 , n68192 , n65371 );
and ( n71399 , n67873 , n65369 );
nor ( n71400 , n71398 , n71399 );
xnor ( n71401 , n71400 , n65168 );
and ( n71402 , n71397 , n71401 );
xor ( n71403 , n71072 , n71076 );
xor ( n71404 , n71403 , n71079 );
and ( n71405 , n71401 , n71404 );
and ( n71406 , n71397 , n71404 );
or ( n71407 , n71402 , n71405 , n71406 );
and ( n71408 , n67307 , n65756 );
and ( n71409 , n67302 , n65754 );
nor ( n71410 , n71408 , n71409 );
xnor ( n71411 , n71410 , n65450 );
and ( n71412 , n71407 , n71411 );
xor ( n71413 , n71082 , n71086 );
xor ( n71414 , n71413 , n71089 );
and ( n71415 , n71411 , n71414 );
and ( n71416 , n71407 , n71414 );
or ( n71417 , n71412 , n71415 , n71416 );
and ( n71418 , n66276 , n66906 );
and ( n71419 , n66142 , n66904 );
nor ( n71420 , n71418 , n71419 );
xnor ( n71421 , n71420 , n66286 );
and ( n71422 , n71417 , n71421 );
xor ( n71423 , n71092 , n71269 );
xor ( n71424 , n71423 , n71272 );
and ( n71425 , n71421 , n71424 );
and ( n71426 , n71417 , n71424 );
or ( n71427 , n71422 , n71425 , n71426 );
and ( n71428 , n65698 , n67498 );
and ( n71429 , n65657 , n67495 );
nor ( n71430 , n71428 , n71429 );
xnor ( n71431 , n71430 , n66511 );
and ( n71432 , n71427 , n71431 );
xor ( n71433 , n71275 , n71279 );
xor ( n71434 , n71433 , n71282 );
and ( n71435 , n71431 , n71434 );
and ( n71436 , n71427 , n71434 );
or ( n71437 , n71432 , n71435 , n71436 );
and ( n71438 , n71373 , n71437 );
xor ( n71439 , n71012 , n71016 );
xor ( n71440 , n71439 , n71019 );
and ( n71441 , n71437 , n71440 );
and ( n71442 , n71373 , n71440 );
or ( n71443 , n71438 , n71441 , n71442 );
xor ( n71444 , n70978 , n70982 );
xor ( n71445 , n71444 , n70985 );
and ( n71446 , n71443 , n71445 );
xor ( n71447 , n71022 , n71026 );
xor ( n71448 , n71447 , n71029 );
and ( n71449 , n71445 , n71448 );
and ( n71450 , n71443 , n71448 );
or ( n71451 , n71446 , n71449 , n71450 );
xor ( n71452 , n70988 , n71032 );
xor ( n71453 , n71452 , n71035 );
and ( n71454 , n71451 , n71453 );
xor ( n71455 , n71327 , n71329 );
xor ( n71456 , n71455 , n71332 );
and ( n71457 , n71453 , n71456 );
and ( n71458 , n71451 , n71456 );
or ( n71459 , n71454 , n71457 , n71458 );
and ( n71460 , n71347 , n71459 );
xor ( n71461 , n71347 , n71459 );
xor ( n71462 , n71451 , n71453 );
xor ( n71463 , n71462 , n71456 );
and ( n71464 , n69095 , n65056 );
and ( n71465 , n68873 , n65054 );
nor ( n71466 , n71464 , n71465 );
xnor ( n71467 , n71466 , n64943 );
and ( n71468 , n69568 , n64897 );
and ( n71469 , n69449 , n64895 );
nor ( n71470 , n71468 , n71469 );
xnor ( n71471 , n71470 , n64850 );
and ( n71472 , n71467 , n71471 );
xor ( n71473 , n71191 , n71225 );
xor ( n71474 , n71473 , n71228 );
and ( n71475 , n71471 , n71474 );
and ( n71476 , n71467 , n71474 );
or ( n71477 , n71472 , n71475 , n71476 );
and ( n71478 , n68439 , n65371 );
and ( n71479 , n68199 , n65369 );
nor ( n71480 , n71478 , n71479 );
xnor ( n71481 , n71480 , n65168 );
and ( n71482 , n71477 , n71481 );
xor ( n71483 , n71106 , n71231 );
xor ( n71484 , n71483 , n71234 );
and ( n71485 , n71481 , n71484 );
and ( n71486 , n71477 , n71484 );
or ( n71487 , n71482 , n71485 , n71486 );
and ( n71488 , n67873 , n65550 );
and ( n71489 , n67833 , n65548 );
nor ( n71490 , n71488 , n71489 );
xnor ( n71491 , n71490 , n65313 );
and ( n71492 , n71487 , n71491 );
and ( n71493 , n68199 , n65371 );
and ( n71494 , n68192 , n65369 );
nor ( n71495 , n71493 , n71494 );
xnor ( n71496 , n71495 , n65168 );
and ( n71497 , n71491 , n71496 );
and ( n71498 , n71487 , n71496 );
or ( n71499 , n71492 , n71497 , n71498 );
and ( n71500 , n67302 , n66016 );
and ( n71501 , n67111 , n66014 );
nor ( n71502 , n71500 , n71501 );
xnor ( n71503 , n71502 , n65650 );
and ( n71504 , n71499 , n71503 );
xor ( n71505 , n71249 , n71253 );
xor ( n71506 , n71505 , n71256 );
and ( n71507 , n71503 , n71506 );
and ( n71508 , n71499 , n71506 );
or ( n71509 , n71504 , n71507 , n71508 );
and ( n71510 , n67111 , n66016 );
and ( n71511 , n66981 , n66014 );
nor ( n71512 , n71510 , n71511 );
xnor ( n71513 , n71512 , n65650 );
and ( n71514 , n71509 , n71513 );
xor ( n71515 , n71259 , n71263 );
xor ( n71516 , n71515 , n71266 );
and ( n71517 , n71513 , n71516 );
and ( n71518 , n71509 , n71516 );
or ( n71519 , n71514 , n71517 , n71518 );
and ( n71520 , n65883 , n67498 );
and ( n71521 , n65698 , n67495 );
nor ( n71522 , n71520 , n71521 );
xnor ( n71523 , n71522 , n66511 );
and ( n71524 , n71519 , n71523 );
and ( n71525 , n66517 , n66657 );
and ( n71526 , n66266 , n66655 );
nor ( n71527 , n71525 , n71526 );
xnor ( n71528 , n71527 , n66130 );
and ( n71529 , n71523 , n71528 );
and ( n71530 , n71519 , n71528 );
or ( n71531 , n71524 , n71529 , n71530 );
and ( n71532 , n66507 , n66657 );
and ( n71533 , n66517 , n66655 );
nor ( n71534 , n71532 , n71533 );
xnor ( n71535 , n71534 , n66130 );
and ( n71536 , n66786 , n66241 );
and ( n71537 , n66781 , n66239 );
nor ( n71538 , n71536 , n71537 );
xnor ( n71539 , n71538 , n65876 );
and ( n71540 , n71535 , n71539 );
xor ( n71541 , n71407 , n71411 );
xor ( n71542 , n71541 , n71414 );
and ( n71543 , n71539 , n71542 );
and ( n71544 , n71535 , n71542 );
or ( n71545 , n71540 , n71543 , n71544 );
and ( n71546 , n66137 , n67160 );
and ( n71547 , n65935 , n67158 );
nor ( n71548 , n71546 , n71547 );
xnor ( n71549 , n71548 , n66514 );
and ( n71550 , n71545 , n71549 );
xor ( n71551 , n71351 , n71355 );
xor ( n71552 , n71551 , n71358 );
and ( n71553 , n71549 , n71552 );
and ( n71554 , n71545 , n71552 );
or ( n71555 , n71550 , n71553 , n71554 );
and ( n71556 , n71531 , n71555 );
xor ( n71557 , n71301 , n71305 );
xor ( n71558 , n71557 , n71308 );
and ( n71559 , n71555 , n71558 );
and ( n71560 , n71531 , n71558 );
or ( n71561 , n71556 , n71559 , n71560 );
xor ( n71562 , n71285 , n71289 );
xor ( n71563 , n71562 , n71294 );
and ( n71564 , n71561 , n71563 );
xor ( n71565 , n71311 , n71315 );
xor ( n71566 , n71565 , n71318 );
and ( n71567 , n71563 , n71566 );
and ( n71568 , n71561 , n71566 );
or ( n71569 , n71564 , n71567 , n71568 );
xor ( n71570 , n71297 , n71321 );
xor ( n71571 , n71570 , n71324 );
and ( n71572 , n71569 , n71571 );
xor ( n71573 , n71443 , n71445 );
xor ( n71574 , n71573 , n71448 );
and ( n71575 , n71571 , n71574 );
and ( n71576 , n71569 , n71574 );
or ( n71577 , n71572 , n71575 , n71576 );
and ( n71578 , n71463 , n71577 );
xor ( n71579 , n71463 , n71577 );
xor ( n71580 , n71569 , n71571 );
xor ( n71581 , n71580 , n71574 );
and ( n71582 , n66781 , n66657 );
and ( n71583 , n66507 , n66655 );
nor ( n71584 , n71582 , n71583 );
xnor ( n71585 , n71584 , n66130 );
and ( n71586 , n66981 , n66241 );
and ( n71587 , n66786 , n66239 );
nor ( n71588 , n71586 , n71587 );
xnor ( n71589 , n71588 , n65876 );
and ( n71590 , n71585 , n71589 );
xor ( n71591 , n71499 , n71503 );
xor ( n71592 , n71591 , n71506 );
and ( n71593 , n71589 , n71592 );
and ( n71594 , n71585 , n71592 );
or ( n71595 , n71590 , n71593 , n71594 );
and ( n71596 , n67833 , n65756 );
and ( n71597 , n67727 , n65754 );
nor ( n71598 , n71596 , n71597 );
xnor ( n71599 , n71598 , n65450 );
and ( n71600 , n68192 , n65550 );
and ( n71601 , n67873 , n65548 );
nor ( n71602 , n71600 , n71601 );
xnor ( n71603 , n71602 , n65313 );
and ( n71604 , n71599 , n71603 );
xor ( n71605 , n71377 , n71381 );
xor ( n71606 , n71605 , n71386 );
and ( n71607 , n71603 , n71606 );
and ( n71608 , n71599 , n71606 );
or ( n71609 , n71604 , n71607 , n71608 );
and ( n71610 , n67727 , n65756 );
and ( n71611 , n67548 , n65754 );
nor ( n71612 , n71610 , n71611 );
xnor ( n71613 , n71612 , n65450 );
and ( n71614 , n71609 , n71613 );
xor ( n71615 , n71389 , n71391 );
xor ( n71616 , n71615 , n71394 );
and ( n71617 , n71613 , n71616 );
and ( n71618 , n71609 , n71616 );
or ( n71619 , n71614 , n71617 , n71618 );
and ( n71620 , n67548 , n65756 );
and ( n71621 , n67307 , n65754 );
nor ( n71622 , n71620 , n71621 );
xnor ( n71623 , n71622 , n65450 );
and ( n71624 , n71619 , n71623 );
xor ( n71625 , n71397 , n71401 );
xor ( n71626 , n71625 , n71404 );
and ( n71627 , n71623 , n71626 );
and ( n71628 , n71619 , n71626 );
or ( n71629 , n71624 , n71627 , n71628 );
and ( n71630 , n71595 , n71629 );
and ( n71631 , n66266 , n66906 );
and ( n71632 , n66276 , n66904 );
nor ( n71633 , n71631 , n71632 );
xnor ( n71634 , n71633 , n66286 );
and ( n71635 , n71629 , n71634 );
and ( n71636 , n71595 , n71634 );
or ( n71637 , n71630 , n71635 , n71636 );
and ( n71638 , n65935 , n67498 );
and ( n71639 , n65883 , n67495 );
nor ( n71640 , n71638 , n71639 );
xnor ( n71641 , n71640 , n66511 );
and ( n71642 , n66142 , n67160 );
and ( n71643 , n66137 , n67158 );
nor ( n71644 , n71642 , n71643 );
xnor ( n71645 , n71644 , n66514 );
and ( n71646 , n71641 , n71645 );
xor ( n71647 , n71509 , n71513 );
xor ( n71648 , n71647 , n71516 );
and ( n71649 , n71645 , n71648 );
and ( n71650 , n71641 , n71648 );
or ( n71651 , n71646 , n71649 , n71650 );
and ( n71652 , n71637 , n71651 );
xor ( n71653 , n71417 , n71421 );
xor ( n71654 , n71653 , n71424 );
and ( n71655 , n71651 , n71654 );
and ( n71656 , n71637 , n71654 );
or ( n71657 , n71652 , n71655 , n71656 );
xor ( n71658 , n71361 , n71365 );
xor ( n71659 , n71658 , n71370 );
and ( n71660 , n71657 , n71659 );
xor ( n71661 , n71427 , n71431 );
xor ( n71662 , n71661 , n71434 );
and ( n71663 , n71659 , n71662 );
and ( n71664 , n71657 , n71662 );
or ( n71665 , n71660 , n71663 , n71664 );
xor ( n71666 , n71373 , n71437 );
xor ( n71667 , n71666 , n71440 );
and ( n71668 , n71665 , n71667 );
xor ( n71669 , n71561 , n71563 );
xor ( n71670 , n71669 , n71566 );
and ( n71671 , n71667 , n71670 );
and ( n71672 , n71665 , n71670 );
or ( n71673 , n71668 , n71671 , n71672 );
and ( n71674 , n71581 , n71673 );
xor ( n71675 , n71581 , n71673 );
and ( n71676 , n69573 , n64897 );
and ( n71677 , n69566 , n64895 );
nor ( n71678 , n71676 , n71677 );
xnor ( n71679 , n71678 , n64850 );
and ( n71680 , n69985 , n64789 );
and ( n71681 , n69979 , n64787 );
nor ( n71682 , n71680 , n71681 );
xnor ( n71683 , n71682 , n64738 );
and ( n71684 , n71679 , n71683 );
xor ( n71685 , n71205 , n71209 );
xor ( n71686 , n71685 , n71212 );
and ( n71687 , n71683 , n71686 );
and ( n71688 , n71679 , n71686 );
or ( n71689 , n71684 , n71687 , n71688 );
and ( n71690 , n69449 , n65056 );
and ( n71691 , n69095 , n65054 );
nor ( n71692 , n71690 , n71691 );
xnor ( n71693 , n71692 , n64943 );
and ( n71694 , n71689 , n71693 );
xor ( n71695 , n71215 , n71219 );
xor ( n71696 , n71695 , n71222 );
and ( n71697 , n71693 , n71696 );
and ( n71698 , n71689 , n71696 );
or ( n71699 , n71694 , n71697 , n71698 );
and ( n71700 , n68444 , n65371 );
and ( n71701 , n68439 , n65369 );
nor ( n71702 , n71700 , n71701 );
xnor ( n71703 , n71702 , n65168 );
and ( n71704 , n71699 , n71703 );
and ( n71705 , n68837 , n65183 );
and ( n71706 , n68625 , n65181 );
nor ( n71707 , n71705 , n71706 );
xnor ( n71708 , n71707 , n64994 );
and ( n71709 , n71703 , n71708 );
and ( n71710 , n71699 , n71708 );
or ( n71711 , n71704 , n71709 , n71710 );
xor ( n71712 , n71110 , n71114 );
and ( n71713 , n70781 , n64709 );
not ( n71714 , n71713 );
and ( n71715 , n71714 , n64682 );
and ( n71716 , n70781 , n64711 );
and ( n71717 , n70786 , n64709 );
nor ( n71718 , n71716 , n71717 );
xnor ( n71719 , n71718 , n64682 );
and ( n71720 , n71715 , n71719 );
and ( n71721 , n70786 , n64711 );
and ( n71722 , n70792 , n64709 );
nor ( n71723 , n71721 , n71722 );
xnor ( n71724 , n71723 , n64682 );
and ( n71725 , n71720 , n71724 );
and ( n71726 , n71724 , n71108 );
and ( n71727 , n71720 , n71108 );
or ( n71728 , n71725 , n71726 , n71727 );
and ( n71729 , n71712 , n71728 );
and ( n71730 , n70792 , n64711 );
and ( n71731 , n70802 , n64709 );
nor ( n71732 , n71730 , n71731 );
xnor ( n71733 , n71732 , n64682 );
and ( n71734 , n71728 , n71733 );
and ( n71735 , n71712 , n71733 );
or ( n71736 , n71729 , n71734 , n71735 );
and ( n71737 , n70802 , n64711 );
and ( n71738 , n70812 , n64709 );
nor ( n71739 , n71737 , n71738 );
xnor ( n71740 , n71739 , n64682 );
and ( n71741 , n71736 , n71740 );
xor ( n71742 , n71115 , n71119 );
xor ( n71743 , n71742 , n70782 );
and ( n71744 , n71740 , n71743 );
and ( n71745 , n71736 , n71743 );
or ( n71746 , n71741 , n71744 , n71745 );
and ( n71747 , n70812 , n64711 );
and ( n71748 , n70822 , n64709 );
nor ( n71749 , n71747 , n71748 );
xnor ( n71750 , n71749 , n64682 );
and ( n71751 , n71746 , n71750 );
xor ( n71752 , n71107 , n71123 );
xor ( n71753 , n71752 , n71128 );
and ( n71754 , n71750 , n71753 );
and ( n71755 , n71746 , n71753 );
or ( n71756 , n71751 , n71754 , n71755 );
and ( n71757 , n70822 , n64711 );
and ( n71758 , n70832 , n64709 );
nor ( n71759 , n71757 , n71758 );
xnor ( n71760 , n71759 , n64682 );
and ( n71761 , n71756 , n71760 );
xor ( n71762 , n71131 , n71135 );
xor ( n71763 , n71762 , n71138 );
and ( n71764 , n71760 , n71763 );
and ( n71765 , n71756 , n71763 );
or ( n71766 , n71761 , n71764 , n71765 );
and ( n71767 , n70832 , n64711 );
and ( n71768 , n70766 , n64709 );
nor ( n71769 , n71767 , n71768 );
xnor ( n71770 , n71769 , n64682 );
and ( n71771 , n71766 , n71770 );
xor ( n71772 , n71141 , n71145 );
xor ( n71773 , n71772 , n71148 );
and ( n71774 , n71770 , n71773 );
and ( n71775 , n71766 , n71773 );
or ( n71776 , n71771 , n71774 , n71775 );
and ( n71777 , n70766 , n64711 );
and ( n71778 , n70266 , n64709 );
nor ( n71779 , n71777 , n71778 );
xnor ( n71780 , n71779 , n64682 );
and ( n71781 , n71776 , n71780 );
xor ( n71782 , n71151 , n71155 );
xor ( n71783 , n71782 , n71158 );
and ( n71784 , n71780 , n71783 );
and ( n71785 , n71776 , n71783 );
or ( n71786 , n71781 , n71784 , n71785 );
and ( n71787 , n69979 , n64897 );
and ( n71788 , n69573 , n64895 );
nor ( n71789 , n71787 , n71788 );
xnor ( n71790 , n71789 , n64850 );
and ( n71791 , n71786 , n71790 );
xor ( n71792 , n71195 , n71199 );
xor ( n71793 , n71792 , n71202 );
and ( n71794 , n71790 , n71793 );
and ( n71795 , n71786 , n71793 );
or ( n71796 , n71791 , n71794 , n71795 );
and ( n71797 , n70238 , n64897 );
and ( n71798 , n69985 , n64895 );
nor ( n71799 , n71797 , n71798 );
xnor ( n71800 , n71799 , n64850 );
and ( n71801 , n70266 , n64789 );
and ( n71802 , n70252 , n64787 );
nor ( n71803 , n71801 , n71802 );
xnor ( n71804 , n71803 , n64738 );
and ( n71805 , n71800 , n71804 );
xor ( n71806 , n71766 , n71770 );
xor ( n71807 , n71806 , n71773 );
and ( n71808 , n71804 , n71807 );
and ( n71809 , n71800 , n71807 );
or ( n71810 , n71805 , n71808 , n71809 );
and ( n71811 , n70252 , n64789 );
and ( n71812 , n70238 , n64787 );
nor ( n71813 , n71811 , n71812 );
xnor ( n71814 , n71813 , n64738 );
and ( n71815 , n71810 , n71814 );
xor ( n71816 , n71776 , n71780 );
xor ( n71817 , n71816 , n71783 );
and ( n71818 , n71814 , n71817 );
and ( n71819 , n71810 , n71817 );
or ( n71820 , n71815 , n71818 , n71819 );
and ( n71821 , n69566 , n65056 );
and ( n71822 , n69568 , n65054 );
nor ( n71823 , n71821 , n71822 );
xnor ( n71824 , n71823 , n64943 );
and ( n71825 , n71820 , n71824 );
xor ( n71826 , n71786 , n71790 );
xor ( n71827 , n71826 , n71793 );
and ( n71828 , n71824 , n71827 );
and ( n71829 , n71820 , n71827 );
or ( n71830 , n71825 , n71828 , n71829 );
and ( n71831 , n71796 , n71830 );
xor ( n71832 , n71679 , n71683 );
xor ( n71833 , n71832 , n71686 );
and ( n71834 , n71830 , n71833 );
and ( n71835 , n71796 , n71833 );
or ( n71836 , n71831 , n71834 , n71835 );
and ( n71837 , n68625 , n65371 );
and ( n71838 , n68444 , n65369 );
nor ( n71839 , n71837 , n71838 );
xnor ( n71840 , n71839 , n65168 );
and ( n71841 , n71836 , n71840 );
and ( n71842 , n68873 , n65183 );
and ( n71843 , n68837 , n65181 );
nor ( n71844 , n71842 , n71843 );
xnor ( n71845 , n71844 , n64994 );
and ( n71846 , n71840 , n71845 );
and ( n71847 , n71836 , n71845 );
or ( n71848 , n71841 , n71846 , n71847 );
and ( n71849 , n68199 , n65550 );
and ( n71850 , n68192 , n65548 );
nor ( n71851 , n71849 , n71850 );
xnor ( n71852 , n71851 , n65313 );
and ( n71853 , n71848 , n71852 );
xor ( n71854 , n71467 , n71471 );
xor ( n71855 , n71854 , n71474 );
and ( n71856 , n71852 , n71855 );
and ( n71857 , n71848 , n71855 );
or ( n71858 , n71853 , n71856 , n71857 );
and ( n71859 , n71711 , n71858 );
xor ( n71860 , n71477 , n71481 );
xor ( n71861 , n71860 , n71484 );
and ( n71862 , n71858 , n71861 );
and ( n71863 , n71711 , n71861 );
or ( n71864 , n71859 , n71862 , n71863 );
and ( n71865 , n67307 , n66016 );
and ( n71866 , n67302 , n66014 );
nor ( n71867 , n71865 , n71866 );
xnor ( n71868 , n71867 , n65650 );
and ( n71869 , n71864 , n71868 );
xor ( n71870 , n71487 , n71491 );
xor ( n71871 , n71870 , n71496 );
and ( n71872 , n71868 , n71871 );
and ( n71873 , n71864 , n71871 );
or ( n71874 , n71869 , n71872 , n71873 );
and ( n71875 , n66276 , n67160 );
and ( n71876 , n66142 , n67158 );
nor ( n71877 , n71875 , n71876 );
xnor ( n71878 , n71877 , n66514 );
and ( n71879 , n71874 , n71878 );
and ( n71880 , n66517 , n66906 );
and ( n71881 , n66266 , n66904 );
nor ( n71882 , n71880 , n71881 );
xnor ( n71883 , n71882 , n66286 );
and ( n71884 , n71878 , n71883 );
and ( n71885 , n71874 , n71883 );
or ( n71886 , n71879 , n71884 , n71885 );
xor ( n71887 , n71595 , n71629 );
xor ( n71888 , n71887 , n71634 );
and ( n71889 , n71886 , n71888 );
xor ( n71890 , n71535 , n71539 );
xor ( n71891 , n71890 , n71542 );
and ( n71892 , n71888 , n71891 );
and ( n71893 , n71886 , n71891 );
or ( n71894 , n71889 , n71892 , n71893 );
xor ( n71895 , n71519 , n71523 );
xor ( n71896 , n71895 , n71528 );
and ( n71897 , n71894 , n71896 );
xor ( n71898 , n71545 , n71549 );
xor ( n71899 , n71898 , n71552 );
and ( n71900 , n71896 , n71899 );
and ( n71901 , n71894 , n71899 );
or ( n71902 , n71897 , n71900 , n71901 );
xor ( n71903 , n71657 , n71659 );
xor ( n71904 , n71903 , n71662 );
and ( n71905 , n71902 , n71904 );
xor ( n71906 , n71531 , n71555 );
xor ( n71907 , n71906 , n71558 );
and ( n71908 , n71904 , n71907 );
and ( n71909 , n71902 , n71907 );
or ( n71910 , n71905 , n71908 , n71909 );
xor ( n71911 , n71665 , n71667 );
xor ( n71912 , n71911 , n71670 );
and ( n71913 , n71910 , n71912 );
xor ( n71914 , n71910 , n71912 );
xor ( n71915 , n71902 , n71904 );
xor ( n71916 , n71915 , n71907 );
and ( n71917 , n66781 , n66906 );
and ( n71918 , n66507 , n66904 );
nor ( n71919 , n71917 , n71918 );
xnor ( n71920 , n71919 , n66286 );
and ( n71921 , n66981 , n66657 );
and ( n71922 , n66786 , n66655 );
nor ( n71923 , n71921 , n71922 );
xnor ( n71924 , n71923 , n66130 );
and ( n71925 , n71920 , n71924 );
and ( n71926 , n69095 , n65183 );
and ( n71927 , n68873 , n65181 );
nor ( n71928 , n71926 , n71927 );
xnor ( n71929 , n71928 , n64994 );
and ( n71930 , n69568 , n65056 );
and ( n71931 , n69449 , n65054 );
nor ( n71932 , n71930 , n71931 );
xnor ( n71933 , n71932 , n64943 );
and ( n71934 , n71929 , n71933 );
xor ( n71935 , n71796 , n71830 );
xor ( n71936 , n71935 , n71833 );
and ( n71937 , n71933 , n71936 );
and ( n71938 , n71929 , n71936 );
or ( n71939 , n71934 , n71937 , n71938 );
and ( n71940 , n68439 , n65550 );
and ( n71941 , n68199 , n65548 );
nor ( n71942 , n71940 , n71941 );
xnor ( n71943 , n71942 , n65313 );
and ( n71944 , n71939 , n71943 );
xor ( n71945 , n71689 , n71693 );
xor ( n71946 , n71945 , n71696 );
and ( n71947 , n71943 , n71946 );
and ( n71948 , n71939 , n71946 );
or ( n71949 , n71944 , n71947 , n71948 );
and ( n71950 , n67873 , n65756 );
and ( n71951 , n67833 , n65754 );
nor ( n71952 , n71950 , n71951 );
xnor ( n71953 , n71952 , n65450 );
and ( n71954 , n71949 , n71953 );
xor ( n71955 , n71699 , n71703 );
xor ( n71956 , n71955 , n71708 );
and ( n71957 , n71953 , n71956 );
and ( n71958 , n71949 , n71956 );
or ( n71959 , n71954 , n71957 , n71958 );
and ( n71960 , n67302 , n66241 );
and ( n71961 , n67111 , n66239 );
nor ( n71962 , n71960 , n71961 );
xnor ( n71963 , n71962 , n65876 );
xor ( n71964 , n71959 , n71963 );
xor ( n71965 , n71599 , n71603 );
xor ( n71966 , n71965 , n71606 );
xor ( n71967 , n71964 , n71966 );
and ( n71968 , n71924 , n71967 );
and ( n71969 , n71920 , n71967 );
or ( n71970 , n71925 , n71968 , n71969 );
and ( n71971 , n69573 , n65056 );
and ( n71972 , n69566 , n65054 );
nor ( n71973 , n71971 , n71972 );
xnor ( n71974 , n71973 , n64943 );
and ( n71975 , n69985 , n64897 );
and ( n71976 , n69979 , n64895 );
nor ( n71977 , n71975 , n71976 );
xnor ( n71978 , n71977 , n64850 );
and ( n71979 , n71974 , n71978 );
xor ( n71980 , n71810 , n71814 );
xor ( n71981 , n71980 , n71817 );
and ( n71982 , n71978 , n71981 );
and ( n71983 , n71974 , n71981 );
or ( n71984 , n71979 , n71982 , n71983 );
and ( n71985 , n68873 , n65371 );
and ( n71986 , n68837 , n65369 );
nor ( n71987 , n71985 , n71986 );
xnor ( n71988 , n71987 , n65168 );
and ( n71989 , n71984 , n71988 );
xor ( n71990 , n71820 , n71824 );
xor ( n71991 , n71990 , n71827 );
and ( n71992 , n71988 , n71991 );
and ( n71993 , n71984 , n71991 );
or ( n71994 , n71989 , n71992 , n71993 );
and ( n71995 , n68444 , n65550 );
and ( n71996 , n68439 , n65548 );
nor ( n71997 , n71995 , n71996 );
xnor ( n71998 , n71997 , n65313 );
and ( n71999 , n71994 , n71998 );
and ( n72000 , n68837 , n65371 );
and ( n72001 , n68625 , n65369 );
nor ( n72002 , n72000 , n72001 );
xnor ( n72003 , n72002 , n65168 );
and ( n72004 , n71998 , n72003 );
and ( n72005 , n71994 , n72003 );
or ( n72006 , n71999 , n72004 , n72005 );
and ( n72007 , n67833 , n66016 );
and ( n72008 , n67727 , n66014 );
nor ( n72009 , n72007 , n72008 );
xnor ( n72010 , n72009 , n65650 );
and ( n72011 , n72006 , n72010 );
xor ( n72012 , n71836 , n71840 );
xor ( n72013 , n72012 , n71845 );
and ( n72014 , n72010 , n72013 );
and ( n72015 , n72006 , n72013 );
or ( n72016 , n72011 , n72014 , n72015 );
and ( n72017 , n67727 , n66016 );
and ( n72018 , n67548 , n66014 );
nor ( n72019 , n72017 , n72018 );
xnor ( n72020 , n72019 , n65650 );
and ( n72021 , n72016 , n72020 );
xor ( n72022 , n71848 , n71852 );
xor ( n72023 , n72022 , n71855 );
and ( n72024 , n72020 , n72023 );
and ( n72025 , n72016 , n72023 );
or ( n72026 , n72021 , n72024 , n72025 );
and ( n72027 , n67548 , n66016 );
and ( n72028 , n67307 , n66014 );
nor ( n72029 , n72027 , n72028 );
xnor ( n72030 , n72029 , n65650 );
and ( n72031 , n72026 , n72030 );
xor ( n72032 , n71711 , n71858 );
xor ( n72033 , n72032 , n71861 );
and ( n72034 , n72030 , n72033 );
and ( n72035 , n72026 , n72033 );
or ( n72036 , n72031 , n72034 , n72035 );
and ( n72037 , n71970 , n72036 );
and ( n72038 , n66266 , n67160 );
and ( n72039 , n66276 , n67158 );
nor ( n72040 , n72038 , n72039 );
xnor ( n72041 , n72040 , n66514 );
and ( n72042 , n72036 , n72041 );
and ( n72043 , n71970 , n72041 );
or ( n72044 , n72037 , n72042 , n72043 );
and ( n72045 , n66507 , n66906 );
and ( n72046 , n66517 , n66904 );
nor ( n72047 , n72045 , n72046 );
xnor ( n72048 , n72047 , n66286 );
and ( n72049 , n66786 , n66657 );
and ( n72050 , n66781 , n66655 );
nor ( n72051 , n72049 , n72050 );
xnor ( n72052 , n72051 , n66130 );
and ( n72053 , n72048 , n72052 );
xor ( n72054 , n71864 , n71868 );
xor ( n72055 , n72054 , n71871 );
and ( n72056 , n72052 , n72055 );
and ( n72057 , n72048 , n72055 );
or ( n72058 , n72053 , n72056 , n72057 );
and ( n72059 , n72044 , n72058 );
xor ( n72060 , n71585 , n71589 );
xor ( n72061 , n72060 , n71592 );
and ( n72062 , n72058 , n72061 );
and ( n72063 , n72044 , n72061 );
or ( n72064 , n72059 , n72062 , n72063 );
and ( n72065 , n71959 , n71963 );
and ( n72066 , n71963 , n71966 );
and ( n72067 , n71959 , n71966 );
or ( n72068 , n72065 , n72066 , n72067 );
and ( n72069 , n67111 , n66241 );
and ( n72070 , n66981 , n66239 );
nor ( n72071 , n72069 , n72070 );
xnor ( n72072 , n72071 , n65876 );
and ( n72073 , n72068 , n72072 );
xor ( n72074 , n71609 , n71613 );
xor ( n72075 , n72074 , n71616 );
and ( n72076 , n72072 , n72075 );
and ( n72077 , n72068 , n72075 );
or ( n72078 , n72073 , n72076 , n72077 );
and ( n72079 , n66137 , n67498 );
and ( n72080 , n65935 , n67495 );
nor ( n72081 , n72079 , n72080 );
xnor ( n72082 , n72081 , n66511 );
and ( n72083 , n72078 , n72082 );
xor ( n72084 , n71619 , n71623 );
xor ( n72085 , n72084 , n71626 );
and ( n72086 , n72082 , n72085 );
and ( n72087 , n72078 , n72085 );
or ( n72088 , n72083 , n72086 , n72087 );
and ( n72089 , n72064 , n72088 );
xor ( n72090 , n71641 , n71645 );
xor ( n72091 , n72090 , n71648 );
and ( n72092 , n72088 , n72091 );
and ( n72093 , n72064 , n72091 );
or ( n72094 , n72089 , n72092 , n72093 );
xor ( n72095 , n71894 , n71896 );
xor ( n72096 , n72095 , n71899 );
and ( n72097 , n72094 , n72096 );
xor ( n72098 , n71637 , n71651 );
xor ( n72099 , n72098 , n71654 );
and ( n72100 , n72096 , n72099 );
and ( n72101 , n72094 , n72099 );
or ( n72102 , n72097 , n72100 , n72101 );
and ( n72103 , n71916 , n72102 );
xor ( n72104 , n71916 , n72102 );
xor ( n72105 , n72094 , n72096 );
xor ( n72106 , n72105 , n72099 );
xor ( n72107 , n71715 , n71719 );
and ( n72108 , n70781 , n64787 );
not ( n72109 , n72108 );
and ( n72110 , n72109 , n64738 );
and ( n72111 , n70781 , n64789 );
and ( n72112 , n70786 , n64787 );
nor ( n72113 , n72111 , n72112 );
xnor ( n72114 , n72113 , n64738 );
and ( n72115 , n72110 , n72114 );
and ( n72116 , n70786 , n64789 );
and ( n72117 , n70792 , n64787 );
nor ( n72118 , n72116 , n72117 );
xnor ( n72119 , n72118 , n64738 );
and ( n72120 , n72115 , n72119 );
and ( n72121 , n72119 , n71713 );
and ( n72122 , n72115 , n71713 );
or ( n72123 , n72120 , n72121 , n72122 );
and ( n72124 , n72107 , n72123 );
and ( n72125 , n70792 , n64789 );
and ( n72126 , n70802 , n64787 );
nor ( n72127 , n72125 , n72126 );
xnor ( n72128 , n72127 , n64738 );
and ( n72129 , n72123 , n72128 );
and ( n72130 , n72107 , n72128 );
or ( n72131 , n72124 , n72129 , n72130 );
and ( n72132 , n70802 , n64789 );
and ( n72133 , n70812 , n64787 );
nor ( n72134 , n72132 , n72133 );
xnor ( n72135 , n72134 , n64738 );
and ( n72136 , n72131 , n72135 );
xor ( n72137 , n71720 , n71724 );
xor ( n72138 , n72137 , n71108 );
and ( n72139 , n72135 , n72138 );
and ( n72140 , n72131 , n72138 );
or ( n72141 , n72136 , n72139 , n72140 );
and ( n72142 , n70812 , n64789 );
and ( n72143 , n70822 , n64787 );
nor ( n72144 , n72142 , n72143 );
xnor ( n72145 , n72144 , n64738 );
and ( n72146 , n72141 , n72145 );
xor ( n72147 , n71712 , n71728 );
xor ( n72148 , n72147 , n71733 );
and ( n72149 , n72145 , n72148 );
and ( n72150 , n72141 , n72148 );
or ( n72151 , n72146 , n72149 , n72150 );
and ( n72152 , n70822 , n64789 );
and ( n72153 , n70832 , n64787 );
nor ( n72154 , n72152 , n72153 );
xnor ( n72155 , n72154 , n64738 );
and ( n72156 , n72151 , n72155 );
xor ( n72157 , n71736 , n71740 );
xor ( n72158 , n72157 , n71743 );
and ( n72159 , n72155 , n72158 );
and ( n72160 , n72151 , n72158 );
or ( n72161 , n72156 , n72159 , n72160 );
and ( n72162 , n70832 , n64789 );
and ( n72163 , n70766 , n64787 );
nor ( n72164 , n72162 , n72163 );
xnor ( n72165 , n72164 , n64738 );
and ( n72166 , n72161 , n72165 );
xor ( n72167 , n71746 , n71750 );
xor ( n72168 , n72167 , n71753 );
and ( n72169 , n72165 , n72168 );
and ( n72170 , n72161 , n72168 );
or ( n72171 , n72166 , n72169 , n72170 );
and ( n72172 , n70766 , n64789 );
and ( n72173 , n70266 , n64787 );
nor ( n72174 , n72172 , n72173 );
xnor ( n72175 , n72174 , n64738 );
and ( n72176 , n72171 , n72175 );
xor ( n72177 , n71756 , n71760 );
xor ( n72178 , n72177 , n71763 );
and ( n72179 , n72175 , n72178 );
and ( n72180 , n72171 , n72178 );
or ( n72181 , n72176 , n72179 , n72180 );
and ( n72182 , n69979 , n65056 );
and ( n72183 , n69573 , n65054 );
nor ( n72184 , n72182 , n72183 );
xnor ( n72185 , n72184 , n64943 );
and ( n72186 , n72181 , n72185 );
xor ( n72187 , n71800 , n71804 );
xor ( n72188 , n72187 , n71807 );
and ( n72189 , n72185 , n72188 );
and ( n72190 , n72181 , n72188 );
or ( n72191 , n72186 , n72189 , n72190 );
and ( n72192 , n70238 , n65056 );
and ( n72193 , n69985 , n65054 );
nor ( n72194 , n72192 , n72193 );
xnor ( n72195 , n72194 , n64943 );
and ( n72196 , n70266 , n64897 );
and ( n72197 , n70252 , n64895 );
nor ( n72198 , n72196 , n72197 );
xnor ( n72199 , n72198 , n64850 );
and ( n72200 , n72195 , n72199 );
xor ( n72201 , n72161 , n72165 );
xor ( n72202 , n72201 , n72168 );
and ( n72203 , n72199 , n72202 );
and ( n72204 , n72195 , n72202 );
or ( n72205 , n72200 , n72203 , n72204 );
and ( n72206 , n70252 , n64897 );
and ( n72207 , n70238 , n64895 );
nor ( n72208 , n72206 , n72207 );
xnor ( n72209 , n72208 , n64850 );
and ( n72210 , n72205 , n72209 );
xor ( n72211 , n72171 , n72175 );
xor ( n72212 , n72211 , n72178 );
and ( n72213 , n72209 , n72212 );
and ( n72214 , n72205 , n72212 );
or ( n72215 , n72210 , n72213 , n72214 );
and ( n72216 , n69566 , n65183 );
and ( n72217 , n69568 , n65181 );
nor ( n72218 , n72216 , n72217 );
xnor ( n72219 , n72218 , n64994 );
and ( n72220 , n72215 , n72219 );
xor ( n72221 , n72181 , n72185 );
xor ( n72222 , n72221 , n72188 );
and ( n72223 , n72219 , n72222 );
and ( n72224 , n72215 , n72222 );
or ( n72225 , n72220 , n72223 , n72224 );
and ( n72226 , n72191 , n72225 );
xor ( n72227 , n71974 , n71978 );
xor ( n72228 , n72227 , n71981 );
and ( n72229 , n72225 , n72228 );
and ( n72230 , n72191 , n72228 );
or ( n72231 , n72226 , n72229 , n72230 );
and ( n72232 , n68625 , n65550 );
and ( n72233 , n68444 , n65548 );
nor ( n72234 , n72232 , n72233 );
xnor ( n72235 , n72234 , n65313 );
and ( n72236 , n72231 , n72235 );
and ( n72237 , n69449 , n65183 );
and ( n72238 , n69095 , n65181 );
nor ( n72239 , n72237 , n72238 );
xnor ( n72240 , n72239 , n64994 );
and ( n72241 , n72235 , n72240 );
and ( n72242 , n72231 , n72240 );
or ( n72243 , n72236 , n72241 , n72242 );
and ( n72244 , n67873 , n66016 );
and ( n72245 , n67833 , n66014 );
nor ( n72246 , n72244 , n72245 );
xnor ( n72247 , n72246 , n65650 );
and ( n72248 , n72243 , n72247 );
xor ( n72249 , n71929 , n71933 );
xor ( n72250 , n72249 , n71936 );
and ( n72251 , n72247 , n72250 );
and ( n72252 , n72243 , n72250 );
or ( n72253 , n72248 , n72251 , n72252 );
and ( n72254 , n68192 , n65756 );
and ( n72255 , n67873 , n65754 );
nor ( n72256 , n72254 , n72255 );
xnor ( n72257 , n72256 , n65450 );
and ( n72258 , n72253 , n72257 );
xor ( n72259 , n71939 , n71943 );
xor ( n72260 , n72259 , n71946 );
and ( n72261 , n72257 , n72260 );
and ( n72262 , n72253 , n72260 );
or ( n72263 , n72258 , n72261 , n72262 );
and ( n72264 , n67307 , n66241 );
and ( n72265 , n67302 , n66239 );
nor ( n72266 , n72264 , n72265 );
xnor ( n72267 , n72266 , n65876 );
and ( n72268 , n72263 , n72267 );
xor ( n72269 , n71949 , n71953 );
xor ( n72270 , n72269 , n71956 );
and ( n72271 , n72267 , n72270 );
and ( n72272 , n72263 , n72270 );
or ( n72273 , n72268 , n72271 , n72272 );
and ( n72274 , n69095 , n65371 );
and ( n72275 , n68873 , n65369 );
nor ( n72276 , n72274 , n72275 );
xnor ( n72277 , n72276 , n65168 );
and ( n72278 , n69568 , n65183 );
and ( n72279 , n69449 , n65181 );
nor ( n72280 , n72278 , n72279 );
xnor ( n72281 , n72280 , n64994 );
and ( n72282 , n72277 , n72281 );
xor ( n72283 , n72191 , n72225 );
xor ( n72284 , n72283 , n72228 );
and ( n72285 , n72281 , n72284 );
and ( n72286 , n72277 , n72284 );
or ( n72287 , n72282 , n72285 , n72286 );
and ( n72288 , n68439 , n65756 );
and ( n72289 , n68199 , n65754 );
nor ( n72290 , n72288 , n72289 );
xnor ( n72291 , n72290 , n65450 );
and ( n72292 , n72287 , n72291 );
xor ( n72293 , n71984 , n71988 );
xor ( n72294 , n72293 , n71991 );
and ( n72295 , n72291 , n72294 );
and ( n72296 , n72287 , n72294 );
or ( n72297 , n72292 , n72295 , n72296 );
and ( n72298 , n68199 , n65756 );
and ( n72299 , n68192 , n65754 );
nor ( n72300 , n72298 , n72299 );
xnor ( n72301 , n72300 , n65450 );
and ( n72302 , n72297 , n72301 );
xor ( n72303 , n71994 , n71998 );
xor ( n72304 , n72303 , n72003 );
and ( n72305 , n72301 , n72304 );
and ( n72306 , n72297 , n72304 );
or ( n72307 , n72302 , n72305 , n72306 );
and ( n72308 , n67548 , n66241 );
and ( n72309 , n67307 , n66239 );
nor ( n72310 , n72308 , n72309 );
xnor ( n72311 , n72310 , n65876 );
and ( n72312 , n72307 , n72311 );
xor ( n72313 , n72006 , n72010 );
xor ( n72314 , n72313 , n72013 );
and ( n72315 , n72311 , n72314 );
and ( n72316 , n72307 , n72314 );
or ( n72317 , n72312 , n72315 , n72316 );
and ( n72318 , n67111 , n66657 );
and ( n72319 , n66981 , n66655 );
nor ( n72320 , n72318 , n72319 );
xnor ( n72321 , n72320 , n66130 );
and ( n72322 , n72317 , n72321 );
xor ( n72323 , n72016 , n72020 );
xor ( n72324 , n72323 , n72023 );
and ( n72325 , n72321 , n72324 );
and ( n72326 , n72317 , n72324 );
or ( n72327 , n72322 , n72325 , n72326 );
and ( n72328 , n72273 , n72327 );
xor ( n72329 , n72026 , n72030 );
xor ( n72330 , n72329 , n72033 );
and ( n72331 , n72327 , n72330 );
and ( n72332 , n72273 , n72330 );
or ( n72333 , n72328 , n72331 , n72332 );
and ( n72334 , n66142 , n67498 );
and ( n72335 , n66137 , n67495 );
nor ( n72336 , n72334 , n72335 );
xnor ( n72337 , n72336 , n66511 );
and ( n72338 , n72333 , n72337 );
xor ( n72339 , n72068 , n72072 );
xor ( n72340 , n72339 , n72075 );
and ( n72341 , n72337 , n72340 );
and ( n72342 , n72333 , n72340 );
or ( n72343 , n72338 , n72341 , n72342 );
xor ( n72344 , n71874 , n71878 );
xor ( n72345 , n72344 , n71883 );
and ( n72346 , n72343 , n72345 );
xor ( n72347 , n72078 , n72082 );
xor ( n72348 , n72347 , n72085 );
and ( n72349 , n72345 , n72348 );
and ( n72350 , n72343 , n72348 );
or ( n72351 , n72346 , n72349 , n72350 );
xor ( n72352 , n71886 , n71888 );
xor ( n72353 , n72352 , n71891 );
and ( n72354 , n72351 , n72353 );
xor ( n72355 , n72064 , n72088 );
xor ( n72356 , n72355 , n72091 );
and ( n72357 , n72353 , n72356 );
and ( n72358 , n72351 , n72356 );
or ( n72359 , n72354 , n72357 , n72358 );
and ( n72360 , n72106 , n72359 );
xor ( n72361 , n72106 , n72359 );
xor ( n72362 , n72351 , n72353 );
xor ( n72363 , n72362 , n72356 );
and ( n72364 , n66276 , n67498 );
and ( n72365 , n66142 , n67495 );
nor ( n72366 , n72364 , n72365 );
xnor ( n72367 , n72366 , n66511 );
and ( n72368 , n66517 , n67160 );
and ( n72369 , n66266 , n67158 );
nor ( n72370 , n72368 , n72369 );
xnor ( n72371 , n72370 , n66514 );
and ( n72372 , n72367 , n72371 );
xor ( n72373 , n71920 , n71924 );
xor ( n72374 , n72373 , n71967 );
and ( n72375 , n72371 , n72374 );
and ( n72376 , n72367 , n72374 );
or ( n72377 , n72372 , n72375 , n72376 );
xor ( n72378 , n71970 , n72036 );
xor ( n72379 , n72378 , n72041 );
and ( n72380 , n72377 , n72379 );
xor ( n72381 , n72048 , n72052 );
xor ( n72382 , n72381 , n72055 );
and ( n72383 , n72379 , n72382 );
and ( n72384 , n72377 , n72382 );
or ( n72385 , n72380 , n72383 , n72384 );
xor ( n72386 , n72044 , n72058 );
xor ( n72387 , n72386 , n72061 );
and ( n72388 , n72385 , n72387 );
xor ( n72389 , n72343 , n72345 );
xor ( n72390 , n72389 , n72348 );
and ( n72391 , n72387 , n72390 );
and ( n72392 , n72385 , n72390 );
or ( n72393 , n72388 , n72391 , n72392 );
and ( n72394 , n72363 , n72393 );
xor ( n72395 , n72363 , n72393 );
and ( n72396 , n66507 , n67160 );
and ( n72397 , n66517 , n67158 );
nor ( n72398 , n72396 , n72397 );
xnor ( n72399 , n72398 , n66514 );
and ( n72400 , n66786 , n66906 );
and ( n72401 , n66781 , n66904 );
nor ( n72402 , n72400 , n72401 );
xnor ( n72403 , n72402 , n66286 );
and ( n72404 , n72399 , n72403 );
xor ( n72405 , n72263 , n72267 );
xor ( n72406 , n72405 , n72270 );
and ( n72407 , n72403 , n72406 );
and ( n72408 , n72399 , n72406 );
or ( n72409 , n72404 , n72407 , n72408 );
and ( n72410 , n69573 , n65183 );
and ( n72411 , n69566 , n65181 );
nor ( n72412 , n72410 , n72411 );
xnor ( n72413 , n72412 , n64994 );
and ( n72414 , n69985 , n65056 );
and ( n72415 , n69979 , n65054 );
nor ( n72416 , n72414 , n72415 );
xnor ( n72417 , n72416 , n64943 );
and ( n72418 , n72413 , n72417 );
xor ( n72419 , n72205 , n72209 );
xor ( n72420 , n72419 , n72212 );
and ( n72421 , n72417 , n72420 );
and ( n72422 , n72413 , n72420 );
or ( n72423 , n72418 , n72421 , n72422 );
and ( n72424 , n69449 , n65371 );
and ( n72425 , n69095 , n65369 );
nor ( n72426 , n72424 , n72425 );
xnor ( n72427 , n72426 , n65168 );
and ( n72428 , n72423 , n72427 );
xor ( n72429 , n72215 , n72219 );
xor ( n72430 , n72429 , n72222 );
and ( n72431 , n72427 , n72430 );
and ( n72432 , n72423 , n72430 );
or ( n72433 , n72428 , n72431 , n72432 );
and ( n72434 , n68444 , n65756 );
and ( n72435 , n68439 , n65754 );
nor ( n72436 , n72434 , n72435 );
xnor ( n72437 , n72436 , n65450 );
and ( n72438 , n72433 , n72437 );
and ( n72439 , n68837 , n65550 );
and ( n72440 , n68625 , n65548 );
nor ( n72441 , n72439 , n72440 );
xnor ( n72442 , n72441 , n65313 );
and ( n72443 , n72437 , n72442 );
and ( n72444 , n72433 , n72442 );
or ( n72445 , n72438 , n72443 , n72444 );
and ( n72446 , n67833 , n66241 );
and ( n72447 , n67727 , n66239 );
nor ( n72448 , n72446 , n72447 );
xnor ( n72449 , n72448 , n65876 );
and ( n72450 , n72445 , n72449 );
xor ( n72451 , n72231 , n72235 );
xor ( n72452 , n72451 , n72240 );
and ( n72453 , n72449 , n72452 );
and ( n72454 , n72445 , n72452 );
or ( n72455 , n72450 , n72453 , n72454 );
and ( n72456 , n67727 , n66241 );
and ( n72457 , n67548 , n66239 );
nor ( n72458 , n72456 , n72457 );
xnor ( n72459 , n72458 , n65876 );
and ( n72460 , n72455 , n72459 );
xor ( n72461 , n72243 , n72247 );
xor ( n72462 , n72461 , n72250 );
and ( n72463 , n72459 , n72462 );
and ( n72464 , n72455 , n72462 );
or ( n72465 , n72460 , n72463 , n72464 );
and ( n72466 , n67302 , n66657 );
and ( n72467 , n67111 , n66655 );
nor ( n72468 , n72466 , n72467 );
xnor ( n72469 , n72468 , n66130 );
and ( n72470 , n72465 , n72469 );
xor ( n72471 , n72253 , n72257 );
xor ( n72472 , n72471 , n72260 );
and ( n72473 , n72469 , n72472 );
and ( n72474 , n72465 , n72472 );
or ( n72475 , n72470 , n72473 , n72474 );
and ( n72476 , n66266 , n67498 );
and ( n72477 , n66276 , n67495 );
nor ( n72478 , n72476 , n72477 );
xnor ( n72479 , n72478 , n66511 );
and ( n72480 , n72475 , n72479 );
xor ( n72481 , n72317 , n72321 );
xor ( n72482 , n72481 , n72324 );
and ( n72483 , n72479 , n72482 );
and ( n72484 , n72475 , n72482 );
or ( n72485 , n72480 , n72483 , n72484 );
and ( n72486 , n72409 , n72485 );
xor ( n72487 , n72273 , n72327 );
xor ( n72488 , n72487 , n72330 );
and ( n72489 , n72485 , n72488 );
and ( n72490 , n72409 , n72488 );
or ( n72491 , n72486 , n72489 , n72490 );
xor ( n72492 , n72377 , n72379 );
xor ( n72493 , n72492 , n72382 );
and ( n72494 , n72491 , n72493 );
xor ( n72495 , n72333 , n72337 );
xor ( n72496 , n72495 , n72340 );
and ( n72497 , n72493 , n72496 );
and ( n72498 , n72491 , n72496 );
or ( n72499 , n72494 , n72497 , n72498 );
xor ( n72500 , n72385 , n72387 );
xor ( n72501 , n72500 , n72390 );
and ( n72502 , n72499 , n72501 );
xor ( n72503 , n72499 , n72501 );
xor ( n72504 , n72491 , n72493 );
xor ( n72505 , n72504 , n72496 );
and ( n72506 , n66781 , n67160 );
and ( n72507 , n66507 , n67158 );
nor ( n72508 , n72506 , n72507 );
xnor ( n72509 , n72508 , n66514 );
and ( n72510 , n66981 , n66906 );
and ( n72511 , n66786 , n66904 );
nor ( n72512 , n72510 , n72511 );
xnor ( n72513 , n72512 , n66286 );
and ( n72514 , n72509 , n72513 );
xor ( n72515 , n72307 , n72311 );
xor ( n72516 , n72515 , n72314 );
and ( n72517 , n72513 , n72516 );
and ( n72518 , n72509 , n72516 );
or ( n72519 , n72514 , n72517 , n72518 );
xor ( n72520 , n72110 , n72114 );
and ( n72521 , n70781 , n64895 );
not ( n72522 , n72521 );
and ( n72523 , n72522 , n64850 );
and ( n72524 , n70781 , n64897 );
and ( n72525 , n70786 , n64895 );
nor ( n72526 , n72524 , n72525 );
xnor ( n72527 , n72526 , n64850 );
and ( n72528 , n72523 , n72527 );
and ( n72529 , n70786 , n64897 );
and ( n72530 , n70792 , n64895 );
nor ( n72531 , n72529 , n72530 );
xnor ( n72532 , n72531 , n64850 );
and ( n72533 , n72528 , n72532 );
and ( n72534 , n72532 , n72108 );
and ( n72535 , n72528 , n72108 );
or ( n72536 , n72533 , n72534 , n72535 );
and ( n72537 , n72520 , n72536 );
and ( n72538 , n70792 , n64897 );
and ( n72539 , n70802 , n64895 );
nor ( n72540 , n72538 , n72539 );
xnor ( n72541 , n72540 , n64850 );
and ( n72542 , n72536 , n72541 );
and ( n72543 , n72520 , n72541 );
or ( n72544 , n72537 , n72542 , n72543 );
and ( n72545 , n70802 , n64897 );
and ( n72546 , n70812 , n64895 );
nor ( n72547 , n72545 , n72546 );
xnor ( n72548 , n72547 , n64850 );
and ( n72549 , n72544 , n72548 );
xor ( n72550 , n72115 , n72119 );
xor ( n72551 , n72550 , n71713 );
and ( n72552 , n72548 , n72551 );
and ( n72553 , n72544 , n72551 );
or ( n72554 , n72549 , n72552 , n72553 );
and ( n72555 , n70812 , n64897 );
and ( n72556 , n70822 , n64895 );
nor ( n72557 , n72555 , n72556 );
xnor ( n72558 , n72557 , n64850 );
and ( n72559 , n72554 , n72558 );
xor ( n72560 , n72107 , n72123 );
xor ( n72561 , n72560 , n72128 );
and ( n72562 , n72558 , n72561 );
and ( n72563 , n72554 , n72561 );
or ( n72564 , n72559 , n72562 , n72563 );
and ( n72565 , n70822 , n64897 );
and ( n72566 , n70832 , n64895 );
nor ( n72567 , n72565 , n72566 );
xnor ( n72568 , n72567 , n64850 );
and ( n72569 , n72564 , n72568 );
xor ( n72570 , n72131 , n72135 );
xor ( n72571 , n72570 , n72138 );
and ( n72572 , n72568 , n72571 );
and ( n72573 , n72564 , n72571 );
or ( n72574 , n72569 , n72572 , n72573 );
and ( n72575 , n70832 , n64897 );
and ( n72576 , n70766 , n64895 );
nor ( n72577 , n72575 , n72576 );
xnor ( n72578 , n72577 , n64850 );
and ( n72579 , n72574 , n72578 );
xor ( n72580 , n72141 , n72145 );
xor ( n72581 , n72580 , n72148 );
and ( n72582 , n72578 , n72581 );
and ( n72583 , n72574 , n72581 );
or ( n72584 , n72579 , n72582 , n72583 );
and ( n72585 , n70766 , n64897 );
and ( n72586 , n70266 , n64895 );
nor ( n72587 , n72585 , n72586 );
xnor ( n72588 , n72587 , n64850 );
and ( n72589 , n72584 , n72588 );
xor ( n72590 , n72151 , n72155 );
xor ( n72591 , n72590 , n72158 );
and ( n72592 , n72588 , n72591 );
and ( n72593 , n72584 , n72591 );
or ( n72594 , n72589 , n72592 , n72593 );
and ( n72595 , n69979 , n65183 );
and ( n72596 , n69573 , n65181 );
nor ( n72597 , n72595 , n72596 );
xnor ( n72598 , n72597 , n64994 );
and ( n72599 , n72594 , n72598 );
xor ( n72600 , n72195 , n72199 );
xor ( n72601 , n72600 , n72202 );
and ( n72602 , n72598 , n72601 );
and ( n72603 , n72594 , n72601 );
or ( n72604 , n72599 , n72602 , n72603 );
and ( n72605 , n69985 , n65183 );
and ( n72606 , n69979 , n65181 );
nor ( n72607 , n72605 , n72606 );
xnor ( n72608 , n72607 , n64994 );
and ( n72609 , n70252 , n65056 );
and ( n72610 , n70238 , n65054 );
nor ( n72611 , n72609 , n72610 );
xnor ( n72612 , n72611 , n64943 );
and ( n72613 , n72608 , n72612 );
xor ( n72614 , n72584 , n72588 );
xor ( n72615 , n72614 , n72591 );
and ( n72616 , n72612 , n72615 );
and ( n72617 , n72608 , n72615 );
or ( n72618 , n72613 , n72616 , n72617 );
and ( n72619 , n69566 , n65371 );
and ( n72620 , n69568 , n65369 );
nor ( n72621 , n72619 , n72620 );
xnor ( n72622 , n72621 , n65168 );
and ( n72623 , n72618 , n72622 );
xor ( n72624 , n72594 , n72598 );
xor ( n72625 , n72624 , n72601 );
and ( n72626 , n72622 , n72625 );
and ( n72627 , n72618 , n72625 );
or ( n72628 , n72623 , n72626 , n72627 );
and ( n72629 , n72604 , n72628 );
xor ( n72630 , n72413 , n72417 );
xor ( n72631 , n72630 , n72420 );
and ( n72632 , n72628 , n72631 );
and ( n72633 , n72604 , n72631 );
or ( n72634 , n72629 , n72632 , n72633 );
and ( n72635 , n68625 , n65756 );
and ( n72636 , n68444 , n65754 );
nor ( n72637 , n72635 , n72636 );
xnor ( n72638 , n72637 , n65450 );
and ( n72639 , n72634 , n72638 );
and ( n72640 , n68873 , n65550 );
and ( n72641 , n68837 , n65548 );
nor ( n72642 , n72640 , n72641 );
xnor ( n72643 , n72642 , n65313 );
and ( n72644 , n72638 , n72643 );
and ( n72645 , n72634 , n72643 );
or ( n72646 , n72639 , n72644 , n72645 );
xor ( n72647 , n72433 , n72437 );
xor ( n72648 , n72647 , n72442 );
and ( n72649 , n72646 , n72648 );
xor ( n72650 , n72277 , n72281 );
xor ( n72651 , n72650 , n72284 );
and ( n72652 , n72648 , n72651 );
and ( n72653 , n72646 , n72651 );
or ( n72654 , n72649 , n72652 , n72653 );
and ( n72655 , n68192 , n66016 );
and ( n72656 , n67873 , n66014 );
nor ( n72657 , n72655 , n72656 );
xnor ( n72658 , n72657 , n65650 );
and ( n72659 , n72654 , n72658 );
xor ( n72660 , n72287 , n72291 );
xor ( n72661 , n72660 , n72294 );
and ( n72662 , n72658 , n72661 );
and ( n72663 , n72654 , n72661 );
or ( n72664 , n72659 , n72662 , n72663 );
and ( n72665 , n67307 , n66657 );
and ( n72666 , n67302 , n66655 );
nor ( n72667 , n72665 , n72666 );
xnor ( n72668 , n72667 , n66130 );
and ( n72669 , n72664 , n72668 );
xor ( n72670 , n72297 , n72301 );
xor ( n72671 , n72670 , n72304 );
and ( n72672 , n72668 , n72671 );
and ( n72673 , n72664 , n72671 );
or ( n72674 , n72669 , n72672 , n72673 );
and ( n72675 , n67302 , n66906 );
and ( n72676 , n67111 , n66904 );
nor ( n72677 , n72675 , n72676 );
xnor ( n72678 , n72677 , n66286 );
and ( n72679 , n67548 , n66657 );
and ( n72680 , n67307 , n66655 );
nor ( n72681 , n72679 , n72680 );
xnor ( n72682 , n72681 , n66130 );
and ( n72683 , n72678 , n72682 );
xor ( n72684 , n72445 , n72449 );
xor ( n72685 , n72684 , n72452 );
and ( n72686 , n72682 , n72685 );
and ( n72687 , n72678 , n72685 );
or ( n72688 , n72683 , n72686 , n72687 );
and ( n72689 , n67111 , n66906 );
and ( n72690 , n66981 , n66904 );
nor ( n72691 , n72689 , n72690 );
xnor ( n72692 , n72691 , n66286 );
and ( n72693 , n72688 , n72692 );
xor ( n72694 , n72455 , n72459 );
xor ( n72695 , n72694 , n72462 );
and ( n72696 , n72692 , n72695 );
and ( n72697 , n72688 , n72695 );
or ( n72698 , n72693 , n72696 , n72697 );
and ( n72699 , n72674 , n72698 );
xor ( n72700 , n72465 , n72469 );
xor ( n72701 , n72700 , n72472 );
and ( n72702 , n72698 , n72701 );
and ( n72703 , n72674 , n72701 );
or ( n72704 , n72699 , n72702 , n72703 );
and ( n72705 , n72519 , n72704 );
xor ( n72706 , n72399 , n72403 );
xor ( n72707 , n72706 , n72406 );
and ( n72708 , n72704 , n72707 );
and ( n72709 , n72519 , n72707 );
or ( n72710 , n72705 , n72708 , n72709 );
xor ( n72711 , n72367 , n72371 );
xor ( n72712 , n72711 , n72374 );
and ( n72713 , n72710 , n72712 );
xor ( n72714 , n72409 , n72485 );
xor ( n72715 , n72714 , n72488 );
and ( n72716 , n72712 , n72715 );
and ( n72717 , n72710 , n72715 );
or ( n72718 , n72713 , n72716 , n72717 );
and ( n72719 , n72505 , n72718 );
xor ( n72720 , n72505 , n72718 );
and ( n72721 , n69095 , n65550 );
and ( n72722 , n68873 , n65548 );
nor ( n72723 , n72721 , n72722 );
xnor ( n72724 , n72723 , n65313 );
and ( n72725 , n69568 , n65371 );
and ( n72726 , n69449 , n65369 );
nor ( n72727 , n72725 , n72726 );
xnor ( n72728 , n72727 , n65168 );
and ( n72729 , n72724 , n72728 );
xor ( n72730 , n72604 , n72628 );
xor ( n72731 , n72730 , n72631 );
and ( n72732 , n72728 , n72731 );
and ( n72733 , n72724 , n72731 );
or ( n72734 , n72729 , n72732 , n72733 );
and ( n72735 , n68439 , n66016 );
and ( n72736 , n68199 , n66014 );
nor ( n72737 , n72735 , n72736 );
xnor ( n72738 , n72737 , n65650 );
and ( n72739 , n72734 , n72738 );
xor ( n72740 , n72423 , n72427 );
xor ( n72741 , n72740 , n72430 );
and ( n72742 , n72738 , n72741 );
and ( n72743 , n72734 , n72741 );
or ( n72744 , n72739 , n72742 , n72743 );
and ( n72745 , n67873 , n66241 );
and ( n72746 , n67833 , n66239 );
nor ( n72747 , n72745 , n72746 );
xnor ( n72748 , n72747 , n65876 );
and ( n72749 , n72744 , n72748 );
and ( n72750 , n68199 , n66016 );
and ( n72751 , n68192 , n66014 );
nor ( n72752 , n72750 , n72751 );
xnor ( n72753 , n72752 , n65650 );
and ( n72754 , n72748 , n72753 );
and ( n72755 , n72744 , n72753 );
or ( n72756 , n72749 , n72754 , n72755 );
and ( n72757 , n70238 , n65183 );
and ( n72758 , n69985 , n65181 );
nor ( n72759 , n72757 , n72758 );
xnor ( n72760 , n72759 , n64994 );
and ( n72761 , n70266 , n65056 );
and ( n72762 , n70252 , n65054 );
nor ( n72763 , n72761 , n72762 );
xnor ( n72764 , n72763 , n64943 );
and ( n72765 , n72760 , n72764 );
xor ( n72766 , n72574 , n72578 );
xor ( n72767 , n72766 , n72581 );
and ( n72768 , n72764 , n72767 );
and ( n72769 , n72760 , n72767 );
or ( n72770 , n72765 , n72768 , n72769 );
and ( n72771 , n69573 , n65371 );
and ( n72772 , n69566 , n65369 );
nor ( n72773 , n72771 , n72772 );
xnor ( n72774 , n72773 , n65168 );
and ( n72775 , n72770 , n72774 );
xor ( n72776 , n72608 , n72612 );
xor ( n72777 , n72776 , n72615 );
and ( n72778 , n72774 , n72777 );
and ( n72779 , n72770 , n72777 );
or ( n72780 , n72775 , n72778 , n72779 );
and ( n72781 , n68873 , n65756 );
and ( n72782 , n68837 , n65754 );
nor ( n72783 , n72781 , n72782 );
xnor ( n72784 , n72783 , n65450 );
and ( n72785 , n72780 , n72784 );
xor ( n72786 , n72618 , n72622 );
xor ( n72787 , n72786 , n72625 );
and ( n72788 , n72784 , n72787 );
and ( n72789 , n72780 , n72787 );
or ( n72790 , n72785 , n72788 , n72789 );
and ( n72791 , n68444 , n66016 );
and ( n72792 , n68439 , n66014 );
nor ( n72793 , n72791 , n72792 );
xnor ( n72794 , n72793 , n65650 );
and ( n72795 , n72790 , n72794 );
and ( n72796 , n68837 , n65756 );
and ( n72797 , n68625 , n65754 );
nor ( n72798 , n72796 , n72797 );
xnor ( n72799 , n72798 , n65450 );
and ( n72800 , n72794 , n72799 );
and ( n72801 , n72790 , n72799 );
or ( n72802 , n72795 , n72800 , n72801 );
and ( n72803 , n68192 , n66241 );
and ( n72804 , n67873 , n66239 );
nor ( n72805 , n72803 , n72804 );
xnor ( n72806 , n72805 , n65876 );
and ( n72807 , n72802 , n72806 );
xor ( n72808 , n72634 , n72638 );
xor ( n72809 , n72808 , n72643 );
and ( n72810 , n72806 , n72809 );
and ( n72811 , n72802 , n72809 );
or ( n72812 , n72807 , n72810 , n72811 );
and ( n72813 , n67727 , n66657 );
and ( n72814 , n67548 , n66655 );
nor ( n72815 , n72813 , n72814 );
xnor ( n72816 , n72815 , n66130 );
and ( n72817 , n72812 , n72816 );
xor ( n72818 , n72646 , n72648 );
xor ( n72819 , n72818 , n72651 );
and ( n72820 , n72816 , n72819 );
and ( n72821 , n72812 , n72819 );
or ( n72822 , n72817 , n72820 , n72821 );
and ( n72823 , n72756 , n72822 );
xor ( n72824 , n72654 , n72658 );
xor ( n72825 , n72824 , n72661 );
and ( n72826 , n72822 , n72825 );
and ( n72827 , n72756 , n72825 );
or ( n72828 , n72823 , n72826 , n72827 );
and ( n72829 , n66507 , n67498 );
and ( n72830 , n66517 , n67495 );
nor ( n72831 , n72829 , n72830 );
xnor ( n72832 , n72831 , n66511 );
and ( n72833 , n72828 , n72832 );
and ( n72834 , n66786 , n67160 );
and ( n72835 , n66781 , n67158 );
nor ( n72836 , n72834 , n72835 );
xnor ( n72837 , n72836 , n66514 );
and ( n72838 , n72832 , n72837 );
and ( n72839 , n72828 , n72837 );
or ( n72840 , n72833 , n72838 , n72839 );
and ( n72841 , n66517 , n67498 );
and ( n72842 , n66266 , n67495 );
nor ( n72843 , n72841 , n72842 );
xnor ( n72844 , n72843 , n66511 );
and ( n72845 , n72840 , n72844 );
xor ( n72846 , n72509 , n72513 );
xor ( n72847 , n72846 , n72516 );
and ( n72848 , n72844 , n72847 );
and ( n72849 , n72840 , n72847 );
or ( n72850 , n72845 , n72848 , n72849 );
xor ( n72851 , n72519 , n72704 );
xor ( n72852 , n72851 , n72707 );
and ( n72853 , n72850 , n72852 );
xor ( n72854 , n72475 , n72479 );
xor ( n72855 , n72854 , n72482 );
and ( n72856 , n72852 , n72855 );
and ( n72857 , n72850 , n72855 );
or ( n72858 , n72853 , n72856 , n72857 );
xor ( n72859 , n72710 , n72712 );
xor ( n72860 , n72859 , n72715 );
and ( n72861 , n72858 , n72860 );
xor ( n72862 , n72858 , n72860 );
xor ( n72863 , n72850 , n72852 );
xor ( n72864 , n72863 , n72855 );
and ( n72865 , n66781 , n67498 );
and ( n72866 , n66507 , n67495 );
nor ( n72867 , n72865 , n72866 );
xnor ( n72868 , n72867 , n66511 );
and ( n72869 , n66981 , n67160 );
and ( n72870 , n66786 , n67158 );
nor ( n72871 , n72869 , n72870 );
xnor ( n72872 , n72871 , n66514 );
and ( n72873 , n72868 , n72872 );
xor ( n72874 , n72678 , n72682 );
xor ( n72875 , n72874 , n72685 );
and ( n72876 , n72872 , n72875 );
and ( n72877 , n72868 , n72875 );
or ( n72878 , n72873 , n72876 , n72877 );
xor ( n72879 , n72664 , n72668 );
xor ( n72880 , n72879 , n72671 );
and ( n72881 , n72878 , n72880 );
xor ( n72882 , n72688 , n72692 );
xor ( n72883 , n72882 , n72695 );
and ( n72884 , n72880 , n72883 );
and ( n72885 , n72878 , n72883 );
or ( n72886 , n72881 , n72884 , n72885 );
xor ( n72887 , n72840 , n72844 );
xor ( n72888 , n72887 , n72847 );
and ( n72889 , n72886 , n72888 );
xor ( n72890 , n72674 , n72698 );
xor ( n72891 , n72890 , n72701 );
and ( n72892 , n72888 , n72891 );
and ( n72893 , n72886 , n72891 );
or ( n72894 , n72889 , n72892 , n72893 );
and ( n72895 , n72864 , n72894 );
xor ( n72896 , n72864 , n72894 );
xor ( n72897 , n72886 , n72888 );
xor ( n72898 , n72897 , n72891 );
xor ( n72899 , n72523 , n72527 );
and ( n72900 , n70781 , n65054 );
not ( n72901 , n72900 );
and ( n72902 , n72901 , n64943 );
and ( n72903 , n70781 , n65056 );
and ( n72904 , n70786 , n65054 );
nor ( n72905 , n72903 , n72904 );
xnor ( n72906 , n72905 , n64943 );
and ( n72907 , n72902 , n72906 );
and ( n72908 , n70786 , n65056 );
and ( n72909 , n70792 , n65054 );
nor ( n72910 , n72908 , n72909 );
xnor ( n72911 , n72910 , n64943 );
and ( n72912 , n72907 , n72911 );
and ( n72913 , n72911 , n72521 );
and ( n72914 , n72907 , n72521 );
or ( n72915 , n72912 , n72913 , n72914 );
and ( n72916 , n72899 , n72915 );
and ( n72917 , n70792 , n65056 );
and ( n72918 , n70802 , n65054 );
nor ( n72919 , n72917 , n72918 );
xnor ( n72920 , n72919 , n64943 );
and ( n72921 , n72915 , n72920 );
and ( n72922 , n72899 , n72920 );
or ( n72923 , n72916 , n72921 , n72922 );
and ( n72924 , n70802 , n65056 );
and ( n72925 , n70812 , n65054 );
nor ( n72926 , n72924 , n72925 );
xnor ( n72927 , n72926 , n64943 );
and ( n72928 , n72923 , n72927 );
xor ( n72929 , n72528 , n72532 );
xor ( n72930 , n72929 , n72108 );
and ( n72931 , n72927 , n72930 );
and ( n72932 , n72923 , n72930 );
or ( n72933 , n72928 , n72931 , n72932 );
and ( n72934 , n70812 , n65056 );
and ( n72935 , n70822 , n65054 );
nor ( n72936 , n72934 , n72935 );
xnor ( n72937 , n72936 , n64943 );
and ( n72938 , n72933 , n72937 );
xor ( n72939 , n72520 , n72536 );
xor ( n72940 , n72939 , n72541 );
and ( n72941 , n72937 , n72940 );
and ( n72942 , n72933 , n72940 );
or ( n72943 , n72938 , n72941 , n72942 );
and ( n72944 , n70822 , n65056 );
and ( n72945 , n70832 , n65054 );
nor ( n72946 , n72944 , n72945 );
xnor ( n72947 , n72946 , n64943 );
and ( n72948 , n72943 , n72947 );
xor ( n72949 , n72544 , n72548 );
xor ( n72950 , n72949 , n72551 );
and ( n72951 , n72947 , n72950 );
and ( n72952 , n72943 , n72950 );
or ( n72953 , n72948 , n72951 , n72952 );
and ( n72954 , n70832 , n65056 );
and ( n72955 , n70766 , n65054 );
nor ( n72956 , n72954 , n72955 );
xnor ( n72957 , n72956 , n64943 );
and ( n72958 , n72953 , n72957 );
xor ( n72959 , n72554 , n72558 );
xor ( n72960 , n72959 , n72561 );
and ( n72961 , n72957 , n72960 );
and ( n72962 , n72953 , n72960 );
or ( n72963 , n72958 , n72961 , n72962 );
and ( n72964 , n70766 , n65056 );
and ( n72965 , n70266 , n65054 );
nor ( n72966 , n72964 , n72965 );
xnor ( n72967 , n72966 , n64943 );
and ( n72968 , n72963 , n72967 );
xor ( n72969 , n72564 , n72568 );
xor ( n72970 , n72969 , n72571 );
and ( n72971 , n72967 , n72970 );
and ( n72972 , n72963 , n72970 );
or ( n72973 , n72968 , n72971 , n72972 );
and ( n72974 , n69979 , n65371 );
and ( n72975 , n69573 , n65369 );
nor ( n72976 , n72974 , n72975 );
xnor ( n72977 , n72976 , n65168 );
and ( n72978 , n72973 , n72977 );
xor ( n72979 , n72760 , n72764 );
xor ( n72980 , n72979 , n72767 );
and ( n72981 , n72977 , n72980 );
and ( n72982 , n72973 , n72980 );
or ( n72983 , n72978 , n72981 , n72982 );
and ( n72984 , n70238 , n65371 );
and ( n72985 , n69985 , n65369 );
nor ( n72986 , n72984 , n72985 );
xnor ( n72987 , n72986 , n65168 );
and ( n72988 , n70266 , n65183 );
and ( n72989 , n70252 , n65181 );
nor ( n72990 , n72988 , n72989 );
xnor ( n72991 , n72990 , n64994 );
and ( n72992 , n72987 , n72991 );
xor ( n72993 , n72953 , n72957 );
xor ( n72994 , n72993 , n72960 );
and ( n72995 , n72991 , n72994 );
and ( n72996 , n72987 , n72994 );
or ( n72997 , n72992 , n72995 , n72996 );
and ( n72998 , n70252 , n65183 );
and ( n72999 , n70238 , n65181 );
nor ( n73000 , n72998 , n72999 );
xnor ( n73001 , n73000 , n64994 );
and ( n73002 , n72997 , n73001 );
xor ( n73003 , n72963 , n72967 );
xor ( n73004 , n73003 , n72970 );
and ( n73005 , n73001 , n73004 );
and ( n73006 , n72997 , n73004 );
or ( n73007 , n73002 , n73005 , n73006 );
and ( n73008 , n69566 , n65550 );
and ( n73009 , n69568 , n65548 );
nor ( n73010 , n73008 , n73009 );
xnor ( n73011 , n73010 , n65313 );
and ( n73012 , n73007 , n73011 );
xor ( n73013 , n72973 , n72977 );
xor ( n73014 , n73013 , n72980 );
and ( n73015 , n73011 , n73014 );
and ( n73016 , n73007 , n73014 );
or ( n73017 , n73012 , n73015 , n73016 );
and ( n73018 , n72983 , n73017 );
xor ( n73019 , n72770 , n72774 );
xor ( n73020 , n73019 , n72777 );
and ( n73021 , n73017 , n73020 );
and ( n73022 , n72983 , n73020 );
or ( n73023 , n73018 , n73021 , n73022 );
and ( n73024 , n68625 , n66016 );
and ( n73025 , n68444 , n66014 );
nor ( n73026 , n73024 , n73025 );
xnor ( n73027 , n73026 , n65650 );
and ( n73028 , n73023 , n73027 );
and ( n73029 , n69449 , n65550 );
and ( n73030 , n69095 , n65548 );
nor ( n73031 , n73029 , n73030 );
xnor ( n73032 , n73031 , n65313 );
and ( n73033 , n73027 , n73032 );
and ( n73034 , n73023 , n73032 );
or ( n73035 , n73028 , n73033 , n73034 );
and ( n73036 , n68199 , n66241 );
and ( n73037 , n68192 , n66239 );
nor ( n73038 , n73036 , n73037 );
xnor ( n73039 , n73038 , n65876 );
and ( n73040 , n73035 , n73039 );
xor ( n73041 , n72724 , n72728 );
xor ( n73042 , n73041 , n72731 );
and ( n73043 , n73039 , n73042 );
and ( n73044 , n73035 , n73042 );
or ( n73045 , n73040 , n73043 , n73044 );
and ( n73046 , n67833 , n66657 );
and ( n73047 , n67727 , n66655 );
nor ( n73048 , n73046 , n73047 );
xnor ( n73049 , n73048 , n66130 );
and ( n73050 , n73045 , n73049 );
xor ( n73051 , n72734 , n72738 );
xor ( n73052 , n73051 , n72741 );
and ( n73053 , n73049 , n73052 );
and ( n73054 , n73045 , n73052 );
or ( n73055 , n73050 , n73053 , n73054 );
and ( n73056 , n67307 , n66906 );
and ( n73057 , n67302 , n66904 );
nor ( n73058 , n73056 , n73057 );
xnor ( n73059 , n73058 , n66286 );
and ( n73060 , n73055 , n73059 );
xor ( n73061 , n72744 , n72748 );
xor ( n73062 , n73061 , n72753 );
and ( n73063 , n73059 , n73062 );
and ( n73064 , n73055 , n73062 );
or ( n73065 , n73060 , n73063 , n73064 );
and ( n73066 , n69095 , n65756 );
and ( n73067 , n68873 , n65754 );
nor ( n73068 , n73066 , n73067 );
xnor ( n73069 , n73068 , n65450 );
and ( n73070 , n69568 , n65550 );
and ( n73071 , n69449 , n65548 );
nor ( n73072 , n73070 , n73071 );
xnor ( n73073 , n73072 , n65313 );
and ( n73074 , n73069 , n73073 );
xor ( n73075 , n72983 , n73017 );
xor ( n73076 , n73075 , n73020 );
and ( n73077 , n73073 , n73076 );
and ( n73078 , n73069 , n73076 );
or ( n73079 , n73074 , n73077 , n73078 );
and ( n73080 , n68439 , n66241 );
and ( n73081 , n68199 , n66239 );
nor ( n73082 , n73080 , n73081 );
xnor ( n73083 , n73082 , n65876 );
and ( n73084 , n73079 , n73083 );
xor ( n73085 , n72780 , n72784 );
xor ( n73086 , n73085 , n72787 );
and ( n73087 , n73083 , n73086 );
and ( n73088 , n73079 , n73086 );
or ( n73089 , n73084 , n73087 , n73088 );
and ( n73090 , n67873 , n66657 );
and ( n73091 , n67833 , n66655 );
nor ( n73092 , n73090 , n73091 );
xnor ( n73093 , n73092 , n66130 );
and ( n73094 , n73089 , n73093 );
xor ( n73095 , n72790 , n72794 );
xor ( n73096 , n73095 , n72799 );
and ( n73097 , n73093 , n73096 );
and ( n73098 , n73089 , n73096 );
or ( n73099 , n73094 , n73097 , n73098 );
and ( n73100 , n67548 , n66906 );
and ( n73101 , n67307 , n66904 );
nor ( n73102 , n73100 , n73101 );
xnor ( n73103 , n73102 , n66286 );
and ( n73104 , n73099 , n73103 );
xor ( n73105 , n72802 , n72806 );
xor ( n73106 , n73105 , n72809 );
and ( n73107 , n73103 , n73106 );
and ( n73108 , n73099 , n73106 );
or ( n73109 , n73104 , n73107 , n73108 );
and ( n73110 , n67111 , n67160 );
and ( n73111 , n66981 , n67158 );
nor ( n73112 , n73110 , n73111 );
xnor ( n73113 , n73112 , n66514 );
and ( n73114 , n73109 , n73113 );
xor ( n73115 , n72812 , n72816 );
xor ( n73116 , n73115 , n72819 );
and ( n73117 , n73113 , n73116 );
and ( n73118 , n73109 , n73116 );
or ( n73119 , n73114 , n73117 , n73118 );
and ( n73120 , n73065 , n73119 );
xor ( n73121 , n72756 , n72822 );
xor ( n73122 , n73121 , n72825 );
and ( n73123 , n73119 , n73122 );
and ( n73124 , n73065 , n73122 );
or ( n73125 , n73120 , n73123 , n73124 );
xor ( n73126 , n72828 , n72832 );
xor ( n73127 , n73126 , n72837 );
and ( n73128 , n73125 , n73127 );
xor ( n73129 , n72878 , n72880 );
xor ( n73130 , n73129 , n72883 );
and ( n73131 , n73127 , n73130 );
and ( n73132 , n73125 , n73130 );
or ( n73133 , n73128 , n73131 , n73132 );
and ( n73134 , n72898 , n73133 );
xor ( n73135 , n72898 , n73133 );
xor ( n73136 , n73125 , n73127 );
xor ( n73137 , n73136 , n73130 );
and ( n73138 , n67833 , n66906 );
and ( n73139 , n67727 , n66904 );
nor ( n73140 , n73138 , n73139 );
xnor ( n73141 , n73140 , n66286 );
and ( n73142 , n68192 , n66657 );
and ( n73143 , n67873 , n66655 );
nor ( n73144 , n73142 , n73143 );
xnor ( n73145 , n73144 , n66130 );
and ( n73146 , n73141 , n73145 );
xor ( n73147 , n73023 , n73027 );
xor ( n73148 , n73147 , n73032 );
and ( n73149 , n73145 , n73148 );
and ( n73150 , n73141 , n73148 );
or ( n73151 , n73146 , n73149 , n73150 );
and ( n73152 , n67727 , n66906 );
and ( n73153 , n67548 , n66904 );
nor ( n73154 , n73152 , n73153 );
xnor ( n73155 , n73154 , n66286 );
and ( n73156 , n73151 , n73155 );
xor ( n73157 , n73035 , n73039 );
xor ( n73158 , n73157 , n73042 );
and ( n73159 , n73155 , n73158 );
and ( n73160 , n73151 , n73158 );
or ( n73161 , n73156 , n73159 , n73160 );
and ( n73162 , n67302 , n67160 );
and ( n73163 , n67111 , n67158 );
nor ( n73164 , n73162 , n73163 );
xnor ( n73165 , n73164 , n66514 );
and ( n73166 , n73161 , n73165 );
xor ( n73167 , n73045 , n73049 );
xor ( n73168 , n73167 , n73052 );
and ( n73169 , n73165 , n73168 );
and ( n73170 , n73161 , n73168 );
or ( n73171 , n73166 , n73169 , n73170 );
and ( n73172 , n66786 , n67498 );
and ( n73173 , n66781 , n67495 );
nor ( n73174 , n73172 , n73173 );
xnor ( n73175 , n73174 , n66511 );
and ( n73176 , n73171 , n73175 );
xor ( n73177 , n73055 , n73059 );
xor ( n73178 , n73177 , n73062 );
and ( n73179 , n73175 , n73178 );
and ( n73180 , n73171 , n73178 );
or ( n73181 , n73176 , n73179 , n73180 );
xor ( n73182 , n72868 , n72872 );
xor ( n73183 , n73182 , n72875 );
and ( n73184 , n73181 , n73183 );
xor ( n73185 , n73065 , n73119 );
xor ( n73186 , n73185 , n73122 );
and ( n73187 , n73183 , n73186 );
and ( n73188 , n73181 , n73186 );
or ( n73189 , n73184 , n73187 , n73188 );
and ( n73190 , n73137 , n73189 );
xor ( n73191 , n73137 , n73189 );
and ( n73192 , n69573 , n65550 );
and ( n73193 , n69566 , n65548 );
nor ( n73194 , n73192 , n73193 );
xnor ( n73195 , n73194 , n65313 );
and ( n73196 , n69985 , n65371 );
and ( n73197 , n69979 , n65369 );
nor ( n73198 , n73196 , n73197 );
xnor ( n73199 , n73198 , n65168 );
and ( n73200 , n73195 , n73199 );
xor ( n73201 , n72997 , n73001 );
xor ( n73202 , n73201 , n73004 );
and ( n73203 , n73199 , n73202 );
and ( n73204 , n73195 , n73202 );
or ( n73205 , n73200 , n73203 , n73204 );
and ( n73206 , n68873 , n66016 );
and ( n73207 , n68837 , n66014 );
nor ( n73208 , n73206 , n73207 );
xnor ( n73209 , n73208 , n65650 );
and ( n73210 , n73205 , n73209 );
xor ( n73211 , n73007 , n73011 );
xor ( n73212 , n73211 , n73014 );
and ( n73213 , n73209 , n73212 );
and ( n73214 , n73205 , n73212 );
or ( n73215 , n73210 , n73213 , n73214 );
and ( n73216 , n68444 , n66241 );
and ( n73217 , n68439 , n66239 );
nor ( n73218 , n73216 , n73217 );
xnor ( n73219 , n73218 , n65876 );
and ( n73220 , n73215 , n73219 );
and ( n73221 , n68837 , n66016 );
and ( n73222 , n68625 , n66014 );
nor ( n73223 , n73221 , n73222 );
xnor ( n73224 , n73223 , n65650 );
and ( n73225 , n73219 , n73224 );
and ( n73226 , n73215 , n73224 );
or ( n73227 , n73220 , n73225 , n73226 );
xor ( n73228 , n72902 , n72906 );
and ( n73229 , n70781 , n65181 );
not ( n73230 , n73229 );
and ( n73231 , n73230 , n64994 );
and ( n73232 , n70781 , n65183 );
and ( n73233 , n70786 , n65181 );
nor ( n73234 , n73232 , n73233 );
xnor ( n73235 , n73234 , n64994 );
and ( n73236 , n73231 , n73235 );
and ( n73237 , n70786 , n65183 );
and ( n73238 , n70792 , n65181 );
nor ( n73239 , n73237 , n73238 );
xnor ( n73240 , n73239 , n64994 );
and ( n73241 , n73236 , n73240 );
and ( n73242 , n73240 , n72900 );
and ( n73243 , n73236 , n72900 );
or ( n73244 , n73241 , n73242 , n73243 );
and ( n73245 , n73228 , n73244 );
and ( n73246 , n70792 , n65183 );
and ( n73247 , n70802 , n65181 );
nor ( n73248 , n73246 , n73247 );
xnor ( n73249 , n73248 , n64994 );
and ( n73250 , n73244 , n73249 );
and ( n73251 , n73228 , n73249 );
or ( n73252 , n73245 , n73250 , n73251 );
and ( n73253 , n70802 , n65183 );
and ( n73254 , n70812 , n65181 );
nor ( n73255 , n73253 , n73254 );
xnor ( n73256 , n73255 , n64994 );
and ( n73257 , n73252 , n73256 );
xor ( n73258 , n72907 , n72911 );
xor ( n73259 , n73258 , n72521 );
and ( n73260 , n73256 , n73259 );
and ( n73261 , n73252 , n73259 );
or ( n73262 , n73257 , n73260 , n73261 );
and ( n73263 , n70812 , n65183 );
and ( n73264 , n70822 , n65181 );
nor ( n73265 , n73263 , n73264 );
xnor ( n73266 , n73265 , n64994 );
and ( n73267 , n73262 , n73266 );
xor ( n73268 , n72899 , n72915 );
xor ( n73269 , n73268 , n72920 );
and ( n73270 , n73266 , n73269 );
and ( n73271 , n73262 , n73269 );
or ( n73272 , n73267 , n73270 , n73271 );
and ( n73273 , n70822 , n65183 );
and ( n73274 , n70832 , n65181 );
nor ( n73275 , n73273 , n73274 );
xnor ( n73276 , n73275 , n64994 );
and ( n73277 , n73272 , n73276 );
xor ( n73278 , n72923 , n72927 );
xor ( n73279 , n73278 , n72930 );
and ( n73280 , n73276 , n73279 );
and ( n73281 , n73272 , n73279 );
or ( n73282 , n73277 , n73280 , n73281 );
and ( n73283 , n70832 , n65183 );
and ( n73284 , n70766 , n65181 );
nor ( n73285 , n73283 , n73284 );
xnor ( n73286 , n73285 , n64994 );
and ( n73287 , n73282 , n73286 );
xor ( n73288 , n72933 , n72937 );
xor ( n73289 , n73288 , n72940 );
and ( n73290 , n73286 , n73289 );
and ( n73291 , n73282 , n73289 );
or ( n73292 , n73287 , n73290 , n73291 );
and ( n73293 , n70766 , n65183 );
and ( n73294 , n70266 , n65181 );
nor ( n73295 , n73293 , n73294 );
xnor ( n73296 , n73295 , n64994 );
and ( n73297 , n73292 , n73296 );
xor ( n73298 , n72943 , n72947 );
xor ( n73299 , n73298 , n72950 );
and ( n73300 , n73296 , n73299 );
and ( n73301 , n73292 , n73299 );
or ( n73302 , n73297 , n73300 , n73301 );
and ( n73303 , n69979 , n65550 );
and ( n73304 , n69573 , n65548 );
nor ( n73305 , n73303 , n73304 );
xnor ( n73306 , n73305 , n65313 );
and ( n73307 , n73302 , n73306 );
xor ( n73308 , n72987 , n72991 );
xor ( n73309 , n73308 , n72994 );
and ( n73310 , n73306 , n73309 );
and ( n73311 , n73302 , n73309 );
or ( n73312 , n73307 , n73310 , n73311 );
and ( n73313 , n70238 , n65550 );
and ( n73314 , n69985 , n65548 );
nor ( n73315 , n73313 , n73314 );
xnor ( n73316 , n73315 , n65313 );
and ( n73317 , n70266 , n65371 );
and ( n73318 , n70252 , n65369 );
nor ( n73319 , n73317 , n73318 );
xnor ( n73320 , n73319 , n65168 );
and ( n73321 , n73316 , n73320 );
xor ( n73322 , n73282 , n73286 );
xor ( n73323 , n73322 , n73289 );
and ( n73324 , n73320 , n73323 );
and ( n73325 , n73316 , n73323 );
or ( n73326 , n73321 , n73324 , n73325 );
and ( n73327 , n70252 , n65371 );
and ( n73328 , n70238 , n65369 );
nor ( n73329 , n73327 , n73328 );
xnor ( n73330 , n73329 , n65168 );
and ( n73331 , n73326 , n73330 );
xor ( n73332 , n73292 , n73296 );
xor ( n73333 , n73332 , n73299 );
and ( n73334 , n73330 , n73333 );
and ( n73335 , n73326 , n73333 );
or ( n73336 , n73331 , n73334 , n73335 );
and ( n73337 , n69566 , n65756 );
and ( n73338 , n69568 , n65754 );
nor ( n73339 , n73337 , n73338 );
xnor ( n73340 , n73339 , n65450 );
and ( n73341 , n73336 , n73340 );
xor ( n73342 , n73302 , n73306 );
xor ( n73343 , n73342 , n73309 );
and ( n73344 , n73340 , n73343 );
and ( n73345 , n73336 , n73343 );
or ( n73346 , n73341 , n73344 , n73345 );
and ( n73347 , n73312 , n73346 );
xor ( n73348 , n73195 , n73199 );
xor ( n73349 , n73348 , n73202 );
and ( n73350 , n73346 , n73349 );
and ( n73351 , n73312 , n73349 );
or ( n73352 , n73347 , n73350 , n73351 );
and ( n73353 , n68625 , n66241 );
and ( n73354 , n68444 , n66239 );
nor ( n73355 , n73353 , n73354 );
xnor ( n73356 , n73355 , n65876 );
and ( n73357 , n73352 , n73356 );
and ( n73358 , n69449 , n65756 );
and ( n73359 , n69095 , n65754 );
nor ( n73360 , n73358 , n73359 );
xnor ( n73361 , n73360 , n65450 );
and ( n73362 , n73356 , n73361 );
and ( n73363 , n73352 , n73361 );
or ( n73364 , n73357 , n73362 , n73363 );
and ( n73365 , n67873 , n66906 );
and ( n73366 , n67833 , n66904 );
nor ( n73367 , n73365 , n73366 );
xnor ( n73368 , n73367 , n66286 );
and ( n73369 , n73364 , n73368 );
xor ( n73370 , n73069 , n73073 );
xor ( n73371 , n73370 , n73076 );
and ( n73372 , n73368 , n73371 );
and ( n73373 , n73364 , n73371 );
or ( n73374 , n73369 , n73372 , n73373 );
and ( n73375 , n73227 , n73374 );
xor ( n73376 , n73079 , n73083 );
xor ( n73377 , n73376 , n73086 );
and ( n73378 , n73374 , n73377 );
and ( n73379 , n73227 , n73377 );
or ( n73380 , n73375 , n73378 , n73379 );
and ( n73381 , n67307 , n67160 );
and ( n73382 , n67302 , n67158 );
nor ( n73383 , n73381 , n73382 );
xnor ( n73384 , n73383 , n66514 );
and ( n73385 , n73380 , n73384 );
xor ( n73386 , n73089 , n73093 );
xor ( n73387 , n73386 , n73096 );
and ( n73388 , n73384 , n73387 );
and ( n73389 , n73380 , n73387 );
or ( n73390 , n73385 , n73388 , n73389 );
and ( n73391 , n66981 , n67498 );
and ( n73392 , n66786 , n67495 );
nor ( n73393 , n73391 , n73392 );
xnor ( n73394 , n73393 , n66511 );
and ( n73395 , n73390 , n73394 );
xor ( n73396 , n73099 , n73103 );
xor ( n73397 , n73396 , n73106 );
and ( n73398 , n73394 , n73397 );
and ( n73399 , n73390 , n73397 );
or ( n73400 , n73395 , n73398 , n73399 );
xor ( n73401 , n73171 , n73175 );
xor ( n73402 , n73401 , n73178 );
and ( n73403 , n73400 , n73402 );
xor ( n73404 , n73109 , n73113 );
xor ( n73405 , n73404 , n73116 );
and ( n73406 , n73402 , n73405 );
and ( n73407 , n73400 , n73405 );
or ( n73408 , n73403 , n73406 , n73407 );
xor ( n73409 , n73181 , n73183 );
xor ( n73410 , n73409 , n73186 );
and ( n73411 , n73408 , n73410 );
xor ( n73412 , n73408 , n73410 );
xor ( n73413 , n73400 , n73402 );
xor ( n73414 , n73413 , n73405 );
and ( n73415 , n69095 , n66016 );
and ( n73416 , n68873 , n66014 );
nor ( n73417 , n73415 , n73416 );
xnor ( n73418 , n73417 , n65650 );
and ( n73419 , n69568 , n65756 );
and ( n73420 , n69449 , n65754 );
nor ( n73421 , n73419 , n73420 );
xnor ( n73422 , n73421 , n65450 );
and ( n73423 , n73418 , n73422 );
xor ( n73424 , n73312 , n73346 );
xor ( n73425 , n73424 , n73349 );
and ( n73426 , n73422 , n73425 );
and ( n73427 , n73418 , n73425 );
or ( n73428 , n73423 , n73426 , n73427 );
and ( n73429 , n68439 , n66657 );
and ( n73430 , n68199 , n66655 );
nor ( n73431 , n73429 , n73430 );
xnor ( n73432 , n73431 , n66130 );
and ( n73433 , n73428 , n73432 );
xor ( n73434 , n73205 , n73209 );
xor ( n73435 , n73434 , n73212 );
and ( n73436 , n73432 , n73435 );
and ( n73437 , n73428 , n73435 );
or ( n73438 , n73433 , n73436 , n73437 );
and ( n73439 , n68199 , n66657 );
and ( n73440 , n68192 , n66655 );
nor ( n73441 , n73439 , n73440 );
xnor ( n73442 , n73441 , n66130 );
and ( n73443 , n73438 , n73442 );
xor ( n73444 , n73215 , n73219 );
xor ( n73445 , n73444 , n73224 );
and ( n73446 , n73442 , n73445 );
and ( n73447 , n73438 , n73445 );
or ( n73448 , n73443 , n73446 , n73447 );
and ( n73449 , n67302 , n67498 );
and ( n73450 , n67111 , n67495 );
nor ( n73451 , n73449 , n73450 );
xnor ( n73452 , n73451 , n66511 );
and ( n73453 , n73448 , n73452 );
and ( n73454 , n67548 , n67160 );
and ( n73455 , n67307 , n67158 );
nor ( n73456 , n73454 , n73455 );
xnor ( n73457 , n73456 , n66514 );
and ( n73458 , n73452 , n73457 );
and ( n73459 , n73448 , n73457 );
or ( n73460 , n73453 , n73458 , n73459 );
and ( n73461 , n67111 , n67498 );
and ( n73462 , n66981 , n67495 );
nor ( n73463 , n73461 , n73462 );
xnor ( n73464 , n73463 , n66511 );
and ( n73465 , n73460 , n73464 );
xor ( n73466 , n73151 , n73155 );
xor ( n73467 , n73466 , n73158 );
and ( n73468 , n73464 , n73467 );
and ( n73469 , n73460 , n73467 );
or ( n73470 , n73465 , n73468 , n73469 );
xor ( n73471 , n73390 , n73394 );
xor ( n73472 , n73471 , n73397 );
and ( n73473 , n73470 , n73472 );
xor ( n73474 , n73161 , n73165 );
xor ( n73475 , n73474 , n73168 );
and ( n73476 , n73472 , n73475 );
and ( n73477 , n73470 , n73475 );
or ( n73478 , n73473 , n73476 , n73477 );
and ( n73479 , n73414 , n73478 );
xor ( n73480 , n73414 , n73478 );
xor ( n73481 , n73470 , n73472 );
xor ( n73482 , n73481 , n73475 );
and ( n73483 , n69573 , n65756 );
and ( n73484 , n69566 , n65754 );
nor ( n73485 , n73483 , n73484 );
xnor ( n73486 , n73485 , n65450 );
and ( n73487 , n69985 , n65550 );
and ( n73488 , n69979 , n65548 );
nor ( n73489 , n73487 , n73488 );
xnor ( n73490 , n73489 , n65313 );
and ( n73491 , n73486 , n73490 );
xor ( n73492 , n73326 , n73330 );
xor ( n73493 , n73492 , n73333 );
and ( n73494 , n73490 , n73493 );
and ( n73495 , n73486 , n73493 );
or ( n73496 , n73491 , n73494 , n73495 );
and ( n73497 , n69449 , n66016 );
and ( n73498 , n69095 , n66014 );
nor ( n73499 , n73497 , n73498 );
xnor ( n73500 , n73499 , n65650 );
and ( n73501 , n73496 , n73500 );
xor ( n73502 , n73336 , n73340 );
xor ( n73503 , n73502 , n73343 );
and ( n73504 , n73500 , n73503 );
and ( n73505 , n73496 , n73503 );
or ( n73506 , n73501 , n73504 , n73505 );
and ( n73507 , n68444 , n66657 );
and ( n73508 , n68439 , n66655 );
nor ( n73509 , n73507 , n73508 );
xnor ( n73510 , n73509 , n66130 );
and ( n73511 , n73506 , n73510 );
and ( n73512 , n68837 , n66241 );
and ( n73513 , n68625 , n66239 );
nor ( n73514 , n73512 , n73513 );
xnor ( n73515 , n73514 , n65876 );
and ( n73516 , n73510 , n73515 );
and ( n73517 , n73506 , n73515 );
or ( n73518 , n73511 , n73516 , n73517 );
and ( n73519 , n67833 , n67160 );
and ( n73520 , n67727 , n67158 );
nor ( n73521 , n73519 , n73520 );
xnor ( n73522 , n73521 , n66514 );
and ( n73523 , n73518 , n73522 );
xor ( n73524 , n73352 , n73356 );
xor ( n73525 , n73524 , n73361 );
and ( n73526 , n73522 , n73525 );
and ( n73527 , n73518 , n73525 );
or ( n73528 , n73523 , n73526 , n73527 );
and ( n73529 , n67727 , n67160 );
and ( n73530 , n67548 , n67158 );
nor ( n73531 , n73529 , n73530 );
xnor ( n73532 , n73531 , n66514 );
and ( n73533 , n73528 , n73532 );
xor ( n73534 , n73364 , n73368 );
xor ( n73535 , n73534 , n73371 );
and ( n73536 , n73532 , n73535 );
and ( n73537 , n73528 , n73535 );
or ( n73538 , n73533 , n73536 , n73537 );
xor ( n73539 , n73141 , n73145 );
xor ( n73540 , n73539 , n73148 );
and ( n73541 , n73538 , n73540 );
xor ( n73542 , n73227 , n73374 );
xor ( n73543 , n73542 , n73377 );
and ( n73544 , n73540 , n73543 );
and ( n73545 , n73538 , n73543 );
or ( n73546 , n73541 , n73544 , n73545 );
xor ( n73547 , n73380 , n73384 );
xor ( n73548 , n73547 , n73387 );
and ( n73549 , n73546 , n73548 );
xor ( n73550 , n73460 , n73464 );
xor ( n73551 , n73550 , n73467 );
and ( n73552 , n73548 , n73551 );
and ( n73553 , n73546 , n73551 );
or ( n73554 , n73549 , n73552 , n73553 );
and ( n73555 , n73482 , n73554 );
xor ( n73556 , n73482 , n73554 );
xor ( n73557 , n73231 , n73235 );
and ( n73558 , n70781 , n65369 );
not ( n73559 , n73558 );
and ( n73560 , n73559 , n65168 );
and ( n73561 , n70781 , n65371 );
and ( n73562 , n70786 , n65369 );
nor ( n73563 , n73561 , n73562 );
xnor ( n73564 , n73563 , n65168 );
and ( n73565 , n73560 , n73564 );
and ( n73566 , n70786 , n65371 );
and ( n73567 , n70792 , n65369 );
nor ( n73568 , n73566 , n73567 );
xnor ( n73569 , n73568 , n65168 );
and ( n73570 , n73565 , n73569 );
and ( n73571 , n73569 , n73229 );
and ( n73572 , n73565 , n73229 );
or ( n73573 , n73570 , n73571 , n73572 );
and ( n73574 , n73557 , n73573 );
and ( n73575 , n70792 , n65371 );
and ( n73576 , n70802 , n65369 );
nor ( n73577 , n73575 , n73576 );
xnor ( n73578 , n73577 , n65168 );
and ( n73579 , n73573 , n73578 );
and ( n73580 , n73557 , n73578 );
or ( n73581 , n73574 , n73579 , n73580 );
and ( n73582 , n70802 , n65371 );
and ( n73583 , n70812 , n65369 );
nor ( n73584 , n73582 , n73583 );
xnor ( n73585 , n73584 , n65168 );
and ( n73586 , n73581 , n73585 );
xor ( n73587 , n73236 , n73240 );
xor ( n73588 , n73587 , n72900 );
and ( n73589 , n73585 , n73588 );
and ( n73590 , n73581 , n73588 );
or ( n73591 , n73586 , n73589 , n73590 );
and ( n73592 , n70812 , n65371 );
and ( n73593 , n70822 , n65369 );
nor ( n73594 , n73592 , n73593 );
xnor ( n73595 , n73594 , n65168 );
and ( n73596 , n73591 , n73595 );
xor ( n73597 , n73228 , n73244 );
xor ( n73598 , n73597 , n73249 );
and ( n73599 , n73595 , n73598 );
and ( n73600 , n73591 , n73598 );
or ( n73601 , n73596 , n73599 , n73600 );
and ( n73602 , n70822 , n65371 );
and ( n73603 , n70832 , n65369 );
nor ( n73604 , n73602 , n73603 );
xnor ( n73605 , n73604 , n65168 );
and ( n73606 , n73601 , n73605 );
xor ( n73607 , n73252 , n73256 );
xor ( n73608 , n73607 , n73259 );
and ( n73609 , n73605 , n73608 );
and ( n73610 , n73601 , n73608 );
or ( n73611 , n73606 , n73609 , n73610 );
and ( n73612 , n70832 , n65371 );
and ( n73613 , n70766 , n65369 );
nor ( n73614 , n73612 , n73613 );
xnor ( n73615 , n73614 , n65168 );
and ( n73616 , n73611 , n73615 );
xor ( n73617 , n73262 , n73266 );
xor ( n73618 , n73617 , n73269 );
and ( n73619 , n73615 , n73618 );
and ( n73620 , n73611 , n73618 );
or ( n73621 , n73616 , n73619 , n73620 );
and ( n73622 , n70766 , n65371 );
and ( n73623 , n70266 , n65369 );
nor ( n73624 , n73622 , n73623 );
xnor ( n73625 , n73624 , n65168 );
and ( n73626 , n73621 , n73625 );
xor ( n73627 , n73272 , n73276 );
xor ( n73628 , n73627 , n73279 );
and ( n73629 , n73625 , n73628 );
and ( n73630 , n73621 , n73628 );
or ( n73631 , n73626 , n73629 , n73630 );
and ( n73632 , n69979 , n65756 );
and ( n73633 , n69573 , n65754 );
nor ( n73634 , n73632 , n73633 );
xnor ( n73635 , n73634 , n65450 );
and ( n73636 , n73631 , n73635 );
xor ( n73637 , n73316 , n73320 );
xor ( n73638 , n73637 , n73323 );
and ( n73639 , n73635 , n73638 );
and ( n73640 , n73631 , n73638 );
or ( n73641 , n73636 , n73639 , n73640 );
and ( n73642 , n70238 , n65756 );
and ( n73643 , n69985 , n65754 );
nor ( n73644 , n73642 , n73643 );
xnor ( n73645 , n73644 , n65450 );
and ( n73646 , n70266 , n65550 );
and ( n73647 , n70252 , n65548 );
nor ( n73648 , n73646 , n73647 );
xnor ( n73649 , n73648 , n65313 );
and ( n73650 , n73645 , n73649 );
xor ( n73651 , n73611 , n73615 );
xor ( n73652 , n73651 , n73618 );
and ( n73653 , n73649 , n73652 );
and ( n73654 , n73645 , n73652 );
or ( n73655 , n73650 , n73653 , n73654 );
and ( n73656 , n70252 , n65550 );
and ( n73657 , n70238 , n65548 );
nor ( n73658 , n73656 , n73657 );
xnor ( n73659 , n73658 , n65313 );
and ( n73660 , n73655 , n73659 );
xor ( n73661 , n73621 , n73625 );
xor ( n73662 , n73661 , n73628 );
and ( n73663 , n73659 , n73662 );
and ( n73664 , n73655 , n73662 );
or ( n73665 , n73660 , n73663 , n73664 );
and ( n73666 , n69566 , n66016 );
and ( n73667 , n69568 , n66014 );
nor ( n73668 , n73666 , n73667 );
xnor ( n73669 , n73668 , n65650 );
and ( n73670 , n73665 , n73669 );
xor ( n73671 , n73631 , n73635 );
xor ( n73672 , n73671 , n73638 );
and ( n73673 , n73669 , n73672 );
and ( n73674 , n73665 , n73672 );
or ( n73675 , n73670 , n73673 , n73674 );
and ( n73676 , n73641 , n73675 );
xor ( n73677 , n73486 , n73490 );
xor ( n73678 , n73677 , n73493 );
and ( n73679 , n73675 , n73678 );
and ( n73680 , n73641 , n73678 );
or ( n73681 , n73676 , n73679 , n73680 );
and ( n73682 , n68625 , n66657 );
and ( n73683 , n68444 , n66655 );
nor ( n73684 , n73682 , n73683 );
xnor ( n73685 , n73684 , n66130 );
and ( n73686 , n73681 , n73685 );
and ( n73687 , n68873 , n66241 );
and ( n73688 , n68837 , n66239 );
nor ( n73689 , n73687 , n73688 );
xnor ( n73690 , n73689 , n65876 );
and ( n73691 , n73685 , n73690 );
and ( n73692 , n73681 , n73690 );
or ( n73693 , n73686 , n73691 , n73692 );
and ( n73694 , n67873 , n67160 );
and ( n73695 , n67833 , n67158 );
nor ( n73696 , n73694 , n73695 );
xnor ( n73697 , n73696 , n66514 );
and ( n73698 , n73693 , n73697 );
xor ( n73699 , n73418 , n73422 );
xor ( n73700 , n73699 , n73425 );
and ( n73701 , n73697 , n73700 );
and ( n73702 , n73693 , n73700 );
or ( n73703 , n73698 , n73701 , n73702 );
and ( n73704 , n68192 , n66906 );
and ( n73705 , n67873 , n66904 );
nor ( n73706 , n73704 , n73705 );
xnor ( n73707 , n73706 , n66286 );
and ( n73708 , n73703 , n73707 );
xor ( n73709 , n73428 , n73432 );
xor ( n73710 , n73709 , n73435 );
and ( n73711 , n73707 , n73710 );
and ( n73712 , n73703 , n73710 );
or ( n73713 , n73708 , n73711 , n73712 );
and ( n73714 , n67307 , n67498 );
and ( n73715 , n67302 , n67495 );
nor ( n73716 , n73714 , n73715 );
xnor ( n73717 , n73716 , n66511 );
and ( n73718 , n73713 , n73717 );
xor ( n73719 , n73438 , n73442 );
xor ( n73720 , n73719 , n73445 );
and ( n73721 , n73717 , n73720 );
and ( n73722 , n73713 , n73720 );
or ( n73723 , n73718 , n73721 , n73722 );
xor ( n73724 , n73448 , n73452 );
xor ( n73725 , n73724 , n73457 );
and ( n73726 , n73723 , n73725 );
xor ( n73727 , n73538 , n73540 );
xor ( n73728 , n73727 , n73543 );
and ( n73729 , n73725 , n73728 );
and ( n73730 , n73723 , n73728 );
or ( n73731 , n73726 , n73729 , n73730 );
xor ( n73732 , n73546 , n73548 );
xor ( n73733 , n73732 , n73551 );
and ( n73734 , n73731 , n73733 );
xor ( n73735 , n73731 , n73733 );
xor ( n73736 , n73723 , n73725 );
xor ( n73737 , n73736 , n73728 );
and ( n73738 , n69095 , n66241 );
and ( n73739 , n68873 , n66239 );
nor ( n73740 , n73738 , n73739 );
xnor ( n73741 , n73740 , n65876 );
and ( n73742 , n69568 , n66016 );
and ( n73743 , n69449 , n66014 );
nor ( n73744 , n73742 , n73743 );
xnor ( n73745 , n73744 , n65650 );
and ( n73746 , n73741 , n73745 );
xor ( n73747 , n73641 , n73675 );
xor ( n73748 , n73747 , n73678 );
and ( n73749 , n73745 , n73748 );
and ( n73750 , n73741 , n73748 );
or ( n73751 , n73746 , n73749 , n73750 );
and ( n73752 , n68439 , n66906 );
and ( n73753 , n68199 , n66904 );
nor ( n73754 , n73752 , n73753 );
xnor ( n73755 , n73754 , n66286 );
and ( n73756 , n73751 , n73755 );
xor ( n73757 , n73496 , n73500 );
xor ( n73758 , n73757 , n73503 );
and ( n73759 , n73755 , n73758 );
and ( n73760 , n73751 , n73758 );
or ( n73761 , n73756 , n73759 , n73760 );
and ( n73762 , n68199 , n66906 );
and ( n73763 , n68192 , n66904 );
nor ( n73764 , n73762 , n73763 );
xnor ( n73765 , n73764 , n66286 );
and ( n73766 , n73761 , n73765 );
xor ( n73767 , n73506 , n73510 );
xor ( n73768 , n73767 , n73515 );
and ( n73769 , n73765 , n73768 );
and ( n73770 , n73761 , n73768 );
or ( n73771 , n73766 , n73769 , n73770 );
and ( n73772 , n67548 , n67498 );
and ( n73773 , n67307 , n67495 );
nor ( n73774 , n73772 , n73773 );
xnor ( n73775 , n73774 , n66511 );
and ( n73776 , n73771 , n73775 );
xor ( n73777 , n73518 , n73522 );
xor ( n73778 , n73777 , n73525 );
and ( n73779 , n73775 , n73778 );
and ( n73780 , n73771 , n73778 );
or ( n73781 , n73776 , n73779 , n73780 );
xor ( n73782 , n73713 , n73717 );
xor ( n73783 , n73782 , n73720 );
and ( n73784 , n73781 , n73783 );
xor ( n73785 , n73528 , n73532 );
xor ( n73786 , n73785 , n73535 );
and ( n73787 , n73783 , n73786 );
and ( n73788 , n73781 , n73786 );
or ( n73789 , n73784 , n73787 , n73788 );
and ( n73790 , n73737 , n73789 );
xor ( n73791 , n73737 , n73789 );
xor ( n73792 , n73781 , n73783 );
xor ( n73793 , n73792 , n73786 );
and ( n73794 , n67833 , n67498 );
and ( n73795 , n67727 , n67495 );
nor ( n73796 , n73794 , n73795 );
xnor ( n73797 , n73796 , n66511 );
and ( n73798 , n68192 , n67160 );
and ( n73799 , n67873 , n67158 );
nor ( n73800 , n73798 , n73799 );
xnor ( n73801 , n73800 , n66514 );
and ( n73802 , n73797 , n73801 );
xor ( n73803 , n73681 , n73685 );
xor ( n73804 , n73803 , n73690 );
and ( n73805 , n73801 , n73804 );
and ( n73806 , n73797 , n73804 );
or ( n73807 , n73802 , n73805 , n73806 );
and ( n73808 , n67727 , n67498 );
and ( n73809 , n67548 , n67495 );
nor ( n73810 , n73808 , n73809 );
xnor ( n73811 , n73810 , n66511 );
and ( n73812 , n73807 , n73811 );
xor ( n73813 , n73693 , n73697 );
xor ( n73814 , n73813 , n73700 );
and ( n73815 , n73811 , n73814 );
and ( n73816 , n73807 , n73814 );
or ( n73817 , n73812 , n73815 , n73816 );
xor ( n73818 , n73771 , n73775 );
xor ( n73819 , n73818 , n73778 );
and ( n73820 , n73817 , n73819 );
xor ( n73821 , n73703 , n73707 );
xor ( n73822 , n73821 , n73710 );
and ( n73823 , n73819 , n73822 );
and ( n73824 , n73817 , n73822 );
or ( n73825 , n73820 , n73823 , n73824 );
and ( n73826 , n73793 , n73825 );
xor ( n73827 , n73793 , n73825 );
xor ( n73828 , n73817 , n73819 );
xor ( n73829 , n73828 , n73822 );
and ( n73830 , n69573 , n66016 );
and ( n73831 , n69566 , n66014 );
nor ( n73832 , n73830 , n73831 );
xnor ( n73833 , n73832 , n65650 );
and ( n73834 , n69985 , n65756 );
and ( n73835 , n69979 , n65754 );
nor ( n73836 , n73834 , n73835 );
xnor ( n73837 , n73836 , n65450 );
and ( n73838 , n73833 , n73837 );
xor ( n73839 , n73655 , n73659 );
xor ( n73840 , n73839 , n73662 );
and ( n73841 , n73837 , n73840 );
and ( n73842 , n73833 , n73840 );
or ( n73843 , n73838 , n73841 , n73842 );
xor ( n73844 , n73560 , n73564 );
and ( n73845 , n70781 , n65548 );
not ( n73846 , n73845 );
and ( n73847 , n73846 , n65313 );
and ( n73848 , n70781 , n65550 );
and ( n73849 , n70786 , n65548 );
nor ( n73850 , n73848 , n73849 );
xnor ( n73851 , n73850 , n65313 );
and ( n73852 , n73847 , n73851 );
and ( n73853 , n70786 , n65550 );
and ( n73854 , n70792 , n65548 );
nor ( n73855 , n73853 , n73854 );
xnor ( n73856 , n73855 , n65313 );
and ( n73857 , n73852 , n73856 );
and ( n73858 , n73856 , n73558 );
and ( n73859 , n73852 , n73558 );
or ( n73860 , n73857 , n73858 , n73859 );
and ( n73861 , n73844 , n73860 );
and ( n73862 , n70792 , n65550 );
and ( n73863 , n70802 , n65548 );
nor ( n73864 , n73862 , n73863 );
xnor ( n73865 , n73864 , n65313 );
and ( n73866 , n73860 , n73865 );
and ( n73867 , n73844 , n73865 );
or ( n73868 , n73861 , n73866 , n73867 );
and ( n73869 , n70802 , n65550 );
and ( n73870 , n70812 , n65548 );
nor ( n73871 , n73869 , n73870 );
xnor ( n73872 , n73871 , n65313 );
and ( n73873 , n73868 , n73872 );
xor ( n73874 , n73565 , n73569 );
xor ( n73875 , n73874 , n73229 );
and ( n73876 , n73872 , n73875 );
and ( n73877 , n73868 , n73875 );
or ( n73878 , n73873 , n73876 , n73877 );
and ( n73879 , n70812 , n65550 );
and ( n73880 , n70822 , n65548 );
nor ( n73881 , n73879 , n73880 );
xnor ( n73882 , n73881 , n65313 );
and ( n73883 , n73878 , n73882 );
xor ( n73884 , n73557 , n73573 );
xor ( n73885 , n73884 , n73578 );
and ( n73886 , n73882 , n73885 );
and ( n73887 , n73878 , n73885 );
or ( n73888 , n73883 , n73886 , n73887 );
and ( n73889 , n70822 , n65550 );
and ( n73890 , n70832 , n65548 );
nor ( n73891 , n73889 , n73890 );
xnor ( n73892 , n73891 , n65313 );
and ( n73893 , n73888 , n73892 );
xor ( n73894 , n73581 , n73585 );
xor ( n73895 , n73894 , n73588 );
and ( n73896 , n73892 , n73895 );
and ( n73897 , n73888 , n73895 );
or ( n73898 , n73893 , n73896 , n73897 );
and ( n73899 , n70832 , n65550 );
and ( n73900 , n70766 , n65548 );
nor ( n73901 , n73899 , n73900 );
xnor ( n73902 , n73901 , n65313 );
and ( n73903 , n73898 , n73902 );
xor ( n73904 , n73591 , n73595 );
xor ( n73905 , n73904 , n73598 );
and ( n73906 , n73902 , n73905 );
and ( n73907 , n73898 , n73905 );
or ( n73908 , n73903 , n73906 , n73907 );
and ( n73909 , n70766 , n65550 );
and ( n73910 , n70266 , n65548 );
nor ( n73911 , n73909 , n73910 );
xnor ( n73912 , n73911 , n65313 );
and ( n73913 , n73908 , n73912 );
xor ( n73914 , n73601 , n73605 );
xor ( n73915 , n73914 , n73608 );
and ( n73916 , n73912 , n73915 );
and ( n73917 , n73908 , n73915 );
or ( n73918 , n73913 , n73916 , n73917 );
and ( n73919 , n69979 , n66016 );
and ( n73920 , n69573 , n66014 );
nor ( n73921 , n73919 , n73920 );
xnor ( n73922 , n73921 , n65650 );
and ( n73923 , n73918 , n73922 );
xor ( n73924 , n73645 , n73649 );
xor ( n73925 , n73924 , n73652 );
and ( n73926 , n73922 , n73925 );
and ( n73927 , n73918 , n73925 );
or ( n73928 , n73923 , n73926 , n73927 );
and ( n73929 , n69985 , n66016 );
and ( n73930 , n69979 , n66014 );
nor ( n73931 , n73929 , n73930 );
xnor ( n73932 , n73931 , n65650 );
and ( n73933 , n70252 , n65756 );
and ( n73934 , n70238 , n65754 );
nor ( n73935 , n73933 , n73934 );
xnor ( n73936 , n73935 , n65450 );
and ( n73937 , n73932 , n73936 );
xor ( n73938 , n73908 , n73912 );
xor ( n73939 , n73938 , n73915 );
and ( n73940 , n73936 , n73939 );
and ( n73941 , n73932 , n73939 );
or ( n73942 , n73937 , n73940 , n73941 );
and ( n73943 , n69566 , n66241 );
and ( n73944 , n69568 , n66239 );
nor ( n73945 , n73943 , n73944 );
xnor ( n73946 , n73945 , n65876 );
and ( n73947 , n73942 , n73946 );
xor ( n73948 , n73918 , n73922 );
xor ( n73949 , n73948 , n73925 );
and ( n73950 , n73946 , n73949 );
and ( n73951 , n73942 , n73949 );
or ( n73952 , n73947 , n73950 , n73951 );
and ( n73953 , n73928 , n73952 );
xor ( n73954 , n73833 , n73837 );
xor ( n73955 , n73954 , n73840 );
and ( n73956 , n73952 , n73955 );
and ( n73957 , n73928 , n73955 );
or ( n73958 , n73953 , n73956 , n73957 );
and ( n73959 , n73843 , n73958 );
xor ( n73960 , n73665 , n73669 );
xor ( n73961 , n73960 , n73672 );
and ( n73962 , n73958 , n73961 );
and ( n73963 , n73843 , n73961 );
or ( n73964 , n73959 , n73962 , n73963 );
and ( n73965 , n68444 , n66906 );
and ( n73966 , n68439 , n66904 );
nor ( n73967 , n73965 , n73966 );
xnor ( n73968 , n73967 , n66286 );
and ( n73969 , n73964 , n73968 );
and ( n73970 , n68837 , n66657 );
and ( n73971 , n68625 , n66655 );
nor ( n73972 , n73970 , n73971 );
xnor ( n73973 , n73972 , n66130 );
and ( n73974 , n73968 , n73973 );
and ( n73975 , n73964 , n73973 );
or ( n73976 , n73969 , n73974 , n73975 );
and ( n73977 , n68625 , n66906 );
and ( n73978 , n68444 , n66904 );
nor ( n73979 , n73977 , n73978 );
xnor ( n73980 , n73979 , n66286 );
and ( n73981 , n68873 , n66657 );
and ( n73982 , n68837 , n66655 );
nor ( n73983 , n73981 , n73982 );
xnor ( n73984 , n73983 , n66130 );
and ( n73985 , n73980 , n73984 );
and ( n73986 , n69449 , n66241 );
and ( n73987 , n69095 , n66239 );
nor ( n73988 , n73986 , n73987 );
xnor ( n73989 , n73988 , n65876 );
and ( n73990 , n73984 , n73989 );
and ( n73991 , n73980 , n73989 );
or ( n73992 , n73985 , n73990 , n73991 );
xor ( n73993 , n73964 , n73968 );
xor ( n73994 , n73993 , n73973 );
and ( n73995 , n73992 , n73994 );
xor ( n73996 , n73741 , n73745 );
xor ( n73997 , n73996 , n73748 );
and ( n73998 , n73994 , n73997 );
and ( n73999 , n73992 , n73997 );
or ( n74000 , n73995 , n73998 , n73999 );
and ( n74001 , n73976 , n74000 );
xor ( n74002 , n73751 , n73755 );
xor ( n74003 , n74002 , n73758 );
and ( n74004 , n74000 , n74003 );
and ( n74005 , n73976 , n74003 );
or ( n74006 , n74001 , n74004 , n74005 );
xor ( n74007 , n73761 , n73765 );
xor ( n74008 , n74007 , n73768 );
and ( n74009 , n74006 , n74008 );
xor ( n74010 , n73807 , n73811 );
xor ( n74011 , n74010 , n73814 );
and ( n74012 , n74008 , n74011 );
and ( n74013 , n74006 , n74011 );
or ( n74014 , n74009 , n74012 , n74013 );
and ( n74015 , n73829 , n74014 );
xor ( n74016 , n73829 , n74014 );
xor ( n74017 , n74006 , n74008 );
xor ( n74018 , n74017 , n74011 );
and ( n74019 , n69095 , n66657 );
and ( n74020 , n68873 , n66655 );
nor ( n74021 , n74019 , n74020 );
xnor ( n74022 , n74021 , n66130 );
and ( n74023 , n69568 , n66241 );
and ( n74024 , n69449 , n66239 );
nor ( n74025 , n74023 , n74024 );
xnor ( n74026 , n74025 , n65876 );
and ( n74027 , n74022 , n74026 );
xor ( n74028 , n73928 , n73952 );
xor ( n74029 , n74028 , n73955 );
and ( n74030 , n74026 , n74029 );
and ( n74031 , n74022 , n74029 );
or ( n74032 , n74027 , n74030 , n74031 );
and ( n74033 , n68439 , n67160 );
and ( n74034 , n68199 , n67158 );
nor ( n74035 , n74033 , n74034 );
xnor ( n74036 , n74035 , n66514 );
and ( n74037 , n74032 , n74036 );
xor ( n74038 , n73843 , n73958 );
xor ( n74039 , n74038 , n73961 );
and ( n74040 , n74036 , n74039 );
and ( n74041 , n74032 , n74039 );
or ( n74042 , n74037 , n74040 , n74041 );
and ( n74043 , n67873 , n67498 );
and ( n74044 , n67833 , n67495 );
nor ( n74045 , n74043 , n74044 );
xnor ( n74046 , n74045 , n66511 );
and ( n74047 , n74042 , n74046 );
and ( n74048 , n68199 , n67160 );
and ( n74049 , n68192 , n67158 );
nor ( n74050 , n74048 , n74049 );
xnor ( n74051 , n74050 , n66514 );
and ( n74052 , n74046 , n74051 );
and ( n74053 , n74042 , n74051 );
or ( n74054 , n74047 , n74052 , n74053 );
xor ( n74055 , n73797 , n73801 );
xor ( n74056 , n74055 , n73804 );
and ( n74057 , n74054 , n74056 );
xor ( n74058 , n73976 , n74000 );
xor ( n74059 , n74058 , n74003 );
and ( n74060 , n74056 , n74059 );
and ( n74061 , n74054 , n74059 );
or ( n74062 , n74057 , n74060 , n74061 );
and ( n74063 , n74018 , n74062 );
xor ( n74064 , n74018 , n74062 );
and ( n74065 , n70238 , n66016 );
and ( n74066 , n69985 , n66014 );
nor ( n74067 , n74065 , n74066 );
xnor ( n74068 , n74067 , n65650 );
and ( n74069 , n70266 , n65756 );
and ( n74070 , n70252 , n65754 );
nor ( n74071 , n74069 , n74070 );
xnor ( n74072 , n74071 , n65450 );
and ( n74073 , n74068 , n74072 );
xor ( n74074 , n73898 , n73902 );
xor ( n74075 , n74074 , n73905 );
and ( n74076 , n74072 , n74075 );
and ( n74077 , n74068 , n74075 );
or ( n74078 , n74073 , n74076 , n74077 );
and ( n74079 , n69573 , n66241 );
and ( n74080 , n69566 , n66239 );
nor ( n74081 , n74079 , n74080 );
xnor ( n74082 , n74081 , n65876 );
and ( n74083 , n74078 , n74082 );
xor ( n74084 , n73932 , n73936 );
xor ( n74085 , n74084 , n73939 );
and ( n74086 , n74082 , n74085 );
and ( n74087 , n74078 , n74085 );
or ( n74088 , n74083 , n74086 , n74087 );
and ( n74089 , n69449 , n66657 );
and ( n74090 , n69095 , n66655 );
nor ( n74091 , n74089 , n74090 );
xnor ( n74092 , n74091 , n66130 );
and ( n74093 , n74088 , n74092 );
xor ( n74094 , n73942 , n73946 );
xor ( n74095 , n74094 , n73949 );
and ( n74096 , n74092 , n74095 );
and ( n74097 , n74088 , n74095 );
or ( n74098 , n74093 , n74096 , n74097 );
and ( n74099 , n68444 , n67160 );
and ( n74100 , n68439 , n67158 );
nor ( n74101 , n74099 , n74100 );
xnor ( n74102 , n74101 , n66514 );
and ( n74103 , n74098 , n74102 );
and ( n74104 , n68837 , n66906 );
and ( n74105 , n68625 , n66904 );
nor ( n74106 , n74104 , n74105 );
xnor ( n74107 , n74106 , n66286 );
and ( n74108 , n74102 , n74107 );
and ( n74109 , n74098 , n74107 );
or ( n74110 , n74103 , n74108 , n74109 );
and ( n74111 , n68192 , n67498 );
and ( n74112 , n67873 , n67495 );
nor ( n74113 , n74111 , n74112 );
xnor ( n74114 , n74113 , n66511 );
and ( n74115 , n74110 , n74114 );
xor ( n74116 , n73980 , n73984 );
xor ( n74117 , n74116 , n73989 );
and ( n74118 , n74114 , n74117 );
and ( n74119 , n74110 , n74117 );
or ( n74120 , n74115 , n74118 , n74119 );
xor ( n74121 , n74042 , n74046 );
xor ( n74122 , n74121 , n74051 );
and ( n74123 , n74120 , n74122 );
xor ( n74124 , n73992 , n73994 );
xor ( n74125 , n74124 , n73997 );
and ( n74126 , n74122 , n74125 );
and ( n74127 , n74120 , n74125 );
or ( n74128 , n74123 , n74126 , n74127 );
xor ( n74129 , n74054 , n74056 );
xor ( n74130 , n74129 , n74059 );
and ( n74131 , n74128 , n74130 );
xor ( n74132 , n74128 , n74130 );
xor ( n74133 , n73847 , n73851 );
and ( n74134 , n70781 , n65754 );
not ( n74135 , n74134 );
and ( n74136 , n74135 , n65450 );
and ( n74137 , n70781 , n65756 );
and ( n74138 , n70786 , n65754 );
nor ( n74139 , n74137 , n74138 );
xnor ( n74140 , n74139 , n65450 );
and ( n74141 , n74136 , n74140 );
and ( n74142 , n70786 , n65756 );
and ( n74143 , n70792 , n65754 );
nor ( n74144 , n74142 , n74143 );
xnor ( n74145 , n74144 , n65450 );
and ( n74146 , n74141 , n74145 );
and ( n74147 , n74145 , n73845 );
and ( n74148 , n74141 , n73845 );
or ( n74149 , n74146 , n74147 , n74148 );
and ( n74150 , n74133 , n74149 );
and ( n74151 , n70792 , n65756 );
and ( n74152 , n70802 , n65754 );
nor ( n74153 , n74151 , n74152 );
xnor ( n74154 , n74153 , n65450 );
and ( n74155 , n74149 , n74154 );
and ( n74156 , n74133 , n74154 );
or ( n74157 , n74150 , n74155 , n74156 );
and ( n74158 , n70802 , n65756 );
and ( n74159 , n70812 , n65754 );
nor ( n74160 , n74158 , n74159 );
xnor ( n74161 , n74160 , n65450 );
and ( n74162 , n74157 , n74161 );
xor ( n74163 , n73852 , n73856 );
xor ( n74164 , n74163 , n73558 );
and ( n74165 , n74161 , n74164 );
and ( n74166 , n74157 , n74164 );
or ( n74167 , n74162 , n74165 , n74166 );
and ( n74168 , n70812 , n65756 );
and ( n74169 , n70822 , n65754 );
nor ( n74170 , n74168 , n74169 );
xnor ( n74171 , n74170 , n65450 );
and ( n74172 , n74167 , n74171 );
xor ( n74173 , n73844 , n73860 );
xor ( n74174 , n74173 , n73865 );
and ( n74175 , n74171 , n74174 );
and ( n74176 , n74167 , n74174 );
or ( n74177 , n74172 , n74175 , n74176 );
and ( n74178 , n70822 , n65756 );
and ( n74179 , n70832 , n65754 );
nor ( n74180 , n74178 , n74179 );
xnor ( n74181 , n74180 , n65450 );
and ( n74182 , n74177 , n74181 );
xor ( n74183 , n73868 , n73872 );
xor ( n74184 , n74183 , n73875 );
and ( n74185 , n74181 , n74184 );
and ( n74186 , n74177 , n74184 );
or ( n74187 , n74182 , n74185 , n74186 );
and ( n74188 , n70832 , n65756 );
and ( n74189 , n70766 , n65754 );
nor ( n74190 , n74188 , n74189 );
xnor ( n74191 , n74190 , n65450 );
and ( n74192 , n74187 , n74191 );
xor ( n74193 , n73878 , n73882 );
xor ( n74194 , n74193 , n73885 );
and ( n74195 , n74191 , n74194 );
and ( n74196 , n74187 , n74194 );
or ( n74197 , n74192 , n74195 , n74196 );
and ( n74198 , n70766 , n65756 );
and ( n74199 , n70266 , n65754 );
nor ( n74200 , n74198 , n74199 );
xnor ( n74201 , n74200 , n65450 );
and ( n74202 , n74197 , n74201 );
xor ( n74203 , n73888 , n73892 );
xor ( n74204 , n74203 , n73895 );
and ( n74205 , n74201 , n74204 );
and ( n74206 , n74197 , n74204 );
or ( n74207 , n74202 , n74205 , n74206 );
and ( n74208 , n69979 , n66241 );
and ( n74209 , n69573 , n66239 );
nor ( n74210 , n74208 , n74209 );
xnor ( n74211 , n74210 , n65876 );
and ( n74212 , n74207 , n74211 );
xor ( n74213 , n74068 , n74072 );
xor ( n74214 , n74213 , n74075 );
and ( n74215 , n74211 , n74214 );
and ( n74216 , n74207 , n74214 );
or ( n74217 , n74212 , n74215 , n74216 );
and ( n74218 , n70238 , n66241 );
and ( n74219 , n69985 , n66239 );
nor ( n74220 , n74218 , n74219 );
xnor ( n74221 , n74220 , n65876 );
and ( n74222 , n70266 , n66016 );
and ( n74223 , n70252 , n66014 );
nor ( n74224 , n74222 , n74223 );
xnor ( n74225 , n74224 , n65650 );
and ( n74226 , n74221 , n74225 );
xor ( n74227 , n74187 , n74191 );
xor ( n74228 , n74227 , n74194 );
and ( n74229 , n74225 , n74228 );
and ( n74230 , n74221 , n74228 );
or ( n74231 , n74226 , n74229 , n74230 );
and ( n74232 , n70252 , n66016 );
and ( n74233 , n70238 , n66014 );
nor ( n74234 , n74232 , n74233 );
xnor ( n74235 , n74234 , n65650 );
and ( n74236 , n74231 , n74235 );
xor ( n74237 , n74197 , n74201 );
xor ( n74238 , n74237 , n74204 );
and ( n74239 , n74235 , n74238 );
and ( n74240 , n74231 , n74238 );
or ( n74241 , n74236 , n74239 , n74240 );
and ( n74242 , n69566 , n66657 );
and ( n74243 , n69568 , n66655 );
nor ( n74244 , n74242 , n74243 );
xnor ( n74245 , n74244 , n66130 );
and ( n74246 , n74241 , n74245 );
xor ( n74247 , n74207 , n74211 );
xor ( n74248 , n74247 , n74214 );
and ( n74249 , n74245 , n74248 );
and ( n74250 , n74241 , n74248 );
or ( n74251 , n74246 , n74249 , n74250 );
and ( n74252 , n74217 , n74251 );
xor ( n74253 , n74078 , n74082 );
xor ( n74254 , n74253 , n74085 );
and ( n74255 , n74251 , n74254 );
and ( n74256 , n74217 , n74254 );
or ( n74257 , n74252 , n74255 , n74256 );
and ( n74258 , n68625 , n67160 );
and ( n74259 , n68444 , n67158 );
nor ( n74260 , n74258 , n74259 );
xnor ( n74261 , n74260 , n66514 );
and ( n74262 , n74257 , n74261 );
and ( n74263 , n68873 , n66906 );
and ( n74264 , n68837 , n66904 );
nor ( n74265 , n74263 , n74264 );
xnor ( n74266 , n74265 , n66286 );
and ( n74267 , n74261 , n74266 );
and ( n74268 , n74257 , n74266 );
or ( n74269 , n74262 , n74267 , n74268 );
and ( n74270 , n68199 , n67498 );
and ( n74271 , n68192 , n67495 );
nor ( n74272 , n74270 , n74271 );
xnor ( n74273 , n74272 , n66511 );
and ( n74274 , n74269 , n74273 );
xor ( n74275 , n74022 , n74026 );
xor ( n74276 , n74275 , n74029 );
and ( n74277 , n74273 , n74276 );
and ( n74278 , n74269 , n74276 );
or ( n74279 , n74274 , n74277 , n74278 );
xor ( n74280 , n74110 , n74114 );
xor ( n74281 , n74280 , n74117 );
and ( n74282 , n74279 , n74281 );
xor ( n74283 , n74032 , n74036 );
xor ( n74284 , n74283 , n74039 );
and ( n74285 , n74281 , n74284 );
and ( n74286 , n74279 , n74284 );
or ( n74287 , n74282 , n74285 , n74286 );
xor ( n74288 , n74120 , n74122 );
xor ( n74289 , n74288 , n74125 );
and ( n74290 , n74287 , n74289 );
xor ( n74291 , n74287 , n74289 );
xor ( n74292 , n74279 , n74281 );
xor ( n74293 , n74292 , n74284 );
and ( n74294 , n69095 , n66906 );
and ( n74295 , n68873 , n66904 );
nor ( n74296 , n74294 , n74295 );
xnor ( n74297 , n74296 , n66286 );
and ( n74298 , n69568 , n66657 );
and ( n74299 , n69449 , n66655 );
nor ( n74300 , n74298 , n74299 );
xnor ( n74301 , n74300 , n66130 );
and ( n74302 , n74297 , n74301 );
xor ( n74303 , n74217 , n74251 );
xor ( n74304 , n74303 , n74254 );
and ( n74305 , n74301 , n74304 );
and ( n74306 , n74297 , n74304 );
or ( n74307 , n74302 , n74305 , n74306 );
and ( n74308 , n68439 , n67498 );
and ( n74309 , n68199 , n67495 );
nor ( n74310 , n74308 , n74309 );
xnor ( n74311 , n74310 , n66511 );
and ( n74312 , n74307 , n74311 );
xor ( n74313 , n74088 , n74092 );
xor ( n74314 , n74313 , n74095 );
and ( n74315 , n74311 , n74314 );
and ( n74316 , n74307 , n74314 );
or ( n74317 , n74312 , n74315 , n74316 );
xor ( n74318 , n74098 , n74102 );
xor ( n74319 , n74318 , n74107 );
and ( n74320 , n74317 , n74319 );
xor ( n74321 , n74269 , n74273 );
xor ( n74322 , n74321 , n74276 );
and ( n74323 , n74319 , n74322 );
and ( n74324 , n74317 , n74322 );
or ( n74325 , n74320 , n74323 , n74324 );
and ( n74326 , n74293 , n74325 );
xor ( n74327 , n74293 , n74325 );
xor ( n74328 , n74317 , n74319 );
xor ( n74329 , n74328 , n74322 );
and ( n74330 , n69573 , n66657 );
and ( n74331 , n69566 , n66655 );
nor ( n74332 , n74330 , n74331 );
xnor ( n74333 , n74332 , n66130 );
and ( n74334 , n69985 , n66241 );
and ( n74335 , n69979 , n66239 );
nor ( n74336 , n74334 , n74335 );
xnor ( n74337 , n74336 , n65876 );
and ( n74338 , n74333 , n74337 );
xor ( n74339 , n74231 , n74235 );
xor ( n74340 , n74339 , n74238 );
and ( n74341 , n74337 , n74340 );
and ( n74342 , n74333 , n74340 );
or ( n74343 , n74338 , n74341 , n74342 );
and ( n74344 , n68873 , n67160 );
and ( n74345 , n68837 , n67158 );
nor ( n74346 , n74344 , n74345 );
xnor ( n74347 , n74346 , n66514 );
and ( n74348 , n74343 , n74347 );
xor ( n74349 , n74241 , n74245 );
xor ( n74350 , n74349 , n74248 );
and ( n74351 , n74347 , n74350 );
and ( n74352 , n74343 , n74350 );
or ( n74353 , n74348 , n74351 , n74352 );
and ( n74354 , n68444 , n67498 );
and ( n74355 , n68439 , n67495 );
nor ( n74356 , n74354 , n74355 );
xnor ( n74357 , n74356 , n66511 );
and ( n74358 , n74353 , n74357 );
and ( n74359 , n68837 , n67160 );
and ( n74360 , n68625 , n67158 );
nor ( n74361 , n74359 , n74360 );
xnor ( n74362 , n74361 , n66514 );
and ( n74363 , n74357 , n74362 );
and ( n74364 , n74353 , n74362 );
or ( n74365 , n74358 , n74363 , n74364 );
xor ( n74366 , n74257 , n74261 );
xor ( n74367 , n74366 , n74266 );
and ( n74368 , n74365 , n74367 );
xor ( n74369 , n74307 , n74311 );
xor ( n74370 , n74369 , n74314 );
and ( n74371 , n74367 , n74370 );
and ( n74372 , n74365 , n74370 );
or ( n74373 , n74368 , n74371 , n74372 );
and ( n74374 , n74329 , n74373 );
xor ( n74375 , n74329 , n74373 );
xor ( n74376 , n74136 , n74140 );
and ( n74377 , n70781 , n66014 );
not ( n74378 , n74377 );
and ( n74379 , n74378 , n65650 );
and ( n74380 , n70781 , n66016 );
and ( n74381 , n70786 , n66014 );
nor ( n74382 , n74380 , n74381 );
xnor ( n74383 , n74382 , n65650 );
and ( n74384 , n74379 , n74383 );
and ( n74385 , n70786 , n66016 );
and ( n74386 , n70792 , n66014 );
nor ( n74387 , n74385 , n74386 );
xnor ( n74388 , n74387 , n65650 );
and ( n74389 , n74384 , n74388 );
and ( n74390 , n74388 , n74134 );
and ( n74391 , n74384 , n74134 );
or ( n74392 , n74389 , n74390 , n74391 );
and ( n74393 , n74376 , n74392 );
and ( n74394 , n70792 , n66016 );
and ( n74395 , n70802 , n66014 );
nor ( n74396 , n74394 , n74395 );
xnor ( n74397 , n74396 , n65650 );
and ( n74398 , n74392 , n74397 );
and ( n74399 , n74376 , n74397 );
or ( n74400 , n74393 , n74398 , n74399 );
and ( n74401 , n70802 , n66016 );
and ( n74402 , n70812 , n66014 );
nor ( n74403 , n74401 , n74402 );
xnor ( n74404 , n74403 , n65650 );
and ( n74405 , n74400 , n74404 );
xor ( n74406 , n74141 , n74145 );
xor ( n74407 , n74406 , n73845 );
and ( n74408 , n74404 , n74407 );
and ( n74409 , n74400 , n74407 );
or ( n74410 , n74405 , n74408 , n74409 );
and ( n74411 , n70812 , n66016 );
and ( n74412 , n70822 , n66014 );
nor ( n74413 , n74411 , n74412 );
xnor ( n74414 , n74413 , n65650 );
and ( n74415 , n74410 , n74414 );
xor ( n74416 , n74133 , n74149 );
xor ( n74417 , n74416 , n74154 );
and ( n74418 , n74414 , n74417 );
and ( n74419 , n74410 , n74417 );
or ( n74420 , n74415 , n74418 , n74419 );
and ( n74421 , n70822 , n66016 );
and ( n74422 , n70832 , n66014 );
nor ( n74423 , n74421 , n74422 );
xnor ( n74424 , n74423 , n65650 );
and ( n74425 , n74420 , n74424 );
xor ( n74426 , n74157 , n74161 );
xor ( n74427 , n74426 , n74164 );
and ( n74428 , n74424 , n74427 );
and ( n74429 , n74420 , n74427 );
or ( n74430 , n74425 , n74428 , n74429 );
and ( n74431 , n70832 , n66016 );
and ( n74432 , n70766 , n66014 );
nor ( n74433 , n74431 , n74432 );
xnor ( n74434 , n74433 , n65650 );
and ( n74435 , n74430 , n74434 );
xor ( n74436 , n74167 , n74171 );
xor ( n74437 , n74436 , n74174 );
and ( n74438 , n74434 , n74437 );
and ( n74439 , n74430 , n74437 );
or ( n74440 , n74435 , n74438 , n74439 );
and ( n74441 , n70766 , n66016 );
and ( n74442 , n70266 , n66014 );
nor ( n74443 , n74441 , n74442 );
xnor ( n74444 , n74443 , n65650 );
and ( n74445 , n74440 , n74444 );
xor ( n74446 , n74177 , n74181 );
xor ( n74447 , n74446 , n74184 );
and ( n74448 , n74444 , n74447 );
and ( n74449 , n74440 , n74447 );
or ( n74450 , n74445 , n74448 , n74449 );
and ( n74451 , n69979 , n66657 );
and ( n74452 , n69573 , n66655 );
nor ( n74453 , n74451 , n74452 );
xnor ( n74454 , n74453 , n66130 );
and ( n74455 , n74450 , n74454 );
xor ( n74456 , n74221 , n74225 );
xor ( n74457 , n74456 , n74228 );
and ( n74458 , n74454 , n74457 );
and ( n74459 , n74450 , n74457 );
or ( n74460 , n74455 , n74458 , n74459 );
and ( n74461 , n69985 , n66657 );
and ( n74462 , n69979 , n66655 );
nor ( n74463 , n74461 , n74462 );
xnor ( n74464 , n74463 , n66130 );
and ( n74465 , n70252 , n66241 );
and ( n74466 , n70238 , n66239 );
nor ( n74467 , n74465 , n74466 );
xnor ( n74468 , n74467 , n65876 );
and ( n74469 , n74464 , n74468 );
xor ( n74470 , n74440 , n74444 );
xor ( n74471 , n74470 , n74447 );
and ( n74472 , n74468 , n74471 );
and ( n74473 , n74464 , n74471 );
or ( n74474 , n74469 , n74472 , n74473 );
and ( n74475 , n69566 , n66906 );
and ( n74476 , n69568 , n66904 );
nor ( n74477 , n74475 , n74476 );
xnor ( n74478 , n74477 , n66286 );
and ( n74479 , n74474 , n74478 );
xor ( n74480 , n74450 , n74454 );
xor ( n74481 , n74480 , n74457 );
and ( n74482 , n74478 , n74481 );
and ( n74483 , n74474 , n74481 );
or ( n74484 , n74479 , n74482 , n74483 );
and ( n74485 , n74460 , n74484 );
xor ( n74486 , n74333 , n74337 );
xor ( n74487 , n74486 , n74340 );
and ( n74488 , n74484 , n74487 );
and ( n74489 , n74460 , n74487 );
or ( n74490 , n74485 , n74488 , n74489 );
and ( n74491 , n68625 , n67498 );
and ( n74492 , n68444 , n67495 );
nor ( n74493 , n74491 , n74492 );
xnor ( n74494 , n74493 , n66511 );
and ( n74495 , n74490 , n74494 );
and ( n74496 , n69449 , n66906 );
and ( n74497 , n69095 , n66904 );
nor ( n74498 , n74496 , n74497 );
xnor ( n74499 , n74498 , n66286 );
and ( n74500 , n74494 , n74499 );
and ( n74501 , n74490 , n74499 );
or ( n74502 , n74495 , n74500 , n74501 );
xor ( n74503 , n74353 , n74357 );
xor ( n74504 , n74503 , n74362 );
and ( n74505 , n74502 , n74504 );
xor ( n74506 , n74297 , n74301 );
xor ( n74507 , n74506 , n74304 );
and ( n74508 , n74504 , n74507 );
and ( n74509 , n74502 , n74507 );
or ( n74510 , n74505 , n74508 , n74509 );
xor ( n74511 , n74365 , n74367 );
xor ( n74512 , n74511 , n74370 );
and ( n74513 , n74510 , n74512 );
xor ( n74514 , n74510 , n74512 );
xor ( n74515 , n74502 , n74504 );
xor ( n74516 , n74515 , n74507 );
and ( n74517 , n69095 , n67160 );
and ( n74518 , n68873 , n67158 );
nor ( n74519 , n74517 , n74518 );
xnor ( n74520 , n74519 , n66514 );
and ( n74521 , n69568 , n66906 );
and ( n74522 , n69449 , n66904 );
nor ( n74523 , n74521 , n74522 );
xnor ( n74524 , n74523 , n66286 );
and ( n74525 , n74520 , n74524 );
xor ( n74526 , n74460 , n74484 );
xor ( n74527 , n74526 , n74487 );
and ( n74528 , n74524 , n74527 );
and ( n74529 , n74520 , n74527 );
or ( n74530 , n74525 , n74528 , n74529 );
xor ( n74531 , n74490 , n74494 );
xor ( n74532 , n74531 , n74499 );
and ( n74533 , n74530 , n74532 );
xor ( n74534 , n74343 , n74347 );
xor ( n74535 , n74534 , n74350 );
and ( n74536 , n74532 , n74535 );
and ( n74537 , n74530 , n74535 );
or ( n74538 , n74533 , n74536 , n74537 );
and ( n74539 , n74516 , n74538 );
xor ( n74540 , n74516 , n74538 );
xor ( n74541 , n74530 , n74532 );
xor ( n74542 , n74541 , n74535 );
and ( n74543 , n70238 , n66657 );
and ( n74544 , n69985 , n66655 );
nor ( n74545 , n74543 , n74544 );
xnor ( n74546 , n74545 , n66130 );
and ( n74547 , n70266 , n66241 );
and ( n74548 , n70252 , n66239 );
nor ( n74549 , n74547 , n74548 );
xnor ( n74550 , n74549 , n65876 );
and ( n74551 , n74546 , n74550 );
xor ( n74552 , n74430 , n74434 );
xor ( n74553 , n74552 , n74437 );
and ( n74554 , n74550 , n74553 );
and ( n74555 , n74546 , n74553 );
or ( n74556 , n74551 , n74554 , n74555 );
and ( n74557 , n69573 , n66906 );
and ( n74558 , n69566 , n66904 );
nor ( n74559 , n74557 , n74558 );
xnor ( n74560 , n74559 , n66286 );
and ( n74561 , n74556 , n74560 );
xor ( n74562 , n74464 , n74468 );
xor ( n74563 , n74562 , n74471 );
and ( n74564 , n74560 , n74563 );
and ( n74565 , n74556 , n74563 );
or ( n74566 , n74561 , n74564 , n74565 );
xor ( n74567 , n74379 , n74383 );
and ( n74568 , n70781 , n66239 );
not ( n74569 , n74568 );
and ( n74570 , n74569 , n65876 );
and ( n74571 , n70781 , n66241 );
and ( n74572 , n70786 , n66239 );
nor ( n74573 , n74571 , n74572 );
xnor ( n74574 , n74573 , n65876 );
and ( n74575 , n74570 , n74574 );
and ( n74576 , n70786 , n66241 );
and ( n74577 , n70792 , n66239 );
nor ( n74578 , n74576 , n74577 );
xnor ( n74579 , n74578 , n65876 );
and ( n74580 , n74575 , n74579 );
and ( n74581 , n74579 , n74377 );
and ( n74582 , n74575 , n74377 );
or ( n74583 , n74580 , n74581 , n74582 );
and ( n74584 , n74567 , n74583 );
and ( n74585 , n70792 , n66241 );
and ( n74586 , n70802 , n66239 );
nor ( n74587 , n74585 , n74586 );
xnor ( n74588 , n74587 , n65876 );
and ( n74589 , n74583 , n74588 );
and ( n74590 , n74567 , n74588 );
or ( n74591 , n74584 , n74589 , n74590 );
and ( n74592 , n70802 , n66241 );
and ( n74593 , n70812 , n66239 );
nor ( n74594 , n74592 , n74593 );
xnor ( n74595 , n74594 , n65876 );
and ( n74596 , n74591 , n74595 );
xor ( n74597 , n74384 , n74388 );
xor ( n74598 , n74597 , n74134 );
and ( n74599 , n74595 , n74598 );
and ( n74600 , n74591 , n74598 );
or ( n74601 , n74596 , n74599 , n74600 );
and ( n74602 , n70812 , n66241 );
and ( n74603 , n70822 , n66239 );
nor ( n74604 , n74602 , n74603 );
xnor ( n74605 , n74604 , n65876 );
and ( n74606 , n74601 , n74605 );
xor ( n74607 , n74376 , n74392 );
xor ( n74608 , n74607 , n74397 );
and ( n74609 , n74605 , n74608 );
and ( n74610 , n74601 , n74608 );
or ( n74611 , n74606 , n74609 , n74610 );
and ( n74612 , n70822 , n66241 );
and ( n74613 , n70832 , n66239 );
nor ( n74614 , n74612 , n74613 );
xnor ( n74615 , n74614 , n65876 );
and ( n74616 , n74611 , n74615 );
xor ( n74617 , n74400 , n74404 );
xor ( n74618 , n74617 , n74407 );
and ( n74619 , n74615 , n74618 );
and ( n74620 , n74611 , n74618 );
or ( n74621 , n74616 , n74619 , n74620 );
and ( n74622 , n70832 , n66241 );
and ( n74623 , n70766 , n66239 );
nor ( n74624 , n74622 , n74623 );
xnor ( n74625 , n74624 , n65876 );
and ( n74626 , n74621 , n74625 );
xor ( n74627 , n74410 , n74414 );
xor ( n74628 , n74627 , n74417 );
and ( n74629 , n74625 , n74628 );
and ( n74630 , n74621 , n74628 );
or ( n74631 , n74626 , n74629 , n74630 );
and ( n74632 , n70766 , n66241 );
and ( n74633 , n70266 , n66239 );
nor ( n74634 , n74632 , n74633 );
xnor ( n74635 , n74634 , n65876 );
and ( n74636 , n74631 , n74635 );
xor ( n74637 , n74420 , n74424 );
xor ( n74638 , n74637 , n74427 );
and ( n74639 , n74635 , n74638 );
and ( n74640 , n74631 , n74638 );
or ( n74641 , n74636 , n74639 , n74640 );
and ( n74642 , n69979 , n66906 );
and ( n74643 , n69573 , n66904 );
nor ( n74644 , n74642 , n74643 );
xnor ( n74645 , n74644 , n66286 );
and ( n74646 , n74641 , n74645 );
xor ( n74647 , n74546 , n74550 );
xor ( n74648 , n74647 , n74553 );
and ( n74649 , n74645 , n74648 );
and ( n74650 , n74641 , n74648 );
or ( n74651 , n74646 , n74649 , n74650 );
and ( n74652 , n70238 , n66906 );
and ( n74653 , n69985 , n66904 );
nor ( n74654 , n74652 , n74653 );
xnor ( n74655 , n74654 , n66286 );
and ( n74656 , n70266 , n66657 );
and ( n74657 , n70252 , n66655 );
nor ( n74658 , n74656 , n74657 );
xnor ( n74659 , n74658 , n66130 );
and ( n74660 , n74655 , n74659 );
xor ( n74661 , n74621 , n74625 );
xor ( n74662 , n74661 , n74628 );
and ( n74663 , n74659 , n74662 );
and ( n74664 , n74655 , n74662 );
or ( n74665 , n74660 , n74663 , n74664 );
and ( n74666 , n70252 , n66657 );
and ( n74667 , n70238 , n66655 );
nor ( n74668 , n74666 , n74667 );
xnor ( n74669 , n74668 , n66130 );
and ( n74670 , n74665 , n74669 );
xor ( n74671 , n74631 , n74635 );
xor ( n74672 , n74671 , n74638 );
and ( n74673 , n74669 , n74672 );
and ( n74674 , n74665 , n74672 );
or ( n74675 , n74670 , n74673 , n74674 );
and ( n74676 , n69566 , n67160 );
and ( n74677 , n69568 , n67158 );
nor ( n74678 , n74676 , n74677 );
xnor ( n74679 , n74678 , n66514 );
and ( n74680 , n74675 , n74679 );
xor ( n74681 , n74641 , n74645 );
xor ( n74682 , n74681 , n74648 );
and ( n74683 , n74679 , n74682 );
and ( n74684 , n74675 , n74682 );
or ( n74685 , n74680 , n74683 , n74684 );
and ( n74686 , n74651 , n74685 );
xor ( n74687 , n74556 , n74560 );
xor ( n74688 , n74687 , n74563 );
and ( n74689 , n74685 , n74688 );
and ( n74690 , n74651 , n74688 );
or ( n74691 , n74686 , n74689 , n74690 );
and ( n74692 , n74566 , n74691 );
xor ( n74693 , n74474 , n74478 );
xor ( n74694 , n74693 , n74481 );
and ( n74695 , n74691 , n74694 );
and ( n74696 , n74566 , n74694 );
or ( n74697 , n74692 , n74695 , n74696 );
and ( n74698 , n68837 , n67498 );
and ( n74699 , n68625 , n67495 );
nor ( n74700 , n74698 , n74699 );
xnor ( n74701 , n74700 , n66511 );
and ( n74702 , n74697 , n74701 );
xor ( n74703 , n74520 , n74524 );
xor ( n74704 , n74703 , n74527 );
and ( n74705 , n74701 , n74704 );
and ( n74706 , n74697 , n74704 );
or ( n74707 , n74702 , n74705 , n74706 );
and ( n74708 , n74542 , n74707 );
xor ( n74709 , n74542 , n74707 );
xor ( n74710 , n74697 , n74701 );
xor ( n74711 , n74710 , n74704 );
and ( n74712 , n68873 , n67498 );
and ( n74713 , n68837 , n67495 );
nor ( n74714 , n74712 , n74713 );
xnor ( n74715 , n74714 , n66511 );
and ( n74716 , n69449 , n67160 );
and ( n74717 , n69095 , n67158 );
nor ( n74718 , n74716 , n74717 );
xnor ( n74719 , n74718 , n66514 );
and ( n74720 , n74715 , n74719 );
xor ( n74721 , n74566 , n74691 );
xor ( n74722 , n74721 , n74694 );
and ( n74723 , n74719 , n74722 );
and ( n74724 , n74715 , n74722 );
or ( n74725 , n74720 , n74723 , n74724 );
and ( n74726 , n74711 , n74725 );
xor ( n74727 , n74711 , n74725 );
and ( n74728 , n69095 , n67498 );
and ( n74729 , n68873 , n67495 );
nor ( n74730 , n74728 , n74729 );
xnor ( n74731 , n74730 , n66511 );
and ( n74732 , n69568 , n67160 );
and ( n74733 , n69449 , n67158 );
nor ( n74734 , n74732 , n74733 );
xnor ( n74735 , n74734 , n66514 );
and ( n74736 , n74731 , n74735 );
xor ( n74737 , n74651 , n74685 );
xor ( n74738 , n74737 , n74688 );
and ( n74739 , n74735 , n74738 );
and ( n74740 , n74731 , n74738 );
or ( n74741 , n74736 , n74739 , n74740 );
xor ( n74742 , n74715 , n74719 );
xor ( n74743 , n74742 , n74722 );
and ( n74744 , n74741 , n74743 );
xor ( n74745 , n74741 , n74743 );
and ( n74746 , n69573 , n67160 );
and ( n74747 , n69566 , n67158 );
nor ( n74748 , n74746 , n74747 );
xnor ( n74749 , n74748 , n66514 );
and ( n74750 , n69985 , n66906 );
and ( n74751 , n69979 , n66904 );
nor ( n74752 , n74750 , n74751 );
xnor ( n74753 , n74752 , n66286 );
and ( n74754 , n74749 , n74753 );
xor ( n74755 , n74665 , n74669 );
xor ( n74756 , n74755 , n74672 );
and ( n74757 , n74753 , n74756 );
and ( n74758 , n74749 , n74756 );
or ( n74759 , n74754 , n74757 , n74758 );
and ( n74760 , n69449 , n67498 );
and ( n74761 , n69095 , n67495 );
nor ( n74762 , n74760 , n74761 );
xnor ( n74763 , n74762 , n66511 );
and ( n74764 , n74759 , n74763 );
xor ( n74765 , n74675 , n74679 );
xor ( n74766 , n74765 , n74682 );
and ( n74767 , n74763 , n74766 );
and ( n74768 , n74759 , n74766 );
or ( n74769 , n74764 , n74767 , n74768 );
xor ( n74770 , n74731 , n74735 );
xor ( n74771 , n74770 , n74738 );
and ( n74772 , n74769 , n74771 );
xor ( n74773 , n74769 , n74771 );
xor ( n74774 , n74759 , n74763 );
xor ( n74775 , n74774 , n74766 );
xor ( n74776 , n74570 , n74574 );
and ( n74777 , n70781 , n66655 );
not ( n74778 , n74777 );
and ( n74779 , n74778 , n66130 );
and ( n74780 , n70781 , n66657 );
and ( n74781 , n70786 , n66655 );
nor ( n74782 , n74780 , n74781 );
xnor ( n74783 , n74782 , n66130 );
and ( n74784 , n74779 , n74783 );
and ( n74785 , n70786 , n66657 );
and ( n74786 , n70792 , n66655 );
nor ( n74787 , n74785 , n74786 );
xnor ( n74788 , n74787 , n66130 );
and ( n74789 , n74784 , n74788 );
and ( n74790 , n74788 , n74568 );
and ( n74791 , n74784 , n74568 );
or ( n74792 , n74789 , n74790 , n74791 );
and ( n74793 , n74776 , n74792 );
and ( n74794 , n70792 , n66657 );
and ( n74795 , n70802 , n66655 );
nor ( n74796 , n74794 , n74795 );
xnor ( n74797 , n74796 , n66130 );
and ( n74798 , n74792 , n74797 );
and ( n74799 , n74776 , n74797 );
or ( n74800 , n74793 , n74798 , n74799 );
and ( n74801 , n70802 , n66657 );
and ( n74802 , n70812 , n66655 );
nor ( n74803 , n74801 , n74802 );
xnor ( n74804 , n74803 , n66130 );
and ( n74805 , n74800 , n74804 );
xor ( n74806 , n74575 , n74579 );
xor ( n74807 , n74806 , n74377 );
and ( n74808 , n74804 , n74807 );
and ( n74809 , n74800 , n74807 );
or ( n74810 , n74805 , n74808 , n74809 );
and ( n74811 , n70812 , n66657 );
and ( n74812 , n70822 , n66655 );
nor ( n74813 , n74811 , n74812 );
xnor ( n74814 , n74813 , n66130 );
and ( n74815 , n74810 , n74814 );
xor ( n74816 , n74567 , n74583 );
xor ( n74817 , n74816 , n74588 );
and ( n74818 , n74814 , n74817 );
and ( n74819 , n74810 , n74817 );
or ( n74820 , n74815 , n74818 , n74819 );
and ( n74821 , n70822 , n66657 );
and ( n74822 , n70832 , n66655 );
nor ( n74823 , n74821 , n74822 );
xnor ( n74824 , n74823 , n66130 );
and ( n74825 , n74820 , n74824 );
xor ( n74826 , n74591 , n74595 );
xor ( n74827 , n74826 , n74598 );
and ( n74828 , n74824 , n74827 );
and ( n74829 , n74820 , n74827 );
or ( n74830 , n74825 , n74828 , n74829 );
and ( n74831 , n70832 , n66657 );
and ( n74832 , n70766 , n66655 );
nor ( n74833 , n74831 , n74832 );
xnor ( n74834 , n74833 , n66130 );
and ( n74835 , n74830 , n74834 );
xor ( n74836 , n74601 , n74605 );
xor ( n74837 , n74836 , n74608 );
and ( n74838 , n74834 , n74837 );
and ( n74839 , n74830 , n74837 );
or ( n74840 , n74835 , n74838 , n74839 );
and ( n74841 , n70766 , n66657 );
and ( n74842 , n70266 , n66655 );
nor ( n74843 , n74841 , n74842 );
xnor ( n74844 , n74843 , n66130 );
and ( n74845 , n74840 , n74844 );
xor ( n74846 , n74611 , n74615 );
xor ( n74847 , n74846 , n74618 );
and ( n74848 , n74844 , n74847 );
and ( n74849 , n74840 , n74847 );
or ( n74850 , n74845 , n74848 , n74849 );
and ( n74851 , n69979 , n67160 );
and ( n74852 , n69573 , n67158 );
nor ( n74853 , n74851 , n74852 );
xnor ( n74854 , n74853 , n66514 );
and ( n74855 , n74850 , n74854 );
xor ( n74856 , n74655 , n74659 );
xor ( n74857 , n74856 , n74662 );
and ( n74858 , n74854 , n74857 );
and ( n74859 , n74850 , n74857 );
or ( n74860 , n74855 , n74858 , n74859 );
and ( n74861 , n70238 , n67160 );
and ( n74862 , n69985 , n67158 );
nor ( n74863 , n74861 , n74862 );
xnor ( n74864 , n74863 , n66514 );
and ( n74865 , n70266 , n66906 );
and ( n74866 , n70252 , n66904 );
nor ( n74867 , n74865 , n74866 );
xnor ( n74868 , n74867 , n66286 );
and ( n74869 , n74864 , n74868 );
xor ( n74870 , n74830 , n74834 );
xor ( n74871 , n74870 , n74837 );
and ( n74872 , n74868 , n74871 );
and ( n74873 , n74864 , n74871 );
or ( n74874 , n74869 , n74872 , n74873 );
and ( n74875 , n70252 , n66906 );
and ( n74876 , n70238 , n66904 );
nor ( n74877 , n74875 , n74876 );
xnor ( n74878 , n74877 , n66286 );
and ( n74879 , n74874 , n74878 );
xor ( n74880 , n74840 , n74844 );
xor ( n74881 , n74880 , n74847 );
and ( n74882 , n74878 , n74881 );
and ( n74883 , n74874 , n74881 );
or ( n74884 , n74879 , n74882 , n74883 );
and ( n74885 , n69566 , n67498 );
and ( n74886 , n69568 , n67495 );
nor ( n74887 , n74885 , n74886 );
xnor ( n74888 , n74887 , n66511 );
and ( n74889 , n74884 , n74888 );
xor ( n74890 , n74850 , n74854 );
xor ( n74891 , n74890 , n74857 );
and ( n74892 , n74888 , n74891 );
and ( n74893 , n74884 , n74891 );
or ( n74894 , n74889 , n74892 , n74893 );
and ( n74895 , n74860 , n74894 );
xor ( n74896 , n74749 , n74753 );
xor ( n74897 , n74896 , n74756 );
and ( n74898 , n74894 , n74897 );
and ( n74899 , n74860 , n74897 );
or ( n74900 , n74895 , n74898 , n74899 );
and ( n74901 , n74775 , n74900 );
xor ( n74902 , n74775 , n74900 );
and ( n74903 , n69568 , n67498 );
and ( n74904 , n69449 , n67495 );
nor ( n74905 , n74903 , n74904 );
xnor ( n74906 , n74905 , n66511 );
xor ( n74907 , n74860 , n74894 );
xor ( n74908 , n74907 , n74897 );
and ( n74909 , n74906 , n74908 );
xor ( n74910 , n74906 , n74908 );
xor ( n74911 , n74884 , n74888 );
xor ( n74912 , n74911 , n74891 );
and ( n74913 , n69573 , n67498 );
and ( n74914 , n69566 , n67495 );
nor ( n74915 , n74913 , n74914 );
xnor ( n74916 , n74915 , n66511 );
and ( n74917 , n69985 , n67160 );
and ( n74918 , n69979 , n67158 );
nor ( n74919 , n74917 , n74918 );
xnor ( n74920 , n74919 , n66514 );
and ( n74921 , n74916 , n74920 );
xor ( n74922 , n74874 , n74878 );
xor ( n74923 , n74922 , n74881 );
and ( n74924 , n74920 , n74923 );
and ( n74925 , n74916 , n74923 );
or ( n74926 , n74921 , n74924 , n74925 );
and ( n74927 , n74912 , n74926 );
xor ( n74928 , n74912 , n74926 );
xor ( n74929 , n74779 , n74783 );
and ( n74930 , n70781 , n66904 );
not ( n74931 , n74930 );
and ( n74932 , n74931 , n66286 );
and ( n74933 , n70781 , n66906 );
and ( n74934 , n70786 , n66904 );
nor ( n74935 , n74933 , n74934 );
xnor ( n74936 , n74935 , n66286 );
and ( n74937 , n74932 , n74936 );
and ( n74938 , n70786 , n66906 );
and ( n74939 , n70792 , n66904 );
nor ( n74940 , n74938 , n74939 );
xnor ( n74941 , n74940 , n66286 );
and ( n74942 , n74937 , n74941 );
and ( n74943 , n74941 , n74777 );
and ( n74944 , n74937 , n74777 );
or ( n74945 , n74942 , n74943 , n74944 );
and ( n74946 , n74929 , n74945 );
and ( n74947 , n70792 , n66906 );
and ( n74948 , n70802 , n66904 );
nor ( n74949 , n74947 , n74948 );
xnor ( n74950 , n74949 , n66286 );
and ( n74951 , n74945 , n74950 );
and ( n74952 , n74929 , n74950 );
or ( n74953 , n74946 , n74951 , n74952 );
and ( n74954 , n70802 , n66906 );
and ( n74955 , n70812 , n66904 );
nor ( n74956 , n74954 , n74955 );
xnor ( n74957 , n74956 , n66286 );
and ( n74958 , n74953 , n74957 );
xor ( n74959 , n74784 , n74788 );
xor ( n74960 , n74959 , n74568 );
and ( n74961 , n74957 , n74960 );
and ( n74962 , n74953 , n74960 );
or ( n74963 , n74958 , n74961 , n74962 );
and ( n74964 , n70812 , n66906 );
and ( n74965 , n70822 , n66904 );
nor ( n74966 , n74964 , n74965 );
xnor ( n74967 , n74966 , n66286 );
and ( n74968 , n74963 , n74967 );
xor ( n74969 , n74776 , n74792 );
xor ( n74970 , n74969 , n74797 );
and ( n74971 , n74967 , n74970 );
and ( n74972 , n74963 , n74970 );
or ( n74973 , n74968 , n74971 , n74972 );
and ( n74974 , n70822 , n66906 );
and ( n74975 , n70832 , n66904 );
nor ( n74976 , n74974 , n74975 );
xnor ( n74977 , n74976 , n66286 );
and ( n74978 , n74973 , n74977 );
xor ( n74979 , n74800 , n74804 );
xor ( n74980 , n74979 , n74807 );
and ( n74981 , n74977 , n74980 );
and ( n74982 , n74973 , n74980 );
or ( n74983 , n74978 , n74981 , n74982 );
and ( n74984 , n70832 , n66906 );
and ( n74985 , n70766 , n66904 );
nor ( n74986 , n74984 , n74985 );
xnor ( n74987 , n74986 , n66286 );
and ( n74988 , n74983 , n74987 );
xor ( n74989 , n74810 , n74814 );
xor ( n74990 , n74989 , n74817 );
and ( n74991 , n74987 , n74990 );
and ( n74992 , n74983 , n74990 );
or ( n74993 , n74988 , n74991 , n74992 );
and ( n74994 , n70766 , n66906 );
and ( n74995 , n70266 , n66904 );
nor ( n74996 , n74994 , n74995 );
xnor ( n74997 , n74996 , n66286 );
and ( n74998 , n74993 , n74997 );
xor ( n74999 , n74820 , n74824 );
xor ( n75000 , n74999 , n74827 );
and ( n75001 , n74997 , n75000 );
and ( n75002 , n74993 , n75000 );
or ( n75003 , n74998 , n75001 , n75002 );
and ( n75004 , n69979 , n67498 );
and ( n75005 , n69573 , n67495 );
nor ( n75006 , n75004 , n75005 );
xnor ( n75007 , n75006 , n66511 );
and ( n75008 , n75003 , n75007 );
xor ( n75009 , n74864 , n74868 );
xor ( n75010 , n75009 , n74871 );
and ( n75011 , n75007 , n75010 );
and ( n75012 , n75003 , n75010 );
or ( n75013 , n75008 , n75011 , n75012 );
xor ( n75014 , n74916 , n74920 );
xor ( n75015 , n75014 , n74923 );
and ( n75016 , n75013 , n75015 );
xor ( n75017 , n75013 , n75015 );
xor ( n75018 , n75003 , n75007 );
xor ( n75019 , n75018 , n75010 );
and ( n75020 , n70238 , n67498 );
and ( n75021 , n69985 , n67495 );
nor ( n75022 , n75020 , n75021 );
xnor ( n75023 , n75022 , n66511 );
and ( n75024 , n70266 , n67160 );
and ( n75025 , n70252 , n67158 );
nor ( n75026 , n75024 , n75025 );
xnor ( n75027 , n75026 , n66514 );
and ( n75028 , n75023 , n75027 );
xor ( n75029 , n74983 , n74987 );
xor ( n75030 , n75029 , n74990 );
and ( n75031 , n75027 , n75030 );
and ( n75032 , n75023 , n75030 );
or ( n75033 , n75028 , n75031 , n75032 );
and ( n75034 , n70252 , n67160 );
and ( n75035 , n70238 , n67158 );
nor ( n75036 , n75034 , n75035 );
xnor ( n75037 , n75036 , n66514 );
and ( n75038 , n75033 , n75037 );
xor ( n75039 , n74993 , n74997 );
xor ( n75040 , n75039 , n75000 );
and ( n75041 , n75037 , n75040 );
and ( n75042 , n75033 , n75040 );
or ( n75043 , n75038 , n75041 , n75042 );
and ( n75044 , n75019 , n75043 );
xor ( n75045 , n75019 , n75043 );
and ( n75046 , n69985 , n67498 );
and ( n75047 , n69979 , n67495 );
nor ( n75048 , n75046 , n75047 );
xnor ( n75049 , n75048 , n66511 );
xor ( n75050 , n75033 , n75037 );
xor ( n75051 , n75050 , n75040 );
and ( n75052 , n75049 , n75051 );
xor ( n75053 , n75049 , n75051 );
xor ( n75054 , n75023 , n75027 );
xor ( n75055 , n75054 , n75030 );
xor ( n75056 , n74932 , n74936 );
and ( n75057 , n70781 , n67158 );
not ( n75058 , n75057 );
and ( n75059 , n75058 , n66514 );
and ( n75060 , n70781 , n67160 );
and ( n75061 , n70786 , n67158 );
nor ( n75062 , n75060 , n75061 );
xnor ( n75063 , n75062 , n66514 );
and ( n75064 , n75059 , n75063 );
and ( n75065 , n70786 , n67160 );
and ( n75066 , n70792 , n67158 );
nor ( n75067 , n75065 , n75066 );
xnor ( n75068 , n75067 , n66514 );
and ( n75069 , n75064 , n75068 );
and ( n75070 , n75068 , n74930 );
and ( n75071 , n75064 , n74930 );
or ( n75072 , n75069 , n75070 , n75071 );
and ( n75073 , n75056 , n75072 );
and ( n75074 , n70792 , n67160 );
and ( n75075 , n70802 , n67158 );
nor ( n75076 , n75074 , n75075 );
xnor ( n75077 , n75076 , n66514 );
and ( n75078 , n75072 , n75077 );
and ( n75079 , n75056 , n75077 );
or ( n75080 , n75073 , n75078 , n75079 );
and ( n75081 , n70802 , n67160 );
and ( n75082 , n70812 , n67158 );
nor ( n75083 , n75081 , n75082 );
xnor ( n75084 , n75083 , n66514 );
and ( n75085 , n75080 , n75084 );
xor ( n75086 , n74937 , n74941 );
xor ( n75087 , n75086 , n74777 );
and ( n75088 , n75084 , n75087 );
and ( n75089 , n75080 , n75087 );
or ( n75090 , n75085 , n75088 , n75089 );
and ( n75091 , n70812 , n67160 );
and ( n75092 , n70822 , n67158 );
nor ( n75093 , n75091 , n75092 );
xnor ( n75094 , n75093 , n66514 );
and ( n75095 , n75090 , n75094 );
xor ( n75096 , n74929 , n74945 );
xor ( n75097 , n75096 , n74950 );
and ( n75098 , n75094 , n75097 );
and ( n75099 , n75090 , n75097 );
or ( n75100 , n75095 , n75098 , n75099 );
and ( n75101 , n70822 , n67160 );
and ( n75102 , n70832 , n67158 );
nor ( n75103 , n75101 , n75102 );
xnor ( n75104 , n75103 , n66514 );
and ( n75105 , n75100 , n75104 );
xor ( n75106 , n74953 , n74957 );
xor ( n75107 , n75106 , n74960 );
and ( n75108 , n75104 , n75107 );
and ( n75109 , n75100 , n75107 );
or ( n75110 , n75105 , n75108 , n75109 );
and ( n75111 , n70832 , n67160 );
and ( n75112 , n70766 , n67158 );
nor ( n75113 , n75111 , n75112 );
xnor ( n75114 , n75113 , n66514 );
and ( n75115 , n75110 , n75114 );
xor ( n75116 , n74963 , n74967 );
xor ( n75117 , n75116 , n74970 );
and ( n75118 , n75114 , n75117 );
and ( n75119 , n75110 , n75117 );
or ( n75120 , n75115 , n75118 , n75119 );
and ( n75121 , n70766 , n67160 );
and ( n75122 , n70266 , n67158 );
nor ( n75123 , n75121 , n75122 );
xnor ( n75124 , n75123 , n66514 );
and ( n75125 , n75120 , n75124 );
xor ( n75126 , n74973 , n74977 );
xor ( n75127 , n75126 , n74980 );
and ( n75128 , n75124 , n75127 );
and ( n75129 , n75120 , n75127 );
or ( n75130 , n75125 , n75128 , n75129 );
and ( n75131 , n75055 , n75130 );
xor ( n75132 , n75055 , n75130 );
and ( n75133 , n70252 , n67498 );
and ( n75134 , n70238 , n67495 );
nor ( n75135 , n75133 , n75134 );
xnor ( n75136 , n75135 , n66511 );
xor ( n75137 , n75120 , n75124 );
xor ( n75138 , n75137 , n75127 );
and ( n75139 , n75136 , n75138 );
xor ( n75140 , n75136 , n75138 );
and ( n75141 , n70266 , n67498 );
and ( n75142 , n70252 , n67495 );
nor ( n75143 , n75141 , n75142 );
xnor ( n75144 , n75143 , n66511 );
xor ( n75145 , n75110 , n75114 );
xor ( n75146 , n75145 , n75117 );
and ( n75147 , n75144 , n75146 );
xor ( n75148 , n75144 , n75146 );
and ( n75149 , n70766 , n67498 );
and ( n75150 , n70266 , n67495 );
nor ( n75151 , n75149 , n75150 );
xnor ( n75152 , n75151 , n66511 );
xor ( n75153 , n75100 , n75104 );
xor ( n75154 , n75153 , n75107 );
and ( n75155 , n75152 , n75154 );
xor ( n75156 , n75152 , n75154 );
and ( n75157 , n70832 , n67498 );
and ( n75158 , n70766 , n67495 );
nor ( n75159 , n75157 , n75158 );
xnor ( n75160 , n75159 , n66511 );
xor ( n75161 , n75090 , n75094 );
xor ( n75162 , n75161 , n75097 );
and ( n75163 , n75160 , n75162 );
xor ( n75164 , n75160 , n75162 );
and ( n75165 , n70822 , n67498 );
and ( n75166 , n70832 , n67495 );
nor ( n75167 , n75165 , n75166 );
xnor ( n75168 , n75167 , n66511 );
xor ( n75169 , n75080 , n75084 );
xor ( n75170 , n75169 , n75087 );
and ( n75171 , n75168 , n75170 );
xor ( n75172 , n75168 , n75170 );
and ( n75173 , n70812 , n67498 );
and ( n75174 , n70822 , n67495 );
nor ( n75175 , n75173 , n75174 );
xnor ( n75176 , n75175 , n66511 );
xor ( n75177 , n75056 , n75072 );
xor ( n75178 , n75177 , n75077 );
and ( n75179 , n75176 , n75178 );
xor ( n75180 , n75176 , n75178 );
and ( n75181 , n70802 , n67498 );
and ( n75182 , n70812 , n67495 );
nor ( n75183 , n75181 , n75182 );
xnor ( n75184 , n75183 , n66511 );
xor ( n75185 , n75064 , n75068 );
xor ( n75186 , n75185 , n74930 );
and ( n75187 , n75184 , n75186 );
xor ( n75188 , n75184 , n75186 );
and ( n75189 , n70792 , n67498 );
and ( n75190 , n70802 , n67495 );
nor ( n75191 , n75189 , n75190 );
xnor ( n75192 , n75191 , n66511 );
xor ( n75193 , n75059 , n75063 );
and ( n75194 , n75192 , n75193 );
xor ( n75195 , n75192 , n75193 );
and ( n75196 , n70786 , n67498 );
and ( n75197 , n70792 , n67495 );
nor ( n75198 , n75196 , n75197 );
xnor ( n75199 , n75198 , n66511 );
and ( n75200 , n75199 , n75057 );
xor ( n75201 , n75199 , n75057 );
and ( n75202 , n70781 , n67498 );
and ( n75203 , n70786 , n67495 );
nor ( n75204 , n75202 , n75203 );
xnor ( n75205 , n75204 , n66511 );
and ( n75206 , n70781 , n67495 );
not ( n75207 , n75206 );
and ( n75208 , n75207 , n66511 );
and ( n75209 , n75205 , n75208 );
and ( n75210 , n75201 , n75209 );
or ( n75211 , n75200 , n75210 );
and ( n75212 , n75195 , n75211 );
or ( n75213 , n75194 , n75212 );
and ( n75214 , n75188 , n75213 );
or ( n75215 , n75187 , n75214 );
and ( n75216 , n75180 , n75215 );
or ( n75217 , n75179 , n75216 );
and ( n75218 , n75172 , n75217 );
or ( n75219 , n75171 , n75218 );
and ( n75220 , n75164 , n75219 );
or ( n75221 , n75163 , n75220 );
and ( n75222 , n75156 , n75221 );
or ( n75223 , n75155 , n75222 );
and ( n75224 , n75148 , n75223 );
or ( n75225 , n75147 , n75224 );
and ( n75226 , n75140 , n75225 );
or ( n75227 , n75139 , n75226 );
and ( n75228 , n75132 , n75227 );
or ( n75229 , n75131 , n75228 );
and ( n75230 , n75053 , n75229 );
or ( n75231 , n75052 , n75230 );
and ( n75232 , n75045 , n75231 );
or ( n75233 , n75044 , n75232 );
and ( n75234 , n75017 , n75233 );
or ( n75235 , n75016 , n75234 );
and ( n75236 , n74928 , n75235 );
or ( n75237 , n74927 , n75236 );
and ( n75238 , n74910 , n75237 );
or ( n75239 , n74909 , n75238 );
and ( n75240 , n74902 , n75239 );
or ( n75241 , n74901 , n75240 );
and ( n75242 , n74773 , n75241 );
or ( n75243 , n74772 , n75242 );
and ( n75244 , n74745 , n75243 );
or ( n75245 , n74744 , n75244 );
and ( n75246 , n74727 , n75245 );
or ( n75247 , n74726 , n75246 );
and ( n75248 , n74709 , n75247 );
or ( n75249 , n74708 , n75248 );
and ( n75250 , n74540 , n75249 );
or ( n75251 , n74539 , n75250 );
and ( n75252 , n74514 , n75251 );
or ( n75253 , n74513 , n75252 );
and ( n75254 , n74375 , n75253 );
or ( n75255 , n74374 , n75254 );
and ( n75256 , n74327 , n75255 );
or ( n75257 , n74326 , n75256 );
and ( n75258 , n74291 , n75257 );
or ( n75259 , n74290 , n75258 );
and ( n75260 , n74132 , n75259 );
or ( n75261 , n74131 , n75260 );
and ( n75262 , n74064 , n75261 );
or ( n75263 , n74063 , n75262 );
and ( n75264 , n74016 , n75263 );
or ( n75265 , n74015 , n75264 );
and ( n75266 , n73827 , n75265 );
or ( n75267 , n73826 , n75266 );
and ( n75268 , n73791 , n75267 );
or ( n75269 , n73790 , n75268 );
and ( n75270 , n73735 , n75269 );
or ( n75271 , n73734 , n75270 );
and ( n75272 , n73556 , n75271 );
or ( n75273 , n73555 , n75272 );
and ( n75274 , n73480 , n75273 );
or ( n75275 , n73479 , n75274 );
and ( n75276 , n73412 , n75275 );
or ( n75277 , n73411 , n75276 );
and ( n75278 , n73191 , n75277 );
or ( n75279 , n73190 , n75278 );
and ( n75280 , n73135 , n75279 );
or ( n75281 , n73134 , n75280 );
and ( n75282 , n72896 , n75281 );
or ( n75283 , n72895 , n75282 );
and ( n75284 , n72862 , n75283 );
or ( n75285 , n72861 , n75284 );
and ( n75286 , n72720 , n75285 );
or ( n75287 , n72719 , n75286 );
and ( n75288 , n72503 , n75287 );
or ( n75289 , n72502 , n75288 );
and ( n75290 , n72395 , n75289 );
or ( n75291 , n72394 , n75290 );
and ( n75292 , n72361 , n75291 );
or ( n75293 , n72360 , n75292 );
and ( n75294 , n72104 , n75293 );
or ( n75295 , n72103 , n75294 );
and ( n75296 , n71914 , n75295 );
or ( n75297 , n71913 , n75296 );
and ( n75298 , n71675 , n75297 );
or ( n75299 , n71674 , n75298 );
and ( n75300 , n71579 , n75299 );
or ( n75301 , n71578 , n75300 );
and ( n75302 , n71461 , n75301 );
or ( n75303 , n71460 , n75302 );
and ( n75304 , n71345 , n75303 );
or ( n75305 , n71344 , n75304 );
and ( n75306 , n71056 , n75305 );
or ( n75307 , n71055 , n75306 );
and ( n75308 , n70754 , n75307 );
or ( n75309 , n70753 , n75308 );
and ( n75310 , n70608 , n75309 );
or ( n75311 , n70607 , n75310 );
and ( n75312 , n70428 , n75311 );
or ( n75313 , n70427 , n75312 );
and ( n75314 , n70396 , n75313 );
or ( n75315 , n70395 , n75314 );
and ( n75316 , n70146 , n75315 );
or ( n75317 , n70145 , n75316 );
and ( n75318 , n69958 , n75317 );
or ( n75319 , n69957 , n75318 );
and ( n75320 , n69767 , n75319 );
or ( n75321 , n69766 , n75320 );
and ( n75322 , n69559 , n75321 );
or ( n75323 , n69558 , n75322 );
and ( n75324 , n69371 , n75323 );
or ( n75325 , n69370 , n75324 );
and ( n75326 , n69223 , n75325 );
or ( n75327 , n69222 , n75326 );
and ( n75328 , n69023 , n75327 );
or ( n75329 , n69022 , n75328 );
and ( n75330 , n68979 , n75329 );
or ( n75331 , n68978 , n75330 );
and ( n75332 , n68795 , n75331 );
or ( n75333 , n68794 , n75332 );
and ( n75334 , n68532 , n75333 );
or ( n75335 , n68531 , n75334 );
and ( n75336 , n68399 , n75335 );
or ( n75337 , n68398 , n75336 );
and ( n75338 , n68185 , n75337 );
or ( n75339 , n68184 , n75338 );
and ( n75340 , n68049 , n75339 );
or ( n75341 , n68048 , n75340 );
and ( n75342 , n68011 , n75341 );
or ( n75343 , n68010 , n75342 );
and ( n75344 , n67675 , n75343 );
or ( n75345 , n67674 , n75344 );
and ( n75346 , n67492 , n75345 );
or ( n75347 , n67491 , n75346 );
and ( n75348 , n67401 , n75347 );
or ( n75349 , n67400 , n75348 );
and ( n75350 , n67298 , n75349 );
or ( n75351 , n67297 , n75350 );
and ( n75352 , n67075 , n75351 );
or ( n75353 , n67074 , n75352 );
and ( n75354 , n66975 , n75353 );
or ( n75355 , n66974 , n75354 );
and ( n75356 , n66698 , n75355 );
or ( n75357 , n66697 , n75356 );
and ( n75358 , n66504 , n75357 );
or ( n75359 , n66503 , n75358 );
and ( n75360 , n66464 , n75359 );
or ( n75361 , n66463 , n75360 );
and ( n75362 , n66203 , n75361 );
or ( n75363 , n66202 , n75362 );
and ( n75364 , n66075 , n75363 );
or ( n75365 , n66074 , n75364 );
and ( n75366 , n66053 , n75365 );
or ( n75367 , n66052 , n75366 );
and ( n75368 , n65853 , n75367 );
or ( n75369 , n65852 , n75368 );
and ( n75370 , n65750 , n75369 );
or ( n75371 , n65749 , n75370 );
and ( n75372 , n65585 , n75371 );
or ( n75373 , n65584 , n75372 );
and ( n75374 , n65512 , n75373 );
or ( n75375 , n65511 , n75374 );
and ( n75376 , n65404 , n75375 );
or ( n75377 , n65403 , n75376 );
and ( n75378 , n65303 , n75377 );
or ( n75379 , n65302 , n75378 );
and ( n75380 , n65214 , n75379 );
or ( n75381 , n65213 , n75380 );
and ( n75382 , n65101 , n75381 );
or ( n75383 , n65100 , n75382 );
and ( n75384 , n65050 , n75383 );
or ( n75385 , n65049 , n75384 );
and ( n75386 , n64936 , n75385 );
or ( n75387 , n64935 , n75386 );
and ( n75388 , n64877 , n75387 );
or ( n75389 , n64876 , n75388 );
and ( n75390 , n64818 , n75389 );
or ( n75391 , n64817 , n75390 );
and ( n75392 , n64768 , n75391 );
or ( n75393 , n64767 , n75392 );
and ( n75394 , n64731 , n75393 );
or ( n75395 , n64730 , n75394 );
and ( n75396 , n64675 , n75395 );
or ( n75397 , n64674 , n75396 );
xor ( n75398 , n64646 , n75397 );
buf ( n75399 , n75398 );
xor ( n75400 , n64675 , n75395 );
buf ( n75401 , n75400 );
xor ( n75402 , n64731 , n75393 );
buf ( n75403 , n75402 );
xor ( n75404 , n64768 , n75391 );
buf ( n75405 , n75404 );
xor ( n75406 , n64818 , n75389 );
buf ( n75407 , n75406 );
xor ( n75408 , n64877 , n75387 );
buf ( n75409 , n75408 );
xor ( n75410 , n64936 , n75385 );
buf ( n75411 , n75410 );
xor ( n75412 , n65050 , n75383 );
buf ( n75413 , n75412 );
xor ( n75414 , n65101 , n75381 );
buf ( n75415 , n75414 );
xor ( n75416 , n65214 , n75379 );
buf ( n75417 , n75416 );
xor ( n75418 , n65303 , n75377 );
buf ( n75419 , n75418 );
xor ( n75420 , n65404 , n75375 );
buf ( n75421 , n75420 );
xor ( n75422 , n65512 , n75373 );
buf ( n75423 , n75422 );
xor ( n75424 , n65585 , n75371 );
buf ( n75425 , n75424 );
xor ( n75426 , n65750 , n75369 );
buf ( n75427 , n75426 );
xor ( n75428 , n65853 , n75367 );
buf ( n75429 , n75428 );
xor ( n75430 , n66053 , n75365 );
buf ( n75431 , n75430 );
xor ( n75432 , n66075 , n75363 );
buf ( n75433 , n75432 );
xor ( n75434 , n66203 , n75361 );
buf ( n75435 , n75434 );
xor ( n75436 , n66464 , n75359 );
buf ( n75437 , n75436 );
xor ( n75438 , n66504 , n75357 );
buf ( n75439 , n75438 );
xor ( n75440 , n66698 , n75355 );
buf ( n75441 , n75440 );
xor ( n75442 , n66975 , n75353 );
buf ( n75443 , n75442 );
xor ( n75444 , n67075 , n75351 );
buf ( n75445 , n75444 );
xor ( n75446 , n67298 , n75349 );
buf ( n75447 , n75446 );
xor ( n75448 , n67401 , n75347 );
buf ( n75449 , n75448 );
xor ( n75450 , n67492 , n75345 );
buf ( n75451 , n75450 );
xor ( n75452 , n67675 , n75343 );
buf ( n75453 , n75452 );
xor ( n75454 , n68011 , n75341 );
buf ( n75455 , n75454 );
xor ( n75456 , n68049 , n75339 );
buf ( n75457 , n75456 );
xor ( n75458 , n68185 , n75337 );
buf ( n75459 , n75458 );
xor ( n75460 , n68399 , n75335 );
buf ( n75461 , n75460 );
xor ( n75462 , n68532 , n75333 );
buf ( n75463 , n75462 );
xor ( n75464 , n68795 , n75331 );
buf ( n75465 , n75464 );
xor ( n75466 , n68979 , n75329 );
buf ( n75467 , n75466 );
xor ( n75468 , n69023 , n75327 );
buf ( n75469 , n75468 );
xor ( n75470 , n69223 , n75325 );
buf ( n75471 , n75470 );
xor ( n75472 , n69371 , n75323 );
buf ( n75473 , n75472 );
xor ( n75474 , n69559 , n75321 );
buf ( n75475 , n75474 );
xor ( n75476 , n69767 , n75319 );
buf ( n75477 , n75476 );
xor ( n75478 , n69958 , n75317 );
buf ( n75479 , n75478 );
xor ( n75480 , n70146 , n75315 );
buf ( n75481 , n75480 );
xor ( n75482 , n70396 , n75313 );
buf ( n75483 , n75482 );
xor ( n75484 , n70428 , n75311 );
buf ( n75485 , n75484 );
xor ( n75486 , n70608 , n75309 );
buf ( n75487 , n75486 );
xor ( n75488 , n70754 , n75307 );
buf ( n75489 , n75488 );
xor ( n75490 , n71056 , n75305 );
buf ( n75491 , n75490 );
xor ( n75492 , n71345 , n75303 );
buf ( n75493 , n75492 );
xor ( n75494 , n71461 , n75301 );
buf ( n75495 , n75494 );
xor ( n75496 , n71579 , n75299 );
buf ( n75497 , n75496 );
xor ( n75498 , n71675 , n75297 );
buf ( n75499 , n75498 );
xor ( n75500 , n71914 , n75295 );
buf ( n75501 , n75500 );
xor ( n75502 , n72104 , n75293 );
buf ( n75503 , n75502 );
xor ( n75504 , n72361 , n75291 );
buf ( n75505 , n75504 );
xor ( n75506 , n72395 , n75289 );
buf ( n75507 , n75506 );
xor ( n75508 , n72503 , n75287 );
buf ( n75509 , n75508 );
xor ( n75510 , n72720 , n75285 );
buf ( n75511 , n75510 );
xor ( n75512 , n72862 , n75283 );
buf ( n75513 , n75512 );
xor ( n75514 , n72896 , n75281 );
buf ( n75515 , n75514 );
xor ( n75516 , n73135 , n75279 );
buf ( n75517 , n75516 );
xor ( n75518 , n73191 , n75277 );
buf ( n75519 , n75518 );
xor ( n75520 , n73412 , n75275 );
buf ( n75521 , n75520 );
xor ( n75522 , n73480 , n75273 );
buf ( n75523 , n75522 );
xor ( n75524 , n73556 , n75271 );
buf ( n75525 , n75524 );
xor ( n75526 , n73735 , n75269 );
buf ( n75527 , n75526 );
xor ( n75528 , n73791 , n75267 );
buf ( n75529 , n75528 );
xor ( n75530 , n73827 , n75265 );
buf ( n75531 , n75530 );
xor ( n75532 , n74016 , n75263 );
buf ( n75533 , n75532 );
xor ( n75534 , n74064 , n75261 );
buf ( n75535 , n75534 );
xor ( n75536 , n74132 , n75259 );
buf ( n75537 , n75536 );
xor ( n75538 , n74291 , n75257 );
buf ( n75539 , n75538 );
xor ( n75540 , n74327 , n75255 );
buf ( n75541 , n75540 );
xor ( n75542 , n74375 , n75253 );
buf ( n75543 , n75542 );
xor ( n75544 , n74514 , n75251 );
buf ( n75545 , n75544 );
xor ( n75546 , n74540 , n75249 );
buf ( n75547 , n75546 );
xor ( n75548 , n74709 , n75247 );
buf ( n75549 , n75548 );
xor ( n75550 , n74727 , n75245 );
buf ( n75551 , n75550 );
xor ( n75552 , n74745 , n75243 );
buf ( n75553 , n75552 );
xor ( n75554 , n74773 , n75241 );
buf ( n75555 , n75554 );
xor ( n75556 , n74902 , n75239 );
buf ( n75557 , n75556 );
xor ( n75558 , n74910 , n75237 );
buf ( n75559 , n75558 );
xor ( n75560 , n74928 , n75235 );
buf ( n75561 , n75560 );
xor ( n75562 , n75017 , n75233 );
buf ( n75563 , n75562 );
xor ( n75564 , n75045 , n75231 );
buf ( n75565 , n75564 );
xor ( n75566 , n75053 , n75229 );
buf ( n75567 , n75566 );
xor ( n75568 , n75132 , n75227 );
buf ( n75569 , n75568 );
xor ( n75570 , n75140 , n75225 );
buf ( n75571 , n75570 );
xor ( n75572 , n75148 , n75223 );
buf ( n75573 , n75572 );
xor ( n75574 , n75156 , n75221 );
buf ( n75575 , n75574 );
xor ( n75576 , n75164 , n75219 );
buf ( n75577 , n75576 );
xor ( n75578 , n75172 , n75217 );
buf ( n75579 , n75578 );
xor ( n75580 , n75180 , n75215 );
buf ( n75581 , n75580 );
xor ( n75582 , n75188 , n75213 );
buf ( n75583 , n75582 );
xor ( n75584 , n75195 , n75211 );
buf ( n75585 , n75584 );
xor ( n75586 , n75201 , n75209 );
buf ( n75587 , n75586 );
xor ( n75588 , n75205 , n75208 );
buf ( n75589 , n75588 );
buf ( n75590 , n75206 );
buf ( n75591 , n75590 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
endmodule
