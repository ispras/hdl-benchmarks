module s5378_bench(
  blif_clk_net,
  blif_reset_net,
  n3065gat,
  n3066gat,
  n3067gat,
  n3068gat,
  n3069gat,
  n3070gat,
  n3071gat,
  n3072gat,
  n3073gat,
  n3074gat,
  n3075gat,
  n3076gat,
  n3077gat,
  n3078gat,
  n3079gat,
  n3080gat,
  n3081gat,
  n3082gat,
  n3083gat,
  n3084gat,
  n3085gat,
  n3086gat,
  n3087gat,
  n3088gat,
  n3089gat,
  n3090gat,
  n3091gat,
  n3092gat,
  n3093gat,
  n3094gat,
  n3095gat,
  n3097gat,
  n3098gat,
  n3099gat,
  n3100gat,
  n3104gat,
  n3105gat,
  n3106gat,
  n3107gat,
  n3108gat,
  n3109gat,
  n3110gat,
  n3111gat,
  n3112gat,
  n3113gat,
  n3114gat,
  n3115gat,
  n3116gat,
  n3117gat,
  n3118gat,
  n3119gat,
  n3120gat,
  n3121gat,
  n3122gat,
  n3123gat,
  n3124gat,
  n3125gat,
  n3126gat,
  n3127gat,
  n3128gat,
  n3129gat,
  n3130gat,
  n3131gat,
  n3132gat,
  n3133gat,
  n3134gat,
  n3135gat,
  n3136gat,
  n3137gat,
  n3138gat,
  n3139gat,
  n3140gat,
  n3141gat,
  n3142gat,
  n3143gat,
  n3144gat,
  n3145gat,
  n3146gat,
  n3147gat,
  n3148gat,
  n3149gat,
  n3150gat,
  n3151gat,
  n3152gat);
input blif_clk_net;
input blif_reset_net;
input n3065gat;
input n3066gat;
input n3067gat;
input n3068gat;
input n3069gat;
input n3070gat;
input n3071gat;
input n3072gat;
input n3073gat;
input n3074gat;
input n3075gat;
input n3076gat;
input n3077gat;
input n3078gat;
input n3079gat;
input n3080gat;
input n3081gat;
input n3082gat;
input n3083gat;
input n3084gat;
input n3085gat;
input n3086gat;
input n3087gat;
input n3088gat;
input n3089gat;
input n3090gat;
input n3091gat;
input n3092gat;
input n3093gat;
input n3094gat;
input n3095gat;
input n3097gat;
input n3098gat;
input n3099gat;
input n3100gat;
output n3104gat;
output n3105gat;
output n3106gat;
output n3107gat;
output n3108gat;
output n3109gat;
output n3110gat;
output n3111gat;
output n3112gat;
output n3113gat;
output n3114gat;
output n3115gat;
output n3116gat;
output n3117gat;
output n3118gat;
output n3119gat;
output n3120gat;
output n3121gat;
output n3122gat;
output n3123gat;
output n3124gat;
output n3125gat;
output n3126gat;
output n3127gat;
output n3128gat;
output n3129gat;
output n3130gat;
output n3131gat;
output n3132gat;
output n3133gat;
output n3134gat;
output n3135gat;
output n3136gat;
output n3137gat;
output n3138gat;
output n3139gat;
output n3140gat;
output n3141gat;
output n3142gat;
output n3143gat;
output n3144gat;
output n3145gat;
output n3146gat;
output n3147gat;
output n3148gat;
output n3149gat;
output n3150gat;
output n3151gat;
output n3152gat;
reg n673gat;
reg n398gat;
reg n402gat;
reg n919gat;
reg n846gat;
reg n2510gat;
reg n271gat;
reg n160gat;
reg n337gat;
reg n842gat;
reg n341gat;
reg n2522gat;
reg n2472gat;
reg n2319gat;
reg n1821gat;
reg n2029gat;
reg n1829gat;
reg n2476gat;
reg n1068gat;
reg n957gat;
reg n861gat;
reg n1294gat;
reg n1241gat;
reg n865gat;
reg n1080gat;
reg n1148gat;
reg n2468gat;
reg n834gat;
reg n707gat;
reg n838gat;
reg n830gat;
reg n614gat;
reg n2526gat;
reg n680gat;
reg n816gat;
reg n580gat;
reg n824gat;
reg n820gat;
reg n883gat;
reg n584gat;
reg n684gat;
reg n699gat;
reg n2464gat;
reg n2399gat;
reg n2343gat;
reg n2203gat;
reg n2562gat;
reg n2207gat;
reg n2626gat;
reg n2490gat;
reg n2622gat;
reg n2630gat;
reg n2543gat;
reg n2102gat;
reg n1880gat;
reg n1763gat;
reg n2155gat;
reg n1035gat;
reg n1121gat;
reg n1072gat;
reg n1282gat;
reg n1226gat;
reg n931gat;
reg n1135gat;
reg n1045gat;
reg n1197gat;
reg n2518gat;
reg n667gat;
reg n659gat;
reg n553gat;
reg n777gat;
reg n561gat;
reg n366gat;
reg n322gat;
reg n318gat;
reg n314gat;
reg n2599gat;
reg n2588gat;
reg n2640gat;
reg n2658gat;
reg n2495gat;
reg n2390gat;
reg n2270gat;
reg n2339gat;
reg n2502gat;
reg n2634gat;
reg n2506gat;
reg n1834gat;
reg n1767gat;
reg n2084gat;
reg n2143gat;
reg n2061gat;
reg n2139gat;
reg n1899gat;
reg n1850gat;
reg n2403gat;
reg n2394gat;
reg n2440gat;
reg n2407gat;
reg n2347gat;
reg n1389gat;
reg n2021gat;
reg n1394gat;
reg n1496gat;
reg n2091gat;
reg n1332gat;
reg n1740gat;
reg n2179gat;
reg n2190gat;
reg n2135gat;
reg n2262gat;
reg n2182gat;
reg n1433gat;
reg n1316gat;
reg n1363gat;
reg n1312gat;
reg n1775gat;
reg n1871gat;
reg n2592gat;
reg n1508gat;
reg n1678gat;
reg n2309gat;
reg n2450gat;
reg n2446gat;
reg n2095gat;
reg n2176gat;
reg n2169gat;
reg n2454gat;
reg n2040gat;
reg n2044gat;
reg n2037gat;
reg n2025gat;
reg n2099gat;
reg n2266gat;
reg n2033gat;
reg n2110gat;
reg n2125gat;
reg n2121gat;
reg n2117gat;
reg n1975gat;
reg n2644gat;
reg n156gat;
reg n152gat;
reg n331gat;
reg n388gat;
reg n463gat;
reg n327gat;
reg n384gat;
reg n256gat;
reg n470gat;
reg n148gat;
reg n2458gat;
reg n2514gat;
reg n1771gat;
reg n1336gat;
reg n1748gat;
reg n1675gat;
reg n1807gat;
reg n1340gat;
reg n1456gat;
reg n1525gat;
reg n1462gat;
reg n1596gat;
reg n1588gat;
wire n43gat;
wire n1967gat;
wire II1344;
wire n911gat;
wire n2167gat;
wire n2612gat;
wire n1706gat;
wire n419gat;
wire n1724gat;
wire II4690;
wire II476;
wire II4518;
wire II880;
wire n3044gat;
wire n2791gat;
wire n221gat;
wire II2915;
wire n1202gat;
wire II1416;
wire n588gat;
wire II2232;
wire n1358gat;
wire n974gat;
wire n194gat;
wire n702gat;
wire n696gat;
wire n1719gat;
wire n443gat;
wire n952gat;
wire II4783;
wire n2577gat;
wire n499gat;
wire n1175gat;
wire n2023gat;
wire II4212;
wire n1790gat;
wire n1656gat;
wire II2394;
wire n2845gat;
wire n1225gat;
wire II2344;
wire n1172gat;
wire n63gat;
wire n878gat;
wire n2050gat;
wire n17gat;
wire n2683gat;
wire n2746gat;
wire n782gat;
wire II2263;
wire n2655gat;
wire n2661gat;
wire n757gat;
wire n1303gat;
wire n2652gat;
wire n1002gat;
wire n2850gat;
wire n1291gat;
wire n2607gat;
wire n721gat;
wire n2418gat;
wire n1219gat;
wire n2621gat;
wire n2433gat;
wire n786gat;
wire n1050gat;
wire n3001gat;
wire II2934;
wire II985;
wire II437;
wire II227;
wire n1008gat;
wire II4699;
wire II1007;
wire n1584gat;
wire II4777;
wire II846;
wire n813gat;
wire n632gat;
wire n2832gat;
wire II726;
wire n2046gat;
wire n1215gat;
wire n1423gat;
wire n1361gat;
wire n2488gat;
wire n508gat;
wire II1708;
wire n2942gat;
wire n2355gat;
wire n1212gat;
wire II4642;
wire II3509;
wire n1161gat;
wire n2223gat;
wire n410gat;
wire II2847;
wire n746gat;
wire II2385;
wire n766gat;
wire II2324;
wire n1701gat;
wire n2741gat;
wire n960gat;
wire n1221gat;
wire n2913gat;
wire n2452gat;
wire n386gat;
wire II3342;
wire n2186gat;
wire n351gat;
wire n2237gat;
wire n1606gat;
wire n2243gat;
wire n1444gat;
wire n212gat;
wire n955gat;
wire n136gat;
wire n1480gat;
wire n2944gat;
wire n2694gat;
wire n1670gat;
wire n1694gat;
wire n2151gat;
wire n3019gat;
wire n1163gat;
wire II3954;
wire II1067;
wire II311;
wire II2885;
wire n2149gat;
wire n2733gat;
wire n855gat;
wire n1174gat;
wire n1164gat;
wire n2486gat;
wire II4657;
wire n688gat;
wire n1838gat;
wire n910gat;
wire n2749gat;
wire n2860gat;
wire n490gat;
wire n1792gat;
wire n2421gat;
wire n127gat;
wire II1360;
wire n2852gat;
wire n1263gat;
wire n959gat;
wire n1729gat;
wire n2702gat;
wire II359;
wire n1448gat;
wire n2863gat;
wire II3923;
wire II512;
wire n2500gat;
wire n1555gat;
wire n646gat;
wire n692gat;
wire n2325gat;
wire n1532gat;
wire n2148gat;
wire n1502gat;
wire n1014gat;
wire n453gat;
wire II4429;
wire n925gat;
wire II2153;
wire II4135;
wire n2910gat;
wire II149;
wire n1104gat;
wire n2672gat;
wire II2084;
wire n1859gat;
wire n1945gat;
wire n1619gat;
wire n2660gat;
wire n2689gat;
wire n1548gat;
wire II3235;
wire n996gat;
wire n2795gat;
wire n1989gat;
wire n923gat;
wire II2242;
wire n1193gat;
wire n947gat;
wire n2693gat;
wire II4217;
wire n857gat;
wire n2986gat;
wire II2831;
wire n1879gat;
wire n40gat;
wire II111;
wire n2238gat;
wire n779gat;
wire n756gat;
wire n1878gat;
wire n1550gat;
wire n2449gat;
wire n219gat;
wire n1067gat;
wire n1173gat;
wire II4792;
wire n1925gat;
wire n1223gat;
wire n277gat;
wire II902;
wire n1330gat;
wire n2534gat;
wire n415gat;
wire n907gat;
wire n3009gat;
wire n683gat;
wire n370gat;
wire n513gat;
wire n874gat;
wire n2814gat;
wire n178gat;
wire n2052gat;
wire n2709gat;
wire n2133gat;
wire II4475;
wire n2213gat;
wire n2955gat;
wire n22gat;
wire n807gat;
wire II62;
wire n990gat;
wire n2018gat;
wire n1309gat;
wire II583;
wire n653gat;
wire II2174;
wire n875gat;
wire n733gat;
wire n523gat;
wire n2932gat;
wire n53gat;
wire n1524gat;
wire n1485gat;
wire n3036gat;
wire n1324gat;
wire n1887gat;
wire n247gat;
wire II3691;
wire II1082;
wire n1099gat;
wire n1123gat;
wire n172gat;
wire n1270gat;
wire n1690gat;
wire II4687;
wire n2939gat;
wire n916gat;
wire II637;
wire II3143;
wire n1610gat;
wire n3045gat;
wire n1636gat;
wire n1436gat;
wire n2128gat;
wire n2697gat;
wire n1495gat;
wire n1214gat;
wire n880gat;
wire II97;
wire n2553gat;
wire II65;
wire n649gat;
wire n992gat;
wire n1095gat;
wire n1115gat;
wire n1917gat;
wire n573gat;
wire n2350gat;
wire n1551gat;
wire n1015gat;
wire II320;
wire n2456gat;
wire n2035gat;
wire II842;
wire II721;
wire n1613gat;
wire n1158gat;
wire II4660;
wire n899gat;
wire II395;
wire n2753gat;
wire II1724;
wire n2775gat;
wire II4489;
wire II220;
wire n2962gat;
wire n1788gat;
wire n71gat;
wire n270gat;
wire n748gat;
wire n1271gat;
wire II4309;
wire n1441gat;
wire II3867;
wire n1420gat;
wire n1479gat;
wire n1483gat;
wire n520gat;
wire n267gat;
wire n1685gat;
wire n2269gat;
wire II2044;
wire II2035;
wire II4499;
wire n507gat;
wire n1662gat;
wire II4630;
wire n2777gat;
wire n1605gat;
wire II4020;
wire n775gat;
wire n2981gat;
wire n809gat;
wire n769gat;
wire n930gat;
wire n635gat;
wire II3394;
wire n1096gat;
wire n2948gat;
wire II340;
wire n571gat;
wire n2115gat;
wire n1382gat;
wire n3047gat;
wire n864gat;
wire n2591gat;
wire n926gat;
wire n897gat;
wire n293gat;
wire n2907gat;
wire II4389;
wire n344gat;
wire II678;
wire n986gat;
wire n1326gat;
wire n170gat;
wire n1955gat;
wire II4723;
wire II378;
wire n253gat;
wire n2539gat;
wire II3387;
wire n783gat;
wire n1934gat;
wire n175gat;
wire n1960gat;
wire II1723;
wire n694gat;
wire n983gat;
wire n1023gat;
wire II253;
wire n1393gat;
wire n144gat;
wire n2637gat;
wire n2359gat;
wire n3017gat;
wire n771gat;
wire n2908gat;
wire n1920gat;
wire n2216gat;
wire n582gat;
wire n2789gat;
wire n56gat;
wire n679gat;
wire II456;
wire n502gat;
wire n204gat;
wire II4412;
wire n2547gat;
wire II1374;
wire II363;
wire n1836gat;
wire n2487gat;
wire n647gat;
wire n1250gat;
wire II4732;
wire n2896gat;
wire n2613gat;
wire n1845gat;
wire n794gat;
wire n691gat;
wire n1842gat;
wire n1602gat;
wire n2079gat;
wire n2959gat;
wire II440;
wire n1007gat;
wire n1417gat;
wire n1563gat;
wire n709gat;
wire II837;
wire II199;
wire n1666gat;
wire n2735gat;
wire n1580gat;
wire n1519gat;
wire II1201;
wire n1077gat;
wire n2212gat;
wire n2009gat;
wire II980;
wire n2388gat;
wire n1734gat;
wire n591gat;
wire n921gat;
wire n2516gat;
wire n1866gat;
wire n933gat;
wire n793gat;
wire n1974gat;
wire n229gat;
wire n2919gat;
wire n2259gat;
wire II2812;
wire n182gat;
wire n879gat;
wire n3028gat;
wire II92;
wire n2917gat;
wire n812gat;
wire n2877gat;
wire n969gat;
wire n2794gat;
wire n1113gat;
wire n2662gat;
wire II1927;
wire n2992gat;
wire n167gat;
wire n1373gat;
wire II3504;
wire n1112gat;
wire n705gat;
wire n273gat;
wire n47gat;
wire n2604gat;
wire n1737gat;
wire n1179gat;
wire II3312;
wire n343gat;
wire n3013gat;
wire n111gat;
wire II620;
wire n2605gat;
wire n2731gat;
wire n828gat;
wire II480;
wire II4654;
wire n1978gat;
wire n244gat;
wire n2357gat;
wire n2880gat;
wire II2721;
wire n1963gat;
wire II5;
wire n662gat;
wire n11gat;
wire n2257gat;
wire n1574gat;
wire n334gat;
wire n1884gat;
wire II3742;
wire n1700gat;
wire II2225;
wire n773gat;
wire n189gat;
wire n2858gat;
wire n2215gat;
wire II2389;
wire n1199gat;
wire II3713;
wire n2934gat;
wire II423;
wire II1236;
wire n2969gat;
wire II2832;
wire II4372;
wire n1696gat;
wire n2696gat;
wire n1097gat;
wire n2881gat;
wire II3297;
wire n1415gat;
wire n891gat;
wire n979gat;
wire n1006gat;
wire n1054gat;
wire n1279gat;
wire II2014;
wire n2439gat;
wire n1970gat;
wire n1564gat;
wire n1082gat;
wire n1994gat;
wire n1839gat;
wire n290gat;
wire n2210gat;
wire II1411;
wire n645gat;
wire n2422gat;
wire n447gat;
wire n3002gat;
wire n2201gat;
wire n1818gat;
wire n2869gat;
wire n1786gat;
wire n1484gat;
wire n1231gat;
wire n38gat;
wire n1277gat;
wire n2820gat;
wire n792gat;
wire n2205gat;
wire n199gat;
wire n147gat;
wire n1409gat;
wire II977;
wire n2960gat;
wire n295gat;
wire n2798gat;
wire II1516;
wire n439gat;
wire n1024gat;
wire n1954gat;
wire n510gat;
wire n1287gat;
wire n2941gat;
wire n1603gat;
wire n2429gat;
wire n2965gat;
wire n1684gat;
wire n2185gat;
wire n479gat;
wire II877;
wire n2829gat;
wire n246gat;
wire n2878gat;
wire n2752gat;
wire n2101gat;
wire n2146gat;
wire n961gat;
wire II3315;
wire n1000gat;
wire II1439;
wire n1421gat;
wire n1247gat;
wire n2957gat;
wire n2575gat;
wire n196gat;
wire n2952gat;
wire n501gat;
wire n2671gat;
wire n262gat;
wire n2916gat;
wire n1533gat;
wire n1152gat;
wire II4717;
wire II23;
wire n3040gat;
wire n1266gat;
wire n1918gat;
wire n2681gat;
wire II3148;
wire n1798gat;
wire II712;
wire n312gat;
wire n2692gat;
wire n2162gat;
wire n64gat;
wire n1762gat;
wire II1035;
wire n2894gat;
wire n228gat;
wire n978gat;
wire n2150gat;
wire n1787gat;
wire n2853gat;
wire n689gat;
wire II3801;
wire n240gat;
wire n2883gat;
wire n2413gat;
wire n1888gat;
wire II2953;
wire n2430gat;
wire n729gat;
wire II259;
wire n965gat;
wire II337;
wire n521gat;
wire II1476;
wire n1075gat;
wire n1609gat;
wire II2181;
wire n2718gat;
wire n968gat;
wire n79gat;
wire II206;
wire n1334gat;
wire n2674gat;
wire II4678;
wire n989gat;
wire n128gat;
wire n2564gat;
wire n2342gat;
wire n141gat;
wire n1861gat;
wire II4626;
wire n1185gat;
wire n741gat;
wire n526gat;
wire n1468gat;
wire n1305gat;
wire n2387gat;
wire n975gat;
wire n356gat;
wire n2286gat;
wire n795gat;
wire n1105gat;
wire n2923gat;
wire n181gat;
wire n1778gat;
wire II1894;
wire n405gat;
wire n1530gat;
wire n2793gat;
wire n732gat;
wire n2570gat;
wire II675;
wire n803gat;
wire II2316;
wire n1769gat;
wire n2292gat;
wire II2040;
wire n76gat;
wire II4747;
wire II4485;
wire n2574gat;
wire n2603gat;
wire n2874gat;
wire n1500gat;
wire II3056;
wire n324gat;
wire n1018gat;
wire II634;
wire n1372gat;
wire n498gat;
wire n3018gat;
wire n62gat;
wire n1642gat;
wire n2949gat;
wire n2338gat;
wire n2688gat;
wire n808gat;
wire n2904gat;
wire n800gat;
wire n1849gat;
wire n1378gat;
wire n2673gat;
wire n2548gat;
wire II812;
wire n814gat;
wire n1369gat;
wire n2470gat;
wire II4623;
wire n1471gat;
wire II2109;
wire II2177;
wire n2199gat;
wire II4194;
wire II3513;
wire II3831;
wire II1115;
wire n2719gat;
wire n1264gat;
wire n1447gat;
wire n2809gat;
wire n2392gat;
wire n1055gat;
wire II1243;
wire II999;
wire n145gat;
wire II473;
wire n739gat;
wire n1280gat;
wire II2837;
wire n2042gat;
wire n2805gat;
wire II4023;
wire n34gat;
wire n3054gat;
wire n82gat;
wire II1174;
wire n1244gat;
wire n249gat;
wire n2253gat;
wire n818gat;
wire n2891gat;
wire n289gat;
wire n1546gat;
wire II1807;
wire n382gat;
wire n2953gat;
wire n565gat;
wire n759gat;
wire n2747gat;
wire n1201gat;
wire n287gat;
wire n1239gat;
wire n909gat;
wire n1608gat;
wire n1855gat;
wire n2317gat;
wire II4530;
wire II1138;
wire n1446gat;
wire n2677gat;
wire n737gat;
wire n1431gat;
wire n2402gat;
wire n1160gat;
wire n1159gat;
wire n2252gat;
wire II4753;
wire n392gat;
wire n948gat;
wire II4105;
wire II3412;
wire n1070gat;
wire n2862gat;
wire n1232gat;
wire n3011gat;
wire n1017gat;
wire n2925gat;
wire n1705gat;
wire II1248;
wire n51gat;
wire n677gat;
wire n1773gat;
wire n2924gat;
wire n2895gat;
wire n664gat;
wire II851;
wire n1091gat;
wire II936;
wire n1359gat;
wire II1121;
wire n2921gat;
wire n1707gat;
wire n1794gat;
wire n3062gat;
wire II2400;
wire n354gat;
wire n84gat;
wire n743gat;
wire II2890;
wire II230;
wire n1819gat;
wire n1571gat;
wire n69gat;
wire n1738gat;
wire n1699gat;
wire n888gat;
wire n938gat;
wire n776gat;
wire II1399;
wire n2727gat;
wire II3303;
wire II300;
wire n1253gat;
wire n2899gat;
wire n524gat;
wire II2145;
wire n2734gat;
wire n517gat;
wire n2840gat;
wire n578gat;
wire n3059gat;
wire n2843gat;
wire n840gat;
wire n2354gat;
wire n1216gat;
wire n3057gat;
wire n2436gat;
wire n1507gat;
wire n1760gat;
wire n1543gat;
wire n1590gat;
wire II3765;
wire n954gat;
wire II1899;
wire n2405gat;
wire n2897gat;
wire n143gat;
wire II443;
wire II834;
wire n2785gat;
wire n2937gat;
wire n1235gat;
wire II1683;
wire n1677gat;
wire n2758gat;
wire n1051gat;
wire II426;
wire II3891;
wire n949gat;
wire n44gat;
wire II1031;
wire n2763gat;
wire n2704gat;
wire II3465;
wire n735gat;
wire n2926gat;
wire n333gat;
wire n987gat;
wire n2048gat;
wire n2406gat;
wire n3060gat;
wire n231gat;
wire n1189gat;
wire II4554;
wire n929gat;
wire II815;
wire n829gat;
wire n1598gat;
wire n503gat;
wire n2572gat;
wire II4349;
wire n1311gat;
wire n620gat;
wire n1968gat;
wire II1402;
wire n1248gat;
wire n1717gat;
wire II30;
wire n634gat;
wire II1481;
wire n408gat;
wire n1742gat;
wire n1114gat;
wire II1155;
wire n2988gat;
wire II958;
wire n1757gat;
wire n321gat;
wire n1593gat;
wire n1505gat;
wire n150gat;
wire n1269gat;
wire n59gat;
wire n1031gat;
wire n1101gat;
wire n1059gat;
wire n1487gat;
wire n863gat;
wire n3000gat;
wire n329gat;
wire n2819gat;
wire n2202gat;
wire n459gat;
wire n1567gat;
wire II1023;
wire n3037gat;
wire n2158gat;
wire n1411gat;
wire n3023gat;
wire n2189gat;
wire II368;
wire n767gat;
wire n484gat;
wire n1338gat;
wire n1630gat;
wire n2781gat;
wire n164gat;
wire n200gat;
wire n760gat;
wire n877gat;
wire n1182gat;
wire n2695gat;
wire n1629gat;
wire II1999;
wire II4524;
wire n2956gat;
wire n2601gat;
wire n1576gat;
wire II4332;
wire n2060gat;
wire n2738gat;
wire n1011gat;
wire n2002gat;
wire n2595gat;
wire n1557gat;
wire n420gat;
wire II1;
wire n1318gat;
wire II4506;
wire n195gat;
wire n1647gat;
wire n2767gat;
wire n2097gat;
wire II1786;
wire n2625gat;
wire n1710gat;
wire n142gat;
wire II4798;
wire n1566gat;
wire n1016gat;
wire n2493gat;
wire n1783gat;
wire n2432gat;
wire n2868gat;
wire n1357gat;
wire n1490gat;
wire n2211gat;
wire n264gat;
wire II734;
wire n1614gat;
wire n3063gat;
wire II1496;
wire n2964gat;
wire II863;
wire n1624gat;
wire n2410gat;
wire n1923gat;
wire n1403gat;
wire II3904;
wire n1268gat;
wire II1791;
wire n2760gat;
wire n2682gat;
wire n2284gat;
wire n92gat;
wire II1923;
wire n2779gat;
wire n1274gat;
wire n576gat;
wire n1846gat;
wire n1257gat;
wire n2855gat;
wire n2750gat;
wire n197gat;
wire n1782gat;
wire n514gat;
wire II2873;
wire II1874;
wire n1618gat;
wire n421gat;
wire II4222;
wire n1732gat;
wire n1556gat;
wire n325gat;
wire n355gat;
wire n509gat;
wire n2836gat;
wire n469gat;
wire n1414gat;
wire II3882;
wire II776;
wire II651;
wire II76;
wire n2699gat;
wire n2220gat;
wire n1587gat;
wire n736gat;
wire n468gat;
wire n2414gat;
wire n2931gat;
wire n1155gat;
wire II2213;
wire II4681;
wire n815gat;
wire n449gat;
wire n2291gat;
wire n587gat;
wire II749;
wire n1356gat;
wire II381;
wire n738gat;
wire n1714gat;
wire II1833;
wire n2736gat;
wire n49gat;
wire n2670gat;
wire II1961;
wire n1578gat;
wire n789gat;
wire n656gat;
wire n2345gat;
wire II240;
wire n2668gat;
wire n2890gat;
wire n1774gat;
wire n184gat;
wire n1207gat;
wire II4580;
wire n1350gat;
wire n2073gat;
wire n2332gat;
wire n1726gat;
wire n2780gat;
wire n1306gat;
wire n943gat;
wire II3336;
wire n1921gat;
wire n1260gat;
wire n266gat;
wire n476gat;
wire n849gat;
wire n313gat;
wire II1488;
wire II1348;
wire II2672;
wire n1200gat;
wire n423gat;
wire II1464;
wire II4768;
wire n1004gat;
wire II1472;
wire n397gat;
wire II3178;
wire n1460gat;
wire n377gat;
wire n1581gat;
wire II1085;
wire n2823gat;
wire n1103gat;
wire n1595gat;
wire II1857;
wire n2936gat;
wire n2124gat;
wire II1339;
wire n380gat;
wire n86gat;
wire n2401gat;
wire n1653gat;
wire II2433;
wire n1208gat;
wire n2846gat;
wire n362gat;
wire n2905gat;
wire n1367gat;
wire n678gat;
wire II4774;
wire n2246gat;
wire n2397gat;
wire n396gat;
wire II2254;
wire n1929gat;
wire n2751gat;
wire II1584;
wire n939gat;
wire n1328gat;
wire n2826gat;
wire n1800gat;
wire n1211gat;
wire II3300;
wire II351;
wire II3290;
wire n2554gat;
wire n1302gat;
wire n2861gat;
wire n1228gat;
wire n2650gat;
wire n981gat;
wire n806gat;
wire II715;
wire n2195gat;
wire n2492gat;
wire n984gat;
wire n2892gat;
wire n2426gat;
wire n2792gat;
wire n461gat;
wire II4145;
wire II4573;
wire n1988gat;
wire n712gat;
wire n506gat;
wire II3948;
wire II2720;
wire n1523gat;
wire n2545gat;
wire n407gat;
wire n1186gat;
wire n752gat;
wire n2283gat;
wire n687gat;
wire II2417;
wire n903gat;
wire II796;
wire n1366gat;
wire n1028gat;
wire n2730gat;
wire n1368gat;
wire II3494;
wire II4352;
wire n1669gat;
wire n269gat;
wire n2724gat;
wire n2576gat;
wire II237;
wire n2691gat;
wire II1515;
wire n630gat;
wire n2967gat;
wire n785gat;
wire II1209;
wire n1553gat;
wire II4409;
wire n1001gat;
wire n2293gat;
wire n3014gat;
wire n906gat;
wire n2147gat;
wire n1607gat;
wire n361gat;
wire n867gat;
wire n2206gat;
wire n1562gat;
wire n177gat;
wire II2731;
wire n455gat;
wire n2797gat;
wire n1599gat;
wire n1083gat;
wire n512gat;
wire n1641gat;
wire II3941;
wire n2762gat;
wire II1322;
wire n1827gat;
wire n2737gat;
wire n1898gat;
wire n2460gat;
wire n1673gat;
wire n1922gat;
wire n255gat;
wire n1632gat;
wire n1785gat;
wire n2520gat;
wire II1630;
wire n294gat;
wire n2163gat;
wire n2830gat;
wire n2615gat;
wire n2768gat;
wire n924gat;
wire n633gat;
wire n291gat;
wire II3539;
wire n1869gat;
wire n1840gat;
wire n1865gat;
wire II1336;
wire n1646gat;
wire n1568gat;
wire n373gat;
wire n966gat;
wire n1549gat;
wire n1841gat;
wire n583gat;
wire n1709gat;
wire n485gat;
wire n522gat;
wire II4756;
wire n701gat;
wire n2686gat;
wire n2996gat;
wire n1379gat;
wire II282;
wire n187gat;
wire n2027gat;
wire n35gat;
wire n2141gat;
wire n2642gat;
wire n1635gat;
wire n2893gat;
wire II790;
wire n1686gat;
wire n1651gat;
wire n853gat;
wire n1205gat;
wire n928gat;
wire n1466gat;
wire n1897gat;
wire II4496;
wire n1736gat;
wire II4122;
wire n1467gat;
wire n1961gat;
wire n3015gat;
wire n2130gat;
wire n444gat;
wire II4789;
wire n448gat;
wire n915gat;
wire n1721gat;
wire n1806gat;
wire II50;
wire n881gat;
wire n2337gat;
wire n2947gat;
wire n1285gat;
wire n2008gat;
wire n1183gat;
wire II3621;
wire n1419gat;
wire n2918gat;
wire n1249gat;
wire n651gat;
wire n2728gat;
wire n406gat;
wire n369gat;
wire n956gat;
wire n788gat;
wire n1019gat;
wire II1667;
wire II4478;
wire n1894gat;
wire n3049gat;
wire n2427gat;
wire n2886gat;
wire n2417gat;
wire n1831gat;
wire n452gat;
wire n1365gat;
wire n625gat;
wire n3042gat;
wire n1780gat;
wire n2679gat;
wire n1424gat;
wire n2053gat;
wire n1486gat;
wire n1314gat;
wire n1723gat;
wire II4684;
wire n1351gat;
wire n1442gat;
wire n1520gat;
wire n3020gat;
wire II1255;
wire n586gat;
wire II3957;
wire n2629gat;
wire n222gat;
wire II4726;
wire n2632gat;
wire II3635;
wire n1408gat;
wire n2684gat;
wire n2582gat;
wire n1482gat;
wire n2578gat;
wire n400gat;
wire n2244gat;
wire n850gat;
wire n393gat;
wire n1374gat;
wire n3025gat;
wire II1795;
wire n2483gat;
wire n1754gat;
wire II2049;
wire n1153gat;
wire n1315gat;
wire n856gat;
wire II4227;
wire n1969gat;
wire n774gat;
wire II3520;
wire n2200gat;
wire n2055gat;
wire n263gat;
wire n345gat;
wire II1002;
wire n555gat;
wire n2815gat;
wire n2938gat;
wire II4329;
wire II3339;
wire n1882gat;
wire n2057gat;
wire II672;
wire n1352gat;
wire n1416gat;
wire n2841gat;
wire II3808;
wire n375gat;
wire n2571gat;
wire n666gat;
wire n1320gat;
wire n2616gat;
wire n3035gat;
wire n2933gat;
wire n1458gat;
wire n2131gat;
wire n1259gat;
wire n1010gat;
wire n2987gat;
wire n2193gat;
wire II243;
wire n563gat;
wire n1376gat;
wire n89gat;
wire n1848gat;
wire n1348gat;
wire n1727gat;
wire n78gat;
wire n2129gat;
wire n1308gat;
wire n2054gat;
wire II4024;
wire n1134gat;
wire n2218gat;
wire II698;
wire n2776gat;
wire n1060gat;
wire n1428gat;
wire n1052gat;
wire n1392gat;
wire n2783gat;
wire n2885gat;
wire n1251gat;
wire n2983gat;
wire n1625gat;
wire n976gat;
wire n364gat;
wire n944gat;
wire n905gat;
wire n2194gat;
wire n819gat;
wire n169gat;
wire n73gat;
wire n1816gat;
wire n2804gat;
wire n574gat;
wire n2565gat;
wire II317;
wire n1412gat;
wire n274gat;
wire n1111gat;
wire n1310gat;
wire n1236gat;
wire II899;
wire n1972gat;
wire II4666;
wire n848gat;
wire n226gat;
wire II4067;
wire n2423gat;
wire n230gat;
wire II44;
wire II2238;
wire n188gat;
wire n2597gat;
wire n690gat;
wire n2610gat;
wire n2847gat;
wire n1889gat;
wire n2556gat;
wire n3056gat;
wire n927gat;
wire II4651;
wire II2428;
wire n551gat;
wire n871gat;
wire n180gat;
wire n2499gat;
wire n223gat;
wire n42gat;
wire n1573gat;
wire n2609gat;
wire n572gat;
wire n2844gat;
wire n414gat;
wire n2982gat;
wire n1703gat;
wire n997gat;
wire II4720;
wire II1216;
wire n39gat;
wire n710gat;
wire n235gat;
wire n993gat;
wire n519gat;
wire n1301gat;
wire n1387gat;
wire II572;
wire n357gat;
wire II3754;
wire n353gat;
wire II2017;
wire n1430gat;
wire n2990gat;
wire n1494gat;
wire n589gat;
wire II921;
wire n2951gat;
wire n1090gat;
wire n964gat;
wire n2740gat;
wire n1094gat;
wire II3174;
wire n751gat;
wire n2930gat;
wire II941;
wire n1528gat;
wire n2596gat;
wire n2537gat;
wire n1674gat;
wire n1671gat;
wire n1973gat;
wire n885gat;
wire II591;
wire n52gat;
wire n65gat;
wire n962gat;
wire II4702;
wire n1722gat;
wire II4744;
wire n2867gat;
wire n2602gat;
wire n2748gat;
wire n1087gat;
wire II3149;
wire II4452;
wire n1864gat;
wire n988gat;
wire n1210gat;
wire n1781gat;
wire n896gat;
wire n2766gat;
wire II1783;
wire II1908;
wire n750gat;
wire n2352gat;
wire II4669;
wire n460gat;
wire n1400gat;
wire II3191;
wire n590gat;
wire II768;
wire II1436;
wire n2729gat;
wire n638gat;
wire n1498gat;
wire n2812gat;
wire II3211;
wire n1281gat;
wire n2573gat;
wire n446gat;
wire II171;
wire II771;
wire II1467;
wire II2989;
wire n1120gat;
wire n2946gat;
wire n1617gat;
wire n441gat;
wire II1407;
wire n2903gat;
wire n2014gat;
wire n50gat;
wire n2633gat;
wire n2531gat;
wire n3050gat;
wire n1029gat;
wire n3003gat;
wire n2985gat;
wire n1150gat;
wire n2119gat;
wire n753gat;
wire n1117gat;
wire II2032;
wire n1450gat;
wire II741;
wire n2419gat;
wire n2389gat;
wire n2197gat;
wire n2541gat;
wire n893gat;
wire n297gat;
wire n282gat;
wire II858;
wire n1100gat;
wire n2720gat;
wire n1477gat;
wire n762gat;
wire n913gat;
wire II409;
wire II2112;
wire II1538;
wire n2646gat;
wire II2696;
wire II4672;
wire II1891;
wire II3951;
wire n365gat;
wire II4449;
wire n3055gat;
wire n1410gat;
wire n890gat;
wire n1246gat;
wire n2808gat;
wire n2011gat;
wire n1234gat;
wire n2909gat;
wire II2257;
wire n886gat;
wire n2557gat;
wire n2217gat;
wire n852gat;
wire n1461gat;
wire n991gat;
wire n629gat;
wire n168gat;
wire n1157gat;
wire n451gat;
wire n860gat;
wire II4432;
wire n2363gat;
wire n2219gat;
wire n2667gat;
wire n1919gat;
wire n2725gat;
wire n1643gat;
wire n162gat;
wire n1203gat;
wire II4108;
wire n2732gat;
wire II4117;
wire II4000;
wire n1151gat;
wire n1860gat;
wire n2560gat;
wire n1777gat;
wire n1521gat;
wire II1996;
wire n134gat;
wire n2687gat;
wire II4765;
wire II1719;
wire n2428gat;
wire n648gat;
wire II414;
wire II264;
wire II420;
wire n1147gat;
wire n1893gat;
wire n1089gat;
wire n755gat;
wire n1162gat;
wire n2538gat;
wire n1558gat;
wire n1402gat;
wire II1124;
wire n2482gat;
wire n48gat;
wire n2639gat;
wire n2997gat;
wire II3703;
wire n1559gat;
wire n158gat;
wire n2214gat;
wire n1252gat;
wire n2282gat;
wire n2385gat;
wire II4735;
wire n804gat;
wire n898gat;
wire n1791gat;
wire n811gat;
wire II3306;
wire n922gat;
wire II3273;
wire n1577gat;
wire II3461;
wire n876gat;
wire II4216;
wire n292gat;
wire n2159gat;
wire II1079;
wire n2261gat;
wire n1154gat;
wire II2130;
wire n13gat;
wire n2665gat;
wire n2184gat;
wire n2620gat;
wire II1028;
wire n2137gat;
wire n2707gat;
wire n2349gat;
wire n2384gat;
wire II1769;
wire n1891gat;
wire n72gat;
wire n2580gat;
wire n715gat;
wire n731gat;
wire n1655gat;
wire n2606gat;
wire n336gat;
wire n2530gat;
wire n1513gat;
wire n2579gat;
wire n2945gat;
wire n2786gat;
wire n278gat;
wire II1230;
wire n241gat;
wire n2935gat;
wire n2409gat;
wire n2818gat;
wire II1091;
wire II1204;
wire n1779gat;
wire n3034gat;
wire II683;
wire n640gat;
wire II642;
wire n917gat;
wire n1043gat;
wire n146gat;
wire n2664gat;
wire n1586gat;
wire n1439gat;
wire n2744gat;
wire n2974gat;
wire n1885gat;
wire n2966gat;
wire n2828gat;
wire II178;
wire n643gat;
wire n418gat;
wire n457gat;
wire n445gat;
wire n2249gat;
wire n2168gat;
wire n122gat;
wire n1554gat;
wire n1278gat;
wire n67gat;
wire II331;
wire n982gat;
wire n2132gat;
wire n173gat;
wire n1958gat;
wire n2255gat;
wire n1381gat;
wire n728gat;
wire n1592gat;
wire II729;
wire n754gat;
wire n637gat;
wire n2722gat;
wire n1681gat;
wire n347gat;
wire II4620;
wire n934gat;
wire n68gat;
wire n1660gat;
wire II2403;
wire n494gat;
wire n1957gat;
wire n892gat;
wire n1025gat;
wire n1759gat;
wire n346gat;
wire n658gat;
wire II4129;
wire II3677;
wire n2078gat;
wire n2922gat;
wire n2082gat;
wire n3064gat;
wire n493gat;
wire II4714;
wire n617gat;
wire n963gat;
wire n2705gat;
wire n1823gat;
wire n2416gat;
wire II4548;
wire n2743gat;
wire II579;
wire n372gat;
wire n970gat;
wire n2504gat;
wire n1012gat;
wire II2735;
wire n46gat;
wire n422gat;
wire n2059gat;
wire II203;
wire n1435gat;
wire n1116gat;
wire n1863gat;
wire n568gat;
wire n234gat;
wire n3032gat;
wire n1102gat;
wire n1634gat;
wire n745gat;
wire n3006gat;
wire n1935gat;
wire n716gat;
wire n2536gat;
wire II4536;
wire n2950gat;
wire n121gat;
wire n2778gat;
wire n3030gat;
wire n3010gat;
wire n1529gat;
wire n2443gat;
wire n259gat;
wire II1166;
wire II1585;
wire n2993gat;
wire II1837;
wire n2480gat;
wire n159gat;
wire II2813;
wire II1453;
wire n2494gat;
wire n1591gat;
wire II4705;
wire n1353gat;
wire n530gat;
wire n2984gat;
wire II4512;
wire II1319;
wire n2016gat;
wire n3004gat;
wire n764gat;
wire n945gat;
wire n810gat;
wire II81;
wire n1765gat;
wire n2726gat;
wire n1713gat;
wire n2353gat;
wire II248;
wire n120gat;
wire n3027gat;
wire n1451gat;
wire n1399gat;
wire n1220gat;
wire n1693gat;
wire n887gat;
wire II4663;
wire II3179;
wire n2739gat;
wire n3043gat;
wire n805gat;
wire n655gat;
wire II278;
wire n496gat;
wire n2811gat;
wire II4081;
wire n1725gat;
wire n3052gat;
wire II4594;
wire n260gat;
wire n594gat;
wire n577gat;
wire n2822gat;
wire n532gat;
wire n631gat;
wire n2717gat;
wire n1254gat;
wire n130gat;
wire n1354gat;
wire II930;
wire n125gat;
wire n1986gat;
wire n1886gat;
wire II1860;
wire n1565gat;
wire n3053gat;
wire n516gat;
wire II406;
wire n2821gat;
wire n477gat;
wire II1278;
wire n2649gat;
wire II1227;
wire n1718gat;
wire n740gat;
wire n481gat;
wire n1476gat;
wire n791gat;
wire n1615gat;
wire II746;
wire II4144;
wire n12gat;
wire n139gat;
wire n2174gat;
wire n765gat;
wire n1053gat;
wire n1924gat;
wire n2991gat;
wire n1377gat;
wire II1877;
wire n2663gat;
wire II446;
wire n2712gat;
wire n2998gat;
wire II2380;
wire II398;
wire n1322gat;
wire n747gat;
wire n951gat;
wire n2358gat;
wire II1493;
wire n3039gat;
wire n946gat;
wire II1251;
wire n2810gat;
wire n686gat;
wire n1222gat;
wire n1999gat;
wire n2093gat;
wire n1418gat;
wire II100;
wire II576;
wire n935gat;
wire II4786;
wire n1323gat;
wire n1398gat;
wire n593gat;
wire n941gat;
wire n1704gat;
wire n1501gat;
wire n980gat;
wire n2558gat;
wire n2329gat;
wire n2251gat;
wire n58gat;
wire n1030gat;
wire n841gat;
wire II4392;
wire n2192gat;
wire n1927gat;
wire n1659gat;
wire n2328gat;
wire n1275gat;
wire II1920;
wire n2698gat;
wire n2138gat;
wire II192;
wire n2839gat;
wire n2256gat;
wire n2927gat;
wire n1991gat;
wire n2978gat;
wire n2569gat;
wire n596gat;
wire II1016;
wire n2039gat;
wire n2977gat;
wire n2209gat;
wire n1784gat;
wire n151gat;
wire n2685gat;
wire n330gat;
wire II1152;
wire II3549;
wire n1380gat;
wire n801gat;
wire n1858gat;
wire II606;
wire n54gat;
wire II3472;
wire n552gat;
wire II2094;
wire n1375gat;
wire n2512gat;
wire n1021gat;
wire n1321gat;
wire n2590gat;
wire II401;
wire n2583gat;
wire n286gat;
wire n2444gat;
wire n2049gat;
wire n2239gat;
wire n387gat;
wire n2906gat;
wire n1582gat;
wire n1230gat;
wire n37gat;
wire II793;
wire II3401;
wire n409gat;
wire II1947;
wire n1469gat;
wire n1180gat;
wire n1146gat;
wire n2181gat;
wire n1702gat;
wire II3163;
wire n2943gat;
wire n381gat;
wire n1649gat;
wire n2462gat;
wire n559gat;
wire n1013gat;
wire n1190gat;
wire n129gat;
wire n1600gat;
wire n2617gat;
wire n358gat;
wire n225gat;
wire n2330gat;
wire II646;
wire II4492;
wire n698gat;
wire n1761gat;
wire n1531gat;
wire n1218gat;
wire n2289gat;
wire n2281gat;
wire II1118;
wire n2624gat;
wire n1204gat;
wire n2790gat;
wire n2437gat;
wire II256;
wire n348gat;
wire n719gat;
wire II2260;
wire n525gat;
wire II1733;
wire n2970gat;
wire II4138;
wire n2550gat;
wire n999gat;
wire n1663gat;
wire n2827gat;
wire n2882gat;
wire n1735gat;
wire n790gat;
wire II468;
wire n133gat;
wire n1262gat;
wire n2108gat;
wire n2854gat;
wire n1452gat;
wire II4236;
wire n1078gat;
wire II913;
wire n1728gat;
wire n15gat;
wire n458gat;
wire II3945;
wire II3457;
wire n1194gat;
wire n242gat;
wire II3999;
wire n1422gat;
wire n2708gat;
wire II3293;
wire n2248gat;
wire n1391gat;
wire n3016gat;
wire n1371gat;
wire n2706gat;
wire II314;
wire II11;
wire n1650gat;
wire n2801gat;
wire n1964gat;
wire II687;
wire n2474gat;
wire n2975gat;
wire n1296gat;
wire II1422;
wire n998gat;
wire n1915gat;
wire n2879gat;
wire n714gat;
wire n288gat;
wire II2148;
wire n967gat;
wire II3483;
wire n1276gat;
wire n2857gat;
wire II4696;
wire n2154gat;
wire n1628gat;
wire n132gat;
wire n1074gat;
wire n2742gat;
wire n3007gat;
wire n2915gat;
wire n1224gat;
wire n1623gat;
wire n2755gat;
wire n2859gat;
wire n2555gat;
wire n2710gat;
wire II3736;
wire n1745gat;
wire n368gat;
wire II963;
wire n1425gat;
wire n21gat;
wire n85gat;
wire n140gat;
wire n2721gat;
wire n2178gat;
wire n901gat;
wire n2628gat;
wire n889gat;
wire n3026gat;
wire n2759gat;
wire n252gat;
wire n1195gat;
wire n93gat;
wire n2995gat;
wire n724gat;
wire II375;
wire n718gat;
wire n339gat;
wire n2806gat;
wire n237gat;
wire n940gat;
wire n1847gat;
wire II3660;
wire n2911gat;
wire n2757gat;
wire n2004gat;
wire n1267gat;
wire n2508gat;
wire II925;
wire n413gat;
wire n254gat;
wire n1743gat;
wire n758gat;
wire n2594gat;
wire n1739gat;
wire n317gat;
wire n483gat;
wire n1698gat;
wire II2414;
wire n504gat;
wire n2461gat;
wire n1360gat;
wire II1371;
wire n595gat;
wire n224gat;
wire n768gat;
wire n1962gat;
wire n2127gat;
wire n836gat;
wire n569gat;
wire n527gat;
wire II4729;
wire n2288gat;
wire n985gat;
wire n2264gat;
wire II2251;
wire n179gat;
wire n784gat;
wire II4601;
wire II2127;
wire n1890gat;
wire n299gat;
wire II47;
wire n2586gat;
wire n2764gat;
wire II1385;
wire n2648gat;
wire n711gat;
wire n832gat;
wire II509;
wire n725gat;
wire n624gat;
wire n2900gat;
wire n1178gat;
wire n2498gat;
wire II217;
wire n1570gat;
wire n2901gat;
wire n1572gat;
wire n2656gat;
wire n1066gat;
wire II4558;
wire n1057gat;
wire n1733gat;
wire n749gat;
wire n2411gat;
wire n3008gat;
wire n2666gat;
wire n243gat;
wire n2051gat;
wire n1716gat;
wire n1256gat;
wire n3021gat;
wire n2647gat;
wire n1297gat;
wire n1971gat;
wire II609;
wire n360gat;
wire n1499gat;
wire n1438gat;
wire II3429;
wire n1472gat;
wire n1440gat;
wire n1756gat;
wire n827gat;
wire n2551gat;
wire n1009gat;
wire n904gat;
wire II18;
wire II1353;
wire II2349;
wire II1450;
wire n2442gat;
wire n697gat;
wire n1916gat;
wire n1079gat;
wire II4587;
wire II210;
wire II4771;
wire II4708;
wire n1797gat;
wire n2800gat;
wire n2398gat;
wire II2926;
wire n1370gat;
wire n45gat;
wire n1209gat;
wire II1752;
wire n1561gat;
wire II658;
wire n859gat;
wire n2415gat;
wire n16gat;
wire n2187gat;
wire n416gat;
wire n1668gat;
wire II2978;
wire n1708gat;
wire II3935;
wire II4741;
wire n1594gat;
wire n2898gat;
wire n2351gat;
wire II692;
wire n1648gat;
wire n2884gat;
wire n2478gat;
wire n1233gat;
wire n174gat;
wire n851gat;
wire n505gat;
wire II4711;
wire n2005gat;
wire n1455gat;
wire n2153gat;
wire n2013gat;
wire n482gat;
wire n1355gat;
wire II1183;
wire n515gat;
wire n2876gat;
wire n1058gat;
wire n1560gat;
wire n1292gat;
wire n2842gat;
wire II2425;
wire n2356gat;
wire n1639gat;
wire n2608gat;
wire n1181gat;
wire n1033gat;
wire II4369;
wire n1453gat;
wire II3016;
wire n401gat;
wire n2700gat;
wire n1552gat;
wire n612gat;
wire II449;
wire n2802gat;
wire II4233;
wire n391gat;
wire II1698;
wire n556gat;
wire n654gat;
wire n873gat;
wire n186gat;
wire II2372;
wire n1300gat;
wire n2333gat;
wire n1261gat;
wire n1213gat;
wire n1626gat;
wire n2346gat;
wire n2636gat;
wire n734gat;
wire n227gat;
wire n2056gat;
wire II354;
wire n1184gat;
wire n575gat;
wire n2081gat;
wire n1229gat;
wire n1667gat;
wire n636gat;
wire n1407gat;
wire n1517gat;
wire n2716gat;
wire n2540gat;
wire II3436;
wire n2940gat;
wire n1098gat;
wire n2123gat;
wire II27;
wire n2914gat;
wire n858gat;
wire n3058gat;
wire n1449gat;
wire n176gat;
wire n1516gat;
wire n2816gat;
wire n869gat;
wire II661;
wire n1478gat;
wire n1413gat;
wire II2439;
wire n1620gat;
wire n531gat;
wire n3046gat;
wire n672gat;
wire n2196gat;
wire II2275;
wire n1106gat;
wire n2745gat;
wire II3587;
wire n261gat;
wire n2831gat;
wire n2999gat;
wire n1329gat;
wire n2856gat;
wire n781gat;
wire n2134gat;
wire n2532gat;
wire n1076gat;
wire n1034gat;
wire n1459gat;
wire n2393gat;
wire n57gat;
wire n2285gat;
wire n644gat;
wire n124gat;
wire n937gat;
wire n579gat;
wire n1796gat;
wire II753;
wire n3041gat;
wire II2420;
wire n1245gat;
wire II1749;
wire n2723gat;
wire n2838gat;
wire n1437gat;
wire n1086gat;
wire n440gat;
wire n1406gat;
wire II3287;
wire II3817;
wire n1396gat;
wire n3048gat;
wire n411gat;
wire II334;
wire n730gat;
wire n2561gat;
wire n378gat;
wire II3558;
wire n207gat;
wire n2619gat;
wire II2228;
wire n1470gat;
wire n1071gat;
wire n1691gat;
wire II2736;
wire n412gat;
wire n557gat;
wire n1481gat;
wire II2889;
wire n1575gat;
wire n2784gat;
wire n1238gat;
wire n2920gat;
wire n2568gat;
wire n1397gat;
wire II1703;
wire n2524gat;
wire n2566gat;
wire II3610;
wire n450gat;
wire n2533gat;
wire n2542gat;
wire n163gat;
wire n2015gat;
wire II2684;
wire n833gat;
wire n2559gat;
wire II1127;
wire n390gat;
wire II1915;
wire n763gat;
wire II1766;
wire n914gat;
wire n2567gat;
wire II3876;
wire II2235;
wire n641gat;
wire II4157;
wire n2864gat;
wire n442gat;
wire n872gat;
wire n1661gat;
wire n2258gat;
wire II384;
wire II4738;
wire n717gat;
wire n171gat;
wire n895gat;
wire n942gat;
wire n2825gat;
wire n706gat;
wire n497gat;
wire n1092gat;
wire n296gat;
wire II1617;
wire II885;
wire n2711gat;
wire II2248;
wire II1103;
wire n797gat;
wire n564gat;
wire n1206gat;
wire n60gat;
wire n1349gat;
wire n2817gat;
wire n1327gat;
wire n2979gat;
wire II1800;
wire n1730gat;
wire n1384gat;
wire n383gat;
wire n1383gat;
wire n787gat;
wire n2364gat;
wire n1665gat;
wire n155gat;
wire II4608;
wire n2994gat;
wire n2761gat;
wire n1022gat;
wire n1621gat;
wire II1088;
wire n1005gat;
wire II4185;
wire n845gat;
wire II1178;
wire n844gat;
wire n2306gat;
wire n567gat;
wire n2611gat;
wire n995gat;
wire n1003gat;
wire n2958gat;
wire II4693;
wire II3914;
wire n2690gat;
wire II3318;
wire n2963gat;
wire n250gat;
wire n2973gat;
wire n1515gat;
wire n973gat;
wire n1633gat;
wire n1731gat;
wire n1255gat;
wire n1176gat;
wire n650gat;
wire II2354;
wire n500gat;
wire n1237gat;
wire n495gat;
wire n1640gat;
wire n2929gat;
wire II955;
wire n349gat;
wire n1692gat;
wire II1550;
wire n1711gat;
wire n2928gat;
wire n2961gat;
wire II3962;
wire II709;
wire II4615;
wire n2290gat;
wire n2638gat;
wire n1088gat;
wire n2001gat;
wire n2000gat;
wire II818;
wire n2954gat;
wire n657gat;
wire n1347gat;
wire II270;
wire n1171gat;
wire n2614gat;
wire n77gat;
wire n1544gat;
wire n1793gat;
wire n1510gat;
wire n2307gat;
wire II1734;
wire n1622gat;
wire II214;
wire II2162;
wire n359gat;
wire n2581gat;
wire n2968gat;
wire n3031gat;
wire n478gat;
wire II2056;
wire n87gat;
wire n2396gat;
wire n1272gat;
wire n462gat;
wire n936gat;
wire n2701gat;
wire n2912gat;
wire n320gat;
wire n796gat;
wire n2851gat;
wire n1156gat;
wire n3033gat;
wire n854gat;
wire n2412gat;
wire n837gat;
wire II3646;
wire II3390;
wire II297;
wire n2341gat;
wire n335gat;
wire n1569gat;
wire n2250gat;
wire n3051gat;
wire n1044gat;
wire II1981;
wire n1504gat;
wire n2047gat;
wire n88gat;
wire n371gat;
wire n882gat;
wire II2925;
wire n3038gat;
wire II3491;
wire n2971gat;
wire n908gat;
wire n1652gat;
wire n1747gat;
wire n1258gat;
wire n2245gat;
wire n1959gat;
wire n3022gat;
wire n316gat;
wire n55gat;
wire n2152gat;
wire n902gat;
wire n1196gat;
wire n2837gat;
wire n1657gat;
wire n3061gat;
wire n1284gat;
wire n994gat;
wire II1011;
wire II4482;
wire II1903;
wire n2669gat;
wire n528gat;
wire n1896gat;
wire II223;
wire n489gat;
wire II2376;
wire n566gat;
wire n1056gat;
wire n560gat;
wire n2902gat;
wire n1286gat;
wire II4312;
wire n1503gat;
wire n41gat;
wire n2260gat;
wire n2090gat;
wire II2843;
wire II623;
wire n126gat;
wire n870gat;
wire n1645gat;
wire n1758gat;
wire II4542;
wire II4675;
wire n3024gat;
wire II4055;
wire II275;
wire n823gat;
wire II1277;
wire II1302;
wire n2549gat;
wire n1339gat;
wire n1828gat;
wire n2680gat;
wire n1616gat;
wire n511gat;
wire n592gat;
wire n265gat;
wire II2935;
wire n350gat;
wire n529gat;
wire II4780;
wire n2782gat;
wire n3005gat;
wire n1832gat;
wire II1655;
wire n780gat;
wire n1427gat;
wire n639gat;
wire II2319;
wire II4014;
wire II461;
wire n374gat;
wire n1133gat;
wire n1926gat;
wire n326gat;
wire n1093gat;
wire n66gat;
wire n110gat;
wire n1188gat;
wire II2088;
wire n1644gat;
wire n695gat;
wire n2438gat;
wire n2188gat;
wire n972gat;
wire II3309;
wire II4566;
wire n1177gat;
wire II916;
wire n480gat;
wire n1601gat;
wire n1304gat;
wire n2643gat;
wire II4795;
wire n1307gat;
wire n2799gat;
wire n894gat;
wire n1862gat;
wire n475gat;
wire n663gat;
wire II2169;
wire n2807gat;
wire n900gat;
wire n1319gat;
wire II3168;
wire n822gat;
wire n971gat;
wire n238gat;
wire n1240gat;
wire II3000;
wire n693gat;
wire n621gat;
wire II2785;
wire n245gat;
wire n417gat;
wire II1305;
wire n248gat;
wire n613gat;
wire n1658gat;
wire II718;
wire n2031gat;
wire n682gat;
wire n2980gat;
wire n2715gat;
wire II14;
wire n2796gat;
wire n918gat;
wire n1654gat;
wire n2813gat;
wire n628gat;
wire n1273gat;
wire n912gat;
wire n2888gat;
wire II1141;
wire n1243gat;
wire n2331gat;
wire n2466gat;
wire n2012gat;
wire II3777;
wire n14gat;
wire n1518gat;
wire II1500;
wire n1895gat;
wire n268gat;
wire II2281;
wire n642gat;
wire n1817gat;
wire II2771;
wire n977gat;
wire n665gat;
wire n1085gat;
wire II4762;
wire n1631gat;
wire n61gat;
wire n671gat;
wire n2058gat;
wire II196;
wire n1443gat;
wire n518gat;
wire n1454gat;
wire n1020gat;
wire n404gat;
wire n2989gat;
wire n1265gat;
wire n720gat;
wire n2889gat;
wire n570gat;
wire n123gat;
wire II2157;
wire n137gat;
wire n1712gat;
wire n281gat;
wire n1401gat;
wire n2754gat;
wire n713gat;
wire n652gat;
wire n3029gat;
wire n1627gat;
wire II2268;
wire n772gat;
wire n1084gat;
wire n2268gat;
wire n1683gat;
wire n2019gat;
wire n2678gat;
wire II4750;
wire II4759;
wire n456gat;
wire n340gat;
wire II2271;
wire II1190;
wire II1843;
wire n953gat;
wire n1118gat;
wire n1892gat;
wire n258gat;
wire n2142gat;
wire n2824gat;
wire II594;
wire n1187gat;
wire n2448gat;
wire n1604gat;
wire II3530;
wire n352gat;
wire II1169;
wire n2703gat;
wire n2489gat;
wire n1217gat;
wire n2552gat;
wire n670gat;
wire n1695gat;
wire n2803gat;
wire n1755gat;
wire n661gat;
wire n2756gat;
wire n70gat;
wire n1032gat;
wire n2265gat;
wire n2585gat;
wire n2546gat;
wire n558gat;
wire n1956gat;
wire II1388;
wire n1426gat;
wire n1801gat;
wire II3841;
wire n950gat;
wire n2887gat;
wire n1293gat;
wire II453;
wire n1191gat;
wire n2875gat;
wire n1990gat;
wire n154gat;
wire n2017gat;
wire n616gat;
wire n761gat;
wire II4633;
wire n868gat;
wire II1606;
wire n2198gat;
wire n1192gat;
wire n251gat;
wire n2765gat;
wire n802gat;
wire n233gat;
wire n1119gat;
wire n1870gat;
wire n1325gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n673gat <= 1;
  else
    n673gat <= n2897gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n398gat <= 1;
  else
    n398gat <= n2782gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n402gat <= 1;
  else
    n402gat <= n2790gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n919gat <= 1;
  else
    n919gat <= n2670gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n846gat <= 1;
  else
    n846gat <= n2793gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2510gat <= 1;
  else
    n2510gat <= n748gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n271gat <= 1;
  else
    n271gat <= n2732gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n160gat <= 1;
  else
    n160gat <= n2776gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n337gat <= 1;
  else
    n337gat <= n2735gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n842gat <= 1;
  else
    n842gat <= n2673gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n341gat <= 1;
  else
    n341gat <= n2779gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2522gat <= 1;
  else
    n2522gat <= n43gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2472gat <= 1;
  else
    n2472gat <= n1620gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2319gat <= 1;
  else
    n2319gat <= n2470gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1821gat <= 1;
  else
    n1821gat <= n1827gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2029gat <= 1;
  else
    n2029gat <= n1816gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1829gat <= 1;
  else
    n1829gat <= n2027gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2476gat <= 1;
  else
    n2476gat <= n55gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1068gat <= 1;
  else
    n1068gat <= n2914gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n957gat <= 1;
  else
    n957gat <= n2928gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n861gat <= 1;
  else
    n861gat <= n2927gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1294gat <= 1;
  else
    n1294gat <= n2896gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1241gat <= 1;
  else
    n1241gat <= n2922gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n865gat <= 1;
  else
    n865gat <= n2894gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1080gat <= 1;
  else
    n1080gat <= n2921gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1148gat <= 1;
  else
    n1148gat <= n2895gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2468gat <= 1;
  else
    n2468gat <= n933gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n834gat <= 1;
  else
    n834gat <= n3064gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n707gat <= 1;
  else
    n707gat <= n3055gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n838gat <= 1;
  else
    n838gat <= n3063gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n830gat <= 1;
  else
    n830gat <= n3062gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n614gat <= 1;
  else
    n614gat <= n3056gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2526gat <= 1;
  else
    n2526gat <= n504gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n680gat <= 1;
  else
    n680gat <= n2913gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n816gat <= 1;
  else
    n816gat <= n2920gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n580gat <= 1;
  else
    n580gat <= n2905gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n824gat <= 1;
  else
    n824gat <= n3057gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n820gat <= 1;
  else
    n820gat <= n3059gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n883gat <= 1;
  else
    n883gat <= n3058gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n584gat <= 1;
  else
    n584gat <= n2898gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n684gat <= 1;
  else
    n684gat <= n3060gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n699gat <= 1;
  else
    n699gat <= n3061gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2464gat <= 1;
  else
    n2464gat <= n567gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2399gat <= 1;
  else
    n2399gat <= n3048gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2343gat <= 1;
  else
    n2343gat <= n3049gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2203gat <= 1;
  else
    n2203gat <= n3051gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2562gat <= 1;
  else
    n2562gat <= n3047gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2207gat <= 1;
  else
    n2207gat <= n3050gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2626gat <= 1;
  else
    n2626gat <= n3040gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2490gat <= 1;
  else
    n2490gat <= n3044gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2622gat <= 1;
  else
    n2622gat <= n3042gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2630gat <= 1;
  else
    n2630gat <= n3037gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2543gat <= 1;
  else
    n2543gat <= n3041gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2102gat <= 1;
  else
    n2102gat <= n1606gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1880gat <= 1;
  else
    n1880gat <= n3052gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1763gat <= 1;
  else
    n1763gat <= n1610gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2155gat <= 1;
  else
    n2155gat <= n1858gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1035gat <= 1;
  else
    n1035gat <= n2918gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1121gat <= 1;
  else
    n1121gat <= n2952gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1072gat <= 1;
  else
    n1072gat <= n2919gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1282gat <= 1;
  else
    n1282gat <= n2910gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1226gat <= 1;
  else
    n1226gat <= n2907gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n931gat <= 1;
  else
    n931gat <= n2911gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1135gat <= 1;
  else
    n1135gat <= n2912gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1045gat <= 1;
  else
    n1045gat <= n2909gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1197gat <= 1;
  else
    n1197gat <= n2908gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2518gat <= 1;
  else
    n2518gat <= n2971gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n667gat <= 1;
  else
    n667gat <= n2904gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n659gat <= 1;
  else
    n659gat <= n2891gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n553gat <= 1;
  else
    n553gat <= n2903gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n777gat <= 1;
  else
    n777gat <= n2915gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n561gat <= 1;
  else
    n561gat <= n2901gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n366gat <= 1;
  else
    n366gat <= n2890gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n322gat <= 1;
  else
    n322gat <= n2888gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n318gat <= 1;
  else
    n318gat <= n2887gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n314gat <= 1;
  else
    n314gat <= n2886gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2599gat <= 1;
  else
    n2599gat <= n3010gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2588gat <= 1;
  else
    n2588gat <= n3016gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2640gat <= 1;
  else
    n2640gat <= n3054gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2658gat <= 1;
  else
    n2658gat <= n2579gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2495gat <= 1;
  else
    n2495gat <= n3036gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2390gat <= 1;
  else
    n2390gat <= n3034gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2270gat <= 1;
  else
    n2270gat <= n3031gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2339gat <= 1;
  else
    n2339gat <= n3035gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2502gat <= 1;
  else
    n2502gat <= n2646gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2634gat <= 1;
  else
    n2634gat <= n3053gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2506gat <= 1;
  else
    n2506gat <= n2613gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1834gat <= 1;
  else
    n1834gat <= n1625gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1767gat <= 1;
  else
    n1767gat <= n1626gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2084gat <= 1;
  else
    n2084gat <= n1603gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2143gat <= 1;
  else
    n2143gat <= n2541gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2061gat <= 1;
  else
    n2061gat <= n2557gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2139gat <= 1;
  else
    n2139gat <= n2487gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1899gat <= 1;
  else
    n1899gat <= n2532gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1850gat <= 1;
  else
    n1850gat <= n2628gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2403gat <= 1;
  else
    n2403gat <= n2397gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2394gat <= 1;
  else
    n2394gat <= n2341gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2440gat <= 1;
  else
    n2440gat <= n2560gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2407gat <= 1;
  else
    n2407gat <= n2205gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2347gat <= 1;
  else
    n2347gat <= n2201gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1389gat <= 1;
  else
    n1389gat <= n1793gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2021gat <= 1;
  else
    n2021gat <= n1781gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1394gat <= 1;
  else
    n1394gat <= n1516gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1496gat <= 1;
  else
    n1496gat <= n1392gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2091gat <= 1;
  else
    n2091gat <= n1685gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1332gat <= 1;
  else
    n1332gat <= n1565gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1740gat <= 1;
  else
    n1740gat <= n1330gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2179gat <= 1;
  else
    n2179gat <= n1945gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2190gat <= 1;
  else
    n2190gat <= n2268gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2135gat <= 1;
  else
    n2135gat <= n2337gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2262gat <= 1;
  else
    n2262gat <= n2388gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2182gat <= 1;
  else
    n2182gat <= n1836gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1433gat <= 1;
  else
    n1433gat <= n2983gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1316gat <= 1;
  else
    n1316gat <= n1431gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1363gat <= 1;
  else
    n1363gat <= n1314gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1312gat <= 1;
  else
    n1312gat <= n1361gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1775gat <= 1;
  else
    n1775gat <= n1696gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1871gat <= 1;
  else
    n1871gat <= n2009gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2592gat <= 1;
  else
    n2592gat <= n1773gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1508gat <= 1;
  else
    n1508gat <= n1636gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1678gat <= 1;
  else
    n1678gat <= n1712gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2309gat <= 1;
  else
    n2309gat <= n3000gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2450gat <= 1;
  else
    n2450gat <= n2307gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2446gat <= 1;
  else
    n2446gat <= n2661gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2095gat <= 1;
  else
    n2095gat <= n827gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2176gat <= 1;
  else
    n2176gat <= n2093gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2169gat <= 1;
  else
    n2169gat <= n2174gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2454gat <= 1;
  else
    n2454gat <= n2163gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2040gat <= 1;
  else
    n2040gat <= n1777gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2044gat <= 1;
  else
    n2044gat <= n2015gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2037gat <= 1;
  else
    n2037gat <= n2042gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2025gat <= 1;
  else
    n2025gat <= n2017gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2099gat <= 1;
  else
    n2099gat <= n2023gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2266gat <= 1;
  else
    n2266gat <= n2493gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2033gat <= 1;
  else
    n2033gat <= n2035gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2110gat <= 1;
  else
    n2110gat <= n2031gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2125gat <= 1;
  else
    n2125gat <= n2108gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2121gat <= 1;
  else
    n2121gat <= n2123gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2117gat <= 1;
  else
    n2117gat <= n2119gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1975gat <= 1;
  else
    n1975gat <= n2632gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2644gat <= 1;
  else
    n2644gat <= n2638gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n156gat <= 1;
  else
    n156gat <= n612gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n152gat <= 1;
  else
    n152gat <= n705gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n331gat <= 1;
  else
    n331gat <= n822gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n388gat <= 1;
  else
    n388gat <= n881gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n463gat <= 1;
  else
    n463gat <= n818gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n327gat <= 1;
  else
    n327gat <= n682gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n384gat <= 1;
  else
    n384gat <= n697gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n256gat <= 1;
  else
    n256gat <= n836gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n470gat <= 1;
  else
    n470gat <= n828gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n148gat <= 1;
  else
    n148gat <= n832gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2458gat <= 1;
  else
    n2458gat <= n2590gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n2514gat <= 1;
  else
    n2514gat <= n2456gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1771gat <= 1;
  else
    n1771gat <= n1613gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1336gat <= 1;
  else
    n1336gat <= n1391gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1748gat <= 1;
  else
    n1748gat <= n1927gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1675gat <= 1;
  else
    n1675gat <= n1713gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1807gat <= 1;
  else
    n1807gat <= n1717gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1340gat <= 1;
  else
    n1340gat <= n1567gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1456gat <= 1;
  else
    n1456gat <= n1564gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1525gat <= 1;
  else
    n1525gat <= n1632gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1462gat <= 1;
  else
    n1462gat <= n1915gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1596gat <= 1;
  else
    n1596gat <= n1800gat;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    n1588gat <= 1;
  else
    n1588gat <= n1593gat;
assign n43gat = (n44gat)|(n45gat)|(n46gat)|(n47gat);
assign n1967gat = ((~n1893gat)&(~n1968gat));
assign II1344 = ((~n814gat));
assign n911gat = ((~II661));
assign n2167gat = ((~n2169gat));
assign n2612gat = ((~n2620gat));
assign n1706gat = ((~n1622gat));
assign n419gat = ((~n409gat)&(~n291gat));
assign n1724gat = ((~n1732gat));
assign II4690 = ((~n2685gat));
assign n3144gat = ((~II4774));
assign II476 = ((~n475gat));
assign II4518 = ((~n2761gat));
assign II880 = ((~n1293gat));
assign n3044gat = ((~II3504));
assign n2791gat = ((~II62));
assign n221gat = (n222gat)|(n223gat)|(n224gat)|(n225gat);
assign n1202gat = ((~n1206gat)&(~n1207gat)&(~n1208gat));
assign II2915 = ((~n1740gat));
assign II1416 = ((~n822gat));
assign n588gat = ((~n591gat)&(~n594gat)&(~n595gat));
assign II2232 = ((~n2640gat));
assign n1358gat = ((~n1425gat)&(~n1105gat));
assign n974gat = ((~n2844gat)&(~n111gat));
assign n194gat = ((~n187gat));
assign n702gat = ((~II149));
assign n696gat = ((~II1481));
assign n1719gat = ((~n1548gat));
assign n443gat = ((~n2778gat)&(~n373gat));
assign n952gat = ((~II842));
assign II4783 = ((~n2827gat));
assign n2577gat = ((~II2238));
assign n499gat = ((~II1085));
assign n1175gat = ((~n621gat)&(~n1006gat));
assign n2023gat = ((~n2025gat));
assign II4212 = ((~n1588gat));
assign n1790gat = ((~n1726gat));
assign n1656gat = ((~n1655gat));
assign II2394 = ((~n2557gat));
assign n2845gat = ((~II23));
assign n1225gat = ((~II1833));
assign II2344 = ((~n2339gat));
assign n1172gat = ((~n2961gat)&(~n1200gat));
assign n63gat = ((~II746));
assign n878gat = ((~n2879gat));
assign n2050gat = ((~n2146gat));
assign n17gat = ((~n564gat));
assign n2683gat = ((~II3951));
assign n2746gat = ((~II4536));
assign n782gat = ((~n789gat)&(~n785gat)&(~n788gat));
assign II2263 = ((~n2202gat));
assign n2655gat = ((~n2508gat)&(~n2656gat)&(~n2500gat)&(~n2504gat));
assign n2661gat = ((~n2662gat));
assign n757gat = ((~II278));
assign n1303gat = ((~n1247gat)&(~n1355gat));
assign n2652gat = ((~II2354));
assign n1002gat = ((~n2946gat));
assign n2850gat = ((~II579));
assign n1291gat = ((~n1603gat)&(~n579gat));
assign n2607gat = ((~II2376));
assign n721gat = ((~II178));
assign n2418gat = ((~II2271));
assign n2621gat = ((~II1617));
assign n1219gat = ((~II203));
assign n2433gat = ((~n2432gat)&(~n2154gat));
assign n786gat = ((~II2035));
assign n1050gat = (n1051gat)|(n1052gat)|(n1053gat)|(n1054gat);
assign II2934 = (n1784gat)|(n1839gat)|(n1788gat);
assign n3001gat = (n2132gat)|(n2130gat);
assign II985 = ((~n3078gat));
assign II437 = ((~n341gat));
assign II227 = ((~n2856gat));
assign n1008gat = ((~n2942gat)&(~n1254gat));
assign II4699 = ((~n2745gat));
assign n1584gat = ((~n2989gat));
assign II1007 = ((~n1078gat));
assign II4777 = ((~n2699gat));
assign II846 = ((~n859gat));
assign n813gat = ((~II1353));
assign n632gat = ((~n414gat)&(~n523gat)&(~n633gat));
assign n2832gat = ((~II768));
assign II726 = ((~n400gat));
assign n2046gat = ((~n2269gat));
assign n1215gat = ((~n1218gat)&(~n1221gat)&(~n1222gat));
assign n1423gat = ((~n2162gat)&(~n1530gat));
assign n1361gat = ((~n1363gat));
assign n2488gat = ((~n2490gat));
assign n508gat = ((~n514gat)&(~n512gat)&(~n511gat));
assign II1708 = ((~n2543gat));
assign n2942gat = (n904gat)|(n903gat);
assign n2355gat = ((~n2341gat));
assign n1212gat = ((~n1123gat)&(~n1034gat));
assign II4642 = ((~n2812gat));
assign II3509 = ((~n2438gat));
assign n1161gat = ((~n583gat)&(~n1603gat));
assign n2223gat = ((~n2354gat)&(~n2217gat));
assign n410gat = ((~n417gat)&(~n413gat)&(~n412gat)&(~n406gat));
assign II2847 = ((~n2394gat));
assign n746gat = ((~n2716gat)&(~n2723gat));
assign n766gat = ((~n93gat)&(~n2734gat));
assign II2385 = ((~n2536gat));
assign II2324 = ((~n3014gat));
assign n1701gat = ((~n1617gat));
assign n960gat = ((~n2734gat)&(~n852gat));
assign n2741gat = (n1182gat)|(n2385gat);
assign n1221gat = ((~II217));
assign n2913gat = (n767gat)|(n653gat);
assign n2452gat = ((~n2454gat));
assign n386gat = ((~n388gat));
assign II3342 = ((~n1316gat));
assign n2186gat = ((~n2613gat));
assign n351gat = ((~II726));
assign n2237gat = ((~n2646gat));
assign n1606gat = ((~n3020gat)&(~n270gat));
assign n2243gat = ((~n55gat));
assign n1444gat = ((~n1442gat));
assign n212gat = ((~n182gat)&(~n78gat));
assign n955gat = ((~n957gat));
assign n136gat = ((~n253gat)&(~n154gat));
assign n1480gat = ((~n2292gat));
assign n2944gat = (n977gat)|(n976gat);
assign n2694gat = (n1381gat)|(n1384gat);
assign n1670gat = ((~n1667gat));
assign n1694gat = ((~II2813));
assign n2151gat = ((~n2193gat));
assign n3019gat = ((~II3235));
assign n1163gat = ((~n882gat)&(~n1603gat));
assign II3954 = ((~n2683gat));
assign II1067 = ((~n616gat));
assign II311 = ((~n271gat));
assign II2885 = ((~n2091gat));
assign n2149gat = ((~n2193gat)&(~n2346gat));
assign n2733gat = ((~II297));
assign n855gat = ((~n2148gat));
assign n1174gat = ((~n845gat)&(~n1007gat));
assign n1164gat = ((~n2953gat));
assign II4657 = ((~n2809gat));
assign n2486gat = ((~n2629gat));
assign n688gat = ((~n691gat)&(~n694gat)&(~n695gat));
assign n910gat = ((~n916gat)&(~n914gat)&(~n913gat));
assign n1838gat = ((~n1898gat));
assign n2749gat = (n1010gat)|(n2246gat);
assign n2860gat = ((~II214));
assign n490gat = ((~II1088));
assign n1792gat = ((~n1794gat)&(~n1796gat));
assign n2421gat = ((~n1601gat)&(~n1704gat));
assign n127gat = ((~II2169));
assign II1360 = ((~n677gat));
assign n2852gat = ((~n2853gat));
assign n1263gat = ((~n1212gat)&(~n2968gat));
assign n959gat = ((~n373gat)&(~n2734gat));
assign n1729gat = ((~n1658gat)&(~n1797gat)&(~n1568gat));
assign n2702gat = (n925gat)|(n1452gat);
assign II359 = ((~n158gat));
assign n1448gat = ((~n1376gat));
assign n2863gat = ((~II220));
assign II3923 = ((~n2710gat));
assign II512 = ((~n2730gat));
assign n2500gat = ((~n2502gat));
assign n1555gat = ((~n1616gat)&(~n1559gat)&(~n1499gat));
assign n646gat = ((~n93gat)&(~n2669gat));
assign n692gat = ((~II1453));
assign n2325gat = ((~n3010gat));
assign n1532gat = ((~n1677gat)&(~n1458gat));
assign n2148gat = ((~II1734));
assign n1502gat = ((~n1607gat)&(~n1449gat));
assign n1014gat = ((~n1018gat)&(~n1019gat)&(~n1020gat));
assign n453gat = ((~n372gat)&(~n452gat));
assign II4429 = ((~n2936gat));
assign n925gat = ((~n927gat));
assign II2153 = ((~n316gat));
assign II4135 = ((~n3098gat));
assign n2910gat = (n645gat)|(n644gat);
assign II149 = ((~n402gat));
assign n1104gat = ((~n1079gat)&(~n1590gat));
assign n2672gat = ((~n2674gat));
assign n1859gat = ((~n1717gat));
assign II2084 = ((~n366gat));
assign n1945gat = ((~n1690gat));
assign n1619gat = ((~n1447gat)&(~n1446gat));
assign n2660gat = ((~n2655gat));
assign n2689gat = ((~II4573));
assign n1548gat = ((~II2721));
assign II3235 = ((~n2238gat));
assign n996gat = ((~n1603gat)&(~n823gat));
assign n2795gat = ((~II4615));
assign n1989gat = ((~n2401gat));
assign n3121gat = ((~II4705));
assign n923gat = ((~n1043gat));
assign II2242 = ((~n2341gat));
assign n1193gat = ((~II1795));
assign n947gat = ((~n954gat)&(~n950gat)&(~n953gat));
assign n2693gat = (n1451gat)|(n1453gat);
assign II4217 = (n1392gat)|(n2989gat)|(II4216);
assign n857gat = ((~n944gat));
assign n2986gat = (n1650gat)|(n1649gat)|(n1563gat);
assign II2831 = (n1839gat)|(n1786gat)|(n1788gat);
assign n1879gat = ((~II1667));
assign n40gat = ((~n325gat)&(~n383gat));
assign n3140gat = ((~II4762));
assign II111 = ((~n846gat));
assign n2238gat = ((~n2448gat)&(~n2444gat));
assign n779gat = (n780gat)|(n781gat)|(n782gat)|(n783gat);
assign n756gat = ((~II275));
assign n1878gat = ((~n1880gat));
assign n1550gat = ((~II2890));
assign n2449gat = ((~II3957));
assign n219gat = ((~n78gat));
assign n1067gat = ((~II790));
assign n1173gat = ((~n1007gat)&(~n1025gat));
assign II4792 = ((~n2680gat));
assign n1925gat = ((~n1920gat));
assign n1223gat = ((~II230));
assign n277gat = ((~n337gat));
assign II902 = ((~n1240gat));
assign n1330gat = ((~n1332gat));
assign n2534gat = ((~n2624gat)&(~n2489gat)&(~n2621gat));
assign n415gat = ((~n2723gat)&(~n740gat));
assign n907gat = ((~n911gat)&(~n912gat)&(~n913gat));
assign n3009gat = (n2350gat)|(n2282gat);
assign n3142gat = ((~II4768));
assign n370gat = ((~n1725gat));
assign n683gat = ((~II1450));
assign n513gat = ((~II1251));
assign n874gat = ((~n559gat)&(~n365gat));
assign n2814gat = ((~II4309));
assign n178gat = ((~n343gat));
assign n2052gat = ((~n2393gat));
assign n2709gat = (n739gat)|(n1841gat);
assign n2133gat = ((~n2135gat));
assign II4475 = ((~n2951gat));
assign n2213gat = ((~n2402gat)&(~n2151gat)&(~n2345gat));
assign n2955gat = (n1177gat)|(n1115gat);
assign n22gat = ((~n92gat)&(~n21gat));
assign n807gat = ((~n813gat)&(~n811gat)&(~n810gat));
assign II62 = ((~n3070gat));
assign n990gat = ((~n841gat)&(~n741gat));
assign n2018gat = ((~n2016gat)&(~n2097gat));
assign n1309gat = ((~n2959gat));
assign II583 = ((~n2786gat));
assign n653gat = ((~n2718gat)&(~n111gat));
assign II2174 = ((~n133gat));
assign n875gat = ((~n559gat));
assign n733gat = ((~II1121));
assign n523gat = ((~n522gat)&(~n356gat));
assign n2932gat = (n1098gat)|(n1090gat)|(n986gat)|(n885gat);
assign n53gat = ((~II480));
assign n1524gat = ((~II4157));
assign n1485gat = ((~n1482gat)&(~n2162gat));
assign n3036gat = ((~II3436));
assign n1324gat = ((~n164gat)&(~n1007gat));
assign n1887gat = ((~n2138gat));
assign n247gat = ((~n334gat)&(~n387gat)&(~n330gat));
assign II3691 = ((~n152gat));
assign II1082 = ((~n402gat));
assign n1099gat = ((~n1111gat)&(~n1293gat));
assign n1123gat = ((~n632gat));
assign n172gat = ((~II609));
assign n1270gat = ((~n1274gat)&(~n1275gat)&(~n1276gat));
assign II4687 = ((~n2690gat));
assign n1690gat = ((~n1700gat)&(~n1702gat));
assign n2939gat = (n1091gat)|(n1088gat)|(n992gat)|(n987gat);
assign n916gat = ((~II692));
assign II637 = ((~n278gat));
assign II3143 = ((~n2592gat));
assign n1610gat = ((~n1698gat)&(~n1543gat));
assign n3045gat = ((~II3509));
assign n1636gat = ((~n1584gat)&(~n1718gat));
assign n1436gat = ((~n1435gat));
assign n2128gat = ((~n2129gat));
assign n1214gat = ((~n1218gat)&(~n1219gat)&(~n1220gat));
assign n2697gat = ((~II4587));
assign n1495gat = ((~II2873));
assign n880gat = ((~n926gat)&(~n566gat));
assign II97 = ((~n3071gat));
assign n2553gat = ((~II2425));
assign II65 = ((~n2791gat));
assign n649gat = ((~n2778gat)&(~n852gat));
assign n992gat = ((~n815gat)&(~n1112gat));
assign n1095gat = ((~n1240gat)&(~n1111gat));
assign n1115gat = ((~n1263gat)&(~n419gat));
assign n1917gat = ((~n1921gat));
assign n573gat = ((~II1422));
assign n2350gat = ((~n2405gat)&(~n2349gat));
assign n1551gat = ((~n1549gat));
assign n1015gat = ((~n1018gat)&(~n1021gat)&(~n1022gat));
assign II320 = ((~n2777gat));
assign n2035gat = ((~n2037gat));
assign n2456gat = ((~n2458gat));
assign II842 = ((~n955gat));
assign II721 = ((~n397gat));
assign n1613gat = ((~n1544gat)&(~n1698gat));
assign n1158gat = ((~n983gat)&(~n1157gat));
assign II4660 = ((~n2801gat));
assign n899gat = ((~n419gat)&(~n1172gat));
assign II395 = ((~n842gat));
assign n2753gat = ((~II4530));
assign II1724 = (n2355gat)|(n2443gat)|(II1723);
assign n2775gat = ((~n2777gat));
assign II4489 = ((~n2046gat));
assign II220 = ((~n2864gat));
assign n2962gat = (n1176gat)|(n1173gat);
assign n1788gat = ((~n2142gat));
assign n71gat = ((~n180gat));
assign n270gat = ((~II311));
assign n748gat = (n749gat)|(n750gat)|(n751gat)|(n752gat);
assign n3120gat = ((~II4702));
assign n1271gat = ((~n1274gat)&(~n1277gat)&(~n1278gat));
assign II4309 = ((~n2941gat));
assign n1441gat = ((~n1437gat)&(~n1378gat));
assign II3867 = ((~n470gat));
assign n1420gat = ((~n1410gat)&(~n2162gat));
assign n1479gat = ((~n2291gat));
assign n1483gat = ((~n2081gat)&(~n1482gat));
assign n520gat = ((~n374gat)&(~n2862gat));
assign n267gat = ((~II363));
assign n1685gat = ((~n1604gat));
assign n2269gat = ((~II2349));
assign II2044 = ((~n775gat));
assign II2035 = ((~n776gat));
assign II4499 = ((~n2688gat));
assign n507gat = ((~n514gat)&(~n510gat)&(~n513gat));
assign n1662gat = ((~n1663gat));
assign II4630 = ((~n1086gat));
assign n2777gat = ((~II317));
assign n1605gat = ((~n1614gat)&(~n1616gat)&(~n1499gat)&(~n396gat));
assign II4020 = ((~n2800gat));
assign n775gat = ((~n777gat));
assign n2981gat = (n1413gat)|(n1408gat)|(n1407gat);
assign n809gat = ((~II1322));
assign n769gat = ((~n93gat)&(~n2731gat));
assign n930gat = ((~II1857));
assign n635gat = ((~n639gat)&(~n634gat)&(~n414gat));
assign II3394 = ((~n2260gat));
assign n1096gat = ((~n819gat)&(~n1112gat));
assign n2948gat = (n1097gat)|(n1089gat)|(n1087gat)|(n991gat);
assign II340 = ((~n2736gat));
assign n571gat = ((~n577gat)&(~n575gat)&(~n574gat));
assign n2115gat = ((~n2117gat));
assign n1382gat = ((~n1280gat));
assign n3047gat = ((~II3520));
assign n864gat = ((~II955));
assign n2591gat = ((~II3143));
assign n926gat = ((~n632gat));
assign n897gat = ((~n2939gat));
assign n293gat = ((~n361gat));
assign n2907gat = (n646gat)|(n641gat);
assign n344gat = ((~n348gat)&(~n349gat)&(~n350gat));
assign II4389 = ((~n2956gat));
assign II678 = ((~n918gat));
assign n986gat = ((~n985gat)&(~n926gat));
assign n1326gat = ((~n1007gat)&(~n282gat));
assign n170gat = ((~n177gat)&(~n173gat)&(~n176gat));
assign n1955gat = ((~n1956gat));
assign II4723 = ((~n2677gat));
assign II378 = ((~n725gat));
assign n253gat = ((~n1702gat));
assign n2539gat = ((~n2048gat)&(~n2437gat));
assign II3387 = ((~n2194gat));
assign n783gat = ((~n789gat)&(~n787gat)&(~n786gat));
assign n1934gat = ((~n2470gat)&(~n1935gat)&(~n2239gat));
assign n175gat = ((~II642));
assign n1960gat = ((~n3043gat));
assign II1723 = (n2354gat)|(n2353gat)|(n2214gat);
assign n694gat = ((~II1472));
assign n983gat = ((~n320gat));
assign II253 = ((~n2906gat));
assign n1023gat = ((~II414));
assign n1393gat = ((~II3168));
assign n144gat = ((~n247gat));
assign n2637gat = ((~n3015gat)&(~n2199gat));
assign n2359gat = ((~n2358gat));
assign n3017gat = ((~II1961));
assign n771gat = ((~n2838gat)&(~n111gat));
assign n2908gat = (n763gat)|(n642gat);
assign n1920gat = ((~n1864gat)&(~n1921gat)&(~n1798gat));
assign n2216gat = ((~n2406gat));
assign n582gat = ((~n584gat));
assign n56gat = ((~n60gat)&(~n61gat)&(~n62gat));
assign n2789gat = ((~n2791gat));
assign n679gat = ((~II1302));
assign II456 = ((~n392gat));
assign n204gat = ((~n200gat)&(~n196gat));
assign n502gat = ((~II1079));
assign n2547gat = ((~n2550gat)&(~n2553gat)&(~n2554gat));
assign II4412 = ((~n2823gat));
assign II1374 = ((~n823gat));
assign II363 = ((~n335gat));
assign n1836gat = ((~n1695gat));
assign n647gat = ((~n2792gat)&(~n373gat));
assign n2487gat = ((~n2489gat));
assign n1250gat = ((~n1603gat)&(~n815gat));
assign II4732 = ((~n2825gat));
assign n2896gat = (n647gat)|(n441gat);
assign n2613gat = (n2614gat)|(n2615gat);
assign n1845gat = ((~n2141gat));
assign n794gat = ((~n852gat)&(~n2775gat));
assign n691gat = ((~II1439));
assign n1602gat = ((~n1594gat)&(~n1587gat)&(~n2989gat));
assign n2079gat = ((~n2078gat)&(~n2178gat)&(~n1990gat)&(~n2128gat));
assign n1842gat = ((~n1711gat));
assign n3135gat = ((~II4747));
assign n2959gat = (n1305gat)|(n1162gat);
assign II440 = ((~n340gat));
assign n1007gat = ((~n635gat));
assign n1417gat = ((~n2162gat)&(~n1480gat));
assign n1563gat = ((~n1561gat)&(~n1562gat)&(~n1659gat));
assign n709gat = (n710gat)|(n711gat)|(n712gat)|(n713gat);
assign II837 = ((~n860gat));
assign II199 = ((~n3085gat));
assign n1666gat = ((~n1986gat)&(~n2212gat)&(~n1991gat));
assign n2735gat = ((~II340));
assign n1580gat = ((~n1577gat));
assign n1519gat = ((~n1584gat)&(~n1339gat)&(~n1600gat));
assign II1201 = ((~n830gat));
assign n1077gat = ((~n110gat)&(~n2672gat));
assign n2212gat = ((~n2402gat));
assign n2009gat = ((~n2016gat)&(~n2664gat)&(~n2004gat));
assign II980 = ((~n1079gat));
assign n2388gat = ((~n2390gat));
assign n1734gat = ((~n1988gat)&(~n2212gat));
assign n591gat = ((~II1374));
assign n921gat = ((~n923gat));
assign n2516gat = ((~n2518gat));
assign n1866gat = ((~n1865gat));
assign n933gat = (n934gat)|(n935gat)|(n936gat)|(n937gat);
assign n793gat = ((~n2852gat)&(~n851gat));
assign n1974gat = ((~II3621));
assign n229gat = ((~II2153));
assign n2919gat = (n766gat)|(n760gat);
assign II2812 = (n1703gat)|(n1704gat)|(n1778gat);
assign n2259gat = ((~n3046gat));
assign n182gat = ((~n72gat)&(~n2720gat));
assign n879gat = ((~n2931gat)&(~n801gat));
assign n3028gat = ((~II3312));
assign II92 = ((~n919gat));
assign n2917gat = (n1074gat)|(n872gat);
assign n812gat = ((~II1348));
assign n969gat = ((~n219gat)&(~n2672gat));
assign n2877gat = (n139gat)|(n136gat);
assign n2794gat = ((~II97));
assign n2662gat = ((~n2660gat)&(~n2586gat));
assign n3104gat = ((~II4654));
assign n1113gat = ((~n393gat)&(~n701gat));
assign II1927 = ((~n1184gat));
assign n2992gat = (n1723gat)|(n1647gat)|(n1646gat);
assign n167gat = (n168gat)|(n169gat)|(n170gat)|(n171gat);
assign n1373gat = ((~n833gat)&(~n1442gat));
assign II3504 = ((~n2330gat));
assign n1112gat = ((~n630gat));
assign n705gat = ((~n707gat));
assign n47gat = ((~n53gat)&(~n51gat)&(~n50gat));
assign n273gat = ((~n341gat));
assign n2604gat = ((~n2611gat)&(~n2607gat)&(~n2610gat));
assign n1737gat = ((~n2212gat)&(~n2152gat));
assign n1179gat = ((~n2947gat));
assign n3115gat = ((~II4687));
assign II3312 = ((~n1699gat));
assign n343gat = (n344gat)|(n345gat)|(n346gat)|(n347gat);
assign n3013gat = (n2461gat)|(n2421gat);
assign n111gat = ((~n182gat));
assign II620 = ((~n160gat));
assign n2605gat = ((~n2611gat)&(~n2609gat)&(~n2608gat));
assign n2731gat = ((~n2733gat));
assign n828gat = ((~n830gat));
assign II480 = ((~n258gat));
assign II4654 = ((~n2819gat));
assign n1978gat = ((~n2286gat));
assign n244gat = ((~n334gat)&(~n386gat));
assign n2357gat = ((~n2285gat)&(~n2355gat)&(~n2443gat));
assign n2880gat = (n299gat)|(n207gat);
assign II2721 = (n1884gat)|(n1783gat)|(II2720);
assign n1963gat = ((~n2137gat));
assign n662gat = ((~n1725gat));
assign II5 = ((~n3087gat));
assign n11gat = ((~n12gat));
assign n2257gat = ((~n2189gat));
assign n1574gat = ((~n1719gat)&(~n1673gat)&(~n1444gat));
assign n334gat = ((~n1700gat));
assign n1884gat = ((~n1897gat));
assign II3742 = ((~n331gat));
assign n1700gat = ((~n1701gat)&(~n3023gat));
assign II2225 = ((~n2638gat));
assign n773gat = ((~n851gat)&(~n2838gat));
assign n189gat = ((~n286gat));
assign n3117gat = ((~II4693));
assign n2858gat = ((~II4129));
assign n2215gat = ((~n2346gat)&(~n2151gat)&(~n2402gat));
assign II2389 = ((~n2487gat));
assign n1199gat = ((~n1123gat)&(~n1284gat));
assign II3713 = ((~n2892gat));
assign n2934gat = (n1104gat)|(n887gat);
assign II423 = ((~n3068gat));
assign II1236 = ((~n612gat));
assign n2969gat = (n1323gat)|(n1264gat);
assign II2832 = (n1884gat)|(n1784gat)|(II2831);
assign n3112gat = ((~II4678));
assign II4372 = ((~n2817gat));
assign n1696gat = ((~n1707gat)&(~n1698gat));
assign n2696gat = ((~II3945));
assign n1097gat = ((~n270gat)&(~n741gat));
assign n2881gat = (n324gat)|(n238gat)|(n237gat);
assign II3297 = ((~n1699gat));
assign n1415gat = ((~n2081gat)&(~n2359gat));
assign n891gat = ((~n420gat)&(~n888gat));
assign n3129gat = ((~II4729));
assign n979gat = ((~n1601gat)&(~n926gat));
assign n1006gat = ((~n630gat));
assign n1054gat = ((~n1060gat)&(~n1058gat)&(~n1057gat));
assign n1279gat = ((~II1927));
assign II2014 = ((~n553gat));
assign n2439gat = ((~II2771));
assign n1970gat = ((~n1896gat));
assign n1564gat = ((~n1584gat)&(~n1719gat)&(~n1790gat)&(~n1576gat));
assign n1994gat = ((~n1719gat)&(~n1922gat));
assign n1082gat = ((~n375gat)&(~n380gat));
assign n1839gat = ((~n2138gat));
assign n3125gat = ((~II4717));
assign n2210gat = ((~n2401gat)&(~n2151gat));
assign n290gat = ((~n525gat));
assign n645gat = ((~n2792gat)&(~n93gat));
assign II1411 = ((~n881gat));
assign n2422gat = ((~n3013gat));
assign n447gat = ((~n2836gat)&(~n111gat));
assign n3002gat = (n2213gat)|(n2150gat)|(n2149gat);
assign n2201gat = ((~n2203gat));
assign n1818gat = ((~n1823gat)&(~n2005gat));
assign n2869gat = ((~II243));
assign n1786gat = ((~n2060gat));
assign n1231gat = ((~n1238gat)&(~n1234gat)&(~n1237gat));
assign n1484gat = ((~n2081gat)&(~n1528gat));
assign n38gat = ((~n151gat)&(~n233gat));
assign n1277gat = ((~II1920));
assign n792gat = ((~n2852gat)&(~n856gat));
assign n2820gat = ((~II4412));
assign n2205gat = ((~n2207gat));
assign n199gat = ((~n87gat));
assign n147gat = ((~II3904));
assign n1409gat = ((~n1476gat));
assign II977 = ((~n1080gat));
assign n2960gat = (n1175gat)|(n1174gat);
assign n295gat = ((~n357gat));
assign n2798gat = (n1032gat)|(n2054gat);
assign II1516 = (n2466gat)|(n2462gat)|(II1515);
assign n439gat = ((~n856gat)&(~n2836gat));
assign n1024gat = ((~n842gat));
assign n1954gat = ((~n3038gat));
assign n1287gat = ((~n1284gat)&(~n1195gat));
assign n510gat = ((~II1216));
assign n2941gat = (n1003gat)|(n902gat);
assign n1603gat = ((~n1831gat));
assign n2429gat = ((~n2541gat));
assign n2965gat = (n1267gat)|(n1257gat);
assign n1684gat = ((~n1759gat));
assign n2185gat = ((~n2261gat)&(~n2189gat));
assign n479gat = ((~n485gat)&(~n483gat)&(~n482gat));
assign II877 = ((~n1294gat));
assign n2829gat = ((~II4429));
assign n246gat = ((~n330gat)&(~n325gat)&(~n334gat));
assign n2878gat = (n234gat)|(n137gat);
assign n2752gat = ((~II4122));
assign n2101gat = ((~II1655));
assign n961gat = ((~n219gat)&(~n2734gat));
assign n2146gat = ((~n3002gat));
assign II3315 = ((~n1869gat));
assign n1000gat = ((~n419gat)&(~n1252gat));
assign II1439 = ((~n583gat));
assign n1421gat = ((~n2162gat)&(~n2359gat));
assign n1247gat = ((~n2958gat));
assign n2957gat = (n1159gat)|(n1158gat)|(n1156gat)|(n1155gat);
assign n2575gat = ((~II2228));
assign n196gat = ((~n297gat)&(~n195gat));
assign n2952gat = (n1076gat)|(n1075gat);
assign n501gat = ((~II1067));
assign n2671gat = ((~II18));
assign n262gat = ((~n268gat)&(~n266gat)&(~n265gat));
assign n2916gat = (n971gat)|(n970gat)|(n968gat);
assign n3111gat = ((~II4675));
assign n1152gat = ((~n926gat)&(~n1150gat));
assign n1533gat = ((~n1524gat)&(~n1403gat));
assign II4717 = ((~n2763gat));
assign II23 = ((~n3081gat));
assign n3040gat = ((~II3472));
assign n1266gat = ((~n2965gat)&(~n1253gat));
assign n1918gat = ((~n2392gat));
assign II3148 = (n1839gat)|(n1884gat)|(n1784gat);
assign n2681gat = ((~II4489));
assign n1798gat = ((~n1739gat)&(~n1673gat));
assign II712 = ((~n274gat));
assign n312gat = ((~n314gat));
assign n2692gat = ((~II3948));
assign n2162gat = ((~n2220gat));
assign n64gat = ((~II749));
assign n1762gat = ((~II1683));
assign II1035 = ((~n944gat));
assign n2894gat = (n443gat)|(n439gat);
assign n228gat = ((~II2148));
assign n978gat = ((~n2944gat)&(~n2945gat));
assign n2150gat = ((~n2401gat)&(~n2346gat));
assign n1787gat = ((~n2141gat));
assign n2853gat = ((~II885));
assign n689gat = ((~n696gat)&(~n692gat)&(~n695gat));
assign II3801 = ((~n2925gat));
assign n240gat = ((~n255gat)&(~n140gat));
assign n2883gat = (n251gat)|(n244gat);
assign n2413gat = ((~n2419gat)&(~n2417gat)&(~n2416gat));
assign n1888gat = ((~n3039gat));
assign II2953 = ((~n2179gat));
assign n729gat = ((~n733gat)&(~n734gat)&(~n735gat));
assign n2430gat = ((~n2533gat)&(~n2486gat)&(~n2429gat));
assign n965gat = ((~n2711gat)&(~n851gat));
assign II259 = ((~n3086gat));
assign II337 = ((~n3066gat));
assign n521gat = ((~n740gat)&(~n2715gat));
assign n1075gat = ((~n855gat));
assign II1476 = ((~n697gat));
assign n1609gat = ((~n1503gat)&(~n3025gat));
assign II2181 = ((~n779gat));
assign n2718gat = ((~n2719gat));
assign n3126gat = ((~II4720));
assign n968gat = ((~n2789gat)&(~n219gat));
assign n79gat = ((~n86gat));
assign II206 = ((~n3084gat));
assign n1334gat = ((~n1336gat));
assign n2674gat = ((~II381));
assign II4678 = ((~n2697gat));
assign n989gat = ((~n721gat)&(~n741gat));
assign n128gat = ((~II2174));
assign n2564gat = ((~n2352gat));
assign n2342gat = ((~II1550));
assign n141gat = ((~n155gat)&(~n253gat)&(~n150gat));
assign n1861gat = ((~n1866gat)&(~n2216gat)&(~n1988gat));
assign n1185gat = ((~n1189gat)&(~n1190gat)&(~n1191gat));
assign II4626 = ((~n1871gat));
assign n526gat = ((~n2859gat)&(~n740gat));
assign n1305gat = ((~n1147gat)&(~n1590gat));
assign n741gat = ((~n629gat));
assign n1468gat = ((~n1519gat));
assign n2387gat = ((~n2056gat)&(~n2437gat));
assign n975gat = ((~n111gat)&(~n2852gat));
assign n795gat = ((~n2731gat)&(~n852gat));
assign n356gat = ((~n2726gat)&(~n740gat));
assign n2286gat = ((~II1585));
assign n1105gat = ((~n2934gat));
assign n2923gat = (n1082gat)|(n796gat);
assign n181gat = ((~n286gat)&(~n179gat)&(~n188gat));
assign n1778gat = ((~n3026gat)&(~n1779gat));
assign II1894 = ((~n1044gat));
assign n405gat = ((~n728gat));
assign n1530gat = ((~n2364gat));
assign n2793gat = ((~II100));
assign n732gat = ((~n738gat)&(~n736gat)&(~n735gat));
assign n2570gat = ((~n2573gat)&(~n2576gat)&(~n2577gat));
assign II675 = ((~n1025gat));
assign n803gat = (n804gat)|(n805gat)|(n806gat)|(n807gat);
assign II2316 = ((~n2390gat));
assign n1769gat = ((~n1771gat));
assign n2292gat = ((~n2443gat)&(~n2284gat)&(~n2285gat));
assign II2040 = ((~n551gat));
assign II4747 = ((~n2816gat));
assign n76gat = ((~n82gat));
assign II4485 = ((~n2682gat));
assign n2574gat = ((~II2225));
assign n2603gat = ((~n2606gat)&(~n2609gat)&(~n2610gat));
assign n2874gat = (n141gat)|(n38gat)|(n37gat);
assign n1500gat = ((~n1113gat));
assign II3056 = ((~n1312gat));
assign n324gat = ((~n255gat)&(~n146gat)&(~n241gat));
assign n1018gat = ((~II378));
assign II634 = ((~n337gat));
assign n1372gat = ((~n282gat)&(~n1444gat));
assign n498gat = ((~II1230));
assign n3018gat = ((~II3211));
assign n62gat = ((~II741));
assign n1642gat = ((~n1559gat)&(~n1616gat)&(~n1645gat));
assign n2949gat = (n1101gat)|(n996gat);
assign n2338gat = ((~II2344));
assign n2688gat = ((~II4496));
assign n808gat = ((~II1305));
assign n2904gat = (n793gat)|(n664gat)|(n556gat);
assign n800gat = ((~n2874gat));
assign n1849gat = ((~II2731));
assign n1378gat = ((~n2975gat));
assign n2673gat = ((~II384));
assign n2548gat = ((~n2555gat)&(~n2551gat)&(~n2554gat));
assign II812 = ((~n957gat));
assign n814gat = ((~n816gat));
assign n1369gat = ((~n2966gat));
assign n2470gat = ((~n2472gat));
assign II4623 = ((~n2806gat));
assign n1471gat = ((~n1334gat)&(~n1858gat)&(~n1604gat));
assign II2109 = ((~n322gat));
assign II2177 = ((~n221gat));
assign n2199gat = ((~n2147gat));
assign II4194 = ((~n1462gat));
assign II3513 = ((~n2439gat));
assign II3831 = ((~n384gat));
assign II1115 = ((~n624gat));
assign n2719gat = ((~II776));
assign n1264gat = ((~n1006gat)&(~n617gat));
assign n1447gat = ((~n1117gat));
assign n2809gat = ((~II4642));
assign n2392gat = ((~n2394gat));
assign n1055gat = ((~II958));
assign II1243 = ((~n404gat));
assign II999 = ((~n1148gat));
assign n145gat = ((~n144gat)&(~n325gat));
assign II473 = ((~n162gat));
assign n739gat = ((~n850gat));
assign n1280gat = ((~n1282gat));
assign II2837 = ((~n2347gat));
assign n2042gat = ((~n2044gat));
assign II4023 = (n2443gat)|(n2290gat)|(n2214gat);
assign n2805gat = ((~II4630));
assign n34gat = ((~n221gat));
assign n3054gat = ((~II3660));
assign n82gat = ((~n16gat)&(~n295gat)&(~n637gat));
assign II1174 = ((~n705gat));
assign n1244gat = ((~n1123gat)&(~n1134gat));
assign n249gat = ((~n386gat)&(~n330gat));
assign n2253gat = ((~n2189gat));
assign n818gat = ((~n820gat));
assign n2891gat = (n795gat)|(n656gat)|(n368gat);
assign n289gat = ((~n563gat));
assign n1546gat = ((~n2980gat));
assign II1807 = ((~n1183gat));
assign n382gat = ((~n384gat));
assign n2953gat = (n1163gat)|(n1102gat);
assign n565gat = ((~n586gat));
assign n759gat = ((~n855gat));
assign n2747gat = ((~n2751gat));
assign n909gat = ((~n916gat)&(~n912gat)&(~n915gat));
assign n1239gat = ((~n1241gat));
assign n287gat = ((~n289gat)&(~n2715gat));
assign n1201gat = (n1202gat)|(n1203gat)|(n1204gat)|(n1205gat);
assign n1608gat = ((~n1704gat)&(~n1703gat));
assign n1855gat = ((~n2014gat));
assign n2317gat = ((~n2319gat));
assign II4530 = ((~n2756gat));
assign II1138 = ((~n834gat));
assign n1446gat = ((~n1318gat));
assign n2677gat = ((~II4492));
assign n737gat = ((~II1115));
assign n1431gat = ((~n1433gat));
assign n2402gat = ((~II2843));
assign n1160gat = ((~n1484gat));
assign n1159gat = ((~n1160gat)&(~n1084gat));
assign n2252gat = ((~n2260gat));
assign II4753 = ((~n2811gat));
assign n392gat = ((~n398gat));
assign n948gat = ((~n954gat)&(~n952gat)&(~n951gat));
assign II4105 = ((~n1456gat));
assign II3412 = ((~n2057gat));
assign n2862gat = ((~n2864gat));
assign n1070gat = ((~n1072gat));
assign n1232gat = ((~n1238gat)&(~n1236gat)&(~n1235gat));
assign n3011gat = (n2333gat)|(n2331gat);
assign n1017gat = ((~n1023gat)&(~n1021gat)&(~n1020gat));
assign n2925gat = (n975gat)|(n972gat)|(n969gat);
assign n1705gat = ((~n1619gat));
assign n51gat = ((~II473));
assign II1248 = ((~n405gat));
assign n677gat = ((~n803gat));
assign n1773gat = ((~n1775gat));
assign n2924gat = (n871gat)|(n797gat);
assign n2895gat = (n444gat)|(n440gat);
assign n664gat = ((~n1725gat));
assign II851 = ((~n1066gat));
assign n1091gat = ((~n1111gat)&(~n956gat));
assign II936 = ((~n1228gat));
assign n1359gat = ((~n1436gat)&(~n1106gat));
assign n2921gat = (n966gat)|(n790gat);
assign II1121 = ((~n621gat));
assign n1707gat = ((~n1626gat));
assign n1794gat = ((~n1673gat)&(~n1719gat));
assign n3062gat = ((~II3876));
assign II2400 = ((~n2601gat));
assign n354gat = ((~n411gat)&(~n522gat));
assign n84gat = ((~n296gat)&(~n17gat)&(~n294gat));
assign n743gat = ((~n746gat));
assign II2890 = (n1788gat)|(n1786gat)|(II2889);
assign II230 = ((~n2855gat));
assign n1819gat = ((~n1821gat));
assign n1571gat = ((~n1670gat)&(~n1658gat)&(~n1797gat));
assign n69gat = ((~n68gat));
assign n1738gat = ((~n1740gat));
assign n1699gat = ((~n2452gat));
assign n888gat = ((~n2933gat));
assign n938gat = ((~II858));
assign n776gat = ((~II2032));
assign II1399 = ((~n883gat));
assign n2727gat = ((~II264));
assign II3303 = ((~n1691gat));
assign II300 = ((~n2733gat));
assign n1253gat = ((~n930gat)&(~n1123gat));
assign n2899gat = (n772gat)|(n451gat)|(n446gat);
assign n524gat = ((~n414gat));
assign II2145 = ((~n314gat));
assign n2734gat = ((~n2736gat));
assign n517gat = ((~n518gat));
assign n2840gat = ((~n2841gat));
assign n3059gat = ((~II3801));
assign n578gat = ((~n580gat));
assign n840gat = ((~n842gat));
assign n2843gat = ((~II985));
assign n1216gat = ((~n1223gat)&(~n1219gat)&(~n1222gat));
assign n2354gat = ((~n2201gat));
assign n3057gat = ((~II3754));
assign n2436gat = ((~n2437gat)&(~n1892gat));
assign n1507gat = ((~II3163));
assign n1760gat = ((~n1681gat)&(~n1602gat)&(~n2985gat));
assign n1543gat = ((~n1606gat));
assign II3765 = ((~n2929gat));
assign n1590gat = ((~n1603gat));
assign n954gat = ((~II851));
assign II1899 = ((~n1133gat));
assign n2405gat = ((~n2407gat));
assign n2897gat = (n648gat)|(n442gat);
assign n143gat = ((~n326gat)&(~n247gat));
assign II443 = ((~n702gat));
assign n2785gat = ((~II583));
assign II834 = ((~n861gat));
assign n2937gat = (n900gat)|(n895gat);
assign n1235gat = ((~II916));
assign II1683 = ((~n1763gat));
assign n1677gat = ((~II3191));
assign n2758gat = ((~II4117));
assign n1051gat = ((~n1055gat)&(~n1056gat)&(~n1057gat));
assign II3891 = ((~n2924gat));
assign II426 = ((~n2780gat));
assign n949gat = ((~II793));
assign n44gat = ((~n48gat)&(~n49gat)&(~n50gat));
assign II1031 = ((~n1050gat));
assign n2763gat = ((~II4506));
assign n2704gat = (n11gat)|(n1889gat);
assign II3465 = ((~n1886gat));
assign n3146gat = ((~II4780));
assign n735gat = ((~II1127));
assign n2926gat = (n1083gat)|(n1077gat);
assign n333gat = ((~n2883gat));
assign n987gat = ((~n741gat)&(~n159gat));
assign n2048gat = ((~n2994gat));
assign n2406gat = ((~II2785));
assign n3060gat = ((~II3817));
assign n231gat = ((~II2162));
assign n1189gat = ((~II1752));
assign II4554 = ((~n2741gat));
assign II815 = ((~n956gat));
assign n929gat = ((~n931gat));
assign n829gat = ((~II1201));
assign n1598gat = ((~n1592gat)&(~n2422gat));
assign n503gat = ((~II1236));
assign n2572gat = ((~n2578gat)&(~n2576gat)&(~n2575gat));
assign II4349 = ((~n2935gat));
assign n1311gat = ((~II3056));
assign n620gat = ((~n846gat));
assign n1968gat = ((~n1958gat));
assign II1402 = ((~n882gat));
assign n1248gat = ((~n2954gat));
assign n1717gat = ((~II2926));
assign II30 = ((~n2668gat));
assign n634gat = ((~n418gat)&(~n521gat));
assign II1481 = ((~n582gat));
assign n408gat = ((~n516gat)&(~n407gat));
assign n1742gat = ((~n2216gat));
assign n1114gat = ((~n725gat)&(~n721gat));
assign II1155 = ((~n706gat));
assign n2988gat = (n1733gat)|(n1581gat);
assign II958 = ((~n864gat));
assign n1757gat = ((~n1773gat)&(~n1769gat));
assign n321gat = ((~II2109));
assign n1593gat = ((~n1551gat)&(~n1310gat));
assign n1505gat = ((~n2980gat));
assign n150gat = ((~n152gat));
assign n1269gat = (n1270gat)|(n1271gat)|(n1272gat)|(n1273gat);
assign n59gat = ((~n65gat)&(~n63gat)&(~n62gat));
assign n1031gat = ((~n1002gat)&(~n455gat));
assign n1101gat = ((~n1590gat)&(~n1293gat));
assign n1059gat = ((~II1011));
assign n1487gat = ((~n1485gat));
assign n863gat = ((~n865gat));
assign n3000gat = (n2000gat)|(n1999gat);
assign n329gat = ((~n331gat));
assign n2819gat = ((~II4651));
assign n2202gat = ((~II2260));
assign n459gat = ((~n457gat)&(~n461gat));
assign n1567gat = ((~n1634gat)&(~n1735gat));
assign II1023 = ((~n928gat));
assign n3037gat = ((~II3457));
assign n2158gat = ((~n1412gat));
assign n1411gat = ((~n1154gat)&(~n1608gat));
assign n3023gat = ((~II3297));
assign n2189gat = ((~II2978));
assign II368 = ((~n269gat));
assign n767gat = ((~n219gat)&(~n2731gat));
assign n484gat = ((~II456));
assign n1338gat = ((~n1340gat));
assign n1630gat = ((~n1895gat)&(~n1631gat));
assign n164gat = ((~II620));
assign n2781gat = ((~n2783gat));
assign n200gat = ((~n199gat)&(~n92gat));
assign n760gat = ((~n855gat));
assign n877gat = ((~n875gat)&(~n876gat));
assign n1182gat = ((~n1180gat)&(~n455gat));
assign n2695gat = (n1586gat)|(n1791gat);
assign n1629gat = ((~n1895gat));
assign II1999 = ((~n658gat));
assign II4524 = ((~n2757gat));
assign n2956gat = (n1178gat)|(n1116gat);
assign n1576gat = ((~n2351gat)&(~n1988gat)&(~n1661gat));
assign n2601gat = (n2602gat)|(n2603gat)|(n2604gat)|(n2605gat);
assign II4332 = ((~n2813gat));
assign n2060gat = ((~II2684));
assign n1011gat = ((~n455gat)&(~n898gat));
assign n2738gat = ((~II4548));
assign n2002gat = ((~n2008gat));
assign n2595gat = ((~n2594gat));
assign n1557gat = ((~n1553gat)&(~n1645gat)&(~n1614gat));
assign n420gat = ((~n408gat)&(~n359gat));
assign II1 = ((~n3088gat));
assign n1318gat = ((~n392gat)&(~n701gat));
assign II4506 = ((~n2764gat));
assign n195gat = ((~n184gat));
assign n1647gat = ((~n1656gat)&(~n1659gat)&(~n1554gat));
assign n2767gat = ((~II14));
assign n2097gat = ((~n2099gat));
assign n2625gat = ((~II1703));
assign II1786 = ((~n1071gat));
assign n1710gat = ((~n1709gat)&(~n1629gat));
assign n142gat = ((~n382gat)&(~n326gat)&(~n144gat));
assign n1016gat = ((~n1023gat)&(~n1019gat)&(~n1022gat));
assign II4798 = ((~n2707gat));
assign n1566gat = ((~n1605gat));
assign n2493gat = ((~n2495gat));
assign n1783gat = ((~n1848gat));
assign n2868gat = ((~II248));
assign n2432gat = ((~n2430gat));
assign n1357gat = ((~n1424gat)&(~n1309gat));
assign n1490gat = ((~n1430gat));
assign n2211gat = ((~n2193gat)&(~n2402gat));
assign n264gat = ((~II334));
assign II734 = ((~n273gat));
assign n1614gat = ((~n396gat)&(~n845gat));
assign n3063gat = ((~II3891));
assign II1496 = ((~n686gat));
assign n2964gat = (n1304gat)|(n1249gat);
assign II863 = ((~n3080gat));
assign n1624gat = ((~n1319gat)&(~n1379gat));
assign n2410gat = ((~n2414gat)&(~n2415gat)&(~n2416gat));
assign n1923gat = ((~n1864gat));
assign n1403gat = ((~n1402gat));
assign II3904 = ((~n148gat));
assign II1791 = ((~n1119gat));
assign n1268gat = ((~n1201gat));
assign n2760gat = ((~II4512));
assign n2682gat = ((~II4482));
assign n92gat = ((~n2785gat));
assign n2284gat = ((~n2342gat));
assign n2779gat = ((~II426));
assign II1923 = ((~n1201gat));
assign n1274gat = ((~II1807));
assign n3138gat = ((~II4756));
assign n576gat = ((~II1496));
assign n1846gat = ((~n1845gat)&(~n1893gat));
assign n1257gat = ((~n1007gat)&(~n274gat));
assign n2855gat = ((~II227));
assign n2750gat = (n1181gat)|(n2243gat);
assign n197gat = ((~n194gat)&(~n297gat));
assign n1782gat = ((~n2971gat));
assign n514gat = ((~II1255));
assign II2873 = ((~n1496gat));
assign II1874 = ((~n1135gat));
assign n1618gat = ((~n1319gat)&(~n1447gat));
assign n421gat = ((~n2715gat)&(~n2723gat));
assign II4222 = ((~n1761gat));
assign n1732gat = ((~n1515gat)&(~n1736gat)&(~n1658gat));
assign n1556gat = ((~n1614gat)&(~n1645gat)&(~n1616gat));
assign n325gat = ((~n327gat));
assign n355gat = ((~n517gat)&(~n410gat)&(~n354gat));
assign n509gat = ((~II1190));
assign n2836gat = ((~n2837gat));
assign n469gat = ((~II3867));
assign n1414gat = ((~n1415gat));
assign II3882 = ((~n256gat));
assign II776 = ((~n3074gat));
assign II651 = ((~n281gat));
assign II76 = ((~n402gat));
assign n2699gat = ((~n2703gat));
assign n2220gat = ((~n2290gat)&(~n2217gat));
assign n1587gat = ((~II4212));
assign n736gat = ((~II1209));
assign n468gat = ((~n470gat));
assign n2414gat = ((~II2254));
assign n2931gat = (n1100gat)|(n994gat)|(n989gat)|(n880gat);
assign n1155gat = ((~n1085gat)&(~n1348gat));
assign II4681 = ((~n2698gat));
assign II2213 = ((~n2342gat));
assign n815gat = ((~II1319));
assign n449gat = ((~n2836gat)&(~n851gat));
assign n587gat = ((~n591gat)&(~n592gat)&(~n593gat));
assign n2291gat = ((~n2353gat)&(~n2355gat)&(~n2443gat));
assign II749 = ((~n343gat));
assign n1356gat = ((~n1354gat));
assign n3145gat = ((~II4777));
assign II381 = ((~n3073gat));
assign n738gat = ((~II1103));
assign n1714gat = ((~II3149));
assign n3116gat = ((~II4690));
assign n2736gat = ((~II337));
assign n49gat = ((~II420));
assign II1833 = ((~n1226gat));
assign n2670gat = ((~II81));
assign II1961 = ((~n2516gat));
assign n1578gat = ((~n2152gat)&(~n2351gat)&(~n1665gat));
assign n789gat = ((~II2049));
assign n656gat = ((~n851gat)&(~n2718gat));
assign n2345gat = ((~n2347gat));
assign II240 = ((~n2717gat));
assign n2668gat = ((~II27));
assign n2890gat = (n654gat)|(n557gat)|(n371gat);
assign n1774gat = ((~II3339));
assign n184gat = ((~n189gat)&(~n188gat)&(~n179gat));
assign n1207gat = ((~II1877));
assign II4580 = ((~n2702gat));
assign n1350gat = ((~n1831gat));
assign n2073gat = ((~n2078gat)&(~n1990gat)&(~n2181gat));
assign n2332gat = ((~n3045gat));
assign n1726gat = ((~n2992gat)&(~n2986gat)&(~n2991gat));
assign n2780gat = ((~II423));
assign n1306gat = ((~n2964gat));
assign n943gat = ((~II1035));
assign II3336 = ((~n2040gat));
assign n1921gat = ((~n1738gat)&(~n1673gat));
assign n1260gat = ((~n1007gat)&(~n278gat));
assign n476gat = ((~n480gat)&(~n481gat)&(~n482gat));
assign n266gat = ((~II359));
assign n849gat = ((~n924gat));
assign n3123gat = ((~II4711));
assign n313gat = ((~II2145));
assign II1488 = ((~n456gat));
assign II1348 = ((~n578gat));
assign II2672 = ((~n2143gat));
assign n1200gat = ((~n1120gat)&(~n1123gat));
assign n423gat = ((~n2724gat)&(~n2726gat));
assign II1464 = ((~n699gat));
assign II4768 = ((~n2755gat));
assign n1004gat = ((~n978gat)&(~n420gat));
assign n397gat = ((~II718));
assign II1472 = ((~n682gat));
assign II3178 = (n1838gat)|(n1785gat)|(n1788gat);
assign n1460gat = ((~n1462gat));
assign n377gat = ((~n110gat)&(~n2778gat));
assign n1581gat = ((~n1858gat)&(~n1580gat));
assign II1085 = ((~n617gat));
assign n2823gat = ((~II4409));
assign n1103gat = ((~n956gat)&(~n1590gat));
assign n1595gat = ((~II4185));
assign II1857 = ((~n931gat));
assign n2936gat = (n901gat)|(n893gat);
assign n2124gat = ((~II3587));
assign II1339 = ((~n579gat));
assign n380gat = ((~n2881gat));
assign n86gat = ((~n743gat)&(~n294gat)&(~n17gat));
assign n2401gat = ((~n2403gat));
assign n1653gat = ((~n1651gat)&(~n1652gat)&(~n1659gat));
assign II2433 = ((~n2628gat));
assign n1208gat = ((~II1894));
assign n2846gat = ((~n2847gat));
assign n362gat = ((~n2723gat)&(~n2727gat));
assign n2905gat = (n964gat)|(n961gat);
assign n1367gat = ((~n1366gat)&(~n1374gat));
assign n678gat = ((~n680gat));
assign II4774 = ((~n2740gat));
assign n2246gat = ((~n933gat));
assign n396gat = ((~n398gat));
assign n2397gat = ((~n2399gat));
assign II2254 = ((~n2206gat));
assign n1929gat = ((~n1758gat)&(~n1790gat));
assign II1584 = (n2353gat)|(n2284gat)|(n2354gat);
assign n2751gat = ((~II4222));
assign n939gat = ((~II936));
assign n1328gat = ((~n1224gat));
assign n2826gat = ((~II4432));
assign n1800gat = ((~n1635gat)&(~n1919gat));
assign n3132gat = ((~II4738));
assign n1211gat = ((~II1908));
assign II3300 = ((~n1699gat));
assign II351 = ((~n337gat));
assign II3290 = ((~n1691gat));
assign n2554gat = ((~II2428));
assign n3136gat = ((~II4750));
assign n1302gat = ((~n1300gat)&(~n1487gat));
assign n2861gat = ((~II199));
assign n1228gat = (n1229gat)|(n1230gat)|(n1231gat)|(n1232gat);
assign n2650gat = ((~n2649gat)&(~n2652gat));
assign n981gat = ((~n926gat)&(~n873gat));
assign n806gat = ((~n813gat)&(~n809gat)&(~n812gat));
assign II715 = ((~n401gat));
assign n2195gat = ((~n2200gat)&(~n1855gat));
assign n2492gat = ((~n2329gat));
assign n984gat = ((~n926gat)&(~n983gat));
assign n2892gat = (n378gat)|(n377gat);
assign n2792gat = ((~n2794gat));
assign n2426gat = ((~n2480gat));
assign n461gat = ((~n463gat));
assign II4145 = (n1788gat)|(n1784gat)|(II4144);
assign II4573 = ((~n2693gat));
assign n506gat = ((~n509gat)&(~n512gat)&(~n513gat));
assign n712gat = ((~n719gat)&(~n715gat)&(~n718gat));
assign n1988gat = ((~n2345gat));
assign II2720 = (n1788gat)|(n1786gat)|(n1839gat);
assign II3948 = ((~n2696gat));
assign n1523gat = ((~n2219gat));
assign n2545gat = (n2546gat)|(n2547gat)|(n2548gat)|(n2549gat);
assign n1186gat = ((~n1189gat)&(~n1192gat)&(~n1193gat));
assign n752gat = ((~n758gat)&(~n756gat)&(~n755gat));
assign n407gat = ((~n355gat));
assign n687gat = ((~n691gat)&(~n692gat)&(~n693gat));
assign n2283gat = ((~n2438gat));
assign II2417 = ((~n2633gat));
assign n903gat = ((~n1007gat)&(~n397gat));
assign II796 = ((~n3076gat));
assign n1366gat = ((~n1365gat));
assign n1028gat = ((~n455gat)&(~n879gat));
assign n2730gat = ((~II509));
assign n1368gat = ((~n1442gat)&(~n613gat));
assign II3494 = ((~n1963gat));
assign II4352 = ((~n2818gat));
assign n1669gat = ((~n1668gat)&(~n1742gat)&(~n1670gat));
assign n269gat = ((~n271gat));
assign n2724gat = ((~II256));
assign n2576gat = ((~II2235));
assign II237 = ((~n640gat));
assign n2691gat = ((~n2695gat));
assign II1515 = (n2474gat)|(n2524gat)|(n2831gat);
assign n630gat = ((~n634gat)&(~n523gat)&(~n524gat));
assign n3131gat = ((~II4735));
assign n2967gat = (n1262gat)|(n1260gat);
assign n785gat = ((~II2017));
assign II1209 = ((~n828gat));
assign n1553gat = ((~n1616gat));
assign n1001gat = ((~n420gat)&(~n1002gat));
assign II4409 = ((~n2938gat));
assign n2293gat = ((~n2353gat)&(~n2284gat)&(~n2443gat));
assign n3014gat = (n2567gat)|(n2499gat);
assign n906gat = (n907gat)|(n908gat)|(n909gat)|(n910gat);
assign n2147gat = ((~n2988gat)&(~n1855gat));
assign n1607gat = ((~n2082gat)&(~n1609gat));
assign n361gat = ((~n2859gat)&(~n2726gat));
assign n867gat = ((~n219gat)&(~n2775gat));
assign n2206gat = ((~II2251));
assign n177gat = ((~II651));
assign n1562gat = ((~n1556gat));
assign II2731 = ((~n1850gat));
assign n1599gat = ((~n1691gat)&(~n336gat));
assign n455gat = ((~n291gat));
assign n2797gat = ((~II4020));
assign n1083gat = ((~n381gat)&(~n375gat));
assign n512gat = ((~II1248));
assign n1641gat = ((~n1645gat)&(~n1553gat)&(~n1559gat));
assign II3941 = ((~n2684gat));
assign n2762gat = (n1028gat)|(n1782gat);
assign n1827gat = ((~n2729gat)&(~n2317gat));
assign II1322 = ((~n815gat));
assign n2737gat = ((~II4554));
assign n2460gat = ((~n666gat)&(~n120gat));
assign n1898gat = ((~II3174));
assign n1673gat = ((~n2989gat));
assign n1922gat = ((~n1798gat));
assign n255gat = ((~II3882));
assign n1632gat = ((~II4145));
assign n1785gat = ((~n2059gat));
assign n2520gat = ((~n2522gat));
assign II1630 = ((~n2630gat));
assign n294gat = ((~n360gat));
assign n2163gat = ((~n1790gat)&(~n1310gat)&(~n2664gat)&(~n2168gat));
assign n2615gat = ((~n2617gat)&(~n2619gat));
assign n2830gat = (n2444gat)|(n1754gat);
assign n2768gat = ((~II11));
assign n3124gat = ((~II4714));
assign n924gat = ((~n1070gat));
assign n633gat = ((~n634gat));
assign n291gat = ((~n290gat)&(~n292gat));
assign II3539 = ((~n2198gat));
assign n1869gat = ((~n1871gat));
assign n1840gat = ((~n1892gat));
assign n1865gat = ((~n1989gat)&(~n1918gat)&(~n1986gat));
assign II1336 = ((~n580gat));
assign n1646gat = ((~n1569gat)&(~n1659gat)&(~n1566gat));
assign n1568gat = ((~n1575gat));
assign n373gat = ((~n2767gat));
assign n966gat = ((~n2789gat)&(~n373gat));
assign n1549gat = ((~II2832));
assign n1841gat = ((~n2058gat));
assign n583gat = ((~II1436));
assign n1709gat = ((~n1849gat));
assign n485gat = ((~II461));
assign n522gat = ((~n374gat)&(~n2859gat));
assign II4756 = ((~n2804gat));
assign n701gat = ((~n402gat));
assign n2686gat = ((~II4499));
assign n2996gat = (n1960gat)|(n1959gat)|(n1957gat);
assign n1379gat = ((~n1377gat));
assign II282 = ((~n1213gat));
assign n2027gat = ((~n2029gat));
assign n187gat = ((~n189gat)&(~n287gat)&(~n188gat));
assign n35gat = ((~n779gat));
assign n2141gat = ((~n2143gat));
assign n2642gat = ((~n2644gat));
assign n1635gat = ((~n1716gat));
assign n2893gat = (n391gat)|(n390gat);
assign II790 = ((~n1068gat));
assign n1686gat = ((~n1774gat)&(~n1869gat)&(~n1684gat));
assign n1651gat = ((~n1642gat));
assign n853gat = ((~n740gat)&(~n2148gat));
assign n1205gat = ((~n1211gat)&(~n1209gat)&(~n1208gat));
assign n928gat = ((~n1050gat));
assign n1466gat = ((~n1392gat)&(~n1461gat)&(~n1396gat));
assign n1897gat = ((~n1899gat));
assign II4496 = ((~n1708gat));
assign n1736gat = ((~n1737gat));
assign II4122 = ((~n1546gat));
assign n1467gat = ((~n2289gat)&(~n1468gat));
assign n1961gat = ((~n2996gat));
assign n3015gat = (n2566gat)|(n2565gat);
assign n2130gat = ((~n2134gat)&(~n2185gat));
assign n444gat = ((~n373gat)&(~n2781gat));
assign II4789 = ((~n2692gat));
assign n448gat = ((~n111gat)&(~n2846gat));
assign n915gat = ((~II687));
assign n1721gat = ((~n2442gat)&(~n1690gat)&(~n1978gat));
assign n1806gat = ((~II4081));
assign II50 = ((~n2783gat));
assign n881gat = ((~n883gat));
assign n2337gat = ((~n2339gat));
assign n2947gat = (n1094gat)|(n1093gat)|(n988gat)|(n984gat);
assign n1285gat = ((~n1196gat)&(~n1269gat));
assign n2008gat = ((~n2012gat)&(~n1774gat));
assign n1183gat = ((~n1184gat));
assign II3621 = ((~n1975gat));
assign n1419gat = ((~n2162gat)&(~n1479gat));
assign n2918gat = (n769gat)|(n759gat);
assign n1249gat = ((~n679gat)&(~n1603gat));
assign n651gat = ((~n93gat)&(~n2778gat));
assign n2728gat = ((~II259));
assign n406gat = ((~n516gat));
assign n369gat = ((~n1725gat));
assign n956gat = ((~II812));
assign n788gat = ((~II2044));
assign n1019gat = ((~II398));
assign II1667 = ((~n1880gat));
assign II4478 = ((~n2807gat));
assign n1894gat = ((~n1968gat)&(~n1891gat)&(~n1969gat));
assign n3049gat = ((~II3539));
assign n2427gat = ((~n2426gat)&(~n2153gat));
assign n2886gat = (n774gat)|(n764gat)|(n369gat);
assign n1831gat = ((~n1832gat)&(~n1765gat)&(~n1878gat));
assign n2417gat = ((~II2268));
assign n452gat = ((~n2885gat));
assign n1365gat = ((~n1479gat)&(~n1591gat));
assign n625gat = ((~II1124));
assign n3042gat = ((~II3491));
assign n1780gat = ((~n1777gat)&(~n1625gat)&(~n1626gat));
assign n2679gat = ((~II3954));
assign n1424gat = ((~n1420gat));
assign n2053gat = ((~n2393gat)&(~n2438gat));
assign n1486gat = ((~n1482gat)&(~n1591gat));
assign n1314gat = ((~n1316gat));
assign n1723gat = ((~n1659gat)&(~n1722gat)&(~n1724gat));
assign II4684 = ((~n2689gat));
assign n1351gat = ((~n1306gat)&(~n1353gat));
assign n1442gat = ((~n1831gat));
assign n1520gat = ((~n1582gat));
assign n3150gat = ((~II4792));
assign n3020gat = ((~II3287));
assign II1255 = ((~n709gat));
assign n586gat = (n587gat)|(n588gat)|(n589gat)|(n590gat);
assign II3957 = ((~n2450gat));
assign n2629gat = ((~II1630));
assign n222gat = ((~n226gat)&(~n227gat)&(~n228gat));
assign II4726 = ((~n2678gat));
assign II3635 = ((~n2558gat));
assign n2632gat = ((~n2634gat));
assign n1408gat = ((~n1507gat)&(~n1396gat)&(~n1393gat));
assign n2684gat = (n1599gat)|(n2051gat);
assign n2582gat = ((~II2248));
assign n1482gat = ((~n2363gat));
assign n2578gat = ((~II2242));
assign n400gat = ((~n402gat));
assign n2244gat = ((~n567gat));
assign n850gat = ((~n929gat));
assign n393gat = ((~II446));
assign n1374gat = ((~n2979gat));
assign n3025gat = ((~II3303));
assign II1795 = ((~n1070gat));
assign n2483gat = ((~n2537gat)&(~n2482gat)&(~n2486gat));
assign n1754gat = ((~n2449gat));
assign II2049 = ((~n657gat));
assign n1153gat = ((~n1414gat)&(~n566gat));
assign n1315gat = ((~II3342));
assign n856gat = ((~n2667gat));
assign II4227 = ((~n1760gat));
assign n1969gat = ((~n2142gat));
assign n774gat = ((~n2842gat)&(~n851gat));
assign II3520 = ((~n2498gat));
assign n2200gat = ((~n2078gat));
assign n2055gat = ((~n1891gat)&(~n1958gat));
assign n345gat = ((~n348gat)&(~n351gat)&(~n352gat));
assign n263gat = ((~II314));
assign II1002 = ((~n1147gat));
assign n555gat = ((~n852gat)&(~n2792gat));
assign n2815gat = ((~II4372));
assign n2938gat = (n899gat)|(n896gat);
assign II4329 = ((~n2950gat));
assign II3339 = ((~n1775gat));
assign n1882gat = ((~n2124gat)&(~n2115gat)&(~n2239gat));
assign n2057gat = ((~n2049gat)&(~n1855gat));
assign II672 = ((~n842gat));
assign n1352gat = ((~n1248gat)&(~n1418gat));
assign n1416gat = ((~n2081gat)&(~n1480gat));
assign n2841gat = ((~II963));
assign II3808 = ((~n327gat));
assign n375gat = ((~n110gat));
assign n2571gat = ((~n2578gat)&(~n2574gat)&(~n2577gat));
assign n666gat = ((~II1981));
assign n1320gat = ((~n1444gat)&(~n278gat));
assign n2616gat = ((~II2400));
assign n3035gat = ((~II3412));
assign n2933gat = (n981gat)|(n890gat)|(n889gat)|(n886gat);
assign n1458gat = ((~n1510gat)&(~n1459gat));
assign n2131gat = ((~n2185gat));
assign n1259gat = ((~n2967gat)&(~n1251gat));
assign n1010gat = ((~n897gat)&(~n455gat));
assign n2987gat = (n1574gat)|(n1573gat);
assign n2193gat = ((~n2393gat)&(~n2439gat));
assign II243 = ((~n3089gat));
assign n1376gat = ((~n724gat)&(~n720gat));
assign n563gat = ((~II1278));
assign n89gat = ((~n88gat)&(~n2784gat));
assign n1848gat = ((~n1850gat));
assign n1348gat = ((~n1349gat));
assign n1727gat = ((~n1728gat));
assign n78gat = ((~n2784gat)&(~n79gat));
assign n2129gat = ((~n2189gat)&(~n2134gat)&(~n2261gat));
assign n1308gat = ((~n2081gat)&(~n1530gat));
assign n2054gat = ((~n2281gat));
assign II4024 = (n2353gat)|(n2284gat)|(II4023);
assign n1134gat = ((~II1874));
assign n2218gat = ((~n2214gat)&(~n2290gat));
assign II698 = ((~n906gat));
assign n2776gat = ((~II320));
assign n1060gat = ((~II1016));
assign n1428gat = ((~n2978gat)&(~n2982gat)&(~n2973gat)&(~n2977gat));
assign n1052gat = ((~n1055gat)&(~n1058gat)&(~n1059gat));
assign n1392gat = ((~n1394gat));
assign n2783gat = ((~II47));
assign n2885gat = (n250gat)|(n249gat)|(n248gat);
assign n1251gat = ((~n1123gat)&(~n1071gat));
assign n2983gat = (n2079gat)|(n2073gat);
assign n1625gat = ((~n3021gat)&(~n1628gat));
assign n976gat = ((~n628gat));
assign n364gat = ((~n366gat));
assign n944gat = (n945gat)|(n946gat)|(n947gat)|(n948gat);
assign n905gat = ((~n625gat)&(~n1006gat));
assign n2194gat = ((~n2187gat)&(~n1855gat));
assign n819gat = ((~II1385));
assign n169gat = ((~n172gat)&(~n175gat)&(~n176gat));
assign n73gat = ((~n67gat)&(~n2784gat));
assign n1816gat = ((~n1817gat));
assign n2804gat = ((~II4236));
assign n574gat = ((~II1488));
assign n2565gat = ((~n2352gat)&(~n2642gat));
assign II317 = ((~n3067gat));
assign n1412gat = ((~n1411gat)&(~n1406gat)&(~n2981gat));
assign n274gat = ((~II709));
assign n1111gat = ((~n635gat));
assign n1310gat = ((~n1312gat));
assign n1236gat = ((~II921));
assign II899 = ((~n1241gat));
assign n1972gat = ((~n1974gat)&(~n1970gat));
assign II4666 = ((~n2795gat));
assign n848gat = ((~n922gat));
assign n226gat = ((~II2112));
assign II4067 = ((~n1675gat));
assign n2423gat = ((~n665gat)&(~n1601gat));
assign n230gat = ((~II2157));
assign II44 = ((~n673gat));
assign II2238 = ((~n2560gat));
assign n188gat = ((~n288gat));
assign n690gat = ((~n696gat)&(~n694gat)&(~n693gat));
assign n2597gat = ((~n2599gat));
assign n2610gat = ((~II2389));
assign n2847gat = ((~II863));
assign n1889gat = ((~n1961gat));
assign n2556gat = ((~n1711gat)&(~n2437gat));
assign n3056gat = ((~II3713));
assign n927gat = ((~n1133gat));
assign II4651 = ((~n2822gat));
assign II2428 = ((~n2541gat));
assign n551gat = ((~n553gat));
assign n871gat = ((~n802gat)&(~n375gat));
assign n180gat = ((~n286gat)&(~n188gat)&(~n287gat));
assign n2499gat = ((~n2389gat)&(~n2494gat));
assign n223gat = ((~n226gat)&(~n229gat)&(~n230gat));
assign n42gat = ((~n475gat));
assign n1573gat = ((~n1444gat)&(~n1858gat)&(~n1635gat));
assign n2609gat = ((~II2385));
assign n2844gat = ((~n2845gat));
assign n572gat = ((~II1360));
assign n414gat = ((~n411gat)&(~n415gat));
assign n1703gat = ((~n1705gat)&(~n3028gat));
assign n2982gat = (n1504gat)|(n1502gat);
assign n997gat = ((~n741gat)&(~n393gat));
assign II4720 = ((~n2686gat));
assign II1216 = ((~n728gat));
assign n39gat = ((~n383gat)&(~n247gat));
assign n710gat = ((~n714gat)&(~n715gat)&(~n716gat));
assign n235gat = ((~n2878gat));
assign n993gat = ((~n1112gat)&(~n698gat));
assign n519gat = ((~n2854gat)&(~n374gat));
assign n1301gat = ((~n1416gat));
assign n1387gat = ((~n1389gat));
assign II572 = ((~n1829gat));
assign n357gat = ((~n2726gat)&(~n2860gat));
assign n353gat = ((~II734));
assign II3754 = ((~n2900gat));
assign II2017 = ((~n552gat));
assign n3143gat = ((~II4771));
assign n2990gat = (n1710gat)|(n1630gat);
assign n1430gat = ((~n1700gat));
assign n1494gat = ((~n1528gat)&(~n2162gat));
assign n589gat = ((~n596gat)&(~n592gat)&(~n595gat));
assign II921 = ((~n1239gat));
assign n1090gat = ((~n1111gat)&(~n860gat));
assign n964gat = ((~n111gat)&(~n2711gat));
assign n2951gat = (n1004gat)|(n1000gat);
assign n2740gat = ((~II4014));
assign n1094gat = ((~n1112gat)&(~n583gat));
assign II3174 = ((~n1899gat));
assign n751gat = ((~n758gat)&(~n754gat)&(~n757gat));
assign n2930gat = (n1153gat)|(n1151gat)|(n982gat)|(n877gat);
assign II941 = ((~n3077gat));
assign n1528gat = ((~n2293gat));
assign n2596gat = ((~n2665gat));
assign n2537gat = ((~n2538gat));
assign n1674gat = ((~II4067));
assign n1671gat = ((~n1669gat));
assign n1973gat = ((~n1975gat));
assign n885gat = ((~n579gat)&(~n1112gat));
assign II591 = ((~n3094gat));
assign n52gat = ((~II476));
assign n65gat = ((~II753));
assign n962gat = ((~n856gat)&(~n2711gat));
assign II4702 = ((~n2746gat));
assign n1722gat = ((~n1558gat));
assign II4744 = ((~n2815gat));
assign n2867gat = ((~n2869gat));
assign n2602gat = ((~n2606gat)&(~n2607gat)&(~n2608gat));
assign n2748gat = ((~n2752gat));
assign n1087gat = ((~n926gat)&(~n1084gat));
assign II3149 = (n1786gat)|(n1787gat)|(II3148);
assign n1864gat = ((~n1858gat)&(~n1495gat)&(~n2090gat));
assign II4452 = ((~n2828gat));
assign n988gat = ((~n340gat)&(~n741gat));
assign n1210gat = ((~II1903));
assign n1781gat = ((~n1780gat));
assign n896gat = ((~n897gat)&(~n420gat));
assign II1783 = ((~n1072gat));
assign n2766gat = ((~II4135));
assign II1908 = ((~n929gat));
assign n750gat = ((~n753gat)&(~n756gat)&(~n757gat));
assign n2352gat = ((~n3011gat)&(~n2215gat));
assign II4669 = ((~n2796gat));
assign n460gat = ((~n462gat)&(~n2884gat));
assign n1400gat = ((~n1674gat)&(~n1403gat));
assign II3191 = ((~n1678gat));
assign n590gat = ((~n596gat)&(~n594gat)&(~n593gat));
assign II768 = ((~n3090gat));
assign II1436 = ((~n584gat));
assign n2729gat = ((~II512));
assign n638gat = ((~n2715gat)&(~n2868gat));
assign n1498gat = ((~n1609gat)&(~n1427gat));
assign n2812gat = (n73gat)|(n70gat)|(n1840gat);
assign n1281gat = ((~II1837));
assign II3211 = ((~n2663gat));
assign n2573gat = ((~II2213));
assign n446gat = ((~n219gat)&(~n2781gat));
assign II171 = ((~n846gat));
assign II771 = ((~n2832gat));
assign II1467 = ((~n698gat));
assign II2989 = ((~n2135gat));
assign n1120gat = ((~II1766));
assign n1617gat = ((~n1319gat)&(~n1448gat));
assign n2946gat = (n1099gat)|(n998gat)|(n995gat)|(n980gat);
assign n441gat = ((~n856gat)&(~n2846gat));
assign II1407 = ((~n818gat));
assign n2903gat = (n794gat)|(n773gat)|(n662gat);
assign n50gat = ((~II468));
assign n2014gat = ((~n2035gat)&(~n2093gat)&(~n2018gat)&(~n2664gat));
assign n2633gat = ((~II2414));
assign n2531gat = ((~n2488gat)&(~n2625gat)&(~n2621gat));
assign n3050gat = ((~II3549));
assign n1029gat = ((~n978gat)&(~n455gat));
assign n3003gat = (n2256gat)|(n2251gat);
assign n2985gat = (n1686gat)|(n1533gat)|(n1532gat)|(n1531gat);
assign n1150gat = ((~n312gat));
assign n2119gat = ((~n2121gat));
assign n753gat = ((~II237));
assign n1117gat = ((~n720gat)&(~n725gat));
assign II2032 = ((~n777gat));
assign n1450gat = ((~n1423gat));
assign II741 = ((~n178gat));
assign n2419gat = ((~II2275));
assign n2389gat = ((~II2316));
assign n2197gat = ((~n2199gat)&(~n2281gat));
assign n2541gat = ((~n2543gat));
assign n893gat = ((~n894gat)&(~n420gat));
assign n297gat = ((~n2721gat));
assign n282gat = ((~II606));
assign II858 = ((~n857gat));
assign n1100gat = ((~n1297gat)&(~n1111gat));
assign n2720gat = ((~n2722gat));
assign n1477gat = ((~n2984gat));
assign n762gat = ((~n855gat));
assign n913gat = ((~II678));
assign II409 = ((~n720gat));
assign II2112 = ((~n321gat));
assign II1538 = ((~n2399gat));
assign n2646gat = (n2647gat)|(n2648gat);
assign II2696 = ((~n2139gat));
assign II4672 = ((~n2705gat));
assign II1891 = ((~n1045gat));
assign n365gat = ((~II2084));
assign II3951 = ((~n2448gat));
assign n3055gat = ((~II3703));
assign n1410gat = ((~n2357gat));
assign II4449 = ((~n2955gat));
assign n890gat = ((~n741gat)&(~n702gat));
assign n1246gat = ((~n864gat)&(~n1590gat));
assign n2011gat = ((~n2306gat));
assign n2808gat = ((~II4233));
assign n1234gat = ((~II902));
assign n2909gat = (n765gat)|(n643gat);
assign II2257 = ((~n2398gat));
assign n886gat = ((~n683gat)&(~n1112gat));
assign n2557gat = ((~n2621gat));
assign n2217gat = ((~n2206gat));
assign n852gat = ((~n854gat));
assign n1461gat = ((~II4194));
assign n991gat = ((~n1112gat)&(~n679gat));
assign n629gat = ((~n414gat)&(~n634gat)&(~n523gat));
assign n168gat = ((~n172gat)&(~n173gat)&(~n174gat));
assign n1157gat = ((~n1483gat));
assign n451gat = ((~n134gat)&(~n372gat));
assign n860gat = ((~II834));
assign II4432 = ((~n2829gat));
assign n2363gat = ((~n2353gat)&(~n2356gat)&(~n2355gat));
assign n2219gat = ((~n2354gat)&(~n2214gat));
assign n2667gat = ((~II30));
assign n1919gat = ((~n1860gat));
assign n2725gat = ((~II5));
assign n1203gat = ((~n1206gat)&(~n1209gat)&(~n1210gat));
assign n1643gat = ((~n1641gat));
assign n162gat = ((~n1013gat));
assign n3118gat = ((~II4696));
assign II4108 = ((~n1340gat));
assign n3130gat = ((~II4732));
assign n2732gat = ((~II300));
assign II4000 = (n2108gat)|(n2093gat)|(n2035gat)|(II3999);
assign II4117 = ((~n1505gat));
assign n1151gat = ((~n1301gat)&(~n1150gat));
assign n1860gat = ((~n1988gat)&(~n2216gat)&(~n1862gat));
assign n2560gat = ((~n2562gat));
assign n1777gat = ((~n1694gat));
assign n1521gat = ((~n2283gat)&(~n1991gat));
assign II1996 = ((~n659gat));
assign n134gat = ((~n2875gat));
assign II4765 = ((~n2748gat));
assign n2687gat = ((~II4558));
assign II1719 = ((~n2562gat));
assign n2428gat = ((~n2433gat)&(~n2427gat));
assign n648gat = ((~n373gat)&(~n2669gat));
assign II414 = ((~n724gat));
assign II264 = ((~n2728gat));
assign II420 = ((~n1013gat));
assign n1147gat = ((~II999));
assign n1893gat = ((~n2060gat));
assign n1089gat = ((~n1067gat)&(~n1111gat));
assign n755gat = ((~II270));
assign n1162gat = ((~n698gat)&(~n1603gat));
assign n1558gat = ((~n1614gat)&(~n1553gat)&(~n1499gat));
assign n2538gat = ((~n2620gat)&(~n2625gat)&(~n2488gat));
assign n1402gat = ((~n1858gat)&(~n1393gat)&(~n1604gat));
assign II1124 = ((~n919gat));
assign n2482gat = ((~n2542gat));
assign n48gat = ((~II375));
assign n2639gat = ((~II2232));
assign n2997gat = (n2053gat)|(n2052gat)|(n1964gat);
assign II3703 = ((~n2917gat));
assign n1559gat = ((~n1614gat));
assign n158gat = ((~n160gat));
assign n2214gat = ((~n2205gat));
assign n1252gat = ((~n1199gat)&(~n2962gat));
assign n2282gat = ((~n2406gat)&(~n2215gat));
assign n804gat = ((~n808gat)&(~n809gat)&(~n810gat));
assign II4735 = ((~n2826gat));
assign n2385gat = ((~n748gat));
assign n898gat = ((~n2940gat));
assign n811gat = ((~II1344));
assign n1791gat = ((~n2013gat));
assign II3306 = ((~n1699gat));
assign n922gat = ((~n1119gat));
assign II3273 = ((~n2169gat));
assign n1577gat = ((~n1520gat)&(~n2351gat)&(~n1988gat));
assign II3461 = ((~n1956gat));
assign n876gat = ((~n1347gat));
assign II4216 = (n1427gat)|(n1595gat)|(n1677gat);
assign n292gat = ((~n415gat)&(~n356gat));
assign n2159gat = ((~n1412gat));
assign II1079 = ((~n489gat));
assign n2261gat = ((~II3000));
assign n1154gat = ((~n1598gat)&(~n2930gat)&(~n2957gat));
assign II2130 = ((~n317gat));
assign n13gat = ((~n2720gat)&(~n14gat));
assign n2665gat = ((~II1516));
assign n2184gat = ((~n3003gat));
assign n2620gat = ((~n2622gat));
assign II1028 = ((~n858gat));
assign n2137gat = ((~n2139gat));
assign n2349gat = ((~n2215gat));
assign n2707gat = ((~II3923));
assign n2384gat = ((~n43gat));
assign II1769 = ((~n1120gat));
assign n72gat = ((~n181gat));
assign n1891gat = ((~n2059gat));
assign n2580gat = ((~n2582gat)&(~n2583gat));
assign n731gat = ((~n738gat)&(~n734gat)&(~n737gat));
assign n715gat = ((~II1155));
assign n1655gat = ((~n1736gat)&(~n1662gat)&(~n1658gat));
assign n2606gat = ((~II2372));
assign n336gat = ((~II351));
assign n2530gat = ((~n2531gat));
assign n1513gat = ((~n2288gat));
assign n2579gat = (n2580gat)|(n2581gat);
assign n2945gat = (n1096gat)|(n1095gat)|(n990gat)|(n979gat);
assign n2786gat = (n3091gat)|(n3092gat);
assign n278gat = ((~II634));
assign II1230 = ((~n613gat));
assign n241gat = ((~n140gat));
assign n2409gat = (n2410gat)|(n2411gat)|(n2412gat)|(n2413gat);
assign n2935gat = (n892gat)|(n891gat);
assign II1091 = ((~n490gat));
assign n2818gat = ((~II4349));
assign II1204 = ((~n829gat));
assign n1779gat = ((~n1623gat));
assign n3034gat = ((~II3401));
assign II683 = ((~n1024gat));
assign n640gat = ((~n1213gat));
assign II642 = ((~n163gat));
assign n917gat = ((~n919gat));
assign n1043gat = ((~n1045gat));
assign n146gat = ((~n148gat));
assign n2664gat = ((~n2850gat)&(~n3018gat));
assign n1586gat = ((~n1869gat)&(~n1683gat));
assign n1439gat = ((~n1486gat));
assign n2744gat = (n2159gat)|(n2478gat);
assign n2974gat = (n1321gat)|(n1320gat);
assign n1885gat = ((~n2048gat));
assign n2966gat = (n1368gat)|(n1258gat);
assign n2828gat = ((~II4449));
assign II178 = ((~n919gat));
assign n643gat = ((~n855gat));
assign n3114gat = ((~II4684));
assign n418gat = ((~n374gat)&(~n2723gat));
assign n457gat = ((~n2884gat));
assign n445gat = ((~n2778gat)&(~n219gat));
assign n2249gat = ((~n2265gat)&(~n3006gat));
assign n2168gat = ((~II3273));
assign n122gat = ((~n125gat)&(~n128gat)&(~n129gat));
assign n1554gat = ((~n1555gat));
assign n1278gat = ((~II1923));
assign n67gat = ((~n85gat));
assign II331 = ((~n160gat));
assign n2132gat = ((~n2133gat)&(~n2131gat));
assign n982gat = ((~n873gat)&(~n1478gat));
assign n173gat = ((~II623));
assign n3134gat = ((~II4744));
assign n2255gat = ((~n2261gat)&(~n2188gat));
assign n1958gat = ((~n1963gat)&(~n1886gat));
assign n1381gat = ((~n1328gat));
assign n728gat = (n729gat)|(n730gat)|(n731gat)|(n732gat);
assign n1592gat = ((~n1529gat));
assign II729 = ((~n396gat));
assign n754gat = ((~II253));
assign n637gat = ((~n529gat));
assign n2722gat = ((~II591));
assign n347gat = ((~n353gat)&(~n351gat)&(~n350gat));
assign n1681gat = ((~II4217));
assign II4620 = ((~n1745gat));
assign n934gat = ((~n938gat)&(~n939gat)&(~n940gat));
assign n68gat = ((~n85gat)&(~n180gat));
assign n1660gat = ((~n1918gat)&(~n1986gat)&(~n2212gat));
assign II2403 = ((~n2629gat));
assign n494gat = ((~n498gat)&(~n499gat)&(~n500gat));
assign n1957gat = ((~n1886gat)&(~n1887gat));
assign n892gat = ((~n419gat)&(~n1265gat));
assign n1025gat = ((~II672));
assign n1759gat = ((~n1818gat)&(~n1935gat)&(~n2765gat));
assign n346gat = ((~n353gat)&(~n349gat)&(~n352gat));
assign n658gat = ((~II1996));
assign n2078gat = ((~n1926gat)&(~n1916gat)&(~n1994gat)&(~n1924gat));
assign II3677 = ((~n156gat));
assign II4129 = ((~n3097gat));
assign n2922gat = (n967gat)|(n792gat);
assign n2082gat = ((~n2084gat));
assign n3064gat = ((~II3914));
assign n493gat = (n494gat)|(n495gat)|(n496gat)|(n497gat);
assign II4714 = ((~n2760gat));
assign n617gat = ((~II1082));
assign n963gat = ((~n856gat)&(~n2838gat));
assign n2705gat = ((~II4601));
assign n1823gat = ((~n1821gat));
assign n2416gat = ((~II2263));
assign II4548 = ((~n2742gat));
assign n2743gat = ((~II4227));
assign II579 = ((~n2851gat));
assign n372gat = ((~n212gat));
assign n970gat = ((~n372gat)&(~n878gat));
assign n2504gat = ((~n2506gat));
assign n1012gat = ((~n1007gat)&(~n918gat));
assign II2735 = (n1788gat)|(n1884gat)|(n1633gat);
assign n46gat = ((~n53gat)&(~n49gat)&(~n52gat));
assign n422gat = ((~n2889gat));
assign n2059gat = ((~n2061gat));
assign II203 = ((~n2859gat));
assign n1435gat = ((~n1591gat)&(~n1528gat));
assign n1116gat = ((~n419gat)&(~n1266gat));
assign n1863gat = ((~n1991gat)&(~n2283gat)&(~n1989gat));
assign n568gat = ((~n572gat)&(~n573gat)&(~n574gat));
assign n234gat = ((~n155gat)&(~n233gat));
assign n1102gat = ((~n1297gat)&(~n1590gat));
assign n3032gat = ((~II3390));
assign n745gat = ((~n2716gat)&(~n2867gat));
assign n1634gat = ((~n1712gat));
assign n1935gat = ((~n1816gat)&(~n1828gat));
assign n3006gat = (n2253gat)|(n2252gat);
assign n3149gat = ((~II4789));
assign n716gat = ((~II1169));
assign n2536gat = ((~n2624gat));
assign II4536 = ((~n2750gat));
assign n121gat = ((~n125gat)&(~n126gat)&(~n127gat));
assign n2950gat = (n1001gat)|(n999gat);
assign n2778gat = ((~n2780gat));
assign n3030gat = ((~II3318));
assign n3010gat = (n2460gat)|(n2423gat);
assign n1529gat = ((~n1528gat)&(~n1523gat));
assign n2443gat = ((~n2561gat));
assign n259gat = ((~n263gat)&(~n264gat)&(~n265gat));
assign II1166 = ((~n838gat));
assign II1585 = (n2356gat)|(n2214gat)|(II1584);
assign n2993gat = (n1894gat)|(n1847gat)|(n1846gat);
assign II1837 = ((~n1282gat));
assign n2480gat = ((~n2530gat)&(~n2482gat)&(~n2486gat));
assign n159gat = ((~II331));
assign II2813 = (n1609gat)|(n1702gat)|(n1700gat)|(II2812);
assign II1453 = ((~n683gat));
assign n2494gat = ((~II2319));
assign n1591gat = ((~n2223gat));
assign II4705 = ((~n2753gat));
assign n1353gat = ((~n1419gat));
assign n530gat = ((~n2862gat)&(~n740gat));
assign n2984gat = (n1467gat)|(n1466gat);
assign n3139gat = ((~II4759));
assign II1319 = ((~n816gat));
assign II4512 = ((~n2762gat));
assign n2016gat = ((~n2019gat)&(~n1878gat));
assign n3004gat = (n2258gat)|(n2257gat)|(n2255gat);
assign n764gat = ((~n852gat)&(~n2781gat));
assign n3122gat = ((~II4708));
assign n945gat = ((~n949gat)&(~n950gat)&(~n951gat));
assign n810gat = ((~II1339));
assign II81 = ((~n2671gat));
assign n3107gat = ((~II4663));
assign n1765gat = ((~n1767gat));
assign n2726gat = ((~n2728gat));
assign n1713gat = ((~II2935));
assign n2353gat = ((~n2398gat));
assign II248 = ((~n2869gat));
assign n120gat = (n121gat)|(n122gat)|(n123gat)|(n124gat);
assign n3027gat = ((~II3309));
assign n1451gat = ((~n1382gat));
assign n1399gat = ((~n1806gat)&(~n1338gat)&(~n1584gat));
assign n1220gat = ((~II210));
assign n1693gat = ((~n2101gat));
assign n887gat = ((~n1603gat)&(~n683gat));
assign II4663 = ((~n2802gat));
assign II3179 = (n1839gat)|(n1784gat)|(II3178);
assign n3151gat = ((~II4795));
assign n2739gat = ((~n2743gat));
assign n3043gat = ((~II3494));
assign n805gat = ((~n808gat)&(~n811gat)&(~n812gat));
assign n655gat = ((~n856gat)&(~n2718gat));
assign II278 = ((~n2889gat));
assign n496gat = ((~n503gat)&(~n499gat)&(~n502gat));
assign n2811gat = ((~II4312));
assign II4081 = ((~n1807gat));
assign n1725gat = ((~n2148gat));
assign n3137gat = ((~II4753));
assign n3052gat = ((~II3610));
assign n260gat = ((~n263gat)&(~n266gat)&(~n267gat));
assign II4594 = ((~n2709gat));
assign n594gat = ((~II1407));
assign n577gat = ((~II1500));
assign n2822gat = (n77gat)|(n13gat)|(n1842gat);
assign n532gat = ((~n527gat)&(~n416gat)&(~n528gat));
assign n2717gat = ((~II1));
assign n631gat = ((~n523gat)&(~n633gat)&(~n524gat));
assign n1254gat = ((~n1123gat)&(~n1044gat));
assign n130gat = ((~II2181));
assign n1354gat = ((~n1591gat)&(~n1530gat));
assign II930 = ((~n1292gat));
assign n125gat = ((~II2056));
assign n1986gat = ((~n2439gat));
assign n1886gat = ((~n1897gat));
assign n3152gat = ((~II4798));
assign II1860 = ((~n930gat));
assign n1565gat = ((~n1735gat)&(~n1552gat));
assign n3053gat = ((~II3635));
assign n516gat = ((~n374gat)&(~n2715gat));
assign II406 = ((~n840gat));
assign n2821gat = ((~II4392));
assign n477gat = ((~n480gat)&(~n483gat)&(~n484gat));
assign II1278 = (n740gat)|(n3030gat)|(II1277);
assign n2649gat = ((~II2324));
assign II1227 = ((~n614gat));
assign n1718gat = ((~n1714gat));
assign n740gat = ((~n2667gat));
assign n481gat = ((~II443));
assign n1476gat = ((~n1858gat)&(~n1590gat));
assign n791gat = ((~n851gat)&(~n2840gat));
assign n1615gat = ((~n1624gat));
assign II746 = ((~n66gat));
assign II4144 = (n1633gat)|(n1838gat)|(n1786gat);
assign n12gat = ((~n186gat)&(~n82gat));
assign n139gat = ((~n253gat)&(~n151gat)&(~n254gat));
assign n2174gat = ((~n2176gat));
assign n765gat = ((~n2781gat)&(~n93gat));
assign n1053gat = ((~n1060gat)&(~n1056gat)&(~n1059gat));
assign n1924gat = ((~n1743gat)&(~n1923gat));
assign n2991gat = (n1654gat)|(n1653gat)|(n1644gat);
assign n1377gat = ((~n724gat)&(~n721gat));
assign II1877 = ((~n1134gat));
assign II446 = ((~n398gat));
assign n2712gat = ((~II818));
assign n2663gat = ((~n2586gat)&(~n2660gat)&(~n2307gat));
assign II2380 = ((~n2540gat));
assign n2998gat = (n2055gat)|(n1967gat);
assign II398 = ((~n841gat));
assign n1322gat = ((~n2974gat));
assign n747gat = ((~n2906gat));
assign n951gat = ((~II837));
assign n2358gat = ((~n2285gat)&(~n2356gat)&(~n2355gat));
assign II1493 = ((~n565gat));
assign n946gat = ((~n949gat)&(~n952gat)&(~n953gat));
assign II1251 = ((~n493gat));
assign n3039gat = ((~II3465));
assign n686gat = (n687gat)|(n688gat)|(n689gat)|(n690gat);
assign n2810gat = ((~II4332));
assign n1222gat = ((~II223));
assign n1999gat = ((~n2001gat));
assign n3108gat = ((~II4666));
assign n2093gat = ((~n2095gat));
assign n1418gat = ((~n1417gat));
assign II100 = ((~n2794gat));
assign II576 = ((~n3100gat));
assign n935gat = ((~n938gat)&(~n941gat)&(~n942gat));
assign II4786 = ((~n2679gat));
assign n1323gat = ((~n1007gat)&(~n401gat));
assign n1398gat = ((~n1455gat)&(~n1397gat));
assign n3110gat = ((~II4672));
assign n593gat = ((~II1402));
assign n941gat = ((~II1028));
assign n1704gat = ((~n3027gat)&(~n1706gat));
assign n1501gat = ((~n1448gat)&(~n1500gat));
assign n980gat = ((~n875gat)&(~n926gat));
assign n2558gat = ((~n2559gat));
assign n58gat = ((~n65gat)&(~n61gat)&(~n64gat));
assign n2251gat = ((~n3033gat));
assign n2329gat = ((~n1855gat)&(~n3007gat));
assign n1030gat = ((~n455gat)&(~n888gat));
assign n841gat = ((~II395));
assign n2192gat = ((~n2184gat)&(~n1855gat));
assign II4392 = ((~n2824gat));
assign n1927gat = ((~n1790gat)&(~n1635gat));
assign n1659gat = ((~n2987gat));
assign n1275gat = ((~II1843));
assign n2328gat = ((~n3008gat));
assign II1920 = ((~n1329gat));
assign n2698gat = ((~II4580));
assign n2138gat = ((~II2696));
assign II192 = ((~n3083gat));
assign n2839gat = ((~II796));
assign n2927gat = (n962gat)|(n959gat);
assign n2256gat = ((~n3032gat));
assign n1991gat = ((~n2393gat));
assign n2978gat = (n1441gat)|(n1440gat)|(n1371gat)|(n1367gat);
assign n3147gat = ((~II4783));
assign n2569gat = ((~n2573gat)&(~n2574gat)&(~n2575gat));
assign n596gat = ((~II1416));
assign II1016 = ((~n863gat));
assign n2039gat = ((~II3336));
assign n2977gat = (n1360gat)|(n1359gat)|(n1358gat)|(n1357gat);
assign n2209gat = ((~n3005gat));
assign n1784gat = ((~n1849gat));
assign n151gat = ((~II3691));
assign n2685gat = ((~n2687gat));
assign II1152 = ((~n707gat));
assign n330gat = ((~II3742));
assign II3549 = ((~n2197gat));
assign n1380gat = ((~n1114gat));
assign n801gat = ((~n672gat)&(~n670gat));
assign n54gat = ((~n167gat));
assign II606 = ((~n271gat));
assign n1858gat = ((~n1673gat));
assign II3472 = ((~n2539gat));
assign n3106gat = ((~II4660));
assign n552gat = ((~II2014));
assign II2094 = ((~n2876gat));
assign n1375gat = ((~n1006gat)&(~n706gat));
assign n1321gat = ((~n1442gat)&(~n837gat));
assign n1021gat = ((~II406));
assign n2512gat = ((~n2514gat));
assign n2590gat = ((~n2592gat));
assign II401 = ((~n721gat));
assign n2583gat = ((~n2582gat)&(~n2585gat));
assign n286gat = ((~n289gat)&(~n2723gat));
assign n2444gat = ((~n2446gat));
assign n2049gat = ((~n3001gat));
assign n2239gat = ((~n2850gat)&(~n3019gat));
assign n2906gat = (n745gat)|(n638gat);
assign n1582gat = ((~n2283gat)&(~n1991gat)&(~n2212gat));
assign n387gat = ((~II3736));
assign n1230gat = ((~n1233gat)&(~n1236gat)&(~n1237gat));
assign n37gat = ((~n151gat)&(~n154gat));
assign II793 = ((~n1067gat));
assign II3401 = ((~n2192gat));
assign n409gat = ((~n406gat)&(~n407gat));
assign II1947 = ((~n1197gat));
assign n1469gat = ((~n1858gat)&(~n1608gat));
assign n1180gat = ((~n2948gat));
assign n1146gat = ((~n1148gat));
assign n2181gat = ((~II3016));
assign II3163 = ((~n1508gat));
assign n1702gat = ((~n3024gat)&(~n1615gat));
assign n2943gat = (n1012gat)|(n905gat);
assign n381gat = ((~n2893gat));
assign n1649gat = ((~n1560gat)&(~n1659gat)&(~n1730gat));
assign n2462gat = ((~n2464gat));
assign n559gat = ((~n561gat));
assign n1013gat = (n1014gat)|(n1015gat)|(n1016gat)|(n1017gat);
assign n1190gat = ((~II1769));
assign n129gat = ((~II2177));
assign n1600gat = ((~n1685gat)&(~n1427gat));
assign n2617gat = ((~n2616gat)&(~n2619gat));
assign n225gat = ((~n231gat)&(~n229gat)&(~n228gat));
assign n358gat = ((~n532gat));
assign II646 = ((~n277gat));
assign n2330gat = ((~n2437gat)&(~n1961gat));
assign II4492 = ((~n2681gat));
assign n698gat = ((~II1464));
assign n1761gat = ((~n2985gat)&(~n1602gat)&(~n1681gat));
assign n1531gat = ((~n1507gat)&(~n1477gat));
assign n1218gat = ((~II196));
assign n2289gat = ((~II1724));
assign II1118 = ((~n846gat));
assign n2624gat = ((~n2626gat));
assign n2281gat = ((~n3009gat));
assign n1204gat = ((~n1211gat)&(~n1207gat)&(~n1210gat));
assign n2790gat = ((~II65));
assign n2437gat = ((~n2195gat));
assign II256 = ((~n2725gat));
assign n348gat = ((~II712));
assign n719gat = ((~II1183));
assign II2260 = ((~n2203gat));
assign n525gat = ((~n526gat)&(~n531gat)&(~n530gat));
assign II1733 = (n2286gat)|(n2428gat)|(n2289gat);
assign n2970gat = (n1383gat)|(n1327gat);
assign n2550gat = ((~II2403));
assign II4138 = ((~n2766gat));
assign n999gat = ((~n419gat)&(~n1171gat));
assign n1663gat = ((~n1986gat)&(~n1918gat));
assign n2827gat = ((~II3962));
assign n2882gat = (n242gat)|(n240gat);
assign n1735gat = ((~n1861gat));
assign n790gat = ((~n856gat)&(~n2840gat));
assign II468 = ((~n42gat));
assign n133gat = ((~n2876gat));
assign n1262gat = ((~n837gat)&(~n1006gat));
assign n2854gat = ((~n2856gat));
assign n2108gat = ((~n2110gat));
assign n1452gat = ((~n2049gat));
assign II4236 = ((~n2808gat));
assign n1078gat = ((~n1080gat));
assign II913 = ((~n673gat));
assign n1728gat = ((~n1568gat)&(~n1736gat)&(~n1658gat));
assign n15gat = ((~n637gat)&(~n17gat)&(~n293gat));
assign n458gat = ((~n2902gat));
assign II3945 = ((~n1350gat));
assign II3457 = ((~n2556gat));
assign n1194gat = ((~II1800));
assign n242gat = ((~n254gat)&(~n241gat));
assign II3999 = (n2167gat)|(n2031gat)|(n2174gat);
assign n1422gat = ((~n2011gat)&(~n2162gat));
assign n2708gat = (n848gat)|(n2047gat);
assign II3293 = ((~n1691gat));
assign n1391gat = ((~n1513gat)&(~n2442gat));
assign n2248gat = ((~n3006gat));
assign n3016gat = (n2596gat)|(n2595gat);
assign n1371gat = ((~n1370gat)&(~n1369gat));
assign n2706gat = ((~II4594));
assign II314 = ((~n270gat));
assign II11 = ((~n3093gat));
assign n1964gat = ((~n2392gat)&(~n2439gat));
assign n1650gat = ((~n1727gat)&(~n1659gat)&(~n1640gat));
assign n2801gat = ((~II4633));
assign II687 = ((~n917gat));
assign n2474gat = ((~n2476gat));
assign n2975gat = (n1443gat)|(n1325gat);
assign n1296gat = ((~n673gat));
assign II1422 = ((~n586gat));
assign n998gat = ((~n725gat)&(~n741gat));
assign n1915gat = ((~n1859gat)&(~n1919gat));
assign n714gat = ((~II1141));
assign n2879gat = (n145gat)|(n143gat);
assign n288gat = ((~n289gat)&(~n2726gat));
assign II2148 = ((~n313gat));
assign n967gat = ((~n373gat)&(~n2672gat));
assign II3483 = ((~n2436gat));
assign n1276gat = ((~II1915));
assign II4696 = ((~n2738gat));
assign n2154gat = ((~II1698));
assign n2857gat = ((~n2858gat));
assign n132gat = ((~n560gat)&(~n364gat));
assign n1628gat = ((~n1621gat));
assign n1074gat = ((~n2775gat)&(~n110gat));
assign n3007gat = (n2250gat)|(n2249gat);
assign n2742gat = (n1005gat)|(n2384gat);
assign n2915gat = (n965gat)|(n960gat)|(n661gat);
assign n1224gat = ((~n1226gat));
assign n1623gat = ((~n1379gat)&(~n1446gat));
assign n2859gat = ((~n2861gat));
assign n2555gat = ((~II2433));
assign n2755gat = ((~n2758gat));
assign II3736 = ((~n388gat));
assign n2710gat = (n69gat)|(n1885gat);
assign n1745gat = ((~n1869gat)&(~n1757gat));
assign II963 = ((~n3079gat));
assign n368gat = ((~n1725gat));
assign n1425gat = ((~n1421gat));
assign n21gat = ((~n15gat));
assign n85gat = ((~n17gat)&(~n294gat)&(~n637gat));
assign n140gat = ((~n151gat)&(~n253gat)&(~n155gat));
assign n2721gat = ((~II594));
assign n2178gat = ((~II2953));
assign n901gat = ((~n419gat)&(~n1259gat));
assign n2628gat = ((~n2630gat));
assign n889gat = ((~n1111gat)&(~n1079gat));
assign n3026gat = ((~II3306));
assign n252gat = ((~n2877gat));
assign n2759gat = ((~II4518));
assign n1195gat = ((~n1197gat));
assign n93gat = ((~n197gat)&(~n22gat));
assign n2995gat = (n1962gat)|(n1955gat);
assign n724gat = ((~n846gat));
assign II375 = ((~n41gat));
assign n718gat = ((~II1178));
assign n339gat = ((~n341gat));
assign n237gat = ((~n140gat)&(~n147gat));
assign n2806gat = ((~II4620));
assign n940gat = ((~II1023));
assign n1847gat = ((~n1958gat)&(~n1845gat));
assign II3660 = ((~n2636gat));
assign n2911gat = (n761gat)|(n651gat);
assign n2757gat = (n1030gat)|(n2245gat);
assign n3127gat = ((~II4723));
assign n2004gat = ((~n1929gat));
assign n1267gat = ((~n613gat)&(~n1006gat));
assign n2508gat = ((~n2510gat));
assign II925 = ((~n1296gat));
assign n413gat = ((~n411gat));
assign n254gat = ((~n256gat));
assign n1743gat = ((~n1713gat));
assign n758gat = ((~II282));
assign n2594gat = ((~n3017gat)&(~n2520gat)&(~n2597gat));
assign n1739gat = ((~II2915));
assign n317gat = ((~II2127));
assign n483gat = ((~II453));
assign n1698gat = ((~n1934gat));
assign II2414 = ((~n2634gat));
assign n2461gat = ((~n120gat)&(~n2666gat));
assign n504gat = (n505gat)|(n506gat)|(n507gat)|(n508gat);
assign n1360gat = ((~n1164gat)&(~n1356gat));
assign n595gat = ((~II1411));
assign II1371 = ((~n824gat));
assign n3141gat = ((~II4765));
assign n224gat = ((~n231gat)&(~n227gat)&(~n230gat));
assign n768gat = ((~n373gat)&(~n2731gat));
assign n1962gat = ((~n1963gat)&(~n1893gat));
assign n2127gat = ((~n2389gat));
assign n836gat = ((~n838gat));
assign n569gat = ((~n572gat)&(~n575gat)&(~n576gat));
assign n527gat = ((~n356gat));
assign II4729 = ((~n2803gat));
assign n2288gat = ((~II4024));
assign n985gat = ((~n775gat));
assign II2251 = ((~n2207gat));
assign n2264gat = ((~n2266gat));
assign n179gat = ((~n287gat));
assign n784gat = ((~II1999));
assign II4601 = ((~n2708gat));
assign II2127 = ((~n318gat));
assign n1890gat = ((~n2328gat));
assign n299gat = ((~n2268gat)&(~n2338gat));
assign II47 = ((~n3069gat));
assign n2586gat = ((~n2588gat));
assign n2764gat = (n1029gat)|(n2237gat);
assign II1385 = ((~n820gat));
assign n2648gat = ((~n2650gat)&(~n2652gat));
assign n711gat = ((~n714gat)&(~n717gat)&(~n718gat));
assign n832gat = ((~n834gat));
assign II509 = ((~n3099gat));
assign n725gat = ((~II171));
assign n624gat = ((~n919gat));
assign n2900gat = (n869gat)|(n453gat)|(n448gat);
assign n1178gat = ((~n420gat)&(~n1179gat));
assign II217 = ((~n2860gat));
assign n1570gat = ((~n1736gat)&(~n1658gat)&(~n1670gat));
assign n2498gat = ((~n2199gat)&(~n2328gat));
assign n2901gat = (n558gat)|(n555gat)|(n450gat);
assign n1572gat = ((~n1576gat));
assign n2656gat = ((~n2658gat));
assign n1066gat = ((~n1068gat));
assign n1733gat = ((~n1673gat)&(~n1572gat));
assign II4558 = ((~n1286gat));
assign n1057gat = ((~II1002));
assign n2411gat = ((~n2414gat)&(~n2417gat)&(~n2418gat));
assign n749gat = ((~n753gat)&(~n754gat)&(~n755gat));
assign n3008gat = (n2332gat)|(n2259gat);
assign n2666gat = ((~n1704gat));
assign n243gat = ((~n1702gat));
assign n2051gat = ((~n2056gat));
assign n1716gat = ((~II2736));
assign n1256gat = ((~n392gat)&(~n702gat));
assign n2647gat = ((~n2649gat)&(~n2650gat));
assign n3021gat = ((~II3290));
assign n1297gat = ((~II913));
assign n1971gat = ((~n1896gat)&(~n1973gat));
assign n360gat = ((~n2859gat)&(~n2727gat));
assign II609 = ((~n282gat));
assign n1499gat = ((~n396gat)&(~n401gat));
assign n1438gat = ((~n1591gat)&(~n1480gat));
assign II3429 = ((~n2266gat));
assign n1472gat = ((~n1476gat)&(~n1471gat)&(~n1469gat));
assign n1440gat = ((~n1322gat)&(~n1439gat));
assign n1756gat = ((~n2512gat)&(~n1769gat)&(~n1773gat));
assign n827gat = ((~n204gat));
assign n2551gat = ((~II2417));
assign n1009gat = ((~n1255gat)&(~n2943gat));
assign n904gat = ((~n1006gat)&(~n490gat));
assign II1353 = ((~n678gat));
assign II18 = ((~n3072gat));
assign II2349 = ((~n2270gat));
assign II1450 = ((~n684gat));
assign n2442gat = ((~n2483gat));
assign n3109gat = ((~II4669));
assign n697gat = ((~n699gat));
assign n1916gat = ((~n1917gat)&(~n1859gat));
assign n1079gat = ((~II977));
assign II4771 = ((~n2797gat));
assign II4708 = ((~n2754gat));
assign II4587 = ((~n2701gat));
assign II210 = ((~n2862gat));
assign n1797gat = ((~n1801gat));
assign n2800gat = (n2158gat)|(n2186gat);
assign n2398gat = ((~II1538));
assign n1370gat = ((~n1426gat));
assign II2926 = (n1884gat)|(n1787gat)|(II2925);
assign n45gat = ((~n48gat)&(~n51gat)&(~n52gat));
assign n1209gat = ((~II1899));
assign II1752 = ((~n1034gat));
assign n1561gat = ((~n1571gat));
assign n859gat = ((~n861gat));
assign II658 = ((~n54gat));
assign n2415gat = ((~II2257));
assign n3148gat = ((~II4786));
assign n2187gat = ((~n3004gat));
assign n16gat = ((~n564gat));
assign n1668gat = ((~n1734gat));
assign n416gat = ((~n415gat));
assign II2978 = ((~n2190gat));
assign n1708gat = ((~n2338gat));
assign II3935 = ((~n2704gat));
assign II4741 = ((~n2821gat));
assign n1594gat = ((~n1596gat));
assign n2898gat = (n447gat)|(n445gat);
assign n2351gat = ((~n2405gat));
assign II692 = ((~n844gat));
assign n1648gat = ((~n1729gat));
assign n2884gat = (n246gat)|(n245gat);
assign n2478gat = ((~n2579gat));
assign n1233gat = ((~II880));
assign n174gat = ((~II637));
assign n851gat = ((~n853gat));
assign n505gat = ((~n509gat)&(~n510gat)&(~n511gat));
assign II4711 = ((~n2759gat));
assign n3128gat = ((~II4726));
assign n2005gat = ((~n2002gat)&(~n2857gat));
assign n1455gat = ((~II4105));
assign n2153gat = ((~n2155gat));
assign n2013gat = ((~II4000));
assign n482gat = ((~II449));
assign n1355gat = ((~n1422gat));
assign II1183 = ((~n832gat));
assign n515gat = ((~n709gat));
assign n2876gat = (n874gat)|(n132gat);
assign n1058gat = ((~II1007));
assign n1292gat = ((~n1294gat));
assign n1560gat = ((~n1557gat));
assign n2842gat = ((~n2843gat));
assign II2425 = ((~n2632gat));
assign n2356gat = ((~n2560gat));
assign n1639gat = ((~n1499gat)&(~n1559gat)&(~n1553gat));
assign n2608gat = ((~II2380));
assign n1181gat = ((~n455gat)&(~n1179gat));
assign n1033gat = ((~n1035gat));
assign II4369 = ((~n2937gat));
assign n1453gat = ((~n2187gat));
assign II3016 = ((~n2182gat));
assign n401gat = ((~II76));
assign n2700gat = ((~II3935));
assign n1552gat = ((~n1550gat));
assign n612gat = ((~n614gat));
assign II449 = ((~n393gat));
assign n2802gat = ((~II4623));
assign II4233 = ((~n1721gat));
assign n391gat = ((~n252gat)&(~n468gat));
assign II1698 = ((~n2155gat));
assign n556gat = ((~n2672gat)&(~n852gat));
assign n654gat = ((~n851gat)&(~n2844gat));
assign n873gat = ((~n316gat));
assign n186gat = ((~n189gat)&(~n287gat)&(~n288gat));
assign II2372 = ((~n2612gat));
assign n1300gat = ((~n2963gat));
assign n2333gat = ((~n2438gat));
assign n1261gat = ((~n833gat)&(~n1006gat));
assign n1213gat = (n1214gat)|(n1215gat)|(n1216gat)|(n1217gat);
assign n1626gat = ((~n1627gat)&(~n3022gat));
assign n2346gat = ((~II2837));
assign n2636gat = ((~n2637gat));
assign n734gat = ((~II1204));
assign n227gat = ((~II2130));
assign n1184gat = (n1185gat)|(n1186gat)|(n1187gat)|(n1188gat);
assign II354 = ((~n336gat));
assign n2056gat = ((~n2998gat));
assign n575gat = ((~II1493));
assign n2081gat = ((~n2218gat));
assign n1229gat = ((~n1233gat)&(~n1234gat)&(~n1235gat));
assign n1667gat = ((~n1991gat)&(~n1986gat));
assign n636gat = ((~n414gat)&(~n633gat)&(~n639gat));
assign n1407gat = ((~n1393gat)&(~n1409gat)&(~n1677gat));
assign n1517gat = ((~n1578gat));
assign n2716gat = ((~II240));
assign n2540gat = ((~n2488gat));
assign II3436 = ((~n2492gat));
assign n2940gat = (n1152gat)|(n1092gat)|(n997gat)|(n993gat);
assign n1098gat = ((~n336gat)&(~n741gat));
assign n2123gat = ((~n2125gat));
assign n858gat = ((~n1228gat));
assign n2914gat = (n768gat)|(n655gat);
assign II27 = ((~n3095gat));
assign n3058gat = ((~II3765));
assign n1449gat = ((~n1494gat));
assign n176gat = ((~II646));
assign n1516gat = ((~n1551gat)&(~n1517gat));
assign n869gat = ((~n219gat)&(~n2792gat));
assign n2816gat = ((~II4352));
assign II661 = ((~n845gat));
assign n1478gat = ((~n1481gat));
assign n1413gat = ((~n1869gat)&(~n672gat)&(~n2591gat));
assign II2439 = ((~n2545gat));
assign n1620gat = ((~n1448gat)&(~n1446gat));
assign n531gat = ((~n740gat)&(~n2854gat));
assign n672gat = ((~II44));
assign n3046gat = ((~II3513));
assign II2275 = ((~n2205gat));
assign n2196gat = ((~n2199gat)&(~n2146gat));
assign n1106gat = ((~n2949gat));
assign n2745gat = ((~II4542));
assign n261gat = ((~n268gat)&(~n264gat)&(~n267gat));
assign n2831gat = ((~II771));
assign II3587 = ((~n2125gat));
assign n2999gat = (n1972gat)|(n1971gat);
assign n1329gat = ((~n2970gat));
assign n781gat = ((~n784gat)&(~n787gat)&(~n788gat));
assign n2856gat = ((~II192));
assign n2134gat = ((~II2989));
assign n2532gat = ((~n2625gat));
assign n1076gat = ((~n93gat)&(~n2775gat));
assign n1034gat = ((~II1749));
assign n1459gat = ((~n1595gat)&(~n1454gat));
assign n2393gat = ((~II2847));
assign n57gat = ((~n60gat)&(~n63gat)&(~n64gat));
assign n2285gat = ((~n2397gat));
assign n124gat = ((~n130gat)&(~n128gat)&(~n127gat));
assign n644gat = ((~n855gat));
assign n937gat = ((~n943gat)&(~n941gat)&(~n940gat));
assign n579gat = ((~II1336));
assign n1796gat = ((~n1858gat)&(~n1635gat));
assign II753 = ((~n167gat));
assign n3041gat = ((~II3483));
assign II2420 = ((~n2542gat));
assign n1245gat = ((~n1590gat)&(~n860gat));
assign II1749 = ((~n1035gat));
assign n2723gat = ((~n2725gat));
assign n2838gat = ((~n2839gat));
assign n1437gat = ((~n1438gat));
assign n1086gat = ((~n1870gat));
assign n440gat = ((~n856gat)&(~n2842gat));
assign n1406gat = ((~n1428gat)&(~n1387gat));
assign n1396gat = ((~n1401gat));
assign II3287 = ((~n1691gat));
assign II3817 = ((~n2916gat));
assign n3048gat = ((~II3530));
assign II334 = ((~n159gat));
assign n411gat = ((~n374gat)&(~n2726gat));
assign n730gat = ((~n733gat)&(~n736gat)&(~n737gat));
assign n2561gat = ((~II1719));
assign n378gat = ((~n375gat)&(~n235gat));
assign II3558 = ((~n2196gat));
assign n207gat = ((~n2337gat)&(~n2269gat));
assign n2619gat = ((~II2439));
assign II2228 = ((~n2561gat));
assign n1470gat = ((~n1472gat)&(~n1747gat));
assign n1071gat = ((~II1783));
assign II2736 = (n1785gat)|(n1784gat)|(II2735);
assign n1691gat = ((~n2452gat));
assign II2889 = (n1784gat)|(n1633gat)|(n1884gat);
assign n557gat = ((~n2669gat)&(~n852gat));
assign n1481gat = ((~n2081gat)&(~n2011gat));
assign n412gat = ((~n522gat));
assign n1575gat = ((~n1918gat)&(~n2283gat));
assign n2784gat = ((~n2786gat));
assign n1238gat = ((~II930));
assign n2920gat = (n867gat)|(n771gat);
assign n2568gat = (n2569gat)|(n2570gat)|(n2571gat)|(n2572gat);
assign n1397gat = ((~n1519gat)&(~n1401gat));
assign II1703 = ((~n2626gat));
assign n2524gat = ((~n2526gat));
assign n2566gat = ((~n2643gat)&(~n2564gat));
assign II3610 = ((~n1882gat));
assign n450gat = ((~n851gat)&(~n2846gat));
assign n2533gat = ((~n2534gat));
assign n2542gat = ((~II1708));
assign n163gat = ((~n160gat));
assign n2015gat = ((~n2039gat)&(~n1774gat)&(~n1315gat));
assign II2684 = ((~n2061gat));
assign n833gat = ((~II1138));
assign II1127 = ((~n625gat));
assign n2559gat = ((~n2999gat)&(~n2437gat));
assign n390gat = ((~n469gat)&(~n2877gat));
assign II1915 = ((~n1268gat));
assign n763gat = ((~n2672gat)&(~n93gat));
assign II1766 = ((~n1121gat));
assign n2567gat = ((~n2493gat)&(~n2388gat));
assign n914gat = ((~II683));
assign II2235 = ((~n2639gat));
assign II3876 = ((~n2926gat));
assign n641gat = ((~n855gat));
assign II4157 = ((~n1525gat));
assign n442gat = ((~n2844gat)&(~n856gat));
assign n2864gat = ((~II206));
assign n872gat = ((~n375gat)&(~n800gat));
assign n1661gat = ((~n1660gat));
assign n2258gat = ((~n2260gat)&(~n2189gat));
assign II4738 = ((~n2820gat));
assign n717gat = ((~II1174));
assign II384 = ((~n2674gat));
assign n171gat = ((~n177gat)&(~n175gat)&(~n174gat));
assign n895gat = ((~n420gat)&(~n898gat));
assign n942gat = ((~II1031));
assign n706gat = ((~II1152));
assign n2825gat = ((~II4452));
assign n497gat = ((~n503gat)&(~n501gat)&(~n500gat));
assign n1092gat = ((~n1147gat)&(~n1111gat));
assign II1617 = ((~n2622gat));
assign n296gat = ((~n421gat));
assign II885 = ((~n3082gat));
assign n2711gat = ((~n2712gat));
assign II2248 = ((~n2568gat));
assign II1103 = ((~n620gat));
assign n797gat = ((~n110gat)&(~n2734gat));
assign n564gat = ((~n3029gat)&(~n2863gat)&(~n2855gat)&(~n374gat));
assign n1206gat = ((~II1860));
assign n60gat = ((~II658));
assign n1349gat = ((~n1479gat)&(~n2081gat));
assign n1327gat = ((~n1281gat)&(~n1224gat));
assign n2979gat = (n1373gat)|(n1372gat);
assign n2817gat = ((~II4369));
assign II1800 = ((~n1033gat));
assign n1730gat = ((~n1731gat));
assign n1384gat = ((~n2184gat));
assign n1383gat = ((~n1280gat)&(~n1225gat));
assign n787gat = ((~II2040));
assign n2364gat = ((~n2353gat)&(~n2284gat)&(~n2356gat));
assign n383gat = ((~II3831));
assign n1665gat = ((~n1666gat));
assign n155gat = ((~II3677));
assign II4608 = ((~n2799gat));
assign n2994gat = (n1954gat)|(n1888gat);
assign n1022gat = ((~II409));
assign n1621gat = ((~n1319gat)&(~n1380gat));
assign n2761gat = (n1031gat)|(n2325gat);
assign II1088 = ((~n398gat));
assign n1005gat = ((~n894gat)&(~n455gat));
assign n845gat = ((~II111));
assign II4185 = ((~n1596gat));
assign II1178 = ((~n836gat));
assign n844gat = ((~n846gat));
assign n2306gat = ((~n2356gat)&(~n2284gat)&(~n2285gat));
assign n567gat = (n568gat)|(n569gat)|(n570gat)|(n571gat);
assign n2611gat = ((~II2394));
assign n3133gat = ((~II4741));
assign n995gat = ((~n823gat)&(~n1112gat));
assign n1003gat = ((~n420gat)&(~n879gat));
assign n2958gat = (n1246gat)|(n1161gat);
assign II4693 = ((~n2737gat));
assign II3914 = ((~n2923gat));
assign n2690gat = ((~II4566));
assign II3318 = ((~n1869gat));
assign n2963gat = (n1291gat)|(n1245gat);
assign n250gat = ((~n329gat)&(~n387gat)&(~n334gat));
assign n2973gat = (n1352gat)|(n1351gat)|(n1303gat)|(n1302gat);
assign n1515gat = ((~n1521gat));
assign n973gat = ((~n372gat)&(~n333gat));
assign n1633gat = ((~n2137gat));
assign n1731gat = ((~n1658gat)&(~n1515gat)&(~n1797gat));
assign n1255gat = ((~n1123gat)&(~n1225gat));
assign n1176gat = ((~n829gat)&(~n1006gat));
assign n650gat = ((~n852gat)&(~n2789gat));
assign II2354 = ((~n2880gat));
assign n500gat = ((~II1091));
assign n1237gat = ((~II925));
assign n495gat = ((~n498gat)&(~n501gat)&(~n502gat));
assign n1640gat = ((~n1639gat));
assign n2929gat = (n974gat)|(n973gat)|(n870gat);
assign II955 = ((~n865gat));
assign n1692gat = ((~n1879gat)&(~n1762gat));
assign n349gat = ((~II715));
assign II1550 = ((~n2343gat));
assign n2928gat = (n963gat)|(n868gat);
assign n1711gat = ((~n2990gat));
assign n2961gat = (n1375gat)|(n1324gat);
assign II3962 = ((~n2830gat));
assign II709 = ((~n341gat));
assign II4615 = ((~n2798gat));
assign n2290gat = ((~n2202gat));
assign n2638gat = ((~n2640gat));
assign n1088gat = ((~n1085gat)&(~n926gat));
assign n2000gat = ((~n1412gat));
assign n2001gat = ((~n1412gat));
assign II818 = ((~n3075gat));
assign n2954gat = (n1250gat)|(n1103gat);
assign n657gat = ((~n659gat));
assign n1347gat = ((~n2081gat)&(~n1410gat));
assign II270 = ((~n422gat));
assign n1171gat = ((~n2960gat)&(~n1243gat));
assign n2614gat = ((~n2616gat)&(~n2617gat));
assign n77gat = ((~n76gat)&(~n2784gat));
assign n1544gat = ((~n1625gat));
assign n1793gat = ((~n1792gat)&(~n1735gat));
assign n1510gat = ((~n1584gat)&(~n1460gat));
assign n2307gat = ((~n2309gat));
assign II1734 = (n1604gat)|(n2214gat)|(II1733);
assign n1622gat = ((~n1380gat)&(~n1446gat));
assign II214 = ((~n2861gat));
assign II2162 = ((~n320gat));
assign n359gat = ((~n290gat)&(~n358gat));
assign n2581gat = ((~n2583gat)&(~n2585gat));
assign n2968gat = (n1326gat)|(n1261gat);
assign n3031gat = ((~II3387));
assign n478gat = ((~n485gat)&(~n481gat)&(~n484gat));
assign II2056 = ((~n35gat));
assign n87gat = ((~n743gat)&(~n17gat)&(~n293gat));
assign n2396gat = ((~n2199gat)&(~n2209gat));
assign n1272gat = ((~n1279gat)&(~n1275gat)&(~n1278gat));
assign n462gat = ((~II3777));
assign n936gat = ((~n943gat)&(~n939gat)&(~n942gat));
assign n2701gat = (n921gat)|(n1890gat);
assign n2912gat = (n762gat)|(n652gat);
assign n320gat = ((~n322gat));
assign n796gat = ((~n2731gat)&(~n110gat));
assign n2851gat = ((~II576));
assign n1156gat = ((~n985gat)&(~n1307gat));
assign n3033gat = ((~II3394));
assign n854gat = ((~n2148gat)&(~n374gat));
assign n2412gat = ((~n2419gat)&(~n2415gat)&(~n2418gat));
assign n837gat = ((~II1166));
assign II3646 = ((~n2644gat));
assign II3390 = ((~n2261gat));
assign II297 = ((~n3065gat));
assign n2341gat = ((~n2343gat));
assign n335gat = ((~n337gat));
assign n1569gat = ((~n1570gat));
assign n2250gat = ((~n2248gat)&(~n2264gat));
assign n3051gat = ((~II3558));
assign n1044gat = ((~II1891));
assign II1981 = ((~n667gat));
assign n1504gat = ((~n1450gat)&(~n1498gat));
assign n2047gat = ((~n2209gat));
assign n88gat = ((~n84gat));
assign n371gat = ((~n1725gat));
assign n882gat = ((~II1399));
assign II2925 = (n1784gat)|(n1785gat)|(n1633gat);
assign n3038gat = ((~II3461));
assign n2971gat = (n1287gat)|(n1285gat);
assign II3491 = ((~n2387gat));
assign n908gat = ((~n911gat)&(~n914gat)&(~n915gat));
assign n1652gat = ((~n1657gat));
assign n1747gat = ((~II4055));
assign n1258gat = ((~n274gat)&(~n1444gat));
assign n1959gat = ((~n1956gat)&(~n1963gat));
assign n2245gat = ((~n504gat));
assign n316gat = ((~n318gat));
assign n3022gat = ((~II3293));
assign n55gat = (n56gat)|(n57gat)|(n58gat)|(n59gat);
assign n2152gat = ((~n2346gat));
assign n902gat = ((~n1009gat)&(~n419gat));
assign n1196gat = ((~II1947));
assign n2837gat = ((~II941));
assign n1657gat = ((~n1662gat)&(~n1797gat)&(~n1658gat));
assign n1284gat = ((~n1269gat));
assign n3061gat = ((~II3841));
assign n994gat = ((~n1112gat)&(~n882gat));
assign II1011 = ((~n1146gat));
assign II1903 = ((~n1043gat));
assign II4482 = ((~n2127gat));
assign n2669gat = ((~n2671gat));
assign n528gat = ((~n521gat));
assign II223 = ((~n2863gat));
assign n1896gat = ((~n2995gat)&(~n1895gat));
assign n489gat = ((~n398gat));
assign II2376 = ((~n2532gat));
assign n566gat = ((~n364gat));
assign n1056gat = ((~II980));
assign n560gat = ((~II2088));
assign n2902gat = (n460gat)|(n459gat);
assign n1286gat = ((~n1269gat));
assign II4312 = ((~n2814gat));
assign n41gat = ((~n258gat));
assign n1503gat = ((~n1501gat));
assign n2260gat = ((~n2262gat));
assign n2090gat = ((~II2885));
assign II2843 = ((~n2403gat));
assign II623 = ((~n164gat));
assign n126gat = ((~II2094));
assign n870gat = ((~n2669gat)&(~n219gat));
assign n1645gat = ((~n1499gat));
assign n1758gat = ((~n1311gat)&(~n1773gat));
assign II4542 = ((~n2749gat));
assign II4675 = ((~n2706gat));
assign n3024gat = ((~II3300));
assign II275 = ((~n747gat));
assign II4055 = ((~n1748gat));
assign n823gat = ((~II1371));
assign n2549gat = ((~n2555gat)&(~n2553gat)&(~n2552gat));
assign II1277 = (n2860gat)|(n2855gat)|(n2863gat);
assign II1302 = ((~n680gat));
assign n1339gat = ((~II4108));
assign n1828gat = ((~II572));
assign n2680gat = ((~II3941));
assign n1616gat = ((~n918gat)&(~n396gat));
assign n511gat = ((~II1243));
assign n592gat = ((~II1388));
assign n265gat = ((~II354));
assign II2935 = (n1785gat)|(n1884gat)|(II2934);
assign n350gat = ((~II721));
assign II4780 = ((~n2691gat));
assign n529gat = ((~n2724gat)&(~n2715gat));
assign n2782gat = ((~II50));
assign n3005gat = (n2211gat)|(n2210gat);
assign n1832gat = ((~n1834gat));
assign n780gat = ((~n784gat)&(~n785gat)&(~n786gat));
assign II1655 = ((~n2102gat));
assign n1427gat = ((~n1608gat));
assign n639gat = ((~n523gat));
assign II2319 = ((~n2495gat));
assign II4014 = ((~n2744gat));
assign n374gat = ((~n2767gat));
assign II461 = ((~n339gat));
assign n1133gat = ((~n1135gat));
assign n1926gat = ((~n1925gat)&(~n1635gat));
assign n326gat = ((~II3808));
assign n1093gat = ((~n1111gat)&(~n864gat));
assign n66gat = ((~n906gat));
assign n1188gat = ((~n1194gat)&(~n1192gat)&(~n1191gat));
assign II2088 = ((~n561gat));
assign n110gat = ((~n182gat)&(~n89gat));
assign n1644gat = ((~n1643gat)&(~n1648gat)&(~n1659gat));
assign n695gat = ((~II1476));
assign n2438gat = ((~n2440gat));
assign n2188gat = ((~n2190gat));
assign n972gat = ((~n372gat)&(~n458gat));
assign II3309 = ((~n1699gat));
assign II4566 = ((~n2694gat));
assign n1177gat = ((~n1180gat)&(~n420gat));
assign II916 = ((~n1297gat));
assign n1304gat = ((~n1590gat)&(~n1067gat));
assign n480gat = ((~II440));
assign n1601gat = ((~n120gat));
assign II4795 = ((~n2700gat));
assign n2643gat = ((~II3646));
assign n3113gat = ((~II4681));
assign n1307gat = ((~n1308gat));
assign n2799gat = (n849gat)|(n2050gat);
assign n894gat = ((~n2932gat));
assign n475gat = (n476gat)|(n477gat)|(n478gat)|(n479gat);
assign n663gat = ((~n1725gat));
assign n1862gat = ((~n1863gat));
assign II2169 = ((~n34gat));
assign n900gat = ((~n419gat)&(~n1008gat));
assign n2807gat = ((~II4475));
assign n1319gat = ((~n1256gat));
assign II3168 = ((~n1394gat));
assign n822gat = ((~n824gat));
assign n971gat = ((~n111gat)&(~n2840gat));
assign n238gat = ((~n147gat)&(~n254gat));
assign n1240gat = ((~II899));
assign II3000 = ((~n2262gat));
assign n693gat = ((~II1467));
assign n621gat = ((~II1118));
assign II2785 = ((~n2407gat));
assign n245gat = ((~n386gat)&(~n334gat));
assign II1305 = ((~n679gat));
assign n417gat = ((~n418gat));
assign n248gat = ((~n330gat)&(~n1490gat));
assign n613gat = ((~II1227));
assign n1658gat = ((~n2216gat));
assign II718 = ((~n398gat));
assign n2031gat = ((~n2033gat));
assign n682gat = ((~n684gat));
assign n2980gat = (n1470gat)|(n1400gat)|(n1399gat)|(n1398gat);
assign n2715gat = ((~n2717gat));
assign II14 = ((~n2768gat));
assign n2796gat = ((~II4608));
assign n918gat = ((~II92));
assign n1654gat = ((~n1671gat)&(~n1659gat));
assign n2813gat = ((~II4329));
assign n628gat = ((~n631gat));
assign n1273gat = ((~n1279gat)&(~n1277gat)&(~n1276gat));
assign n912gat = ((~II675));
assign n2888gat = (n663gat)|(n649gat)|(n449gat);
assign II1141 = ((~n833gat));
assign n1243gat = ((~n1281gat)&(~n1123gat));
assign n2331gat = ((~n2393gat)&(~n2401gat));
assign n2466gat = ((~n2468gat));
assign II3777 = ((~n463gat));
assign n2012gat = ((~n2016gat));
assign n14gat = ((~n186gat));
assign II1500 = ((~n803gat));
assign n1518gat = ((~n1694gat));
assign n268gat = ((~II368));
assign II2281 = ((~n2409gat));
assign n1895gat = ((~n1845gat)&(~n1891gat)&(~n1968gat));
assign n642gat = ((~n855gat));
assign n1817gat = ((~n1819gat)&(~n1823gat));
assign II2771 = ((~n2440gat));
assign n977gat = ((~n670gat)&(~n671gat));
assign n665gat = ((~n667gat));
assign n1085gat = ((~n551gat));
assign II4762 = ((~n2747gat));
assign n1631gat = ((~n1848gat));
assign n61gat = ((~II698));
assign n1443gat = ((~n1442gat)&(~n706gat));
assign II196 = ((~n2854gat));
assign n2058gat = ((~n2997gat));
assign n671gat = ((~n673gat));
assign n1020gat = ((~II401));
assign n1454gat = ((~n1469gat));
assign n518gat = ((~n520gat)&(~n519gat));
assign n404gat = ((~n493gat));
assign n2989gat = (n1693gat)|(n1692gat);
assign n1265gat = ((~n1244gat)&(~n2969gat));
assign n720gat = ((~n919gat));
assign n123gat = ((~n130gat)&(~n126gat)&(~n129gat));
assign n570gat = ((~n577gat)&(~n573gat)&(~n576gat));
assign n2889gat = (n423gat)|(n362gat);
assign II2157 = ((~n312gat));
assign n137gat = ((~n154gat)&(~n253gat));
assign n1712gat = ((~II3179));
assign n281gat = ((~n271gat));
assign n1401gat = ((~n1584gat)&(~n1590gat));
assign n713gat = ((~n719gat)&(~n717gat)&(~n716gat));
assign n2754gat = ((~II4524));
assign n652gat = ((~n2789gat)&(~n93gat));
assign n3029gat = ((~II3315));
assign n1627gat = ((~n1618gat));
assign II2268 = ((~n2397gat));
assign n772gat = ((~n111gat)&(~n2842gat));
assign n1084gat = ((~n657gat));
assign n2268gat = ((~n2270gat));
assign n1683gat = ((~n1756gat));
assign n2019gat = ((~n2021gat));
assign n2678gat = ((~II4485));
assign II4750 = ((~n2810gat));
assign II4759 = ((~n2739gat));
assign n456gat = ((~n686gat));
assign n340gat = ((~II437));
assign II2271 = ((~n2201gat));
assign II1843 = ((~n2970gat));
assign II1190 = ((~n515gat));
assign n953gat = ((~II846));
assign n1118gat = ((~n1033gat));
assign n1892gat = ((~n2993gat));
assign n258gat = (n259gat)|(n260gat)|(n261gat)|(n262gat);
assign n2142gat = ((~II2672));
assign n1187gat = ((~n1194gat)&(~n1190gat)&(~n1193gat));
assign II594 = ((~n2722gat));
assign n2824gat = ((~II4389));
assign n2448gat = ((~n2450gat));
assign n3119gat = ((~II4699));
assign n1604gat = ((~n1778gat)&(~n1609gat)&(~n1702gat)&(~n1700gat));
assign II3530 = ((~n2396gat));
assign II1169 = ((~n837gat));
assign n352gat = ((~II729));
assign n2489gat = ((~II1606));
assign n2703gat = (n1755gat)|(n1518gat);
assign n1217gat = ((~n1223gat)&(~n1221gat)&(~n1220gat));
assign n3105gat = ((~II4657));
assign n2552gat = ((~II2420));
assign n670gat = ((~n636gat));
assign n1695gat = ((~n1609gat)&(~n1778gat)&(~n1704gat)&(~n1703gat));
assign n2803gat = ((~II4478));
assign n1755gat = ((~n1769gat)&(~n1773gat)&(~n2512gat));
assign n661gat = ((~n1725gat));
assign n2756gat = (n1011gat)|(n2244gat);
assign n70gat = ((~n71gat)&(~n2720gat));
assign n1032gat = ((~n1118gat));
assign n2546gat = ((~n2550gat)&(~n2551gat)&(~n2552gat));
assign n2585gat = ((~II2281));
assign n2265gat = ((~II3429));
assign n558gat = ((~n1725gat));
assign II1388 = ((~n819gat));
assign n1956gat = ((~n1898gat));
assign n1426gat = ((~n2011gat)&(~n1591gat));
assign n1801gat = ((~n2152gat)&(~n1989gat));
assign n950gat = ((~II815));
assign II3841 = ((~n2899gat));
assign n1293gat = ((~II877));
assign n2887gat = (n791gat)|(n650gat)|(n370gat);
assign II453 = ((~n701gat));
assign n1191gat = ((~II1786));
assign n2875gat = (n142gat)|(n40gat)|(n39gat);
assign n1990gat = ((~n2988gat));
assign n154gat = ((~n156gat));
assign n616gat = ((~n402gat));
assign n2017gat = ((~n1790gat)&(~n2016gat));
assign n761gat = ((~n855gat));
assign n868gat = ((~n2775gat)&(~n373gat));
assign II4633 = ((~n2805gat));
assign II1606 = ((~n2490gat));
assign n2198gat = ((~n2199gat)&(~n2058gat));
assign n1192gat = ((~II1791));
assign n251gat = ((~n1490gat)&(~n387gat));
assign n802gat = ((~n2882gat));
assign n2765gat = ((~II4138));
assign n233gat = ((~n243gat));
assign n1119gat = ((~n1121gat));
assign n1870gat = ((~II4626));
assign n1325gat = ((~n1444gat)&(~n164gat));
endmodule
