//NOTE: no-implementation module stub

module REG16LC (
    input DSPCLK,
    input MMR_web,
    input CKR_we,
    input [15:0] DMD,
    output [15:0] CKR,
    input PRST
);

endmodule
