module lcell (gnd, marker_bep_outwire);
  input gnd;
  output marker_bep_outwire;
endmodule