//NOTE: no-implementation module stub

module REG9LC (
    input DSPCLK,
    input MMR_web,
    input TSR_we,
    input [15:0] DMD,
    input [8:0] CLKsel,
    output [7:0] TSR,
    input T_RST
);
endmodule
