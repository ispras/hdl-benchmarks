//NOTE: no-implementation module stub

module coplogic (
    input wire SYSCLK,
    input wire TMODE,
    input wire RESET_D1_R_N,
    output wire EXCEPTION,
    input wire COPNO,
    input wire INSTSF,
    input wire INSTM32_S_R_N,
    output wire RHOLD,
    output wire DLOAD,
    input wire CMEMOPM_R,
    input wire CONDINN,
    input wire CPCONDN_R,
    input wire CRDADDR,
    output wire CRDGEN,
    output wire CRDCON,
    output wire CRDDATA,
    input wire CWRADDR_R,
    output wire CWRGEN_R,
    output wire CWRCON_R,
    output wire CWRDATA_R,
    output wire CDRIVERM_R,
    input wire CIDBUSINM,
    output wire CRDDATAM_R
);

endmodule
