// IWLS benchmark module "i10" printed on Wed May 29 16:34:21 2002
module i10(\V32(0) , \V32(1) , \V32(2) , \V32(3) , \V56(0) , \V289(0) , \V10(0) , \V13(0) , \V35(0) , \V203(0) , \V288(6) , \V288(7) , \V248(0) , \V249(0) , \V62(0) , \V59(0) , \V174(0) , \V215(0) , \V66(0) , \V70(0) , \V43(0) , \V214(0) , \V37(0) , \V271(0) , \V40(0) , \V45(0) , \V149(7) , \V149(6) , \V149(5) , \V149(4) , \V1(0) , \V7(0) , \V34(0) , \V243(0) , \V244(0) , \V245(0) , \V246(0) , \V247(0) , \V293(0) , \V302(0) , \V270(0) , \V269(0) , \V274(0) , \V202(0) , \V275(0) , \V257(7) , \V257(5) , \V257(3) , \V257(1) , \V257(2) , \V257(4) , \V257(6) , \V9(0) , \V149(0) , \V149(1) , \V149(2) , \V149(3) , \V169(1) , \V165(0) , \V165(2) , \V165(4) , \V165(5) , \V165(6) , \V165(7) , \V165(1) , \V88(2) , \V88(3) , \V55(0) , \V169(0) , \V52(0) , \V5(0) , \V6(0) , \V12(0) , \V11(0) , \V4(0) , \V165(3) , \V51(0) , \V65(0) , \V290(0) , \V279(0) , \V280(0) , \V288(4) , \V288(2) , \V288(0) , \V258(0) , \V229(5) , \V229(4) , \V229(3) , \V229(2) , \V229(1) , \V229(0) , \V223(5) , \V223(4) , \V223(3) , \V223(2) , \V223(1) , \V223(0) , \V189(5) , \V189(4) , \V189(3) , \V189(2) , \V189(1) , \V189(0) , \V183(5) , \V183(4) , \V183(3) , \V183(2) , \V183(1) , \V183(0) , \V239(4) , \V239(3) , \V239(2) , \V239(1) , \V239(0) , \V234(4) , \V234(3) , \V234(2) , \V234(1) , \V234(0) , \V199(4) , \V199(3) , \V199(2) , \V199(1) , \V199(0) , \V194(4) , \V194(3) , \V194(2) , \V194(1) , \V194(0) , \V257(0) , \V32(8) , \V32(7) , \V32(6) , \V32(5) , \V32(4) , \V32(11) , \V32(10) , \V32(9) , \V88(1) , \V88(0) , \V84(5) , \V84(4) , \V84(3) , \V84(2) , \V84(1) , \V84(0) , \V78(5) , \V78(4) , \V2(0) , \V3(0) , \V14(0) , \V213(0) , \V213(5) , \V213(4) , \V213(3) , \V213(2) , \V213(1) , \V268(5) , \V268(3) , \V268(1) , \V268(2) , \V268(4) , \V8(0) , \V60(0) , \V53(0) , \V57(0) , \V109(0) , \V277(0) , \V278(0) , \V259(0) , \V260(0) , \V67(0) , \V68(0) , \V69(0) , \V216(0) , \V175(0) , \V177(0) , \V172(0) , \V171(0) , \V50(0) , \V63(0) , \V71(0) , \V292(0) , \V291(0) , \V91(0) , \V91(1) , \V294(0) , \V207(0) , \V295(0) , \V204(0) , \V205(0) , \V261(0) , \V262(0) , \V100(0) , \V100(5) , \V100(4) , \V100(3) , \V100(2) , \V100(1) , \V240(0) , \V242(0) , \V241(0) , \V33(0) , \V16(0) , \V15(0) , \V101(0) , \V268(0) , \V288(1) , \V288(3) , \V288(5) , \V301(0) , \V108(0) , \V108(1) , \V108(2) , \V108(3) , \V108(4) , \V108(5) , \V124(5) , \V124(4) , \V124(3) , \V124(2) , \V124(1) , \V124(0) , \V132(7) , \V132(6) , \V132(5) , \V132(4) , \V132(3) , \V132(2) , \V132(1) , \V132(0) , \V118(5) , \V118(4) , \V118(3) , \V118(2) , \V118(1) , \V118(0) , \V118(7) , \V118(6) , \V46(0) , \V48(0) , \V102(0) , \V110(0) , \V134(1) , \V134(0) , \V272(0) , \V78(2) , \V78(3) , \V39(0) , \V38(0) , \V42(0) , \V44(0) , \V41(0) , \V78(1) , \V78(0) , \V94(0) , \V94(1) , \V321(2) , V356, V357, V373, \V375(0) , V377, \V393(0) , \V398(0) , \V410(0) , \V423(0) , V432, \V435(0) , \V500(0) , \V508(0) , \V511(0) , V512, V527, V537, V538, V539, V540, V541, V542, V543, V544, V545, V546, V547, V548, \V572(9) , \V572(8) , \V572(7) , \V572(6) , \V572(5) , \V572(4) , \V572(3) , \V572(2) , \V572(1) , \V572(0) , \V585(0) , V587, \V591(0) , \V597(0) , \V603(0) , \V609(0) , V620, V621, V630, \V634(0) , \V640(0) , V657, V707, V763, V775, V778, V779, V780, V781, V782, V783, V784, V787, V789, \V798(0) , V801, \V802(0) , \V821(0) , \V826(0) , V966, V986, \V1213(11) , \V1213(10) , \V1213(9) , \V1213(8) , \V1213(7) , \V1213(6) , \V1213(5) , \V1213(4) , \V1213(3) , \V1213(2) , \V1213(1) , \V1213(0) , \V1243(9) , \V1243(8) , \V1243(7) , \V1243(6) , \V1243(5) , \V1243(4) , \V1243(3) , \V1243(2) , \V1243(1) , \V1243(0) , V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263, V1264, V1265, V1266, V1267, \V1274(0) , \V1281(0) , \V1297(4) , \V1297(3) , \V1297(2) , \V1297(1) , \V1297(0) , V1365, V1375, V1378, V1380, V1382, V1384, V1386, V1387, \V1392(0) , V1423, V1426, V1428, V1429, V1431, V1432, \V1439(0) , \V1440(0) , \V1451(0) , \V1459(0) , \V1467(0) , V1470, \V1480(0) , \V1481(0) , \V1492(0) , \V1495(0) , \V1512(3) , \V1512(2) , \V1512(1) , \V1536(0) , V1537, V1539, \V1552(1) , \V1552(0) , \V1613(0) , \V1613(1) , \V1620(0) , \V1629(0) , \V1645(0) , \V1652(0) , V1669, \V1671(0) , \V1679(0) , \V1693(0) , \V1709(4) , \V1709(3) , \V1709(2) , \V1709(1) , \V1709(0) , \V1717(0) , V1719, \V1726(0) , V1736, \V1741(0) , \V1745(0) , \V1757(0) , \V1758(0) , \V1759(0) , \V1760(0) , \V1771(1) , \V1771(0) , \V1781(1) , \V1781(0) , \V1829(9) , \V1829(8) , \V1829(7) , \V1829(6) , \V1829(5) , \V1829(4) , \V1829(3) , \V1829(2) , \V1829(1) , \V1829(0) , V1832, \V1833(0) , \V1863(0) , \V1864(0) , \V1896(0) , \V1897(0) , \V1898(0) , \V1899(0) , \V1900(0) , \V1901(0) , \V1921(5) , \V1921(4) , \V1921(3) , \V1921(2) , \V1921(1) , \V1921(0) , \V1953(1) , \V1953(7) , \V1953(6) , \V1953(5) , \V1953(4) , \V1953(3) , \V1953(2) , \V1953(0) , \V1960(1) , \V1960(0) , \V1968(0) , \V1992(1) , \V1992(0) , V650, V651, V652, V653, V654, V655, V656, V1370, V1371, V1372, V1373, V1374);
input
  \V223(1) ,
  \V223(0) ,
  \V100(3) ,
  \V100(2) ,
  \V100(5) ,
  \V100(4) ,
  \V100(1) ,
  \V100(0) ,
  \V60(0) ,
  \V247(0) ,
  \V7(0) ,
  \V124(3) ,
  \V124(2) ,
  \V124(5) ,
  \V124(4) ,
  \V11(0) ,
  \V124(1) ,
  \V124(0) ,
  \V259(0) ,
  \V84(0) ,
  \V84(1) ,
  \V84(2) ,
  \V84(3) ,
  \V84(4) ,
  \V84(5) ,
  \V35(0) ,
  \V302(0) ,
  \V59(0) ,
  \V240(0) ,
  \V203(0) ,
  \V288(3) ,
  \V215(0) ,
  \V288(2) ,
  \V288(5) ,
  \V288(4) ,
  \V40(0) ,
  \V288(1) ,
  \V288(0) ,
  \V165(3) ,
  \V165(2) ,
  \V165(5) ,
  \V165(4) ,
  \V239(3) ,
  \V288(7) ,
  \V239(2) ,
  \V288(6) ,
  \V52(0) ,
  \V165(1) ,
  \V239(4) ,
  \V165(0) ,
  \V239(1) ,
  \V239(0) ,
  \V165(7) ,
  \V165(6) ,
  \V177(0) ,
  \V189(3) ,
  \V189(2) ,
  \V189(5) ,
  \V189(4) ,
  \V189(1) ,
  \V189(0) ,
  \V15(0) ,
  \V88(0) ,
  \V88(1) ,
  \V88(2) ,
  \V88(3) ,
  \V39(0) ,
  \V293(0) ,
  \V244(0) ,
  \V4(0) ,
  \V194(3) ,
  \V194(2) ,
  \V194(4) ,
  \V268(3) ,
  \V268(2) ,
  \V268(5) ,
  \V194(1) ,
  \V268(4) ,
  \V194(0) ,
  \V268(1) ,
  \V268(0) ,
  \V207(0) ,
  \V32(0) ,
  \V32(1) ,
  \V32(2) ,
  \V32(3) ,
  \V32(4) ,
  \V32(5) ,
  \V32(6) ,
  \V32(7) ,
  \V32(8) ,
  \V44(0) ,
  \V32(9) ,
  \V108(3) ,
  \V108(2) ,
  \V56(0) ,
  \V108(5) ,
  \V108(4) ,
  \V169(1) ,
  \V169(0) ,
  \V108(1) ,
  \V108(0) ,
  \V68(0) ,
  \V261(0) ,
  \V101(0) ,
  \V174(0) ,
  \V248(0) ,
  \V8(0) ,
  \V12(0) ,
  \V149(3) ,
  \V149(2) ,
  \V149(5) ,
  \V149(4) ,
  \V149(1) ,
  \V149(0) ,
  \V149(7) ,
  \V149(6) ,
  \V48(0) ,
  \V290(0) ,
  \V32(11) ,
  \V32(10) ,
  \V241(0) ,
  \V1(0) ,
  \V204(0) ,
  \V277(0) ,
  \V216(0) ,
  \V41(0) ,
  \V289(0) ,
  \V53(0) ,
  \V65(0) ,
  \V16(0) ,
  \V270(0) ,
  \V294(0) ,
  \V171(0) ,
  \V183(3) ,
  \V110(0) ,
  \V183(2) ,
  \V245(0) ,
  \V183(5) ,
  \V5(0) ,
  \V183(4) ,
  \V257(3) ,
  \V257(2) ,
  \V70(0) ,
  \V257(5) ,
  \V183(1) ,
  \V257(4) ,
  \V183(0) ,
  \V257(1) ,
  \V257(0) ,
  \V257(7) ,
  \V257(6) ,
  \V134(1) ,
  \V134(0) ,
  \V269(0) ,
  \V94(0) ,
  \V94(1) ,
  \V33(0) ,
  \V45(0) ,
  \V57(0) ,
  \V109(0) ,
  \V69(0) ,
  \V262(0) ,
  \V213(3) ,
  \V213(2) ,
  \V213(5) ,
  \V213(4) ,
  \V274(0) ,
  \V213(1) ,
  \V213(0) ,
  \V50(0) ,
  \V102(0) ,
  \V62(0) ,
  \V175(0) ,
  \V249(0) ,
  \V9(0) ,
  \V13(0) ,
  \V199(3) ,
  \V199(2) ,
  \V199(4) ,
  \V199(1) ,
  \V199(0) ,
  \V37(0) ,
  \V291(0) ,
  \V242(0) ,
  \V2(0) ,
  \V205(0) ,
  \V91(0) ,
  \V91(1) ,
  \V278(0) ,
  \V229(3) ,
  \V229(2) ,
  \V42(0) ,
  \V229(5) ,
  \V229(4) ,
  \V229(1) ,
  \V229(0) ,
  \V118(3) ,
  \V118(2) ,
  \V66(0) ,
  \V118(5) ,
  \V118(4) ,
  \V118(1) ,
  \V118(0) ,
  \V78(0) ,
  \V78(1) ,
  \V118(7) ,
  \V78(2) ,
  \V118(6) ,
  \V78(3) ,
  \V78(4) ,
  \V78(5) ,
  \V271(0) ,
  \V234(3) ,
  \V234(2) ,
  \V234(4) ,
  \V295(0) ,
  \V234(1) ,
  \V234(0) ,
  \V172(0) ,
  \V246(0) ,
  \V6(0) ,
  \V71(0) ,
  \V10(0) ,
  \V258(0) ,
  \V34(0) ,
  \V46(0) ,
  \V301(0) ,
  \V202(0) ,
  \V275(0) ,
  \V214(0) ,
  \V51(0) ,
  \V63(0) ,
  \V14(0) ,
  \V38(0) ,
  \V280(0) ,
  \V292(0) ,
  \V243(0) ,
  \V3(0) ,
  \V132(3) ,
  \V132(2) ,
  \V132(5) ,
  \V132(4) ,
  \V132(1) ,
  \V132(0) ,
  \V132(7) ,
  \V132(6) ,
  \V279(0) ,
  \V43(0) ,
  \V55(0) ,
  \V67(0) ,
  \V260(0) ,
  \V272(0) ,
  \V223(3) ,
  \V223(2) ,
  \V223(5) ,
  \V223(4) ;
output
  \V1243(7) ,
  \V500(0) ,
  \V1243(6) ,
  \V1243(9) ,
  \V1243(8) ,
  \V1243(1) ,
  \V1243(0) ,
  \V1717(0) ,
  \V1243(3) ,
  \V1243(2) ,
  \V1243(5) ,
  \V1243(4) ,
  \V585(0) ,
  \V597(0) ,
  \V1679(0) ,
  \V1833(0) ,
  \V1968(0) ,
  \V1771(1) ,
  \V1771(0) ,
  \V640(0) ,
  \V375(0) ,
  \V603(0) ,
  \V1758(0) ,
  \V1900(0) ,
  \V1709(1) ,
  \V1709(0) ,
  \V1709(3) ,
  \V1709(2) ,
  \V1709(4) ,
  \V1512(1) ,
  \V1512(3) ,
  \V1512(2) ,
  \V1536(0) ,
  \V1898(0) ,
  \V1652(0) ,
  \V1726(0) ,
  \V1953(7) ,
  \V1953(6) ,
  \V410(0) ,
  \V1953(1) ,
  \V1953(0) ,
  \V1953(3) ,
  \V1953(2) ,
  \V1953(5) ,
  \V1953(4) ,
  \V508(0) ,
  \V1392(0) ,
  \V1829(7) ,
  \V1829(6) ,
  \V1829(9) ,
  \V1829(8) ,
  \V1281(0) ,
  \V1620(0) ,
  \V1829(1) ,
  \V1829(0) ,
  \V1829(3) ,
  \V1829(2) ,
  \V1693(0) ,
  \V1829(5) ,
  \V1829(4) ,
  \V1921(1) ,
  \V1921(0) ,
  \V1921(3) ,
  \V1921(2) ,
  \V1921(5) ,
  \V1921(4) ,
  \V802(0) ,
  \V826(0) ,
  \V1213(10) ,
  \V1213(11) ,
  \V1760(0) ,
  \V1495(0) ,
  \V591(0) ,
  \V1759(0) ,
  \V1901(0) ,
  \V1297(1) ,
  \V1297(0) ,
  \V1297(3) ,
  \V1297(2) ,
  \V1297(4) ,
  \V1451(0) ,
  \V1863(0) ,
  \V393(0) ,
  \V1899(0) ,
  \V1480(0) ,
  \V423(0) ,
  \V1492(0) ,
  \V435(0) ,
  \V1781(1) ,
  \V1781(0) ,
  V1256,
  V1257,
  V1258,
  V1259,
  V1260,
  V1261,
  V1262,
  V1263,
  V1264,
  V1265,
  V1266,
  V1267,
  \V1467(0) ,
  V1365,
  V1370,
  V1371,
  V1372,
  V1373,
  V1374,
  V1375,
  V1378,
  V1380,
  V1382,
  V1384,
  V1386,
  V1387,
  V1423,
  V1426,
  V1428,
  V1429,
  V1431,
  V1432,
  V1470,
  \V1645(0) ,
  V1537,
  V1539,
  V1669,
  V1719,
  \V1896(0) ,
  V1736,
  V1832,
  \V1459(0) ,
  \V1213(7) ,
  \V1213(6) ,
  \V1213(9) ,
  \V1213(8) ,
  \V1613(1) ,
  \V1274(0) ,
  \V1613(0) ,
  \V1213(1) ,
  \V1213(0) ,
  \V1213(3) ,
  \V1213(2) ,
  \V1213(5) ,
  \V1213(4) ,
  \V1440(0) ,
  \V321(2) ,
  \V1864(0) ,
  \V1741(0) ,
  \V572(3) ,
  \V572(2) ,
  \V634(0) ,
  \V572(5) ,
  \V572(4) ,
  \V1439(0) ,
  \V572(1) ,
  \V572(0) ,
  \V511(0) ,
  \V572(7) ,
  \V572(6) ,
  \V572(9) ,
  \V572(8) ,
  \V1992(1) ,
  \V1992(0) ,
  \V609(0) ,
  \V1481(0) ,
  \V1629(0) ,
  \V798(0) ,
  \V398(0) ,
  \V1671(0) ,
  \V1745(0) ,
  \V1757(0) ,
  \V1960(1) ,
  \V1960(0) ,
  V356,
  V357,
  V373,
  V377,
  \V1897(0) ,
  V432,
  V512,
  V527,
  V537,
  V538,
  V539,
  V540,
  V541,
  V542,
  V543,
  V544,
  V545,
  V546,
  V547,
  V548,
  V587,
  V620,
  V621,
  V630,
  V650,
  V651,
  V652,
  V653,
  V654,
  V655,
  V656,
  V657,
  \V821(0) ,
  \V1552(1) ,
  \V1552(0) ,
  V707,
  V763,
  V775,
  V778,
  V779,
  V780,
  V781,
  V782,
  V783,
  V784,
  V787,
  V789,
  V801,
  V966,
  V986;
wire
  \V758(0) ,
  \V1354(0) ,
  \V1631(0) ,
  \V985(0) ,
  \V450(0) ,
  \V1255(1) ,
  \V1255(0) ,
  \V1255(3) ,
  \V1255(2) ,
  \V536(0) ,
  \[200] ,
  \[201] ,
  \[202] ,
  \[203] ,
  \V1124(12) ,
  \[204] ,
  \V1124(13) ,
  \[205] ,
  \V813(0) ,
  \[206] ,
  \[207] ,
  \V413(0) ,
  \[208] ,
  \[209] ,
  \V1124(10) ,
  \V1124(11) ,
  \V1421(0) ,
  \[210] ,
  \[211] ,
  \V2033(0) ,
  \[212] ,
  \[213] ,
  \[214] ,
  \[215] ,
  \[216] ,
  \[217] ,
  \[218] ,
  \[219] ,
  \[220] ,
  \[221] ,
  \[222] ,
  \[223] ,
  \V1069(7) ,
  \V1069(6) ,
  \V1069(9) ,
  \V1069(8) ,
  \V1395(0) ,
  \V1334(0) ,
  \V1069(5) ,
  \V1069(4) ,
  \V1623(0) ,
  \V965(0) ,
  \V504(0) ,
  \V1647(0) ,
  \V1124(7) ,
  \V1124(6) ,
  \V1124(9) ,
  \V1124(8) ,
  \V380(0) ,
  \V1124(3) ,
  \V731(0) ,
  \V1124(2) ,
  \V1124(5) ,
  \V1597(0) ,
  \V1124(4) ,
  \V405(0) ,
  \V817(0) ,
  \V1351(0) ,
  \V1086(1) ,
  \V1086(0) ,
  \V1086(3) ,
  \V1086(2) ,
  \V1437(0) ,
  \V982(0) ,
  \V1399(0) ,
  \V1553(0) ,
  \V1177(7) ,
  \V1177(6) ,
  \V1177(9) ,
  \V1177(8) ,
  \[10] ,
  \[11] ,
  \V1977(0) ,
  \[12] ,
  \[13] ,
  \[14] ,
  \[15] ,
  \V1177(1) ,
  \[16] ,
  \V1177(0) ,
  \[17] ,
  \V1177(3) ,
  \[18] ,
  \V1177(2) ,
  \[19] ,
  \V1177(5) ,
  \V1854(0) ,
  \V1177(4) ,
  \V384(0) ,
  \[20] ,
  \[21] ,
  \[22] ,
  \[23] ,
  \V396(0) ,
  \[24] ,
  \[25] ,
  \V1331(0) ,
  \[26] ,
  \V2078(0) ,
  \[27] ,
  \[28] ,
  \[29] ,
  \V612(0) ,
  \[30] ,
  \[31] ,
  \V1417(0) ,
  \V1681(0) ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \V759(0) ,
  \[36] ,
  \[37] ,
  \[38] ,
  \[39] ,
  \V1632(0) ,
  \[40] ,
  \[41] ,
  \[42] ,
  \V1306(0) ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ,
  \[59] ,
  \V1268(0) ,
  \V1471(0) ,
  \V1069(10) ,
  \[60] ,
  \V1069(11) ,
  \[61] ,
  \V414(0) ,
  \[62] ,
  \[63] ,
  \[64] ,
  \[65] ,
  \[66] ,
  \[67] ,
  \V487(0) ,
  \[68] ,
  \[69] ,
  \V1422(0) ,
  \V1360(0) ,
  \[70] ,
  \[71] ,
  \[72] ,
  \[73] ,
  \[74] ,
  \[75] ,
  \[76] ,
  \[77] ,
  \[78] ,
  \V1711(0) ,
  \[79] ,
  \V376(0) ,
  \V1311(0) ,
  \V2058(0) ,
  \V788(0) ,
  \[80] ,
  \[81] ,
  \[82] ,
  \[83] ,
  \[84] ,
  \[85] ,
  \[86] ,
  \[87] ,
  \[88] ,
  \[89] ,
  \V1396(0) ,
  \[90] ,
  \V1409(0) ,
  \[91] ,
  \[92] ,
  \[93] ,
  \[94] ,
  \[95] ,
  \[96] ,
  \[97] ,
  \[98] ,
  \[99] ,
  \V2002(0) ,
  \V1463(0) ,
  \V467(0) ,
  \V1340(0) ,
  \V1475(0) ,
  \V2087(0) ,
  \V2038(0) ,
  \V633(0) ,
  \V1641(0) ,
  \V1653(0) ,
  V1000,
  V1002,
  V1004,
  V1006,
  V1008,
  V1010,
  V1012,
  V1014,
  V1016,
  V1018,
  V1020,
  V1022,
  V1024,
  V1025,
  V1026,
  V1027,
  V1028,
  V1029,
  V1030,
  V1031,
  V1032,
  V1033,
  V1034,
  V1036,
  V1038,
  V1040,
  V1042,
  V1044,
  V1046,
  V1048,
  V1050,
  V1052,
  V1054,
  V1055,
  V1056,
  V1057,
  V1058,
  V1059,
  V1060,
  V1061,
  \V1554(0) ,
  V1070,
  V1071,
  V1072,
  V1073,
  V1074,
  V1075,
  V1076,
  V1077,
  V1078,
  V1079,
  V1081,
  V1083,
  V1085,
  V1087,
  V1088,
  V1089,
  V1090,
  V1092,
  V1093,
  V1094,
  V1095,
  V1096,
  V1097,
  V1098,
  V1099,
  \V1831(0) ,
  \V496(0) ,
  V1100,
  V1101,
  V1103,
  V1105,
  V1107,
  V1109,
  V1111,
  V1113,
  V1115,
  V1117,
  V1119,
  V1121,
  V1123,
  V1125,
  V1127,
  V1128,
  V1129,
  V1130,
  V1131,
  V1132,
  V1133,
  V1134,
  V1136,
  V1138,
  V1140,
  V1142,
  V1144,
  V1146,
  V1148,
  V1149,
  V1150,
  V1151,
  V1152,
  V1153,
  V1154,
  V1155,
  V1156,
  V1157,
  V1158,
  V1160,
  V1162,
  V1164,
  V1166,
  V1168,
  V1170,
  V1172,
  V1174,
  V1176,
  V1178,
  V1179,
  V1180,
  V1181,
  V1182,
  V1183,
  V1184,
  V1185,
  V1186,
  V1187,
  V1188,
  V1189,
  V1190,
  V1192,
  V1194,
  V1196,
  V1198,
  \V1855(0) ,
  \V385(0) ,
  V1200,
  V1202,
  V1204,
  V1206,
  V1208,
  V1210,
  V1212,
  V1214,
  V1215,
  V1216,
  V1217,
  V1218,
  V1219,
  \V1455(0) ,
  V1220,
  V1221,
  V1222,
  V1223,
  V1224,
  V1226,
  V1228,
  \V2067(0) ,
  V1230,
  V1232,
  V1234,
  V1236,
  V1238,
  V1240,
  V1242,
  V1244,
  V1245,
  V1246,
  V1247,
  V1248,
  V1250,
  V1252,
  V1254,
  V1272,
  V1273,
  V1276,
  V1279,
  V1280,
  V1283,
  V1284,
  V1285,
  V1286,
  V1287,
  V1288,
  V1290,
  V1292,
  V1294,
  V1296,
  V1298,
  V1299,
  \V336(0) ,
  \V2018(0) ,
  V1300,
  V1301,
  V1302,
  V1303,
  V1304,
  V1305,
  V1307,
  V1308,
  V1309,
  V1310,
  V1312,
  V1316,
  V1317,
  V1318,
  V1319,
  V1320,
  V1324,
  V1325,
  V1326,
  V1327,
  V1328,
  V1329,
  V1330,
  V1332,
  V1333,
  V1335,
  V1336,
  V1338,
  V1339,
  V1344,
  V1345,
  V1346,
  V1347,
  V1348,
  V1349,
  V1350,
  V1352,
  V1353,
  V1355,
  V1356,
  V1358,
  V1359,
  V1366,
  V1367,
  V1368,
  V1369,
  V1390,
  V1391,
  V1393,
  V1402,
  V1403,
  V1404,
  V1406,
  V1407,
  V1411,
  V1412,
  V1413,
  V1414,
  V1416,
  V1418,
  V1425,
  V1427,
  V1435,
  V1436,
  V1438,
  V1443,
  V1445,
  V1448,
  V1450,
  V1453,
  V1454,
  V1456,
  V1458,
  V1461,
  V1462,
  V1464,
  V1466,
  V1473,
  V1474,
  V1476,
  V1478,
  V1479,
  V1486,
  V1490,
  V1491,
  V1494,
  V1497,
  \V1983(0) ,
  V1501,
  V1503,
  V1504,
  V1505,
  V1507,
  V1509,
  V1511,
  V1513,
  V1516,
  V1517,
  V1518,
  V1524,
  V1526,
  V1527,
  V1532,
  V1535,
  V1545,
  V1547,
  V1548,
  V1549,
  V1551,
  V1555,
  V1557,
  V1558,
  V1564,
  V1568,
  V1569,
  V1570,
  V1571,
  V1572,
  V1579,
  V1580,
  V1581,
  V1582,
  V1583,
  V1584,
  V1585,
  V1586,
  V1587,
  V1588,
  V1589,
  V1590,
  V1591,
  V1592,
  V1593,
  V1594,
  V1598,
  V1599,
  \V2011(0) ,
  V1600,
  V1601,
  V1602,
  V1603,
  V1604,
  V1605,
  V1606,
  V1607,
  V1608,
  V1609,
  V1610,
  V1611,
  V1614,
  V1615,
  V1616,
  V1621,
  V1622,
  V1624,
  V1628,
  \V1472(0) ,
  V1633,
  V1634,
  V1635,
  V1636,
  V1637,
  V1638,
  V1639,
  V1640,
  \V476(0) ,
  V1643,
  V1644,
  V1646,
  \V2084(0) ,
  V1648,
  V1651,
  V1656,
  V1660,
  V1662,
  V1663,
  \V1546(0) ,
  V1664,
  \V1023(7) ,
  V1672,
  V1673,
  V1675,
  V1678,
  \V1023(6) ,
  V1683,
  V1686,
  V1688,
  \V1023(9) ,
  V1691,
  V1692,
  V1695,
  V1696,
  V1697,
  V1698,
  V1699,
  \V1023(8) ,
  \V1023(10) ,
  \V1023(11) ,
  V1700,
  V1702,
  V1704,
  V1706,
  V1708,
  \V1023(1) ,
  V1710,
  V1712,
  V1716,
  \V1023(0) ,
  V1721,
  V1723,
  V1725,
  V1729,
  \V1023(3) ,
  V1730,
  V1731,
  V1732,
  V1733,
  V1735,
  V1738,
  V1739,
  \V1023(2) ,
  V1740,
  V1744,
  V1748,
  V1749,
  \V1023(5) ,
  V1750,
  V1751,
  V1752,
  V1754,
  V1755,
  V1756,
  \V1835(0) ,
  \V1023(4) ,
  V1764,
  V1765,
  V1768,
  V1770,
  V1774,
  V1775,
  V1778,
  V1780,
  V1792,
  V1793,
  V1794,
  V1795,
  V1796,
  V1797,
  V1798,
  V1799,
  \V777(0) ,
  V1800,
  V1801,
  \V1447(0) ,
  V1810,
  V1812,
  V1814,
  V1816,
  V1818,
  V1820,
  V1822,
  V1824,
  V1826,
  V1828,
  V1830,
  V1834,
  V1836,
  V1838,
  V1839,
  V1840,
  V1842,
  V1844,
  V1846,
  V1848,
  V1850,
  V1852,
  V1867,
  V1868,
  V1869,
  V1870,
  V1871,
  V1872,
  V1873,
  V1874,
  V1875,
  V1876,
  V1877,
  V1878,
  V1879,
  V1880,
  V1881,
  V1882,
  V1883,
  V1885,
  V1886,
  V1887,
  \[0] ,
  V1889,
  V1890,
  V1891,
  V1892,
  V1893,
  V1895,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \[5] ,
  \[6] ,
  \[7] ,
  \V1397(0) ,
  V1902,
  V1904,
  V1905,
  V1906,
  V1907,
  V1908,
  \[8] ,
  V1909,
  V1910,
  V1912,
  V1914,
  V1916,
  V1918,
  \[9] ,
  V1920,
  V1922,
  V1923,
  V1924,
  V1925,
  V1926,
  V1927,
  V1928,
  V1929,
  V1930,
  V1931,
  V1932,
  V1933,
  V1934,
  V1935,
  V1936,
  V1937,
  V1938,
  V1940,
  V1941,
  V1943,
  V1945,
  V1947,
  V1949,
  V1951,
  V1954,
  V1955,
  V1956,
  V1957,
  V1959,
  \V1674(0) ,
  V1961,
  V1962,
  V1966,
  V1967,
  V1972,
  V1973,
  V1974,
  V1978,
  V1979,
  V1981,
  V1982,
  V1986,
  V1987,
  V1988,
  V1989,
  V1991,
  V1994,
  V1995,
  V1996,
  V1997,
  \V629(0) ,
  \V1963(0) ,
  \V493(0) ,
  \V382(0) ,
  \V2064(0) ,
  \V1999(0) ,
  \V807(0) ,
  \V1538(0) ,
  \V1415(0) ,
  \V1642(0) ,
  \V1728(0) ,
  \[100] ,
  \[101] ,
  \[102] ,
  \[103] ,
  \[104] ,
  \V473(0) ,
  \[105] ,
  \V2081(0) ,
  \V812(0) ,
  \[106] ,
  \[107] ,
  \V412(0) ,
  \[108] ,
  \[109] ,
  V2000,
  V2001,
  V2003,
  V2005,
  V2006,
  V2009,
  V2012,
  V2013,
  V2014,
  V2015,
  V2021,
  V2023,
  V2025,
  V2026,
  V2027,
  V2028,
  V2029,
  V2030,
  V2031,
  V2032,
  V2034,
  V2035,
  V2036,
  V2037,
  V2039,
  V2043,
  V2044,
  V2045,
  V2046,
  V2047,
  V2051,
  V2052,
  V2053,
  V2054,
  V2055,
  V2056,
  V2057,
  V2059,
  V2060,
  V2062,
  V2063,
  V2065,
  V2066,
  \[110] ,
  V2071,
  V2072,
  V2073,
  V2074,
  V2075,
  V2076,
  V2077,
  V2079,
  \V424(0) ,
  \[111] ,
  V2080,
  V2082,
  V2083,
  V2085,
  V2086,
  \[112] ,
  \[113] ,
  \[114] ,
  \V762(0) ,
  \[115] ,
  \[116] ,
  \[117] ,
  \[118] ,
  \[119] ,
  V2104,
  V2106,
  V2107,
  V2109,
  V2115,
  V2116,
  V2119,
  V2122,
  V2157,
  \[120] ,
  \[121] ,
  V2188,
  V2189,
  \[122] ,
  \[123] ,
  \[124] ,
  \[125] ,
  \[126] ,
  \[127] ,
  \[128] ,
  \V1856(0) ,
  \V386(0) ,
  \[129] ,
  V2208,
  V2209,
  V2212,
  V2213,
  V2216,
  V2217,
  V2220,
  V2221,
  V2224,
  V2225,
  V2228,
  V2229,
  V2232,
  V2233,
  V2236,
  V2237,
  V2240,
  V2241,
  V2244,
  V2245,
  V2248,
  V2249,
  V2252,
  V2253,
  V2256,
  V2257,
  \V2007(0) ,
  V2260,
  V2261,
  V2264,
  V2265,
  V2268,
  V2269,
  \[130] ,
  V2272,
  V2273,
  V2276,
  V2277,
  \V1394(0) ,
  \[131] ,
  V2280,
  V2281,
  V2284,
  V2285,
  V2288,
  V2289,
  \[132] ,
  V2292,
  V2293,
  V2296,
  V2297,
  \[133] ,
  \[134] ,
  \[135] ,
  \[136] ,
  \[137] ,
  \V2019(0) ,
  \[138] ,
  \[139] ,
  V2300,
  V2301,
  V2304,
  V2305,
  V2308,
  V2309,
  V2312,
  V2313,
  V2316,
  V2317,
  V2320,
  V2321,
  V2324,
  V2325,
  V2328,
  V2329,
  V2332,
  V2333,
  V2336,
  V2337,
  V2340,
  V2341,
  V2344,
  V2345,
  V2348,
  V2349,
  V2352,
  V2353,
  V2356,
  V2357,
  V2360,
  V2361,
  V2364,
  V2365,
  V2368,
  V2369,
  \[140] ,
  V2372,
  V2373,
  V2376,
  V2377,
  \[141] ,
  V2380,
  V2381,
  V2384,
  V2385,
  V2388,
  V2389,
  \[142] ,
  V2392,
  V2393,
  V2396,
  V2397,
  \[143] ,
  \[144] ,
  \[145] ,
  \V1357(0) ,
  \[146] ,
  \V490(0) ,
  \[147] ,
  \[148] ,
  \[149] ,
  V2400,
  V2401,
  V2404,
  V2405,
  V2408,
  V2409,
  V2412,
  V2413,
  V2416,
  V2417,
  V2420,
  V2421,
  V2424,
  V2425,
  V2428,
  V2429,
  V2432,
  V2433,
  V2436,
  \V503(0) ,
  V2437,
  V2440,
  V2441,
  V2444,
  V2445,
  V2448,
  V2449,
  V2452,
  V2453,
  V2456,
  V2457,
  V2460,
  V2461,
  V2464,
  V2465,
  V2468,
  V2469,
  \[150] ,
  V2472,
  V2473,
  V2476,
  V2477,
  \[151] ,
  V2480,
  V2481,
  V2484,
  V2485,
  V2488,
  V2489,
  \[152] ,
  V2492,
  V2493,
  V2496,
  V2497,
  \[153] ,
  \[154] ,
  \[155] ,
  \[156] ,
  \[157] ,
  \V1984(0) ,
  \[158] ,
  \[159] ,
  V2500,
  V2501,
  V2504,
  V2505,
  V2508,
  V2509,
  V2512,
  V2513,
  V2516,
  V2517,
  V2520,
  V2521,
  V2524,
  V2525,
  V2528,
  \V2061(0) ,
  V2529,
  V2532,
  V2533,
  V2536,
  V2537,
  V2540,
  V2541,
  V2544,
  V2545,
  V2548,
  V2549,
  V2552,
  V2553,
  V2556,
  V2557,
  V2560,
  V2561,
  V2564,
  V2565,
  V2568,
  V2569,
  \[160] ,
  V2572,
  V2573,
  V2576,
  V2577,
  \[161] ,
  V2580,
  V2581,
  \V391(0) ,
  V2584,
  V2585,
  \V730(0) ,
  V2588,
  V2589,
  \[162] ,
  V2592,
  V2593,
  V2596,
  V2597,
  \[163] ,
  \[164] ,
  \[165] ,
  \[166] ,
  \V1147(7) ,
  \[167] ,
  \V404(0) ,
  \V1147(6) ,
  \[168] ,
  \V1147(9) ,
  \[169] ,
  V2600,
  V2601,
  V2604,
  V2605,
  V2608,
  V2609,
  \V1147(8) ,
  V2612,
  V2613,
  V2616,
  V2617,
  V2620,
  V2621,
  V2624,
  V2625,
  V2628,
  V2629,
  V2632,
  V2633,
  V2636,
  V2637,
  V2640,
  V2641,
  V323,
  V2644,
  V324,
  V2645,
  V325,
  V326,
  V2648,
  V2649,
  V329,
  V2652,
  V332,
  V2653,
  V335,
  V2656,
  V2657,
  V339,
  V2660,
  V340,
  V2661,
  V341,
  V2664,
  V2665,
  V345,
  V347,
  V2668,
  V348,
  V2669,
  V349,
  \[170] ,
  V350,
  V351,
  V2672,
  V352,
  V2673,
  V353,
  V354,
  V355,
  V2676,
  V2677,
  V358,
  V359,
  \[171] ,
  V2680,
  V360,
  V2681,
  V2684,
  V2685,
  V2688,
  V2689,
  \[172] ,
  V2692,
  V372,
  V2693,
  V2696,
  V2697,
  V379,
  \[173] ,
  V387,
  V388,
  V389,
  \[174] ,
  V390,
  V392,
  V395,
  V397,
  \V1147(5) ,
  \[175] ,
  \[176] ,
  \[177] ,
  \[178] ,
  \[179] ,
  V2700,
  V2701,
  V2704,
  V2705,
  V2708,
  V2709,
  V2712,
  V2713,
  V2716,
  V2717,
  V2720,
  V400,
  V2721,
  V401,
  V402,
  V2724,
  V2725,
  V406,
  V407,
  V2728,
  V2729,
  V409,
  V411,
  V2732,
  V2733,
  V415,
  V2736,
  V416,
  V2737,
  V417,
  V419,
  V2740,
  V420,
  V2741,
  V421,
  V422,
  V2744,
  V2745,
  V425,
  V2748,
  V2749,
  V2752,
  V2753,
  V433,
  V2756,
  V2757,
  V437,
  V438,
  V439,
  V2760,
  V440,
  V2761,
  V441,
  V442,
  V443,
  V2764,
  V444,
  V2765,
  V446,
  V447,
  V2768,
  V448,
  V2769,
  V449,
  \[180] ,
  V451,
  V2772,
  V452,
  V2773,
  V453,
  V454,
  V455,
  V2776,
  V456,
  V2777,
  \[181] ,
  V2780,
  V460,
  V2781,
  V461,
  V462,
  V463,
  V2784,
  V464,
  V2785,
  V465,
  V466,
  V2788,
  V468,
  V2789,
  V469,
  \[182] ,
  V471,
  V2792,
  V472,
  V2793,
  V474,
  V475,
  V2796,
  V2797,
  \[183] ,
  V480,
  V481,
  V482,
  V483,
  V484,
  V485,
  V486,
  V488,
  V489,
  \[184] ,
  V491,
  V492,
  V494,
  V495,
  V499,
  \[185] ,
  \[186] ,
  \V1147(10) ,
  \[187] ,
  \V1147(11) ,
  \V378(0) ,
  \[188] ,
  \[189] ,
  V2800,
  V2801,
  V2804,
  V2805,
  V2808,
  V2809,
  V2812,
  V2813,
  V2816,
  V2817,
  V501,
  V502,
  V505,
  V506,
  V507,
  V509,
  V513,
  V514,
  V515,
  V516,
  V517,
  V518,
  V525,
  V529,
  V530,
  V531,
  V534,
  V535,
  V549,
  \[190] ,
  V550,
  V551,
  V552,
  V553,
  V555,
  V557,
  V559,
  \[191] ,
  \V729(0) ,
  V561,
  V563,
  V565,
  V567,
  V569,
  \[192] ,
  V571,
  V573,
  V574,
  V575,
  V576,
  V577,
  V578,
  V579,
  \[193] ,
  V580,
  V581,
  V582,
  V589,
  \[194] ,
  V590,
  V593,
  V594,
  V596,
  V599,
  \[195] ,
  \[196] ,
  \[197] ,
  \[198] ,
  \V1398(0) ,
  \[199] ,
  V600,
  V602,
  V605,
  V606,
  V608,
  \V1337(0) ,
  V611,
  V613,
  V614,
  V615,
  V616,
  \V470(0) ,
  V623,
  V626,
  V627,
  V628,
  V631,
  V632,
  V637,
  V638,
  V644,
  V645,
  V646,
  V647,
  V648,
  V649,
  V687,
  V695,
  V696,
  V697,
  V698,
  \V1687(0) ,
  V700,
  V701,
  V702,
  V703,
  V704,
  V706,
  V710,
  V711,
  V712,
  V713,
  V714,
  V715,
  V716,
  V717,
  V718,
  V719,
  V720,
  V721,
  V722,
  V723,
  V724,
  V725,
  V726,
  V727,
  V728,
  V734,
  V735,
  V736,
  V737,
  V738,
  V739,
  V740,
  V741,
  V742,
  V743,
  V744,
  V745,
  V746,
  V747,
  V748,
  V749,
  V750,
  V751,
  V755,
  V756,
  V757,
  V761,
  V766,
  V767,
  V768,
  V769,
  V774,
  V776,
  V790,
  V794,
  V797,
  V799,
  \V1053(7) ,
  \V445(0) ,
  \V1053(6) ,
  V806,
  V808,
  \V1053(9) ,
  V811,
  V814,
  V815,
  V816,
  V818,
  \V1053(8) ,
  V820,
  V823,
  V824,
  V825,
  V828,
  V829,
  V830,
  V831,
  V836,
  V838,
  V839,
  V840,
  V841,
  V846,
  V848,
  V849,
  \V1853(0) ,
  V850,
  V851,
  \V383(0) ,
  V856,
  V858,
  V859,
  V860,
  V861,
  V866,
  V868,
  V869,
  V870,
  V871,
  V876,
  V878,
  V879,
  V880,
  V881,
  V886,
  V888,
  V889,
  \V1053(1) ,
  V890,
  V891,
  V896,
  V898,
  V899,
  \V1053(0) ,
  \V1053(3) ,
  \V1053(2) ,
  \V1053(5) ,
  \V1053(4) ,
  V900,
  V901,
  V906,
  V908,
  V909,
  V910,
  V911,
  V916,
  V918,
  V919,
  V920,
  V921,
  V926,
  V928,
  V929,
  V930,
  V931,
  V936,
  V938,
  V939,
  V940,
  V941,
  \V408(0) ,
  V946,
  V952,
  V953,
  V954,
  V955,
  V960,
  V961,
  V962,
  V963,
  V968,
  V976,
  V978,
  V981,
  V983,
  V984,
  V988,
  V989,
  V990,
  V991,
  V992,
  V993,
  V994,
  V995,
  V996,
  V997,
  V998,
  V999;
assign
  \V758(0)  = V756 | (V755 | V757),
  \V1354(0)  = V1353 | V1352,
  \V1631(0)  = V766 | V769,
  \V1243(7)  = \[84] ,
  \V500(0)  = \[12] ,
  \V1243(6)  = \[85] ,
  \V1243(9)  = \[82] ,
  \V1243(8)  = \[83] ,
  \V1243(1)  = \[90] ,
  \V1243(0)  = \[91] ,
  \V1717(0)  = \[159] ,
  \V1243(3)  = \[88] ,
  \V985(0)  = V983 | (V978 | V984),
  \V1243(2)  = \[89] ,
  \V1243(5)  = \[86] ,
  \V1243(4)  = \[87] ,
  \V450(0)  = V448 | (V447 | V449),
  \V585(0)  = \[39] ,
  \V1255(1)  = V1252 | V1246,
  \V1255(0)  = V1254 | V1247,
  \V1255(3)  = V1248 | V1244,
  \V1255(2)  = V1250 | V1245,
  \V597(0)  = \[42] ,
  \V536(0)  = V534 | V535,
  \[200]  = V1941 | V1933,
  \[201]  = V1943 | V1934,
  \[202]  = V1945 | V1935,
  \[203]  = V1947 | V1936,
  \V1124(12)  = V1103 | V1093,
  \[204]  = V1949 | V1937,
  \V1124(13)  = V1101 | V1092,
  \[205]  = V1951 | V1938,
  \V813(0)  = \V807(0)  | V697,
  \[206]  = V1954 | V1940,
  \[207]  = V1957 | V1955,
  \V1679(0)  = \[152] ,
  \V413(0)  = \V174(0)  | (V502 | (V411 | \V404(0) )),
  \[208]  = V1959 | V1956,
  \[209]  = V1966 | V1967,
  \V1124(10)  = V1107 | V1095,
  \V1124(11)  = V1105 | V1094,
  \V1421(0)  = V1404 | (V1403 | V1418),
  \[210]  = V1989 | V1987,
  \[211]  = V1991 | V1988,
  \V2033(0)  = V2031 | (V2030 | V2032),
  \[212]  = V2293 | V2292,
  \[213]  = V2297 | V2296,
  \[214]  = V2301 | V2300,
  \[215]  = V2305 | V2304,
  \[216]  = V2309 | V2308,
  \V1833(0)  = \[184] ,
  \V1968(0)  = \[209] ,
  \[217]  = V2313 | V2312,
  \[218]  = V2317 | V2316,
  \[219]  = V2573 | V2572,
  \V1771(1)  = \[169] ,
  \V1771(0)  = \[170] ,
  \V640(0)  = \[49] ,
  \V375(0)  = \[4] ,
  \[220]  = V2577 | V2576,
  \[221]  = V2581 | V2580,
  \[222]  = V2585 | V2584,
  \[223]  = V2589 | V2588,
  \V1069(7)  = V1074 | V1058,
  \V1069(6)  = V1075 | V1059,
  \V1069(9)  = V1072 | V1056,
  \V1069(8)  = V1073 | V1057,
  \V1395(0)  = V700 | V701,
  \V603(0)  = \[43] ,
  \V1334(0)  = V1333 | V1332,
  \V1069(5)  = V1076 | V1060,
  \V1069(4)  = V1077 | V1061,
  \V1623(0)  = V1621 | V1622,
  \V1758(0)  = \[166] ,
  \V965(0)  = V962 | (V960 | (V961 | V963)),
  \V1900(0)  = \[191] ,
  \V504(0)  = V740 | V741,
  \V1709(1)  = \[157] ,
  \V1709(0)  = \[158] ,
  \V1709(3)  = \[155] ,
  \V1709(2)  = \[156] ,
  \V1709(4)  = \[154] ,
  \V1512(1)  = \[138] ,
  \V1647(0)  = V727 | (V769 | V726),
  \V1124(7)  = V1113 | V1098,
  \V1512(3)  = \[136] ,
  \V1124(6)  = V1115 | V1099,
  \V1512(2)  = \[137] ,
  \V1124(9)  = V1109 | V1096,
  \V1124(8)  = V1111 | V1097,
  \V380(0)  = V379 | V721,
  \V1124(3)  = V1402 | V1121,
  \V731(0)  = V723 | (V722 | V724),
  \V1124(2)  = V1402 | V1123,
  \V1124(5)  = V1117 | V1100,
  \V1597(0)  = ~V1594 | ~V1593,
  \V1124(4)  = V1402 | V1119,
  \V1536(0)  = \[139] ,
  \V405(0)  = V734 | (V515 | \V731(0) ),
  \V817(0)  = V696 | (\V214(0)  | (V815 | (V814 | (\V289(0)  | (\V302(0)  | V816))))),
  \V1351(0)  = V1350 | V1349,
  \V1086(1)  = V1083 | V1089,
  \V1086(0)  = V1090 | (V1085 | V1078),
  \V1086(3)  = V1079 | V1087,
  \V1086(2)  = V1081 | V1088,
  \V1898(0)  = \[189] ,
  \V1437(0)  = V1436 | ~\V278(0) ,
  \V982(0)  = V501 | (\V2011(0)  | V721),
  \V1652(0)  = \[149] ,
  \V1726(0)  = \[161] ,
  \V1399(0)  = V721 | V769,
  \V1953(7)  = \[200] ,
  \V1953(6)  = \[201] ,
  \V410(0)  = \[8] ,
  \V1953(1)  = \[199] ,
  \V1953(0)  = \[206] ,
  \V1953(3)  = \[204] ,
  \V1953(2)  = \[205] ,
  \V1553(0)  = \V60(0)  | \V63(0) ,
  \V1953(5)  = \[202] ,
  \V1953(4)  = \[203] ,
  \V1177(7)  = V1162 | V1150,
  \V1177(6)  = V1164 | V1151,
  \V1177(9)  = V1158 | V1148,
  \V1177(8)  = V1160 | V1149,
  \V508(0)  = \[13] ,
  \[10]  = ~V1570 & (~V1569 & (~V1568 & (~V1491 & (~V1646 & (~V1643 & (~V425 & (~\V1681(0)  & (~V1571 & (~V1572 & (~V392 & (~V1476 & (~\[165]  & (\[9]  & (~\V214(0)  & ~\V43(0) )))))))))))))),
  \[11]  = \[10]  | \[47] ,
  \V1977(0)  = V700 | V702,
  \[12]  = ~V499,
  \[13]  = V506 | (V613 | (V505 | V507)),
  \[14]  = \V40(0)  | V529,
  \[15]  = ~V530 & ~V509,
  \V1177(1)  = V1174 | V1156,
  \[16]  = ~V525 & (~V1646 & (~V695 & (~\V214(0)  & ~\V43(0) ))),
  \V1177(0)  = V1176 | V1157,
  \[17]  = V769 & \[81] ,
  \V1177(3)  = V1170 | V1154,
  \[18]  = V769 & \[80] ,
  \V1177(2)  = V1172 | V1155,
  \[19]  = V769 & \[79] ,
  \V1177(5)  = V1166 | V1152,
  \V1854(0)  = \V288(2)  | \V288(3) ,
  \V1177(4)  = V1168 | V1153,
  \V384(0)  = ~V351 | ~V350,
  \[20]  = V769 & \[78] ,
  \[21]  = V769 & \[77] ,
  \[22]  = V769 & \[76] ,
  \V1392(0)  = \[119] ,
  \[23]  = V769 & \[75] ,
  \V396(0)  = V395 | \[9] ,
  \[24]  = V769 & \[74] ,
  \[25]  = V769 & \[73] ,
  \V1331(0)  = V1330 | V1329,
  \[26]  = V769 & \[72] ,
  \V2078(0)  = V2077 | V2076,
  \[27]  = V769 & \[71] ,
  \[28]  = V769 & \[70] ,
  \[29]  = V553 | V573,
  \V612(0)  = V611 | V502,
  \V1829(7)  = \[175] ,
  \V1829(6)  = \[176] ,
  \V1829(9)  = \[173] ,
  \V1829(8)  = \[174] ,
  \[30]  = V555 | V574,
  \[31]  = V557 | V575,
  \V1417(0)  = V1416 | (V1406 | V745),
  \V1681(0)  = \V262(0)  | \V1674(0) ,
  \[32]  = V559 | V576,
  \[33]  = V561 | V577,
  \[34]  = V563 | V578,
  \V1281(0)  = \[105] ,
  \V1620(0)  = \[146] ,
  \[35]  = V579 | (V565 | V549),
  \V759(0)  = V747 | V748,
  \[36]  = V580 | (V567 | V550),
  \V1829(1)  = \[181] ,
  \[37]  = V581 | (V569 | V551),
  \V1829(0)  = \[182] ,
  \[38]  = V582 | (V571 | V552),
  \V1829(3)  = \[179] ,
  \[39]  = ~\V34(0) ,
  \V1829(2)  = \[180] ,
  \V1693(0)  = \[153] ,
  \V1829(5)  = \[177] ,
  \V1829(4)  = \[178] ,
  \V1632(0)  = V739 | (V741 | (V740 | V768)),
  \[40]  = ~V341 & ~\V243(0) ,
  \[41]  = V589 | V590,
  \[42]  = V594 | V596,
  \V1306(0)  = V1304 | (V1303 | V1305),
  \[43]  = V600 | V602,
  \[44]  = V606 | V608,
  \[45]  = ~V616 & (~V615 & ~V614),
  \[46]  = ~V531 & \V293(0) ,
  \[47]  = \V629(0)  & (~V623 & ~\V302(0) ),
  \[48]  = ~\V633(0) ,
  \[49]  = ~V638,
  \V1921(1)  = \[197] ,
  \V1921(0)  = \[198] ,
  \V1921(3)  = \[195] ,
  \V1921(2)  = \[196] ,
  \V1921(5)  = \[193] ,
  \[50]  = ~\V257(7) ,
  \V1921(4)  = \[194] ,
  \[51]  = V766 & ~\V149(3) ,
  \[52]  = ~V799 & (\V762(0)  & (~\V291(0)  & (~\V292(0)  & \V169(0) ))),
  \[53]  = ~\V807(0)  & (\V1674(0)  & (\[52]  & (\V14(0)  & \V70(0) ))),
  \[54]  = \V9(0)  & \V5(0) ,
  \[55]  = \V6(0)  & V372,
  \[56]  = \V6(0)  & \V9(0) ,
  \V802(0)  = \[65] ,
  \[57]  = \V6(0)  & (\V12(0)  & \V777(0) ),
  \[58]  = \V7(0)  & V372,
  \[59]  = \V11(0)  & \V5(0) ,
  \V1268(0)  = V721 | (V726 | (V400 | (V501 | (V769 | (V727 | V728))))),
  \V1471(0)  = V769 | (V766 | V701),
  \V1069(10)  = V1071 | V1055,
  \[60]  = \V11(0)  & \V7(0) ,
  \V1069(11)  = V1070 | V1054,
  \[61]  = \V9(0)  & \V7(0) ,
  \V414(0)  = \V1681(0)  | \V405(0) ,
  \[62]  = \V4(0)  & (\V788(0)  & \V9(0) ),
  \[63]  = ~V797,
  \[64]  = V799 & ~\V759(0) ,
  \[65]  = \V51(0)  | \V52(0) ,
  \[66]  = V818 | V820,
  \[67]  = V824 | (V823 | V825),
  \V487(0)  = V486 | V485,
  \[68]  = \V965(0)  & (~\V807(0)  & \V14(0) ),
  \V826(0)  = \[67] ,
  \[69]  = \V985(0)  & (~\V807(0)  & \V14(0) ),
  \V1422(0)  = V1407 | ~\V1417(0) ,
  \V1213(10)  = \[71] ,
  \V1213(11)  = \[70] ,
  \V1760(0)  = \[168] ,
  \V1360(0)  = V1359 | V1358,
  \V1495(0)  = \[135] ,
  \[70]  = V1190 | V1178,
  \[71]  = V1192 | V1179,
  \[72]  = V1194 | V1180,
  \[73]  = V1196 | V1181,
  \[74]  = V1198 | V1182,
  \[75]  = V1200 | V1183,
  \[76]  = V1202 | V1184,
  \[77]  = V1204 | V1185,
  \[78]  = V1206 | V1186,
  \V1711(0)  = V421 | V721,
  \[79]  = V1208 | V1187,
  \V376(0)  = V697 | \V35(0) ,
  \V1311(0)  = V1309 | (V1308 | V1310),
  \V2058(0)  = V2057 | V2056,
  \V788(0)  = ~V1564 | \V13(0) ,
  \[80]  = V1210 | V1188,
  \[81]  = V1212 | V1189,
  \[82]  = V1224 | V1214,
  \[83]  = V1226 | V1215,
  \[84]  = V1228 | V1216,
  \[85]  = V1230 | V1217,
  \V591(0)  = \[41] ,
  \[86]  = V1232 | V1218,
  \[87]  = V1234 | V1219,
  \[88]  = V1236 | V1220,
  \[89]  = V1238 | V1221,
  \V1396(0)  = \V60(0)  | \V59(0) ,
  \[90]  = V1240 | V1222,
  \V1409(0)  = V726 | (\V1395(0)  | V769),
  \[91]  = V1242 | V1223,
  \[92]  = V372 & \V2(0) ,
  \[93]  = ~V1558 & (~V1557 & (~V1555 & (\V2(0)  & (\V12(0)  & (~\V174(0)  & ~\V35(0) ))))),
  \[94]  = \V9(0)  & \V2(0) ,
  \[95]  = \V9(0)  & \V3(0) ,
  \[96]  = \V11(0)  & \V3(0) ,
  \[97]  = \[96]  & ~\V62(0) ,
  \[98]  = V372 & \V4(0) ,
  \[99]  = \V9(0)  & \V4(0) ,
  \V1759(0)  = \[167] ,
  \V1901(0)  = \[192] ,
  \V1297(1)  = \[109] ,
  \V1297(0)  = \[110] ,
  \V1297(3)  = \[107] ,
  \V1297(2)  = \[108] ,
  \V1297(4)  = \[106] ,
  \V1451(0)  = \[128] ,
  \V2002(0)  = V2001 | (V1996 | (V2000 | (\V1999(0)  | V1997))),
  \V1863(0)  = \[185] ,
  \V393(0)  = \[6] ,
  \V1463(0)  = V1461 | V1462,
  \V467(0)  = V466 | V465,
  \V1340(0)  = V1339 | V1338,
  \V1475(0)  = V1473 | V1474,
  \V2087(0)  = V2086 | V2085,
  \V2038(0)  = V2036 | (V2035 | V2037),
  \V1899(0)  = \[190] ,
  \V633(0)  = V631 | V632,
  \V1641(0)  = V1636 | (V1634 | (V1633 | (V1635 | V1637))),
  \V1653(0)  = V746 | (V743 | (V736 | (V735 | (V742 | (V744 | \V1687(0) ))))),
  V1000 = ~\V1395(0)  & (\V2011(0)  & \V189(5) ),
  V1002 = ~\V1395(0)  & (\V2011(0)  & \V189(4) ),
  V1004 = ~\V1395(0)  & (\V2011(0)  & \V189(3) ),
  V1006 = ~\V1395(0)  & (\V2011(0)  & \V189(2) ),
  V1008 = ~\V1395(0)  & (\V2011(0)  & \V189(1) ),
  V1010 = ~\V1395(0)  & (\V2011(0)  & \V189(0) ),
  V1012 = ~\V1395(0)  & (\V2011(0)  & \V183(5) ),
  V1014 = ~\V1395(0)  & (\V2011(0)  & \V183(4) ),
  V1016 = ~\V1395(0)  & (\V2011(0)  & \V183(3) ),
  V1018 = ~\V1395(0)  & (\V2011(0)  & \V183(2) ),
  V1020 = ~\V1395(0)  & (\V2011(0)  & \V183(1) ),
  V1022 = ~\V1395(0)  & (\V2011(0)  & \V183(0) ),
  V1024 = \V1395(0)  & (~\V2011(0)  & \V239(4) ),
  V1025 = \V1395(0)  & (~\V2011(0)  & \V239(3) ),
  V1026 = \V1395(0)  & (~\V2011(0)  & \V239(2) ),
  V1027 = \V1395(0)  & (~\V2011(0)  & \V239(1) ),
  V1028 = \V1395(0)  & (~\V2011(0)  & \V239(0) ),
  V1029 = \V1395(0)  & (~\V2011(0)  & \V234(4) ),
  V1030 = \V1395(0)  & (~\V2011(0)  & \V234(3) ),
  V1031 = \V1395(0)  & (~\V2011(0)  & \V234(2) ),
  V1032 = \V1395(0)  & (~\V2011(0)  & \V234(1) ),
  V1033 = \V1395(0)  & (~\V2011(0)  & \V234(0) ),
  V1034 = ~\V1395(0)  & (\V2011(0)  & \V199(4) ),
  V1036 = ~\V1395(0)  & (\V2011(0)  & \V199(3) ),
  V1038 = ~\V1395(0)  & (\V2011(0)  & \V199(2) ),
  \V1480(0)  = \[132] ,
  V1040 = ~\V1395(0)  & (\V2011(0)  & \V199(1) ),
  V1042 = ~\V1395(0)  & (\V2011(0)  & \V199(0) ),
  V1044 = ~\V1395(0)  & (\V2011(0)  & \V194(4) ),
  V1046 = ~\V1395(0)  & (\V2011(0)  & \V194(3) ),
  V1048 = ~\V1395(0)  & (\V2011(0)  & \V194(2) ),
  V1050 = ~\V1395(0)  & (\V2011(0)  & \V194(1) ),
  V1052 = ~\V1395(0)  & (\V2011(0)  & \V194(0) ),
  V1054 = ~\V1421(0)  & (V2115 & (\V1681(0)  & \V257(6) )),
  V1055 = ~\V1421(0)  & (V2115 & (\V1681(0)  & \V257(5) )),
  V1056 = ~\V1421(0)  & (V2115 & (\V1681(0)  & \V257(4) )),
  V1057 = ~\V1421(0)  & (V2115 & (\V1681(0)  & \V257(3) )),
  V1058 = ~\V1421(0)  & (V2115 & (\V1681(0)  & \V257(2) )),
  V1059 = ~\V1421(0)  & (V2115 & (\V1681(0)  & \V257(1) )),
  V1060 = ~\V1421(0)  & (V2115 & (\V1681(0)  & \V257(0) )),
  V1061 = ~\V1421(0)  & (V2115 & (\V1681(0)  & \V257(6) )),
  \V1554(0)  = V769 | (\V731(0)  | (V710 | (\V729(0)  | (V721 | \V730(0) )))),
  V1070 = \V1421(0)  & (V2116 & (\V1023(11)  & ~\V1681(0) )),
  V1071 = \V1421(0)  & (V2116 & (\V1023(10)  & ~\V1681(0) )),
  V1072 = \V1421(0)  & (V2116 & (\V1023(9)  & ~\V1681(0) )),
  V1073 = \V1421(0)  & (V2116 & (\V1023(8)  & ~\V1681(0) )),
  V1074 = \V1421(0)  & (V2116 & (\V1023(7)  & ~\V1681(0) )),
  V1075 = \V1421(0)  & (V2116 & (\V1023(6)  & ~\V1681(0) )),
  V1076 = \V1421(0)  & (V2116 & (\V1023(5)  & ~\V1681(0) )),
  V1077 = \V1421(0)  & (V2116 & (\V1023(4)  & ~\V1681(0) )),
  V1078 = V2119 & (~\V1421(0)  & (\V1681(0)  & \V257(7) )),
  V1079 = ~\V1421(0)  & (~V1445 & (V727 & (~\V1681(0)  & (\V149(7)  & ~\V59(0) )))),
  \V423(0)  = \[9] ,
  V1081 = ~\V1421(0)  & (~V1445 & (V727 & (~\V1681(0)  & (\V149(6)  & ~\V59(0) )))),
  V1083 = ~\V1421(0)  & (~V1445 & (V727 & (~\V1681(0)  & (\V149(5)  & ~\V59(0) )))),
  V1085 = ~\V1421(0)  & (~V1445 & (V727 & (~\V1681(0)  & (\V149(4)  & ~\V59(0) )))),
  V1087 = V2122 & (\V1421(0)  & (\V1053(3)  & ~\V1681(0) )),
  V1088 = V2122 & (\V1421(0)  & (\V1053(2)  & ~\V1681(0) )),
  V1089 = V2122 & (\V1421(0)  & (\V1053(1)  & ~\V1681(0) )),
  V1090 = V2122 & (\V1421(0)  & (\V1053(0)  & ~\V1681(0) )),
  V1092 = V1402 & \V32(8) ,
  V1093 = V1402 & \V32(7) ,
  V1094 = V1402 & \V32(6) ,
  V1095 = V1402 & \V32(5) ,
  V1096 = V1402 & \V32(4) ,
  V1097 = V1402 & \V32(3) ,
  V1098 = V1402 & \V32(2) ,
  V1099 = V1402 & \V32(1) ,
  \V1492(0)  = \[134] ,
  \V1831(0)  = V1830 | V1834,
  \V496(0)  = V495 | V494,
  V1100 = V1402 & \V32(0) ,
  V1101 = ~V1402 & \V32(11) ,
  V1103 = ~V1402 & \V32(10) ,
  V1105 = ~V1402 & \V32(9) ,
  V1107 = ~V1402 & \V32(8) ,
  V1109 = ~V1402 & \V32(7) ,
  \V435(0)  = \[11] ,
  V1111 = ~V1402 & \V32(6) ,
  V1113 = ~V1402 & \V32(5) ,
  V1115 = ~V1402 & \V32(4) ,
  V1117 = ~V1402 & \V32(3) ,
  V1119 = ~V1402 & \V32(2) ,
  V1121 = ~V1402 & \V32(1) ,
  V1123 = ~V1402 & \V32(0) ,
  V1125 = ~\V1681(0)  & \[52] ,
  V1127 = ~V1125 & \V1069(11) ,
  V1128 = ~V1125 & \V1069(10) ,
  V1129 = ~V1125 & \V1069(9) ,
  V1130 = ~V1125 & \V1069(8) ,
  V1131 = ~V1125 & \V1069(7) ,
  V1132 = ~V1125 & \V1069(6) ,
  V1133 = ~V1125 & \V1069(5) ,
  V1134 = V1125 & \V1124(6) ,
  V1136 = V1125 & \V1124(5) ,
  V1138 = V1125 & \V1124(4) ,
  V1140 = V1125 & \V1124(3) ,
  V1142 = V1125 & \V1124(2) ,
  V1144 = V1402 & V1125,
  V1146 = ~V1402 & V1125,
  V1148 = ~V1125 & (V2122 & (\V1421(0)  & (\V1053(9)  & ~\V1681(0) ))),
  V1149 = ~V1125 & (V2122 & (\V1421(0)  & (\V1053(8)  & ~\V1681(0) ))),
  V1150 = ~V1125 & (V2122 & (\V1421(0)  & (\V1053(7)  & ~\V1681(0) ))),
  V1151 = ~V1125 & (V2122 & (\V1421(0)  & (\V1053(6)  & ~\V1681(0) ))),
  V1152 = ~V1125 & (V2122 & (\V1421(0)  & (\V1053(5)  & ~\V1681(0) ))),
  V1153 = ~V1125 & (V2122 & (\V1421(0)  & (\V1053(4)  & ~\V1681(0) ))),
  V1154 = ~V1125 & \V1086(3) ,
  V1155 = ~V1125 & \V1086(2) ,
  V1156 = ~V1125 & \V1086(1) ,
  V1157 = ~V1125 & \V1086(0) ,
  V1158 = V1402 & (V1125 & \V32(11) ),
  V1160 = V1402 & (V1125 & \V32(10) ),
  V1162 = V1402 & (V1125 & \V32(9) ),
  V1164 = V1125 & \V1124(13) ,
  V1166 = V1125 & \V1124(12) ,
  V1168 = V1125 & \V1124(11) ,
  V1170 = V1125 & \V1124(10) ,
  V1172 = V1125 & \V1124(9) ,
  V1174 = V1125 & \V1124(8) ,
  V1176 = V1125 & \V1124(7) ,
  V1178 = ~\V1417(0)  & (\V1422(0)  & \V1147(11) ),
  V1179 = ~\V1417(0)  & (\V1422(0)  & \V1147(10) ),
  V1180 = ~\V1417(0)  & (\V1422(0)  & \V1147(9) ),
  V1181 = ~\V1417(0)  & (\V1422(0)  & \V1147(8) ),
  V1182 = ~\V1417(0)  & (\V1422(0)  & \V1147(7) ),
  V1183 = ~\V1417(0)  & (\V1422(0)  & \V1147(6) ),
  V1184 = ~\V1417(0)  & (\V1422(0)  & \V1147(5) ),
  V1185 = ~\V1417(0)  & (\V1422(0)  & (~V1125 & \V1069(4) )),
  V1186 = ~\V1417(0)  & (\V1422(0)  & (~V1125 & (\V1421(0)  & (V2116 & (\V1023(3)  & ~\V1681(0) ))))),
  V1187 = ~\V1417(0)  & (\V1422(0)  & (~V1125 & (\V1421(0)  & (V2116 & (\V1023(2)  & ~\V1681(0) ))))),
  V1188 = ~\V1417(0)  & (\V1422(0)  & (~V1125 & (\V1421(0)  & (V2116 & (\V1023(1)  & ~\V1681(0) ))))),
  V1189 = ~\V1417(0)  & (\V1422(0)  & (~V1125 & (\V1421(0)  & (V2116 & (\V1023(0)  & ~\V1681(0) ))))),
  V1190 = \V1417(0)  & (~\V1422(0)  & \V32(11) ),
  V1192 = \V1417(0)  & (~\V1422(0)  & \V32(10) ),
  V1194 = \V1417(0)  & (~\V1422(0)  & \V32(9) ),
  V1196 = \V1417(0)  & (~\V1422(0)  & \V32(8) ),
  V1198 = \V1417(0)  & (~\V1422(0)  & \V32(7) ),
  \V1781(1)  = \[171] ,
  \V1781(0)  = \[172] ,
  \V1855(0)  = \V288(4)  | \V288(5) ,
  \V385(0)  = ~V353 | ~V352,
  V1200 = \V1417(0)  & (~\V1422(0)  & \V32(6) ),
  V1202 = \V1417(0)  & (~\V1422(0)  & \V32(5) ),
  V1204 = \V1417(0)  & (~\V1422(0)  & \V32(4) ),
  V1206 = \V1417(0)  & (~\V1422(0)  & \V32(3) ),
  V1208 = \V1417(0)  & (~\V1422(0)  & \V32(2) ),
  V1210 = \V1417(0)  & (~\V1422(0)  & \V32(1) ),
  V1212 = \V1417(0)  & (~\V1422(0)  & \V32(0) ),
  V1214 = ~\V1417(0)  & (\V1422(0)  & \V1177(9) ),
  V1215 = ~\V1417(0)  & (\V1422(0)  & \V1177(8) ),
  V1216 = ~\V1417(0)  & (\V1422(0)  & \V1177(7) ),
  V1217 = ~\V1417(0)  & (\V1422(0)  & \V1177(6) ),
  V1218 = ~\V1417(0)  & (\V1422(0)  & \V1177(5) ),
  V1219 = ~\V1417(0)  & (\V1422(0)  & \V1177(4) ),
  \V1455(0)  = V1453 | V1454,
  V1220 = ~\V1417(0)  & (\V1422(0)  & \V1177(3) ),
  V1221 = ~\V1417(0)  & (\V1422(0)  & \V1177(2) ),
  V1222 = ~\V1417(0)  & (\V1422(0)  & \V1177(1) ),
  V1223 = ~\V1417(0)  & (\V1422(0)  & \V1177(0) ),
  V1224 = \V1417(0)  & (~\V1422(0)  & \V88(1) ),
  V1226 = \V1417(0)  & (~\V1422(0)  & \V88(0) ),
  V1228 = \V1417(0)  & (~\V1422(0)  & \V84(5) ),
  \V2067(0)  = V2066 | V2065,
  V1230 = \V1417(0)  & (~\V1422(0)  & \V84(4) ),
  V1232 = \V1417(0)  & (~\V1422(0)  & \V84(3) ),
  V1234 = \V1417(0)  & (~\V1422(0)  & \V84(2) ),
  V1236 = \V1417(0)  & (~\V1422(0)  & \V84(1) ),
  V1238 = \V1417(0)  & (~\V1422(0)  & \V84(0) ),
  V1240 = \V1417(0)  & (~\V1422(0)  & \V78(5) ),
  V1242 = \V1417(0)  & (~\V1422(0)  & \V78(4) ),
  V1244 = ~\V1417(0)  & (\V1422(0)  & (~V1125 & (\V1421(0)  & (V2116 & (\V1023(3)  & ~\V1681(0) ))))),
  V1245 = ~\V1417(0)  & (\V1422(0)  & (~V1125 & (\V1421(0)  & (V2116 & (\V1023(2)  & ~\V1681(0) ))))),
  V1246 = ~\V1417(0)  & (\V1422(0)  & (~V1125 & (\V1421(0)  & (V2116 & (\V1023(1)  & ~\V1681(0) ))))),
  V1247 = ~\V1417(0)  & (\V1422(0)  & (~V1125 & (\V1421(0)  & (V2116 & (\V1023(0)  & ~\V1681(0) ))))),
  V1248 = \V1417(0)  & (~\V1422(0)  & \V32(3) ),
  V1250 = \V1417(0)  & (~\V1422(0)  & \V32(2) ),
  V1252 = \V1417(0)  & (~\V1422(0)  & \V32(1) ),
  V1254 = \V1417(0)  & (~\V1422(0)  & \V32(0) ),
  V1256 = \[92] ,
  V1257 = \[93] ,
  V1258 = \[94] ,
  V1259 = \[95] ,
  V1260 = \[96] ,
  V1261 = \[97] ,
  V1262 = \[98] ,
  V1263 = \[99] ,
  V1264 = \[100] ,
  V1265 = \[101] ,
  V1266 = \[102] ,
  V1267 = \[103] ,
  V1272 = ~\V807(0)  & (V502 & (\V14(0)  & \V62(0) )),
  V1273 = ~\V1268(0)  & (~\V807(0)  & (~V768 & (~V767 & (~V749 & (~\[160]  & (\V14(0)  & \V59(0) )))))),
  V1276 = \V56(0)  & V735,
  V1279 = ~\V1984(0)  & (~V1276 & (\V213(0)  & \V14(0) )),
  V1280 = \V1546(0)  & \V1984(0) ,
  V1283 = ~V1979 & (~V1276 & (\V213(5)  & \V14(0) )),
  V1284 = ~V1979 & (~V1276 & (\V213(4)  & \V14(0) )),
  V1285 = ~V1979 & (~V1276 & (\V213(3)  & \V14(0) )),
  V1286 = ~V1979 & (~V1276 & (\V213(2)  & \V14(0) )),
  V1287 = ~V1979 & (~V1276 & (\V213(1)  & \V14(0) )),
  V1288 = V1979 & \V165(7) ,
  V1290 = V1979 & \V165(6) ,
  V1292 = V1979 & \V165(5) ,
  V1294 = V1979 & \V165(4) ,
  V1296 = V1979 & \V165(3) ,
  V1298 = V2513 | V2512,
  V1299 = V2025 & V1846,
  \V1467(0)  = \[130] ,
  \V336(0)  = V332 | (V323 | (V329 | V335)),
  \V2018(0)  = V2013 | (V2012 | V2014),
  V1300 = V2517 | V2516,
  V1301 = V2521 | V2520,
  V1302 = V2525 | V2524,
  V1303 = V1299 & V1848,
  V1304 = V1299 & V2029,
  V1305 = V1848 & V2029,
  V1307 = V2529 | V2528,
  V1308 = \V1306(0)  & V1839,
  V1309 = \V1306(0)  & V2034,
  V1310 = V1839 & V2034,
  V1312 = V2533 | V2532,
  V1316 = V2537 | V2536,
  V1317 = ~V1302 & ~V1298,
  V1318 = V2541 | V2540,
  V1319 = V1317 & ~V1307,
  V1320 = V2545 | V2544,
  V1324 = V2549 | V2548,
  V1325 = ~V1316 & V1298,
  V1326 = V2553 | V2552,
  V1327 = V1325 & ~V1318,
  V1328 = V2557 | V2556,
  V1329 = V1312 & V1848,
  V1330 = V1328 & ~V1848,
  V1332 = V1848 & V1307,
  V1333 = V1326 & ~V1848,
  V1335 = V1848 & V1302,
  V1336 = V1324 & ~V1848,
  V1338 = V1848 & V1298,
  V1339 = ~V1848 & V1298,
  V1344 = V2561 | V2560,
  V1345 = ~\V1340(0)  & ~\V1337(0) ,
  V1346 = V2565 | V2564,
  V1347 = V1345 & ~\V1334(0) ,
  V1348 = V2569 | V2568,
  V1349 = V1312 & V1846,
  V1350 = V1348 & ~V1846,
  V1352 = V1846 & V1307,
  V1353 = V1346 & ~V1846,
  V1355 = V1846 & V1302,
  V1356 = V1344 & ~V1846,
  V1358 = V1846 & V1298,
  V1359 = ~\V1340(0)  & ~V1846,
  V1365 = \[111] ,
  V1366 = \V268(4)  & (\V268(2)  & (\V268(1)  & (\V268(3)  & \V268(5) ))),
  V1367 = \V268(4)  & (\V268(2)  & (\V268(3)  & \V268(5) )),
  V1368 = \V268(4)  & (\V268(3)  & \V268(5) ),
  V1369 = \V268(4)  & \V268(5) ,
  V1370 = \[219] ,
  V1371 = \[220] ,
  V1372 = \[221] ,
  V1373 = \[222] ,
  V1374 = \[223] ,
  V1375 = \[112] ,
  V1378 = \[113] ,
  V1380 = \[114] ,
  V1382 = \[115] ,
  V1384 = \[116] ,
  V1386 = \[117] ,
  V1387 = \[118] ,
  V1390 = ~\V807(0)  & (~V401 & (~V741 & (\V14(0)  & \V65(0) ))),
  V1391 = ~\V807(0)  & (\[52]  & (\V14(0)  & (\V165(3)  & (\V165(6)  & (~\V165(5)  & (~\V165(4)  & \V70(0) )))))),
  V1393 = ~V1445 & V769,
  V1402 = \V1394(0)  & \[52] ,
  V1403 = V1445 & V727,
  V1404 = \V1396(0)  & (~V1445 & V727),
  V1406 = ~\V1415(0)  & (\V1398(0)  & \V1397(0) ),
  V1407 = \V1399(0)  & \V60(0) ,
  V1411 = V502 & \V56(0) ,
  V1412 = V502 & \V60(0) ,
  V1413 = V411 & \V56(0) ,
  V1414 = V411 & \V60(0) ,
  V1416 = ~V726 & (~V727 & (~\V1681(0)  & (\V53(0)  & ~\V56(0) ))),
  V1418 = \V1409(0)  & ~\V174(0) ,
  V1423 = \[120] ,
  V1425 = \V9(0)  & \V1(0) ,
  V1426 = \[121] ,
  V1427 = \V109(0)  & ~\V13(0) ,
  V1428 = \[122] ,
  V1429 = \[123] ,
  V1431 = \[124] ,
  V1432 = \[125] ,
  V1435 = ~V769 & (\V277(0)  & \V14(0) ),
  V1436 = V769 & \V277(0) ,
  V1438 = \V1437(0)  & \V14(0) ,
  V1443 = \V277(0)  & V769,
  V1445 = ~V1443 & \V278(0) ,
  V1448 = \V1447(0)  & (\V14(0)  & ~\V258(0) ),
  V1450 = ~\V1447(0)  & (\V14(0)  & \V258(0) ),
  V1453 = \V258(0)  & V1830,
  V1454 = V1836 & ~\V258(0) ,
  V1456 = \V1455(0)  & (~\V259(0)  & \V14(0) ),
  V1458 = ~\V1455(0)  & (\V259(0)  & \V14(0) ),
  V1461 = \V259(0)  & V1453,
  V1462 = V1454 & ~\V259(0) ,
  V1464 = \V1463(0)  & (~\V260(0)  & \V14(0) ),
  V1466 = ~\V1463(0)  & (\V260(0)  & \V14(0) ),
  V1470 = \[131] ,
  V1473 = \V1471(0)  & \[65] ,
  V1474 = \V1472(0)  & \V56(0) ,
  V1476 = \V1475(0)  & \V1597(0) ,
  V1478 = ~V701 & \[165] ,
  V1479 = V701 & (\[165]  & \[65] ),
  V1486 = ~\V69(0)  & (~\V68(0)  & (~\V70(0)  & ~\V66(0) )),
  V1490 = ~\V1999(0)  & (~V1486 & (\V14(0)  & \V215(0) )),
  V1491 = \V66(0)  & \V215(0) ,
  V1494 = \V216(0)  & ~\V214(0) ,
  V1497 = ~\V2002(0)  & (\V536(0)  & ~V345),
  \V1645(0)  = \[148] ,
  \V1983(0)  = V1981 | V1978,
  V1501 = ~\V2002(0)  & V345,
  V1503 = ~V1535 & ~\V2002(0) ,
  V1504 = ~V1535 & ~V1497,
  V1505 = ~V1535 & ~V1501,
  V1507 = V1535 & ~V360,
  V1509 = V1535 & ~V359,
  V1511 = V1535 & ~V358,
  V1513 = \V278(0)  & \V2011(0) ,
  V1516 = ~\V274(0)  & ~\V271(0) ,
  V1517 = \V172(0)  & \V56(0) ,
  V1518 = \V171(0)  & (\V1395(0)  & \V56(0) ),
  V1524 = ~V1518 & (~V1517 & (~V1513 & (\V177(0)  & ~\V248(0) ))),
  V1526 = V406 & ~\V172(0) ,
  V1527 = V515 & \V59(0) ,
  V1532 = ~V1527 & (~V1526 & (~V1524 & ~V1516)),
  V1535 = ~V1532 & (~\V2002(0)  & ~\V536(0) ),
  V1537 = \[140] ,
  V1539 = \[141] ,
  V1545 = ~\V165(3)  & (~\V165(7)  & (~\V165(6)  & (~\V165(5)  & ~\V165(4) ))),
  V1547 = ~V379 & (V721 & (~\[65]  & ~\V239(4) )),
  V1548 = V1986 & (~V379 & (V721 & ~\[65] )),
  V1549 = V379 & (V2157 & \[82] ),
  V1551 = V379 & (V2157 & \[83] ),
  V1555 = \V1554(0)  & \V57(0) ,
  V1557 = V739 & ~\V57(0) ,
  V1558 = V745 & \V1553(0) ,
  V1564 = \V71(0)  & \V202(0) ,
  V1568 = \[160]  & \V302(0) ,
  V1569 = V697 & \[160] ,
  V1570 = \[160]  & V698,
  V1571 = V1867 & (\[160]  & ~\V248(0) ),
  V1572 = V605 & (\[160]  & (\V247(0)  & ~\V248(0) )),
  V1579 = V2593 | V2592,
  V1580 = V2597 | V2596,
  V1581 = V2601 | V2600,
  V1582 = V2605 | V2604,
  V1583 = V2609 | V2608,
  V1584 = V2613 | V2612,
  V1585 = V2617 | V2616,
  V1586 = V2621 | V2620,
  V1587 = V2625 | V2624,
  V1588 = V2629 | V2628,
  V1589 = V2633 | V2632,
  V1590 = V2637 | V2636,
  V1591 = V2641 | V2640,
  V1592 = V2645 | V2644,
  V1593 = V2649 | V2648,
  V1594 = V2653 | V2652,
  V1598 = V2657 | V2656,
  V1599 = V2661 | V2660,
  \V2011(0)  = \V2007(0)  | V726,
  V1600 = V2665 | V2664,
  V1601 = V2669 | V2668,
  V1602 = V2673 | V2672,
  V1603 = V2677 | V2676,
  V1604 = V2681 | V2680,
  V1605 = V2685 | V2684,
  V1606 = V2689 | V2688,
  V1607 = V2693 | V2692,
  V1608 = V2697 | V2696,
  V1609 = V2701 | V2700,
  V1610 = V2705 | V2704,
  V1611 = V2709 | V2708,
  V1614 = \V292(0)  & ~\V302(0) ,
  V1615 = \V174(0)  & V695,
  V1616 = \V174(0)  & \V2002(0) ,
  V1621 = \V91(0)  & \V59(0) ,
  V1622 = \V91(1)  & \V62(0) ,
  V1624 = \V1623(0)  & V739,
  V1628 = ~V611 & (~V741 & ~\V294(0) ),
  \V1472(0)  = V744 | (V745 | V739),
  V1633 = \V1631(0)  & (\[65]  & ~\[52] ),
  V1634 = \[65]  & V701,
  V1635 = V737 & \V66(0) ,
  V1636 = \V1632(0)  & \V56(0) ,
  V1637 = \V66(0)  & \[52] ,
  V1638 = \V149(7)  & (V701 & \[65] ),
  V1639 = V766 & V687,
  V1640 = V701 & ~\V302(0) ,
  \V476(0)  = V475 | V474,
  V1643 = \V1641(0)  & \V336(0) ,
  V1644 = \V1642(0)  & (V1646 & (~V695 & (\V14(0)  & ~\V289(0) ))),
  V1646 = ~V1517 & \V207(0) ,
  \V2084(0)  = V2083 | V2082,
  V1648 = \V1647(0)  & V1445,
  V1651 = ~V1648 & (~\V1681(0)  & (\V295(0)  & (~\V290(0)  & (~\V249(0)  & ~\V289(0) )))),
  V1656 = ~\V1653(0)  & (~\V1687(0)  & (~V739 & (~V740 & ~V741))),
  V1660 = ~V1656 & (~\V812(0)  & (~\V2002(0)  & (~V696 & ~\V289(0) ))),
  V1662 = ~\V1653(0)  & (\[163]  & ~\V289(0) ),
  V1663 = V698 & (~\[65]  & ~\V289(0) ),
  \V1546(0)  = V1545 | V1646,
  V1664 = \V66(0)  & V737,
  V1669 = \[150] ,
  \V1023(7)  = V1008 | V992,
  V1672 = \V261(0)  & (~\V204(0)  & (\V165(3)  & (\V165(1)  & (\V165(7)  & (\V165(6)  & (\V165(5)  & (\V165(4)  & (\V165(2)  & \V165(0) )))))))),
  V1673 = \[52]  & (\V165(2)  & (\V165(1)  & (\V165(0)  & (\V165(6)  & (\V165(4)  & (\V165(3)  & (\V165(5)  & (\V261(0)  & (\V165(7)  & \V70(0) ))))))))),
  V1675 = ~\V260(0)  & (~\V259(0)  & (\V258(0)  & ~\V59(0) )),
  V1678 = ~V1675 & (\V262(0)  & \V14(0) ),
  \V1023(6)  = V1010 | V993,
  V1683 = \V1835(0)  & (~V1678 & \V262(0) ),
  V1686 = \V262(0)  & V1678,
  V1688 = \V56(0)  & V736,
  \V1023(9)  = V1004 | V990,
  V1691 = ~\V1983(0)  & (~V1688 & (\V100(0)  & \V14(0) )),
  V1692 = \V1983(0)  & \V1546(0) ,
  V1695 = ~V1978 & (~V1688 & (\V100(5)  & \V14(0) )),
  V1696 = ~V1978 & (~V1688 & (\V100(4)  & \V14(0) )),
  V1697 = ~V1978 & (~V1688 & (\V100(3)  & \V14(0) )),
  V1698 = ~V1978 & (~V1688 & (\V100(2)  & \V14(0) )),
  V1699 = ~V1978 & (~V1688 & (\V100(1)  & \V14(0) )),
  \V1023(8)  = V1006 | V991,
  \V1023(10)  = V1002 | V989,
  \V1023(11)  = V1000 | V988,
  V1700 = V1978 & \V165(7) ,
  V1702 = V1978 & \V165(6) ,
  V1704 = V1978 & \V165(5) ,
  V1706 = V1978 & \V165(4) ,
  V1708 = V1978 & \V165(3) ,
  \V1023(1)  = V1020 | V998,
  V1710 = V721 & ~\V280(0) ,
  V1712 = \V1711(0)  & \[65] ,
  V1716 = ~V1710 & (~\V807(0)  & (~V697 & (~V695 & (\V240(0)  & ~\V172(0) )))),
  V1719 = \[160] ,
  \V1023(0)  = V1022 | V999,
  V1721 = V1867 & \V194(0) ,
  V1723 = V1721 & (V1535 & \V2011(0) ),
  V1725 = ~\V2007(0)  & (\V242(0)  & \V14(0) ),
  \V1896(0)  = \[187] ,
  V1729 = \V1728(0)  & \V241(0) ,
  \V1023(3)  = V1016 | V996,
  V1730 = ~V768 & (~V738 & (V1646 & (~V687 & ~V701))),
  V1731 = V1646 & (V687 & (~V701 & \V59(0) )),
  V1732 = V768 & (V1646 & (~V701 & \V59(0) )),
  V1733 = V738 & (V1646 & (~V701 & \V62(0) )),
  V1735 = ~V1729 & ~V726,
  V1736 = \[162] ,
  V1738 = V1730 & ~V695,
  V1739 = V1731 & ~V695,
  \V1023(2)  = V1018 | V997,
  V1740 = V1732 & ~V695,
  V1744 = ~V747 & (~V725 & (\V33(0)  & \V289(0) )),
  V1748 = \V290(0)  & V695,
  V1749 = V751 & \V56(0) ,
  \V1023(5)  = V1012 | V994,
  V1750 = \V15(0)  & \V16(0) ,
  V1751 = \V15(0)  & ~\V16(0) ,
  V1752 = ~\V15(0)  & \V16(0) ,
  V1754 = V1752 & V700,
  V1755 = ~V1749 & (\V101(0)  & \V14(0) ),
  V1756 = V1752 & V725,
  \V1835(0)  = \V62(0)  | (\V56(0)  | \V50(0) ),
  \V1023(4)  = V1014 | V995,
  V1764 = V745 & ~\V88(3) ,
  V1765 = V745 & ~\V88(2) ,
  V1768 = ~V745 & ~\V134(1) ,
  V1770 = ~V745 & ~\V134(0) ,
  V1774 = ~V745 & ~\[70] ,
  V1775 = ~V745 & ~\[71] ,
  V1778 = V745 & ~\V78(3) ,
  V1780 = V745 & ~\V78(2) ,
  V1792 = ~\[82]  & \V37(0) ,
  V1793 = ~\[83]  & \V37(0) ,
  V1794 = ~\[84]  & \V37(0) ,
  V1795 = ~\[85]  & \V37(0) ,
  V1796 = ~\[86]  & \V37(0) ,
  V1797 = ~\[87]  & \V37(0) ,
  V1798 = ~\[88]  & \V37(0) ,
  V1799 = ~\[89]  & \V37(0) ,
  \V777(0)  = \V52(0)  | V776,
  V1800 = ~\[90]  & \V37(0) ,
  V1801 = ~\[79]  & \V37(0) ,
  \V1447(0)  = V1830 | V1836,
  V1810 = ~\[91]  & ~\V37(0) ,
  V1812 = ~\[70]  & ~\V37(0) ,
  V1814 = ~\[71]  & ~\V37(0) ,
  V1816 = ~\[72]  & ~\V37(0) ,
  V1818 = ~\[73]  & ~\V37(0) ,
  V1820 = ~\[74]  & ~\V37(0) ,
  V1822 = ~\[75]  & ~\V37(0) ,
  V1824 = ~\[76]  & ~\V37(0) ,
  V1826 = ~\[77]  & ~\V37(0) ,
  V1828 = ~\[91]  & ~\V37(0) ,
  V1830 = V1366 & \V268(0) ,
  V1832 = \[183] ,
  V1834 = ~V1683 & \V261(0) ,
  V1836 = \V1835(0)  & \V1681(0) ,
  V1838 = \V288(0)  & \V288(1) ,
  V1839 = \V288(2)  & \V288(3) ,
  V1840 = \V288(4)  & \V288(5) ,
  V1842 = \V288(5)  & ~\V288(4) ,
  V1844 = ~\V288(5)  & \V288(4) ,
  V1846 = \V288(3)  & ~\V288(2) ,
  V1848 = ~\V288(3)  & \V288(2) ,
  V1850 = \V288(1)  & ~\V288(0) ,
  V1852 = ~\V288(1)  & \V288(0) ,
  V1867 = \V199(3)  & (\V199(1)  & (\V194(4)  & (\V194(2)  & (\V194(1)  & (\V194(3)  & (\V199(0)  & (\V199(2)  & \V199(4) ))))))),
  V1868 = \V199(3)  & (\V199(1)  & (\V194(4)  & (\V194(2)  & (\V194(3)  & (\V199(0)  & (\V199(2)  & \V199(4) )))))),
  V1869 = \V199(3)  & (\V199(1)  & (\V194(4)  & (\V194(3)  & (\V199(0)  & (\V199(2)  & \V199(4) ))))),
  V1870 = \V199(3)  & (\V199(1)  & (\V194(4)  & (\V199(0)  & (\V199(2)  & \V199(4) )))),
  V1871 = \V199(3)  & (\V199(1)  & (\V199(0)  & (\V199(2)  & \V199(4) ))),
  V1872 = \V199(3)  & (\V199(1)  & (\V199(2)  & \V199(4) )),
  V1873 = \V199(3)  & (\V199(2)  & \V199(4) ),
  V1874 = \V199(3)  & \V199(4) ,
  V1875 = V2713 | V2712,
  V1876 = V2717 | V2716,
  V1877 = V2721 | V2720,
  V1878 = V2725 | V2724,
  V1879 = V2729 | V2728,
  V1880 = V2733 | V2732,
  V1881 = V2737 | V2736,
  V1882 = V2741 | V2740,
  V1883 = V2745 | V2744,
  V1885 = V1476 & V769,
  V1886 = V1995 & V725,
  V1887 = V1995 & V700,
  \[0]  = ~\[91] ,
  V1889 = ~V1902 & \V108(0) ,
  V1890 = ~V1902 & \V108(1) ,
  V1891 = ~V1902 & \V108(2) ,
  V1892 = ~V1902 & \V108(3) ,
  V1893 = ~V1902 & \V108(4) ,
  V1895 = ~V1749 & \V108(5) ,
  \[1]  = ~V954 & (~V952 & (~V936 & (~V916 & (~V896 & (~V876 & (~V856 & (~V836 & V347))))))),
  \V1459(0)  = \[129] ,
  \[2]  = ~V955 & (~V953 & (~V946 & (~V926 & (~V906 & (~V886 & (~V866 & (~V846 & ~\V1681(0) ))))))),
  \[3]  = \V10(0)  & \V13(0) ,
  \[4]  = \[120]  | (V1425 | (\[94]  | (\[124]  | (\[61]  | (\[54]  | (\[56]  | (\[118]  | (\[95]  | (\[99]  | \[62] ))))))))),
  \[5]  = \V376(0)  & \V203(0) ,
  \[6]  = V1571 | (V392 | V1572),
  \[7]  = ~V397,
  \V1397(0)  = V721 | (\V729(0)  | (V710 | (\V731(0)  | V1393))),
  V1902 = V750 & \V56(0) ,
  V1904 = ~V750 & (~V742 & (V736 & (~V735 & \V100(5) ))),
  V1905 = ~V750 & (~V742 & (V736 & (~V735 & \V100(4) ))),
  V1906 = ~V750 & (~V742 & (V736 & (~V735 & \V100(3) ))),
  V1907 = ~V750 & (~V742 & (V736 & (~V735 & \V100(2) ))),
  \V1213(7)  = \[74] ,
  V1908 = ~V750 & (~V742 & (V736 & (~V735 & \V100(1) ))),
  \[8]  = ~V409,
  V1909 = ~V750 & (~V742 & (V736 & (~V735 & \V100(0) ))),
  V1910 = ~V750 & (~V742 & (~V736 & (V735 & \V213(5) ))),
  V1912 = ~V750 & (~V742 & (~V736 & (V735 & \V213(4) ))),
  V1914 = ~V750 & (~V742 & (~V736 & (V735 & \V213(3) ))),
  V1916 = ~V750 & (~V742 & (~V736 & (V735 & \V213(2) ))),
  \V1213(6)  = \[75] ,
  V1918 = ~V750 & (~V742 & (~V736 & (V735 & \V213(1) ))),
  \[9]  = V420 | (V402 | (V417 | (V415 | (V416 | (V419 | (\[160]  | V422)))))),
  V1920 = ~V750 & (~V742 & (~V736 & (V735 & \V213(0) ))),
  V1922 = ~V750 & (V742 & (~V736 & (~V735 & \V124(5) ))),
  V1923 = ~V750 & (V742 & (~V736 & (~V735 & \V124(4) ))),
  V1924 = ~V750 & (V742 & (~V736 & (~V735 & \V124(3) ))),
  V1925 = ~V750 & (V742 & (~V736 & (~V735 & \V124(2) ))),
  V1926 = ~V750 & (V742 & (~V736 & (~V735 & \V124(1) ))),
  V1927 = ~V750 & (V742 & (~V736 & (~V735 & \V124(0) ))),
  \V1213(9)  = \[72] ,
  V1928 = V750 & (~V742 & (~V736 & (~V735 & \V108(4) ))),
  V1929 = V750 & (~V742 & (~V736 & (~V735 & \V108(3) ))),
  V1930 = V750 & (~V742 & (~V736 & (~V735 & \V108(2) ))),
  V1931 = V750 & (~V742 & (~V736 & (~V735 & \V108(1) ))),
  V1932 = V750 & (~V742 & (~V736 & (~V735 & \V108(0) ))),
  V1933 = ~V751 & (~V743 & (V742 & \V132(7) )),
  V1934 = ~V751 & (~V743 & (V742 & \V132(6) )),
  V1935 = ~V751 & (~V743 & (V742 & \V132(5) )),
  V1936 = ~V751 & (~V743 & (V742 & \V132(4) )),
  V1937 = ~V751 & (~V743 & (V742 & \V132(3) )),
  \V1213(8)  = \[73] ,
  V1938 = ~V751 & (~V743 & (V742 & \V132(2) )),
  V1940 = ~V751 & (~V743 & (V742 & \V132(0) )),
  V1941 = ~V751 & (V743 & (~V742 & \V118(5) )),
  V1943 = ~V751 & (V743 & (~V742 & \V118(4) )),
  V1945 = ~V751 & (V743 & (~V742 & \V118(3) )),
  V1947 = ~V751 & (V743 & (~V742 & \V118(2) )),
  V1949 = ~V751 & (V743 & (~V742 & \V118(1) )),
  V1951 = ~V751 & (V743 & (~V742 & \V118(0) )),
  V1954 = V751 & (~V743 & (~V742 & \V108(5) )),
  V1955 = V743 & (~\V382(0)  & \V118(7) ),
  V1956 = V743 & (~\V382(0)  & \V118(6) ),
  V1957 = ~V743 & (\V382(0)  & \V46(0) ),
  V1959 = ~V743 & (\V382(0)  & \V48(0) ),
  \V1674(0)  = V1672 | V1673,
  V1961 = V743 & \V56(0) ,
  V1962 = V1751 & (~\V108(4)  & \V101(0) ),
  V1966 = \V1963(0)  & (V700 & ~\V110(0) ),
  V1967 = ~V1962 & (~V1961 & (\V110(0)  & \V14(0) )),
  V1972 = ~\V288(7)  & ~\V288(6) ,
  V1973 = V2749 | V2748,
  V1974 = \V288(7)  & ~\V288(6) ,
  V1978 = \V290(0)  & (\V1977(0)  & V695),
  V1979 = V725 & (\V290(0)  & V695),
  \V1613(1)  = \[145] ,
  V1981 = \V1977(0)  & (~V1644 & (~V747 & (V1646 & ~V695))),
  V1982 = ~V1644 & (~V747 & (V725 & (V1646 & ~V695))),
  V1986 = V2753 | V2752,
  V1987 = ~V2009 & (V2188 & (V2006 & ~\V134(1) )),
  V1988 = ~V2009 & (V1994 & (V2188 & V2006)),
  \V1274(0)  = \[104] ,
  V1989 = ~V2009 & (V2189 & (~V2006 & \V134(1) )),
  \V1613(0)  = \[144] ,
  V1991 = ~V2009 & (V2189 & (~V2006 & \V134(0) )),
  V1994 = V2757 | V2756,
  V1995 = \V215(0)  & (\V172(0)  & \V67(0) ),
  V1996 = ~V1735 & (~V1445 & (~\[65]  & \V261(0) )),
  V1997 = ~V1735 & (V1445 & (~\[65]  & (\V272(0)  & (\V261(0)  & ~\V275(0) )))),
  \V1213(1)  = \[80] ,
  \V1213(0)  = \[81] ,
  \V1213(3)  = \[78] ,
  \V1213(2)  = \[79] ,
  \V1213(5)  = \[76] ,
  \V1213(4)  = \[77] ,
  \V629(0)  = \V270(0)  | (V626 | (V627 | V628)),
  \V1963(0)  = \[166]  | \V102(0) ,
  \V493(0)  = V492 | V491,
  \V1440(0)  = \[127] ,
  \V321(2)  = \[0] ,
  \V382(0)  = V740 | V741,
  \V2064(0)  = V2063 | V2062,
  \V1864(0)  = \[186] ,
  \V1999(0)  = V1732 | (V1730 | (V1995 | (\V214(0)  | (V1731 | V1733)))),
  \V807(0)  = \V2002(0)  | (V698 | (\V302(0)  | V696)),
  \V1538(0)  = \V69(0)  | \V50(0) ,
  \V1741(0)  = \[163] ,
  \V1415(0)  = V1413 | (V1411 | (V1412 | V1414)),
  \V572(3)  = \[35] ,
  \V572(2)  = \[36] ,
  \V634(0)  = \[48] ,
  \V572(5)  = \[33] ,
  \V572(4)  = \[34] ,
  \V1439(0)  = \[126] ,
  \V572(1)  = \[37] ,
  \V572(0)  = \[38] ,
  \V1642(0)  = V738 | (V1639 | (V768 | V1640)),
  \V511(0)  = \[14] ,
  \V572(7)  = \[31] ,
  \V572(6)  = \[32] ,
  \V572(9)  = \[29] ,
  \V572(8)  = \[30] ,
  \V1992(1)  = \[210] ,
  \V1728(0)  = V769 | V727,
  \V1992(0)  = \[211] ,
  \[100]  = \V12(0)  & \V4(0) ,
  \[101]  = \[100]  & \V52(0) ,
  \[102]  = \V11(0)  & \V4(0) ,
  \V609(0)  = \[44] ,
  \[103]  = \V11(0)  & \V2(0) ,
  \[104]  = V1273 | V1272,
  \V473(0)  = V472 | V471,
  \[105]  = V1280 | V1279,
  \V2081(0)  = V2080 | V2079,
  \V812(0)  = V811 | (V808 | V981),
  \[106]  = V1288 | V1283,
  \[107]  = V1290 | V1284,
  \V412(0)  = V721 | (\V729(0)  | (V710 | (\V1681(0)  | \V731(0) ))),
  \[108]  = V1292 | V1285,
  \[109]  = V1294 | V1286,
  V2000 = ~V2003 & (~V1445 & (\V2011(0)  & (~\[65]  & \V242(0) ))),
  V2001 = V1445 & (~\[65]  & (\V272(0)  & (\V134(0)  & (\V134(1)  & (\V242(0)  & ~\V275(0) ))))),
  V2003 = \V56(0)  & \V2007(0) ,
  V2005 = V1445 & ~\[65] ,
  V2006 = ~V745 & (~\V274(0)  & \V271(0) ),
  V2009 = \V2007(0)  & \[65] ,
  V2012 = ~V2023 & (~V2021 & (~V2005 & (~V1996 & \V2007(0) ))),
  V2013 = ~V2023 & (~V1996 & (~V1721 & (V726 & (~V1445 & ~\[65] )))),
  V2014 = V2006 & (~V1721 & (V1445 & (\V134(0)  & \V134(1) ))),
  V2015 = ~V1445 & (\V2011(0)  & ~\[65] ),
  V2021 = V1721 & ~\[65] ,
  V2023 = ~\[65]  & \V248(0) ,
  V2025 = V2761 | V2760,
  V2026 = ~V1974 & V1842,
  V2027 = V2765 | V2764,
  V2028 = V2769 | V2768,
  V2029 = V2773 | V2772,
  V2030 = V2026 & V1844,
  V2031 = V2026 & ~V1973,
  V2032 = ~V1973 & V1844,
  V2034 = V2777 | V2776,
  V2035 = \V2033(0)  & V1840,
  V2036 = \V2033(0)  & V1972,
  V2037 = V1840 & V1972,
  V2039 = V2781 | V2780,
  \V1481(0)  = \[133] ,
  V2043 = V2785 | V2784,
  V2044 = ~V2029 & ~V2025,
  V2045 = V2789 | V2788,
  V2046 = V2044 & ~V2034,
  V2047 = V2793 | V2792,
  V2051 = V2797 | V2796,
  V2052 = ~V2043 & V2025,
  V2053 = V2801 | V2800,
  V2054 = V2052 & ~V2045,
  V2055 = V2805 | V2804,
  V2056 = V2039 & V1844,
  V2057 = V2055 & ~V1844,
  V2059 = V1844 & V2034,
  V2060 = V2053 & ~V1844,
  V2062 = V1844 & V2029,
  V2063 = V2051 & ~V1844,
  V2065 = V1844 & V2025,
  V2066 = ~V1844 & V2025,
  \[110]  = V1296 | V1287,
  V2071 = V2809 | V2808,
  V2072 = ~\V2067(0)  & ~\V2064(0) ,
  V2073 = V2813 | V2812,
  V2074 = V2072 & ~\V2061(0) ,
  V2075 = V2817 | V2816,
  V2076 = V2039 & V1842,
  V2077 = V2075 & ~V1842,
  V2079 = V1842 & V2034,
  \V424(0)  = \[52]  | V687,
  \[111]  = ~\V807(0)  & (~V738 & (~V739 & (~\V1681(0)  & (~V734 & (~V515 & (~\V731(0)  & (~V740 & (\V14(0)  & \V62(0) )))))))),
  V2080 = V2073 & ~V1842,
  V2082 = V1842 & V2029,
  V2083 = V2071 & ~V1842,
  V2085 = V1842 & V2025,
  V2086 = ~\V2067(0)  & ~V1842,
  \[112]  = ~\V268(5) ,
  \[113]  = V2009 & (V372 & \V7(0) ),
  \V1629(0)  = \[147] ,
  \[114]  = \V2018(0)  & (V372 & \V7(0) ),
  \V762(0)  = V761 | (V700 | V725),
  \[115]  = \V380(0)  & (V372 & \V7(0) ),
  \[116]  = V372 & (V339 & \V7(0) ),
  \[117]  = V1836 & (V372 & \V7(0) ),
  \[118]  = \V8(0)  & \V9(0) ,
  \[119]  = V1390 | V1391,
  V2104 = ~\[65]  | ~V769,
  V2106 = ~\[65]  | ~V769,
  V2107 = ~\[65]  | ~V727,
  V2109 = ~\[65]  | ~V727,
  V2115 = V1445 | (~V727 | \V59(0) ),
  V2116 = V1445 | (~V727 | \V59(0) ),
  V2119 = V1445 | (~V727 | \V59(0) ),
  V2122 = V1445 | (~V727 | \V59(0) ),
  V2157 = ~V721 | \[65] ,
  \[120]  = \V9(0)  & \V1(0) ,
  \[121]  = V372 & \V1(0) ,
  V2188 = V2009 | V2006,
  V2189 = V2009 | ~V2006,
  \[122]  = \V1(0)  & \V11(0) ,
  \[123]  = \V1(0)  & \V12(0) ,
  \[124]  = ~V1427 & (\V9(0)  & \V1(0) ),
  \[125]  = ~\V807(0)  & (\V14(0)  & \V66(0) ),
  \[126]  = V1435 | V746,
  \[127]  = ~V1438,
  \[128]  = V1448 | V1450,
  \V1856(0)  = \V288(6)  | \V288(7) ,
  \V386(0)  = ~V355 | ~V354,
  \[129]  = V1456 | V1458,
  V2208 = V451 & ~\V32(0) ,
  V2209 = ~V451 & \V32(0) ,
  V2212 = V446 & ~\V32(1) ,
  V2213 = ~V446 & \V32(1) ,
  V2216 = V441 & ~\V32(2) ,
  V2217 = ~V441 & \V32(2) ,
  V2220 = ~V1298 & V1850,
  V2221 = V1298 & ~V1850,
  V2224 = ~V1302 & V1852,
  V2225 = V1302 & ~V1852,
  V2228 = ~V1307 & V1838,
  V2229 = V1307 & ~V1838,
  V2232 = V439 & ~V438,
  V2233 = ~V439 & V438,
  V2236 = ~V440 & \V445(0) ,
  V2237 = V440 & ~\V445(0) ,
  V2240 = V1312 & ~\V450(0) ,
  V2241 = ~V1312 & \V450(0) ,
  V2244 = V437 & V441,
  V2245 = ~V437 & ~V441,
  V2248 = ~V453 & V446,
  V2249 = V453 & ~V446,
  V2252 = ~V455 & V451,
  V2253 = V455 & ~V451,
  V2256 = V452 & ~V437,
  V2257 = ~V452 & V437,
  \V2007(0)  = V769 | V727,
  \V798(0)  = \[63] ,
  V2260 = ~V461 & V454,
  V2261 = V461 & ~V454,
  V2264 = V456 & ~V463,
  V2265 = ~V456 & V463,
  V2268 = \V476(0)  & \V473(0) ,
  V2269 = ~\V476(0)  & ~\V473(0) ,
  \[130]  = V1464 | V1466,
  V2272 = ~V481 & \V470(0) ,
  V2273 = V481 & ~\V470(0) ,
  V2276 = ~V483 & \V467(0) ,
  V2277 = V483 & ~\V467(0) ,
  \V1394(0)  = \V60(0)  | (\V56(0)  | \V59(0) ),
  \[131]  = ~\V807(0)  & (~V737 & (\V67(0)  & \V14(0) )),
  V2280 = ~\V38(0)  & \V39(0) ,
  V2281 = \V38(0)  & ~\V39(0) ,
  V2284 = ~\V44(0)  & \V42(0) ,
  V2285 = \V44(0)  & ~\V42(0) ,
  \V398(0)  = \[7] ,
  V2288 = \V41(0)  & ~\V45(0) ,
  V2289 = ~\V41(0)  & \V45(0) ,
  \[132]  = V1478 | (V1476 | V1479),
  V2292 = ~V644 & \V257(0) ,
  V2293 = V644 & ~\V257(0) ,
  V2296 = ~V645 & \V257(1) ,
  V2297 = V645 & ~\V257(1) ,
  \[133]  = ~\V214(0) ,
  \[134]  = V1490 | V1494,
  \[135]  = ~\V175(0) ,
  \[136]  = V1507 | V1503,
  \V1671(0)  = \[151] ,
  \[137]  = V1509 | V1504,
  \V2019(0)  = V2014 | V2015,
  \[138]  = V1511 | V1505,
  \[139]  = ~V1535,
  V2300 = ~V646 & \V257(2) ,
  V2301 = V646 & ~\V257(2) ,
  V2304 = ~V647 & \V257(3) ,
  V2305 = V647 & ~\V257(3) ,
  V2308 = ~V648 & \V257(4) ,
  V2309 = V648 & ~\V257(4) ,
  \V1745(0)  = \[164] ,
  V2312 = ~V649 & \V257(5) ,
  V2313 = V649 & ~\V257(5) ,
  V2316 = \V257(6)  & ~\V257(7) ,
  V2317 = ~\V257(6)  & \V257(7) ,
  V2320 = \V2078(0)  & ~\V1255(0) ,
  V2321 = ~\V2078(0)  & \V1255(0) ,
  V2324 = \V2081(0)  & ~\V1255(1) ,
  V2325 = ~\V2081(0)  & \V1255(1) ,
  V2328 = \V2084(0)  & ~\V1255(2) ,
  V2329 = ~\V2084(0)  & \V1255(2) ,
  V2332 = \V2087(0)  & ~\V1255(3) ,
  V2333 = ~\V2087(0)  & \V1255(3) ,
  V2336 = \V2058(0)  & ~\V1255(0) ,
  V2337 = ~\V2058(0)  & \V1255(0) ,
  V2340 = \V2061(0)  & ~\V1255(1) ,
  V2341 = ~\V2061(0)  & \V1255(1) ,
  V2344 = \V2064(0)  & ~\V1255(2) ,
  V2345 = ~\V2064(0)  & \V1255(2) ,
  V2348 = \V2067(0)  & ~\V1255(3) ,
  V2349 = ~\V2067(0)  & \V1255(3) ,
  V2352 = V2047 & ~\V1255(0) ,
  V2353 = ~V2047 & \V1255(0) ,
  V2356 = V2045 & ~\V1255(1) ,
  V2357 = ~V2045 & \V1255(1) ,
  V2360 = V2043 & ~\V1255(2) ,
  V2361 = ~V2043 & \V1255(2) ,
  V2364 = ~V2025 & ~\V1255(3) ,
  V2365 = V2025 & \V1255(3) ,
  V2368 = V2039 & ~\V1255(0) ,
  V2369 = ~V2039 & \V1255(0) ,
  \[140]  = ~\V807(0)  & (\V68(0)  & \V14(0) ),
  V2372 = V2034 & ~\V1255(1) ,
  V2373 = ~V2034 & \V1255(1) ,
  V2376 = V2029 & ~\V1255(2) ,
  V2377 = ~V2029 & \V1255(2) ,
  \[141]  = \V1538(0)  & (~\V807(0)  & \V14(0) ),
  V2380 = V2025 & ~\V1255(3) ,
  V2381 = ~V2025 & \V1255(3) ,
  V2384 = \V1351(0)  & ~\V1255(0) ,
  V2385 = ~\V1351(0)  & \V1255(0) ,
  V2388 = \V1354(0)  & ~\V1255(1) ,
  V2389 = ~\V1354(0)  & \V1255(1) ,
  \[142]  = V1549 | V1547,
  V2392 = \V1357(0)  & ~\V1255(2) ,
  V2393 = ~\V1357(0)  & \V1255(2) ,
  V2396 = \V1360(0)  & ~\V1255(3) ,
  V2397 = ~\V1360(0)  & \V1255(3) ,
  \V1757(0)  = \[165] ,
  \[143]  = V1551 | V1548,
  \[144]  = ~V1610,
  \[145]  = ~V1611,
  \V1960(1)  = \[207] ,
  \V1357(0)  = V1356 | V1355,
  \[146]  = V1616 | (V1614 | (V1615 | V799)),
  \V1960(0)  = \[208] ,
  \V490(0)  = V489 | V488,
  \[147]  = V1628 | (V1624 | V531),
  \[148]  = V1643 | (V1644 | V1638),
  \[149]  = ~V1651,
  V2400 = \V1331(0)  & ~\V1255(0) ,
  V2401 = ~\V1331(0)  & \V1255(0) ,
  V2404 = \V1334(0)  & ~\V1255(1) ,
  V2405 = ~\V1334(0)  & \V1255(1) ,
  V2408 = \V1337(0)  & ~\V1255(2) ,
  V2409 = ~\V1337(0)  & \V1255(2) ,
  V2412 = \V1340(0)  & ~\V1255(3) ,
  V2413 = ~\V1340(0)  & \V1255(3) ,
  V2416 = V1320 & ~\V1255(0) ,
  V2417 = ~V1320 & \V1255(0) ,
  V2420 = V1318 & ~\V1255(1) ,
  V2421 = ~V1318 & \V1255(1) ,
  V2424 = V1316 & ~\V1255(2) ,
  V2425 = ~V1316 & \V1255(2) ,
  V2428 = ~\V1255(3)  & ~V1298,
  V2429 = \V1255(3)  & V1298,
  V2432 = V1312 & ~\V1255(0) ,
  V2433 = ~V1312 & \V1255(0) ,
  V2436 = ~\V1255(1)  & V1307,
  \V503(0)  = V727 | (V721 | (V501 | (V769 | V611))),
  V2437 = \V1255(1)  & ~V1307,
  V2440 = ~\V1255(2)  & V1302,
  V2441 = \V1255(2)  & ~V1302,
  V2444 = ~\V1255(3)  & V1298,
  V2445 = \V1255(3)  & ~V1298,
  V2448 = ~\V1255(0)  & \V487(0) ,
  V2449 = \V1255(0)  & ~\V487(0) ,
  V2452 = ~\V1255(1)  & \V490(0) ,
  V2453 = \V1255(1)  & ~\V490(0) ,
  V2456 = ~\V1255(2)  & \V493(0) ,
  V2457 = \V1255(2)  & ~\V493(0) ,
  V2460 = ~\V1255(3)  & \V496(0) ,
  V2461 = \V1255(3)  & ~\V496(0) ,
  V2464 = ~\V1255(0)  & \V467(0) ,
  V2465 = \V1255(0)  & ~\V467(0) ,
  V2468 = ~\V1255(1)  & \V470(0) ,
  V2469 = \V1255(1)  & ~\V470(0) ,
  \[150]  = ~V1664 & (~V1663 & (~V1662 & ~V1660)),
  V2472 = ~\V1255(2)  & \V473(0) ,
  V2473 = \V1255(2)  & ~\V473(0) ,
  V2476 = ~\V1255(3)  & \V476(0) ,
  V2477 = \V1255(3)  & ~\V476(0) ,
  \[151]  = ~\V205(0) ,
  V2480 = V456 & ~\V1255(0) ,
  V2481 = ~V456 & \V1255(0) ,
  V2484 = ~\V1255(1)  & V454,
  V2485 = \V1255(1)  & ~V454,
  V2488 = ~\V1255(2)  & V452,
  V2489 = \V1255(2)  & ~V452,
  \[152]  = \V1674(0)  | V1678,
  V2492 = ~\V1255(3)  & ~V437,
  V2493 = \V1255(3)  & V437,
  V2496 = ~\V1255(0)  & V451,
  V2497 = \V1255(0)  & ~V451,
  \[153]  = V1692 | V1691,
  \[154]  = V1700 | V1695,
  \[155]  = V1702 | V1696,
  \[156]  = V1704 | V1697,
  \[157]  = V1706 | V1698,
  \V1984(0)  = V1979 | V1982,
  \[158]  = V1708 | V1699,
  \[159]  = V1712 | V1716,
  V2500 = ~\V1255(1)  & V446,
  V2501 = \V1255(1)  & ~V446,
  V2504 = ~\V1255(2)  & V441,
  V2505 = \V1255(2)  & ~V441,
  V2508 = ~\V1255(3)  & V437,
  V2509 = \V1255(3)  & ~V437,
  V2512 = ~V2025 & V1846,
  V2513 = V2025 & ~V1846,
  V2516 = ~V2029 & V1848,
  V2517 = V2029 & ~V1848,
  V2520 = ~V2034 & V1839,
  V2521 = V2034 & ~V1839,
  V2524 = V1300 & ~V1299,
  V2525 = ~V1300 & V1299,
  V2528 = ~V1301 & \V1306(0) ,
  \V2061(0)  = V2060 | V2059,
  V2529 = V1301 & ~\V1306(0) ,
  V2532 = V2039 & ~\V1311(0) ,
  V2533 = ~V2039 & \V1311(0) ,
  V2536 = V1302 & V1298,
  V2537 = ~V1302 & ~V1298,
  V2540 = ~V1317 & V1307,
  V2541 = V1317 & ~V1307,
  V2544 = V1312 & ~V1319,
  V2545 = ~V1312 & V1319,
  V2548 = V1316 & ~V1298,
  V2549 = ~V1316 & V1298,
  V2552 = ~V1325 & V1318,
  V2553 = V1325 & ~V1318,
  V2556 = V1320 & ~V1327,
  V2557 = ~V1320 & V1327,
  V2560 = \V1340(0)  & \V1337(0) ,
  V2561 = ~\V1340(0)  & ~\V1337(0) ,
  V2564 = ~V1345 & \V1334(0) ,
  V2565 = V1345 & ~\V1334(0) ,
  V2568 = ~V1347 & \V1331(0) ,
  V2569 = V1347 & ~\V1331(0) ,
  \[160]  = ~V695 & (\V240(0)  & ~\V172(0) ),
  V2572 = ~V1366 & \V268(0) ,
  V2573 = V1366 & ~\V268(0) ,
  V2576 = ~V1367 & \V268(1) ,
  V2577 = V1367 & ~\V268(1) ,
  \[161]  = V1723 | V1725,
  V2580 = ~V1368 & \V268(2) ,
  V2581 = V1368 & ~\V268(2) ,
  \V391(0)  = V389 | (V387 | (V388 | V390)),
  V2584 = ~V1369 & \V268(3) ,
  V2585 = V1369 & ~\V268(3) ,
  \V730(0)  = V719 | V720,
  V2588 = \V268(4)  & ~\V268(5) ,
  V2589 = ~\V268(4)  & \V268(5) ,
  \[162]  = V1735 & (V698 & (~\[65]  & (~\V290(0)  & ~\V289(0) ))),
  V2592 = ~\V78(0)  & \V78(1) ,
  V2593 = \V78(0)  & ~\V78(1) ,
  V2596 = \V78(3)  & ~\V78(2) ,
  V2597 = ~\V78(3)  & \V78(2) ,
  \[163]  = V1740 | (V1738 | (V1748 | (V1739 | V1733))),
  \[164]  = ~V1744,
  \[165]  = V1750 | V1751,
  \[166]  = V1751 | V1752,
  \V1147(7)  = V1142 | V1131,
  \[167]  = V1755 | (V1754 | V1756),
  \V404(0)  = V400 | V728,
  \V1147(6)  = V1144 | V1132,
  \[168]  = ~\V101(0) ,
  \V1147(9)  = V1138 | V1129,
  \[169]  = V1768 | V1764,
  V2600 = ~\V78(4)  & \V78(5) ,
  V2601 = \V78(4)  & ~\V78(5) ,
  V2604 = ~\V84(0)  & \V84(1) ,
  V2605 = \V84(0)  & ~\V84(1) ,
  V2608 = ~\V84(2)  & \V84(3) ,
  V2609 = \V84(2)  & ~\V84(3) ,
  \V1147(8)  = V1140 | V1130,
  V2612 = ~\V84(4)  & \V84(5) ,
  V2613 = \V84(4)  & ~\V84(5) ,
  V2616 = ~\V88(0)  & \V88(1) ,
  V2617 = \V88(0)  & ~\V88(1) ,
  V2620 = \V88(3)  & ~\V88(2) ,
  V2621 = ~\V88(3)  & \V88(2) ,
  V2624 = V1580 & ~V1579,
  V2625 = ~V1580 & V1579,
  V2628 = V1582 & ~V1581,
  V2629 = ~V1582 & V1581,
  V2632 = V1584 & ~V1583,
  V2633 = ~V1584 & V1583,
  V2636 = V1586 & ~V1585,
  V2637 = ~V1586 & V1585,
  V2640 = V1588 & ~V1587,
  V2641 = ~V1588 & V1587,
  V323 = ~V451 & \V32(0) ,
  V2644 = V1590 & ~V1589,
  V324 = V2209 | V2208,
  V2645 = ~V1590 & V1589,
  V325 = V2213 | V2212,
  V326 = V2217 | V2216,
  V2648 = ~V1591 & \V94(0) ,
  V2649 = V1591 & ~\V94(0) ,
  V329 = ~V324 & (~V446 & \V32(1) ),
  V2652 = ~V1592 & \V94(1) ,
  V332 = ~V325 & (~V441 & (~V324 & \V32(2) )),
  V2653 = V1592 & ~\V94(1) ,
  V335 = ~V326 & (~V437 & (~V325 & (~V324 & \V32(3) ))),
  V2656 = ~\[198]  & \[197] ,
  V2657 = \[198]  & ~\[197] ,
  V339 = V744 & (~V695 & (~V1476 & \V56(0) )),
  V2660 = ~\[196]  & \[195] ,
  V340 = V721 & \[65] ,
  V2661 = \[196]  & ~\[195] ,
  V341 = \[65]  & \V2011(0) ,
  V2664 = ~\[194]  & \[193] ,
  V2665 = \[194]  & ~\[193] ,
  V345 = \V759(0)  & \V56(0) ,
  V347 = ~V433 & ~\V1681(0) ,
  V2668 = ~\[206]  & \[199] ,
  V348 = ~V946 & (~V936 & ~\V1681(0) ),
  V2669 = \[206]  & ~\[199] ,
  V349 = ~V926 & (~V916 & ~\V1681(0) ),
  \[170]  = V1770 | V1765,
  V350 = ~V906 & (~V896 & ~\V1681(0) ),
  V351 = ~V886 & (~V876 & ~\V1681(0) ),
  V2672 = ~\[205]  & \[204] ,
  V352 = ~V866 & (~V856 & ~\V1681(0) ),
  V2673 = \[205]  & ~\[204] ,
  V353 = ~V846 & (~V836 & ~\V1681(0) ),
  V354 = ~V955 & (~V954 & ~\V1681(0) ),
  V355 = ~V953 & (~V952 & ~\V1681(0) ),
  V2676 = ~\[203]  & \[202] ,
  V356 = \[1] ,
  V2677 = \[203]  & ~\[202] ,
  V357 = \[2] ,
  V358 = ~V946 & (~V936 & (~V926 & (~V916 & (~V906 & (~V896 & (~V886 & ~V876)))))),
  V359 = ~V946 & (~V936 & (~V926 & (~V916 & (~V866 & (~V856 & (~V846 & ~V836)))))),
  \[171]  = V1778 | V1774,
  V2680 = ~\[201]  & \[200] ,
  V360 = ~V955 & (~V954 & (~V946 & (~V936 & (~V906 & (~V896 & (~V866 & ~V856)))))),
  V2681 = \[201]  & ~\[200] ,
  V2684 = ~\[208]  & \[207] ,
  V2685 = \[208]  & ~\[207] ,
  V2688 = V1599 & ~V1598,
  V2689 = ~V1599 & V1598,
  \[172]  = V1780 | V1775,
  V2692 = V1601 & ~V1600,
  V372 = ~\V13(0)  & \V10(0) ,
  V2693 = ~V1601 & V1600,
  V373 = \[3] ,
  V2696 = V1603 & ~V1602,
  V2697 = ~V1603 & V1602,
  V377 = \[5] ,
  V379 = \V378(0)  & \[65] ,
  \[173]  = V1810 | V1792,
  V387 = V1838 & \V383(0) ,
  V388 = V1839 & \V384(0) ,
  V389 = V1840 & \V385(0) ,
  \[174]  = V1812 | V1793,
  V390 = \V288(7)  & (\V288(6)  & \V386(0) ),
  V392 = \V391(0)  & (\[160]  & (\[84]  & (\[83]  & (\[82]  & ~\V248(0) )))),
  V395 = \V248(0)  & \[160] ,
  V397 = ~V1570 & (~V1569 & (~V1568 & (~V425 & (\V396(0)  & (~V1571 & (~V1572 & (~V392 & (~\V214(0)  & ~\V43(0) )))))))),
  \V1147(5)  = V1146 | V1133,
  \[175]  = V1814 | V1794,
  \[176]  = V1816 | V1795,
  \[177]  = V1818 | V1796,
  \[178]  = V1820 | V1797,
  \[179]  = V1822 | V1798,
  V2700 = V1605 & ~V1604,
  V2701 = ~V1605 & V1604,
  V2704 = V1607 & ~V1606,
  V2705 = ~V1607 & V1606,
  V2708 = V1609 & ~V1608,
  V2709 = ~V1609 & V1608,
  V2712 = ~V1867 & \V194(0) ,
  V2713 = V1867 & ~\V194(0) ,
  V2716 = ~V1868 & \V194(1) ,
  V2717 = V1868 & ~\V194(1) ,
  V2720 = ~V1869 & \V194(2) ,
  V400 = ~V687 & \V730(0) ,
  V2721 = V1869 & ~\V194(2) ,
  V401 = \V729(0)  & V687,
  V402 = V401 & \V62(0) ,
  V2724 = ~V1870 & \V194(3) ,
  V2725 = V1870 & ~\V194(3) ,
  V406 = \V404(0)  & \V56(0) ,
  \V1897(0)  = \[188] ,
  V407 = \V405(0)  & \V59(0) ,
  V2728 = ~V1871 & \V194(4) ,
  V2729 = V1871 & ~\V194(4) ,
  V409 = \V408(0)  & (~V695 & ~\[165] ),
  V411 = V687 & \V729(0) ,
  V2732 = ~V1872 & \V199(0) ,
  V2733 = V1872 & ~\V199(0) ,
  V415 = \V412(0)  & \[65] ,
  V2736 = ~V1873 & \V199(1) ,
  V416 = \V413(0)  & \V56(0) ,
  V2737 = V1873 & ~\V199(1) ,
  V417 = \V414(0)  & \V59(0) ,
  V419 = ~V695 & (\[52]  & (\V66(0)  & ~\V215(0) )),
  V2740 = ~V1874 & \V199(2) ,
  V420 = \V1681(0)  & \V70(0) ,
  V2741 = V1874 & ~\V199(2) ,
  V421 = ~V1445 & \V2011(0) ,
  V422 = V421 & \[65] ,
  V2744 = \V199(3)  & ~\V199(4) ,
  V2745 = ~\V199(3)  & \V199(4) ,
  V425 = \V424(0)  & \[65] ,
  V2748 = \V288(7)  & ~\V288(6) ,
  V2749 = ~\V288(7)  & \V288(6) ,
  V2752 = ~\V239(3)  & \V239(4) ,
  V432 = \[10] ,
  V2753 = \V239(3)  & ~\V239(4) ,
  V433 = V749 & ~\[65] ,
  V2756 = ~\V134(0)  & \V134(1) ,
  V2757 = \V134(0)  & ~\V134(1) ,
  V437 = V2221 | V2220,
  V438 = V1298 & V1850,
  V439 = V2225 | V2224,
  V2760 = V1974 & V1842,
  V440 = V2229 | V2228,
  V2761 = ~V1974 & ~V1842,
  V441 = V2233 | V2232,
  V442 = V438 & V1852,
  V443 = V438 & V1302,
  V2764 = V1973 & V1844,
  V444 = V1852 & V1302,
  V2765 = ~V1973 & ~V1844,
  V446 = V2237 | V2236,
  V447 = \V445(0)  & V1838,
  V2768 = ~V1972 & V1840,
  V448 = \V445(0)  & V1307,
  V2769 = V1972 & ~V1840,
  V449 = V1838 & V1307,
  \[180]  = V1824 | V1799,
  V451 = V2241 | V2240,
  V2772 = V2027 & ~V2026,
  V452 = V2245 | V2244,
  V2773 = ~V2027 & V2026,
  V453 = ~V437 & ~V441,
  V454 = V2249 | V2248,
  V455 = V453 & ~V446,
  V2776 = ~V2028 & \V2033(0) ,
  V456 = V2253 | V2252,
  V2777 = V2028 & ~\V2033(0) ,
  \[181]  = V1826 | V1800,
  V2780 = ~\V2038(0)  & V1972,
  V460 = V2257 | V2256,
  V2781 = \V2038(0)  & ~V1972,
  V461 = ~V452 & V437,
  V462 = V2261 | V2260,
  V463 = V461 & ~V454,
  V2784 = V2029 & V2025,
  V464 = V2265 | V2264,
  V2785 = ~V2029 & ~V2025,
  V465 = V1852 & V451,
  V466 = V464 & ~V1852,
  V2788 = ~V2044 & V2034,
  V468 = V1852 & V446,
  V2789 = V2044 & ~V2034,
  V469 = V462 & ~V1852,
  \[182]  = V1828 | V1801,
  V471 = V1852 & V441,
  V2792 = V2039 & ~V2046,
  V472 = V460 & ~V1852,
  V2793 = ~V2039 & V2046,
  V474 = V1852 & V437,
  V475 = ~V1852 & V437,
  V2796 = V2043 & ~V2025,
  V2797 = ~V2043 & V2025,
  \[183]  = \V1831(0)  & \V14(0) ,
  V480 = V2269 | V2268,
  V481 = ~\V476(0)  & ~\V473(0) ,
  V482 = V2273 | V2272,
  V483 = V481 & ~\V470(0) ,
  V484 = V2277 | V2276,
  V485 = V1850 & V451,
  V486 = V484 & ~V1850,
  V488 = V1850 & V446,
  V489 = V482 & ~V1850,
  \[184]  = ~\V261(0) ,
  V491 = V1850 & V441,
  V492 = V480 & ~V1850,
  V494 = V1850 & V437,
  V495 = ~\V476(0)  & ~V1850,
  V499 = \V14(0)  & ~\V271(0) ,
  \[185]  = ~\V301(0) ,
  \[186]  = ~\V302(0) ,
  \V1147(10)  = V1136 | V1128,
  \[187]  = V1750 | (V1476 | V1889),
  \V1147(11)  = V1134 | V1127,
  \V378(0)  = V766 | V701,
  \[188]  = V1890 | V1885,
  \[189]  = V1891 | V1886,
  V2800 = ~V2052 & V2045,
  V2801 = V2052 & ~V2045,
  V2804 = V2047 & ~V2054,
  V2805 = ~V2047 & V2054,
  V2808 = \V2067(0)  & \V2064(0) ,
  V2809 = ~\V2067(0)  & ~\V2064(0) ,
  V2812 = ~V2072 & \V2061(0) ,
  V2813 = V2072 & ~\V2061(0) ,
  V2816 = ~V2074 & \V2058(0) ,
  V2817 = V2074 & ~\V2058(0) ,
  V501 = V710 & ~V687,
  V502 = V710 & V687,
  V505 = \V503(0)  & \V56(0) ,
  V506 = \V504(0)  & \V56(0) ,
  V507 = \V59(0)  & V502,
  V509 = V2281 | V2280,
  V512 = \[15] ,
  V513 = V400 & \V56(0) ,
  V514 = \V56(0)  & V728,
  V515 = \V730(0)  & V687,
  V516 = V515 & \V59(0) ,
  V517 = \V729(0)  & (~V687 & \V59(0) ),
  V518 = \V59(0)  & \V731(0) ,
  V525 = ~V518 & (~V517 & (~V516 & (~V514 & (~V513 & ~V402)))),
  V527 = \[16] ,
  V529 = \V45(0)  & ~\V43(0) ,
  V530 = V2285 | V2284,
  V531 = V2289 | V2288,
  V534 = \V149(7)  & (V701 & \V56(0) ),
  V535 = V701 & V1646,
  V537 = \[17] ,
  V538 = \[18] ,
  V539 = \[19] ,
  V540 = \[20] ,
  V541 = \[21] ,
  V542 = \[22] ,
  V543 = \[23] ,
  V544 = \[24] ,
  V545 = \[25] ,
  V546 = \[26] ,
  V547 = \[27] ,
  V548 = \[28] ,
  V549 = ~\V2019(0)  & (V2104 & (V727 & (\[65]  & \V149(7) ))),
  \[190]  = V1892 | V1887,
  V550 = ~\V2019(0)  & (V2104 & (V727 & (\[65]  & \V149(6) ))),
  V551 = ~\V2019(0)  & (V2104 & (V727 & (\[65]  & \V149(5) ))),
  V552 = ~\V2019(0)  & (V2104 & (V727 & (\[65]  & \V149(4) ))),
  V553 = V2106 & (\V2019(0)  & (V2107 & ~\V199(4) )),
  V555 = V2106 & (\V2019(0)  & (V2107 & V1883)),
  V557 = V2106 & (\V2019(0)  & (V2107 & V1882)),
  V559 = V2106 & (\V2019(0)  & (V2107 & V1881)),
  \[191]  = V1893 | V1751,
  \V729(0)  = V717 | (V715 | (V713 | (V711 | (V712 | (V714 | (V716 | V718)))))),
  V561 = V2106 & (\V2019(0)  & (V2107 & V1880)),
  V563 = V2106 & (\V2019(0)  & (V2107 & V1879)),
  V565 = V2106 & (\V2019(0)  & (V2107 & V1878)),
  V567 = V2106 & (\V2019(0)  & (V2107 & V1877)),
  V569 = V2106 & (\V2019(0)  & (V2107 & V1876)),
  \[192]  = V1895 | V1752,
  V571 = V2106 & (\V2019(0)  & (V2107 & V1875)),
  V573 = V2109 & (~\V2019(0)  & (V769 & (\[82]  & \[65] ))),
  V574 = V2109 & (~\V2019(0)  & (V769 & (\[83]  & \[65] ))),
  V575 = V2109 & (~\V2019(0)  & (V769 & (\[84]  & \[65] ))),
  V576 = V2109 & (~\V2019(0)  & (V769 & (\[85]  & \[65] ))),
  V577 = V2109 & (~\V2019(0)  & (V769 & (\[86]  & \[65] ))),
  V578 = V2109 & (~\V2019(0)  & (V769 & (\[87]  & \[65] ))),
  V579 = V2109 & (~\V2019(0)  & (V769 & (\[88]  & \[65] ))),
  \[193]  = V1922 | (V1910 | V1904),
  V580 = V2109 & (~\V2019(0)  & (V769 & (\[89]  & \[65] ))),
  V581 = V2109 & (~\V2019(0)  & (V769 & (\[90]  & \[65] ))),
  V582 = V2109 & (~\V2019(0)  & (V769 & (\[91]  & \[65] ))),
  V587 = \[40] ,
  V589 = ~V341 & (~\V244(0)  & \V243(0) ),
  \[194]  = V1928 | (V1923 | (V1912 | V1905)),
  V590 = ~V341 & (\V244(0)  & ~\V243(0) ),
  V593 = \V244(0)  & \V243(0) ,
  V594 = V593 & (~V341 & ~\V245(0) ),
  V596 = ~V593 & (~V341 & \V245(0) ),
  V599 = \V245(0)  & V593,
  \[195]  = V1929 | (V1924 | (V1914 | V1906)),
  \[196]  = V1930 | (V1925 | (V1916 | V1907)),
  \[197]  = V1931 | (V1926 | (V1918 | V1908)),
  \[198]  = V1932 | (V1927 | (V1920 | V1909)),
  \V1398(0)  = \V57(0)  | (\V53(0)  | \V56(0) ),
  \[199]  = ~V751 & (~V743 & (V742 & \V132(1) )),
  V600 = V599 & (~V341 & ~\V246(0) ),
  V602 = ~V599 & (~V341 & \V246(0) ),
  V605 = \V246(0)  & V599,
  V606 = V605 & (~V341 & ~\V247(0) ),
  V608 = ~V605 & (~V341 & \V247(0) ),
  \V1337(0)  = V1336 | V1335,
  V611 = V739 & ~V1476,
  V613 = \V62(0)  & V741,
  V614 = V505 & (~V1646 & (~V695 & ~\V214(0) )),
  V615 = \V612(0)  & (~V695 & (~\V214(0)  & \V59(0) )),
  V616 = V741 & (~V695 & (~\V214(0)  & \V62(0) )),
  \V470(0)  = V469 | V468,
  V620 = \[45] ,
  V621 = \[46] ,
  V623 = \V62(0)  & V745,
  V626 = \[65]  & (\V1647(0)  & V1445),
  V627 = ~V1735 & (V1445 & \V59(0) ),
  V628 = \V56(0)  & V745,
  V630 = \[47] ,
  V631 = ~V637 & (\V269(0)  & \V271(0) ),
  V632 = ~V637 & (\V274(0)  & ~\V271(0) ),
  V637 = ~\V202(0)  & (\V274(0)  & ~\V271(0) ),
  V638 = ~V637 & ~\V271(0) ,
  V644 = \V257(6)  & (\V257(4)  & (\V257(2)  & (\V257(1)  & (\V257(3)  & (\V257(5)  & \V257(7) ))))),
  V645 = \V257(6)  & (\V257(4)  & (\V257(2)  & (\V257(3)  & (\V257(5)  & \V257(7) )))),
  V646 = \V257(6)  & (\V257(4)  & (\V257(3)  & (\V257(5)  & \V257(7) ))),
  V647 = \V257(6)  & (\V257(4)  & (\V257(5)  & \V257(7) )),
  V648 = \V257(6)  & (\V257(5)  & \V257(7) ),
  V649 = \V257(6)  & \V257(7) ,
  V650 = \[212] ,
  V651 = \[213] ,
  V652 = \[214] ,
  V653 = \[215] ,
  V654 = \[216] ,
  V655 = \[217] ,
  V656 = \[218] ,
  V657 = \[50] ,
  V687 = \V169(1)  & \V1395(0) ,
  V695 = \V165(1)  & (~\V165(2)  & \V165(0) ),
  V696 = V695 & (~\V290(0)  & \V165(7) ),
  V697 = \V165(1)  & (\V165(2)  & (~\V165(0)  & \V203(0) )),
  V698 = V695 & ~\V165(7) ,
  \V821(0)  = \[66] ,
  \V1552(1)  = \[142] ,
  \V1552(0)  = \[143] ,
  \V1687(0)  = V1686 | \V1674(0) ,
  V700 = ~\V149(2)  & (~\V149(1)  & ~\V149(0) ),
  V701 = \V149(2)  & (~\V149(1)  & ~\V149(0) ),
  V702 = ~\V149(2)  & (\V149(1)  & ~\V149(0) ),
  V703 = \V149(2)  & (~\V149(1)  & \V149(0) ),
  V704 = \V149(1)  & (\V149(0)  & \V149(2) ),
  V706 = ~\V149(2)  & (\V149(1)  & \V149(0) ),
  V707 = \[51] ,
  V710 = V766 & \V149(3) ,
  V711 = \[51]  & (\V149(4)  & ~\V149(5) ),
  V712 = \V149(4)  & (\[51]  & \V149(5) ),
  V713 = \[51]  & (\V88(3)  & (~\V88(2)  & (~\V149(4)  & ~\V149(5) ))),
  V714 = \[51]  & (~\V88(3)  & (\V88(2)  & (~\V149(4)  & ~\V149(5) ))),
  V715 = \[51]  & (\V88(3)  & (\V88(2)  & (~\V149(4)  & ~\V149(5) ))),
  V716 = V766 & (~\V88(3)  & (~\V88(2)  & (~\V149(3)  & (~\V149(4)  & \V149(5) )))),
  V717 = V766 & (\V88(3)  & (~\V88(2)  & (~\V149(3)  & (~\V149(4)  & \V149(5) )))),
  V718 = V766 & (~\V88(3)  & (\V88(2)  & (~\V149(3)  & (~\V149(4)  & \V149(5) )))),
  V719 = \[51]  & (~\V88(3)  & (~\V88(2)  & (~\V149(4)  & ~\V149(5) ))),
  V720 = V766 & (\V88(3)  & (\V88(2)  & (~\V149(3)  & (~\V149(4)  & \V149(5) )))),
  V721 = V701 & \V149(3) ,
  V722 = V701 & (~\V149(3)  & (~\V149(4)  & ~\V149(5) )),
  V723 = V701 & (~\V149(3)  & (~\V149(4)  & \V149(5) )),
  V724 = V701 & (~\V149(3)  & (\V149(4)  & ~\V149(5) )),
  V725 = ~\V149(3)  & (\V149(2)  & (\V149(1)  & (~\V149(0)  & \V149(4) ))),
  V726 = ~\V149(3)  & (\V149(2)  & (\V149(1)  & (~\V149(0)  & ~\V149(4) ))),
  V727 = \V149(3)  & (\V149(2)  & (\V149(1)  & ~\V149(0) )),
  V728 = V701 & (~\V149(3)  & (\V149(4)  & \V149(5) )),
  V734 = \V729(0)  & ~V687,
  V735 = V702 & (~\V149(3)  & (~\V149(4)  & (~\V149(5)  & (~\V149(6)  & \V149(7) )))),
  V736 = V702 & (~\V149(3)  & (~\V149(4)  & (~\V149(5)  & (\V149(6)  & ~\V149(7) )))),
  V737 = V702 & (~\V149(3)  & (~\V149(4)  & (~\V149(5)  & (\V149(6)  & \V149(7) )))),
  V738 = V702 & (~\V149(3)  & (~\V149(4)  & (\V149(5)  & (~\V149(6)  & ~\V149(7) )))),
  V739 = V702 & (~\V149(3)  & (~\V149(4)  & (\V149(5)  & (~\V149(6)  & \V149(7) )))),
  V740 = V702 & (~\V149(3)  & (~\V149(4)  & (\V149(5)  & (\V149(6)  & ~\V149(7) )))),
  V741 = V702 & (~\V149(3)  & (~\V149(4)  & (\V149(5)  & (\V149(6)  & \V149(7) )))),
  V742 = V702 & (~\V149(3)  & (\V149(4)  & (~\V149(5)  & (~\V149(6)  & ~\V149(7) )))),
  V743 = V702 & (~\V149(3)  & (\V149(4)  & (~\V149(5)  & (~\V149(6)  & \V149(7) )))),
  V744 = V702 & (~\V149(3)  & (\V149(4)  & (~\V149(5)  & (\V149(6)  & ~\V149(7) )))),
  V745 = V702 & (~\V149(3)  & (\V149(4)  & (~\V149(5)  & (\V149(6)  & \V149(7) )))),
  V746 = V702 & (~\V149(3)  & (\V149(4)  & (\V149(5)  & (~\V149(6)  & \V149(7) )))),
  V747 = V702 & (~\V149(3)  & (\V149(4)  & (\V149(5)  & (\V149(6)  & ~\V149(7) )))),
  V748 = V702 & (~\V149(3)  & (\V149(4)  & (\V149(5)  & (\V149(6)  & \V149(7) )))),
  V749 = V702 & (\V149(3)  & (~\V149(4)  & (~\V149(5)  & (~\V149(6)  & ~\V149(7) )))),
  V750 = V702 & (\V149(3)  & (~\V149(4)  & (~\V149(5)  & (~\V149(6)  & \V149(7) )))),
  V751 = V702 & (\V149(3)  & (~\V149(4)  & (~\V149(5)  & (\V149(6)  & ~\V149(7) )))),
  V755 = ~V751 & (~V750 & (V702 & (~V749 & \V149(3) ))),
  V756 = V702 & (~\V149(3)  & (~\V149(4)  & (~\V149(5)  & (~\V149(6)  & ~\V149(7) )))),
  V757 = V702 & (~\V149(3)  & (\V149(4)  & (\V149(5)  & (~\V149(6)  & ~\V149(7) )))),
  V761 = \V759(0)  & (~\[65]  & ~\V55(0) ),
  V763 = \[52] ,
  V766 = V700 & ~\V174(0) ,
  V767 = V747 & ~\V174(0) ,
  V768 = V748 & ~\V174(0) ,
  V769 = V725 & ~\V174(0) ,
  V774 = ~\V758(0)  & (~V706 & (~V704 & ~V703)),
  V775 = \[53] ,
  V776 = V345 & ~\V174(0) ,
  V778 = \[54] ,
  V779 = \[55] ,
  V780 = \[56] ,
  V781 = \[57] ,
  V782 = \[58] ,
  V783 = \[59] ,
  V784 = \[60] ,
  V787 = \[61] ,
  V789 = \[62] ,
  V790 = \V758(0)  & ~\V302(0) ,
  V794 = ~V790 & (~V774 & ~\V1681(0) ),
  V797 = ~\V817(0)  & (~V794 & \V14(0) ),
  V799 = \V165(3)  & (~\V165(6)  & (~\V165(5)  & (~\V165(4)  & \V70(0) ))),
  \V1053(7)  = V1038 | V1026,
  \V445(0)  = V443 | (V442 | V444),
  \V1053(6)  = V1040 | V1027,
  V801 = \[64] ,
  V806 = ~V739 & ~V740,
  V808 = V741 & \V65(0) ,
  \V1053(9)  = V1034 | V1024,
  V811 = ~V806 & \V62(0) ,
  V814 = \V812(0)  & (~V698 & ~\[163] ),
  V815 = ~V1735 & \V813(0) ,
  V816 = ~V695 & \V290(0) ,
  V818 = V340 & \V149(5) ,
  \V1053(8)  = V1036 | V1025,
  V820 = ~V340 & ~\V279(0) ,
  V823 = V340 & \V149(4) ,
  V824 = V820 & ~\V280(0) ,
  V825 = ~V340 & (\V280(0)  & \V279(0) ),
  V828 = V2321 | V2320,
  V829 = V2325 | V2324,
  V830 = V2329 | V2328,
  V831 = V2333 | V2332,
  V836 = \V1855(0)  & (~V831 & (~V830 & (~V829 & (~V828 & ~V433)))),
  V838 = V2337 | V2336,
  V839 = V2341 | V2340,
  V840 = V2345 | V2344,
  V841 = V2349 | V2348,
  V846 = ~V841 & (~V840 & (~V839 & (~V838 & (~V433 & \V288(4) )))),
  V848 = V2353 | V2352,
  V849 = V2357 | V2356,
  \V1853(0)  = \V288(0)  | \V288(1) ,
  V850 = V2361 | V2360,
  V851 = V2365 | V2364,
  \V383(0)  = ~V349 | ~V348,
  V856 = ~V851 & (~V850 & (~V849 & (~V848 & (~V433 & V1840)))),
  V858 = V2369 | V2368,
  V859 = V2373 | V2372,
  V860 = V2377 | V2376,
  V861 = V2381 | V2380,
  V866 = ~V861 & (~V860 & (~V859 & (~V858 & (~V433 & V1840)))),
  V868 = V2385 | V2384,
  V869 = V2389 | V2388,
  V870 = V2393 | V2392,
  V871 = V2397 | V2396,
  V876 = \V1854(0)  & (~V871 & (~V870 & (~V869 & (~V868 & ~V433)))),
  V878 = V2401 | V2400,
  V879 = V2405 | V2404,
  V880 = V2409 | V2408,
  V881 = V2413 | V2412,
  V886 = ~V881 & (~V880 & (~V879 & (~V878 & (~V433 & \V288(2) )))),
  V888 = V2417 | V2416,
  V889 = V2421 | V2420,
  \V1053(1)  = V1050 | V1032,
  V890 = V2425 | V2424,
  V891 = V2429 | V2428,
  V896 = ~V891 & (~V890 & (~V889 & (~V888 & (~V433 & V1839)))),
  V898 = V2433 | V2432,
  V899 = V2437 | V2436,
  \V1053(0)  = V1052 | V1033,
  \V1053(3)  = V1046 | V1030,
  \V1053(2)  = V1048 | V1031,
  \V1053(5)  = V1042 | V1028,
  \V1053(4)  = V1044 | V1029,
  V900 = V2441 | V2440,
  V901 = V2445 | V2444,
  V906 = ~V901 & (~V900 & (~V899 & (~V898 & (~V433 & V1839)))),
  V908 = V2449 | V2448,
  V909 = V2453 | V2452,
  V910 = V2457 | V2456,
  V911 = V2461 | V2460,
  V916 = \V1853(0)  & (~V911 & (~V910 & (~V909 & (~V908 & ~V433)))),
  V918 = V2465 | V2464,
  V919 = V2469 | V2468,
  V920 = V2473 | V2472,
  V921 = V2477 | V2476,
  V926 = ~V921 & (~V920 & (~V919 & (~V918 & (~V433 & \V288(0) )))),
  V928 = V2481 | V2480,
  V929 = V2485 | V2484,
  V930 = V2489 | V2488,
  V931 = V2493 | V2492,
  V936 = ~V931 & (~V930 & (~V929 & (~V928 & (~V433 & V1838)))),
  V938 = V2497 | V2496,
  V939 = V2501 | V2500,
  V940 = V2505 | V2504,
  V941 = V2509 | V2508,
  \V408(0)  = V407 | (V406 | V402),
  V946 = ~V941 & (~V940 & (~V939 & (~V938 & (~V433 & V1838)))),
  V952 = \V1856(0)  & (~\V1255(3)  & (~\V1255(2)  & (~\V1255(1)  & (~\V1255(0)  & ~V433)))),
  V953 = \V1255(3)  & (~\V1255(2)  & (~\V1255(1)  & (~\V1255(0)  & (~V433 & \V288(6) )))),
  V954 = ~\V1255(3)  & (\V1255(2)  & (~\V1255(1)  & (~\V1255(0)  & (~V433 & (\V288(7)  & \V288(6) ))))),
  V955 = \V1255(3)  & (\V1255(2)  & (~\V1255(1)  & (~\V1255(0)  & (~V433 & (\V288(7)  & \V288(6) ))))),
  V960 = ~V794 & \[65] ,
  V961 = \V777(0)  & (\V759(0)  & (\[52]  & \V56(0) )),
  V962 = \V758(0)  & \V56(0) ,
  V963 = \V759(0)  & V799,
  V966 = \[68] ,
  V968 = \V1681(0)  & (~\V260(0)  & (~\V259(0)  & (\V258(0)  & ~\V59(0) ))),
  V976 = ~V968 & (~V746 & (~V743 & (~V742 & (~V736 & (~V735 & ~V744))))),
  V978 = V976 & (~V961 & (~\V758(0)  & \V56(0) )),
  V981 = ~V976 & \V56(0) ,
  V983 = \V982(0)  & \V59(0) ,
  V984 = \V1681(0)  & \V62(0) ,
  V986 = \[69] ,
  V988 = \V1395(0)  & (~\V2011(0)  & \V229(5) ),
  V989 = \V1395(0)  & (~\V2011(0)  & \V229(4) ),
  V990 = \V1395(0)  & (~\V2011(0)  & \V229(3) ),
  V991 = \V1395(0)  & (~\V2011(0)  & \V229(2) ),
  V992 = \V1395(0)  & (~\V2011(0)  & \V229(1) ),
  V993 = \V1395(0)  & (~\V2011(0)  & \V229(0) ),
  V994 = \V1395(0)  & (~\V2011(0)  & \V223(5) ),
  V995 = \V1395(0)  & (~\V2011(0)  & \V223(4) ),
  V996 = \V1395(0)  & (~\V2011(0)  & \V223(3) ),
  V997 = \V1395(0)  & (~\V2011(0)  & \V223(2) ),
  V998 = \V1395(0)  & (~\V2011(0)  & \V223(1) ),
  V999 = \V1395(0)  & (~\V2011(0)  & \V223(0) );
endmodule

