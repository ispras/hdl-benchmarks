// IWLS benchmark module "MultiplierB_16" printed on Wed May 29 22:12:33 2002
module MultiplierB_16(\1 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \13 , \14 , \15 , \16 , \17 , \18 , \50 );
input
  \1 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ,
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ;
output
  \50 ;
reg
  \2 ,
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ,
  \34 ,
  \35 ,
  \36 ,
  \37 ,
  \38 ,
  \39 ,
  \40 ,
  \41 ,
  \42 ,
  \43 ,
  \44 ,
  \45 ,
  \46 ,
  \47 ,
  \48 ;
wire
  \164 ,
  \168 ,
  \169 ,
  \[45] ,
  \173 ,
  \174 ,
  \178 ,
  \179 ,
  \[70] ,
  \[46] ,
  \183 ,
  \184 ,
  \188 ,
  \191 ,
  \[71] ,
  \[47] ,
  \194 ,
  \197 ,
  \[72] ,
  \[48] ,
  \[73] ,
  \[49] ,
  \[74] ,
  \[75] ,
  \200 ,
  \203 ,
  \206 ,
  \209 ,
  \212 ,
  \215 ,
  \218 ,
  \221 ,
  \[50] ,
  \224 ,
  \227 ,
  \230 ,
  \[51] ,
  \233 ,
  \235 ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ,
  \[59] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \[60] ,
  \[36] ,
  \[61] ,
  \[37] ,
  \[62] ,
  \[38] ,
  \[63] ,
  \[39] ,
  \[64] ,
  \[65] ,
  \[66] ,
  \[67] ,
  \[68] ,
  \[69] ,
  \114 ,
  \118 ,
  \119 ,
  \[40] ,
  \123 ,
  \124 ,
  \128 ,
  \129 ,
  \[41] ,
  \133 ,
  \134 ,
  \138 ,
  \139 ,
  \[42] ,
  \143 ,
  \144 ,
  \148 ,
  \149 ,
  \[43] ,
  \153 ,
  \154 ,
  \158 ,
  \159 ,
  \[44] ,
  \163 ;
assign
  \164  = (~\[71]  & ~\221 ) | (\[71]  & \221 ),
  \168  = (~\164  & \221 ) | (~\221  & \44 ),
  \169  = (~\[72]  & ~\224 ) | (\[72]  & \224 ),
  \[45]  = \184 ,
  \173  = (~\169  & \224 ) | (~\224  & \45 ),
  \174  = (~\[73]  & ~\227 ) | (\[73]  & \227 ),
  \178  = (~\174  & \227 ) | (~\227  & \46 ),
  \179  = (~\[74]  & ~\230 ) | (\[74]  & \230 ),
  \[70]  = ~\12  | ~\1 ,
  \[46]  = \118 ,
  \183  = (~\179  & \230 ) | (~\230  & \47 ),
  \184  = (~\[75]  & ~\233 ) | (\[75]  & \233 ),
  \188  = (~\184  & \233 ) | (~\233  & \48 ),
  \191  = (~\20  & \34 ) | (\20  & ~\34 ),
  \[71]  = ~\13  | ~\1 ,
  \[47]  = \123 ,
  \194  = (~\21  & \35 ) | (\21  & ~\35 ),
  \197  = (~\22  & \36 ) | (\22  & ~\36 ),
  \[72]  = ~\14  | ~\1 ,
  \[48]  = \128 ,
  \[73]  = ~\15  | ~\1 ,
  \[49]  = \133 ,
  \[74]  = ~\16  | ~\1 ,
  \[75]  = ~\17  | ~\1 ,
  \200  = (~\23  & \37 ) | (\23  & ~\37 ),
  \203  = (~\24  & \38 ) | (\24  & ~\38 ),
  \206  = (~\25  & \39 ) | (\25  & ~\39 ),
  \209  = (~\26  & \40 ) | (\26  & ~\40 ),
  \212  = (~\27  & \41 ) | (\27  & ~\41 ),
  \215  = (~\28  & \42 ) | (\28  & ~\42 ),
  \218  = (~\29  & \43 ) | (\29  & ~\43 ),
  \221  = (~\30  & \44 ) | (\30  & ~\44 ),
  \[50]  = \138 ,
  \224  = (~\31  & \45 ) | (\31  & ~\45 ),
  \227  = (~\32  & \46 ) | (\32  & ~\46 ),
  \230  = (~\33  & \47 ) | (\33  & ~\47 ),
  \[51]  = \143 ,
  \233  = (~\2  & \48 ) | (\2  & ~\48 ),
  \235  = \18  & \1 ,
  \[52]  = \148 ,
  \50  = \114 ,
  \[53]  = \153 ,
  \[54]  = \158 ,
  \[55]  = \163 ,
  \[56]  = \168 ,
  \[57]  = \173 ,
  \[58]  = \178 ,
  \[59]  = \183 ,
  \[31]  = \235 ,
  \[32]  = \119 ,
  \[33]  = \124 ,
  \[34]  = \129 ,
  \[35]  = \134 ,
  \[60]  = \188 ,
  \[36]  = \139 ,
  \[61]  = ~\3  | ~\1 ,
  \[37]  = \144 ,
  \[62]  = ~\4  | ~\1 ,
  \[38]  = \149 ,
  \[63]  = ~\5  | ~\1 ,
  \[39]  = \154 ,
  \[64]  = ~\6  | ~\1 ,
  \[65]  = ~\7  | ~\1 ,
  \[66]  = ~\8  | ~\1 ,
  \[67]  = ~\9  | ~\1 ,
  \[68]  = ~\10  | ~\1 ,
  \[69]  = ~\11  | ~\1 ,
  \114  = (~\[61]  & ~\191 ) | (\[61]  & \191 ),
  \118  = (~\114  & \191 ) | (~\191  & \34 ),
  \119  = (~\[62]  & ~\194 ) | (\[62]  & \194 ),
  \[40]  = \159 ,
  \123  = (~\119  & \194 ) | (~\194  & \35 ),
  \124  = (~\[63]  & ~\197 ) | (\[63]  & \197 ),
  \128  = (~\124  & \197 ) | (~\197  & \36 ),
  \129  = (~\[64]  & ~\200 ) | (\[64]  & \200 ),
  \[41]  = \164 ,
  \133  = (~\129  & \200 ) | (~\200  & \37 ),
  \134  = (~\[65]  & ~\203 ) | (\[65]  & \203 ),
  \138  = (~\134  & \203 ) | (~\203  & \38 ),
  \139  = (~\[66]  & ~\206 ) | (\[66]  & \206 ),
  \[42]  = \169 ,
  \143  = (~\139  & \206 ) | (~\206  & \39 ),
  \144  = (~\[67]  & ~\209 ) | (\[67]  & \209 ),
  \148  = (~\144  & \209 ) | (~\209  & \40 ),
  \149  = (~\[68]  & ~\212 ) | (\[68]  & \212 ),
  \[43]  = \174 ,
  \153  = (~\149  & \212 ) | (~\212  & \41 ),
  \154  = (~\[69]  & ~\215 ) | (\[69]  & \215 ),
  \158  = (~\154  & \215 ) | (~\215  & \42 ),
  \159  = (~\[70]  & ~\218 ) | (\[70]  & \218 ),
  \[44]  = \179 ,
  \163  = (~\159  & \218 ) | (~\218  & \43 );
always begin
  \2  = \[31] ;
  \20  = \[32] ;
  \21  = \[33] ;
  \22  = \[34] ;
  \23  = \[35] ;
  \24  = \[36] ;
  \25  = \[37] ;
  \26  = \[38] ;
  \27  = \[39] ;
  \28  = \[40] ;
  \29  = \[41] ;
  \30  = \[42] ;
  \31  = \[43] ;
  \32  = \[44] ;
  \33  = \[45] ;
  \34  = \[46] ;
  \35  = \[47] ;
  \36  = \[48] ;
  \37  = \[49] ;
  \38  = \[50] ;
  \39  = \[51] ;
  \40  = \[52] ;
  \41  = \[53] ;
  \42  = \[54] ;
  \43  = \[55] ;
  \44  = \[56] ;
  \45  = \[57] ;
  \46  = \[58] ;
  \47  = \[59] ;
  \48  = \[60] ;
end
initial begin
  \2  = 0;
  \20  = 0;
  \21  = 0;
  \22  = 0;
  \23  = 0;
  \24  = 0;
  \25  = 0;
  \26  = 0;
  \27  = 0;
  \28  = 0;
  \29  = 0;
  \30  = 0;
  \31  = 0;
  \32  = 0;
  \33  = 0;
  \34  = 0;
  \35  = 0;
  \36  = 0;
  \37  = 0;
  \38  = 0;
  \39  = 0;
  \40  = 0;
  \41  = 0;
  \42  = 0;
  \43  = 0;
  \44  = 0;
  \45  = 0;
  \46  = 0;
  \47  = 0;
  \48  = 0;
end
endmodule

