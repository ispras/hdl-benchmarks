//NOTE: no-implementation module stub

module lmi_watchd (
    input wire CLK,
    input wire TMODE,
    input wire RESET_D1_R_N,
    input wire X_HALT_R,
    input wire C_IADDR_A,
    input wire IX_MISS_S_R,
    input wire IX_VAL,
    input wire DC_MISS_W_R,
    input wire DC_VAL,
    input wire LW_IADDR_S_R,
    input wire anyIMiss_S,
    input wire anyIVal,
    input wire anyDMiss_W,
    input wire anyDVal,
    input wire anyIBusy,
    input wire anyDBusy
);

endmodule
