// IWLS benchmark module "cordic" printed on Wed May 29 16:31:29 2002
module cordic(a6, a4, a3, a2, a5, v, x0, x1, x2, x3, y0, y1, y2, y3, z0, z1, z2, ex0, ex1, ex2, ey0, ey1, ey2, d, dn);
input
  ex0,
  ex1,
  ex2,
  ey0,
  ey1,
  ey2,
  v,
  x0,
  x1,
  x2,
  x3,
  y0,
  y1,
  y2,
  y3,
  z0,
  z1,
  z2,
  a2,
  a3,
  a4,
  a5,
  a6;
output
  dn,
  d;
wire
  \[157] ,
  \[646] ,
  \[574] ,
  \[123] ,
  \[540] ,
  \[90] ,
  \[526] ,
  \[124] ,
  \[367] ,
  \[590] ,
  \[91] ,
  \[576] ,
  \[614] ,
  \[77] ,
  \[368] ,
  \[542] ,
  \[78] ,
  \[592] ,
  \[630] ,
  \[578] ,
  \[616] ,
  \[350] ,
  \[544] ,
  \[128] ,
  \[594] ,
  \[632] ,
  \[129] ,
  \[618] ,
  \[511] ,
  \[546] ,
  \[596] ,
  \[634] ,
  \[0] ,
  \[514] ,
  \[598] ,
  \[636] ,
  \[321] ,
  \[1] ,
  \[516] ,
  \[250] ,
  \[638] ,
  \[580] ,
  \[237] ,
  \[130] ,
  \[582] ,
  \[568] ,
  \[117] ,
  \[375] ,
  \[118] ,
  \[584] ,
  \[376] ,
  \[119] ,
  \[608] ,
  \[586] ,
  \[503] ,
  \[552] ,
  \[640] ,
  \[588] ,
  \[626] ,
  \[360] ,
  \[505] ,
  \[554] ,
  \[642] ,
  \[347] ,
  \[628] ,
  \[570] ,
  \[522] ,
  \[120] ,
  \[363] ,
  \[508] ,
  \[644] ,
  \[572] ,
  \[524] ;
assign
  \[157]  = ~\[90]  & ~\[91] ,
  \[646]  = ~y1 | y0,
  \[574]  = ~\[554]  | z0,
  \[123]  = ~\[77]  & ex1,
  \[540]  = ~\[570]  | (~\[508]  | ~\[505] ),
  dn = \[1] ,
  \[90]  = ~\[118]  & ~\[117] ,
  \[526]  = ~\[628]  | (~\[626]  | (~\[630]  | ~\[250] )),
  \[124]  = ~\[78]  & ~ex1,
  \[367]  = ~\[598]  | ~\[596] ,
  \[590]  = ~\[368]  | \[367] ,
  \[91]  = ~\[120]  & ~\[119] ,
  \[576]  = \[376]  | ~\[375] ,
  \[614]  = ~ey1 | ~\[522] ,
  \[77]  = ex2 & ex0,
  \[368]  = ~\[594]  | ~\[592] ,
  \[542]  = ~\[574]  | ~\[572] ,
  \[78]  = ~ex2 & ~ex0,
  \[592]  = x3 | ~x2,
  \[630]  = \[360]  | ~\[363] ,
  \[578]  = ~\[376]  | \[375] ,
  \[616]  = ~\[524]  | ey1,
  \[350]  = ~\[634]  | ~\[632] ,
  \[544]  = ~\[578]  | ~\[576] ,
  \[128]  = ~z2 & (~z1 & z0),
  d = \[0] ,
  \[594]  = ~x3 | x2,
  \[632]  = y3 | ~y2,
  \[129]  = z2 & (z1 & ~z0),
  \[618]  = ~\[526]  | ~\[508] ,
  \[511]  = ~\[321]  | (a3 | (a4 | a6)),
  \[546]  = ~\[590]  | ~\[588] ,
  \[596]  = x1 | x0,
  \[634]  = ~y3 | y2,
  \[0]  = ~\[503] ,
  \[514]  = ~\[608]  | v,
  \[598]  = ~x1 | ~x0,
  \[636]  = x3 | ~x2,
  \[321]  = ~a5 & ~a2,
  \[1]  = ~\[568]  | ~\[511] ,
  \[516]  = ~\[618]  | (~\[616]  | (~\[237]  | ~\[614] )),
  \[250]  = ~\[129]  & (~\[128]  & ~\[130] ),
  \[638]  = ~x3 | x2,
  \[580]  = y3 | ~y2,
  \[237]  = ~\[124]  & ~\[123] ,
  \[130]  = ~\[350]  & \[347] ,
  \[582]  = ~y3 | y2,
  \[568]  = ~\[540]  | v,
  \[117]  = ~ey1 & (~ey0 & ~ey2),
  \[375]  = ~\[586]  | ~\[584] ,
  \[118]  = ey2 & (ey1 & ey0),
  \[584]  = y1 | y0,
  \[376]  = ~\[582]  | ~\[580] ,
  \[119]  = ~ex1 & (~ex0 & ~ex2),
  \[608]  = ~\[516]  | ~\[505] ,
  \[586]  = ~y1 | ~y0,
  \[503]  = ~\[514]  | ~\[511] ,
  \[552]  = z2 | z1,
  \[640]  = x1 | ~x0,
  \[588]  = \[368]  | ~\[367] ,
  \[626]  = ~\[350]  | \[347] ,
  \[360]  = ~\[642]  | ~\[640] ,
  \[505]  = a2 | (a3 | (~a4 | ~a6)),
  \[554]  = ~z1 | ~z2,
  \[642]  = ~x1 | x0,
  \[347]  = ~\[646]  | ~\[644] ,
  \[628]  = ~\[360]  | \[363] ,
  \[570]  = ~\[542]  | (~\[544]  | (~\[157]  | ~\[546] )),
  \[522]  = ~ey2 | ~ey0,
  \[120]  = ex2 & (ex1 & ex0),
  \[363]  = ~\[638]  | ~\[636] ,
  \[508]  = a2 | (~a3 | (a4 | ~a6)),
  \[644]  = y1 | ~y0,
  \[572]  = ~z0 | ~\[552] ,
  \[524]  = ey2 | ey0;
endmodule

