//NOTE: no-implementation module stub

module lmi_icache (
    input wire CLK,
    input wire TMODE,
    input wire RESET_D1_R_N,
    input wire DISABLEC,
    input wire INVALIDATE,
    input wire MEMSEQUENTIAL,
    input wire MEMZEROFIRST,
    input wire EXT_ICREQRAM_R,
    input wire IC_GNTRAM_R,
    input wire NEXTADDR,
    input wire RDOP_N,
    output wire IS_VAL,
    output wire IC_VAL,
    output wire LACK,
    output wire X_HALT_R,
    output wire IC_MISS_P,
    output wire IC_MISS_R,
    output wire IC_HALT_S_R,
    input wire IC_TAGINDEX,
    input wire ICR_TAGRD0,
    input wire IC_TAGWR0,
    input wire IC_TAG0WE,
    input wire IC_TAG0WEN,
    input wire IC_TAG0RE,
    input wire IC_TAG0REN,
    input wire IC_TAG0CS,
    input wire IC_TAG0CSN,
    input wire IC_DATAINDEX,
    input wire IC_DATA0WE,
    input wire IC_DATA0WEN,
    input wire IC_DATA0RE,
    input wire IC_DATA0REN,
    input wire IC_DATA0CS,
    input wire IC_DATA0CSN,
    output wire IC_DATAOE,
    output wire IC_LBCOE,
    input wire ICC_TAGMASK,
    output wire IC_TAG0COMPARE
);

endmodule
