//NOTE: no-implementation module stub

module pcont_cop0 (
    input wire [31:0] INST_S_R,
    input wire SYSCLK,
    input wire TMODE,
    input wire RESET_D1_R_N,
    input wire [31:0] INST_I,
    input wire CP0_INSTM32_I_R_N,
    input wire CP0_M16IADDRB1_I,
    input wire CLMI_RHOLD,
    input wire CLMI_SELINST_S_P
);

endmodule
