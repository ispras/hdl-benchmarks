//NOTE: no-implementation module stub

module INVGSS (
    output O,
    input I
);
endmodule

module XOSCAHB (
    inout wire IO,
    input wire I,
    input wire E,
    output wire O,
    input wire FEB,
    input wire EB,
    input wire S0,
    input wire S1
);
endmodule

module XFMB (
    output O,
    input I,
    input PU,
    input PD,
    input SMT
);
endmodule

module BUFJSS (
    output O,
    input I
);
endmodule

module YFA28SB (
    output O,
    input I,
    input E,
    input E2,
    input E4,
    input SR
);
endmodule

module OR2HSS (
    output wire O,
    input wire I1,
    input wire I2
);
endmodule

module AO12JSS (
    output wire O,
    input wire A1,
    input wire B1,
    input wire B2
);
endmodule

module ZFMA28SB (
    inout wire IO,
    output wire O,
    input wire I,
    input wire E,
    input wire E4,
    input wire E2,
    input wire SMT,
    input wire PU,
    input wire PD,
    input wire SR
);
endmodule

module INVHSS (
    output wire O,
    input wire I
);
endmodule
