//NOTE: no-implementation module stub

module REG11LC (
    input wire DSPCLK,
    input wire MMR_web,
    input wire MWORD_we_PSET,
    input wire [10:0] DMD_MW,
    output reg [10:0] MW_OUT,
    input wire RST
);

endmodule
