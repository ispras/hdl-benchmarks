module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 ;
output g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( g17 , n18 );
buf ( g18 , n19 );
buf ( g19 , n20 );
buf ( g20 , n21 );
buf ( g21 , n22 );
buf ( g22 , n23 );
buf ( g23 , n24 );
buf ( g24 , n25 );
buf ( g25 , n26 );
buf ( g26 , n27 );
buf ( g27 , n28 );
buf ( g28 , n29 );
buf ( g29 , n30 );
buf ( g30 , n31 );
buf ( g31 , n32 );
buf ( n18 , n993 );
buf ( n19 , n953 );
buf ( n20 , n971 );
buf ( n21 , n702 );
buf ( n22 , n893 );
buf ( n23 , n800 );
buf ( n24 , n620 );
buf ( n25 , n991 );
buf ( n26 , n991 );
buf ( n27 , n987 );
buf ( n28 , n978 );
buf ( n29 , n405 );
buf ( n30 , n927 );
buf ( n31 , n522 );
buf ( n32 , n867 );
not ( n35 , n13 );
nand ( n36 , n35 , n12 );
not ( n37 , n15 );
nand ( n38 , n37 , n16 );
not ( n39 , n38 );
not ( n40 , n17 );
nand ( n41 , n39 , n40 , n10 );
not ( n42 , n41 );
nor ( n43 , n9 , n11 );
nor ( n44 , n8 , n14 );
nand ( n45 , n43 , n44 );
not ( n46 , n45 );
nand ( n47 , n42 , n46 );
nor ( n48 , n36 , n47 );
nand ( n49 , n48 , n1 );
not ( n50 , n8 );
nor ( n51 , n14 , n11 );
nand ( n52 , n50 , n51 , n9 );
not ( n53 , n52 );
and ( n54 , n16 , n17 );
nor ( n55 , n54 , n15 );
nor ( n56 , n55 , n10 );
and ( n57 , n53 , n56 );
not ( n58 , n1 );
nor ( n59 , n58 , n3 );
buf ( n60 , n59 );
nand ( n61 , n57 , n60 );
and ( n62 , n49 , n61 );
not ( n63 , n5 );
nor ( n64 , n63 , n2 );
not ( n65 , n4 );
nand ( n66 , n64 , n65 );
not ( n67 , n66 );
buf ( n68 , n67 );
not ( n69 , n68 );
nor ( n70 , n62 , n69 );
nor ( n71 , n15 , n16 );
not ( n72 , n14 );
nand ( n73 , n71 , n72 );
not ( n74 , n73 );
nand ( n75 , n74 , n40 );
not ( n76 , n75 );
or ( n77 , n6 , n7 );
not ( n78 , n77 );
nand ( n79 , n76 , n78 );
not ( n80 , n79 );
not ( n81 , n80 );
not ( n82 , n3 );
nor ( n83 , n82 , n1 );
nor ( n84 , n2 , n5 );
and ( n85 , n83 , n84 );
nand ( n86 , n85 , n4 );
not ( n87 , n86 );
not ( n88 , n87 );
or ( n89 , n81 , n88 );
not ( n90 , n15 );
not ( n91 , n16 );
nand ( n92 , n90 , n91 , n72 , n17 );
not ( n93 , n92 );
not ( n94 , n2 );
nand ( n95 , n94 , n4 );
not ( n96 , n5 );
nor ( n97 , n95 , n96 );
not ( n98 , n1 );
nand ( n99 , n97 , n98 );
not ( n100 , n99 );
nand ( n101 , n93 , n100 );
nand ( n102 , n2 , n4 );
not ( n103 , n102 );
and ( n104 , n103 , n5 );
nand ( n105 , n1 , n3 );
buf ( n106 , n105 );
not ( n107 , n106 );
nand ( n108 , n104 , n107 );
and ( n109 , n101 , n108 );
nand ( n110 , n89 , n109 );
nor ( n111 , n70 , n110 );
not ( n112 , n9 );
not ( n113 , n12 );
nand ( n114 , n113 , n13 );
nand ( n115 , n36 , n114 );
nor ( n116 , n10 , n11 );
and ( n117 , n115 , n116 );
not ( n118 , n117 );
not ( n119 , n16 );
nand ( n120 , n119 , n15 );
nor ( n121 , n120 , n40 );
not ( n122 , n121 );
or ( n123 , n118 , n122 );
nand ( n124 , n39 , n17 );
not ( n125 , n124 );
not ( n126 , n13 );
nor ( n127 , n10 , n12 );
nand ( n128 , n126 , n127 );
not ( n129 , n128 );
not ( n130 , n11 );
nand ( n131 , n125 , n129 , n130 );
nand ( n132 , n123 , n131 );
not ( n133 , n132 );
or ( n134 , n112 , n133 );
not ( n135 , n11 );
not ( n136 , n129 );
or ( n137 , n135 , n136 );
nand ( n138 , n12 , n13 );
not ( n139 , n138 );
and ( n140 , n139 , n116 );
not ( n141 , n9 );
nor ( n142 , n140 , n141 );
nand ( n143 , n137 , n142 );
nand ( n144 , n39 , n40 );
not ( n145 , n144 );
nand ( n146 , n143 , n145 );
nand ( n147 , n134 , n146 );
not ( n148 , n4 );
nand ( n149 , n148 , n2 );
not ( n150 , n5 );
nor ( n151 , n149 , n150 );
not ( n152 , n6 );
nand ( n153 , n152 , n8 );
not ( n154 , n153 );
nand ( n155 , n154 , n14 );
not ( n156 , n155 );
and ( n157 , n151 , n156 , n3 );
nand ( n158 , n147 , n157 );
not ( n159 , n45 );
nand ( n160 , n159 , n129 );
not ( n161 , n160 );
nor ( n162 , n1 , n3 );
and ( n163 , n162 , n5 );
and ( n164 , n163 , n78 );
buf ( n165 , n71 );
and ( n166 , n161 , n164 , n165 );
buf ( n167 , n103 );
nand ( n168 , n166 , n167 );
not ( n169 , n14 );
nand ( n170 , n7 , n6 , n8 );
nor ( n171 , n169 , n170 );
not ( n172 , n171 );
not ( n173 , n172 );
not ( n174 , n9 );
nor ( n175 , n174 , n11 );
not ( n176 , n10 );
nor ( n177 , n176 , n8 );
nor ( n178 , n12 , n13 );
nand ( n179 , n175 , n177 , n178 );
not ( n180 , n15 );
not ( n181 , n16 );
nand ( n182 , n180 , n181 );
nand ( n183 , n182 , n72 );
or ( n184 , n179 , n183 );
not ( n185 , n184 );
or ( n186 , n173 , n185 );
not ( n187 , n105 );
and ( n188 , n187 , n4 );
not ( n189 , n188 );
not ( n190 , n5 );
nor ( n191 , n189 , n190 );
nand ( n192 , n186 , n191 );
nand ( n193 , n9 , n14 );
nor ( n194 , n153 , n193 );
not ( n195 , n120 );
and ( n196 , n194 , n195 );
buf ( n197 , n83 );
not ( n198 , n197 );
not ( n199 , n198 );
not ( n200 , n149 );
buf ( n201 , n200 );
nand ( n202 , n196 , n199 , n201 );
and ( n203 , n192 , n202 );
or ( n204 , n99 , n141 );
nand ( n205 , n197 , n64 );
nand ( n206 , n204 , n205 );
not ( n207 , n73 );
not ( n208 , n170 );
and ( n209 , n207 , n208 );
nand ( n210 , n206 , n209 );
nand ( n211 , n158 , n168 , n203 , n210 );
not ( n212 , n2 );
not ( n213 , n17 );
nor ( n214 , n213 , n14 );
not ( n215 , n10 );
nand ( n216 , n214 , n43 , n215 );
nor ( n217 , n8 , n13 );
not ( n218 , n12 );
nand ( n219 , n71 , n217 , n218 );
nor ( n220 , n216 , n219 );
not ( n221 , n7 );
and ( n222 , n220 , n221 );
buf ( n223 , n163 );
nand ( n224 , n222 , n223 );
not ( n225 , n224 );
not ( n226 , n225 );
or ( n227 , n212 , n226 );
or ( n228 , n15 , n16 );
nand ( n229 , n228 , n10 );
or ( n230 , n229 , n45 );
not ( n231 , n230 );
not ( n232 , n15 );
not ( n233 , n17 );
and ( n234 , n232 , n233 );
nor ( n235 , n234 , n128 );
nand ( n236 , n53 , n235 );
not ( n237 , n236 );
or ( n238 , n231 , n237 );
not ( n239 , n197 );
nor ( n240 , n239 , n66 );
nand ( n241 , n238 , n240 );
nor ( n242 , n52 , n55 );
not ( n243 , n127 );
nor ( n244 , n2 , n4 );
nand ( n245 , n59 , n244 );
nor ( n246 , n243 , n245 );
nand ( n247 , n242 , n246 );
nand ( n248 , n241 , n247 );
not ( n249 , n230 );
nand ( n250 , n249 , n60 );
not ( n251 , n95 );
nor ( n252 , n251 , n64 );
nor ( n253 , n250 , n252 );
nor ( n254 , n248 , n253 );
nand ( n255 , n227 , n254 );
nor ( n256 , n211 , n255 );
buf ( n257 , n120 );
nand ( n258 , n124 , n257 );
buf ( n259 , n194 );
nand ( n260 , n258 , n259 );
not ( n261 , n260 );
nand ( n262 , n97 , n197 );
not ( n263 , n262 );
and ( n264 , n261 , n263 );
nand ( n265 , n4 , n5 );
nor ( n266 , n265 , n1 );
nor ( n267 , n2 , n3 );
nand ( n268 , n266 , n267 );
not ( n269 , n268 );
nor ( n270 , n8 , n14 );
not ( n271 , n270 );
nor ( n272 , n271 , n141 );
buf ( n273 , n182 );
and ( n274 , n269 , n272 , n273 );
nor ( n275 , n264 , n274 );
not ( n276 , n7 );
nand ( n277 , n276 , n3 );
nor ( n278 , n277 , n1 );
nand ( n279 , n278 , n17 );
not ( n280 , n279 );
not ( n281 , n2 );
nor ( n282 , n281 , n5 );
buf ( n283 , n282 );
buf ( n284 , n178 );
nand ( n285 , n280 , n46 , n283 , n284 );
not ( n286 , n285 );
nor ( n287 , n144 , n138 );
nand ( n288 , n270 , n141 );
nor ( n289 , n288 , n130 );
not ( n290 , n64 );
nor ( n291 , n106 , n290 );
nand ( n292 , n287 , n289 , n291 );
not ( n293 , n292 );
or ( n294 , n286 , n293 );
nor ( n295 , n4 , n10 );
nand ( n296 , n294 , n295 );
nand ( n297 , n275 , n296 );
nand ( n298 , n200 , n150 );
not ( n299 , n298 );
not ( n300 , n299 );
not ( n301 , n183 );
and ( n302 , n301 , n197 );
not ( n303 , n302 );
not ( n304 , n303 );
not ( n305 , n304 );
or ( n306 , n300 , n305 );
nand ( n307 , n171 , n187 );
not ( n308 , n4 );
nand ( n309 , n308 , n84 );
or ( n310 , n307 , n309 );
nand ( n311 , n306 , n310 );
not ( n312 , n100 );
nand ( n313 , n125 , n259 , n116 );
nor ( n314 , n313 , n139 );
not ( n315 , n314 );
or ( n316 , n312 , n315 );
or ( n317 , n92 , n205 );
nand ( n318 , n316 , n317 );
not ( n319 , n60 );
nor ( n320 , n7 , n15 );
nor ( n321 , n6 , n16 );
not ( n322 , n8 );
nor ( n323 , n322 , n17 , n14 );
nand ( n324 , n320 , n321 , n323 );
nor ( n325 , n319 , n324 , n309 );
nor ( n326 , n297 , n311 , n318 , n325 );
and ( n327 , n111 , n256 , n326 );
buf ( n328 , n162 );
not ( n329 , n328 );
and ( n330 , n145 , n156 );
not ( n331 , n330 );
or ( n332 , n329 , n331 );
not ( n333 , n229 );
nand ( n334 , n333 , n289 , n284 );
not ( n335 , n334 );
nand ( n336 , n335 , n98 );
nand ( n337 , n332 , n336 );
nand ( n338 , n337 , n299 );
and ( n339 , n220 , n7 );
not ( n340 , n3 );
nand ( n341 , n339 , n340 );
not ( n342 , n341 );
not ( n343 , n97 );
buf ( n344 , n343 );
not ( n345 , n344 );
nand ( n346 , n342 , n345 );
and ( n347 , n338 , n346 );
not ( n348 , n167 );
not ( n349 , n335 );
or ( n350 , n348 , n349 );
not ( n351 , n92 );
nand ( n352 , n351 , n201 );
nand ( n353 , n350 , n352 );
nand ( n354 , n353 , n223 );
not ( n355 , n151 );
not ( n356 , n355 );
nand ( n357 , n342 , n356 );
and ( n358 , n354 , n357 );
not ( n359 , n299 );
nand ( n360 , n40 , n162 );
not ( n361 , n360 );
and ( n362 , n361 , n78 );
and ( n363 , n362 , n129 , n46 , n165 );
not ( n364 , n363 );
or ( n365 , n359 , n364 );
not ( n366 , n52 );
not ( n367 , n229 );
nand ( n368 , n366 , n367 );
not ( n369 , n368 );
not ( n370 , n60 );
nand ( n371 , n282 , n4 );
nor ( n372 , n370 , n371 );
nand ( n373 , n369 , n372 );
nand ( n374 , n365 , n373 );
not ( n375 , n114 );
nand ( n376 , n42 , n375 );
nor ( n377 , n376 , n271 );
nand ( n378 , n269 , n377 );
nor ( n379 , n130 , n378 );
nor ( n380 , n374 , n379 );
not ( n381 , n15 );
nand ( n382 , n381 , n16 );
nand ( n383 , n382 , n120 );
nand ( n384 , n156 , n383 );
nor ( n385 , n384 , n198 );
and ( n386 , n385 , n356 );
not ( n387 , n386 );
nor ( n388 , n190 , n4 );
nand ( n389 , n60 , n388 );
or ( n390 , n47 , n389 );
nand ( n391 , n387 , n390 );
not ( n392 , n339 );
not ( n393 , n309 );
and ( n394 , n393 , n1 );
and ( n395 , n107 , n244 );
nor ( n396 , n394 , n395 );
nor ( n397 , n392 , n396 );
nor ( n398 , n391 , n397 );
nand ( n399 , n380 , n398 );
and ( n400 , n339 , n60 );
not ( n401 , n400 );
not ( n402 , n167 );
nor ( n403 , n401 , n402 );
nor ( n404 , n399 , n403 );
nand ( n405 , n327 , n347 , n358 , n404 );
not ( n406 , n184 );
nand ( n407 , n406 , n60 );
not ( n408 , n407 );
nand ( n409 , n190 , n4 );
not ( n410 , n409 );
and ( n411 , n408 , n410 );
not ( n412 , n355 );
not ( n413 , n196 );
not ( n414 , n117 );
nor ( n415 , n413 , n414 );
nand ( n416 , n412 , n415 , n361 );
not ( n417 , n416 );
nor ( n418 , n411 , n417 );
nand ( n419 , n406 , n107 );
not ( n420 , n419 );
not ( n421 , n344 );
and ( n422 , n420 , n421 );
nor ( n423 , n324 , n309 , n3 );
nor ( n424 , n307 , n290 );
nor ( n425 , n423 , n424 );
not ( n426 , n307 );
nand ( n427 , n426 , n244 );
nand ( n428 , n425 , n427 );
nor ( n429 , n422 , n428 );
nand ( n430 , n418 , n429 );
nand ( n431 , n351 , n251 );
not ( n432 , n431 );
nand ( n433 , n432 , n98 );
nand ( n434 , n207 , n78 );
or ( n435 , n434 , n268 );
or ( n436 , n303 , n298 );
nand ( n437 , n435 , n436 );
nor ( n438 , n434 , n86 );
nor ( n439 , n437 , n438 );
nand ( n440 , n433 , n439 );
nor ( n441 , n430 , n440 );
nand ( n442 , n340 , n97 );
nand ( n443 , n396 , n442 );
and ( n444 , n443 , n339 );
and ( n445 , n289 , n287 );
not ( n446 , n66 );
and ( n447 , n446 , n187 );
nand ( n448 , n445 , n447 , n215 );
nand ( n449 , n390 , n448 );
nor ( n450 , n444 , n449 );
and ( n451 , n441 , n354 , n450 );
not ( n452 , n70 );
nand ( n453 , n87 , n53 , n273 , n284 );
nand ( n454 , n452 , n453 );
and ( n455 , n415 , n17 );
and ( n456 , n209 , n141 );
nor ( n457 , n455 , n456 );
nor ( n458 , n457 , n99 );
nor ( n459 , n454 , n458 );
and ( n460 , n44 , n130 );
not ( n461 , n460 );
nor ( n462 , n461 , n229 );
nand ( n463 , n139 , n462 );
not ( n464 , n463 );
nand ( n465 , n367 , n284 );
not ( n466 , n465 );
not ( n467 , n288 );
and ( n468 , n466 , n467 );
buf ( n469 , n42 );
nor ( n470 , n271 , n12 );
and ( n471 , n469 , n470 );
nor ( n472 , n468 , n471 );
not ( n473 , n272 );
not ( n474 , n145 );
or ( n475 , n473 , n474 );
nand ( n476 , n475 , n230 );
not ( n477 , n476 );
nand ( n478 , n53 , n273 , n127 );
and ( n479 , n472 , n477 , n478 );
not ( n480 , n479 );
or ( n481 , n464 , n480 );
nand ( n482 , n481 , n87 );
not ( n483 , n255 );
nand ( n484 , n482 , n483 );
and ( n485 , n2 , n5 );
nand ( n486 , n400 , n485 );
not ( n487 , n486 );
nor ( n488 , n484 , n487 );
not ( n489 , n401 );
not ( n490 , n201 );
not ( n491 , n490 );
and ( n492 , n489 , n491 );
not ( n493 , n147 );
and ( n494 , n151 , n107 );
nand ( n495 , n494 , n156 );
nor ( n496 , n493 , n495 );
not ( n497 , n371 );
and ( n498 , n369 , n497 , n1 );
nor ( n499 , n496 , n498 );
and ( n500 , n166 , n4 );
not ( n501 , n309 );
not ( n502 , n328 );
not ( n503 , n502 );
and ( n504 , n501 , n503 );
nor ( n505 , n371 , n106 );
nor ( n506 , n504 , n505 );
nand ( n507 , n317 , n506 );
nor ( n508 , n500 , n507 );
not ( n509 , n371 );
nand ( n510 , n509 , n3 );
or ( n511 , n510 , n324 );
and ( n512 , n154 , n9 );
not ( n513 , n257 );
nand ( n514 , n299 , n512 , n199 , n513 );
not ( n515 , n262 );
nand ( n516 , n209 , n515 );
nand ( n517 , n511 , n514 , n516 );
not ( n518 , n275 );
nor ( n519 , n517 , n518 );
nand ( n520 , n499 , n508 , n519 );
nor ( n521 , n492 , n520 );
nand ( n522 , n451 , n459 , n488 , n521 );
and ( n523 , n201 , n304 );
buf ( n524 , n301 );
not ( n525 , n524 );
not ( n526 , n104 );
nor ( n527 , n525 , n526 , n277 );
nor ( n528 , n523 , n527 );
nand ( n529 , n196 , n98 );
not ( n530 , n529 );
nand ( n531 , n530 , n299 );
and ( n532 , n84 , n4 );
nand ( n533 , n532 , n3 );
not ( n534 , n533 );
and ( n535 , n42 , n460 );
nand ( n536 , n534 , n535 );
and ( n537 , n528 , n531 , n536 );
nor ( n538 , n47 , n12 );
nor ( n539 , n343 , n98 );
nand ( n540 , n538 , n539 );
buf ( n541 , n196 );
nand ( n542 , n541 , n223 , n167 );
and ( n543 , n540 , n542 , n390 );
nand ( n544 , n537 , n543 , n486 );
not ( n545 , n240 );
nor ( n546 , n545 , n79 );
or ( n547 , n160 , n279 , n355 );
nand ( n548 , n547 , n108 );
nor ( n549 , n546 , n548 );
or ( n550 , n224 , n65 );
nor ( n551 , n368 , n533 );
not ( n552 , n551 );
not ( n553 , n139 );
or ( n554 , n552 , n553 );
nand ( n555 , n554 , n101 );
not ( n556 , n87 );
not ( n557 , n476 );
or ( n558 , n556 , n557 );
nand ( n559 , n377 , n87 );
nand ( n560 , n558 , n559 );
nor ( n561 , n555 , n560 );
not ( n562 , n448 );
nor ( n563 , n250 , n290 );
nor ( n564 , n562 , n563 );
nand ( n565 , n549 , n550 , n561 , n564 );
nand ( n566 , n259 , n39 );
and ( n567 , n92 , n566 );
nor ( n568 , n567 , n298 );
nor ( n569 , n334 , n402 );
nor ( n570 , n568 , n569 );
or ( n571 , n570 , n502 );
and ( n572 , n384 , n324 );
not ( n573 , n199 );
nor ( n574 , n572 , n573 );
nand ( n575 , n497 , n574 );
buf ( n576 , n84 );
buf ( n577 , n576 );
not ( n578 , n577 );
nor ( n579 , n578 , n419 );
nand ( n580 , n406 , n1 );
nor ( n581 , n580 , n95 );
nor ( n582 , n579 , n581 );
nand ( n583 , n571 , n575 , n582 );
nor ( n584 , n544 , n565 , n583 );
not ( n585 , n85 );
nor ( n586 , n585 , n4 );
not ( n587 , n586 );
not ( n588 , n351 );
or ( n589 , n587 , n588 );
buf ( n590 , n220 );
not ( n591 , n278 );
nor ( n592 , n591 , n371 );
nand ( n593 , n590 , n592 );
nand ( n594 , n589 , n593 );
and ( n595 , n188 , n576 );
and ( n596 , n595 , n171 );
nor ( n597 , n594 , n596 );
and ( n598 , n338 , n597 );
not ( n599 , n172 );
not ( n600 , n392 );
or ( n601 , n599 , n600 );
nand ( n602 , n601 , n447 );
not ( n603 , n75 );
nand ( n604 , n603 , n208 );
not ( n605 , n604 );
not ( n606 , n251 );
not ( n607 , n199 );
or ( n608 , n606 , n607 );
nand ( n609 , n608 , n205 );
and ( n610 , n605 , n609 );
nand ( n611 , n369 , n595 );
not ( n612 , n611 );
nor ( n613 , n610 , n612 );
nand ( n614 , n369 , n188 );
or ( n615 , n614 , n2 , n13 );
nand ( n616 , n602 , n613 , n615 );
not ( n617 , n346 );
nor ( n618 , n616 , n617 );
not ( n619 , n454 );
nand ( n620 , n584 , n598 , n618 , n619 );
not ( n621 , n47 );
not ( n622 , n36 );
nand ( n623 , n621 , n447 , n622 );
nor ( n624 , n370 , n298 );
nand ( n625 , n538 , n624 );
nand ( n626 , n535 , n595 );
nand ( n627 , n448 , n626 );
not ( n628 , n627 );
not ( n629 , n4 );
nand ( n630 , n629 , n258 , n512 );
and ( n631 , n92 , n630 );
nor ( n632 , n631 , n585 );
nor ( n633 , n64 , n4 );
not ( n634 , n633 );
not ( n635 , n302 );
or ( n636 , n634 , n635 );
nand ( n637 , n77 , n170 );
nand ( n638 , n207 , n85 , n637 );
nand ( n639 , n636 , n638 );
nor ( n640 , n632 , n639 );
and ( n641 , n623 , n625 , n628 , n640 );
not ( n642 , n336 );
not ( n643 , n298 );
and ( n644 , n642 , n643 );
buf ( n645 , n154 );
not ( n646 , n591 );
not ( n647 , n75 );
and ( n648 , n645 , n646 , n647 );
and ( n649 , n648 , n485 );
nor ( n650 , n644 , n649 );
not ( n651 , n419 );
not ( n652 , n244 );
not ( n653 , n652 );
and ( n654 , n651 , n653 );
and ( n655 , n166 , n2 );
nor ( n656 , n654 , n655 );
nand ( n657 , n641 , n650 , n656 );
not ( n658 , n328 );
nand ( n659 , n658 , n341 );
not ( n660 , n659 );
nor ( n661 , n660 , n69 );
nor ( n662 , n657 , n661 );
and ( n663 , n353 , n328 );
not ( n664 , n663 );
nand ( n665 , n605 , n494 );
and ( n666 , n664 , n665 );
not ( n667 , n407 );
nand ( n668 , n667 , n251 );
not ( n669 , n580 );
nand ( n670 , n669 , n68 );
nand ( n671 , n668 , n670 , n224 );
nand ( n672 , n433 , n427 );
not ( n673 , n85 );
not ( n674 , n335 );
or ( n675 , n673 , n674 );
nor ( n676 , n1 , n17 );
nand ( n677 , n541 , n497 , n676 );
nand ( n678 , n675 , n677 );
and ( n679 , n574 , n167 );
nor ( n680 , n671 , n672 , n678 , n679 );
nor ( n681 , n189 , n2 );
not ( n682 , n681 );
not ( n683 , n538 );
or ( n684 , n682 , n683 );
and ( n685 , n590 , n646 , n190 );
not ( n686 , n576 );
or ( n687 , n686 , n307 );
nand ( n688 , n151 , n383 , n645 , n197 );
nand ( n689 , n687 , n688 );
nor ( n690 , n685 , n689 );
nand ( n691 , n684 , n690 );
and ( n692 , n345 , n339 , n3 );
nor ( n693 , n691 , n692 );
not ( n694 , n604 );
nand ( n695 , n68 , n98 );
not ( n696 , n695 );
and ( n697 , n694 , n696 );
and ( n698 , n222 , n98 , n201 );
nor ( n699 , n697 , n698 );
and ( n700 , n158 , n611 );
and ( n701 , n693 , n699 , n700 );
nand ( n702 , n662 , n666 , n680 , n701 );
not ( n703 , n3 );
not ( n704 , n48 );
or ( n705 , n704 , n69 );
nand ( n706 , n406 , n393 );
nand ( n707 , n705 , n706 );
not ( n708 , n707 );
or ( n709 , n703 , n708 );
not ( n710 , n604 );
nand ( n711 , n244 , n197 );
and ( n712 , n711 , n585 );
not ( n713 , n712 );
and ( n714 , n710 , n713 );
nor ( n715 , n714 , n318 );
nand ( n716 , n709 , n715 );
buf ( n717 , n415 );
nand ( n718 , n717 , n356 , n676 );
nand ( n719 , n550 , n718 );
not ( n720 , n269 );
not ( n721 , n377 );
or ( n722 , n720 , n721 );
and ( n723 , n67 , n59 );
and ( n724 , n532 , n1 );
nor ( n725 , n723 , n724 );
or ( n726 , n184 , n725 );
nand ( n727 , n722 , n726 );
not ( n728 , n727 );
nand ( n729 , n577 , n1 );
or ( n730 , n392 , n729 );
nand ( n731 , n207 , n637 );
or ( n732 , n731 , n268 );
nand ( n733 , n728 , n730 , n732 );
or ( n734 , n392 , n245 );
nor ( n735 , n309 , n3 , n12 );
and ( n736 , n57 , n735 );
and ( n737 , n462 , n269 );
nor ( n738 , n736 , n737 );
and ( n739 , n145 , n251 );
and ( n740 , n273 , n576 );
nor ( n741 , n739 , n740 );
nand ( n742 , n46 , n340 , n1 , n10 );
nor ( n743 , n741 , n742 );
not ( n744 , n743 );
nand ( n745 , n734 , n738 , n744 );
nor ( n746 , n716 , n719 , n733 , n745 );
nor ( n747 , n4 , n5 );
not ( n748 , n747 );
not ( n749 , n337 );
or ( n750 , n748 , n749 );
not ( n751 , n672 );
nand ( n752 , n750 , n751 );
not ( n753 , n16 );
and ( n754 , n217 , n753 , n1 , n7 );
and ( n755 , n43 , n215 );
nor ( n756 , n3 , n5 , n12 , n15 );
and ( n757 , n754 , n755 , n756 , n214 );
nor ( n758 , n752 , n757 );
and ( n759 , n242 , n129 );
nor ( n760 , n759 , n249 );
or ( n761 , n760 , n711 );
or ( n762 , n572 , n510 );
nand ( n763 , n761 , n762 );
not ( n764 , n763 );
and ( n765 , n3 , n251 , n339 );
not ( n766 , n415 );
nor ( n767 , n766 , n99 );
nor ( n768 , n765 , n767 );
nand ( n769 , n764 , n768 );
not ( n770 , n678 );
not ( n771 , n614 );
not ( n772 , n5 );
and ( n773 , n771 , n772 );
not ( n774 , n747 );
or ( n775 , n303 , n774 );
nand ( n776 , n258 , n393 , n512 , n98 );
nand ( n777 , n775 , n776 );
nor ( n778 , n773 , n777 );
not ( n779 , n283 );
nand ( n780 , n779 , n490 );
and ( n781 , n780 , n363 );
and ( n782 , n328 , n747 );
and ( n783 , n782 , n383 , n259 );
nor ( n784 , n781 , n783 );
nand ( n785 , n770 , n778 , n784 );
nor ( n786 , n769 , n785 );
buf ( n787 , n540 );
and ( n788 , n524 , n104 , n646 );
and ( n789 , n72 , n676 );
and ( n790 , n393 , n789 , n78 );
nor ( n791 , n788 , n790 );
and ( n792 , n425 , n791 , n506 );
nand ( n793 , n787 , n792 , n542 );
not ( n794 , n356 );
not ( n795 , n574 );
or ( n796 , n794 , n795 );
not ( n797 , n297 );
nand ( n798 , n796 , n797 );
nor ( n799 , n793 , n798 );
nand ( n800 , n746 , n758 , n786 , n799 );
nand ( n801 , n659 , n244 );
nand ( n802 , n623 , n296 );
not ( n803 , n802 );
not ( n804 , n184 );
nand ( n805 , n67 , n340 );
not ( n806 , n805 );
and ( n807 , n804 , n806 );
not ( n808 , n260 );
and ( n809 , n808 , n782 );
nor ( n810 , n807 , n809 );
nor ( n811 , n4 , n17 );
nand ( n812 , n166 , n811 );
not ( n813 , n431 );
nand ( n814 , n813 , n199 );
nand ( n815 , n810 , n812 , n814 );
not ( n816 , n167 );
not ( n817 , n225 );
or ( n818 , n816 , n817 );
nand ( n819 , n743 , n12 );
nand ( n820 , n818 , n819 );
nor ( n821 , n815 , n820 );
and ( n822 , n801 , n803 , n821 );
nand ( n823 , n648 , n356 );
not ( n824 , n551 );
not ( n825 , n824 );
not ( n826 , n115 );
and ( n827 , n825 , n826 );
not ( n828 , n283 );
not ( n829 , n361 );
or ( n830 , n828 , n829 );
or ( n831 , n360 , n4 );
nand ( n832 , n64 , n162 );
nand ( n833 , n831 , n832 );
nand ( n834 , n833 , n622 , n116 );
nand ( n835 , n830 , n834 );
and ( n836 , n835 , n541 );
nor ( n837 , n827 , n836 );
or ( n838 , n313 , n13 );
or ( n839 , n230 , n218 );
nand ( n840 , n838 , n839 );
not ( n841 , n832 );
nand ( n842 , n840 , n841 );
nand ( n843 , n823 , n837 , n842 );
not ( n844 , n498 );
not ( n845 , n376 );
nand ( n846 , n845 , n289 );
not ( n847 , n846 );
not ( n848 , n79 );
or ( n849 , n847 , n848 );
nand ( n850 , n849 , n841 );
not ( n851 , n409 );
nand ( n852 , n851 , n669 );
and ( n853 , n393 , n637 , n789 );
nor ( n854 , n853 , n505 );
nand ( n855 , n844 , n850 , n852 , n854 );
not ( n856 , n393 );
and ( n857 , n339 , n1 );
not ( n858 , n857 );
or ( n859 , n856 , n858 );
nand ( n860 , n859 , n778 );
nor ( n861 , n843 , n855 , n860 );
nor ( n862 , n479 , n585 );
nor ( n863 , n336 , n774 );
and ( n864 , n605 , n841 , n141 );
nor ( n865 , n862 , n863 , n864 , n692 );
nand ( n866 , n400 , n577 );
nand ( n867 , n822 , n861 , n865 , n866 );
not ( n868 , n515 );
not ( n869 , n335 );
or ( n870 , n868 , n869 );
nand ( n871 , n870 , n625 );
or ( n872 , n407 , n344 );
nand ( n873 , n621 , n595 );
nand ( n874 , n406 , n447 );
nand ( n875 , n872 , n873 , n874 );
or ( n876 , n434 , n1 );
nand ( n877 , n876 , n502 );
and ( n878 , n877 , n68 );
or ( n879 , n711 , n92 );
nand ( n880 , n171 , n281 );
or ( n881 , n880 , n189 );
nand ( n882 , n879 , n881 );
nor ( n883 , n878 , n882 );
nand ( n884 , n574 , n104 );
nand ( n885 , n647 , n87 , n637 );
nand ( n886 , n883 , n884 , n885 );
nor ( n887 , n871 , n875 , n886 );
not ( n888 , n363 );
or ( n889 , n888 , n402 );
nand ( n890 , n222 , n98 , n388 );
nand ( n891 , n889 , n890 );
nor ( n892 , n891 , n496 , n325 );
nand ( n893 , n887 , n664 , n892 , n665 );
not ( n894 , n338 );
or ( n895 , n604 , n545 );
not ( n896 , n497 );
not ( n897 , n896 );
nand ( n898 , n897 , n648 );
nand ( n899 , n895 , n898 );
not ( n900 , n328 );
not ( n901 , n431 );
not ( n902 , n901 );
or ( n903 , n900 , n902 );
or ( n904 , n442 , n47 );
nand ( n905 , n904 , n427 );
nor ( n906 , n905 , n386 );
nand ( n907 , n903 , n906 );
nor ( n908 , n894 , n899 , n907 );
nand ( n909 , n249 , n269 );
and ( n910 , n623 , n296 , n909 );
not ( n911 , n910 );
or ( n912 , n250 , n309 );
not ( n913 , n288 );
nand ( n914 , n845 , n269 , n913 );
nand ( n915 , n912 , n914 );
nor ( n916 , n915 , n437 );
not ( n917 , n109 );
nand ( n918 , n622 , n5 );
nor ( n919 , n614 , n918 );
nor ( n920 , n917 , n919 );
nand ( n921 , n916 , n550 , n920 , n718 );
nor ( n922 , n911 , n921 );
not ( n923 , n457 );
nand ( n924 , n923 , n269 );
and ( n925 , n314 , n269 );
nor ( n926 , n925 , n757 );
nand ( n927 , n908 , n922 , n924 , n926 );
not ( n928 , n311 );
nand ( n929 , n928 , n101 );
nand ( n930 , n665 , n738 );
not ( n931 , n269 );
not ( n932 , n717 );
or ( n933 , n931 , n932 );
nand ( n934 , n933 , n730 );
not ( n935 , n465 );
nand ( n936 , n935 , n532 , n460 , n60 );
or ( n937 , n510 , n384 );
nand ( n938 , n936 , n732 , n506 , n937 );
nor ( n939 , n929 , n930 , n934 , n938 );
nand ( n940 , n744 , n416 );
nor ( n941 , n802 , n940 );
not ( n942 , n419 );
and ( n943 , n942 , n393 );
not ( n944 , n343 );
and ( n945 , n369 , n944 , n107 , n622 );
nor ( n946 , n943 , n945 );
nand ( n947 , n946 , n787 );
not ( n948 , n378 );
nor ( n949 , n948 , n274 );
nand ( n950 , n363 , n747 );
nand ( n951 , n949 , n823 , n950 );
nor ( n952 , n947 , n951 );
nand ( n953 , n939 , n941 , n952 , n926 );
not ( n954 , n87 );
not ( n955 , n605 );
or ( n956 , n954 , n955 );
nand ( n957 , n956 , n597 );
nor ( n958 , n871 , n957 );
not ( n959 , n385 );
nand ( n960 , n646 , n645 , n72 , n40 );
and ( n961 , n959 , n529 , n960 );
nor ( n962 , n961 , n526 );
nor ( n963 , n875 , n962 );
nand ( n964 , n663 , n190 );
not ( n965 , n547 );
or ( n966 , n303 , n355 );
nand ( n967 , n524 , n646 , n485 );
nand ( n968 , n966 , n967 );
nor ( n969 , n896 , n888 );
nor ( n970 , n965 , n968 , n969 , n546 );
nand ( n971 , n958 , n963 , n964 , n970 );
nand ( n972 , n107 , n577 );
nor ( n973 , n392 , n972 );
nor ( n974 , n260 , n414 , n268 );
nor ( n975 , n929 , n973 , n940 , n974 );
nand ( n976 , n400 , n283 );
nand ( n977 , n857 , n532 );
nand ( n978 , n975 , n910 , n976 , n977 );
not ( n979 , n101 );
not ( n980 , n538 );
nand ( n981 , n944 , n107 );
nor ( n982 , n980 , n981 );
nor ( n983 , n979 , n982 );
nand ( n984 , n161 , n280 , n299 );
not ( n985 , n984 );
nor ( n986 , n985 , n311 );
nand ( n987 , n983 , n946 , n986 );
and ( n988 , n385 , n497 );
and ( n989 , n351 , n269 );
nor ( n990 , n988 , n989 );
nand ( n991 , n928 , n990 , n984 );
nand ( n992 , n87 , n57 , n375 );
nand ( n993 , n373 , n992 );
endmodule
