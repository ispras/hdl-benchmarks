module lut_input (in1, in2);
  input in1;
  input in2;
endmodule