module sub_6_2(a, b, c);
  input [5:0] a;
  input [1:0] b;
  output [6:0] c;
  assign c = a - b;
endmodule
