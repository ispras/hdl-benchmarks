module s838_1_bench(
  blif_clk_net,
  blif_reset_net,
  P_0,
  C_32,
  C_31,
  C_30,
  C_29,
  C_28,
  C_27,
  C_26,
  C_25,
  C_24,
  C_23,
  C_22,
  C_21,
  C_20,
  C_19,
  C_18,
  C_17,
  C_16,
  C_15,
  C_14,
  C_13,
  C_12,
  C_11,
  C_10,
  C_9,
  C_8,
  C_7,
  C_6,
  C_5,
  C_4,
  C_3,
  C_2,
  C_1,
  C_0,
  Z);
input blif_clk_net;
input blif_reset_net;
input P_0;
input C_32;
input C_31;
input C_30;
input C_29;
input C_28;
input C_27;
input C_26;
input C_25;
input C_24;
input C_23;
input C_22;
input C_21;
input C_20;
input C_19;
input C_18;
input C_17;
input C_16;
input C_15;
input C_14;
input C_13;
input C_12;
input C_11;
input C_10;
input C_9;
input C_8;
input C_7;
input C_6;
input C_5;
input C_4;
input C_3;
input C_2;
input C_1;
input C_0;
output Z;
reg X_4;
reg X_3;
reg X_2;
reg X_1;
reg X_8;
reg X_7;
reg X_6;
reg X_5;
reg X_12;
reg X_11;
reg X_10;
reg X_9;
reg X_16;
reg X_15;
reg X_14;
reg X_13;
reg X_20;
reg X_19;
reg X_18;
reg X_17;
reg X_24;
reg X_23;
reg X_22;
reg X_21;
reg X_28;
reg X_27;
reg X_26;
reg X_25;
reg X_32;
reg X_31;
reg X_30;
reg X_29;
wire I949;
wire I1_5;
wire I1194;
wire I658_1;
wire P_7;
wire I1155_1;
wire I752;
wire I105_4;
wire I661_1;
wire I701;
wire I1_6;
wire I497_3;
wire I816;
wire I1106;
wire I1061_5;
wire I556;
wire I465_1;
wire I1243;
wire I578_2;
wire I407;
wire I363;
wire I244;
wire I15;
wire I1083_2;
wire I503;
wire I265;
wire P_16;
wire I1218;
wire I799_7;
wire I193_1;
wire I1061_2;
wire I894;
wire I804_4;
wire I442;
wire I480_3;
wire I699;
wire I874;
wire I595_2;
wire I209;
wire I1150;
wire I269_2;
wire I291_1;
wire I865;
wire P_24;
wire I1062_4;
wire I838;
wire I1159_2;
wire I602;
wire I946;
wire I112;
wire P_30;
wire I578_4;
wire I208;
wire I578_1;
wire I804_3;
wire I801_4;
wire I800_7;
wire I269_1;
wire I595_1;
wire I1195;
wire I186_1;
wire I804_5;
wire I661_2;
wire I801_8;
wire I799_8;
wire I803_2;
wire I683_1;
wire I110;
wire I803_1;
wire I809;
wire I636;
wire I462_1;
wire I1083_1;
wire I164;
wire I389_1;
wire P_14;
wire I1151;
wire I802_7;
wire I504;
wire I111;
wire I1123;
wire I358;
wire I203_1;
wire I497_4;
wire P_25;
wire I1061_4;
wire I864;
wire I306;
wire I844;
wire I1062_3;
wire I804_2;
wire I753;
wire I66;
wire I1_4;
wire I563_3;
wire I7_3;
wire I693_1;
wire I441;
wire I367_1;
wire I601;
wire I465_4;
wire I956;
wire I301_1;
wire I676_3;
wire I1203_1;
wire I1079;
wire I246;
wire I947;
wire I836;
wire I1002;
wire I113;
wire I799_5;
wire I342;
wire I872;
wire I776_1;
wire I69;
wire I1103;
wire I800_2;
wire I652;
wire I921;
wire I950;
wire P_1;
wire I364_1;
wire I7_1;
wire I1146;
wire I801_3;
wire P_2;
wire I676_2;
wire I1207_2;
wire I2_7;
wire I693_2;
wire I770_1;
wire I1_3;
wire I1062_6;
wire I1013;
wire I747;
wire I750;
wire I661_3;
wire I171_4;
wire I803_4;
wire I167;
wire I902;
wire I480_1;
wire I284_2;
wire I502;
wire I258;
wire I978;
wire I105_1;
wire I13;
wire I1_2;
wire I168_1;
wire I301_2;
wire I186_3;
wire I1178;
wire I600;
wire P_22;
wire I1222;
wire I88_2;
wire I654;
wire I73_3;
wire I563_4;
wire I367_4;
wire I203_2;
wire I309;
wire I269_4;
wire P_23;
wire I920;
wire I892;
wire I12;
wire P_9;
wire I1087_2;
wire I497_1;
wire I7_2;
wire I1203_2;
wire I505;
wire I1078;
wire I928;
wire I1003;
wire I800_4;
wire I382_3;
wire I1111_2;
wire I1251_1;
wire I799_4;
wire I801_6;
wire I62;
wire I404;
wire I802_6;
wire I171_3;
wire I186_2;
wire I480_2;
wire I751;
wire I1062_5;
wire I637;
wire I595_3;
wire I803_3;
wire I866;
wire I563_1;
wire I770_2;
wire I264;
wire I1251_2;
wire I356;
wire I1130;
wire I269_3;
wire I578_3;
wire I749;
wire I162;
wire I837;
wire I1061_3;
wire I458;
wire I497_2;
wire I676_1;
wire I1087_1;
wire I540;
wire I203_3;
wire I14;
wire I343;
wire I661_4;
wire P_15;
wire I73_4;
wire I465_3;
wire I88_1;
wire I262;
wire I802_2;
wire P_28;
wire I203_4;
wire I1179_2;
wire I308;
wire I1255_2;
wire I835;
wire I987;
wire I846;
wire I650;
wire I2_6;
wire I903;
wire I977;
wire I922;
wire I88_4;
wire I799_3;
wire I211;
wire I959;
wire I2_2;
wire I801_5;
wire I456;
wire I890;
wire I803_5;
wire P_4;
wire I1131_1;
wire I399_4;
wire I147;
wire I1226;
wire P_11;
wire I554;
wire P_20;
wire I806;
wire I1250;
wire I146;
wire I770_3;
wire I563_2;
wire I810;
wire I405;
wire I461;
wire I1242;
wire I1062_8;
wire I700;
wire I382_2;
wire I693_4;
wire I73_1;
wire P_6;
wire I105_3;
wire I1004;
wire I560_1;
wire I367_2;
wire I918;
wire I1247;
wire P_3;
wire I803_6;
wire I1255_1;
wire I160;
wire I307;
wire I171_1;
wire I1159_1;
wire I2_3;
wire I863;
wire I800_6;
wire I284_1;
wire I930;
wire I559;
wire I693_3;
wire I1199;
wire I245;
wire I799_2;
wire I847;
wire I1231_2;
wire I552;
wire I1207_1;
wire I976;
wire I755_1;
wire P_29;
wire I1135_1;
wire I1135_2;
wire I802_3;
wire I802_8;
wire I1155_2;
wire I595_4;
wire I539;
wire I900;
wire I1102;
wire P_21;
wire I1111_1;
wire I367_3;
wire I406;
wire I360;
wire I958;
wire I1062_7;
wire I382_1;
wire I1147;
wire I1_8;
wire I1126;
wire I984;
wire I893;
wire I1014;
wire I399_3;
wire P_13;
wire I105_2;
wire I818;
wire I171_2;
wire I1154;
wire I399_1;
wire I1005;
wire I1223;
wire I800_3;
wire I808;
wire P_26;
wire I758_1;
wire I1122;
wire I487_1;
wire I1062_2;
wire I1061_1;
wire I88_3;
wire I465_2;
wire P_10;
wire I50;
wire I73_2;
wire I803_7;
wire I1006;
wire I399_2;
wire I440;
wire I801_7;
wire I301_3;
wire I538;
wire I480_4;
wire I802_4;
wire I1183_1;
wire I1075;
wire I779_1;
wire I800_8;
wire I1198;
wire I770_4;
wire P_17;
wire I657;
wire I1174;
wire I1107_2;
wire I186_4;
wire I585_1;
wire I1062_9;
wire I737;
wire I975;
wire I49;
wire I64;
wire I1127;
wire I558;
wire I804_6;
wire I260;
wire I382_4;
wire I148;
wire P_31;
wire I1061_7;
wire I1231_1;
wire I931;
wire I948;
wire I301_4;
wire I1227_2;
wire P_18;
wire I1171;
wire I95_1;
wire I284_4;
wire I166;
wire I7_4;
wire I986;
wire I1_7;
wire I1061_8;
wire I1175;
wire I1011;
wire P_8;
wire I801_2;
wire I1107_1;
wire I676_4;
wire I1098;
wire I2_5;
wire I819;
wire I807;
wire I68;
wire I638;
wire I1246;
wire I834;
wire I1074;
wire I891;
wire I799_6;
wire I1131_2;
wire I1183_2;
wire I656;
wire I460;
wire P_27;
wire I362;
wire I802_5;
wire I344;
wire P_12;
wire I875;
wire I1170;
wire I736;
wire I2_4;
wire I919;
wire I1061_6;
wire I210;
wire I70_1;
wire I804_7;
wire I454;
wire I1179_1;
wire I1219;
wire I800_5;
wire I284_3;
wire I2_1;
wire I266_1;
wire I1227_1;
wire P_32;
wire I1099;
wire I1082;
wire I1202;
wire I603;
wire I698;
wire P_19;
wire P_5;
wire I974;
wire I862;
wire I48;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_4 <= 0;
  else
    X_4 <= I12;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_3 <= 0;
  else
    X_3 <= I13;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_2 <= 0;
  else
    X_2 <= I14;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_1 <= 0;
  else
    X_1 <= I15;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_8 <= 0;
  else
    X_8 <= I110;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_7 <= 0;
  else
    X_7 <= I111;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_6 <= 0;
  else
    X_6 <= I112;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_5 <= 0;
  else
    X_5 <= I113;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_12 <= 0;
  else
    X_12 <= I208;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_11 <= 0;
  else
    X_11 <= I209;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_10 <= 0;
  else
    X_10 <= I210;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_9 <= 0;
  else
    X_9 <= I211;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_16 <= 0;
  else
    X_16 <= I306;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_15 <= 0;
  else
    X_15 <= I307;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_14 <= 0;
  else
    X_14 <= I308;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_13 <= 0;
  else
    X_13 <= I309;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_20 <= 0;
  else
    X_20 <= I404;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_19 <= 0;
  else
    X_19 <= I405;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_18 <= 0;
  else
    X_18 <= I406;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_17 <= 0;
  else
    X_17 <= I407;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_24 <= 0;
  else
    X_24 <= I502;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_23 <= 0;
  else
    X_23 <= I503;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_22 <= 0;
  else
    X_22 <= I504;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_21 <= 0;
  else
    X_21 <= I505;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_28 <= 0;
  else
    X_28 <= I600;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_27 <= 0;
  else
    X_27 <= I601;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_26 <= 0;
  else
    X_26 <= I602;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_25 <= 0;
  else
    X_25 <= I603;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_32 <= 0;
  else
    X_32 <= I698;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_31 <= 0;
  else
    X_31 <= I699;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_30 <= 0;
  else
    X_30 <= I700;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    X_29 <= 0;
  else
    X_29 <= I701;
assign I465_3 = (I461&I465_2);
assign I949 = ((~X_23));
assign I1_5 = (I2_4&I1_4);
assign I1194 = ((~P_22));
assign I262 = ((~X_9))|((~I1_3));
assign I88_1 = ((~X_1));
assign P_28 = (I804_6&I802_7);
assign I802_2 = ((~X_7)&(~I844)&(~I838));
assign I1179_2 = (I1170)|(I1174);
assign I203_4 = (X_10&I203_1);
assign I658_1 = (I656)|(X_28)|(I638);
assign P_7 = (I803_1&I801_2);
assign I308 = ((~I301_3)&(~I301_4));
assign I1155_1 = (I1147)|(I1151);
assign I1255_2 = (P_28&C_28);
assign I752 = ((~I751));
assign I835 = ((~X_5));
assign I987 = ((~I986));
assign I105_4 = (X_6&I105_1);
assign I661_1 = ((~I657));
assign I701 = (I770_3)|(I770_4);
assign I1_6 = (I2_5&I1_5);
assign I846 = ((~I835))|((~P_0));
assign I650 = ((~I683_1))|((~X_28));
assign I497_3 = (I556&I497_2);
assign I816 = ((~I819))|((~I808));
assign I2_6 = ((~I554)&(~I539)&(~I540));
assign I903 = ((~I902));
assign I1106 = ((~I1111_1)&(~I1111_2));
assign I1061_5 = ((~I1179_1))|((~I1179_2))|((~I1178));
assign I977 = ((~X_27));
assign I556 = ((~X_21))|((~I1_6));
assign I465_1 = ((~I461));
assign I922 = ((~X_20));
assign I88_4 = (P_0&I88_1);
assign I799_3 = ((~I862)&(~I863));
assign I1243 = ((~P_31));
assign I578_2 = ((~I1_6));
assign I211 = (I284_3)|(I284_4);
assign I959 = ((~I958));
assign I407 = (I480_3)|(I480_4);
assign I363 = ((~I358)&(~I342));
assign I2_2 = ((~I162)&(~I147)&(~I148));
assign I244 = ((~I1_3));
assign I15 = (I88_3)|(I88_4);
assign I801_5 = ((~I921)&(~I928));
assign I456 = ((~X_17))|((~X_18));
assign I1083_2 = (I1074)|(I1078);
assign I803_5 = ((~X_20)&(~X_18)&(~X_19)&(~X_17));
assign I890 = ((~P_0));
assign I503 = (I563_3)|(I563_4);
assign I1131_1 = (I1123)|(I1127);
assign P_4 = ((~X_3)&(~I816)&(~I810));
assign I399_4 = (X_18&I399_1);
assign I147 = ((~X_8));
assign I1226 = ((~I1231_1)&(~I1231_2));
assign I265 = ((~I260)&(~I244));
assign P_16 = (I804_3&I802_4);
assign P_11 = (I804_2&I801_3);
assign I554 = ((~X_21))|((~X_22));
assign I1218 = ((~P_26));
assign I799_7 = ((~I974)&(~I975));
assign Z = (I1062_8)|(I1062_9);
assign I193_1 = (I162)|(I148)|(I146);
assign P_20 = (I804_4&I802_5);
assign I1250 = ((~I1255_1)&(~I1255_2));
assign I806 = ((~P_0));
assign I1061_2 = ((~I1107_1))|((~I1107_2))|((~I1106));
assign I894 = ((~X_16));
assign I146 = ((~I1_2));
assign I804_4 = (I804_3&I803_4);
assign I770_3 = (X_29&I770_2);
assign I480_3 = (X_17&I480_2);
assign I810 = ((~X_4));
assign I563_2 = ((~X_23));
assign I442 = ((~X_19));
assign I1242 = ((~P_30));
assign I461 = ((~I456)&(~I440));
assign I405 = (I465_3)|(I465_4);
assign I1062_8 = (I1062_7)|(I1061_8);
assign I699 = ((~I758_1))|((~I749));
assign I382_2 = ((~I1_4));
assign I700 = ((~I693_3)&(~I693_4));
assign I693_4 = (X_30&I693_1);
assign I874 = ((~I863))|((~P_0));
assign I595_2 = ((~X_26));
assign I209 = (I269_3)|(I269_4);
assign I1150 = ((~C_14));
assign I269_2 = ((~X_11));
assign I73_1 = ((~I69));
assign I291_1 = (I260)|(I246)|(I244);
assign P_6 = (I803_1&I800_2);
assign I865 = ((~X_11));
assign I105_3 = (I164&I105_2);
assign P_24 = (I804_5&I802_6);
assign I1062_4 = (I1062_3)|(I1061_4);
assign I838 = ((~X_8));
assign I1004 = ((~X_30));
assign I1159_2 = (P_12&C_12);
assign I602 = ((~I595_3)&(~I595_4));
assign I560_1 = (I558)|(X_24)|(I540);
assign I946 = ((~P_0));
assign I367_2 = ((~X_15));
assign I918 = ((~P_0));
assign I112 = ((~I105_3)&(~I105_4));
assign I1247 = ((~C_31));
assign I578_4 = (I1_6&I578_1);
assign P_30 = (I804_7&I800_8);
assign I803_6 = ((~X_24)&(~X_22)&(~X_23)&(~X_21));
assign P_3 = ((~I809)&(~I816));
assign I1255_1 = (P_29&C_29);
assign I208 = ((~I266_1))|((~I258));
assign I160 = ((~I193_1))|((~X_8));
assign I307 = (I367_3)|(I367_4);
assign I171_1 = ((~I167));
assign I1159_1 = (P_13&C_13);
assign I578_1 = ((~X_21));
assign I804_3 = (I804_2&I803_3);
assign I801_4 = ((~I893)&(~I900));
assign I2_3 = ((~I260)&(~I245)&(~I246));
assign I863 = ((~X_9));
assign I800_7 = ((~I976)&(~I986));
assign I800_6 = ((~I948)&(~I958));
assign I269_1 = ((~I265));
assign I595_1 = ((~I654));
assign I930 = ((~I919))|((~P_0));
assign I284_1 = ((~X_9));
assign I1195 = ((~P_23));
assign I186_1 = ((~X_5));
assign I559 = ((~I554)&(~I538));
assign I693_3 = (I751&I693_2);
assign I1199 = ((~C_23));
assign I245 = ((~X_12));
assign I804_5 = (I804_4&I803_5);
assign I799_2 = ((~I834)&(~I835));
assign I1231_2 = (P_24&C_24);
assign I847 = ((~I846));
assign I661_2 = ((~X_27));
assign I801_8 = ((~I1005)&(~I1011));
assign I799_8 = ((~I1002)&(~I1003));
assign I803_2 = ((~X_8)&(~X_6)&(~X_7)&(~X_5));
assign I552 = ((~I585_1))|((~X_24));
assign I683_1 = (I652)|(I638)|(I636);
assign I1207_1 = (P_21&C_21);
assign I110 = ((~I168_1))|((~I160));
assign I803_1 = ((~X_4)&(~X_2)&(~X_3)&(~X_1));
assign I976 = ((~X_26));
assign I809 = ((~X_3));
assign I636 = ((~I1_7));
assign I755_1 = (I753)|(X_32)|(I736);
assign I462_1 = (I460)|(X_20)|(I442);
assign P_29 = (I804_7&I799_8);
assign I1083_1 = (I1075)|(I1079);
assign I1135_1 = (P_9&C_9);
assign I1135_2 = (P_8&C_8);
assign I802_8 = ((~X_31)&(~I1011)&(~I1006));
assign I802_3 = ((~X_11)&(~I872)&(~I866));
assign I164 = ((~X_5))|((~I1_2));
assign I389_1 = (I358)|(I344)|(I342);
assign I1155_2 = (I1146)|(I1150);
assign P_14 = (I804_3&I800_4);
assign I1151 = ((~C_15));
assign I900 = ((~I903))|((~I892));
assign I802_7 = ((~X_27)&(~I984)&(~I978));
assign I595_4 = (X_26&I595_1);
assign I539 = ((~X_24));
assign I504 = ((~I497_3)&(~I497_4));
assign I1102 = ((~C_6));
assign I111 = (I171_3)|(I171_4);
assign I1123 = ((~P_11));
assign P_21 = (I804_5&I799_6);
assign I1111_1 = (P_5&C_5);
assign I358 = ((~X_13))|((~X_14));
assign I367_3 = (I363&I367_2);
assign I203_1 = ((~I262));
assign I406 = ((~I399_3)&(~I399_4));
assign I1062_7 = (I1062_6)|(I1061_7);
assign I958 = ((~I947))|((~P_0));
assign I360 = ((~X_13))|((~I1_4));
assign I497_4 = (X_22&I497_1);
assign I1147 = ((~P_15));
assign I382_1 = ((~X_13));
assign P_25 = (I804_6&I799_7);
assign I1061_4 = ((~I1155_1))|((~I1155_2))|((~I1154));
assign I984 = ((~I987))|((~I976));
assign I1126 = ((~C_10));
assign I1_8 = (I2_7&I1_7);
assign I893 = ((~X_15));
assign I864 = ((~X_10));
assign I1014 = ((~I1013));
assign I306 = ((~I364_1))|((~I356));
assign I844 = ((~I847))|((~I836));
assign P_13 = (I804_3&I799_4);
assign I399_3 = (I458&I399_2);
assign I818 = ((~I807))|((~P_0));
assign I105_2 = ((~X_6));
assign I1062_3 = (I1062_2)|(I1061_3);
assign I804_2 = (I803_1&I803_2);
assign I753 = ((~I752))|((~X_30));
assign I66 = ((~X_1))|((~P_0));
assign I1154 = ((~I1159_1)&(~I1159_2));
assign I563_3 = (I559&I563_2);
assign I171_2 = ((~X_7));
assign I1_4 = (I2_3&I1_3);
assign I7_3 = (I66&I7_2);
assign I693_1 = ((~I751));
assign I1005 = ((~X_31));
assign I399_1 = ((~I458));
assign I367_1 = ((~I363));
assign I441 = ((~X_20));
assign I601 = (I661_3)|(I661_4);
assign I465_4 = (X_19&I465_1);
assign I1223 = ((~C_27));
assign I800_3 = ((~I864)&(~I874));
assign I956 = ((~I959))|((~I948));
assign I301_1 = ((~I360));
assign I676_3 = (X_25&I676_2);
assign I1203_1 = (I1195)|(I1199);
assign I808 = ((~X_2));
assign P_26 = (I804_6&I800_7);
assign I758_1 = (I753)|(X_31);
assign I487_1 = (I456)|(I442)|(I440);
assign I1122 = ((~P_10));
assign I1062_2 = (I1061_1)|(I1061_2);
assign I1079 = ((~C_3));
assign I246 = ((~X_11));
assign I1061_1 = ((~I1083_1))|((~I1083_2))|((~I1082));
assign I88_3 = (X_1&I88_2);
assign I465_2 = ((~X_19));
assign I947 = ((~X_21));
assign I836 = ((~X_6));
assign I113 = (I186_3)|(I186_4);
assign I1002 = ((~P_0));
assign I799_5 = ((~I918)&(~I919));
assign I342 = ((~I1_4));
assign P_10 = (I804_2&I800_3);
assign I872 = ((~I875))|((~I864));
assign I50 = ((~X_3));
assign I776_1 = (I751)|(I737)|(I736);
assign I69 = ((~I64)&(~I48));
assign I803_7 = ((~X_28)&(~X_26)&(~X_27)&(~X_25));
assign I73_2 = ((~X_3));
assign I1006 = ((~X_32));
assign I1103 = ((~C_7));
assign I801_7 = ((~I977)&(~I984));
assign I399_2 = ((~X_18));
assign I440 = ((~I1_5));
assign I652 = ((~X_25))|((~X_26));
assign I800_2 = ((~I836)&(~I846));
assign I921 = ((~X_19));
assign I301_3 = (I360&I301_2);
assign I950 = ((~X_24));
assign I1183_1 = (P_17&C_17);
assign P_1 = ((~I806)&(~I807));
assign I802_4 = ((~X_15)&(~I900)&(~I894));
assign I480_4 = (I1_5&I480_1);
assign I538 = ((~I1_6));
assign I1075 = ((~P_3));
assign I364_1 = (I362)|(X_16)|(I344);
assign I779_1 = (I752&X_30);
assign I800_8 = ((~I1004)&(~I1013));
assign I7_1 = ((~I66));
assign I801_3 = ((~I865)&(~I872));
assign I1146 = ((~P_14));
assign I1198 = ((~C_22));
assign I770_4 = (I1_8&I770_1);
assign P_2 = ((~I808)&(~I818));
assign P_17 = (I804_4&I799_5);
assign I657 = ((~I652)&(~I636));
assign I1174 = ((~C_18));
assign I1107_2 = (I1098)|(I1102);
assign I585_1 = (I554)|(I540)|(I538);
assign I186_4 = (I1_2&I186_1);
assign I1062_9 = (P_32&C_32);
assign I676_2 = ((~I1_7));
assign I737 = ((~X_30));
assign I1207_2 = (P_20&C_20);
assign I2_7 = ((~I652)&(~I637)&(~I638));
assign I693_2 = ((~X_30));
assign I1_3 = (I2_2&I1_2);
assign I770_1 = ((~X_29));
assign I975 = ((~X_25));
assign I49 = ((~X_4));
assign I747 = ((~I776_1))|((~X_32));
assign I1062_6 = (I1062_5)|(I1061_6);
assign I1013 = ((~I1003))|((~P_0));
assign I64 = ((~X_1))|((~X_2));
assign I661_3 = (I657&I661_2);
assign I750 = ((~I736)&(~I779_1));
assign I1127 = ((~C_11));
assign I171_4 = (X_7&I171_1);
assign I804_6 = (I804_5&I803_6);
assign I803_4 = ((~X_16)&(~X_14)&(~X_15)&(~X_13));
assign I167 = ((~I162)&(~I146));
assign I558 = ((~I559));
assign I260 = ((~X_9))|((~X_10));
assign I382_4 = (I1_4&I382_1);
assign I148 = ((~X_7));
assign I1061_7 = ((~I1227_1))|((~I1227_2))|((~I1226));
assign I902 = ((~I891))|((~P_0));
assign P_31 = (I804_7&I801_8);
assign I480_1 = ((~X_17));
assign I1231_1 = (P_25&C_25);
assign I284_2 = ((~I1_3));
assign I931 = ((~I930));
assign I258 = ((~I291_1))|((~X_12));
assign I502 = ((~I560_1))|((~I552));
assign I948 = ((~X_22));
assign I1227_2 = (I1218)|(I1222);
assign I301_4 = (X_14&I301_1);
assign P_18 = (I804_4&I800_5);
assign I1171 = ((~P_19));
assign I105_1 = ((~I164));
assign I978 = ((~X_28));
assign I95_1 = (I64)|(I50)|(I48);
assign I1_2 = (I2_1&P_0);
assign I13 = (I73_3)|(I73_4);
assign I284_4 = (I1_3&I284_1);
assign I168_1 = (I166)|(X_8)|(I148);
assign I166 = ((~I167));
assign I301_2 = ((~X_14));
assign I186_3 = (X_5&I186_2);
assign I1178 = ((~I1183_1)&(~I1183_2));
assign I600 = ((~I658_1))|((~I650));
assign I7_4 = (X_2&I7_1);
assign P_22 = (I804_5&I800_6);
assign I88_2 = ((~P_0));
assign I1222 = ((~C_26));
assign I654 = ((~X_25))|((~I1_7));
assign I986 = ((~I975))|((~P_0));
assign I563_4 = (X_23&I563_1);
assign I73_3 = (I69&I73_2);
assign I1_7 = (I2_6&I1_6);
assign I1061_8 = ((~I1251_1))|((~I1251_2))|((~I1250));
assign I367_4 = (X_15&I367_1);
assign I203_2 = ((~X_10));
assign I309 = (I382_3)|(I382_4);
assign I269_4 = (X_11&I269_1);
assign I892 = ((~X_14));
assign I920 = ((~X_18));
assign P_23 = (I804_5&I801_6);
assign I12 = ((~I70_1))|((~I62));
assign P_9 = (I804_2&I799_3);
assign I1175 = ((~C_19));
assign I1087_2 = (P_0&C_0);
assign I1011 = ((~I1014))|((~I1004));
assign I497_1 = ((~I556));
assign P_8 = (I803_1&I802_2);
assign I7_2 = ((~X_2));
assign I1203_2 = (I1194)|(I1198);
assign I801_2 = ((~I837)&(~I844));
assign I1107_1 = (I1099)|(I1103);
assign I505 = (I578_3)|(I578_4);
assign I1078 = ((~C_2));
assign I676_4 = (I1_7&I676_1);
assign I928 = ((~I931))|((~I920));
assign I1098 = ((~P_6));
assign I1003 = ((~X_29));
assign I2_5 = ((~I456)&(~I441)&(~I442));
assign I819 = ((~I818));
assign I800_4 = ((~I892)&(~I902));
assign I807 = ((~X_1));
assign I382_3 = (X_13&I382_2);
assign I638 = ((~X_27));
assign I68 = ((~I69));
assign I1246 = ((~C_30));
assign I834 = ((~P_0));
assign I1074 = ((~P_2));
assign I891 = ((~X_13));
assign I1131_2 = (I1122)|(I1126);
assign I1111_2 = (P_4&C_4);
assign I799_6 = ((~I946)&(~I947));
assign I1251_1 = (I1243)|(I1247);
assign I1183_2 = (P_16&C_16);
assign I799_4 = ((~I890)&(~I891));
assign I656 = ((~I657));
assign I801_6 = ((~I949)&(~I956));
assign I460 = ((~I461));
assign P_27 = (I804_6&I801_7);
assign I362 = ((~I363));
assign I62 = ((~I95_1))|((~X_4));
assign I404 = ((~I462_1))|((~I454));
assign I802_6 = ((~X_23)&(~I956)&(~I950));
assign I802_5 = ((~X_19)&(~I928)&(~I922));
assign I171_3 = (I167&I171_2);
assign I344 = ((~X_15));
assign P_12 = (I804_2&I802_3);
assign I186_2 = ((~I1_2));
assign I480_2 = ((~I1_5));
assign I875 = ((~I874));
assign I1170 = ((~P_18));
assign I751 = ((~X_29))|((~I1_8));
assign I1062_5 = (I1062_4)|(I1061_5);
assign I736 = ((~X_31));
assign I637 = ((~X_28));
assign I595_3 = (I654&I595_2);
assign I803_3 = ((~X_12)&(~X_10)&(~X_11)&(~X_9));
assign I2_4 = ((~I358)&(~I343)&(~I344));
assign I866 = ((~X_12));
assign I919 = ((~X_17));
assign I1061_6 = ((~I1203_1))|((~I1203_2))|((~I1202));
assign I563_1 = ((~I559));
assign I210 = ((~I203_3)&(~I203_4));
assign I70_1 = (I68)|(X_4)|(I50);
assign I770_2 = ((~I1_8));
assign I264 = ((~I265));
assign I804_7 = (I804_6&I803_7);
assign I454 = ((~I487_1))|((~X_20));
assign I1251_2 = (I1242)|(I1246);
assign I1179_1 = (I1171)|(I1175);
assign I356 = ((~I389_1))|((~X_16));
assign I1219 = ((~P_27));
assign I1130 = ((~I1135_1)&(~I1135_2));
assign I800_5 = ((~I920)&(~I930));
assign I578_3 = (X_21&I578_2);
assign I269_3 = (I265&I269_2);
assign I162 = ((~X_5))|((~X_6));
assign I749 = ((~I750));
assign I284_3 = (X_9&I284_2);
assign I1227_1 = (I1219)|(I1223);
assign I266_1 = (I264)|(X_12)|(I246);
assign I2_1 = ((~I64)&(~I49)&(~I50));
assign P_32 = (I804_7&I802_8);
assign I837 = ((~X_7));
assign I1061_3 = ((~I1131_1))|((~I1131_2))|((~I1130));
assign I497_2 = ((~X_22));
assign I458 = ((~X_17))|((~I1_5));
assign I1082 = ((~I1087_1)&(~I1087_2));
assign I676_1 = ((~X_25));
assign I1099 = ((~P_7));
assign I1202 = ((~I1207_1)&(~I1207_2));
assign I603 = (I676_3)|(I676_4);
assign I1087_1 = (P_1&C_1);
assign I540 = ((~X_23));
assign I203_3 = (I262&I203_2);
assign I14 = ((~I7_3)&(~I7_4));
assign I343 = ((~X_16));
assign I698 = ((~I755_1))|((~I747));
assign P_5 = (I803_1&I799_2);
assign I661_4 = (X_27&I661_1);
assign P_19 = (I804_4&I801_5);
assign I974 = ((~P_0));
assign I862 = ((~P_0));
assign P_15 = (I804_3&I801_4);
assign I73_4 = (X_3&I73_1);
assign I48 = ((~P_0));
endmodule
