module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 ;
output n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
 n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
 n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
 n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
 n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
 n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
 n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
 n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
 n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
 n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
 n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
 n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
 n220 , n221 , n222 , n223 , n224 , n225 , n226 ;
wire n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , 
 n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , 
 n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , 
 n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , 
 n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , 
 n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , 
 n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , 
 n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , 
 n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , 
 n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , 
 n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , 
 n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , 
 n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , 
 n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , 
 n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , 
 n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , 
 n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , 
 n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , 
 n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , 
 n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , 
 n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , 
 n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , 
 n675 , n676 , n677 , n678 , n679 , n680 , n29489 , n29490 , n29491 , n29492 , 
 n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , 
 n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , 
 n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , 
 n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , 
 n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , 
 n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , 
 n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , 
 n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , 
 n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , 
 n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , 
 n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , 
 n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , 
 n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , 
 n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , 
 n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , 
 n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , 
 n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , 
 n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , 
 n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , 
 n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , 
 n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , 
 n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , 
 n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , 
 n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , 
 n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , 
 n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , 
 n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , 
 n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , 
 n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , 
 n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , 
 n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , 
 n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , 
 n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , 
 n29823 , n29824 , n684 , n29826 , n686 , n687 , n29829 , n29830 , n690 , n29832 , 
 n29833 , n693 , n29835 , n695 , n29837 , n29838 , n698 , n29840 , n29841 , n701 , 
 n29843 , n703 , n29845 , n29846 , n29847 , n707 , n29849 , n29850 , n29851 , n29852 , 
 n29853 , n29854 , n714 , n29856 , n716 , n717 , n718 , n719 , n720 , n721 , 
 n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , 
 n732 , n733 , n734 , n735 , n736 , n29878 , n741 , n29880 , n743 , n29882 , 
 n745 , n29884 , n29885 , n748 , n29887 , n750 , n29889 , n752 , n29891 , n29892 , 
 n758 , n29894 , n29895 , n761 , n29897 , n763 , n29899 , n765 , n29901 , n770 , 
 n29903 , n772 , n29905 , n29906 , n775 , n776 , n777 , n778 , n782 , n29912 , 
 n784 , n29914 , n786 , n29916 , n788 , n789 , n790 , n791 , n29921 , n29922 , 
 n29923 , n795 , n29925 , n797 , n798 , n799 , n29929 , n801 , n29931 , n29932 , 
 n804 , n29934 , n29935 , n807 , n29937 , n29938 , n29939 , n29940 , n815 , n29942 , 
 n29943 , n818 , n29945 , n29946 , n29947 , n822 , n29949 , n824 , n29951 , n29952 , 
 n827 , n29954 , n29955 , n830 , n29957 , n832 , n833 , n834 , n29961 , n29962 , 
 n29963 , n29964 , n842 , n29966 , n29967 , n845 , n29969 , n29970 , n848 , n29972 , 
 n850 , n851 , n852 , n29976 , n854 , n29978 , n856 , n857 , n29981 , n859 , 
 n29983 , n29984 , n29985 , n863 , n29987 , n29988 , n869 , n29990 , n29991 , n872 , 
 n29993 , n29994 , n875 , n876 , n29997 , n878 , n879 , n30000 , n881 , n882 , 
 n30003 , n884 , n885 , n30006 , n887 , n30008 , n30009 , n30010 , n891 , n30012 , 
 n30013 , n894 , n30015 , n30016 , n30017 , n898 , n30019 , n30020 , n901 , n30022 , 
 n30023 , n904 , n30025 , n30026 , n907 , n30028 , n909 , n910 , n30031 , n30032 , 
 n30033 , n30034 , n30035 , n919 , n30037 , n30038 , n922 , n30040 , n30041 , n925 , 
 n926 , n927 , n928 , n929 , n30047 , n931 , n932 , n933 , n30051 , n30052 , 
 n936 , n30054 , n30055 , n939 , n30057 , n30058 , n942 , n30060 , n30061 , n945 , 
 n30063 , n30064 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n30072 , 
 n959 , n960 , n961 , n30076 , n963 , n30078 , n30079 , n966 , n30081 , n30082 , 
 n969 , n970 , n971 , n972 , n973 , n30088 , n975 , n30090 , n30091 , n978 , 
 n979 , n30094 , n981 , n30096 , n30097 , n984 , n30099 , n986 , n30101 , n30102 , 
 n989 , n30104 , n30105 , n30106 , n996 , n30108 , n998 , n30110 , n1000 , n1001 , 
 n30113 , n30114 , n1004 , n30116 , n30117 , n1007 , n30119 , n30120 , n1010 , n30122 , 
 n1012 , n30124 , n30125 , n1015 , n30127 , n30128 , n1018 , n30130 , n30131 , n1024 , 
 n30133 , n30134 , n1027 , n1028 , n30137 , n1030 , n30139 , n30140 , n30141 , n30142 , 
 n1035 , n30144 , n30145 , n1038 , n1039 , n30148 , n1041 , n30150 , n30151 , n30152 , 
 n1045 , n30154 , n30155 , n1048 , n30157 , n30158 , n30159 , n1052 , n30161 , n1054 , 
 n30163 , n1056 , n30165 , n1058 , n1059 , n30168 , n1061 , n30170 , n30171 , n30172 , 
 n1065 , n30174 , n30175 , n1068 , n30177 , n30178 , n30179 , n30180 , n1073 , n1074 , 
 n30183 , n30184 , n1077 , n30186 , n30187 , n1080 , n30189 , n1085 , n30191 , n30192 , 
 n1088 , n1089 , n1090 , n1091 , n30197 , n1093 , n1094 , n1095 , n1096 , n1097 , 
 n1098 , n1099 , n30205 , n30206 , n1102 , n30208 , n30209 , n1105 , n30211 , n1107 , 
 n1108 , n30214 , n1110 , n30216 , n1112 , n1113 , n30219 , n30220 , n1116 , n30222 , 
 n30223 , n1119 , n30225 , n30226 , n30227 , n1126 , n30229 , n30230 , n1129 , n30232 , 
 n1131 , n30234 , n1133 , n30236 , n1135 , n30238 , n30239 , n1138 , n30241 , n1140 , 
 n1141 , n30244 , n1143 , n30246 , n30247 , n30248 , n1147 , n30250 , n30251 , n1150 , 
 n30253 , n30254 , n30255 , n1154 , n30257 , n30258 , n1157 , n30260 , n1159 , n1160 , 
 n1161 , n1162 , n1163 , n30266 , n30267 , n1166 , n30269 , n1168 , n30271 , n30272 , 
 n30273 , n30274 , n1173 , n30276 , n1175 , n30278 , n30279 , n1178 , n30281 , n30282 , 
 n30283 , n1182 , n30285 , n1187 , n30287 , n1189 , n1190 , n30290 , n30291 , n1193 , 
 n30293 , n30294 , n1196 , n30296 , n30297 , n1199 , n1200 , n30300 , n30301 , n1203 , 
 n30303 , n30304 , n1206 , n30306 , n30307 , n1209 , n30309 , n30310 , n1212 , n30312 , 
 n30313 , n1215 , n1216 , n30316 , n1221 , n1222 , n30319 , n30320 , n1225 , n1226 , 
 n30323 , n30324 , n1229 , n30326 , n30327 , n1232 , n30329 , n1234 , n1235 , n30332 , 
 n30333 , n30334 , n1239 , n1240 , n30337 , n30338 , n1243 , n30340 , n30341 , n1246 , 
 n30343 , n1248 , n30345 , n1250 , n30347 , n1252 , n1253 , n1254 , n1255 , n30352 , 
 n1257 , n30354 , n1259 , n1260 , n30357 , n30358 , n1263 , n30360 , n30361 , n1266 , 
 n30363 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , 
 n30373 , n30374 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , 
 n1287 , n1288 , n1289 , n1290 , n1291 , n30388 , n1293 , n30390 , n30391 , n1296 , 
 n30393 , n30394 , n1299 , n30396 , n1301 , n1302 , n1303 , n1304 , n1305 , n1309 , 
 n30403 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n30411 , n1319 , 
 n30413 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
 n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n30429 , n1337 , n30431 , n30432 , 
 n1343 , n1344 , n1345 , n30436 , n30437 , n30438 , n1349 , n1350 , n1351 , n1352 , 
 n1353 , n1354 , n1355 , n1356 , n30447 , n30448 , n1359 , n30450 , n30451 , n1362 , 
 n30453 , n30454 , n1365 , n1366 , n30457 , n30458 , n30459 , n1370 , n30461 , n30462 , 
 n1373 , n30464 , n30465 , n1376 , n30467 , n30468 , n30469 , n30470 , n30471 , n1382 , 
 n30473 , n30474 , n1385 , n30476 , n30477 , n1388 , n1389 , n1390 , n1391 , n30482 , 
 n1393 , n30484 , n30485 , n1396 , n30487 , n1398 , n1399 , n1400 , n1401 , n1402 , 
 n1403 , n30494 , n1405 , n30496 , n30497 , n1411 , n1412 , n30500 , n30501 , n1415 , 
 n30503 , n30504 , n1418 , n30506 , n30507 , n30508 , n1422 , n30510 , n30511 , n1425 , 
 n30513 , n30514 , n30515 , n1429 , n30517 , n1431 , n30519 , n30520 , n30521 , n1435 , 
 n30523 , n1437 , n30525 , n1439 , n30527 , n30528 , n1442 , n30530 , n30531 , n1445 , 
 n30533 , n30534 , n1448 , n30536 , n30537 , n1451 , n1452 , n1453 , n30541 , n30542 , 
 n30543 , n1460 , n30545 , n1462 , n30547 , n1464 , n1465 , n30550 , n1467 , n30552 , 
 n1469 , n1470 , n30555 , n30556 , n1473 , n30558 , n30559 , n1476 , n30561 , n30562 , 
 n30563 , n1480 , n30565 , n30566 , n1483 , n30568 , n30569 , n30570 , n30571 , n1488 , 
 n30573 , n30574 , n1491 , n1492 , n1493 , n1494 , n1495 , n30580 , n1497 , n30582 , 
 n30583 , n1500 , n30585 , n30586 , n1503 , n30588 , n1505 , n30590 , n1507 , n30592 , 
 n30593 , n1510 , n1511 , n30596 , n30597 , n1514 , n30599 , n30600 , n1517 , n30602 , 
 n30603 , n1520 , n30605 , n30606 , n1523 , n1524 , n30609 , n1526 , n30611 , n1528 , 
 n1529 , n30614 , n30615 , n1532 , n30617 , n30618 , n1535 , n30620 , n30621 , n30622 , 
 n1539 , n30624 , n30625 , n1542 , n30627 , n30628 , n1545 , n30630 , n1547 , n30632 , 
 n1549 , n1550 , n30635 , n30636 , n1553 , n30638 , n1555 , n1556 , n30641 , n30642 , 
 n1559 , n30644 , n30645 , n1562 , n30647 , n30648 , n1565 , n30650 , n30651 , n1568 , 
 n30653 , n30654 , n30655 , n30656 , n30657 , n1577 , n30659 , n1579 , n1580 , n1581 , 
 n1582 , n1583 , n30665 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , 
 n1592 , n1593 , n1594 , n30676 , n1596 , n30678 , n1598 , n30680 , n30681 , n30682 , 
 n1605 , n30684 , n30685 , n30686 , n1609 , n30688 , n30689 , n1612 , n30691 , n30692 , 
 n30693 , n30694 , n1617 , n30696 , n1619 , n30698 , n30699 , n30700 , n30701 , n1624 , 
 n30703 , n30704 , n30705 , n1628 , n30707 , n30708 , n1631 , n30710 , n30711 , n1634 , 
 n1635 , n1636 , n1637 , n30716 , n30717 , n1640 , n30719 , n1642 , n30721 , n1644 , 
 n1645 , n30724 , n30725 , n1648 , n30727 , n30728 , n30729 , n1652 , n30731 , n30732 , 
 n1655 , n30734 , n30735 , n30736 , n1659 , n1660 , n30739 , n1662 , n30741 , n30742 , 
 n1665 , n30744 , n30745 , n30746 , n1669 , n30748 , n30749 , n1675 , n30751 , n1677 , 
 n30753 , n30754 , n1680 , n30756 , n30757 , n1683 , n30759 , n30760 , n1686 , n30762 , 
 n30763 , n1689 , n1690 , n1691 , n30767 , n1693 , n30769 , n30770 , n1696 , n1697 , 
 n1698 , n30774 , n1700 , n30776 , n1702 , n30778 , n30779 , n1705 , n30781 , n30782 , 
 n1708 , n30784 , n30785 , n1711 , n30787 , n1713 , n30789 , n1715 , n1716 , n30792 , 
 n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , 
 n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n30811 , n1740 , 
 n30813 , n30814 , n1743 , n30816 , n1745 , n30818 , n1747 , n1748 , n1749 , n1750 , 
 n1751 , n30824 , n1753 , n30826 , n1755 , n30828 , n1757 , n1758 , n30831 , n30832 , 
 n1761 , n30834 , n30835 , n30836 , n1765 , n30838 , n30839 , n1768 , n30841 , n30842 , 
 n30843 , n30844 , n1773 , n30846 , n30847 , n30848 , n1777 , n30850 , n30851 , n1780 , 
 n30853 , n1782 , n30855 , n1784 , n1785 , n1786 , n30859 , n1788 , n30861 , n1790 , 
 n30863 , n30864 , n1793 , n30866 , n30867 , n1796 , n30869 , n30870 , n1799 , n1800 , 
 n1801 , n1802 , n30875 , n30876 , n1805 , n30878 , n1807 , n30880 , n1809 , n1810 , 
 n30883 , n30884 , n30885 , n1814 , n30887 , n30888 , n30889 , n30890 , n30891 , n1820 , 
 n30893 , n30894 , n30895 , n30896 , n1825 , n30898 , n30899 , n1828 , n30901 , n30902 , 
 n1831 , n30904 , n30905 , n1834 , n30907 , n1836 , n1837 , n30910 , n1839 , n30912 , 
 n30913 , n30914 , n1843 , n1844 , n30917 , n30918 , n1847 , n30920 , n30921 , n1850 , 
 n30923 , n1852 , n1853 , n1854 , n1855 , n30928 , n1857 , n1858 , n1859 , n1860 , 
 n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1870 , n30940 , n1872 , n1873 , 
 n1874 , n1875 , n1876 , n30946 , n1878 , n30948 , n1880 , n1881 , n1882 , n1883 , 
 n30953 , n1885 , n1886 , n30956 , n30957 , n1889 , n30959 , n30960 , n1892 , n30962 , 
 n30963 , n1895 , n1896 , n30966 , n30967 , n1899 , n30969 , n30970 , n1905 , n30972 , 
 n30973 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n30981 , n1916 , 
 n30983 , n1918 , n1919 , n30986 , n1921 , n30988 , n1923 , n1924 , n30991 , n1926 , 
 n30993 , n1928 , n30995 , n30996 , n1931 , n30998 , n30999 , n1934 , n31001 , n31002 , 
 n1937 , n31004 , n31005 , n1940 , n1941 , n31008 , n31009 , n1944 , n31011 , n31012 , 
 n1947 , n31014 , n1949 , n1950 , n1951 , n31018 , n1953 , n31020 , n1955 , n1956 , 
 n31023 , n1958 , n1959 , n1960 , n1961 , n31028 , n31029 , n1964 , n31031 , n1966 , 
 n31033 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n31040 , n31041 , n1976 , 
 n31043 , n31044 , n1979 , n31046 , n31047 , n31048 , n1983 , n31050 , n1985 , n31052 , 
 n1987 , n1991 , n31055 , n31056 , n1994 , n31058 , n31059 , n1997 , n31061 , n31062 , 
 n2000 , n2001 , n31065 , n31066 , n2004 , n31068 , n31069 , n2007 , n31071 , n31072 , 
 n2010 , n31074 , n31075 , n2013 , n31077 , n31078 , n2016 , n31080 , n31081 , n2019 , 
 n31083 , n2021 , n2022 , n2023 , n2024 , n31088 , n2026 , n2027 , n2028 , n2029 , 
 n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n31101 , n2039 , 
 n31103 , n2041 , n2042 , n31106 , n31107 , n2045 , n31109 , n2047 , n2048 , n2049 , 
 n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n31122 , 
 n2063 , n2064 , n2065 , n2066 , n31127 , n2068 , n31129 , n31130 , n2071 , n31132 , 
 n31133 , n2074 , n31135 , n31136 , n31137 , n31138 , n2079 , n31140 , n31141 , n31142 , 
 n31143 , n2084 , n31145 , n31146 , n2087 , n31148 , n31149 , n2090 , n31151 , n31152 , 
 n2093 , n31154 , n31155 , n31156 , n31157 , n31158 , n2099 , n31160 , n31161 , n31162 , 
 n31163 , n31164 , n2105 , n31166 , n31167 , n2108 , n31169 , n31170 , n2111 , n31172 , 
 n31173 , n2114 , n31175 , n31176 , n31177 , n31178 , n2119 , n31180 , n31181 , n2122 , 
 n31183 , n31184 , n2125 , n31186 , n31187 , n2128 , n2129 , n2130 , n31191 , n31192 , 
 n2133 , n31194 , n31195 , n2136 , n31197 , n31198 , n31199 , n31200 , n31201 , n2142 , 
 n31203 , n31204 , n2145 , n31206 , n31207 , n31208 , n2149 , n31210 , n2151 , n31212 , 
 n31213 , n2154 , n2155 , n31216 , n2157 , n31218 , n31219 , n2160 , n2161 , n2162 , 
 n31223 , n31224 , n2165 , n2166 , n2167 , n31228 , n31229 , n2170 , n31231 , n31232 , 
 n2173 , n2174 , n31235 , n31236 , n31237 , n31238 , n2179 , n31240 , n31241 , n31242 , 
 n31243 , n2184 , n31245 , n31246 , n2187 , n2188 , n31249 , n31250 , n2191 , n2192 , 
 n2193 , n31254 , n31255 , n2196 , n31257 , n31258 , n31259 , n31260 , n31261 , n2202 , 
 n31263 , n31264 , n2208 , n31266 , n31267 , n31268 , n31269 , n2213 , n31271 , n31272 , 
 n31273 , n2217 , n31275 , n31276 , n2220 , n31278 , n31279 , n2223 , n31281 , n31282 , 
 n2226 , n2227 , n31285 , n31286 , n2230 , n2231 , n2232 , n31290 , n31291 , n2235 , 
 n2236 , n2237 , n31295 , n31296 , n2240 , n2241 , n2242 , n31300 , n31301 , n2248 , 
 n31303 , n31304 , n2251 , n31306 , n31307 , n2254 , n31309 , n31310 , n2257 , n31312 , 
 n31313 , n2260 , n31315 , n31316 , n2263 , n31318 , n31319 , n2266 , n31321 , n31322 , 
 n2269 , n31324 , n31325 , n31326 , n31327 , n2274 , n31329 , n31330 , n2277 , n2278 , 
 n31333 , n31334 , n2281 , n31336 , n31337 , n2284 , n2285 , n2286 , n2287 , n31342 , 
 n31343 , n2290 , n31345 , n31346 , n31347 , n2294 , n31349 , n31350 , n2297 , n31352 , 
 n31353 , n2300 , n2301 , n2302 , n2303 , n31358 , n31359 , n2306 , n31361 , n31362 , 
 n2309 , n31364 , n31365 , n31366 , n31367 , n2314 , n31369 , n31370 , n2317 , n31372 , 
 n31373 , n2320 , n31375 , n31376 , n2323 , n31378 , n31379 , n2326 , n31381 , n31382 , 
 n2329 , n31384 , n31385 , n2332 , n2333 , n2334 , n2335 , n31390 , n31391 , n2338 , 
 n31393 , n31394 , n31395 , n31396 , n2343 , n31398 , n31399 , n2346 , n31401 , n31402 , 
 n2349 , n2350 , n31405 , n31406 , n2353 , n2354 , n31409 , n2356 , n2357 , n2358 , 
 n2359 , n31414 , n31415 , n31416 , n31417 , n31418 , n2365 , n31420 , n31421 , n2368 , 
 n31423 , n31424 , n2371 , n2372 , n2373 , n2374 , n2375 , n31430 , n31431 , n2378 , 
 n31433 , n31434 , n2381 , n2382 , n2383 , n2384 , n31439 , n31440 , n2387 , n31442 , 
 n31443 , n2390 , n31445 , n31446 , n31447 , n31448 , n2395 , n31450 , n31451 , n2398 , 
 n31453 , n31454 , n2401 , n31456 , n31457 , n2404 , n31459 , n31460 , n31461 , n31462 , 
 n2412 , n31464 , n31465 , n31466 , n31467 , n2417 , n31469 , n31470 , n2420 , n31472 , 
 n31473 , n2423 , n31475 , n31476 , n2426 , n31478 , n31479 , n2429 , n2430 , n2431 , 
 n2432 , n2433 , n31485 , n31486 , n2436 , n31488 , n31489 , n2439 , n31491 , n31492 , 
 n2442 , n2443 , n2444 , n2445 , n31497 , n31498 , n2448 , n31500 , n31501 , n31502 , 
 n31503 , n2453 , n31505 , n31506 , n2456 , n31508 , n31509 , n2459 , n31511 , n2461 , 
 n31513 , n2463 , n2464 , n31516 , n2466 , n31518 , n31519 , n2469 , n2470 , n31522 , 
 n31523 , n2473 , n2474 , n31526 , n2476 , n2477 , n2478 , n2479 , n2480 , n31532 , 
 n31533 , n2483 , n2484 , n2485 , n2486 , n31538 , n31539 , n2489 , n31541 , n31542 , 
 n2492 , n31544 , n31545 , n31546 , n31547 , n2497 , n31549 , n31550 , n2500 , n31552 , 
 n31553 , n2503 , n31555 , n31556 , n2506 , n31558 , n31559 , n2509 , n31561 , n31562 , 
 n2512 , n2513 , n2514 , n2515 , n31567 , n31568 , n2518 , n31570 , n31571 , n2521 , 
 n31573 , n31574 , n31575 , n31576 , n2526 , n31578 , n31579 , n2529 , n31581 , n31582 , 
 n2532 , n31584 , n31585 , n2535 , n31587 , n31588 , n2538 , n2539 , n2540 , n2541 , 
 n31593 , n31594 , n2544 , n31596 , n31597 , n2547 , n31599 , n31600 , n31601 , n31602 , 
 n31603 , n2553 , n31605 , n31606 , n2556 , n31608 , n31609 , n2559 , n2560 , n31612 , 
 n31613 , n2563 , n31615 , n31616 , n2566 , n31618 , n31619 , n31620 , n31621 , n31622 , 
 n2575 , n2576 , n2577 , n2578 , n31627 , n31628 , n2581 , n31630 , n31631 , n31632 , 
 n31633 , n2586 , n31635 , n31636 , n2589 , n31638 , n31639 , n2592 , n31641 , n2594 , 
 n31643 , n2596 , n31645 , n2598 , n2599 , n31648 , n2601 , n31650 , n31651 , n2604 , 
 n2605 , n31654 , n2607 , n31656 , n31657 , n2610 , n2611 , n31660 , n31661 , n2614 , 
 n2615 , n31664 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , 
 n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n31679 , n2632 , n2633 , n2634 , 
 n2635 , n2636 , n2637 , n31686 , n2639 , n2640 , n31689 , n2642 , n31691 , n2644 , 
 n31693 , n31694 , n2647 , n2648 , n31697 , n31698 , n31699 , n31700 , n31701 , n2654 , 
 n31703 , n31704 , n31705 , n2658 , n31707 , n31708 , n2661 , n31710 , n31711 , n31712 , 
 n2665 , n31714 , n2667 , n2668 , n2669 , n2670 , n2671 , n31720 , n2673 , n2674 , 
 n2675 , n2676 , n2677 , n2678 , n2679 , n31728 , n31729 , n2682 , n31731 , n31732 , 
 n2685 , n31734 , n31735 , n2688 , n2689 , n2690 , n2691 , n2692 , n31741 , n31742 , 
 n2695 , n31744 , n31745 , n2698 , n31747 , n2700 , n31749 , n31750 , n2703 , n2704 , 
 n31753 , n2706 , n31755 , n2708 , n31757 , n2710 , n31759 , n2712 , n31761 , n31762 , 
 n2715 , n2716 , n31765 , n2718 , n31767 , n2720 , n2721 , n31770 , n2723 , n2724 , 
 n2725 , n31774 , n2727 , n31776 , n2729 , n31778 , n2731 , n2732 , n31781 , n31782 , 
 n2738 , n31784 , n31785 , n2741 , n31787 , n31788 , n2744 , n31790 , n31791 , n2747 , 
 n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n31800 , n2756 , n31802 , 
 n31803 , n31804 , n2760 , n31806 , n31807 , n2763 , n31809 , n31810 , n2766 , n31812 , 
 n31813 , n2769 , n31815 , n31816 , n2772 , n31818 , n31819 , n31820 , n2776 , n31822 , 
 n2778 , n31824 , n2780 , n31826 , n31827 , n2783 , n31829 , n31830 , n2786 , n2787 , 
 n31833 , n31834 , n2790 , n31836 , n31837 , n2793 , n31839 , n31840 , n2796 , n2797 , 
 n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , 
 n31853 , n2809 , n31855 , n2811 , n31857 , n31858 , n2814 , n31860 , n31861 , n2817 , 
 n31863 , n2819 , n31865 , n2821 , n31867 , n2823 , n2824 , n2825 , n2826 , n2827 , 
 n2828 , n2829 , n2830 , n2831 , n2832 , n31878 , n2834 , n31880 , n31881 , n2837 , 
 n2838 , n31884 , n31885 , n2841 , n2842 , n2843 , n2844 , n2845 , n31891 , n2847 , 
 n2848 , n31894 , n31895 , n2851 , n31897 , n31898 , n2854 , n31900 , n31901 , n2857 , 
 n31903 , n31904 , n2860 , n31906 , n31907 , n2863 , n2864 , n2865 , n31911 , n31912 , 
 n2868 , n31914 , n2870 , n31916 , n2872 , n31918 , n2874 , n2875 , n2876 , n2877 , 
 n2878 , n2879 , n31925 , n2881 , n31927 , n2883 , n2884 , n31930 , n31931 , n2887 , 
 n2888 , n31934 , n31935 , n31936 , n2895 , n31938 , n2897 , n2898 , n2899 , n31942 , 
 n2901 , n31944 , n2903 , n2904 , n31947 , n2906 , n31949 , n2908 , n31951 , n31952 , 
 n2911 , n2912 , n31955 , n31956 , n2915 , n31958 , n31959 , n2918 , n31961 , n31962 , 
 n31963 , n2922 , n31965 , n31966 , n2925 , n31968 , n2927 , n2928 , n31971 , n2930 , 
 n31973 , n2932 , n2933 , n2934 , n31977 , n2936 , n31979 , n2938 , n2939 , n2940 , 
 n2941 , n2942 , n2943 , n2944 , n31987 , n2946 , n2947 , n31990 , n31991 , n2950 , 
 n31993 , n31994 , n2953 , n31996 , n31997 , n2956 , n2957 , n2958 , n2959 , n2960 , 
 n2961 , n32004 , n32005 , n2964 , n32007 , n32008 , n2967 , n32010 , n2969 , n2970 , 
 n32013 , n32014 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n32021 , n2980 , 
 n32023 , n32024 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n32032 , 
 n2991 , n32034 , n2993 , n2994 , n2995 , n2996 , n32039 , n2998 , n32041 , n3000 , 
 n32043 , n3002 , n32045 , n3004 , n3005 , n32048 , n32049 , n3008 , n32051 , n32052 , 
 n3011 , n32054 , n32055 , n3014 , n3015 , n32058 , n32059 , n3018 , n32061 , n32062 , 
 n3021 , n32064 , n32065 , n3024 , n3025 , n3026 , n32069 , n32070 , n3029 , n3030 , 
 n3031 , n32074 , n32075 , n3034 , n3035 , n32078 , n32079 , n3041 , n32081 , n3043 , 
 n3044 , n3045 , n32085 , n3047 , n32087 , n32088 , n3050 , n32090 , n32091 , n32092 , 
 n3054 , n32094 , n3056 , n32096 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , 
 n3064 , n32104 , n3066 , n32106 , n32107 , n3069 , n3070 , n32110 , n3072 , n32112 , 
 n3074 , n32114 , n32115 , n3077 , n32117 , n32118 , n3080 , n32120 , n3082 , n32122 , 
 n3084 , n32124 , n3086 , n32126 , n32127 , n3089 , n3090 , n32130 , n32131 , n3093 , 
 n32133 , n32134 , n3096 , n32136 , n32137 , n3099 , n3100 , n32140 , n32141 , n3103 , 
 n32143 , n32144 , n3106 , n32146 , n32147 , n3109 , n32149 , n32150 , n3112 , n3113 , 
 n32153 , n3115 , n32155 , n3117 , n32157 , n3119 , n3120 , n32160 , n32161 , n3123 , 
 n32163 , n32164 , n3126 , n32166 , n32167 , n3129 , n3130 , n32170 , n3132 , n32172 , 
 n3134 , n3135 , n32175 , n32176 , n3138 , n32178 , n32179 , n3141 , n32181 , n32182 , 
 n3144 , n3145 , n3146 , n32186 , n3148 , n32188 , n32189 , n3151 , n32191 , n3153 , 
 n32193 , n3155 , n32195 , n3157 , n3158 , n32198 , n32199 , n3161 , n32201 , n32202 , 
 n3164 , n32204 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n32211 , n3176 , 
 n3177 , n3178 , n3179 , n32216 , n3181 , n32218 , n3183 , n32220 , n3185 , n3186 , 
 n32223 , n3188 , n32225 , n3190 , n3191 , n32228 , n32229 , n3194 , n32231 , n32232 , 
 n3197 , n32234 , n32235 , n32236 , n3201 , n32238 , n32239 , n3204 , n32241 , n32242 , 
 n3207 , n3208 , n3209 , n3210 , n3211 , n32248 , n3213 , n3214 , n3215 , n3216 , 
 n3217 , n3218 , n3219 , n3220 , n32257 , n32258 , n3223 , n32260 , n32261 , n3226 , 
 n32263 , n32264 , n3229 , n32266 , n32267 , n3232 , n32269 , n3234 , n3235 , n32272 , 
 n32273 , n3238 , n3239 , n32276 , n32277 , n32278 , n3243 , n32280 , n32281 , n3246 , 
 n32283 , n3248 , n32285 , n32286 , n3251 , n3252 , n32289 , n32290 , n3255 , n32292 , 
 n32293 , n3258 , n3259 , n32296 , n3261 , n32298 , n32299 , n3264 , n3265 , n32302 , 
 n32303 , n3268 , n32305 , n32306 , n3271 , n32308 , n3273 , n3274 , n32311 , n32312 , 
 n3277 , n3278 , n3279 , n32316 , n3281 , n3282 , n32319 , n3284 , n32321 , n3286 , 
 n32323 , n3288 , n3289 , n3290 , n3291 , n32328 , n3293 , n32330 , n32331 , n32332 , 
 n3297 , n32334 , n3302 , n32336 , n32337 , n32338 , n3306 , n32340 , n3308 , n32342 , 
 n32343 , n3311 , n3312 , n32346 , n3314 , n32348 , n32349 , n3317 , n32351 , n32352 , 
 n32353 , n3321 , n32355 , n3323 , n3324 , n32358 , n3326 , n3327 , n3328 , n3329 , 
 n32363 , n3331 , n32365 , n32366 , n3334 , n32368 , n32369 , n3337 , n32371 , n32372 , 
 n3340 , n3341 , n32375 , n32376 , n3344 , n3345 , n3346 , n3347 , n32381 , n3349 , 
 n32383 , n3351 , n3352 , n3353 , n3354 , n32388 , n32389 , n32390 , n32391 , n3359 , 
 n32393 , n3361 , n32395 , n3363 , n3364 , n3365 , n3366 , n32400 , n3368 , n32402 , 
 n3370 , n32404 , n3372 , n32406 , n3374 , n3375 , n32409 , n32410 , n3378 , n32412 , 
 n32413 , n3381 , n32415 , n3383 , n3384 , n3385 , n32419 , n3387 , n3388 , n3389 , 
 n32423 , n3391 , n3392 , n3393 , n32427 , n3395 , n3396 , n3397 , n3398 , n3399 , 
 n32433 , n3401 , n32435 , n3403 , n32437 , n32438 , n32439 , n3407 , n32441 , n3409 , 
 n32443 , n3411 , n32445 , n32446 , n3417 , n32448 , n32449 , n3420 , n32451 , n32452 , 
 n32453 , n3424 , n32455 , n3426 , n3427 , n32458 , n3429 , n3430 , n3431 , n3432 , 
 n3433 , n3434 , n32465 , n3436 , n32467 , n32468 , n3439 , n3440 , n32471 , n32472 , 
 n3443 , n32474 , n32475 , n3446 , n32477 , n32478 , n32479 , n3450 , n32481 , n32482 , 
 n3453 , n32484 , n32485 , n3456 , n32487 , n32488 , n3459 , n3460 , n3461 , n3462 , 
 n32493 , n32494 , n3465 , n32496 , n32497 , n32498 , n3469 , n32500 , n32501 , n3472 , 
 n3473 , n32504 , n3475 , n32506 , n3477 , n3478 , n32509 , n3480 , n32511 , n32512 , 
 n3483 , n32514 , n32515 , n3486 , n32517 , n3488 , n3489 , n3490 , n3491 , n32522 , 
 n3493 , n32524 , n3495 , n32526 , n3497 , n32528 , n3499 , n3500 , n32531 , n32532 , 
 n3503 , n32534 , n32535 , n3506 , n32537 , n32538 , n3509 , n3510 , n3511 , n3512 , 
 n32543 , n3514 , n32545 , n3516 , n32547 , n32548 , n32549 , n3523 , n3524 , n32552 , 
 n3526 , n3527 , n32555 , n32556 , n3530 , n3531 , n32559 , n32560 , n3534 , n32562 , 
 n32563 , n32564 , n3538 , n32566 , n3540 , n3541 , n32569 , n32570 , n3544 , n3545 , 
 n32573 , n32574 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n32582 , 
 n3556 , n32584 , n32585 , n3559 , n32587 , n3561 , n3562 , n3563 , n32591 , n3565 , 
 n32593 , n32594 , n3568 , n32596 , n32597 , n3571 , n3572 , n32600 , n3574 , n3575 , 
 n32603 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , 
 n3586 , n3587 , n32615 , n3589 , n32617 , n3591 , n3592 , n3593 , n3594 , n3595 , 
 n3596 , n3597 , n3598 , n3599 , n32627 , n32628 , n3602 , n32630 , n3604 , n3605 , 
 n32633 , n3607 , n32635 , n32636 , n3610 , n32638 , n32639 , n3616 , n32641 , n3618 , 
 n32643 , n3620 , n3621 , n3622 , n32647 , n3624 , n32649 , n32650 , n32651 , n3628 , 
 n3629 , n32654 , n3631 , n32656 , n3633 , n32658 , n3635 , n32660 , n32661 , n3638 , 
 n3639 , n32664 , n32665 , n3642 , n32667 , n32668 , n3645 , n32670 , n32671 , n32672 , 
 n3649 , n32674 , n32675 , n3652 , n3653 , n32678 , n3655 , n3656 , n32681 , n3658 , 
 n3659 , n3660 , n32685 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , 
 n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n32702 , 
 n32703 , n3680 , n32705 , n3682 , n3683 , n32708 , n3685 , n32710 , n3687 , n32712 , 
 n32713 , n3690 , n32715 , n32716 , n3693 , n32718 , n32719 , n3696 , n32721 , n32722 , 
 n32723 , n3703 , n3704 , n32726 , n3706 , n32728 , n3708 , n3709 , n32731 , n3711 , 
 n32733 , n32734 , n32735 , n3715 , n32737 , n3717 , n32739 , n32740 , n3720 , n32742 , 
 n32743 , n3723 , n3724 , n3725 , n32747 , n32748 , n3728 , n3729 , n3730 , n32752 , 
 n32753 , n3733 , n3734 , n3735 , n32757 , n32758 , n3738 , n3739 , n3740 , n32762 , 
 n3742 , n3743 , n32765 , n3745 , n3746 , n3747 , n3748 , n32770 , n32771 , n3751 , 
 n3752 , n3753 , n32775 , n32776 , n3756 , n3757 , n3758 , n32780 , n3760 , n3761 , 
 n3762 , n3763 , n3764 , n3765 , n3766 , n32788 , n3768 , n3769 , n3770 , n32792 , 
 n32793 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , 
 n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , 
 n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , 
 n32823 , n3806 , n32825 , n32826 , n3809 , n32828 , n3811 , n3812 , n32831 , n3814 , 
 n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n32839 , n3822 , n3823 , n32842 , 
 n32843 , n3826 , n3827 , n32846 , n32847 , n3830 , n32849 , n3832 , n3833 , n3834 , 
 n32853 , n32854 , n3837 , n32856 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , 
 n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , 
 n32873 , n32874 , n3860 , n32876 , n32877 , n3863 , n32879 , n32880 , n3866 , n32882 , 
 n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n32889 , n3875 , n3876 , n32892 , 
 n32893 , n3879 , n32895 , n32896 , n3882 , n32898 , n32899 , n3885 , n32901 , n32902 , 
 n3888 , n32904 , n3890 , n3891 , n32907 , n3896 , n3897 , n3898 , n3899 , n3900 , 
 n3901 , n3902 , n32915 , n3904 , n32917 , n3906 , n3907 , n3908 , n3909 , n3910 , 
 n32923 , n32924 , n3913 , n32926 , n3915 , n32928 , n32929 , n3918 , n32931 , n32932 , 
 n3921 , n32934 , n32935 , n32936 , n3925 , n32938 , n3927 , n32940 , n3929 , n3930 , 
 n32943 , n32944 , n3933 , n32946 , n32947 , n3936 , n32949 , n32950 , n3942 , n3943 , 
 n32953 , n3945 , n3946 , n3947 , n3948 , n32958 , n3950 , n32960 , n32961 , n3953 , 
 n32963 , n32964 , n3956 , n32966 , n32967 , n32968 , n3960 , n32970 , n3962 , n3963 , 
 n32973 , n3965 , n32975 , n3967 , n3968 , n3969 , n3970 , n3971 , n32981 , n3976 , 
 n32983 , n3978 , n32985 , n3980 , n3981 , n3982 , n32989 , n32990 , n32991 , n32992 , 
 n3987 , n32994 , n3989 , n3990 , n3991 , n32998 , n32999 , n3994 , n33001 , n3996 , 
 n3997 , n3998 , n33005 , n4000 , n4001 , n33008 , n4003 , n4004 , n4005 , n33012 , 
 n33013 , n33014 , n4009 , n4010 , n4011 , n33018 , n4013 , n4014 , n4015 , n4016 , 
 n4017 , n33024 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n33031 , n4026 , 
 n4027 , n4028 , n33035 , n4030 , n33037 , n4032 , n4033 , n33040 , n4035 , n33042 , 
 n4037 , n4038 , n4039 , n4040 , n33047 , n33048 , n33049 , n4044 , n4045 , n4046 , 
 n4047 , n33054 , n4049 , n33056 , n4051 , n33058 , n4053 , n4054 , n4055 , n4056 , 
 n33063 , n33064 , n4059 , n33066 , n33067 , n4062 , n33069 , n33070 , n4065 , n33072 , 
 n33073 , n4068 , n33075 , n4070 , n33077 , n33078 , n33079 , n33080 , n4075 , n33082 , 
 n33083 , n33084 , n4079 , n33086 , n33087 , n4082 , n33089 , n33090 , n4085 , n4086 , 
 n33093 , n33094 , n4089 , n4090 , n33097 , n33098 , n33099 , n33100 , n4095 , n33102 , 
 n33103 , n33104 , n4099 , n33106 , n33107 , n4102 , n33109 , n4104 , n33111 , n4106 , 
 n4107 , n33114 , n4109 , n33116 , n4111 , n33118 , n33119 , n4114 , n33121 , n33122 , 
 n4117 , n4118 , n33125 , n4120 , n33127 , n33128 , n4123 , n33130 , n33131 , n33132 , 
 n4127 , n33134 , n33135 , n4130 , n33137 , n33138 , n4133 , n33140 , n33141 , n33142 , 
 n4137 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , 
 n33153 , n33154 , n4149 , n33156 , n33157 , n33158 , n4153 , n33160 , n33161 , n4156 , 
 n33163 , n33164 , n33165 , n4160 , n33167 , n4162 , n33169 , n33170 , n4165 , n33172 , 
 n4170 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , 
 n4183 , n33184 , n33185 , n33186 , n33187 , n33188 , n4189 , n33190 , n33191 , n4192 , 
 n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n4199 , n33200 , n33201 , n4202 , 
 n33203 , n33204 , n4205 , n33206 , n4207 , n33208 , n33209 , n4210 , n33211 , n33212 , 
 n4213 , n4214 , n33215 , n4216 , n4217 , n4218 , n33219 , n4220 , n4221 , n33222 , 
 n33223 , n4224 , n33225 , n33226 , n33227 , n4228 , n33229 , n4230 , n33231 , n33232 , 
 n33233 , n4234 , n33235 , n33236 , n33237 , n33238 , n4239 , n33240 , n4241 , n4242 , 
 n33243 , n4244 , n33245 , n4249 , n33247 , n33248 , n4252 , n4253 , n33251 , n33252 , 
 n4259 , n4260 , n33255 , n33256 , n33257 , n4264 , n33259 , n33260 , n4267 , n4268 , 
 n33263 , n33264 , n4271 , n4272 , n33267 , n4274 , n4275 , n4276 , n33271 , n33272 , 
 n33273 , n33274 , n4281 , n33276 , n33277 , n4284 , n33279 , n33280 , n33281 , n33282 , 
 n33283 , n33284 , n4291 , n33286 , n33287 , n4294 , n33289 , n33290 , n4297 , n33292 , 
 n33293 , n4300 , n33295 , n33296 , n33297 , n33298 , n4305 , n33300 , n33301 , n33302 , 
 n33303 , n4310 , n33305 , n33306 , n33307 , n4314 , n33309 , n4316 , n33311 , n33312 , 
 n4319 , n33314 , n4321 , n4322 , n4323 , n33318 , n33319 , n4326 , n33321 , n33322 , 
 n33323 , n33324 , n4331 , n4332 , n33327 , n4334 , n4335 , n4336 , n33331 , n33332 , 
 n33333 , n33334 , n4344 , n33336 , n33337 , n4347 , n4348 , n4349 , n33341 , n33342 , 
 n33343 , n33344 , n33345 , n4358 , n33347 , n33348 , n4361 , n33350 , n33351 , n4364 , 
 n33353 , n33354 , n33355 , n33356 , n33357 , n4370 , n33359 , n4372 , n4373 , n33362 , 
 n33363 , n33364 , n4377 , n33366 , n33367 , n4380 , n33369 , n33370 , n4383 , n33372 , 
 n33373 , n4386 , n4387 , n4388 , n4389 , n33378 , n33379 , n4392 , n33381 , n33382 , 
 n33383 , n33384 , n4397 , n33386 , n33387 , n4400 , n33389 , n4402 , n33391 , n4404 , 
 n33393 , n33394 , n4407 , n33396 , n33397 , n4410 , n33399 , n33400 , n4413 , n33402 , 
 n33403 , n4416 , n33405 , n33406 , n33407 , n4420 , n33409 , n33410 , n4423 , n33412 , 
 n33413 , n4426 , n33415 , n33416 , n33417 , n4430 , n33419 , n33420 , n33421 , n33422 , 
 n4435 , n33424 , n33425 , n33426 , n33427 , n4440 , n33429 , n33430 , n33431 , n33432 , 
 n33433 , n4449 , n33435 , n33436 , n33437 , n4453 , n33439 , n4458 , n4459 , n33442 , 
 n4461 , n33444 , n4463 , n33446 , n33447 , n4466 , n33449 , n4468 , n33451 , n33452 , 
 n4471 , n33454 , n4473 , n33456 , n4475 , n33458 , n33459 , n4478 , n33461 , n33462 , 
 n33463 , n33464 , n33465 , n4484 , n33467 , n4486 , n33469 , n4488 , n4489 , n33472 , 
 n33473 , n4492 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n4500 , 
 n33483 , n33484 , n4503 , n33486 , n33487 , n4506 , n33489 , n33490 , n4509 , n33492 , 
 n33493 , n4512 , n33495 , n4514 , n4515 , n33498 , n33499 , n4518 , n33501 , n33502 , 
 n4521 , n33504 , n33505 , n33506 , n33507 , n4526 , n33509 , n33510 , n4529 , n33512 , 
 n4531 , n4532 , n33515 , n33516 , n4535 , n33518 , n33519 , n4538 , n33521 , n33522 , 
 n4541 , n4542 , n33525 , n4544 , n33527 , n33528 , n33529 , n33530 , n33531 , n4550 , 
 n33533 , n33534 , n4553 , n33536 , n33537 , n4559 , n33539 , n4561 , n33541 , n33542 , 
 n4564 , n4565 , n33545 , n33546 , n33547 , n4572 , n33549 , n33550 , n4575 , n33552 , 
 n4577 , n4578 , n33555 , n33556 , n4581 , n33558 , n4583 , n4584 , n33561 , n33562 , 
 n4587 , n33564 , n4589 , n4590 , n33567 , n33568 , n4593 , n33570 , n4595 , n4596 , 
 n4597 , n33574 , n33575 , n4600 , n33577 , n4602 , n4603 , n33580 , n33581 , n4606 , 
 n33583 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , 
 n4617 , n4618 , n4619 , n4620 , n33597 , n33598 , n4623 , n33600 , n4625 , n33602 , 
 n33603 , n33604 , n4629 , n33606 , n33607 , n4632 , n33609 , n4634 , n4635 , n33612 , 
 n33613 , n4638 , n33615 , n33616 , n4641 , n33618 , n33619 , n33620 , n33621 , n33622 , 
 n33623 , n4648 , n33625 , n33626 , n4651 , n33628 , n33629 , n33630 , n33631 , n33632 , 
 n4657 , n33634 , n33635 , n4660 , n33637 , n33638 , n4663 , n4664 , n4665 , n33642 , 
 n4667 , n33644 , n33645 , n33646 , n4671 , n4672 , n4673 , n33650 , n4675 , n4676 , 
 n33653 , n33654 , n33655 , n4683 , n4684 , n33658 , n33659 , n4690 , n4691 , n4692 , 
 n33663 , n4694 , n4695 , n33666 , n33667 , n4698 , n4699 , n33670 , n4701 , n33672 , 
 n33673 , n4704 , n33675 , n4706 , n33677 , n33678 , n33679 , n33680 , n4711 , n33682 , 
 n33683 , n33684 , n4715 , n33686 , n33687 , n33688 , n4719 , n33690 , n4721 , n33692 , 
 n33693 , n33694 , n4725 , n33696 , n33697 , n4728 , n33699 , n33700 , n4731 , n33702 , 
 n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n33710 , n4741 , n4742 , 
 n33713 , n4744 , n33715 , n4746 , n4747 , n33718 , n33719 , n4750 , n33721 , n33722 , 
 n4753 , n33724 , n33725 , n33726 , n4757 , n33728 , n4759 , n4760 , n33731 , n33732 , 
 n4763 , n33734 , n33735 , n4766 , n33737 , n33738 , n4769 , n33740 , n33741 , n4772 , 
 n4773 , n33744 , n33745 , n4776 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , 
 n4783 , n33754 , n33755 , n4786 , n33757 , n33758 , n4789 , n4790 , n33761 , n33762 , 
 n4793 , n33764 , n33765 , n4796 , n33767 , n33768 , n33769 , n4800 , n4801 , n33772 , 
 n4803 , n4804 , n4805 , n33776 , n4810 , n33778 , n4812 , n33780 , n33781 , n4818 , 
 n4819 , n33784 , n4821 , n33786 , n33787 , n33788 , n4825 , n33790 , n4827 , n4828 , 
 n33793 , n33794 , n4831 , n33796 , n33797 , n4834 , n33799 , n33800 , n4837 , n33802 , 
 n33803 , n4840 , n4841 , n4842 , n4843 , n4844 , n33809 , n33810 , n4847 , n4848 , 
 n4849 , n33814 , n33815 , n4852 , n4853 , n4854 , n33819 , n4856 , n33821 , n4858 , 
 n4859 , n4860 , n4861 , n33826 , n33827 , n4864 , n33829 , n33830 , n33831 , n4868 , 
 n4869 , n4870 , n33835 , n33836 , n4873 , n4874 , n4875 , n33840 , n4877 , n4878 , 
 n4879 , n33844 , n33845 , n4882 , n4883 , n4884 , n33849 , n4886 , n33851 , n4888 , 
 n4889 , n33854 , n4891 , n33856 , n4893 , n4894 , n4895 , n4896 , n4897 , n33862 , 
 n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , 
 n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , 
 n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n33890 , n33891 , n4928 , 
 n4929 , n4930 , n33895 , n33896 , n4933 , n33898 , n4935 , n33900 , n33901 , n33902 , 
 n4939 , n33904 , n33905 , n4942 , n33907 , n4944 , n33909 , n4949 , n33911 , n33912 , 
 n4952 , n33914 , n4957 , n4958 , n4959 , n4960 , n33919 , n4962 , n4963 , n4964 , 
 n4965 , n33924 , n33925 , n4968 , n4969 , n4970 , n4971 , n4972 , n33931 , n33932 , 
 n4975 , n33934 , n33935 , n4978 , n33937 , n33938 , n4981 , n33940 , n33941 , n33942 , 
 n4985 , n33944 , n4987 , n4988 , n33947 , n33948 , n4991 , n33950 , n33951 , n33952 , 
 n4995 , n33954 , n33955 , n4998 , n33957 , n33958 , n5001 , n33960 , n5003 , n33962 , 
 n5005 , n33964 , n33965 , n5008 , n33967 , n33968 , n5011 , n5012 , n33971 , n5014 , 
 n33973 , n33974 , n33975 , n33976 , n5019 , n33978 , n33979 , n5022 , n33981 , n33982 , 
 n33983 , n33984 , n33985 , n5028 , n33987 , n33988 , n5031 , n5032 , n5033 , n33992 , 
 n5035 , n33994 , n5037 , n33996 , n5039 , n5040 , n5041 , n5042 , n5043 , n34002 , 
 n34003 , n34004 , n5047 , n34006 , n34007 , n5050 , n34009 , n5052 , n5053 , n5054 , 
 n5055 , n5056 , n5057 , n5058 , n5059 , n34018 , n34019 , n5062 , n34021 , n5064 , 
 n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n34030 , n5073 , n5074 , 
 n5075 , n5076 , n5077 , n34036 , n34037 , n5080 , n34039 , n34040 , n5083 , n34042 , 
 n34043 , n34044 , n34045 , n5088 , n34047 , n5090 , n5091 , n5092 , n5093 , n34052 , 
 n5098 , n34054 , n5100 , n5101 , n34057 , n5106 , n5107 , n5108 , n5109 , n5110 , 
 n5111 , n34064 , n5113 , n34066 , n5115 , n34068 , n5117 , n34070 , n5119 , n5120 , 
 n5121 , n34074 , n5123 , n34076 , n5125 , n5126 , n34079 , n5128 , n5129 , n34082 , 
 n5131 , n34084 , n34085 , n34086 , n34087 , n5136 , n34089 , n5138 , n34091 , n5140 , 
 n34093 , n5142 , n34095 , n34096 , n5145 , n34098 , n34099 , n34100 , n5149 , n34102 , 
 n5151 , n34104 , n34105 , n5154 , n5155 , n34108 , n5157 , n34110 , n5159 , n34112 , 
 n34113 , n5162 , n34115 , n5164 , n34117 , n5166 , n5167 , n5168 , n5169 , n5170 , 
 n5171 , n5172 , n34125 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , 
 n5181 , n34134 , n5183 , n34136 , n5185 , n34138 , n34139 , n5188 , n34141 , n5190 , 
 n5191 , n34144 , n5193 , n34146 , n5195 , n34148 , n34149 , n5198 , n34151 , n34152 , 
 n5201 , n5202 , n34155 , n5204 , n34157 , n34158 , n5207 , n5208 , n34161 , n34162 , 
 n5211 , n5212 , n5213 , n5214 , n34167 , n34168 , n5217 , n34170 , n34171 , n34172 , 
 n5221 , n34174 , n5223 , n34176 , n34177 , n5226 , n34179 , n5228 , n34181 , n5230 , 
 n34183 , n5232 , n34185 , n5234 , n34187 , n34188 , n5237 , n34190 , n34191 , n5240 , 
 n5241 , n34194 , n5243 , n34196 , n34197 , n34198 , n34199 , n34200 , n5249 , n5250 , 
 n34203 , n34204 , n34205 , n34206 , n34207 , n5259 , n34209 , n34210 , n5265 , n5266 , 
 n5267 , n5268 , n34215 , n34216 , n34217 , n5272 , n5273 , n5274 , n5275 , n34222 , 
 n34223 , n34224 , n5279 , n34226 , n5281 , n5282 , n34229 , n5284 , n34231 , n5286 , 
 n34233 , n34234 , n5289 , n34236 , n34237 , n34238 , n34239 , n5294 , n34241 , n5296 , 
 n34243 , n34244 , n34245 , n34246 , n5301 , n34248 , n34249 , n34250 , n5305 , n34252 , 
 n34253 , n34254 , n5309 , n34256 , n5311 , n5312 , n5313 , n34260 , n34261 , n5316 , 
 n34263 , n34264 , n5319 , n34266 , n34267 , n5322 , n34269 , n34270 , n5325 , n5326 , 
 n5327 , n5328 , n5329 , n34276 , n5331 , n34278 , n34279 , n5334 , n5335 , n5336 , 
 n5337 , n5338 , n34285 , n34286 , n5341 , n34288 , n34289 , n5344 , n34291 , n34292 , 
 n5347 , n5348 , n5349 , n34296 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , 
 n5357 , n5358 , n5359 , n5360 , n5361 , n34308 , n5363 , n5364 , n5365 , n34312 , 
 n34313 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , 
 n5377 , n34324 , n5379 , n5380 , n5381 , n34328 , n34329 , n5384 , n34331 , n5386 , 
 n5387 , n5388 , n5389 , n5390 , n5391 , n34338 , n5393 , n5394 , n5395 , n5396 , 
 n5397 , n5398 , n5399 , n34346 , n34347 , n5402 , n34349 , n5404 , n5405 , n5406 , 
 n34353 , n5408 , n34355 , n34356 , n5411 , n34358 , n34359 , n34360 , n34361 , n5416 , 
 n5417 , n5418 , n5419 , n5420 , n5421 , n34368 , n34369 , n34370 , n34371 , n5429 , 
 n34373 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , 
 n5443 , n34384 , n34385 , n5446 , n5447 , n5448 , n5449 , n5450 , n34391 , n5452 , 
 n5453 , n34394 , n5455 , n34396 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , 
 n34403 , n34404 , n5465 , n34406 , n34407 , n5468 , n34409 , n34410 , n34411 , n5472 , 
 n34413 , n34414 , n34415 , n34416 , n34417 , n5478 , n34419 , n5480 , n34421 , n5482 , 
 n5483 , n34424 , n5485 , n34426 , n5487 , n5488 , n34429 , n34430 , n5491 , n34432 , 
 n34433 , n5494 , n34435 , n34436 , n34437 , n5498 , n34439 , n34440 , n34441 , n34442 , 
 n34443 , n5504 , n34445 , n34446 , n5507 , n34448 , n34449 , n5510 , n5511 , n5512 , 
 n5513 , n34454 , n5515 , n5516 , n5517 , n5518 , n5519 , n34460 , n34461 , n5522 , 
 n34463 , n5524 , n34465 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , 
 n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , 
 n5543 , n5544 , n5545 , n5546 , n34487 , n5548 , n34489 , n5550 , n5551 , n5552 , 
 n5553 , n5554 , n34495 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , 
 n34503 , n34504 , n5565 , n34506 , n34507 , n5568 , n34509 , n34510 , n5571 , n5572 , 
 n5573 , n34514 , n5575 , n34516 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , 
 n34523 , n34524 , n34525 , n5586 , n34527 , n5588 , n34529 , n34530 , n34531 , n34532 , 
 n5596 , n5597 , n34535 , n5602 , n34537 , n34538 , n5605 , n34540 , n5607 , n5608 , 
 n34543 , n5610 , n34545 , n34546 , n5613 , n34548 , n34549 , n5616 , n34551 , n34552 , 
 n5619 , n34554 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n34562 , 
 n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , 
 n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , 
 n5649 , n5650 , n5651 , n5652 , n34587 , n5654 , n5655 , n5656 , n5657 , n5658 , 
 n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n34599 , n34600 , n5667 , n5668 , 
 n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , 
 n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , 
 n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n34630 , n5697 , n5698 , 
 n34633 , n5700 , n34635 , n34636 , n34637 , n5704 , n34639 , n34640 , n5707 , n34642 , 
 n34643 , n5710 , n34645 , n34646 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , 
 n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , 
 n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n34672 , 
 n5739 , n34674 , n5741 , n34676 , n34677 , n5744 , n34679 , n34680 , n5747 , n34682 , 
 n34683 , n5753 , n34685 , n5755 , n5756 , n34688 , n34689 , n5762 , n5763 , n34692 , 
 n5765 , n34694 , n34695 , n5768 , n34697 , n34698 , n5771 , n34700 , n34701 , n5774 , 
 n34703 , n34704 , n34705 , n5778 , n34707 , n34708 , n5781 , n5782 , n5783 , n5784 , 
 n5785 , n5786 , n5787 , n5788 , n5789 , n34718 , n5791 , n5792 , n5793 , n34722 , 
 n5795 , n34724 , n34725 , n34726 , n5799 , n34728 , n5801 , n5802 , n5803 , n5804 , 
 n5805 , n5806 , n5807 , n5808 , n34737 , n5810 , n5811 , n5812 , n5813 , n5814 , 
 n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , 
 n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , 
 n5835 , n5836 , n5837 , n34766 , n5839 , n34768 , n34769 , n34770 , n5843 , n34772 , 
 n34773 , n5846 , n34775 , n34776 , n5849 , n34778 , n34779 , n5852 , n34781 , n34782 , 
 n34783 , n5856 , n34785 , n5858 , n5859 , n34788 , n34789 , n5862 , n34791 , n34792 , 
 n5865 , n34794 , n34795 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , 
 n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , 
 n5885 , n5886 , n34815 , n34816 , n5889 , n34818 , n34819 , n5892 , n34821 , n34822 , 
 n5895 , n34824 , n34825 , n5898 , n5899 , n5900 , n34829 , n5902 , n34831 , n5904 , 
 n34833 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , 
 n5915 , n5916 , n34845 , n34846 , n5919 , n5920 , n34849 , n5925 , n34851 , n5927 , 
 n5928 , n34854 , n5933 , n5934 , n5935 , n34858 , n5937 , n34860 , n34861 , n5940 , 
 n34863 , n5942 , n5943 , n34866 , n5945 , n34868 , n5947 , n34870 , n34871 , n34872 , 
 n5951 , n34874 , n34875 , n5954 , n34877 , n34878 , n34879 , n5958 , n34881 , n34882 , 
 n5961 , n34884 , n5963 , n34886 , n5965 , n34888 , n5967 , n5968 , n5969 , n5970 , 
 n5971 , n5972 , n5973 , n5974 , n34897 , n34898 , n5977 , n34900 , n5979 , n5980 , 
 n5981 , n5982 , n5983 , n34906 , n34907 , n5986 , n34909 , n34910 , n5989 , n34912 , 
 n5991 , n5992 , n5993 , n34916 , n5995 , n34918 , n34919 , n34920 , n5999 , n34922 , 
 n6001 , n6002 , n34925 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , 
 n34933 , n34934 , n34935 , n6014 , n34937 , n34938 , n6017 , n34940 , n34941 , n34942 , 
 n34943 , n34944 , n6023 , n34946 , n34947 , n6026 , n34949 , n34950 , n6029 , n34952 , 
 n34953 , n6032 , n34955 , n34956 , n34957 , n34958 , n6037 , n34960 , n34961 , n6040 , 
 n34963 , n34964 , n6043 , n34966 , n34967 , n6046 , n6047 , n6048 , n34971 , n34972 , 
 n6051 , n6052 , n6053 , n34976 , n34977 , n34978 , n34979 , n6058 , n34981 , n34982 , 
 n34983 , n34984 , n34985 , n6064 , n34987 , n34988 , n6067 , n34990 , n34991 , n6070 , 
 n6071 , n34994 , n34995 , n6074 , n34997 , n34998 , n34999 , n35000 , n35001 , n6080 , 
 n35003 , n35004 , n35005 , n35006 , n6088 , n35008 , n35009 , n6094 , n35011 , n35012 , 
 n6097 , n35014 , n35015 , n6100 , n6101 , n6102 , n35019 , n35020 , n35021 , n35022 , 
 n6107 , n35024 , n35025 , n35026 , n35027 , n6112 , n35029 , n35030 , n6115 , n35032 , 
 n35033 , n6118 , n35035 , n35036 , n6121 , n6122 , n6123 , n35040 , n35041 , n6126 , 
 n35043 , n35044 , n6129 , n35046 , n35047 , n35048 , n35049 , n6134 , n35051 , n35052 , 
 n6137 , n35054 , n35055 , n6140 , n35057 , n35058 , n6143 , n35060 , n6145 , n35062 , 
 n35063 , n6148 , n35065 , n35066 , n6151 , n35068 , n35069 , n6154 , n35071 , n35072 , 
 n6157 , n6158 , n6159 , n6160 , n35077 , n35078 , n6163 , n6164 , n6165 , n35082 , 
 n6167 , n35084 , n35085 , n6170 , n6171 , n6172 , n35089 , n35090 , n35091 , n35092 , 
 n6177 , n35094 , n35095 , n35096 , n35097 , n6182 , n35099 , n35100 , n6185 , n35102 , 
 n35103 , n6188 , n35105 , n35106 , n6191 , n6192 , n6193 , n35110 , n35111 , n6196 , 
 n6197 , n35114 , n35115 , n6200 , n6201 , n6202 , n35119 , n35120 , n6205 , n35122 , 
 n35123 , n6208 , n6209 , n6210 , n35127 , n35128 , n6213 , n6214 , n35131 , n35132 , 
 n6217 , n6218 , n6219 , n6220 , n6221 , n35138 , n35139 , n6224 , n6225 , n6226 , 
 n35143 , n35144 , n6229 , n6230 , n6231 , n35148 , n35149 , n6234 , n6235 , n6236 , 
 n6237 , n6238 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , 
 n35163 , n35164 , n35165 , n35166 , n6257 , n35168 , n35169 , n6260 , n35171 , n35172 , 
 n6263 , n35174 , n35175 , n35176 , n35177 , n6268 , n35179 , n35180 , n35181 , n35182 , 
 n6273 , n35184 , n35185 , n6276 , n35187 , n35188 , n6279 , n35190 , n35191 , n6282 , 
 n35193 , n35194 , n6285 , n35196 , n35197 , n6288 , n35199 , n35200 , n35201 , n35202 , 
 n6293 , n35204 , n35205 , n6296 , n35207 , n35208 , n6299 , n35210 , n35211 , n6302 , 
 n35213 , n35214 , n6305 , n35216 , n35217 , n6308 , n6309 , n6310 , n35221 , n35222 , 
 n35223 , n35224 , n6315 , n35226 , n35227 , n35228 , n35229 , n6320 , n35231 , n35232 , 
 n6323 , n6324 , n35235 , n35236 , n6327 , n6328 , n6329 , n35240 , n35241 , n6332 , 
 n6333 , n6334 , n35245 , n35246 , n6337 , n6338 , n6339 , n35250 , n35251 , n6342 , 
 n35253 , n35254 , n6345 , n35256 , n6347 , n6348 , n35259 , n35260 , n6351 , n6352 , 
 n35263 , n35264 , n6355 , n6356 , n35267 , n35268 , n6359 , n6360 , n6361 , n6362 , 
 n6363 , n35274 , n35275 , n6366 , n6367 , n6368 , n35279 , n35280 , n6371 , n6372 , 
 n6373 , n35284 , n35285 , n6376 , n6377 , n6378 , n35289 , n6380 , n6381 , n6382 , 
 n6383 , n6384 , n6385 , n35296 , n6387 , n6388 , n6389 , n6390 , n35301 , n35302 , 
 n35303 , n6394 , n6395 , n35306 , n35307 , n35308 , n6402 , n6403 , n35311 , n35312 , 
 n6409 , n6410 , n6411 , n6412 , n35317 , n35318 , n6415 , n6416 , n6417 , n6418 , 
 n6419 , n35324 , n35325 , n6422 , n35327 , n35328 , n6425 , n35330 , n35331 , n6428 , 
 n6429 , n6430 , n6431 , n35336 , n35337 , n6434 , n6435 , n6436 , n6437 , n6438 , 
 n35343 , n35344 , n35345 , n35346 , n6443 , n35348 , n35349 , n35350 , n35351 , n6448 , 
 n35353 , n35354 , n6451 , n35356 , n35357 , n6454 , n35359 , n35360 , n6457 , n35362 , 
 n35363 , n6460 , n35365 , n35366 , n6463 , n35368 , n35369 , n35370 , n35371 , n6468 , 
 n35373 , n35374 , n6471 , n35376 , n35377 , n6474 , n35379 , n35380 , n6477 , n35382 , 
 n35383 , n6480 , n35385 , n35386 , n35387 , n35388 , n6485 , n35390 , n35391 , n35392 , 
 n35393 , n6490 , n35395 , n35396 , n6493 , n35398 , n35399 , n6496 , n35401 , n35402 , 
 n6499 , n35404 , n35405 , n6502 , n6503 , n6504 , n6505 , n35410 , n35411 , n6508 , 
 n35413 , n35414 , n6511 , n35416 , n35417 , n35418 , n35419 , n6516 , n35421 , n35422 , 
 n6519 , n35424 , n35425 , n35426 , n6523 , n35428 , n35429 , n6526 , n35431 , n35432 , 
 n6529 , n35434 , n35435 , n6532 , n35437 , n35438 , n6535 , n6536 , n6537 , n35442 , 
 n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n6548 , n35450 , n35451 , n6554 , 
 n6555 , n6556 , n6557 , n35456 , n35457 , n6560 , n6561 , n35460 , n35461 , n6564 , 
 n6565 , n6566 , n6567 , n35466 , n35467 , n6570 , n6571 , n6572 , n35471 , n35472 , 
 n6575 , n6576 , n6577 , n35476 , n35477 , n6580 , n35479 , n35480 , n6583 , n6584 , 
 n6585 , n35484 , n35485 , n6588 , n6589 , n6590 , n6591 , n35490 , n35491 , n6594 , 
 n35493 , n35494 , n6597 , n35496 , n6599 , n35498 , n6601 , n6602 , n35501 , n6604 , 
 n35503 , n35504 , n6607 , n6608 , n35507 , n35508 , n6611 , n35510 , n35511 , n6614 , 
 n35513 , n35514 , n6617 , n6618 , n35517 , n35518 , n6621 , n35520 , n35521 , n6624 , 
 n35523 , n6626 , n6627 , n6628 , n35527 , n35528 , n6631 , n35530 , n6633 , n6634 , 
 n35533 , n35534 , n6637 , n35536 , n6639 , n6640 , n35539 , n6642 , n6643 , n6644 , 
 n6645 , n6646 , n35545 , n35546 , n6649 , n6650 , n6651 , n6652 , n35551 , n35552 , 
 n6655 , n6656 , n6657 , n6658 , n35557 , n35558 , n6661 , n35560 , n35561 , n6664 , 
 n35563 , n35564 , n35565 , n35566 , n6669 , n35568 , n35569 , n6672 , n35571 , n35572 , 
 n6675 , n35574 , n35575 , n6678 , n35577 , n35578 , n6681 , n35580 , n35581 , n6684 , 
 n35583 , n35584 , n6690 , n35586 , n35587 , n35588 , n35589 , n6698 , n35591 , n35592 , 
 n6701 , n35594 , n35595 , n6704 , n35597 , n35598 , n6707 , n35600 , n35601 , n35602 , 
 n35603 , n6712 , n35605 , n35606 , n35607 , n35608 , n6717 , n35610 , n35611 , n6720 , 
 n35613 , n35614 , n6723 , n35616 , n35617 , n6726 , n35619 , n35620 , n6729 , n35622 , 
 n35623 , n6732 , n35625 , n35626 , n35627 , n35628 , n6737 , n35630 , n35631 , n6740 , 
 n35633 , n35634 , n6743 , n35636 , n35637 , n6746 , n35639 , n35640 , n6749 , n35642 , 
 n35643 , n6752 , n35645 , n35646 , n6755 , n6756 , n6757 , n6758 , n35651 , n35652 , 
 n6761 , n6762 , n35655 , n6764 , n6765 , n35658 , n35659 , n6768 , n6769 , n6770 , 
 n6771 , n35664 , n35665 , n6774 , n6775 , n6776 , n6777 , n6778 , n35671 , n35672 , 
 n6781 , n6782 , n6783 , n6784 , n35677 , n35678 , n6787 , n35680 , n35681 , n35682 , 
 n6791 , n35684 , n35685 , n6794 , n35687 , n35688 , n6797 , n35690 , n35691 , n6800 , 
 n6801 , n6802 , n6803 , n6804 , n35697 , n35698 , n6807 , n35700 , n35701 , n6810 , 
 n35703 , n35704 , n6813 , n35706 , n35707 , n6816 , n35709 , n35710 , n35711 , n35712 , 
 n6821 , n6822 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n6836 , 
 n35723 , n35724 , n6839 , n35726 , n35727 , n6842 , n6843 , n35730 , n35731 , n6846 , 
 n6847 , n35734 , n6849 , n6850 , n6851 , n6852 , n6853 , n35740 , n35741 , n6856 , 
 n35743 , n6858 , n6859 , n6860 , n6861 , n6862 , n35749 , n6864 , n35751 , n6866 , 
 n35753 , n6868 , n35755 , n6870 , n6871 , n6872 , n6873 , n35760 , n6875 , n35762 , 
 n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , 
 n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n35782 , 
 n6897 , n6898 , n35785 , n6900 , n35787 , n35788 , n6903 , n35790 , n35791 , n35792 , 
 n6907 , n35794 , n6909 , n35796 , n6911 , n35798 , n6913 , n6914 , n6915 , n6916 , 
 n6917 , n6918 , n6919 , n35806 , n6921 , n6922 , n35809 , n6924 , n6925 , n6926 , 
 n6927 , n35814 , n6929 , n35816 , n6931 , n35818 , n35819 , n6934 , n35821 , n6936 , 
 n6937 , n6938 , n35825 , n6940 , n6941 , n6942 , n6943 , n6944 , n35831 , n35832 , 
 n35833 , n35834 , n35835 , n35836 , n6954 , n35838 , n6956 , n6957 , n35841 , n6962 , 
 n6963 , n6964 , n6965 , n35846 , n6967 , n35848 , n6969 , n6970 , n6971 , n6972 , 
 n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , 
 n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n35871 , n6992 , 
 n35873 , n6994 , n35875 , n35876 , n6997 , n35878 , n6999 , n7000 , n7001 , n7002 , 
 n7003 , n7004 , n7005 , n7006 , n7007 , n35888 , n35889 , n7010 , n35891 , n7012 , 
 n35893 , n7014 , n7015 , n35896 , n35897 , n35898 , n7019 , n7020 , n7021 , n7022 , 
 n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , 
 n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , 
 n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , 
 n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , 
 n35943 , n35944 , n7065 , n7066 , n35947 , n7071 , n35949 , n7073 , n7074 , n35952 , 
 n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , 
 n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , 
 n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , 
 n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , 
 n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , 
 n7129 , n36004 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , 
 n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , 
 n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , 
 n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , 
 n7169 , n36044 , n36045 , n7172 , n7173 , n36048 , n7178 , n36050 , n7180 , n7181 , 
 n36053 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , 
 n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , 
 n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , 
 n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , 
 n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n36099 , n7232 , n7233 , n7234 , 
 n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , 
 n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , 
 n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , 
 n7265 , n7266 , n36135 , n36136 , n7269 , n7270 , n36139 , n7275 , n36141 , n7277 , 
 n7278 , n36144 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , 
 n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , 
 n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , 
 n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , 
 n7321 , n7322 , n7323 , n36186 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , 
 n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , 
 n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , 
 n7351 , n7352 , n7353 , n36216 , n7355 , n36218 , n7360 , n36220 , n7362 , n7363 , 
 n36223 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , 
 n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , 
 n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , 
 n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n36259 , n7404 , n7405 , n7406 , 
 n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n36269 , n7414 , n36271 , n7416 , 
 n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , 
 n7427 , n7428 , n36285 , n7433 , n36287 , n7435 , n7436 , n36290 , n7441 , n7442 , 
 n36293 , n7444 , n36295 , n7446 , n36297 , n7448 , n36299 , n7450 , n36301 , n36302 , 
 n7453 , n36304 , n7455 , n36306 , n7457 , n7458 , n36309 , n7460 , n36311 , n7462 , 
 n36313 , n36314 , n7465 , n36316 , n7467 , n7468 , n36319 , n36320 , n36321 , n36322 , 
 n36323 , n7474 , n7475 , n36326 , n36327 , n36328 , n7479 , n36330 , n36331 , n7482 , 
 n36333 , n7484 , n7485 , n7486 , n36337 , n36338 , n7489 , n36340 , n36341 , n36342 , 
 n7496 , n36344 , n7498 , n7499 , n36347 , n36348 , n7505 , n36350 , n36351 , n7508 , 
 n36353 , n36354 , n7511 , n36356 , n7513 , n36358 , n7515 , n7516 , n36361 , n36362 , 
 n36363 , n7520 , n36365 , n36366 , n7523 , n36368 , n36369 , n7526 , n36371 , n36372 , 
 n36373 , n36374 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n36382 , 
 n7539 , n36384 , n7541 , n36386 , n36387 , n7547 , n36389 , n7549 , n7550 , n36392 , 
 n7555 , n7556 , n36395 , n7558 , n36397 , n7560 , n7561 , n36400 , n7563 , n36402 , 
 n7565 , n36404 , n36405 , n7568 , n36407 , n7570 , n7571 , n7572 , n7573 , n7574 , 
 n7575 , n36414 , n7577 , n7578 , n36417 , n7583 , n7584 , n7585 , n36421 , n7587 , 
 n7588 , n7589 , n7590 , n36426 , n36427 , n7593 , n7594 , n7595 , n7596 , n7597 , 
 n36433 , n36434 , n7603 , n36436 , n36437 , n36438 , n7610 , n36440 , n36441 , n7613 , 
 n36443 , n36444 , n36445 , n7620 , n36447 , n7622 , n7623 , n36450 , n36451 , n36452 , 
 n36453 , n36454 , n36455 , n36456 , n7637 , n7638 , n36459 , n7640 , n36461 , n36462 , 
 n7646 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , 
 n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , 
 n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , 
 n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , 
 n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , 
 n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , 
 n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , 
 n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , 
 n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , 
 n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , 
 n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , 
 n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , 
 n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , 
 n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , 
 n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , 
 n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , 
 n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , 
 n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , 
 n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , 
 n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , 
 n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , 
 n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , 
 n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , 
 n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , 
 n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , 
 n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , 
 n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , 
 n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , 
 n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , 
 n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , 
 n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , 
 n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , 
 n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , 
 n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , 
 n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , 
 n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , 
 n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , 
 n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , 
 n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , 
 n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , 
 n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , 
 n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , 
 n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , 
 n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , 
 n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , 
 n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , 
 n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , 
 n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , 
 n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , 
 n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , 
 n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , 
 n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , 
 n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , 
 n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , 
 n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , 
 n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , 
 n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , 
 n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , 
 n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , 
 n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , 
 n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , 
 n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , 
 n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , 
 n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , 
 n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , 
 n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , 
 n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , 
 n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , 
 n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , 
 n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , 
 n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , 
 n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , 
 n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , 
 n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , 
 n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , 
 n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , 
 n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , 
 n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , 
 n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , 
 n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , 
 n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , 
 n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , 
 n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , 
 n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , 
 n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , 
 n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , 
 n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , 
 n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , 
 n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , 
 n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , 
 n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , 
 n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , 
 n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , 
 n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , 
 n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , 
 n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , 
 n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , 
 n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , 
 n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , 
 n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , 
 n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , 
 n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , 
 n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , 
 n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , 
 n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , 
 n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , 
 n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , 
 n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , 
 n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , 
 n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , 
 n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , 
 n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , 
 n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , 
 n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , 
 n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , 
 n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , 
 n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , 
 n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , 
 n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , 
 n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , 
 n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , 
 n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , 
 n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , 
 n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , 
 n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , 
 n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , 
 n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , 
 n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , 
 n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , 
 n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , 
 n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , 
 n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , 
 n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , 
 n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , 
 n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , 
 n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , 
 n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , 
 n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , 
 n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , 
 n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , 
 n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , 
 n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , 
 n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , 
 n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , 
 n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , 
 n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , 
 n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , 
 n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , 
 n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , 
 n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , 
 n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , 
 n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , 
 n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , 
 n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , 
 n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , 
 n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , 
 n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , 
 n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , 
 n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , 
 n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , 
 n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , 
 n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , 
 n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , 
 n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , 
 n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , 
 n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , 
 n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , 
 n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , 
 n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , 
 n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , 
 n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , 
 n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , 
 n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , 
 n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , 
 n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , 
 n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , 
 n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , 
 n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , 
 n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , 
 n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , 
 n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , 
 n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , 
 n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , 
 n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , 
 n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , 
 n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , 
 n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , 
 n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , 
 n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , 
 n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , 
 n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , 
 n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , 
 n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , 
 n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , 
 n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , 
 n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , 
 n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , 
 n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , 
 n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , 
 n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , 
 n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , 
 n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , 
 n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , 
 n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , 
 n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , 
 n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , 
 n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , 
 n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , 
 n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , 
 n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , 
 n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , 
 n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , 
 n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , 
 n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , 
 n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , 
 n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , 
 n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , 
 n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , 
 n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , 
 n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , 
 n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , 
 n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , 
 n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , 
 n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , 
 n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , 
 n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , 
 n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , 
 n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , 
 n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , 
 n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , 
 n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , 
 n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , 
 n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , 
 n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , 
 n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , 
 n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , 
 n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , 
 n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , 
 n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , 
 n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , 
 n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , 
 n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , 
 n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , 
 n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , 
 n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , 
 n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , 
 n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , 
 n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , 
 n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , 
 n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , 
 n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , 
 n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , 
 n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , 
 n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , 
 n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , 
 n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , 
 n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , 
 n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , 
 n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , 
 n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , 
 n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , 
 n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , 
 n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , 
 n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , 
 n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , 
 n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , 
 n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , 
 n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , 
 n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , 
 n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , 
 n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , 
 n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , 
 n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , 
 n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , 
 n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , 
 n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , 
 n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , 
 n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , 
 n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , 
 n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , 
 n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , 
 n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , 
 n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , 
 n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , 
 n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , 
 n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , 
 n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , 
 n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , 
 n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , 
 n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , 
 n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , 
 n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , 
 n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , 
 n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , 
 n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , 
 n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , 
 n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , 
 n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , 
 n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , 
 n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , 
 n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , 
 n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , 
 n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , 
 n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , 
 n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , 
 n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , 
 n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , 
 n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , 
 n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , 
 n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , 
 n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , 
 n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , 
 n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , 
 n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , 
 n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , 
 n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , 
 n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , 
 n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , 
 n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , 
 n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , 
 n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , 
 n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , 
 n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , 
 n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , 
 n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , 
 n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , 
 n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , 
 n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , 
 n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , 
 n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , 
 n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , 
 n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , 
 n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , 
 n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , 
 n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , 
 n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , 
 n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , 
 n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , 
 n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , 
 n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , 
 n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , 
 n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , 
 n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , 
 n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , 
 n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , 
 n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , 
 n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , 
 n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , 
 n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , 
 n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , 
 n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , 
 n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , 
 n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , 
 n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , 
 n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , 
 n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , 
 n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , 
 n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , 
 n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , 
 n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , 
 n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , 
 n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , 
 n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , 
 n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , 
 n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , 
 n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , 
 n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , 
 n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , 
 n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , 
 n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , 
 n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , 
 n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , 
 n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , 
 n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , 
 n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , 
 n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , 
 n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , 
 n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , 
 n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , 
 n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , 
 n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , 
 n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , 
 n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , 
 n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , 
 n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , 
 n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , 
 n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , 
 n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , 
 n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , 
 n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , 
 n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , 
 n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , 
 n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , 
 n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , 
 n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , 
 n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , 
 n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , 
 n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , 
 n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , 
 n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , 
 n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , 
 n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , 
 n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , 
 n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , 
 n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , 
 n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , 
 n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , 
 n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , 
 n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , 
 n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , 
 n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , 
 n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , 
 n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , 
 n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , 
 n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , 
 n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , 
 n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , 
 n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , 
 n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , 
 n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , 
 n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , 
 n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , 
 n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , 
 n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , 
 n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , 
 n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , 
 n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , 
 n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , 
 n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , 
 n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , 
 n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , 
 n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , 
 n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , 
 n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , 
 n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , 
 n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , 
 n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , 
 n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , 
 n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , 
 n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , 
 n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , 
 n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , 
 n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , 
 n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , 
 n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , 
 n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , 
 n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , 
 n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , 
 n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , 
 n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , 
 n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , 
 n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , 
 n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , 
 n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , 
 n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , 
 n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , 
 n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , 
 n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , 
 n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , 
 n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , 
 n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , 
 n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , 
 n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , 
 n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , 
 n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , 
 n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , 
 n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , 
 n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , 
 n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , 
 n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , 
 n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , 
 n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , 
 n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , 
 n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , 
 n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , 
 n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , 
 n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , 
 n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , 
 n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , 
 n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , 
 n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , 
 n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , 
 n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , 
 n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , 
 n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , 
 n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , 
 n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , 
 n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , 
 n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , 
 n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , 
 n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , 
 n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , 
 n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , 
 n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , 
 n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , 
 n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , 
 n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , 
 n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , 
 n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , 
 n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , 
 n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , 
 n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , 
 n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , 
 n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , 
 n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , 
 n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , 
 n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , 
 n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , 
 n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , 
 n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , 
 n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , 
 n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , 
 n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , 
 n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , 
 n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , 
 n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , 
 n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , 
 n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , 
 n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , 
 n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , 
 n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , 
 n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , 
 n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , 
 n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , 
 n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , 
 n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , 
 n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , 
 n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , 
 n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , 
 n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , 
 n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , 
 n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , 
 n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , 
 n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , 
 n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , 
 n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , 
 n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , 
 n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , 
 n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , 
 n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , 
 n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , 
 n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , 
 n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , 
 n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , 
 n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , 
 n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , 
 n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , 
 n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , 
 n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , 
 n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , 
 n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , 
 n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , 
 n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , 
 n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , 
 n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , 
 n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , 
 n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , 
 n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , 
 n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , 
 n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , 
 n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , 
 n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , 
 n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , 
 n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , 
 n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , 
 n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , 
 n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , 
 n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , 
 n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , 
 n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , 
 n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , 
 n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , 
 n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , 
 n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , 
 n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , 
 n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , 
 n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , 
 n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , 
 n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , 
 n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , 
 n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , 
 n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , 
 n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , 
 n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , 
 n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , 
 n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , 
 n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , 
 n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , 
 n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , 
 n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , 
 n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , 
 n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , 
 n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , 
 n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , 
 n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , 
 n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , 
 n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , 
 n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , 
 n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , 
 n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , 
 n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , 
 n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , 
 n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , 
 n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , 
 n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , 
 n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , 
 n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , 
 n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , 
 n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , 
 n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , 
 n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , 
 n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , 
 n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , 
 n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , 
 n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , 
 n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , 
 n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , 
 n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , 
 n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , 
 n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , 
 n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , 
 n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , 
 n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , 
 n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , 
 n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , 
 n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , 
 n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , 
 n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , 
 n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , 
 n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , 
 n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , 
 n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , 
 n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , 
 n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , 
 n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , 
 n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , 
 n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , 
 n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , 
 n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , 
 n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , 
 n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , 
 n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , 
 n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , 
 n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , 
 n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , 
 n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , 
 n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , 
 n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , 
 n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , 
 n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , 
 n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , 
 n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , 
 n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , 
 n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , 
 n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , 
 n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , 
 n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , 
 n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , 
 n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , 
 n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , 
 n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , 
 n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , 
 n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , 
 n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , 
 n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , 
 n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , 
 n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , 
 n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , 
 n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , 
 n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , 
 n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , 
 n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , 
 n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , 
 n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , 
 n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , 
 n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , 
 n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , 
 n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , 
 n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , 
 n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , 
 n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , 
 n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , 
 n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , 
 n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , 
 n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , 
 n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , 
 n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , 
 n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , 
 n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , 
 n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , 
 n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , 
 n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , 
 n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , 
 n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , 
 n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , 
 n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , 
 n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , 
 n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , 
 n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , 
 n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , 
 n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , 
 n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , 
 n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , 
 n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , 
 n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , 
 n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , 
 n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , 
 n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , 
 n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , 
 n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , 
 n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , 
 n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , 
 n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , 
 n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , 
 n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , 
 n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , 
 n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , 
 n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , 
 n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , 
 n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , 
 n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , 
 n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , 
 n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , 
 n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , 
 n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , 
 n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , 
 n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , 
 n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , 
 n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , 
 n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , 
 n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , 
 n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , 
 n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , 
 n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , 
 n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , 
 n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , 
 n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , 
 n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , 
 n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , 
 n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , 
 n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , 
 n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , 
 n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , 
 n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , 
 n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , 
 n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , 
 n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , 
 n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , 
 n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , 
 n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , 
 n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , 
 n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , 
 n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , 
 n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , 
 n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , 
 n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , 
 n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , 
 n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , 
 n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , 
 n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , 
 n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , 
 n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , 
 n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , 
 n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , 
 n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , 
 n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , 
 n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , 
 n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , 
 n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , 
 n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , 
 n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , 
 n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , 
 n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , 
 n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , 
 n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , 
 n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , 
 n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , 
 n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , 
 n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , 
 n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , 
 n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , 
 n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , 
 n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , 
 n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , 
 n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , 
 n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , 
 n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , 
 n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , 
 n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , 
 n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , 
 n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , 
 n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , 
 n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , 
 n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , 
 n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , 
 n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , 
 n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , 
 n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , 
 n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , 
 n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , 
 n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , 
 n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , 
 n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , 
 n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , 
 n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , 
 n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , 
 n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , 
 n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , 
 n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , 
 n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , 
 n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , 
 n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , 
 n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , 
 n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , 
 n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , 
 n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , 
 n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , 
 n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , 
 n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , 
 n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , 
 n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , 
 n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , 
 n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , 
 n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , 
 n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , 
 n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , 
 n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , 
 n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , 
 n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , 
 n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , 
 n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , 
 n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , 
 n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , 
 n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , 
 n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , 
 n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , 
 n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , 
 n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , 
 n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , 
 n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , 
 n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , 
 n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , 
 n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , 
 n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , 
 n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , 
 n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , 
 n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , 
 n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , 
 n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , 
 n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , 
 n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , 
 n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , 
 n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , 
 n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , 
 n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , 
 n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , 
 n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , 
 n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , 
 n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , 
 n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , 
 n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , 
 n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , 
 n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , 
 n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , 
 n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , 
 n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , 
 n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , 
 n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , 
 n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , 
 n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , 
 n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , 
 n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , 
 n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , 
 n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , 
 n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , 
 n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , 
 n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , 
 n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , 
 n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , 
 n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , 
 n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , 
 n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , 
 n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , 
 n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , 
 n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , 
 n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , 
 n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , 
 n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , 
 n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , 
 n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , 
 n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , 
 n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , 
 n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , 
 n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , 
 n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , 
 n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , 
 n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , 
 n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , 
 n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , 
 n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , 
 n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , 
 n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , 
 n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , 
 n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , 
 n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , 
 n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , 
 n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , 
 n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , 
 n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , 
 n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , 
 n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , 
 n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , 
 n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , 
 n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , 
 n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , 
 n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , 
 n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , 
 n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , 
 n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , 
 n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , 
 n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , 
 n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , 
 n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , 
 n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , 
 n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , 
 n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , 
 n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , 
 n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , 
 n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , 
 n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , 
 n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , 
 n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , 
 n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , 
 n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , 
 n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , 
 n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , 
 n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , 
 n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , 
 n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , 
 n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , 
 n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , 
 n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , 
 n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , 
 n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , 
 n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , 
 n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , 
 n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , 
 n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , 
 n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , 
 n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , 
 n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , 
 n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , 
 n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , 
 n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , 
 n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , 
 n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , 
 n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , 
 n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , 
 n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , 
 n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , 
 n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , 
 n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , 
 n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , 
 n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , 
 n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , 
 n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , 
 n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , 
 n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , 
 n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , 
 n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , 
 n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , 
 n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , 
 n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , 
 n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , 
 n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , 
 n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , 
 n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , 
 n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , 
 n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , 
 n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , 
 n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , 
 n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , 
 n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , 
 n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , 
 n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , 
 n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , 
 n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , 
 n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , 
 n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , 
 n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , 
 n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , 
 n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , 
 n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , 
 n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , 
 n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , 
 n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , 
 n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , 
 n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , 
 n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , 
 n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , 
 n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , 
 n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , 
 n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , 
 n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , 
 n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , 
 n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , 
 n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , 
 n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , 
 n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , 
 n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , 
 n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , 
 n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , 
 n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , 
 n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , 
 n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , 
 n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , 
 n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , 
 n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , 
 n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , 
 n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , 
 n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , 
 n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , 
 n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , 
 n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , C0n , 
 C0 , C1n , C1 ;
buf ( n454 , n0 );
buf ( n455 , n1 );
buf ( n456 , n2 );
buf ( n457 , n3 );
buf ( n458 , n4 );
buf ( n459 , n5 );
buf ( n460 , n6 );
buf ( n461 , n7 );
buf ( n462 , n8 );
buf ( n463 , n9 );
buf ( n464 , n10 );
buf ( n465 , n11 );
buf ( n466 , n12 );
buf ( n467 , n13 );
buf ( n468 , n14 );
buf ( n469 , n15 );
buf ( n470 , n16 );
buf ( n471 , n17 );
buf ( n472 , n18 );
buf ( n473 , n19 );
buf ( n474 , n20 );
buf ( n475 , n21 );
buf ( n476 , n22 );
buf ( n477 , n23 );
buf ( n478 , n24 );
buf ( n479 , n25 );
buf ( n480 , n26 );
buf ( n481 , n27 );
buf ( n482 , n28 );
buf ( n483 , n29 );
buf ( n484 , n30 );
buf ( n485 , n31 );
buf ( n486 , n32 );
buf ( n487 , n33 );
buf ( n488 , n34 );
buf ( n489 , n35 );
buf ( n490 , n36 );
buf ( n491 , n37 );
buf ( n492 , n38 );
buf ( n493 , n39 );
buf ( n494 , n40 );
buf ( n495 , n41 );
buf ( n496 , n42 );
buf ( n497 , n43 );
buf ( n498 , n44 );
buf ( n499 , n45 );
buf ( n500 , n46 );
buf ( n501 , n47 );
buf ( n502 , n48 );
buf ( n503 , n49 );
buf ( n504 , n50 );
buf ( n505 , n51 );
buf ( n506 , n52 );
buf ( n507 , n53 );
buf ( n508 , n54 );
buf ( n509 , n55 );
buf ( n510 , n56 );
buf ( n511 , n57 );
buf ( n512 , n58 );
buf ( n513 , n59 );
buf ( n514 , n60 );
buf ( n515 , n61 );
buf ( n516 , n62 );
buf ( n517 , n63 );
buf ( n518 , n64 );
buf ( n519 , n65 );
buf ( n520 , n66 );
buf ( n521 , n67 );
buf ( n522 , n68 );
buf ( n523 , n69 );
buf ( n524 , n70 );
buf ( n525 , n71 );
buf ( n526 , n72 );
buf ( n527 , n73 );
buf ( n528 , n74 );
buf ( n529 , n75 );
buf ( n530 , n76 );
buf ( n531 , n77 );
buf ( n532 , n78 );
buf ( n533 , n79 );
buf ( n534 , n80 );
buf ( n535 , n81 );
buf ( n536 , n82 );
buf ( n537 , n83 );
buf ( n538 , n84 );
buf ( n539 , n85 );
buf ( n540 , n86 );
buf ( n541 , n87 );
buf ( n542 , n88 );
buf ( n543 , n89 );
buf ( n544 , n90 );
buf ( n545 , n91 );
buf ( n546 , n92 );
buf ( n547 , n93 );
buf ( n548 , n94 );
buf ( n549 , n95 );
buf ( n550 , n96 );
buf ( n551 , n97 );
buf ( n552 , n98 );
buf ( n99 , n553 );
buf ( n100 , n554 );
buf ( n101 , n555 );
buf ( n102 , n556 );
buf ( n103 , n557 );
buf ( n104 , n558 );
buf ( n105 , n559 );
buf ( n106 , n560 );
buf ( n107 , n561 );
buf ( n108 , n562 );
buf ( n109 , n563 );
buf ( n110 , n564 );
buf ( n111 , n565 );
buf ( n112 , n566 );
buf ( n113 , n567 );
buf ( n114 , n568 );
buf ( n115 , n569 );
buf ( n116 , n570 );
buf ( n117 , n571 );
buf ( n118 , n572 );
buf ( n119 , n573 );
buf ( n120 , n574 );
buf ( n121 , n575 );
buf ( n122 , n576 );
buf ( n123 , n577 );
buf ( n124 , n578 );
buf ( n125 , n579 );
buf ( n126 , n580 );
buf ( n127 , n581 );
buf ( n128 , n582 );
buf ( n129 , n583 );
buf ( n130 , n584 );
buf ( n131 , n585 );
buf ( n132 , n586 );
buf ( n133 , n587 );
buf ( n134 , n588 );
buf ( n135 , n589 );
buf ( n136 , n590 );
buf ( n137 , n591 );
buf ( n138 , n592 );
buf ( n139 , n593 );
buf ( n140 , n594 );
buf ( n141 , n595 );
buf ( n142 , n596 );
buf ( n143 , n597 );
buf ( n144 , n598 );
buf ( n145 , n599 );
buf ( n146 , n600 );
buf ( n147 , n601 );
buf ( n148 , n602 );
buf ( n149 , n603 );
buf ( n150 , n604 );
buf ( n151 , n605 );
buf ( n152 , n606 );
buf ( n153 , n607 );
buf ( n154 , n608 );
buf ( n155 , n609 );
buf ( n156 , n610 );
buf ( n157 , n611 );
buf ( n158 , n612 );
buf ( n159 , n613 );
buf ( n160 , n614 );
buf ( n161 , n615 );
buf ( n162 , n616 );
buf ( n163 , n617 );
buf ( n164 , n618 );
buf ( n165 , n619 );
buf ( n166 , n620 );
buf ( n167 , n621 );
buf ( n168 , n622 );
buf ( n169 , n623 );
buf ( n170 , n624 );
buf ( n171 , n625 );
buf ( n172 , n626 );
buf ( n173 , n627 );
buf ( n174 , n628 );
buf ( n175 , n629 );
buf ( n176 , n630 );
buf ( n177 , n631 );
buf ( n178 , n632 );
buf ( n179 , n633 );
buf ( n180 , n634 );
buf ( n181 , n635 );
buf ( n182 , n636 );
buf ( n183 , n637 );
buf ( n184 , n638 );
buf ( n185 , n639 );
buf ( n186 , n640 );
buf ( n187 , n641 );
buf ( n188 , n642 );
buf ( n189 , n643 );
buf ( n190 , n644 );
buf ( n191 , n645 );
buf ( n192 , n646 );
buf ( n193 , n647 );
buf ( n194 , n648 );
buf ( n195 , n649 );
buf ( n196 , n650 );
buf ( n197 , n651 );
buf ( n198 , n652 );
buf ( n199 , n653 );
buf ( n200 , n654 );
buf ( n201 , n655 );
buf ( n202 , n656 );
buf ( n203 , n657 );
buf ( n204 , n658 );
buf ( n205 , n659 );
buf ( n206 , n660 );
buf ( n207 , n661 );
buf ( n208 , n662 );
buf ( n209 , n663 );
buf ( n210 , n664 );
buf ( n211 , n665 );
buf ( n212 , n666 );
buf ( n213 , n667 );
buf ( n214 , n668 );
buf ( n215 , n669 );
buf ( n216 , n670 );
buf ( n217 , n671 );
buf ( n218 , n672 );
buf ( n219 , n673 );
buf ( n220 , n674 );
buf ( n221 , n675 );
buf ( n222 , n676 );
buf ( n223 , n677 );
buf ( n224 , n678 );
buf ( n225 , n679 );
buf ( n226 , n680 );
buf ( n553 , n46573 );
buf ( n554 , n46573 );
buf ( n555 , n46573 );
buf ( n556 , n46573 );
buf ( n557 , n46573 );
buf ( n558 , n46573 );
buf ( n559 , n46573 );
buf ( n560 , n46573 );
buf ( n561 , n46573 );
buf ( n562 , n46573 );
buf ( n563 , n46573 );
buf ( n564 , n46573 );
buf ( n565 , n46573 );
buf ( n566 , n46573 );
buf ( n567 , n46573 );
buf ( n568 , n46573 );
buf ( n569 , n46573 );
buf ( n570 , n46573 );
buf ( n571 , n46573 );
buf ( n572 , n46573 );
buf ( n573 , n46573 );
buf ( n574 , n46573 );
buf ( n575 , n46573 );
buf ( n576 , n46573 );
buf ( n577 , n46573 );
buf ( n578 , n46573 );
buf ( n579 , n46573 );
buf ( n580 , n46573 );
buf ( n581 , n46573 );
buf ( n582 , n46573 );
buf ( n583 , n46573 );
buf ( n584 , n46324 );
buf ( n585 , n46309 );
buf ( n586 , n46315 );
buf ( n587 , n46366 );
buf ( n588 , n46500 );
buf ( n589 , n46258 );
buf ( n590 , n46348 );
buf ( n591 , n46388 );
buf ( n592 , n46440 );
buf ( n593 , n46361 );
buf ( n594 , n46426 );
buf ( n595 , n42171 );
buf ( n596 , n46430 );
buf ( n597 , n40912 );
buf ( n598 , n42881 );
buf ( n599 , n42908 );
buf ( n600 , n42883 );
buf ( n601 , n41080 );
buf ( n602 , n40975 );
buf ( n603 , n36959 );
buf ( n604 , n6851 );
buf ( n605 , n6962 );
buf ( n606 , n44747 );
buf ( n607 , n6884 );
buf ( n608 , n7039 );
buf ( n609 , n6979 );
buf ( n610 , n7022 );
buf ( n611 , n2358 );
buf ( n612 , n43477 );
buf ( n613 , n46644 );
buf ( n614 , n46649 );
buf ( n615 , n46663 );
buf ( n616 , n46658 );
buf ( n617 , C0 );
buf ( n618 , C0 );
buf ( n619 , C0 );
buf ( n620 , C0 );
buf ( n621 , C0 );
buf ( n622 , C0 );
buf ( n623 , C0 );
buf ( n624 , n46652 );
buf ( n625 , n46549 );
buf ( n626 , n46549 );
buf ( n627 , n46549 );
buf ( n628 , n46549 );
buf ( n629 , n46549 );
buf ( n630 , n46549 );
buf ( n631 , n46549 );
buf ( n632 , n46549 );
buf ( n633 , n46549 );
buf ( n634 , n46549 );
buf ( n635 , n46549 );
buf ( n636 , n46549 );
buf ( n637 , n46549 );
buf ( n638 , n46549 );
buf ( n639 , n46549 );
buf ( n640 , n46549 );
buf ( n641 , n46549 );
buf ( n642 , n46549 );
buf ( n643 , n46549 );
buf ( n644 , n46549 );
buf ( n645 , n46549 );
buf ( n646 , n46549 );
buf ( n647 , n46549 );
buf ( n648 , n46549 );
buf ( n649 , n46549 );
buf ( n650 , n46549 );
buf ( n651 , n46677 );
buf ( n652 , n46489 );
buf ( n653 , n46547 );
buf ( n654 , n46379 );
buf ( n655 , n46520 );
buf ( n656 , n46571 );
buf ( n657 , n46562 );
buf ( n658 , n46405 );
buf ( n659 , n46396 );
buf ( n660 , n46455 );
buf ( n661 , n46445 );
buf ( n662 , n46560 );
buf ( n663 , n46613 );
buf ( n664 , n42877 );
buf ( n665 , n46602 );
buf ( n666 , n42905 );
buf ( n667 , n46690 );
buf ( n668 , n42919 );
buf ( n669 , n42931 );
buf ( n670 , n46701 );
buf ( n671 , n46629 );
buf ( n672 , n37044 );
buf ( n673 , n7409 );
buf ( n674 , n46639 );
buf ( n675 , n46634 );
buf ( n676 , n46694 );
buf ( n677 , n43494 );
buf ( n678 , n46618 );
buf ( n679 , n46653 );
buf ( n680 , n46538 );
and ( n29489 , n456 , n461 );
not ( n29490 , n456 );
and ( n29491 , n29490 , n477 );
nor ( n29492 , n29489 , n29491 );
not ( n29493 , n29492 );
buf ( n29494 , n29493 );
not ( n29495 , n464 );
and ( n29496 , n456 , n29495 );
not ( n29497 , n456 );
not ( n29498 , n480 );
and ( n29499 , n29497 , n29498 );
nor ( n29500 , n29496 , n29499 );
buf ( n29501 , n29500 );
buf ( n29502 , n29501 );
and ( n29503 , n456 , n468 );
not ( n29504 , n456 );
and ( n29505 , n29504 , n484 );
nor ( n29506 , n29503 , n29505 );
not ( n29507 , n29506 );
buf ( n29508 , n29507 );
and ( n29509 , n456 , n470 );
not ( n29510 , n456 );
and ( n29511 , n29510 , n486 );
nor ( n29512 , n29509 , n29511 );
not ( n29513 , n29512 );
buf ( n29514 , n29513 );
not ( n29515 , n488 );
or ( n29516 , n29515 , n456 );
nand ( n29517 , n456 , n472 );
nand ( n29518 , n29516 , n29517 );
not ( n29519 , n455 );
not ( n29520 , n29519 );
buf ( n29521 , n499 );
buf ( n29522 , n519 );
xor ( n29523 , n29521 , n29522 );
buf ( n29524 , n29523 );
buf ( n29525 , n29524 );
not ( n29526 , n29525 );
xor ( n29527 , n501 , n500 );
not ( n29528 , n29527 );
not ( n29529 , n500 );
not ( n29530 , n499 );
and ( n29531 , n29529 , n29530 );
and ( n29532 , n500 , n499 );
nor ( n29533 , n29531 , n29532 );
nand ( n29534 , n29528 , n29533 );
not ( n29535 , n29534 );
buf ( n29536 , n29535 );
not ( n29537 , n29536 );
or ( n29538 , n29526 , n29537 );
buf ( n29539 , n500 );
buf ( n29540 , n501 );
xor ( n29541 , n29539 , n29540 );
buf ( n29542 , n29541 );
buf ( n29543 , n29542 );
buf ( n29544 , n29543 );
buf ( n29545 , n518 );
buf ( n29546 , n499 );
xor ( n29547 , n29545 , n29546 );
buf ( n29548 , n29547 );
buf ( n29549 , n29548 );
nand ( n29550 , n29544 , n29549 );
buf ( n29551 , n29550 );
buf ( n29552 , n29551 );
nand ( n29553 , n29538 , n29552 );
buf ( n29554 , n29553 );
buf ( n29555 , n29554 );
buf ( n29556 , n520 );
buf ( n29557 , n500 );
or ( n29558 , n29556 , n29557 );
buf ( n29559 , n501 );
nand ( n29560 , n29558 , n29559 );
buf ( n29561 , n29560 );
buf ( n29562 , n29561 );
buf ( n29563 , n520 );
buf ( n29564 , n500 );
nand ( n29565 , n29563 , n29564 );
buf ( n29566 , n29565 );
buf ( n29567 , n29566 );
buf ( n29568 , n499 );
and ( n29569 , n29562 , n29567 , n29568 );
buf ( n29570 , n29569 );
buf ( n29571 , n29570 );
buf ( n29572 , n516 );
buf ( n29573 , n503 );
xor ( n29574 , n29572 , n29573 );
buf ( n29575 , n29574 );
buf ( n29576 , n29575 );
not ( n29577 , n29576 );
not ( n29578 , n504 );
nand ( n29579 , n29578 , n503 );
buf ( n29580 , n29579 );
not ( n29581 , n29580 );
buf ( n29582 , n29581 );
buf ( n29583 , n29582 );
not ( n29584 , n29583 );
or ( n29585 , n29577 , n29584 );
buf ( n29586 , n515 );
buf ( n29587 , n503 );
xor ( n29588 , n29586 , n29587 );
buf ( n29589 , n29588 );
buf ( n29590 , n29589 );
buf ( n29591 , n504 );
nand ( n29592 , n29590 , n29591 );
buf ( n29593 , n29592 );
buf ( n29594 , n29593 );
nand ( n29595 , n29585 , n29594 );
buf ( n29596 , n29595 );
buf ( n29597 , n29596 );
and ( n29598 , n29571 , n29597 );
buf ( n29599 , n29598 );
buf ( n29600 , n29599 );
xor ( n29601 , n29555 , n29600 );
xor ( n29602 , n498 , n499 );
not ( n29603 , n29602 );
not ( n29604 , n29603 );
buf ( n29605 , n29604 );
buf ( n29606 , n520 );
and ( n29607 , n29605 , n29606 );
buf ( n29608 , n29607 );
buf ( n29609 , n29608 );
buf ( n29610 , n29589 );
not ( n29611 , n29610 );
buf ( n29612 , n29582 );
not ( n29613 , n29612 );
or ( n29614 , n29611 , n29613 );
xor ( n29615 , n503 , n514 );
buf ( n29616 , n29615 );
buf ( n29617 , n504 );
nand ( n29618 , n29616 , n29617 );
buf ( n29619 , n29618 );
buf ( n29620 , n29619 );
nand ( n29621 , n29614 , n29620 );
buf ( n29622 , n29621 );
buf ( n29623 , n29622 );
xor ( n29624 , n29609 , n29623 );
buf ( n29625 , n501 );
buf ( n29626 , n517 );
xor ( n29627 , n29625 , n29626 );
buf ( n29628 , n29627 );
buf ( n29629 , n29628 );
not ( n29630 , n29629 );
buf ( n29631 , n502 );
buf ( n29632 , n503 );
xor ( n29633 , n29631 , n29632 );
buf ( n29634 , n29633 );
buf ( n29635 , n29634 );
not ( n29636 , n29635 );
buf ( n29637 , n29636 );
xor ( n29638 , n502 , n501 );
nand ( n29639 , n29637 , n29638 );
not ( n29640 , n29639 );
buf ( n29641 , n29640 );
not ( n29642 , n29641 );
or ( n29643 , n29630 , n29642 );
buf ( n29644 , n29637 );
not ( n29645 , n29644 );
buf ( n29646 , n29645 );
buf ( n29647 , n29646 );
buf ( n29648 , n29647 );
buf ( n29649 , n29648 );
buf ( n29650 , n29649 );
buf ( n29651 , n516 );
buf ( n29652 , n501 );
xor ( n29653 , n29651 , n29652 );
buf ( n29654 , n29653 );
buf ( n29655 , n29654 );
nand ( n29656 , n29650 , n29655 );
buf ( n29657 , n29656 );
buf ( n29658 , n29657 );
nand ( n29659 , n29643 , n29658 );
buf ( n29660 , n29659 );
buf ( n29661 , n29660 );
xor ( n29662 , n29624 , n29661 );
buf ( n29663 , n29662 );
buf ( n29664 , n29663 );
xor ( n29665 , n29601 , n29664 );
buf ( n29666 , n29665 );
buf ( n29667 , n501 );
buf ( n29668 , n518 );
xor ( n29669 , n29667 , n29668 );
buf ( n29670 , n29669 );
buf ( n29671 , n29670 );
not ( n29672 , n29671 );
buf ( n29673 , n29640 );
not ( n29674 , n29673 );
or ( n29675 , n29672 , n29674 );
buf ( n29676 , n29649 );
buf ( n29677 , n29628 );
nand ( n29678 , n29676 , n29677 );
buf ( n29679 , n29678 );
buf ( n29680 , n29679 );
nand ( n29681 , n29675 , n29680 );
buf ( n29682 , n29681 );
buf ( n29683 , n29682 );
buf ( n29684 , n499 );
buf ( n29685 , n520 );
and ( n29686 , n29684 , n29685 );
not ( n29687 , n29684 );
buf ( n29688 , n520 );
not ( n29689 , n29688 );
buf ( n29690 , n29689 );
buf ( n29691 , n29690 );
and ( n29692 , n29687 , n29691 );
nor ( n29693 , n29686 , n29692 );
buf ( n29694 , n29693 );
buf ( n29695 , n29694 );
not ( n29696 , n29695 );
buf ( n29697 , n29535 );
not ( n29698 , n29697 );
or ( n29699 , n29696 , n29698 );
buf ( n29700 , n29543 );
buf ( n29701 , n29524 );
nand ( n29702 , n29700 , n29701 );
buf ( n29703 , n29702 );
buf ( n29704 , n29703 );
nand ( n29705 , n29699 , n29704 );
buf ( n29706 , n29705 );
buf ( n29707 , n29706 );
xor ( n29708 , n29683 , n29707 );
xor ( n29709 , n29571 , n29597 );
buf ( n29710 , n29709 );
buf ( n29711 , n29710 );
and ( n29712 , n29708 , n29711 );
and ( n29713 , n29683 , n29707 );
or ( n29714 , n29712 , n29713 );
buf ( n29715 , n29714 );
nor ( n29716 , n29666 , n29715 );
not ( n29717 , n29716 );
and ( n29718 , n29666 , n29715 );
not ( n29719 , n29718 );
nand ( n29720 , n29717 , n29719 );
not ( n29721 , n29720 );
buf ( n29722 , n29543 );
buf ( n29723 , n520 );
and ( n29724 , n29722 , n29723 );
buf ( n29725 , n29724 );
buf ( n29726 , n29725 );
buf ( n29727 , n503 );
buf ( n29728 , n517 );
xor ( n29729 , n29727 , n29728 );
buf ( n29730 , n29729 );
buf ( n29731 , n29730 );
not ( n29732 , n29731 );
not ( n29733 , n503 );
nor ( n29734 , n29733 , n504 );
buf ( n29735 , n29734 );
not ( n29736 , n29735 );
or ( n29737 , n29732 , n29736 );
buf ( n29738 , n29575 );
buf ( n29739 , n504 );
nand ( n29740 , n29738 , n29739 );
buf ( n29741 , n29740 );
buf ( n29742 , n29741 );
nand ( n29743 , n29737 , n29742 );
buf ( n29744 , n29743 );
buf ( n29745 , n29744 );
xor ( n29746 , n29726 , n29745 );
buf ( n29747 , n501 );
buf ( n29748 , n519 );
xor ( n29749 , n29747 , n29748 );
buf ( n29750 , n29749 );
buf ( n29751 , n29750 );
not ( n29752 , n29751 );
buf ( n29753 , n29640 );
not ( n29754 , n29753 );
or ( n29755 , n29752 , n29754 );
buf ( n29756 , n29649 );
buf ( n29757 , n29670 );
nand ( n29758 , n29756 , n29757 );
buf ( n29759 , n29758 );
buf ( n29760 , n29759 );
nand ( n29761 , n29755 , n29760 );
buf ( n29762 , n29761 );
buf ( n29763 , n29762 );
and ( n29764 , n29746 , n29763 );
and ( n29765 , n29726 , n29745 );
or ( n29766 , n29764 , n29765 );
buf ( n29767 , n29766 );
xor ( n29768 , n29683 , n29707 );
xor ( n29769 , n29768 , n29711 );
buf ( n29770 , n29769 );
xor ( n29771 , n29767 , n29770 );
xor ( n29772 , n29726 , n29745 );
xor ( n29773 , n29772 , n29763 );
buf ( n29774 , n29773 );
not ( n29775 , n29774 );
buf ( n29776 , n520 );
buf ( n29777 , n502 );
or ( n29778 , n29776 , n29777 );
buf ( n29779 , n503 );
nand ( n29780 , n29778 , n29779 );
buf ( n29781 , n29780 );
buf ( n29782 , n29781 );
buf ( n29783 , n520 );
buf ( n29784 , n502 );
nand ( n29785 , n29783 , n29784 );
buf ( n29786 , n29785 );
buf ( n29787 , n29786 );
buf ( n29788 , n501 );
and ( n29789 , n29782 , n29787 , n29788 );
buf ( n29790 , n29789 );
buf ( n29791 , n29790 );
buf ( n29792 , n503 );
buf ( n29793 , n518 );
xor ( n29794 , n29792 , n29793 );
buf ( n29795 , n29794 );
buf ( n29796 , n29795 );
not ( n29797 , n29796 );
buf ( n29798 , n29734 );
not ( n29799 , n29798 );
or ( n29800 , n29797 , n29799 );
buf ( n29801 , n29730 );
buf ( n29802 , n504 );
nand ( n29803 , n29801 , n29802 );
buf ( n29804 , n29803 );
buf ( n29805 , n29804 );
nand ( n29806 , n29800 , n29805 );
buf ( n29807 , n29806 );
buf ( n29808 , n29807 );
and ( n29809 , n29791 , n29808 );
buf ( n29810 , n29809 );
not ( n29811 , n29810 );
nand ( n29812 , n29775 , n29811 );
not ( n29813 , n29812 );
xor ( n29814 , n29791 , n29808 );
buf ( n29815 , n29814 );
buf ( n29816 , n29750 );
not ( n29817 , n29816 );
buf ( n29818 , n29649 );
not ( n29819 , n29818 );
or ( n29820 , n29817 , n29819 );
buf ( n29821 , n29640 );
buf ( n29822 , n501 );
buf ( n29823 , n520 );
and ( n29824 , n29822 , n29823 );
not ( n684 , n29822 );
buf ( n29826 , n29690 );
and ( n686 , n684 , n29826 );
nor ( n687 , n29824 , n686 );
buf ( n29829 , n687 );
buf ( n29830 , n29829 );
nand ( n690 , n29821 , n29830 );
buf ( n29832 , n690 );
buf ( n29833 , n29832 );
nand ( n693 , n29820 , n29833 );
buf ( n29835 , n693 );
nor ( n695 , n29815 , n29835 );
buf ( n29837 , n503 );
buf ( n29838 , n519 );
xor ( n698 , n29837 , n29838 );
buf ( n29840 , n698 );
buf ( n29841 , n29840 );
not ( n701 , n29841 );
buf ( n29843 , n29582 );
not ( n703 , n29843 );
or ( n29845 , n701 , n703 );
buf ( n29846 , n29795 );
buf ( n29847 , n504 );
nand ( n707 , n29846 , n29847 );
buf ( n29849 , n707 );
buf ( n29850 , n29849 );
nand ( n29851 , n29845 , n29850 );
buf ( n29852 , n29851 );
buf ( n29853 , n29649 );
buf ( n29854 , n520 );
and ( n714 , n29853 , n29854 );
buf ( n29856 , n714 );
or ( n716 , n29852 , n29856 );
or ( n717 , n29734 , n29840 );
and ( n718 , n717 , n29690 , n503 );
and ( n719 , n716 , n718 );
and ( n720 , n29852 , n29856 );
nor ( n721 , n719 , n720 );
or ( n722 , n695 , n721 );
nand ( n723 , n29815 , n29835 );
nand ( n724 , n722 , n723 );
not ( n725 , n724 );
or ( n726 , n29813 , n725 );
nand ( n727 , n29774 , n29810 );
nand ( n728 , n726 , n727 );
and ( n729 , n29771 , n728 );
and ( n730 , n29767 , n29770 );
or ( n731 , n729 , n730 );
not ( n732 , n731 );
or ( n733 , n29721 , n732 );
or ( n734 , n731 , n29720 );
nand ( n735 , n733 , n734 );
not ( n736 , n735 );
or ( n29878 , n29520 , n736 );
and ( n741 , n500 , n501 );
not ( n29880 , n500 );
not ( n743 , n501 );
and ( n29882 , n29880 , n743 );
nor ( n745 , n741 , n29882 );
buf ( n29884 , n745 );
buf ( n29885 , n29884 );
not ( n748 , n29885 );
buf ( n29887 , n499 );
not ( n750 , n29887 );
buf ( n29889 , n29513 );
not ( n752 , n29889 );
buf ( n29891 , n752 );
buf ( n29892 , n29891 );
not ( n758 , n29892 );
or ( n29894 , n750 , n758 );
buf ( n29895 , n29513 );
not ( n761 , n29895 );
buf ( n29897 , n761 );
not ( n763 , n29897 );
buf ( n29899 , n499 );
not ( n765 , n29899 );
buf ( n29901 , n765 );
nand ( n770 , n763 , n29901 );
buf ( n29903 , n770 );
nand ( n772 , n29894 , n29903 );
buf ( n29905 , n772 );
buf ( n29906 , n29905 );
not ( n775 , n29906 );
or ( n776 , n748 , n775 );
and ( n777 , n456 , n471 );
not ( n778 , n456 );
and ( n782 , n778 , n487 );
nor ( n29912 , n777 , n782 );
not ( n784 , n29912 );
buf ( n29914 , n784 );
not ( n786 , n29914 );
buf ( n29916 , n786 );
and ( n788 , n29916 , n499 );
not ( n789 , n29916 );
and ( n790 , n789 , n29901 );
or ( n791 , n788 , n790 );
buf ( n29921 , n791 );
buf ( n29922 , n500 );
buf ( n29923 , n501 );
xnor ( n795 , n29922 , n29923 );
buf ( n29925 , n795 );
xor ( n797 , n500 , n499 );
nand ( n798 , n29925 , n797 );
not ( n799 , n798 );
buf ( n29929 , n799 );
buf ( n801 , n29929 );
buf ( n29931 , n801 );
buf ( n29932 , n29931 );
nand ( n804 , n29921 , n29932 );
buf ( n29934 , n804 );
buf ( n29935 , n29934 );
nand ( n807 , n776 , n29935 );
buf ( n29937 , n807 );
buf ( n29938 , n29937 );
buf ( n29939 , n29518 );
buf ( n29940 , n29939 );
not ( n815 , n29940 );
buf ( n29942 , n815 );
buf ( n29943 , n29942 );
not ( n818 , n29943 );
buf ( n29945 , n818 );
buf ( n29946 , n29945 );
buf ( n29947 , n500 );
or ( n822 , n29946 , n29947 );
buf ( n29949 , n501 );
nand ( n824 , n822 , n29949 );
buf ( n29951 , n824 );
buf ( n29952 , n29939 );
not ( n827 , n29952 );
buf ( n29954 , n827 );
buf ( n29955 , n29954 );
not ( n830 , n29955 );
buf ( n29957 , n830 );
and ( n832 , n29957 , n500 );
nor ( n833 , n832 , n29901 );
and ( n834 , n29951 , n833 );
buf ( n29961 , n834 );
buf ( n29962 , n503 );
not ( n29963 , n29962 );
buf ( n29964 , n504 );
nor ( n842 , n29963 , n29964 );
buf ( n29966 , n842 );
buf ( n29967 , n29966 );
buf ( n845 , n29967 );
buf ( n29969 , n845 );
buf ( n29970 , n29969 );
not ( n848 , n29970 );
buf ( n29972 , n503 );
not ( n850 , n29972 );
and ( n851 , n456 , n468 );
not ( n852 , n456 );
and ( n29976 , n852 , n484 );
nor ( n854 , n851 , n29976 );
buf ( n29978 , n854 );
not ( n856 , n29978 );
or ( n857 , n850 , n856 );
buf ( n29981 , n854 );
not ( n859 , n29981 );
buf ( n29983 , n859 );
buf ( n29984 , n29983 );
buf ( n29985 , n503 );
not ( n863 , n29985 );
buf ( n29987 , n863 );
buf ( n29988 , n29987 );
nand ( n869 , n29984 , n29988 );
buf ( n29990 , n869 );
buf ( n29991 , n29990 );
nand ( n872 , n857 , n29991 );
buf ( n29993 , n872 );
buf ( n29994 , n29993 );
not ( n875 , n29994 );
or ( n876 , n848 , n875 );
buf ( n29997 , n503 );
not ( n878 , n29997 );
and ( n879 , n456 , n467 );
not ( n30000 , n456 );
and ( n881 , n30000 , n483 );
nor ( n882 , n879 , n881 );
buf ( n30003 , n882 );
not ( n884 , n30003 );
or ( n885 , n878 , n884 );
buf ( n30006 , n882 );
not ( n887 , n30006 );
buf ( n30008 , n887 );
buf ( n30009 , n30008 );
buf ( n30010 , n29987 );
nand ( n891 , n30009 , n30010 );
buf ( n30012 , n891 );
buf ( n30013 , n30012 );
nand ( n894 , n885 , n30013 );
buf ( n30015 , n894 );
buf ( n30016 , n30015 );
buf ( n30017 , n504 );
nand ( n898 , n30016 , n30017 );
buf ( n30019 , n898 );
buf ( n30020 , n30019 );
nand ( n901 , n876 , n30020 );
buf ( n30022 , n901 );
buf ( n30023 , n30022 );
and ( n904 , n29961 , n30023 );
buf ( n30025 , n904 );
buf ( n30026 , n30025 );
xor ( n907 , n29938 , n30026 );
buf ( n30028 , n29945 );
xor ( n909 , n498 , n499 );
buf ( n910 , n909 );
buf ( n30031 , n910 );
and ( n30032 , n30028 , n30031 );
buf ( n30033 , n30032 );
buf ( n30034 , n30033 );
buf ( n30035 , n29969 );
not ( n919 , n30035 );
buf ( n30037 , n30015 );
not ( n30038 , n30037 );
or ( n922 , n919 , n30038 );
buf ( n30040 , n504 );
buf ( n30041 , n503 );
not ( n925 , n30041 );
and ( n926 , n456 , n466 );
not ( n927 , n456 );
and ( n928 , n927 , n482 );
nor ( n929 , n926 , n928 );
buf ( n30047 , n929 );
not ( n931 , n30047 );
or ( n932 , n925 , n931 );
not ( n933 , n929 );
buf ( n30051 , n933 );
buf ( n30052 , n29987 );
nand ( n936 , n30051 , n30052 );
buf ( n30054 , n936 );
buf ( n30055 , n30054 );
nand ( n939 , n932 , n30055 );
buf ( n30057 , n939 );
buf ( n30058 , n30057 );
nand ( n942 , n30040 , n30058 );
buf ( n30060 , n942 );
buf ( n30061 , n30060 );
nand ( n945 , n922 , n30061 );
buf ( n30063 , n945 );
buf ( n30064 , n30063 );
xor ( n951 , n30034 , n30064 );
not ( n952 , n503 );
not ( n953 , n502 );
not ( n954 , n953 );
or ( n955 , n952 , n954 );
not ( n956 , n503 );
nand ( n957 , n956 , n502 );
nand ( n30072 , n955 , n957 );
not ( n959 , n30072 );
xor ( n960 , n502 , n501 );
nand ( n961 , n959 , n960 );
buf ( n30076 , n961 );
not ( n963 , n30076 );
buf ( n30078 , n963 );
buf ( n30079 , n30078 );
not ( n966 , n30079 );
buf ( n30081 , n501 );
not ( n30082 , n30081 );
and ( n969 , n456 , n469 );
not ( n970 , n456 );
and ( n971 , n970 , n485 );
nor ( n972 , n969 , n971 );
not ( n973 , n972 );
buf ( n30088 , n973 );
not ( n975 , n30088 );
buf ( n30090 , n975 );
buf ( n30091 , n30090 );
not ( n978 , n30091 );
or ( n979 , n30082 , n978 );
buf ( n30094 , n30090 );
not ( n981 , n30094 );
buf ( n30096 , n981 );
buf ( n30097 , n30096 );
not ( n984 , n501 );
buf ( n30099 , n984 );
nand ( n986 , n30097 , n30099 );
buf ( n30101 , n986 );
buf ( n30102 , n30101 );
nand ( n989 , n979 , n30102 );
buf ( n30104 , n989 );
buf ( n30105 , n30104 );
not ( n30106 , n30105 );
or ( n996 , n966 , n30106 );
buf ( n30108 , n501 );
not ( n998 , n30108 );
buf ( n30110 , n854 );
not ( n1000 , n30110 );
or ( n1001 , n998 , n1000 );
buf ( n30113 , n29983 );
buf ( n30114 , n984 );
nand ( n1004 , n30113 , n30114 );
buf ( n30116 , n1004 );
buf ( n30117 , n30116 );
nand ( n1007 , n1001 , n30117 );
buf ( n30119 , n1007 );
buf ( n30120 , n30119 );
buf ( n1010 , n30072 );
buf ( n30122 , n1010 );
nand ( n1012 , n30120 , n30122 );
buf ( n30124 , n1012 );
buf ( n30125 , n30124 );
nand ( n1015 , n996 , n30125 );
buf ( n30127 , n1015 );
buf ( n30128 , n30127 );
xor ( n1018 , n951 , n30128 );
buf ( n30130 , n1018 );
buf ( n30131 , n30130 );
xor ( n1024 , n907 , n30131 );
buf ( n30133 , n1024 );
not ( n30134 , n29884 );
not ( n1027 , n791 );
or ( n1028 , n30134 , n1027 );
buf ( n30137 , n499 );
not ( n1030 , n30137 );
buf ( n30139 , n29954 );
not ( n30140 , n30139 );
buf ( n30141 , n30140 );
buf ( n30142 , n30141 );
not ( n1035 , n30142 );
buf ( n30144 , n1035 );
buf ( n30145 , n30144 );
not ( n1038 , n30145 );
or ( n1039 , n1030 , n1038 );
buf ( n30148 , n30144 );
not ( n1041 , n30148 );
buf ( n30150 , n1041 );
buf ( n30151 , n30150 );
buf ( n30152 , n29901 );
nand ( n1045 , n30151 , n30152 );
buf ( n30154 , n1045 );
buf ( n30155 , n30154 );
nand ( n1048 , n1039 , n30155 );
buf ( n30157 , n1048 );
buf ( n30158 , n30157 );
buf ( n30159 , n29931 );
nand ( n1052 , n30158 , n30159 );
buf ( n30161 , n1052 );
nand ( n1054 , n1028 , n30161 );
buf ( n30163 , n501 );
not ( n1056 , n30163 );
buf ( n30165 , n29897 );
not ( n1058 , n30165 );
or ( n1059 , n1056 , n1058 );
buf ( n30168 , n29897 );
not ( n1061 , n30168 );
buf ( n30170 , n1061 );
buf ( n30171 , n30170 );
buf ( n30172 , n984 );
nand ( n1065 , n30171 , n30172 );
buf ( n30174 , n1065 );
buf ( n30175 , n30174 );
nand ( n1068 , n1059 , n30175 );
buf ( n30177 , n1068 );
buf ( n30178 , n30177 );
not ( n30179 , n30178 );
buf ( n30180 , n30078 );
not ( n1073 , n30180 );
or ( n1074 , n30179 , n1073 );
buf ( n30183 , n30104 );
buf ( n30184 , n1010 );
nand ( n1077 , n30183 , n30184 );
buf ( n30186 , n1077 );
buf ( n30187 , n30186 );
nand ( n1080 , n1074 , n30187 );
buf ( n30189 , n1080 );
xor ( n1085 , n1054 , n30189 );
xor ( n30191 , n29961 , n30023 );
buf ( n30192 , n30191 );
and ( n1088 , n1085 , n30192 );
and ( n1089 , n1054 , n30189 );
or ( n1090 , n1088 , n1089 );
nor ( n1091 , n30133 , n1090 );
not ( n30197 , n1091 );
and ( n1093 , n30133 , n1090 );
not ( n1094 , n1093 );
nand ( n1095 , n30197 , n1094 );
not ( n1096 , n1095 );
xor ( n1097 , n1054 , n30189 );
xor ( n1098 , n1097 , n30192 );
not ( n1099 , n1098 );
buf ( n30205 , n29945 );
buf ( n30206 , n29884 );
and ( n1102 , n30205 , n30206 );
buf ( n30208 , n1102 );
buf ( n30209 , n504 );
not ( n1105 , n30209 );
buf ( n30211 , n29993 );
not ( n1107 , n30211 );
or ( n1108 , n1105 , n1107 );
buf ( n30214 , n503 );
not ( n1110 , n30214 );
buf ( n30216 , n30090 );
not ( n1112 , n30216 );
or ( n1113 , n1110 , n1112 );
buf ( n30219 , n30096 );
buf ( n30220 , n29987 );
nand ( n1116 , n30219 , n30220 );
buf ( n30222 , n1116 );
buf ( n30223 , n30222 );
nand ( n1119 , n1113 , n30223 );
buf ( n30225 , n1119 );
buf ( n30226 , n30225 );
buf ( n30227 , n29969 );
nand ( n1126 , n30226 , n30227 );
buf ( n30229 , n1126 );
buf ( n30230 , n30229 );
nand ( n1129 , n1108 , n30230 );
buf ( n30232 , n1129 );
xor ( n1131 , n30208 , n30232 );
buf ( n30234 , n1010 );
not ( n1133 , n30234 );
buf ( n30236 , n30177 );
not ( n1135 , n30236 );
or ( n30238 , n1133 , n1135 );
buf ( n30239 , n501 );
not ( n1138 , n30239 );
buf ( n30241 , n29916 );
not ( n1140 , n30241 );
or ( n1141 , n1138 , n1140 );
buf ( n30244 , n29916 );
not ( n1143 , n30244 );
buf ( n30246 , n1143 );
buf ( n30247 , n30246 );
buf ( n30248 , n984 );
nand ( n1147 , n30247 , n30248 );
buf ( n30250 , n1147 );
buf ( n30251 , n30250 );
nand ( n1150 , n1141 , n30251 );
buf ( n30253 , n1150 );
buf ( n30254 , n30253 );
buf ( n30255 , n30078 );
nand ( n1154 , n30254 , n30255 );
buf ( n30257 , n1154 );
buf ( n30258 , n30257 );
nand ( n1157 , n30238 , n30258 );
buf ( n30260 , n1157 );
and ( n1159 , n1131 , n30260 );
and ( n1160 , n30208 , n30232 );
or ( n1161 , n1159 , n1160 );
not ( n1162 , n1161 );
nand ( n1163 , n1099 , n1162 );
buf ( n30266 , n30150 );
buf ( n30267 , n502 );
and ( n1166 , n30266 , n30267 );
buf ( n30269 , n984 );
nor ( n1168 , n1166 , n30269 );
buf ( n30271 , n1168 );
buf ( n30272 , n30271 );
buf ( n30273 , n29957 );
buf ( n30274 , n502 );
or ( n1173 , n30273 , n30274 );
buf ( n30276 , n503 );
nand ( n1175 , n1173 , n30276 );
buf ( n30278 , n1175 );
buf ( n30279 , n30278 );
and ( n1178 , n30272 , n30279 );
buf ( n30281 , n1178 );
buf ( n30282 , n30281 );
buf ( n30283 , n29969 );
not ( n1182 , n30283 );
buf ( n30285 , n503 );
not ( n1187 , n30285 );
buf ( n30287 , n29897 );
not ( n1189 , n30287 );
or ( n1190 , n1187 , n1189 );
buf ( n30290 , n30170 );
buf ( n30291 , n29987 );
nand ( n1193 , n30290 , n30291 );
buf ( n30293 , n1193 );
buf ( n30294 , n30293 );
nand ( n1196 , n1190 , n30294 );
buf ( n30296 , n1196 );
buf ( n30297 , n30296 );
not ( n1199 , n30297 );
or ( n1200 , n1182 , n1199 );
buf ( n30300 , n30225 );
buf ( n30301 , n504 );
nand ( n1203 , n30300 , n30301 );
buf ( n30303 , n1203 );
buf ( n30304 , n30303 );
nand ( n1206 , n1200 , n30304 );
buf ( n30306 , n1206 );
buf ( n30307 , n30306 );
xor ( n1209 , n30282 , n30307 );
buf ( n30309 , n1209 );
buf ( n30310 , n30078 );
not ( n1212 , n30310 );
buf ( n30312 , n984 );
buf ( n30313 , n30144 );
and ( n1215 , n30312 , n30313 );
not ( n1216 , n30312 );
buf ( n30316 , n30150 );
and ( n1221 , n1216 , n30316 );
nor ( n1222 , n1215 , n1221 );
buf ( n30319 , n1222 );
buf ( n30320 , n30319 );
not ( n1225 , n30320 );
or ( n1226 , n1212 , n1225 );
buf ( n30323 , n30253 );
buf ( n30324 , n1010 );
nand ( n1229 , n30323 , n30324 );
buf ( n30326 , n1229 );
buf ( n30327 , n30326 );
nand ( n1232 , n1226 , n30327 );
buf ( n30329 , n1232 );
nor ( n1234 , n30309 , n30329 );
and ( n1235 , n30150 , n1010 );
buf ( n30332 , n503 );
not ( n30333 , n30332 );
buf ( n30334 , n29916 );
not ( n1239 , n30334 );
or ( n1240 , n30333 , n1239 );
buf ( n30337 , n30246 );
buf ( n30338 , n29987 );
nand ( n1243 , n30337 , n30338 );
buf ( n30340 , n1243 );
buf ( n30341 , n30340 );
nand ( n1246 , n1240 , n30341 );
buf ( n30343 , n1246 );
not ( n1248 , n30343 );
buf ( n30345 , n29969 );
not ( n1250 , n30345 );
buf ( n30347 , n1250 );
nand ( n1252 , n1248 , n30347 );
nor ( n1253 , n30150 , n29987 );
and ( n1254 , n1252 , n1253 );
or ( n1255 , n1235 , n1254 );
buf ( n30352 , n504 );
not ( n1257 , n30352 );
buf ( n30354 , n30296 );
not ( n1259 , n30354 );
or ( n1260 , n1257 , n1259 );
buf ( n30357 , n29969 );
buf ( n30358 , n30343 );
nand ( n1263 , n30357 , n30358 );
buf ( n30360 , n1263 );
buf ( n30361 , n30360 );
nand ( n1266 , n1260 , n30361 );
buf ( n30363 , n1266 );
nand ( n1268 , n1255 , n30363 );
or ( n1269 , n1234 , n1268 );
nand ( n1270 , n30309 , n30329 );
nand ( n1271 , n1269 , n1270 );
not ( n1272 , n1271 );
xor ( n1273 , n30208 , n30232 );
xor ( n1274 , n1273 , n30260 );
not ( n1275 , n1274 );
and ( n1276 , n30282 , n30307 );
buf ( n30373 , n1276 );
not ( n30374 , n30373 );
nand ( n1279 , n1275 , n30374 );
not ( n1280 , n1279 );
or ( n1281 , n1272 , n1280 );
nand ( n1282 , n1274 , n30373 );
nand ( n1283 , n1281 , n1282 );
nand ( n1284 , n1163 , n1283 );
nand ( n1285 , n1161 , n1098 );
nand ( n1286 , n1284 , n1285 );
buf ( n1287 , n1286 );
not ( n1288 , n1287 );
or ( n1289 , n1096 , n1288 );
or ( n1290 , n1095 , n1287 );
nand ( n1291 , n1289 , n1290 );
nand ( n30388 , n1291 , n455 );
nand ( n1293 , n29878 , n30388 );
buf ( n30390 , n1293 );
buf ( n30391 , n549 );
or ( n1296 , n30390 , n30391 );
buf ( n30393 , n1296 );
buf ( n30394 , n30393 );
not ( n1299 , n30394 );
buf ( n30396 , n551 );
not ( n1301 , n455 );
nand ( n1302 , n1279 , n1282 );
buf ( n1303 , n1271 );
not ( n1304 , n1303 );
and ( n1305 , n1302 , n1304 );
not ( n1309 , n1302 );
and ( n30403 , n1309 , n1303 );
nor ( n1311 , n1305 , n30403 );
not ( n1312 , n1311 );
or ( n1313 , n1301 , n1312 );
nand ( n1314 , n29812 , n727 );
xnor ( n1315 , n1314 , n724 );
nand ( n1316 , n29519 , n1315 );
nand ( n1317 , n1313 , n1316 );
buf ( n30411 , n1317 );
xor ( n1319 , n30396 , n30411 );
buf ( n30413 , n552 );
not ( n1321 , n29519 );
not ( n1322 , n695 );
nand ( n1323 , n1322 , n723 );
xor ( n1324 , n721 , n1323 );
not ( n1325 , n1324 );
or ( n1326 , n1321 , n1325 );
not ( n1327 , n1234 );
nand ( n1328 , n1327 , n1270 );
and ( n1329 , n1328 , n1268 );
not ( n1330 , n1328 );
not ( n1331 , n1268 );
and ( n1332 , n1330 , n1331 );
nor ( n1333 , n1329 , n1332 );
nand ( n1334 , n1333 , n455 );
nand ( n1335 , n1326 , n1334 );
buf ( n30429 , n1335 );
and ( n1337 , n30413 , n30429 );
buf ( n30431 , n1337 );
buf ( n30432 , n30431 );
and ( n1343 , n1319 , n30432 );
and ( n1344 , n30396 , n30411 );
or ( n1345 , n1343 , n1344 );
buf ( n30436 , n1345 );
buf ( n30437 , n30436 );
not ( n30438 , n29519 );
xor ( n1349 , n29767 , n29770 );
xor ( n1350 , n1349 , n728 );
not ( n1351 , n1350 );
or ( n1352 , n30438 , n1351 );
xor ( n1353 , n1161 , n1098 );
xor ( n1354 , n1353 , n1283 );
nand ( n1355 , n1354 , n455 );
nand ( n1356 , n1352 , n1355 );
buf ( n30447 , n1356 );
buf ( n30448 , n550 );
or ( n1359 , n30447 , n30448 );
buf ( n30450 , n1359 );
buf ( n30451 , n30450 );
and ( n1362 , n30437 , n30451 );
buf ( n30453 , n1362 );
buf ( n30454 , n30453 );
not ( n1365 , n30454 );
or ( n1366 , n1299 , n1365 );
buf ( n30457 , n30393 );
buf ( n30458 , n550 );
buf ( n30459 , n1356 );
nand ( n1370 , n30458 , n30459 );
buf ( n30461 , n1370 );
buf ( n30462 , n30461 );
not ( n1373 , n30462 );
buf ( n30464 , n1373 );
buf ( n30465 , n30464 );
and ( n1376 , n30457 , n30465 );
buf ( n30467 , n1293 );
buf ( n30468 , n549 );
and ( n30469 , n30467 , n30468 );
buf ( n30470 , n30469 );
buf ( n30471 , n30470 );
nor ( n1382 , n1376 , n30471 );
buf ( n30473 , n1382 );
buf ( n30474 , n30473 );
nand ( n1385 , n1366 , n30474 );
buf ( n30476 , n1385 );
buf ( n30477 , n30476 );
not ( n1388 , n30197 );
not ( n1389 , n1287 );
or ( n1390 , n1388 , n1389 );
nand ( n1391 , n1390 , n1094 );
buf ( n30482 , n29969 );
not ( n1393 , n30482 );
buf ( n30484 , n30057 );
not ( n30485 , n30484 );
or ( n1396 , n1393 , n30485 );
buf ( n30487 , n503 );
not ( n1398 , n30487 );
and ( n1399 , n456 , n465 );
not ( n1400 , n456 );
and ( n1401 , n1400 , n481 );
nor ( n1402 , n1399 , n1401 );
not ( n1403 , n1402 );
buf ( n30494 , n1403 );
not ( n1405 , n30494 );
buf ( n30496 , n1405 );
buf ( n30497 , n30496 );
not ( n1411 , n30497 );
or ( n1412 , n1398 , n1411 );
buf ( n30500 , n1403 );
buf ( n30501 , n29987 );
nand ( n1415 , n30500 , n30501 );
buf ( n30503 , n1415 );
buf ( n30504 , n30503 );
nand ( n1418 , n1412 , n30504 );
buf ( n30506 , n1418 );
buf ( n30507 , n30506 );
buf ( n30508 , n504 );
nand ( n1422 , n30507 , n30508 );
buf ( n30510 , n1422 );
buf ( n30511 , n30510 );
nand ( n1425 , n1396 , n30511 );
buf ( n30513 , n1425 );
buf ( n30514 , n30513 );
buf ( n30515 , n498 );
not ( n1429 , n30515 );
buf ( n30517 , n30144 );
nand ( n1431 , n1429 , n30517 );
buf ( n30519 , n1431 );
buf ( n30520 , n30519 );
buf ( n30521 , n499 );
and ( n1435 , n30520 , n30521 );
buf ( n30523 , n498 );
not ( n1437 , n30523 );
buf ( n30525 , n29957 );
not ( n1439 , n30525 );
or ( n30527 , n1437 , n1439 );
buf ( n30528 , n497 );
nand ( n1442 , n30527 , n30528 );
buf ( n30530 , n1442 );
buf ( n30531 , n30530 );
nor ( n1445 , n1435 , n30531 );
buf ( n30533 , n1445 );
buf ( n30534 , n30533 );
xor ( n1448 , n30514 , n30534 );
buf ( n30536 , n1448 );
buf ( n30537 , n30536 );
xor ( n1451 , n30034 , n30064 );
and ( n1452 , n1451 , n30128 );
and ( n1453 , n30034 , n30064 );
or ( n30541 , n1452 , n1453 );
buf ( n30542 , n30541 );
buf ( n30543 , n30542 );
xor ( n1460 , n30537 , n30543 );
buf ( n30545 , n29931 );
not ( n1462 , n30545 );
buf ( n30547 , n29905 );
not ( n1464 , n30547 );
or ( n1465 , n1462 , n1464 );
buf ( n30550 , n499 );
not ( n1467 , n30550 );
buf ( n30552 , n30090 );
not ( n1469 , n30552 );
or ( n1470 , n1467 , n1469 );
buf ( n30555 , n30096 );
buf ( n30556 , n29901 );
nand ( n1473 , n30555 , n30556 );
buf ( n30558 , n1473 );
buf ( n30559 , n30558 );
nand ( n1476 , n1470 , n30559 );
buf ( n30561 , n1476 );
buf ( n30562 , n30561 );
buf ( n30563 , n29884 );
nand ( n1480 , n30562 , n30563 );
buf ( n30565 , n1480 );
buf ( n30566 , n30565 );
nand ( n1483 , n1465 , n30566 );
buf ( n30568 , n1483 );
buf ( n30569 , n30568 );
buf ( n30570 , n497 );
buf ( n30571 , n498 );
xnor ( n1488 , n30570 , n30571 );
buf ( n30573 , n1488 );
buf ( n30574 , n30573 );
not ( n1491 , n499 );
nand ( n1492 , n1491 , n498 );
not ( n1493 , n498 );
nand ( n1494 , n1493 , n499 );
nand ( n1495 , n1492 , n1494 );
buf ( n30580 , n1495 );
nor ( n1497 , n30574 , n30580 );
buf ( n30582 , n1497 );
buf ( n30583 , n30582 );
buf ( n1500 , n30583 );
buf ( n30585 , n1500 );
buf ( n30586 , n30585 );
not ( n1503 , n30586 );
buf ( n30588 , n497 );
not ( n1505 , n30588 );
buf ( n30590 , n29939 );
not ( n1507 , n30590 );
buf ( n30592 , n1507 );
buf ( n30593 , n30592 );
not ( n1510 , n30593 );
or ( n1511 , n1505 , n1510 );
buf ( n30596 , n29945 );
buf ( n30597 , n497 );
not ( n1514 , n30597 );
buf ( n30599 , n1514 );
buf ( n30600 , n30599 );
nand ( n1517 , n30596 , n30600 );
buf ( n30602 , n1517 );
buf ( n30603 , n30602 );
nand ( n1520 , n1511 , n30603 );
buf ( n30605 , n1520 );
buf ( n30606 , n30605 );
not ( n1523 , n30606 );
or ( n1524 , n1503 , n1523 );
buf ( n30609 , n497 );
not ( n1526 , n30609 );
buf ( n30611 , n29916 );
not ( n1528 , n30611 );
or ( n1529 , n1526 , n1528 );
buf ( n30614 , n784 );
buf ( n30615 , n30599 );
nand ( n1532 , n30614 , n30615 );
buf ( n30617 , n1532 );
buf ( n30618 , n30617 );
nand ( n1535 , n1529 , n30618 );
buf ( n30620 , n1535 );
buf ( n30621 , n30620 );
buf ( n30622 , n909 );
nand ( n1539 , n30621 , n30622 );
buf ( n30624 , n1539 );
buf ( n30625 , n30624 );
nand ( n1542 , n1524 , n30625 );
buf ( n30627 , n1542 );
buf ( n30628 , n30627 );
xor ( n1545 , n30569 , n30628 );
buf ( n30630 , n30078 );
not ( n1547 , n30630 );
buf ( n30632 , n30119 );
not ( n1549 , n30632 );
or ( n1550 , n1547 , n1549 );
buf ( n30635 , n1010 );
buf ( n30636 , n501 );
not ( n1553 , n30636 );
buf ( n30638 , n882 );
not ( n1555 , n30638 );
or ( n1556 , n1553 , n1555 );
buf ( n30641 , n30008 );
buf ( n30642 , n984 );
nand ( n1559 , n30641 , n30642 );
buf ( n30644 , n1559 );
buf ( n30645 , n30644 );
nand ( n1562 , n1556 , n30645 );
buf ( n30647 , n1562 );
buf ( n30648 , n30647 );
nand ( n1565 , n30635 , n30648 );
buf ( n30650 , n1565 );
buf ( n30651 , n30650 );
nand ( n1568 , n1550 , n30651 );
buf ( n30653 , n1568 );
buf ( n30654 , n30653 );
xor ( n30655 , n1545 , n30654 );
buf ( n30656 , n30655 );
buf ( n30657 , n30656 );
xor ( n1577 , n1460 , n30657 );
buf ( n30659 , n1577 );
not ( n1579 , n30659 );
xor ( n1580 , n29938 , n30026 );
and ( n1581 , n1580 , n30131 );
and ( n1582 , n29938 , n30026 );
or ( n1583 , n1581 , n1582 );
buf ( n30665 , n1583 );
not ( n1585 , n30665 );
nand ( n1586 , n1579 , n1585 );
nand ( n1587 , n30659 , n30665 );
nand ( n1588 , n1586 , n1587 );
not ( n1589 , n1588 );
and ( n1590 , n1391 , n1589 );
not ( n1591 , n1391 );
and ( n1592 , n1591 , n1588 );
nor ( n1593 , n1590 , n1592 );
nand ( n1594 , n1593 , n455 );
buf ( n30676 , n29615 );
not ( n1596 , n30676 );
buf ( n30678 , n29582 );
not ( n1598 , n30678 );
or ( n30680 , n1596 , n1598 );
buf ( n30681 , n513 );
buf ( n30682 , n503 );
xor ( n1605 , n30681 , n30682 );
buf ( n30684 , n1605 );
buf ( n30685 , n30684 );
buf ( n30686 , n504 );
nand ( n1609 , n30685 , n30686 );
buf ( n30688 , n1609 );
buf ( n30689 , n30688 );
nand ( n1612 , n30680 , n30689 );
buf ( n30691 , n1612 );
buf ( n30692 , n30691 );
buf ( n30693 , n520 );
buf ( n30694 , n498 );
or ( n1617 , n30693 , n30694 );
buf ( n30696 , n499 );
nand ( n1619 , n1617 , n30696 );
buf ( n30698 , n1619 );
buf ( n30699 , n30698 );
buf ( n30700 , n520 );
buf ( n30701 , n498 );
nand ( n1624 , n30700 , n30701 );
buf ( n30703 , n1624 );
buf ( n30704 , n30703 );
buf ( n30705 , n497 );
and ( n1628 , n30699 , n30704 , n30705 );
buf ( n30707 , n1628 );
buf ( n30708 , n30707 );
xor ( n1631 , n30692 , n30708 );
buf ( n30710 , n1631 );
buf ( n30711 , n30710 );
xor ( n1634 , n29609 , n29623 );
and ( n1635 , n1634 , n29661 );
and ( n1636 , n29609 , n29623 );
or ( n1637 , n1635 , n1636 );
buf ( n30716 , n1637 );
buf ( n30717 , n30716 );
xor ( n1640 , n30711 , n30717 );
buf ( n30719 , n29654 );
not ( n1642 , n30719 );
buf ( n30721 , n29640 );
not ( n1644 , n30721 );
or ( n1645 , n1642 , n1644 );
buf ( n30724 , n515 );
buf ( n30725 , n501 );
xor ( n1648 , n30724 , n30725 );
buf ( n30727 , n1648 );
buf ( n30728 , n30727 );
buf ( n30729 , n29649 );
nand ( n1652 , n30728 , n30729 );
buf ( n30731 , n1652 );
buf ( n30732 , n30731 );
nand ( n1655 , n1645 , n30732 );
buf ( n30734 , n1655 );
buf ( n30735 , n30734 );
buf ( n30736 , n29548 );
not ( n1659 , n30736 );
nand ( n1660 , n29528 , n29533 );
buf ( n30739 , n1660 );
not ( n1662 , n30739 );
buf ( n30741 , n1662 );
buf ( n30742 , n30741 );
not ( n1665 , n30742 );
or ( n30744 , n1659 , n1665 );
buf ( n30745 , n517 );
buf ( n30746 , n499 );
xnor ( n1669 , n30745 , n30746 );
buf ( n30748 , n1669 );
buf ( n30749 , n30748 );
not ( n1675 , n30749 );
buf ( n30751 , n29543 );
nand ( n1677 , n1675 , n30751 );
buf ( n30753 , n1677 );
buf ( n30754 , n30753 );
nand ( n1680 , n30744 , n30754 );
buf ( n30756 , n1680 );
buf ( n30757 , n30756 );
xor ( n1683 , n30735 , n30757 );
buf ( n30759 , n520 );
buf ( n30760 , n497 );
xor ( n1686 , n30759 , n30760 );
buf ( n30762 , n1686 );
buf ( n30763 , n30762 );
not ( n1689 , n30763 );
xnor ( n1690 , n497 , n498 );
nor ( n1691 , n1690 , n29602 );
buf ( n30767 , n1691 );
buf ( n1693 , n30767 );
buf ( n30769 , n1693 );
buf ( n30770 , n30769 );
not ( n1696 , n30770 );
or ( n1697 , n1689 , n1696 );
buf ( n1698 , n29604 );
buf ( n30774 , n1698 );
xor ( n1700 , n497 , n519 );
buf ( n30776 , n1700 );
nand ( n1702 , n30774 , n30776 );
buf ( n30778 , n1702 );
buf ( n30779 , n30778 );
nand ( n1705 , n1697 , n30779 );
buf ( n30781 , n1705 );
buf ( n30782 , n30781 );
xor ( n1708 , n1683 , n30782 );
buf ( n30784 , n1708 );
buf ( n30785 , n30784 );
xor ( n1711 , n1640 , n30785 );
buf ( n30787 , n1711 );
xor ( n1713 , n29555 , n29600 );
and ( n30789 , n1713 , n29664 );
and ( n1715 , n29555 , n29600 );
or ( n1716 , n30789 , n1715 );
buf ( n30792 , n1716 );
and ( n1718 , n30787 , n30792 );
not ( n1719 , n1718 );
nor ( n1720 , n30787 , n30792 );
not ( n1721 , n1720 );
nand ( n1722 , n1719 , n1721 );
not ( n1723 , n1722 );
not ( n1724 , n29717 );
not ( n1725 , n731 );
or ( n1726 , n1724 , n1725 );
nand ( n1727 , n1726 , n29719 );
not ( n1728 , n1727 );
or ( n1729 , n1723 , n1728 );
or ( n1730 , n1727 , n1722 );
nand ( n1731 , n1729 , n1730 );
nand ( n1732 , n1731 , n29519 );
nand ( n1733 , n1594 , n1732 );
not ( n1734 , n548 );
nand ( n1735 , n1733 , n1734 );
buf ( n30811 , n1735 );
nand ( n1740 , n30477 , n30811 );
buf ( n30813 , n1740 );
buf ( n30814 , n547 );
not ( n1743 , n30814 );
buf ( n30816 , n1743 );
not ( n1745 , n30816 );
not ( n30818 , n29519 );
not ( n1747 , n731 );
nor ( n1748 , n1720 , n29716 );
not ( n1749 , n1748 );
or ( n1750 , n1747 , n1749 );
and ( n1751 , n1721 , n29718 );
nor ( n30824 , n1751 , n1718 );
nand ( n1753 , n1750 , n30824 );
buf ( n30826 , n30684 );
not ( n1755 , n30826 );
buf ( n30828 , n29734 );
not ( n1757 , n30828 );
or ( n1758 , n1755 , n1757 );
buf ( n30831 , n512 );
buf ( n30832 , n503 );
xor ( n1761 , n30831 , n30832 );
buf ( n30834 , n1761 );
buf ( n30835 , n30834 );
buf ( n30836 , n504 );
nand ( n1765 , n30835 , n30836 );
buf ( n30838 , n1765 );
buf ( n30839 , n30838 );
nand ( n1768 , n1758 , n30839 );
buf ( n30841 , n1768 );
buf ( n30842 , n30841 );
buf ( n30843 , n496 );
buf ( n30844 , n497 );
xor ( n1773 , n30843 , n30844 );
buf ( n30846 , n1773 );
buf ( n30847 , n30846 );
buf ( n30848 , n520 );
and ( n1777 , n30847 , n30848 );
buf ( n30850 , n1777 );
buf ( n30851 , n30850 );
xor ( n1780 , n30842 , n30851 );
buf ( n30853 , n1700 );
not ( n1782 , n30853 );
buf ( n30855 , n30769 );
not ( n1784 , n30855 );
or ( n1785 , n1782 , n1784 );
not ( n1786 , n29603 );
buf ( n30859 , n1786 );
xor ( n1788 , n497 , n518 );
buf ( n30861 , n1788 );
nand ( n1790 , n30859 , n30861 );
buf ( n30863 , n1790 );
buf ( n30864 , n30863 );
nand ( n1793 , n1785 , n30864 );
buf ( n30866 , n1793 );
buf ( n30867 , n30866 );
xor ( n1796 , n1780 , n30867 );
buf ( n30869 , n1796 );
buf ( n30870 , n30869 );
xor ( n1799 , n30735 , n30757 );
and ( n1800 , n1799 , n30782 );
and ( n1801 , n30735 , n30757 );
or ( n1802 , n1800 , n1801 );
buf ( n30875 , n1802 );
buf ( n30876 , n30875 );
xor ( n1805 , n30870 , n30876 );
buf ( n30878 , n30727 );
not ( n1807 , n30878 );
buf ( n30880 , n29640 );
not ( n1809 , n30880 );
or ( n1810 , n1807 , n1809 );
buf ( n30883 , n29649 );
buf ( n30884 , n514 );
buf ( n30885 , n501 );
xor ( n1814 , n30884 , n30885 );
buf ( n30887 , n1814 );
buf ( n30888 , n30887 );
nand ( n30889 , n30883 , n30888 );
buf ( n30890 , n30889 );
buf ( n30891 , n30890 );
nand ( n1820 , n1810 , n30891 );
buf ( n30893 , n1820 );
buf ( n30894 , n30893 );
buf ( n30895 , n30691 );
buf ( n30896 , n30707 );
and ( n1825 , n30895 , n30896 );
buf ( n30898 , n1825 );
buf ( n30899 , n30898 );
xor ( n1828 , n30894 , n30899 );
buf ( n30901 , n516 );
buf ( n30902 , n499 );
xor ( n1831 , n30901 , n30902 );
buf ( n30904 , n1831 );
buf ( n30905 , n30904 );
not ( n1834 , n30905 );
buf ( n30907 , n29543 );
not ( n1836 , n30907 );
or ( n1837 , n1834 , n1836 );
buf ( n30910 , n29535 );
not ( n1839 , n30910 );
buf ( n30912 , n1839 );
buf ( n30913 , n30912 );
buf ( n30914 , n30748 );
or ( n1843 , n30913 , n30914 );
nand ( n1844 , n1837 , n1843 );
buf ( n30917 , n1844 );
buf ( n30918 , n30917 );
xor ( n1847 , n1828 , n30918 );
buf ( n30920 , n1847 );
buf ( n30921 , n30920 );
xor ( n1850 , n1805 , n30921 );
buf ( n30923 , n1850 );
xor ( n1852 , n30711 , n30717 );
and ( n1853 , n1852 , n30785 );
and ( n1854 , n30711 , n30717 );
or ( n1855 , n1853 , n1854 );
buf ( n30928 , n1855 );
nor ( n1857 , n30923 , n30928 );
not ( n1858 , n1857 );
nand ( n1859 , n30923 , n30928 );
nand ( n1860 , n1858 , n1859 );
xnor ( n1861 , n1753 , n1860 );
not ( n1862 , n1861 );
or ( n1863 , n30818 , n1862 );
nor ( n1864 , n30659 , n30665 );
nor ( n1865 , n1864 , n1091 );
not ( n1866 , n1865 );
not ( n1870 , n1286 );
or ( n30940 , n1866 , n1870 );
and ( n1872 , n1586 , n1093 );
not ( n1873 , n1587 );
nor ( n1874 , n1872 , n1873 );
nand ( n1875 , n30940 , n1874 );
not ( n1876 , n1875 );
buf ( n30946 , n504 );
not ( n1878 , n30946 );
buf ( n30948 , n503 );
not ( n1880 , n30948 );
and ( n1881 , n456 , n464 );
nor ( n1882 , n29498 , n456 );
nor ( n1883 , n1881 , n1882 );
buf ( n30953 , n1883 );
not ( n1885 , n30953 );
or ( n1886 , n1880 , n1885 );
buf ( n30956 , n29501 );
buf ( n30957 , n29987 );
nand ( n1889 , n30956 , n30957 );
buf ( n30959 , n1889 );
buf ( n30960 , n30959 );
nand ( n1892 , n1886 , n30960 );
buf ( n30962 , n1892 );
buf ( n30963 , n30962 );
not ( n1895 , n30963 );
or ( n1896 , n1878 , n1895 );
buf ( n30966 , n30506 );
buf ( n30967 , n29969 );
nand ( n1899 , n30966 , n30967 );
buf ( n30969 , n1899 );
buf ( n30970 , n30969 );
nand ( n1905 , n1896 , n30970 );
buf ( n30972 , n1905 );
buf ( n30973 , n29957 );
not ( n1908 , n496 );
not ( n1909 , n497 );
not ( n1910 , n1909 );
or ( n1911 , n1908 , n1910 );
not ( n1912 , n496 );
nand ( n1913 , n1912 , n497 );
nand ( n1914 , n1911 , n1913 );
buf ( n30981 , n1914 );
nand ( n1916 , n30973 , n30981 );
buf ( n30983 , n1916 );
and ( n1918 , n30972 , n30983 );
not ( n1919 , n30972 );
buf ( n30986 , n30983 );
not ( n1921 , n30986 );
buf ( n30988 , n1921 );
and ( n1923 , n1919 , n30988 );
or ( n1924 , n1918 , n1923 );
buf ( n30991 , n909 );
not ( n1926 , n30991 );
buf ( n30993 , n497 );
not ( n1928 , n30993 );
buf ( n30995 , n29897 );
not ( n30996 , n30995 );
or ( n1931 , n1928 , n30996 );
buf ( n30998 , n29514 );
buf ( n30999 , n30599 );
nand ( n1934 , n30998 , n30999 );
buf ( n31001 , n1934 );
buf ( n31002 , n31001 );
nand ( n1937 , n1931 , n31002 );
buf ( n31004 , n1937 );
buf ( n31005 , n31004 );
not ( n1940 , n31005 );
or ( n1941 , n1926 , n1940 );
buf ( n31008 , n30620 );
buf ( n31009 , n30585 );
nand ( n1944 , n31008 , n31009 );
buf ( n31011 , n1944 );
buf ( n31012 , n31011 );
nand ( n1947 , n1941 , n31012 );
buf ( n31014 , n1947 );
buf ( n1949 , n31014 );
and ( n1950 , n1924 , n1949 );
not ( n1951 , n1924 );
buf ( n31018 , n31014 );
not ( n1953 , n31018 );
buf ( n31020 , n1953 );
and ( n1955 , n1951 , n31020 );
nor ( n1956 , n1950 , n1955 );
buf ( n31023 , n1956 );
xor ( n1958 , n30569 , n30628 );
and ( n1959 , n1958 , n30654 );
and ( n1960 , n30569 , n30628 );
or ( n1961 , n1959 , n1960 );
buf ( n31028 , n1961 );
buf ( n31029 , n31028 );
xor ( n1964 , n31023 , n31029 );
buf ( n31031 , n799 );
not ( n1966 , n31031 );
buf ( n31033 , n30561 );
not ( n1968 , n31033 );
or ( n1969 , n1966 , n1968 );
not ( n1970 , n499 );
or ( n1971 , n29507 , n1970 );
nand ( n1972 , n29507 , n29901 );
nand ( n1973 , n1971 , n1972 );
buf ( n31040 , n1973 );
buf ( n31041 , n745 );
nand ( n1976 , n31040 , n31041 );
buf ( n31043 , n1976 );
buf ( n31044 , n31043 );
nand ( n1979 , n1969 , n31044 );
buf ( n31046 , n1979 );
buf ( n31047 , n31046 );
buf ( n31048 , n1010 );
not ( n1983 , n31048 );
buf ( n31050 , n501 );
not ( n1985 , n31050 );
buf ( n31052 , n929 );
not ( n1987 , n31052 );
or ( n1991 , n1985 , n1987 );
buf ( n31055 , n933 );
buf ( n31056 , n984 );
nand ( n1994 , n31055 , n31056 );
buf ( n31058 , n1994 );
buf ( n31059 , n31058 );
nand ( n1997 , n1991 , n31059 );
buf ( n31061 , n1997 );
buf ( n31062 , n31061 );
not ( n2000 , n31062 );
or ( n2001 , n1983 , n2000 );
buf ( n31065 , n30647 );
buf ( n31066 , n30078 );
nand ( n2004 , n31065 , n31066 );
buf ( n31068 , n2004 );
buf ( n31069 , n31068 );
nand ( n2007 , n2001 , n31069 );
buf ( n31071 , n2007 );
buf ( n31072 , n31071 );
xor ( n2010 , n31047 , n31072 );
buf ( n31074 , n30513 );
buf ( n31075 , n30533 );
and ( n2013 , n31074 , n31075 );
buf ( n31077 , n2013 );
buf ( n31078 , n31077 );
xor ( n2016 , n2010 , n31078 );
buf ( n31080 , n2016 );
buf ( n31081 , n31080 );
xor ( n2019 , n1964 , n31081 );
buf ( n31083 , n2019 );
xor ( n2021 , n30537 , n30543 );
and ( n2022 , n2021 , n30657 );
and ( n2023 , n30537 , n30543 );
or ( n2024 , n2022 , n2023 );
buf ( n31088 , n2024 );
nand ( n2026 , n31083 , n31088 );
not ( n2027 , n2026 );
nor ( n2028 , n31083 , n31088 );
buf ( n2029 , n2028 );
nor ( n2030 , n2027 , n2029 );
not ( n2031 , n2030 );
and ( n2032 , n1876 , n2031 );
not ( n2033 , n1876 );
and ( n2034 , n2033 , n2030 );
nor ( n2035 , n2032 , n2034 );
nand ( n2036 , n2035 , n455 );
nand ( n2037 , n1863 , n2036 );
buf ( n31101 , n2037 );
not ( n2039 , n31101 );
buf ( n31103 , n2039 );
not ( n2041 , n31103 );
or ( n2042 , n1745 , n2041 );
buf ( n31106 , n2037 );
buf ( n31107 , n547 );
nand ( n2045 , n31106 , n31107 );
buf ( n31109 , n2045 );
nand ( n2047 , n2042 , n31109 );
not ( n2048 , n1733 );
not ( n2049 , n2048 );
nor ( n2050 , n2047 , n2049 );
not ( n2051 , n2050 );
nand ( n2052 , n2049 , n2047 );
nand ( n2053 , n2048 , n548 );
nand ( n2054 , n30813 , n2051 , n2052 , n2053 );
not ( n2055 , n2054 );
not ( n2056 , n2052 );
not ( n2057 , n2051 );
or ( n2058 , n2056 , n2057 );
nand ( n31122 , n2053 , n30813 );
nand ( n2063 , n2058 , n31122 );
not ( n2064 , n2063 );
or ( n2065 , n2055 , n2064 );
nand ( n2066 , n2065 , n454 );
buf ( n31127 , n469 );
not ( n2068 , n31127 );
buf ( n31129 , n533 );
buf ( n31130 , n552 );
nand ( n2071 , n31129 , n31130 );
buf ( n31132 , n2071 );
buf ( n31133 , n31132 );
nand ( n2074 , n2068 , n31133 );
buf ( n31135 , n2074 );
buf ( n31136 , n31135 );
buf ( n31137 , n534 );
buf ( n31138 , n550 );
and ( n2079 , n31137 , n31138 );
buf ( n31140 , n2079 );
buf ( n31141 , n31140 );
buf ( n31142 , n535 );
buf ( n31143 , n549 );
and ( n2084 , n31142 , n31143 );
buf ( n31145 , n2084 );
buf ( n31146 , n31145 );
xor ( n2087 , n31141 , n31146 );
buf ( n31148 , n533 );
buf ( n31149 , n551 );
and ( n2090 , n31148 , n31149 );
buf ( n31151 , n2090 );
buf ( n31152 , n31151 );
xor ( n2093 , n2087 , n31152 );
buf ( n31154 , n2093 );
buf ( n31155 , n31154 );
xor ( n31156 , n31136 , n31155 );
buf ( n31157 , n536 );
buf ( n31158 , n548 );
and ( n2099 , n31157 , n31158 );
buf ( n31160 , n2099 );
buf ( n31161 , n31160 );
buf ( n31162 , n468 );
buf ( n31163 , n532 );
buf ( n31164 , n552 );
and ( n2105 , n31163 , n31164 );
buf ( n31166 , n2105 );
buf ( n31167 , n31166 );
xor ( n2108 , n31162 , n31167 );
buf ( n31169 , n2108 );
buf ( n31170 , n31169 );
xor ( n2111 , n31161 , n31170 );
buf ( n31172 , n535 );
buf ( n31173 , n550 );
and ( n2114 , n31172 , n31173 );
buf ( n31175 , n2114 );
buf ( n31176 , n31175 );
buf ( n31177 , n536 );
buf ( n31178 , n549 );
and ( n2119 , n31177 , n31178 );
buf ( n31180 , n2119 );
buf ( n31181 , n31180 );
xor ( n2122 , n31176 , n31181 );
buf ( n31183 , n534 );
buf ( n31184 , n551 );
and ( n2125 , n31183 , n31184 );
buf ( n31186 , n2125 );
buf ( n31187 , n31186 );
and ( n2128 , n2122 , n31187 );
and ( n2129 , n31176 , n31181 );
or ( n2130 , n2128 , n2129 );
buf ( n31191 , n2130 );
buf ( n31192 , n31191 );
xor ( n2133 , n2111 , n31192 );
buf ( n31194 , n2133 );
buf ( n31195 , n31194 );
xor ( n2136 , n31156 , n31195 );
buf ( n31197 , n2136 );
buf ( n31198 , n31197 );
buf ( n31199 , n470 );
buf ( n31200 , n534 );
buf ( n31201 , n552 );
and ( n2142 , n31200 , n31201 );
buf ( n31203 , n2142 );
buf ( n31204 , n31203 );
and ( n2145 , n31199 , n31204 );
buf ( n31206 , n2145 );
buf ( n31207 , n31206 );
buf ( n31208 , n469 );
not ( n2149 , n31208 );
buf ( n31210 , n31132 );
not ( n2151 , n31210 );
buf ( n31212 , n2151 );
buf ( n31213 , n31212 );
not ( n2154 , n31213 );
or ( n2155 , n2149 , n2154 );
buf ( n31216 , n31135 );
nand ( n2157 , n2155 , n31216 );
buf ( n31218 , n2157 );
buf ( n31219 , n31218 );
xor ( n2160 , n31207 , n31219 );
xor ( n2161 , n31176 , n31181 );
xor ( n2162 , n2161 , n31187 );
buf ( n31223 , n2162 );
buf ( n31224 , n31223 );
and ( n2165 , n2160 , n31224 );
and ( n2166 , n31207 , n31219 );
or ( n2167 , n2165 , n2166 );
buf ( n31228 , n2167 );
buf ( n31229 , n31228 );
nor ( n2170 , n31198 , n31229 );
buf ( n31231 , n2170 );
buf ( n31232 , n31231 );
xor ( n2173 , n31207 , n31219 );
xor ( n2174 , n2173 , n31224 );
buf ( n31235 , n2174 );
buf ( n31236 , n31235 );
buf ( n31237 , n536 );
buf ( n31238 , n550 );
and ( n2179 , n31237 , n31238 );
buf ( n31240 , n2179 );
buf ( n31241 , n31240 );
buf ( n31242 , n535 );
buf ( n31243 , n551 );
and ( n2184 , n31242 , n31243 );
buf ( n31245 , n2184 );
buf ( n31246 , n31245 );
xor ( n2187 , n31241 , n31246 );
xor ( n2188 , n31199 , n31204 );
buf ( n31249 , n2188 );
buf ( n31250 , n31249 );
and ( n2191 , n2187 , n31250 );
and ( n2192 , n31241 , n31246 );
or ( n2193 , n2191 , n2192 );
buf ( n31254 , n2193 );
buf ( n31255 , n31254 );
or ( n2196 , n31236 , n31255 );
buf ( n31257 , n2196 );
buf ( n31258 , n31257 );
buf ( n31259 , n471 );
buf ( n31260 , n536 );
buf ( n31261 , n551 );
and ( n2202 , n31260 , n31261 );
buf ( n31263 , n2202 );
buf ( n31264 , n31263 );
and ( n2208 , n31259 , n31264 );
buf ( n31266 , n2208 );
buf ( n31267 , n31266 );
buf ( n31268 , n535 );
buf ( n31269 , n552 );
and ( n2213 , n31268 , n31269 );
buf ( n31271 , n2213 );
buf ( n31272 , n31271 );
buf ( n31273 , n472 );
not ( n2217 , n31273 );
buf ( n31275 , n536 );
buf ( n31276 , n552 );
nand ( n2220 , n31275 , n31276 );
buf ( n31278 , n2220 );
buf ( n31279 , n31278 );
nor ( n2223 , n2217 , n31279 );
buf ( n31281 , n2223 );
buf ( n31282 , n31281 );
xor ( n2226 , n31272 , n31282 );
xor ( n2227 , n31259 , n31264 );
buf ( n31285 , n2227 );
buf ( n31286 , n31285 );
and ( n2230 , n2226 , n31286 );
and ( n2231 , n31272 , n31282 );
or ( n2232 , n2230 , n2231 );
buf ( n31290 , n2232 );
buf ( n31291 , n31290 );
xor ( n2235 , n31267 , n31291 );
xor ( n2236 , n31241 , n31246 );
xor ( n2237 , n2236 , n31250 );
buf ( n31295 , n2237 );
buf ( n31296 , n31295 );
and ( n2240 , n2235 , n31296 );
and ( n2241 , n31267 , n31291 );
or ( n2242 , n2240 , n2241 );
buf ( n31300 , n2242 );
buf ( n31301 , n31300 );
and ( n2248 , n31258 , n31301 );
buf ( n31303 , n31235 );
buf ( n31304 , n31254 );
and ( n2251 , n31303 , n31304 );
buf ( n31306 , n2251 );
buf ( n31307 , n31306 );
nor ( n2254 , n2248 , n31307 );
buf ( n31309 , n2254 );
buf ( n31310 , n31309 );
or ( n2257 , n31232 , n31310 );
buf ( n31312 , n31197 );
buf ( n31313 , n31228 );
nand ( n2260 , n31312 , n31313 );
buf ( n31315 , n2260 );
buf ( n31316 , n31315 );
nand ( n2263 , n2257 , n31316 );
buf ( n31318 , n2263 );
buf ( n31319 , n31318 );
not ( n2266 , n31319 );
buf ( n31321 , n535 );
buf ( n31322 , n548 );
and ( n2269 , n31321 , n31322 );
buf ( n31324 , n2269 );
buf ( n31325 , n31324 );
buf ( n31326 , n536 );
buf ( n31327 , n547 );
and ( n2274 , n31326 , n31327 );
buf ( n31329 , n2274 );
buf ( n31330 , n31329 );
xor ( n2277 , n31325 , n31330 );
and ( n2278 , n31162 , n31167 );
buf ( n31333 , n2278 );
buf ( n31334 , n31333 );
xor ( n2281 , n2277 , n31334 );
buf ( n31336 , n2281 );
buf ( n31337 , n31336 );
xor ( n2284 , n31161 , n31170 );
and ( n2285 , n2284 , n31192 );
and ( n2286 , n31161 , n31170 );
or ( n2287 , n2285 , n2286 );
buf ( n31342 , n2287 );
buf ( n31343 , n31342 );
xor ( n2290 , n31337 , n31343 );
buf ( n31345 , n467 );
buf ( n31346 , n531 );
buf ( n31347 , n552 );
and ( n2294 , n31346 , n31347 );
buf ( n31349 , n2294 );
buf ( n31350 , n31349 );
xor ( n2297 , n31345 , n31350 );
buf ( n31352 , n2297 );
buf ( n31353 , n31352 );
xor ( n2300 , n31141 , n31146 );
and ( n2301 , n2300 , n31152 );
and ( n2302 , n31141 , n31146 );
or ( n2303 , n2301 , n2302 );
buf ( n31358 , n2303 );
buf ( n31359 , n31358 );
xor ( n2306 , n31353 , n31359 );
buf ( n31361 , n533 );
buf ( n31362 , n550 );
and ( n2309 , n31361 , n31362 );
buf ( n31364 , n2309 );
buf ( n31365 , n31364 );
buf ( n31366 , n534 );
buf ( n31367 , n549 );
and ( n2314 , n31366 , n31367 );
buf ( n31369 , n2314 );
buf ( n31370 , n31369 );
xor ( n2317 , n31365 , n31370 );
buf ( n31372 , n532 );
buf ( n31373 , n551 );
and ( n2320 , n31372 , n31373 );
buf ( n31375 , n2320 );
buf ( n31376 , n31375 );
xor ( n2323 , n2317 , n31376 );
buf ( n31378 , n2323 );
buf ( n31379 , n31378 );
xor ( n2326 , n2306 , n31379 );
buf ( n31381 , n2326 );
buf ( n31382 , n31381 );
xor ( n2329 , n2290 , n31382 );
buf ( n31384 , n2329 );
buf ( n31385 , n31384 );
xor ( n2332 , n31136 , n31155 );
and ( n2333 , n2332 , n31195 );
and ( n2334 , n31136 , n31155 );
or ( n2335 , n2333 , n2334 );
buf ( n31390 , n2335 );
buf ( n31391 , n31390 );
or ( n2338 , n31385 , n31391 );
buf ( n31393 , n2338 );
buf ( n31394 , n31393 );
buf ( n31395 , n31390 );
buf ( n31396 , n31384 );
nand ( n2343 , n31395 , n31396 );
buf ( n31398 , n2343 );
buf ( n31399 , n31398 );
nand ( n2346 , n31394 , n31399 );
buf ( n31401 , n2346 );
buf ( n31402 , n31401 );
not ( n2349 , n31402 );
or ( n2350 , n2266 , n2349 );
buf ( n31405 , n31401 );
buf ( n31406 , n31318 );
or ( n2353 , n31405 , n31406 );
nand ( n2354 , n2350 , n2353 );
buf ( n31409 , n2354 );
not ( n2356 , n454 );
nand ( n2357 , n31409 , n2356 );
nand ( n2358 , n2066 , n2357 );
and ( n2359 , n31345 , n31350 );
buf ( n31414 , n2359 );
buf ( n31415 , n31414 );
buf ( n31416 , n466 );
buf ( n31417 , n530 );
buf ( n31418 , n552 );
and ( n2365 , n31417 , n31418 );
buf ( n31420 , n2365 );
buf ( n31421 , n31420 );
xor ( n2368 , n31416 , n31421 );
buf ( n31423 , n2368 );
buf ( n31424 , n31423 );
xor ( n2371 , n31415 , n31424 );
xor ( n2372 , n31365 , n31370 );
and ( n2373 , n2372 , n31376 );
and ( n2374 , n31365 , n31370 );
or ( n2375 , n2373 , n2374 );
buf ( n31430 , n2375 );
buf ( n31431 , n31430 );
xor ( n2378 , n2371 , n31431 );
buf ( n31433 , n2378 );
buf ( n31434 , n31433 );
xor ( n2381 , n31353 , n31359 );
and ( n2382 , n2381 , n31379 );
and ( n2383 , n31353 , n31359 );
or ( n2384 , n2382 , n2383 );
buf ( n31439 , n2384 );
buf ( n31440 , n31439 );
xor ( n2387 , n31434 , n31440 );
buf ( n31442 , n531 );
buf ( n31443 , n551 );
and ( n2390 , n31442 , n31443 );
buf ( n31445 , n2390 );
buf ( n31446 , n31445 );
buf ( n31447 , n534 );
buf ( n31448 , n548 );
and ( n2395 , n31447 , n31448 );
buf ( n31450 , n2395 );
buf ( n31451 , n31450 );
xor ( n2398 , n31446 , n31451 );
buf ( n31453 , n535 );
buf ( n31454 , n547 );
and ( n2401 , n31453 , n31454 );
buf ( n31456 , n2401 );
buf ( n31457 , n31456 );
xor ( n2404 , n2398 , n31457 );
buf ( n31459 , n2404 );
buf ( n31460 , n31459 );
buf ( n31461 , n532 );
buf ( n31462 , n550 );
and ( n2412 , n31461 , n31462 );
buf ( n31464 , n2412 );
buf ( n31465 , n31464 );
buf ( n31466 , n536 );
buf ( n31467 , n546 );
and ( n2417 , n31466 , n31467 );
buf ( n31469 , n2417 );
buf ( n31470 , n31469 );
xor ( n2420 , n31465 , n31470 );
buf ( n31472 , n533 );
buf ( n31473 , n549 );
and ( n2423 , n31472 , n31473 );
buf ( n31475 , n2423 );
buf ( n31476 , n31475 );
xor ( n2426 , n2420 , n31476 );
buf ( n31478 , n2426 );
buf ( n31479 , n31478 );
xor ( n2429 , n31460 , n31479 );
xor ( n2430 , n31325 , n31330 );
and ( n2431 , n2430 , n31334 );
and ( n2432 , n31325 , n31330 );
or ( n2433 , n2431 , n2432 );
buf ( n31485 , n2433 );
buf ( n31486 , n31485 );
xor ( n2436 , n2429 , n31486 );
buf ( n31488 , n2436 );
buf ( n31489 , n31488 );
xor ( n2439 , n2387 , n31489 );
buf ( n31491 , n2439 );
buf ( n31492 , n31491 );
xor ( n2442 , n31337 , n31343 );
and ( n2443 , n2442 , n31382 );
and ( n2444 , n31337 , n31343 );
or ( n2445 , n2443 , n2444 );
buf ( n31497 , n2445 );
buf ( n31498 , n31497 );
or ( n2448 , n31492 , n31498 );
buf ( n31500 , n2448 );
buf ( n31501 , n31500 );
buf ( n31502 , n31491 );
buf ( n31503 , n31497 );
nand ( n2453 , n31502 , n31503 );
buf ( n31505 , n2453 );
buf ( n31506 , n31505 );
nand ( n2456 , n31501 , n31506 );
buf ( n31508 , n2456 );
buf ( n31509 , n31508 );
not ( n2459 , n31509 );
buf ( n31511 , n31393 );
not ( n2461 , n31511 );
buf ( n31513 , n31318 );
not ( n2463 , n31513 );
or ( n2464 , n2461 , n2463 );
buf ( n31516 , n31398 );
nand ( n2466 , n2464 , n31516 );
buf ( n31518 , n2466 );
buf ( n31519 , n31518 );
not ( n2469 , n31519 );
or ( n2470 , n2459 , n2469 );
buf ( n31522 , n31518 );
buf ( n31523 , n31508 );
or ( n2473 , n31522 , n31523 );
nand ( n2474 , n2470 , n2473 );
buf ( n31526 , n2474 );
nand ( n2476 , n31526 , n2356 );
xor ( n2477 , n31446 , n31451 );
and ( n2478 , n2477 , n31457 );
and ( n2479 , n31446 , n31451 );
or ( n2480 , n2478 , n2479 );
buf ( n31532 , n2480 );
buf ( n31533 , n31532 );
xor ( n2483 , n31465 , n31470 );
and ( n2484 , n2483 , n31476 );
and ( n2485 , n31465 , n31470 );
or ( n2486 , n2484 , n2485 );
buf ( n31538 , n2486 );
buf ( n31539 , n31538 );
xor ( n2489 , n31533 , n31539 );
buf ( n31541 , n532 );
buf ( n31542 , n549 );
and ( n2492 , n31541 , n31542 );
buf ( n31544 , n2492 );
buf ( n31545 , n31544 );
buf ( n31546 , n530 );
buf ( n31547 , n551 );
and ( n2497 , n31546 , n31547 );
buf ( n31549 , n2497 );
buf ( n31550 , n31549 );
xor ( n2500 , n31545 , n31550 );
buf ( n31552 , n533 );
buf ( n31553 , n548 );
and ( n2503 , n31552 , n31553 );
buf ( n31555 , n2503 );
buf ( n31556 , n31555 );
xor ( n2506 , n2500 , n31556 );
buf ( n31558 , n2506 );
buf ( n31559 , n31558 );
xor ( n2509 , n2489 , n31559 );
buf ( n31561 , n2509 );
buf ( n31562 , n31561 );
xor ( n2512 , n31460 , n31479 );
and ( n2513 , n2512 , n31486 );
and ( n2514 , n31460 , n31479 );
or ( n2515 , n2513 , n2514 );
buf ( n31567 , n2515 );
buf ( n31568 , n31567 );
xor ( n2518 , n31562 , n31568 );
buf ( n31570 , n531 );
buf ( n31571 , n550 );
and ( n2521 , n31570 , n31571 );
buf ( n31573 , n2521 );
buf ( n31574 , n31573 );
buf ( n31575 , n535 );
buf ( n31576 , n546 );
and ( n2526 , n31575 , n31576 );
buf ( n31578 , n2526 );
buf ( n31579 , n31578 );
xor ( n2529 , n31574 , n31579 );
buf ( n31581 , n536 );
buf ( n31582 , n545 );
and ( n2532 , n31581 , n31582 );
buf ( n31584 , n2532 );
buf ( n31585 , n31584 );
xor ( n2535 , n2529 , n31585 );
buf ( n31587 , n2535 );
buf ( n31588 , n31587 );
xor ( n2538 , n31415 , n31424 );
and ( n2539 , n2538 , n31431 );
and ( n2540 , n31415 , n31424 );
or ( n2541 , n2539 , n2540 );
buf ( n31593 , n2541 );
buf ( n31594 , n31593 );
xor ( n2544 , n31588 , n31594 );
buf ( n31596 , n534 );
buf ( n31597 , n547 );
and ( n2547 , n31596 , n31597 );
buf ( n31599 , n2547 );
buf ( n31600 , n31599 );
buf ( n31601 , n465 );
buf ( n31602 , n529 );
buf ( n31603 , n552 );
and ( n2553 , n31602 , n31603 );
buf ( n31605 , n2553 );
buf ( n31606 , n31605 );
xor ( n2556 , n31601 , n31606 );
buf ( n31608 , n2556 );
buf ( n31609 , n31608 );
xor ( n2559 , n31600 , n31609 );
and ( n2560 , n31416 , n31421 );
buf ( n31612 , n2560 );
buf ( n31613 , n31612 );
xor ( n2563 , n2559 , n31613 );
buf ( n31615 , n2563 );
buf ( n31616 , n31615 );
xor ( n2566 , n2544 , n31616 );
buf ( n31618 , n2566 );
buf ( n31619 , n31618 );
xor ( n31620 , n2518 , n31619 );
buf ( n31621 , n31620 );
buf ( n31622 , n31621 );
xor ( n2575 , n31434 , n31440 );
and ( n2576 , n2575 , n31489 );
and ( n2577 , n31434 , n31440 );
or ( n2578 , n2576 , n2577 );
buf ( n31627 , n2578 );
buf ( n31628 , n31627 );
or ( n2581 , n31622 , n31628 );
buf ( n31630 , n2581 );
buf ( n31631 , n31630 );
buf ( n31632 , n31621 );
buf ( n31633 , n31627 );
nand ( n2586 , n31632 , n31633 );
buf ( n31635 , n2586 );
buf ( n31636 , n31635 );
nand ( n2589 , n31631 , n31636 );
buf ( n31638 , n2589 );
buf ( n31639 , n31638 );
not ( n2592 , n31639 );
buf ( n31641 , n31500 );
not ( n2594 , n31641 );
buf ( n31643 , n31393 );
not ( n2596 , n31643 );
buf ( n31645 , n31318 );
not ( n2598 , n31645 );
or ( n2599 , n2596 , n2598 );
buf ( n31648 , n31398 );
nand ( n2601 , n2599 , n31648 );
buf ( n31650 , n2601 );
buf ( n31651 , n31650 );
not ( n2604 , n31651 );
or ( n2605 , n2594 , n2604 );
buf ( n31654 , n31505 );
nand ( n2607 , n2605 , n31654 );
buf ( n31656 , n2607 );
buf ( n31657 , n31656 );
not ( n2610 , n31657 );
or ( n2611 , n2592 , n2610 );
buf ( n31660 , n31656 );
buf ( n31661 , n31638 );
or ( n2614 , n31660 , n31661 );
nand ( n2615 , n2611 , n2614 );
buf ( n31664 , n2615 );
nand ( n2617 , n31664 , n2356 );
not ( n2618 , n454 );
and ( n2619 , n456 , n2618 );
not ( n2620 , n456 );
and ( n2621 , n2620 , n454 );
nor ( n2622 , n2619 , n2621 );
and ( n2623 , n455 , n2622 );
not ( n2624 , n455 );
not ( n2625 , n2622 );
and ( n2626 , n2624 , n2625 );
or ( n2627 , n2623 , n2626 );
not ( n2628 , n2627 );
not ( n2629 , n2628 );
not ( n2630 , n2629 );
buf ( n31679 , n29931 );
not ( n2632 , n31679 );
not ( n2633 , n1402 );
and ( n2634 , n2633 , n29901 );
not ( n2635 , n2633 );
and ( n2636 , n2635 , n499 );
or ( n2637 , n2634 , n2636 );
buf ( n31686 , n2637 );
not ( n2639 , n31686 );
or ( n2640 , n2632 , n2639 );
buf ( n31689 , n499 );
not ( n2642 , n31689 );
buf ( n31691 , n29501 );
not ( n2644 , n31691 );
buf ( n31693 , n2644 );
buf ( n31694 , n31693 );
not ( n2647 , n31694 );
or ( n2648 , n2642 , n2647 );
buf ( n31697 , n29501 );
buf ( n31698 , n29901 );
nand ( n31699 , n31697 , n31698 );
buf ( n31700 , n31699 );
buf ( n31701 , n31700 );
nand ( n2654 , n2648 , n31701 );
buf ( n31703 , n2654 );
buf ( n31704 , n31703 );
buf ( n31705 , n29884 );
nand ( n2658 , n31704 , n31705 );
buf ( n31707 , n2658 );
buf ( n31708 , n31707 );
nand ( n2661 , n2640 , n31708 );
buf ( n31710 , n2661 );
buf ( n31711 , n31710 );
buf ( n31712 , n1010 );
not ( n2665 , n31712 );
buf ( n31714 , n501 );
not ( n2667 , n31714 );
and ( n2668 , n456 , n463 );
not ( n2669 , n456 );
and ( n2670 , n2669 , n479 );
nor ( n2671 , n2668 , n2670 );
buf ( n31720 , n2671 );
not ( n2673 , n31720 );
or ( n2674 , n2667 , n2673 );
and ( n2675 , n456 , n463 );
not ( n2676 , n456 );
and ( n2677 , n2676 , n479 );
nor ( n2678 , n2675 , n2677 );
not ( n2679 , n2678 );
buf ( n31728 , n2679 );
buf ( n31729 , n984 );
nand ( n2682 , n31728 , n31729 );
buf ( n31731 , n2682 );
buf ( n31732 , n31731 );
nand ( n2685 , n2674 , n31732 );
buf ( n31734 , n2685 );
buf ( n31735 , n31734 );
not ( n2688 , n31735 );
or ( n2689 , n2665 , n2688 );
or ( n2690 , n743 , n29501 );
nand ( n2691 , n29501 , n984 );
nand ( n2692 , n2690 , n2691 );
buf ( n31741 , n2692 );
buf ( n31742 , n30078 );
nand ( n2695 , n31741 , n31742 );
buf ( n31744 , n2695 );
buf ( n31745 , n31744 );
nand ( n2698 , n2689 , n31745 );
buf ( n31747 , n2698 );
not ( n2700 , n31747 );
buf ( n31749 , n30141 );
buf ( n31750 , n494 );
and ( n2703 , n31749 , n31750 );
not ( n2704 , n493 );
buf ( n31753 , n2704 );
nor ( n2706 , n2703 , n31753 );
buf ( n31755 , n2706 );
not ( n2708 , n494 );
buf ( n31757 , n2708 );
not ( n2710 , n31757 );
buf ( n31759 , n29939 );
not ( n2712 , n31759 );
buf ( n31761 , n2712 );
buf ( n31762 , n31761 );
not ( n2715 , n31762 );
or ( n2716 , n2710 , n2715 );
buf ( n31765 , n495 );
nand ( n2718 , n2716 , n31765 );
buf ( n31767 , n2718 );
nand ( n2720 , n31755 , n31767 );
nor ( n2721 , n2700 , n2720 );
buf ( n31770 , n2721 );
xor ( n2723 , n31711 , n31770 );
not ( n2724 , n1914 );
not ( n2725 , n2724 );
buf ( n31774 , n2725 );
not ( n2727 , n31774 );
buf ( n31776 , n495 );
not ( n2729 , n31776 );
buf ( n31778 , n30090 );
not ( n2731 , n31778 );
or ( n2732 , n2729 , n2731 );
buf ( n31781 , n973 );
buf ( n31782 , n495 );
not ( n2738 , n31782 );
buf ( n31784 , n2738 );
buf ( n31785 , n31784 );
nand ( n2741 , n31781 , n31785 );
buf ( n31787 , n2741 );
buf ( n31788 , n31787 );
nand ( n2744 , n2732 , n31788 );
buf ( n31790 , n2744 );
buf ( n31791 , n31790 );
not ( n2747 , n31791 );
or ( n2748 , n2727 , n2747 );
not ( n2749 , n31784 );
not ( n2750 , n29513 );
or ( n2751 , n2749 , n2750 );
not ( n2752 , n495 );
or ( n2753 , n29513 , n2752 );
nand ( n2754 , n2751 , n2753 );
buf ( n31800 , n2754 );
xor ( n2756 , n496 , n495 );
buf ( n31802 , n2756 );
buf ( n31803 , n496 );
buf ( n31804 , n497 );
xnor ( n2760 , n31803 , n31804 );
buf ( n31806 , n2760 );
buf ( n31807 , n31806 );
nand ( n2763 , n31802 , n31807 );
buf ( n31809 , n2763 );
buf ( n31810 , n31809 );
not ( n2766 , n31810 );
buf ( n31812 , n2766 );
buf ( n31813 , n31812 );
nand ( n2769 , n31800 , n31813 );
buf ( n31815 , n2769 );
buf ( n31816 , n31815 );
nand ( n2772 , n2748 , n31816 );
buf ( n31818 , n2772 );
buf ( n31819 , n31818 );
buf ( n31820 , n504 );
not ( n2776 , n31820 );
buf ( n31822 , n503 );
not ( n2778 , n31822 );
buf ( n31824 , n29493 );
buf ( n2780 , n31824 );
buf ( n31826 , n2780 );
buf ( n31827 , n31826 );
not ( n2783 , n31827 );
buf ( n31829 , n2783 );
buf ( n31830 , n31829 );
not ( n2786 , n31830 );
or ( n2787 , n2778 , n2786 );
buf ( n31833 , n31826 );
buf ( n31834 , n29987 );
nand ( n2790 , n31833 , n31834 );
buf ( n31836 , n2790 );
buf ( n31837 , n31836 );
nand ( n2793 , n2787 , n31837 );
buf ( n31839 , n2793 );
buf ( n31840 , n31839 );
not ( n2796 , n31840 );
or ( n2797 , n2776 , n2796 );
not ( n2798 , n503 );
not ( n2799 , n478 );
or ( n2800 , n2799 , n456 );
nand ( n2801 , n456 , n462 );
nand ( n2802 , n2800 , n2801 );
buf ( n2803 , n2802 );
not ( n2804 , n2803 );
or ( n2805 , n2798 , n2804 );
or ( n2806 , n2803 , n503 );
nand ( n2807 , n2805 , n2806 );
buf ( n31853 , n2807 );
not ( n2809 , n31853 );
buf ( n31855 , n29969 );
nand ( n2811 , n2809 , n31855 );
buf ( n31857 , n2811 );
buf ( n31858 , n31857 );
nand ( n2814 , n2797 , n31858 );
buf ( n31860 , n2814 );
buf ( n31861 , n31860 );
xor ( n2817 , n31819 , n31861 );
buf ( n31863 , n910 );
not ( n2819 , n31863 );
buf ( n31865 , n497 );
not ( n2821 , n31865 );
buf ( n31867 , n882 );
not ( n2823 , n31867 );
or ( n2824 , n2821 , n2823 );
not ( n2825 , n467 );
and ( n2826 , n456 , n2825 );
not ( n2827 , n456 );
not ( n2828 , n483 );
and ( n2829 , n2827 , n2828 );
nor ( n2830 , n2826 , n2829 );
buf ( n2831 , n2830 );
nand ( n2832 , n2831 , n30599 );
buf ( n31878 , n2832 );
nand ( n2834 , n2824 , n31878 );
buf ( n31880 , n2834 );
buf ( n31881 , n31880 );
not ( n2837 , n31881 );
or ( n2838 , n2819 , n2837 );
buf ( n31884 , n30585 );
buf ( n31885 , n497 );
not ( n2841 , n31885 );
and ( n2842 , n456 , n468 );
not ( n2843 , n456 );
and ( n2844 , n2843 , n484 );
nor ( n2845 , n2842 , n2844 );
buf ( n31891 , n2845 );
not ( n2847 , n31891 );
or ( n2848 , n2841 , n2847 );
buf ( n31894 , n29983 );
buf ( n31895 , n30599 );
nand ( n2851 , n31894 , n31895 );
buf ( n31897 , n2851 );
buf ( n31898 , n31897 );
nand ( n2854 , n2848 , n31898 );
buf ( n31900 , n2854 );
buf ( n31901 , n31900 );
nand ( n2857 , n31884 , n31901 );
buf ( n31903 , n2857 );
buf ( n31904 , n31903 );
nand ( n2860 , n2838 , n31904 );
buf ( n31906 , n2860 );
buf ( n31907 , n31906 );
and ( n2863 , n2817 , n31907 );
and ( n2864 , n31819 , n31861 );
or ( n2865 , n2863 , n2864 );
buf ( n31911 , n2865 );
buf ( n31912 , n31911 );
xor ( n2868 , n2723 , n31912 );
buf ( n31914 , n2868 );
not ( n2870 , n2807 );
buf ( n31916 , n504 );
not ( n2872 , n31916 );
buf ( n31918 , n2872 );
not ( n2874 , n31918 );
and ( n2875 , n2870 , n2874 );
and ( n2876 , n456 , n463 );
not ( n2877 , n456 );
and ( n2878 , n2877 , n479 );
or ( n2879 , n2876 , n2878 );
buf ( n31925 , n2879 );
not ( n2881 , n31925 );
buf ( n31927 , n29987 );
not ( n2883 , n31927 );
and ( n2884 , n2881 , n2883 );
buf ( n31930 , n2879 );
buf ( n31931 , n29987 );
and ( n2887 , n31930 , n31931 );
nor ( n2888 , n2884 , n2887 );
buf ( n31934 , n2888 );
buf ( n31935 , n31934 );
buf ( n31936 , n30347 );
nor ( n2895 , n31935 , n31936 );
buf ( n31938 , n2895 );
nor ( n2897 , n2875 , n31938 );
not ( n2898 , n2897 );
not ( n2899 , n2898 );
buf ( n31942 , n1914 );
not ( n2901 , n31942 );
buf ( n31944 , n2754 );
not ( n2903 , n31944 );
or ( n2904 , n2901 , n2903 );
buf ( n31947 , n495 );
not ( n2906 , n31947 );
buf ( n31949 , n784 );
not ( n2908 , n31949 );
buf ( n31951 , n2908 );
buf ( n31952 , n31951 );
not ( n2911 , n31952 );
or ( n2912 , n2906 , n2911 );
buf ( n31955 , n784 );
buf ( n31956 , n31784 );
nand ( n2915 , n31955 , n31956 );
buf ( n31958 , n2915 );
buf ( n31959 , n31958 );
nand ( n2918 , n2912 , n31959 );
buf ( n31961 , n2918 );
buf ( n31962 , n31961 );
buf ( n31963 , n31812 );
nand ( n2922 , n31962 , n31963 );
buf ( n31965 , n2922 );
buf ( n31966 , n31965 );
nand ( n2925 , n2904 , n31966 );
buf ( n31968 , n2925 );
not ( n2927 , n31968 );
or ( n2928 , n2899 , n2927 );
buf ( n31971 , n31968 );
not ( n2930 , n31971 );
buf ( n31973 , n2930 );
not ( n2932 , n31973 );
not ( n2933 , n2897 );
or ( n2934 , n2932 , n2933 );
buf ( n31977 , n29884 );
not ( n2936 , n31977 );
buf ( n31979 , n499 );
not ( n2938 , n31979 );
not ( n2939 , n466 );
and ( n2940 , n456 , n2939 );
not ( n2941 , n456 );
not ( n2942 , n482 );
and ( n2943 , n2941 , n2942 );
or ( n2944 , n2940 , n2943 );
buf ( n31987 , n2944 );
not ( n2946 , n31987 );
or ( n2947 , n2938 , n2946 );
buf ( n31990 , n933 );
buf ( n31991 , n29901 );
nand ( n2950 , n31990 , n31991 );
buf ( n31993 , n2950 );
buf ( n31994 , n31993 );
nand ( n2953 , n2947 , n31994 );
buf ( n31996 , n2953 );
buf ( n31997 , n31996 );
not ( n2956 , n31997 );
or ( n2957 , n2936 , n2956 );
and ( n2958 , n882 , n499 );
not ( n2959 , n882 );
and ( n2960 , n2959 , n29901 );
or ( n2961 , n2958 , n2960 );
buf ( n32004 , n2961 );
buf ( n32005 , n799 );
nand ( n2964 , n32004 , n32005 );
buf ( n32007 , n2964 );
buf ( n32008 , n32007 );
nand ( n2967 , n2957 , n32008 );
buf ( n32010 , n2967 );
nand ( n2969 , n2934 , n32010 );
nand ( n2970 , n2928 , n2969 );
buf ( n32013 , n2970 );
buf ( n32014 , n30141 );
and ( n2973 , n494 , n495 );
not ( n2974 , n494 );
not ( n2975 , n495 );
and ( n2976 , n2974 , n2975 );
nor ( n2977 , n2973 , n2976 );
buf ( n2978 , n2977 );
buf ( n32021 , n2978 );
and ( n2980 , n32014 , n32021 );
buf ( n32023 , n2980 );
buf ( n32024 , n32023 );
and ( n2983 , n1403 , n501 );
not ( n2984 , n1403 );
and ( n2985 , n2984 , n984 );
nor ( n2986 , n2983 , n2985 );
not ( n2987 , n2986 );
not ( n2988 , n30072 );
nand ( n2989 , n2988 , n960 );
buf ( n32032 , n2989 );
not ( n2991 , n32032 );
buf ( n32034 , n2991 );
not ( n2993 , n32034 );
or ( n2994 , n2987 , n2993 );
nand ( n2995 , n2692 , n1010 );
nand ( n2996 , n2994 , n2995 );
buf ( n32039 , n2996 );
xor ( n2998 , n32024 , n32039 );
buf ( n32041 , n30585 );
not ( n3000 , n32041 );
buf ( n32043 , n497 );
not ( n3002 , n32043 );
buf ( n32045 , n30090 );
not ( n3004 , n32045 );
or ( n3005 , n3002 , n3004 );
buf ( n32048 , n30096 );
buf ( n32049 , n30599 );
nand ( n3008 , n32048 , n32049 );
buf ( n32051 , n3008 );
buf ( n32052 , n32051 );
nand ( n3011 , n3005 , n32052 );
buf ( n32054 , n3011 );
buf ( n32055 , n32054 );
not ( n3014 , n32055 );
or ( n3015 , n3000 , n3014 );
buf ( n32058 , n31900 );
buf ( n32059 , n910 );
nand ( n3018 , n32058 , n32059 );
buf ( n32061 , n3018 );
buf ( n32062 , n32061 );
nand ( n3021 , n3015 , n32062 );
buf ( n32064 , n3021 );
buf ( n32065 , n32064 );
and ( n3024 , n2998 , n32065 );
and ( n3025 , n32024 , n32039 );
or ( n3026 , n3024 , n3025 );
buf ( n32069 , n3026 );
buf ( n32070 , n32069 );
xor ( n3029 , n32013 , n32070 );
xor ( n3030 , n31819 , n31861 );
xor ( n3031 , n3030 , n31907 );
buf ( n32074 , n3031 );
buf ( n32075 , n32074 );
and ( n3034 , n3029 , n32075 );
and ( n3035 , n32013 , n32070 );
or ( n32078 , n3034 , n3035 );
buf ( n32079 , n32078 );
xor ( n3041 , n31914 , n32079 );
buf ( n32081 , n29945 );
xor ( n3043 , n492 , n493 );
not ( n3044 , n3043 );
not ( n3045 , n3044 );
buf ( n32085 , n3045 );
nand ( n3047 , n32081 , n32085 );
buf ( n32087 , n3047 );
buf ( n32088 , n32087 );
not ( n3050 , n32088 );
buf ( n32090 , n3050 );
buf ( n32091 , n32090 );
buf ( n32092 , n910 );
not ( n3054 , n32092 );
buf ( n32094 , n497 );
not ( n3056 , n32094 );
buf ( n32096 , n2944 );
not ( n3058 , n32096 );
or ( n3059 , n3056 , n3058 );
and ( n3060 , n456 , n2939 );
not ( n3061 , n456 );
and ( n3062 , n3061 , n2942 );
nor ( n3063 , n3060 , n3062 );
nand ( n3064 , n3063 , n30599 );
buf ( n32104 , n3064 );
nand ( n3066 , n3059 , n32104 );
buf ( n32106 , n3066 );
buf ( n32107 , n32106 );
not ( n3069 , n32107 );
or ( n3070 , n3054 , n3069 );
buf ( n32110 , n31880 );
nor ( n3072 , n30573 , n1495 );
buf ( n32112 , n3072 );
nand ( n3074 , n32110 , n32112 );
buf ( n32114 , n3074 );
buf ( n32115 , n32114 );
nand ( n3077 , n3070 , n32115 );
buf ( n32117 , n3077 );
buf ( n32118 , n32117 );
xor ( n3080 , n32091 , n32118 );
buf ( n32120 , n1010 );
not ( n3082 , n32120 );
buf ( n32122 , n501 );
not ( n3084 , n32122 );
buf ( n32124 , n2803 );
not ( n3086 , n32124 );
buf ( n32126 , n3086 );
buf ( n32127 , n32126 );
not ( n3089 , n32127 );
or ( n3090 , n3084 , n3089 );
buf ( n32130 , n2803 );
buf ( n32131 , n984 );
nand ( n3093 , n32130 , n32131 );
buf ( n32133 , n3093 );
buf ( n32134 , n32133 );
nand ( n3096 , n3090 , n32134 );
buf ( n32136 , n3096 );
buf ( n32137 , n32136 );
not ( n3099 , n32137 );
or ( n3100 , n3082 , n3099 );
buf ( n32140 , n31734 );
buf ( n32141 , n30078 );
nand ( n3103 , n32140 , n32141 );
buf ( n32143 , n3103 );
buf ( n32144 , n32143 );
nand ( n3106 , n3100 , n32144 );
buf ( n32146 , n3106 );
buf ( n32147 , n32146 );
xor ( n3109 , n3080 , n32147 );
buf ( n32149 , n3109 );
buf ( n32150 , n32149 );
not ( n3112 , n2977 );
not ( n3113 , n3112 );
buf ( n32153 , n3113 );
not ( n3115 , n32153 );
buf ( n32155 , n493 );
not ( n3117 , n32155 );
buf ( n32157 , n29916 );
not ( n3119 , n32157 );
or ( n3120 , n3117 , n3119 );
buf ( n32160 , n784 );
buf ( n32161 , n2704 );
nand ( n3123 , n32160 , n32161 );
buf ( n32163 , n3123 );
buf ( n32164 , n32163 );
nand ( n3126 , n3120 , n32164 );
buf ( n32166 , n3126 );
buf ( n32167 , n32166 );
not ( n3129 , n32167 );
or ( n3130 , n3115 , n3129 );
buf ( n32170 , n493 );
not ( n3132 , n32170 );
buf ( n32172 , n30592 );
not ( n3134 , n32172 );
or ( n3135 , n3132 , n3134 );
buf ( n32175 , n29945 );
buf ( n32176 , n2704 );
nand ( n3138 , n32175 , n32176 );
buf ( n32178 , n3138 );
buf ( n32179 , n32178 );
nand ( n3141 , n3135 , n32179 );
buf ( n32181 , n3141 );
buf ( n32182 , n32181 );
xor ( n3144 , n494 , n493 );
nand ( n3145 , n3112 , n3144 );
not ( n3146 , n3145 );
buf ( n32186 , n3146 );
nand ( n3148 , n32182 , n32186 );
buf ( n32188 , n3148 );
buf ( n32189 , n32188 );
nand ( n3151 , n3130 , n32189 );
buf ( n32191 , n3151 );
not ( n3153 , n32191 );
buf ( n32193 , n29884 );
not ( n3155 , n32193 );
buf ( n32195 , n2637 );
not ( n3157 , n32195 );
or ( n3158 , n3155 , n3157 );
buf ( n32198 , n31996 );
buf ( n32199 , n799 );
nand ( n3161 , n32198 , n32199 );
buf ( n32201 , n3161 );
buf ( n32202 , n32201 );
nand ( n3164 , n3158 , n32202 );
buf ( n32204 , n3164 );
not ( n3166 , n32204 );
or ( n3167 , n3153 , n3166 );
or ( n3168 , n32191 , n32204 );
not ( n3169 , n2720 );
not ( n3170 , n3169 );
not ( n3171 , n2700 );
or ( n32211 , n3170 , n3171 );
nand ( n3176 , n31747 , n2720 );
nand ( n3177 , n32211 , n3176 );
nand ( n3178 , n3168 , n3177 );
nand ( n3179 , n3167 , n3178 );
buf ( n32216 , n3179 );
xor ( n3181 , n32150 , n32216 );
buf ( n32218 , n32166 );
not ( n3183 , n32218 );
buf ( n32220 , n3146 );
not ( n3185 , n32220 );
or ( n3186 , n3183 , n3185 );
buf ( n32223 , n493 );
not ( n3188 , n32223 );
buf ( n32225 , n29512 );
not ( n3190 , n32225 );
or ( n3191 , n3188 , n3190 );
buf ( n32228 , n29513 );
buf ( n32229 , n2704 );
nand ( n3194 , n32228 , n32229 );
buf ( n32231 , n3194 );
buf ( n32232 , n32231 );
nand ( n3197 , n3191 , n32232 );
buf ( n32234 , n3197 );
buf ( n32235 , n32234 );
buf ( n32236 , n2978 );
nand ( n3201 , n32235 , n32236 );
buf ( n32238 , n3201 );
buf ( n32239 , n32238 );
nand ( n3204 , n3186 , n32239 );
buf ( n32241 , n3204 );
buf ( n32242 , n503 );
not ( n3207 , n32242 );
and ( n3208 , n456 , n460 );
not ( n3209 , n456 );
and ( n3210 , n3209 , n476 );
nor ( n3211 , n3208 , n3210 );
buf ( n32248 , n3211 );
not ( n3213 , n32248 );
or ( n3214 , n3207 , n3213 );
not ( n3215 , n460 );
and ( n3216 , n456 , n3215 );
not ( n3217 , n456 );
not ( n3218 , n476 );
and ( n3219 , n3217 , n3218 );
nor ( n3220 , n3216 , n3219 );
buf ( n32257 , n3220 );
buf ( n32258 , n29987 );
nand ( n3223 , n32257 , n32258 );
buf ( n32260 , n3223 );
buf ( n32261 , n32260 );
nand ( n3226 , n3214 , n32261 );
buf ( n32263 , n3226 );
buf ( n32264 , n32263 );
not ( n3229 , n32264 );
buf ( n32266 , n3229 );
buf ( n32267 , n32266 );
not ( n3232 , n32267 );
buf ( n32269 , n31918 );
not ( n3234 , n32269 );
and ( n3235 , n3232 , n3234 );
buf ( n32272 , n31839 );
buf ( n32273 , n29969 );
and ( n3238 , n32272 , n32273 );
nor ( n3239 , n3235 , n3238 );
buf ( n32276 , n3239 );
buf ( n32277 , n32276 );
buf ( n32278 , n31812 );
not ( n3243 , n32278 );
buf ( n32280 , n3243 );
buf ( n32281 , n32280 );
not ( n3246 , n32281 );
buf ( n32283 , n31790 );
not ( n3248 , n32283 );
buf ( n32285 , n3248 );
buf ( n32286 , n32285 );
not ( n3251 , n32286 );
and ( n3252 , n3246 , n3251 );
buf ( n32289 , n495 );
buf ( n32290 , n29507 );
not ( n3255 , n32290 );
buf ( n32292 , n3255 );
buf ( n32293 , n32292 );
and ( n3258 , n32289 , n32293 );
not ( n3259 , n32289 );
buf ( n32296 , n32292 );
not ( n3261 , n32296 );
buf ( n32298 , n3261 );
buf ( n32299 , n32298 );
and ( n3264 , n3259 , n32299 );
nor ( n3265 , n3258 , n3264 );
buf ( n32302 , n3265 );
buf ( n32303 , n32302 );
not ( n3268 , n32303 );
buf ( n32305 , n3268 );
buf ( n32306 , n32305 );
not ( n3271 , n2724 );
buf ( n32308 , n3271 );
and ( n3273 , n32306 , n32308 );
nor ( n3274 , n3252 , n3273 );
buf ( n32311 , n3274 );
buf ( n32312 , n32311 );
and ( n3277 , n32277 , n32312 );
not ( n3278 , n32277 );
not ( n3279 , n32311 );
buf ( n32316 , n3279 );
and ( n3281 , n3278 , n32316 );
nor ( n3282 , n3277 , n3281 );
buf ( n32319 , n3282 );
xor ( n3284 , n32241 , n32319 );
buf ( n32321 , n3284 );
xor ( n3286 , n3181 , n32321 );
buf ( n32323 , n3286 );
xor ( n3288 , n3041 , n32323 );
not ( n3289 , n3288 );
xor ( n3290 , n32191 , n32204 );
xor ( n3291 , n3290 , n3177 );
buf ( n32328 , n31761 );
not ( n3293 , n32328 );
buf ( n32330 , n3293 );
buf ( n32331 , n32330 );
buf ( n32332 , n496 );
and ( n3297 , n32331 , n32332 );
buf ( n32334 , n31784 );
nor ( n3302 , n3297 , n32334 );
buf ( n32336 , n3302 );
buf ( n32337 , n32336 );
buf ( n32338 , n1912 );
not ( n3306 , n32338 );
buf ( n32340 , n29939 );
not ( n3308 , n32340 );
buf ( n32342 , n3308 );
buf ( n32343 , n32342 );
not ( n3311 , n32343 );
or ( n3312 , n3306 , n3311 );
buf ( n32346 , n497 );
nand ( n3314 , n3312 , n32346 );
buf ( n32348 , n3314 );
buf ( n32349 , n32348 );
and ( n3317 , n32337 , n32349 );
buf ( n32351 , n3317 );
buf ( n32352 , n32351 );
buf ( n32353 , n30078 );
not ( n3321 , n32353 );
buf ( n32355 , n31061 );
not ( n3323 , n32355 );
or ( n3324 , n3321 , n3323 );
buf ( n32358 , n1010 );
and ( n3326 , n1403 , n984 );
not ( n3327 , n1403 );
and ( n3328 , n3327 , n501 );
or ( n3329 , n3326 , n3328 );
buf ( n32363 , n3329 );
nand ( n3331 , n32358 , n32363 );
buf ( n32365 , n3331 );
buf ( n32366 , n32365 );
nand ( n3334 , n3324 , n32366 );
buf ( n32368 , n3334 );
buf ( n32369 , n32368 );
and ( n3337 , n32352 , n32369 );
buf ( n32371 , n3337 );
buf ( n32372 , n32371 );
xor ( n3340 , n32024 , n32039 );
xor ( n3341 , n3340 , n32065 );
buf ( n32375 , n3341 );
buf ( n32376 , n32375 );
xor ( n3344 , n32372 , n32376 );
not ( n3345 , n31812 );
and ( n3346 , n31784 , n31761 );
not ( n3347 , n31784 );
buf ( n32381 , n30592 );
not ( n3349 , n32381 );
buf ( n32383 , n3349 );
and ( n3351 , n3347 , n32383 );
nor ( n3352 , n3346 , n3351 );
not ( n3353 , n3352 );
or ( n3354 , n3345 , n3353 );
buf ( n32388 , n31961 );
buf ( n32389 , n1914 );
nand ( n32390 , n32388 , n32389 );
buf ( n32391 , n32390 );
nand ( n3359 , n3354 , n32391 );
buf ( n32393 , n29969 );
not ( n3361 , n32393 );
buf ( n32395 , n30962 );
not ( n3363 , n32395 );
or ( n3364 , n3361 , n3363 );
not ( n3365 , n31934 );
nand ( n3366 , n3365 , n504 );
buf ( n32400 , n3366 );
nand ( n3368 , n3364 , n32400 );
buf ( n32402 , n3368 );
xor ( n3370 , n3359 , n32402 );
buf ( n32404 , n910 );
not ( n3372 , n32404 );
buf ( n32406 , n32054 );
not ( n3374 , n32406 );
or ( n3375 , n3372 , n3374 );
buf ( n32409 , n31004 );
buf ( n32410 , n30585 );
nand ( n3378 , n32409 , n32410 );
buf ( n32412 , n3378 );
buf ( n32413 , n32412 );
nand ( n3381 , n3375 , n32413 );
buf ( n32415 , n3381 );
and ( n3383 , n3370 , n32415 );
and ( n3384 , n3359 , n32402 );
or ( n3385 , n3383 , n3384 );
buf ( n32419 , n3385 );
and ( n3387 , n3344 , n32419 );
and ( n3388 , n32372 , n32376 );
or ( n3389 , n3387 , n3388 );
buf ( n32423 , n3389 );
xor ( n3391 , n3291 , n32423 );
xor ( n3392 , n32013 , n32070 );
xor ( n3393 , n3392 , n32075 );
buf ( n32427 , n3393 );
and ( n3395 , n3391 , n32427 );
and ( n3396 , n3291 , n32423 );
or ( n3397 , n3395 , n3396 );
not ( n3398 , n3397 );
and ( n3399 , n3289 , n3398 );
buf ( n32433 , n492 );
not ( n3401 , n32433 );
buf ( n32435 , n30592 );
nand ( n3403 , n3401 , n32435 );
buf ( n32437 , n3403 );
buf ( n32438 , n32437 );
buf ( n32439 , n493 );
and ( n3407 , n32438 , n32439 );
buf ( n32441 , n492 );
not ( n3409 , n32441 );
buf ( n32443 , n29939 );
not ( n3411 , n32443 );
or ( n32445 , n3409 , n3411 );
buf ( n32446 , n491 );
nand ( n3417 , n32445 , n32446 );
buf ( n32448 , n3417 );
buf ( n32449 , n32448 );
nor ( n3420 , n3407 , n32449 );
buf ( n32451 , n3420 );
buf ( n32452 , n32451 );
buf ( n32453 , n29969 );
not ( n3424 , n32453 );
buf ( n32455 , n32263 );
not ( n3426 , n32455 );
or ( n3427 , n3424 , n3426 );
buf ( n32458 , n503 );
not ( n3429 , n32458 );
and ( n3430 , n456 , n459 );
not ( n3431 , n456 );
and ( n3432 , n3431 , n475 );
nor ( n3433 , n3430 , n3432 );
not ( n3434 , n3433 );
buf ( n32465 , n3434 );
not ( n3436 , n32465 );
buf ( n32467 , n3436 );
buf ( n32468 , n32467 );
not ( n3439 , n32468 );
or ( n3440 , n3429 , n3439 );
buf ( n32471 , n3434 );
buf ( n32472 , n29987 );
nand ( n3443 , n32471 , n32472 );
buf ( n32474 , n3443 );
buf ( n32475 , n32474 );
nand ( n3446 , n3440 , n32475 );
buf ( n32477 , n3446 );
buf ( n32478 , n32477 );
buf ( n32479 , n504 );
nand ( n3450 , n32478 , n32479 );
buf ( n32481 , n3450 );
buf ( n32482 , n32481 );
nand ( n3453 , n3427 , n32482 );
buf ( n32484 , n3453 );
buf ( n32485 , n32484 );
xor ( n3456 , n32452 , n32485 );
buf ( n32487 , n3456 );
buf ( n32488 , n32487 );
xor ( n3459 , n32091 , n32118 );
and ( n3460 , n3459 , n32147 );
and ( n3461 , n32091 , n32118 );
or ( n3462 , n3460 , n3461 );
buf ( n32493 , n3462 );
buf ( n32494 , n32493 );
xor ( n3465 , n32488 , n32494 );
buf ( n32496 , n3279 );
not ( n32497 , n32496 );
buf ( n32498 , n32276 );
not ( n3469 , n32498 );
buf ( n32500 , n3469 );
buf ( n32501 , n32500 );
not ( n3472 , n32501 );
or ( n3473 , n32497 , n3472 );
buf ( n32504 , n32276 );
not ( n3475 , n32504 );
buf ( n32506 , n32311 );
not ( n3477 , n32506 );
or ( n3478 , n3475 , n3477 );
buf ( n32509 , n32241 );
nand ( n3480 , n3478 , n32509 );
buf ( n32511 , n3480 );
buf ( n32512 , n32511 );
nand ( n3483 , n3473 , n32512 );
buf ( n32514 , n3483 );
buf ( n32515 , n32514 );
xor ( n3486 , n3465 , n32515 );
buf ( n32517 , n3486 );
xor ( n3488 , n32150 , n32216 );
and ( n3489 , n3488 , n32321 );
and ( n3490 , n32150 , n32216 );
or ( n3491 , n3489 , n3490 );
buf ( n32522 , n3491 );
xor ( n3493 , n32517 , n32522 );
buf ( n32524 , n2978 );
not ( n3495 , n32524 );
buf ( n32526 , n493 );
not ( n3497 , n32526 );
buf ( n32528 , n30090 );
not ( n3499 , n32528 );
or ( n3500 , n3497 , n3499 );
buf ( n32531 , n973 );
buf ( n32532 , n2704 );
nand ( n3503 , n32531 , n32532 );
buf ( n32534 , n3503 );
buf ( n32535 , n32534 );
nand ( n3506 , n3500 , n32535 );
buf ( n32537 , n3506 );
buf ( n32538 , n32537 );
not ( n3509 , n32538 );
or ( n3510 , n3495 , n3509 );
not ( n3511 , n3145 );
nand ( n3512 , n32234 , n3511 );
buf ( n32543 , n3512 );
nand ( n3514 , n3510 , n32543 );
buf ( n32545 , n3514 );
not ( n3516 , n32545 );
buf ( n32547 , n3043 );
not ( n32548 , n32547 );
buf ( n32549 , n784 );
not ( n3523 , n32549 );
not ( n3524 , n491 );
buf ( n32552 , n3524 );
not ( n3526 , n32552 );
and ( n3527 , n3523 , n3526 );
buf ( n32555 , n784 );
buf ( n32556 , n3524 );
and ( n3530 , n32555 , n32556 );
nor ( n3531 , n3527 , n3530 );
buf ( n32559 , n3531 );
buf ( n32560 , n32559 );
nor ( n3534 , n32548 , n32560 );
buf ( n32562 , n3534 );
buf ( n32563 , n32562 );
buf ( n32564 , n29939 );
not ( n3538 , n32564 );
buf ( n32566 , n3524 );
not ( n3540 , n32566 );
and ( n3541 , n3538 , n3540 );
buf ( n32569 , n29939 );
buf ( n32570 , n3524 );
and ( n3544 , n32569 , n32570 );
nor ( n3545 , n3541 , n3544 );
buf ( n32573 , n3545 );
buf ( n32574 , n32573 );
not ( n3548 , n3043 );
and ( n3549 , n491 , n492 );
not ( n3550 , n491 );
not ( n3551 , n492 );
and ( n3552 , n3550 , n3551 );
nor ( n3553 , n3549 , n3552 );
nand ( n3554 , n3548 , n3553 );
buf ( n32582 , n3554 );
nor ( n3556 , n32574 , n32582 );
buf ( n32584 , n3556 );
buf ( n32585 , n32584 );
nor ( n3559 , n32563 , n32585 );
buf ( n32587 , n3559 );
not ( n3561 , n32587 );
not ( n3562 , n3561 );
or ( n3563 , n3516 , n3562 );
buf ( n32591 , n32545 );
not ( n3565 , n32591 );
buf ( n32593 , n3565 );
nand ( n32594 , n32593 , n32587 );
nand ( n3568 , n3563 , n32594 );
buf ( n32596 , n29901 );
buf ( n32597 , n2679 );
and ( n3571 , n32596 , n32597 );
not ( n3572 , n32596 );
buf ( n32600 , n2671 );
and ( n3574 , n3572 , n32600 );
nor ( n3575 , n3571 , n3574 );
buf ( n32603 , n3575 );
not ( n3577 , n32603 );
not ( n3578 , n745 );
not ( n3579 , n3578 );
and ( n3580 , n3577 , n3579 );
and ( n3581 , n31703 , n799 );
nor ( n3582 , n3580 , n3581 );
and ( n3583 , n3568 , n3582 );
not ( n3584 , n3568 );
not ( n3585 , n3582 );
and ( n3586 , n3584 , n3585 );
nor ( n3587 , n3583 , n3586 );
buf ( n32615 , n30585 );
not ( n3589 , n32615 );
buf ( n32617 , n32106 );
not ( n3591 , n32617 );
or ( n3592 , n3589 , n3591 );
not ( n3593 , n497 );
and ( n3594 , n456 , n465 );
not ( n3595 , n456 );
and ( n3596 , n3595 , n481 );
nor ( n3597 , n3594 , n3596 );
not ( n3598 , n3597 );
or ( n3599 , n3593 , n3598 );
buf ( n32627 , n1403 );
buf ( n32628 , n30599 );
nand ( n3602 , n32627 , n32628 );
buf ( n32630 , n3602 );
nand ( n3604 , n3599 , n32630 );
nand ( n3605 , n3604 , n909 );
buf ( n32633 , n3605 );
nand ( n3607 , n3592 , n32633 );
buf ( n32635 , n3607 );
buf ( n32636 , n31809 );
not ( n3610 , n32636 );
buf ( n32638 , n32302 );
not ( n32639 , n32638 );
and ( n3616 , n3610 , n32639 );
buf ( n32641 , n495 );
not ( n3618 , n32641 );
buf ( n32643 , n882 );
not ( n3620 , n32643 );
or ( n3621 , n3618 , n3620 );
nand ( n3622 , n2831 , n31784 );
buf ( n32647 , n3622 );
nand ( n3624 , n3621 , n32647 );
buf ( n32649 , n3624 );
buf ( n32650 , n32649 );
buf ( n32651 , n3271 );
and ( n3628 , n32650 , n32651 );
nor ( n3629 , n3616 , n3628 );
buf ( n32654 , n3629 );
xor ( n3631 , n32635 , n32654 );
buf ( n32656 , n501 );
not ( n3633 , n32656 );
buf ( n32658 , n29493 );
not ( n3635 , n32658 );
buf ( n32660 , n3635 );
buf ( n32661 , n32660 );
not ( n3638 , n32661 );
or ( n3639 , n3633 , n3638 );
buf ( n32664 , n31826 );
buf ( n32665 , n984 );
nand ( n3642 , n32664 , n32665 );
buf ( n32667 , n3642 );
buf ( n32668 , n32667 );
nand ( n3645 , n3639 , n32668 );
buf ( n32670 , n3645 );
buf ( n32671 , n32670 );
buf ( n32672 , n1010 );
and ( n3649 , n32671 , n32672 );
buf ( n32674 , n32136 );
buf ( n32675 , n30078 );
and ( n3652 , n32674 , n32675 );
nor ( n3653 , n3649 , n3652 );
buf ( n32678 , n3653 );
xor ( n3655 , n3631 , n32678 );
xor ( n3656 , n3587 , n3655 );
xor ( n32681 , n31711 , n31770 );
and ( n3658 , n32681 , n31912 );
and ( n3659 , n31711 , n31770 );
or ( n3660 , n3658 , n3659 );
buf ( n32685 , n3660 );
xor ( n3662 , n3656 , n32685 );
xor ( n3663 , n3493 , n3662 );
not ( n3664 , n3663 );
xor ( n3665 , n31914 , n32079 );
and ( n3666 , n3665 , n32323 );
and ( n3667 , n31914 , n32079 );
or ( n3668 , n3666 , n3667 );
not ( n3669 , n3668 );
and ( n3670 , n3664 , n3669 );
nor ( n3671 , n3399 , n3670 );
not ( n3672 , n3671 );
xor ( n3673 , n3291 , n32423 );
xor ( n3674 , n3673 , n32427 );
not ( n3675 , n3674 );
xor ( n3676 , n31968 , n2898 );
xor ( n3677 , n3676 , n32010 );
buf ( n32702 , n3677 );
buf ( n32703 , n29884 );
not ( n3680 , n32703 );
buf ( n32705 , n2961 );
not ( n3682 , n32705 );
or ( n3683 , n3680 , n3682 );
buf ( n32708 , n798 );
not ( n3685 , n32708 );
buf ( n32710 , n1973 );
nand ( n3687 , n3685 , n32710 );
buf ( n32712 , n3687 );
buf ( n32713 , n32712 );
nand ( n3690 , n3683 , n32713 );
buf ( n32715 , n3690 );
buf ( n32716 , n32715 );
xor ( n3693 , n32352 , n32369 );
buf ( n32718 , n3693 );
buf ( n32719 , n32718 );
xor ( n3696 , n32716 , n32719 );
buf ( n32721 , n30988 );
not ( n32722 , n32721 );
buf ( n32723 , n30972 );
not ( n3703 , n32723 );
or ( n3704 , n32722 , n3703 );
buf ( n32726 , n504 );
not ( n3706 , n32726 );
buf ( n32728 , n30962 );
not ( n3708 , n32728 );
or ( n3709 , n3706 , n3708 );
buf ( n32731 , n30969 );
nand ( n3711 , n3709 , n32731 );
buf ( n32733 , n3711 );
buf ( n32734 , n32733 );
buf ( n32735 , n30988 );
or ( n3715 , n32734 , n32735 );
buf ( n32737 , n31014 );
nand ( n3717 , n3715 , n32737 );
buf ( n32739 , n3717 );
buf ( n32740 , n32739 );
nand ( n3720 , n3704 , n32740 );
buf ( n32742 , n3720 );
buf ( n32743 , n32742 );
and ( n3723 , n3696 , n32743 );
and ( n3724 , n32716 , n32719 );
or ( n3725 , n3723 , n3724 );
buf ( n32747 , n3725 );
buf ( n32748 , n32747 );
xor ( n3728 , n32702 , n32748 );
xor ( n3729 , n32372 , n32376 );
xor ( n3730 , n3729 , n32419 );
buf ( n32752 , n3730 );
buf ( n32753 , n32752 );
and ( n3733 , n3728 , n32753 );
and ( n3734 , n32702 , n32748 );
or ( n3735 , n3733 , n3734 );
buf ( n32757 , n3735 );
not ( n32758 , n32757 );
nand ( n3738 , n3675 , n32758 );
xor ( n3739 , n32702 , n32748 );
xor ( n3740 , n3739 , n32753 );
buf ( n32762 , n3740 );
xor ( n3742 , n3359 , n32402 );
xor ( n3743 , n3742 , n32415 );
buf ( n32765 , n3743 );
xor ( n3745 , n31047 , n31072 );
and ( n3746 , n3745 , n31078 );
and ( n3747 , n31047 , n31072 );
or ( n3748 , n3746 , n3747 );
buf ( n32770 , n3748 );
buf ( n32771 , n32770 );
xor ( n3751 , n32765 , n32771 );
xor ( n3752 , n32716 , n32719 );
xor ( n3753 , n3752 , n32743 );
buf ( n32775 , n3753 );
buf ( n32776 , n32775 );
and ( n3756 , n3751 , n32776 );
and ( n3757 , n32765 , n32771 );
or ( n3758 , n3756 , n3757 );
buf ( n32780 , n3758 );
nor ( n3760 , n32762 , n32780 );
not ( n3761 , n3760 );
not ( n3762 , n2028 );
xor ( n3763 , n31023 , n31029 );
and ( n3764 , n3763 , n31081 );
and ( n3765 , n31023 , n31029 );
or ( n3766 , n3764 , n3765 );
buf ( n32788 , n3766 );
not ( n3768 , n32788 );
xor ( n3769 , n32765 , n32771 );
xor ( n3770 , n3769 , n32776 );
buf ( n32792 , n3770 );
not ( n32793 , n32792 );
nand ( n3776 , n3768 , n32793 );
nand ( n3777 , n3762 , n3776 );
not ( n3778 , n3777 );
nand ( n3779 , n3738 , n1875 , n3761 , n3778 );
nand ( n3780 , n32792 , n32788 );
not ( n3781 , n3780 );
not ( n3782 , n2026 );
or ( n3783 , n3781 , n3782 );
nand ( n3784 , n3783 , n3776 );
nor ( n3785 , n3760 , n3784 );
nand ( n3786 , n3674 , n32757 );
nand ( n3787 , n32762 , n32780 );
nand ( n3788 , n3786 , n3787 );
or ( n3789 , n3785 , n3788 );
nand ( n3790 , n3789 , n3738 );
nand ( n3791 , n3779 , n3790 );
not ( n3792 , n3791 );
or ( n3793 , n3672 , n3792 );
nor ( n3794 , n3668 , n3663 );
nand ( n3795 , n3288 , n3397 );
or ( n3796 , n3794 , n3795 );
nand ( n3797 , n3663 , n3668 );
nand ( n3798 , n3796 , n3797 );
not ( n3799 , n3798 );
nand ( n3800 , n3793 , n3799 );
not ( n3801 , n32635 );
nand ( n3802 , n32678 , n32654 );
not ( n3803 , n3802 );
or ( n3804 , n3801 , n3803 );
buf ( n32823 , n32678 );
not ( n3806 , n32823 );
buf ( n32825 , n3806 );
buf ( n32826 , n32654 );
not ( n3809 , n32826 );
buf ( n32828 , n3809 );
nand ( n3811 , n32825 , n32828 );
nand ( n3812 , n3804 , n3811 );
buf ( n32831 , n3812 );
not ( n3814 , n32831 );
not ( n3815 , n32593 );
not ( n3816 , n3582 );
and ( n3817 , n3815 , n3816 );
and ( n3818 , n32593 , n3582 );
nor ( n3819 , n3818 , n32587 );
nor ( n3820 , n3817 , n3819 );
buf ( n32839 , n3820 );
not ( n3822 , n32839 );
and ( n3823 , n3814 , n3822 );
buf ( n32842 , n3820 );
buf ( n32843 , n3812 );
and ( n3826 , n32842 , n32843 );
nor ( n3827 , n3823 , n3826 );
buf ( n32846 , n3827 );
buf ( n32847 , n29939 );
not ( n3830 , n32847 );
buf ( n32849 , n3830 );
xor ( n3832 , n490 , n491 );
not ( n3833 , n3832 );
nor ( n3834 , n32849 , n3833 );
buf ( n32853 , n3834 );
buf ( n32854 , n29969 );
not ( n3837 , n32854 );
buf ( n32856 , n32477 );
not ( n3842 , n32856 );
or ( n3843 , n3837 , n3842 );
not ( n3844 , n503 );
and ( n3845 , n456 , n458 );
not ( n3846 , n456 );
and ( n3847 , n3846 , n474 );
nor ( n3848 , n3845 , n3847 );
not ( n3849 , n3848 );
or ( n3850 , n3844 , n3849 );
and ( n3851 , n456 , n458 );
not ( n3852 , n456 );
and ( n3853 , n3852 , n474 );
nor ( n3854 , n3851 , n3853 );
not ( n3855 , n3854 );
nand ( n3856 , n3855 , n29987 );
nand ( n3857 , n3850 , n3856 );
buf ( n32873 , n3857 );
buf ( n32874 , n504 );
nand ( n3860 , n32873 , n32874 );
buf ( n32876 , n3860 );
buf ( n32877 , n32876 );
nand ( n3863 , n3843 , n32877 );
buf ( n32879 , n3863 );
buf ( n32880 , n32879 );
xor ( n3866 , n32853 , n32880 );
buf ( n32882 , n1010 );
not ( n3868 , n32882 );
not ( n3869 , n3220 );
not ( n3870 , n984 );
or ( n3871 , n3869 , n3870 );
nand ( n3872 , n501 , n3211 );
nand ( n3873 , n3871 , n3872 );
buf ( n32889 , n3873 );
not ( n3875 , n32889 );
or ( n3876 , n3868 , n3875 );
buf ( n32892 , n32670 );
buf ( n32893 , n30078 );
nand ( n3879 , n32892 , n32893 );
buf ( n32895 , n3879 );
buf ( n32896 , n32895 );
nand ( n3882 , n3876 , n32896 );
buf ( n32898 , n3882 );
buf ( n32899 , n32898 );
xor ( n3885 , n3866 , n32899 );
buf ( n32901 , n3885 );
buf ( n32902 , n32901 );
buf ( n3888 , n32902 );
buf ( n32904 , n3888 );
not ( n3890 , n32904 );
and ( n3891 , n32846 , n3890 );
not ( n32907 , n32846 );
and ( n3896 , n32907 , n32904 );
nor ( n3897 , n3891 , n3896 );
xor ( n3898 , n3587 , n3655 );
and ( n3899 , n3898 , n32685 );
and ( n3900 , n3587 , n3655 );
or ( n3901 , n3899 , n3900 );
xor ( n3902 , n3897 , n3901 );
buf ( n32915 , n3146 );
not ( n3904 , n32915 );
buf ( n32917 , n32537 );
not ( n3906 , n32917 );
or ( n3907 , n3904 , n3906 );
not ( n3908 , n493 );
not ( n3909 , n854 );
or ( n3910 , n3908 , n3909 );
buf ( n32923 , n29507 );
buf ( n32924 , n2704 );
nand ( n3913 , n32923 , n32924 );
buf ( n32926 , n3913 );
nand ( n3915 , n3910 , n32926 );
buf ( n32928 , n3915 );
buf ( n32929 , n3113 );
nand ( n3918 , n32928 , n32929 );
buf ( n32931 , n3918 );
buf ( n32932 , n32931 );
nand ( n3921 , n3907 , n32932 );
buf ( n32934 , n3921 );
buf ( n32935 , n32934 );
buf ( n32936 , n3045 );
not ( n3925 , n32936 );
buf ( n32938 , n491 );
not ( n3927 , n32938 );
buf ( n32940 , n29897 );
not ( n3929 , n32940 );
or ( n3930 , n3927 , n3929 );
buf ( n32943 , n29514 );
buf ( n32944 , n3524 );
nand ( n3933 , n32943 , n32944 );
buf ( n32946 , n3933 );
buf ( n32947 , n32946 );
nand ( n3936 , n3930 , n32947 );
buf ( n32949 , n3936 );
buf ( n32950 , n32949 );
not ( n3942 , n32950 );
or ( n3943 , n3925 , n3942 );
buf ( n32953 , n32559 );
not ( n3945 , n32953 );
not ( n3946 , n3043 );
nand ( n3947 , n3946 , n3553 );
not ( n3948 , n3947 );
buf ( n32958 , n3948 );
nand ( n3950 , n3945 , n32958 );
buf ( n32960 , n3950 );
buf ( n32961 , n32960 );
nand ( n3953 , n3943 , n32961 );
buf ( n32963 , n3953 );
buf ( n32964 , n32963 );
xor ( n3956 , n32935 , n32964 );
and ( n32966 , n32452 , n32485 );
buf ( n32967 , n32966 );
buf ( n32968 , n32967 );
xor ( n3960 , n3956 , n32968 );
buf ( n32970 , n3960 );
not ( n3962 , n745 );
not ( n3963 , n29901 );
buf ( n32973 , n2803 );
not ( n3965 , n32973 );
buf ( n32975 , n3965 );
not ( n3967 , n32975 );
not ( n3968 , n3967 );
or ( n3969 , n3963 , n3968 );
nand ( n3970 , n32126 , n499 );
nand ( n3971 , n3969 , n3970 );
not ( n32981 , n3971 );
or ( n3976 , n3962 , n32981 );
not ( n32983 , n32603 );
nand ( n3978 , n32983 , n799 );
nand ( n32985 , n3976 , n3978 );
not ( n3980 , n32985 );
not ( n3981 , n3271 );
not ( n3982 , n495 );
not ( n32989 , n929 );
or ( n32990 , n3982 , n32989 );
buf ( n32991 , n933 );
buf ( n32992 , n31784 );
nand ( n3987 , n32991 , n32992 );
buf ( n32994 , n3987 );
nand ( n3989 , n32990 , n32994 );
not ( n3990 , n3989 );
or ( n3991 , n3981 , n3990 );
buf ( n32998 , n32649 );
buf ( n32999 , n31812 );
nand ( n3994 , n32998 , n32999 );
buf ( n33001 , n3994 );
nand ( n3996 , n3991 , n33001 );
not ( n3997 , n3996 );
not ( n3998 , n3604 );
not ( n33005 , n3072 );
or ( n4000 , n3998 , n33005 );
and ( n4001 , n29501 , n497 );
not ( n33008 , n29501 );
and ( n4003 , n33008 , n30599 );
nor ( n4004 , n4001 , n4003 );
not ( n4005 , n4004 );
buf ( n33012 , n909 );
not ( n33013 , n33012 );
buf ( n33014 , n33013 );
or ( n4009 , n4005 , n33014 );
nand ( n4010 , n4000 , n4009 );
nand ( n4011 , n3980 , n3997 , n4010 );
not ( n33018 , n4010 );
not ( n4013 , n745 );
not ( n4014 , n3971 );
or ( n4015 , n4013 , n4014 );
nand ( n4016 , n4015 , n3978 );
nand ( n4017 , n33018 , n4016 , n3997 );
not ( n33024 , n33018 );
nand ( n4019 , n33024 , n3996 , n4016 );
not ( n4020 , n3997 );
not ( n4021 , n4016 );
nand ( n4022 , n4020 , n4021 , n33018 );
nand ( n4023 , n4011 , n4017 , n4019 , n4022 );
xor ( n4024 , n32970 , n4023 );
xor ( n33031 , n32488 , n32494 );
and ( n4026 , n33031 , n32515 );
and ( n4027 , n32488 , n32494 );
or ( n4028 , n4026 , n4027 );
buf ( n33035 , n4028 );
xor ( n4030 , n4024 , n33035 );
xor ( n33037 , n3902 , n4030 );
xor ( n4032 , n32517 , n32522 );
and ( n4033 , n4032 , n3662 );
and ( n33040 , n32517 , n32522 );
or ( n4035 , n4033 , n33040 );
or ( n33042 , n33037 , n4035 );
nand ( n4037 , n33037 , n4035 );
nand ( n4038 , n33042 , n4037 );
nand ( n4039 , n3800 , n4038 , n455 );
not ( n4040 , n4039 );
buf ( n33047 , n508 );
not ( n33048 , n33047 );
buf ( n33049 , n33048 );
and ( n4044 , n503 , n33049 );
not ( n4045 , n503 );
and ( n4046 , n4045 , n508 );
or ( n4047 , n4044 , n4046 );
buf ( n33054 , n4047 );
not ( n4049 , n33054 );
buf ( n33056 , n29734 );
not ( n4051 , n33056 );
or ( n33058 , n4049 , n4051 );
and ( n4053 , n507 , n503 );
not ( n4054 , n507 );
and ( n4055 , n4054 , n956 );
nor ( n4056 , n4053 , n4055 );
buf ( n33063 , n4056 );
buf ( n33064 , n504 );
nand ( n4059 , n33063 , n33064 );
buf ( n33066 , n4059 );
buf ( n33067 , n33066 );
nand ( n4062 , n33058 , n33067 );
buf ( n33069 , n4062 );
buf ( n33070 , n33069 );
not ( n4065 , n33070 );
buf ( n33072 , n520 );
buf ( n33073 , n492 );
or ( n4068 , n33072 , n33073 );
buf ( n33075 , n493 );
nand ( n4070 , n4068 , n33075 );
buf ( n33077 , n4070 );
buf ( n33078 , n33077 );
buf ( n33079 , n520 );
buf ( n33080 , n492 );
nand ( n4075 , n33079 , n33080 );
buf ( n33082 , n4075 );
buf ( n33083 , n33082 );
buf ( n33084 , n491 );
and ( n4079 , n33078 , n33083 , n33084 );
buf ( n33086 , n4079 );
buf ( n33087 , n33086 );
not ( n4082 , n33087 );
buf ( n33089 , n4082 );
buf ( n33090 , n33089 );
not ( n4085 , n33090 );
or ( n4086 , n4065 , n4085 );
buf ( n33093 , n33089 );
buf ( n33094 , n33069 );
or ( n4089 , n33093 , n33094 );
nand ( n4090 , n4086 , n4089 );
buf ( n33097 , n4090 );
buf ( n33098 , n33097 );
buf ( n33099 , n492 );
buf ( n33100 , n493 );
xor ( n4095 , n33099 , n33100 );
buf ( n33102 , n4095 );
buf ( n33103 , n33102 );
buf ( n33104 , n520 );
and ( n4099 , n33103 , n33104 );
buf ( n33106 , n4099 );
buf ( n33107 , n33106 );
xor ( n4102 , n497 , n515 );
buf ( n33109 , n4102 );
not ( n4104 , n33109 );
buf ( n33111 , n1691 );
not ( n4106 , n33111 );
or ( n4107 , n4104 , n4106 );
buf ( n33114 , n1786 );
xor ( n4109 , n497 , n514 );
buf ( n33116 , n4109 );
nand ( n4111 , n33114 , n33116 );
buf ( n33118 , n4111 );
buf ( n33119 , n33118 );
nand ( n4114 , n4107 , n33119 );
buf ( n33121 , n4114 );
buf ( n33122 , n33121 );
xor ( n4117 , n33107 , n33122 );
xor ( n4118 , n501 , n511 );
buf ( n33125 , n4118 );
not ( n4120 , n33125 );
buf ( n33127 , n29640 );
not ( n33128 , n33127 );
or ( n4123 , n4120 , n33128 );
buf ( n33130 , n29649 );
buf ( n33131 , n510 );
buf ( n33132 , n501 );
xor ( n4127 , n33131 , n33132 );
buf ( n33134 , n4127 );
buf ( n33135 , n33134 );
nand ( n4130 , n33130 , n33135 );
buf ( n33137 , n4130 );
buf ( n33138 , n33137 );
nand ( n4133 , n4123 , n33138 );
buf ( n33140 , n4133 );
buf ( n33141 , n33140 );
and ( n33142 , n4117 , n33141 );
and ( n4137 , n33107 , n33122 );
or ( n33144 , n33142 , n4137 );
buf ( n33145 , n33144 );
buf ( n33146 , n33145 );
xor ( n33147 , n33098 , n33146 );
buf ( n33148 , n509 );
buf ( n33149 , n503 );
xor ( n33150 , n33148 , n33149 );
buf ( n33151 , n33150 );
buf ( n33152 , n33151 );
not ( n33153 , n33152 );
buf ( n33154 , n29582 );
not ( n4149 , n33154 );
or ( n33156 , n33153 , n4149 );
buf ( n33157 , n4047 );
buf ( n33158 , n504 );
nand ( n4153 , n33157 , n33158 );
buf ( n33160 , n4153 );
buf ( n33161 , n33160 );
nand ( n4156 , n33156 , n33161 );
buf ( n33163 , n4156 );
buf ( n33164 , n33163 );
buf ( n33165 , n30846 );
buf ( n4160 , n33165 );
buf ( n33167 , n4160 );
not ( n4162 , n33167 );
buf ( n33169 , n516 );
buf ( n33170 , n495 );
xor ( n4165 , n33169 , n33170 );
buf ( n33172 , n4165 );
not ( n4170 , n33172 );
or ( n33174 , n4162 , n4170 );
buf ( n33175 , n495 );
buf ( n33176 , n496 );
xor ( n33177 , n33175 , n33176 );
buf ( n33178 , n33177 );
buf ( n33179 , n33178 );
buf ( n33180 , n496 );
not ( n33181 , n33180 );
buf ( n33182 , n497 );
nand ( n4183 , n33181 , n33182 );
buf ( n33184 , n4183 );
buf ( n33185 , n33184 );
buf ( n33186 , n497 );
not ( n33187 , n33186 );
buf ( n33188 , n496 );
nand ( n4189 , n33187 , n33188 );
buf ( n33190 , n4189 );
buf ( n33191 , n33190 );
and ( n4192 , n33179 , n33185 , n33191 );
buf ( n33193 , n4192 );
buf ( n33194 , n33193 );
not ( n33195 , n33194 );
buf ( n33196 , n33195 );
buf ( n33197 , n517 );
buf ( n33198 , n495 );
xor ( n4199 , n33197 , n33198 );
buf ( n33200 , n4199 );
buf ( n33201 , n33200 );
not ( n4202 , n33201 );
buf ( n33203 , n4202 );
or ( n33204 , n33196 , n33203 );
nand ( n4205 , n33174 , n33204 );
buf ( n33206 , n4205 );
xor ( n4207 , n33164 , n33206 );
buf ( n33208 , n518 );
buf ( n33209 , n493 );
xor ( n4210 , n33208 , n33209 );
buf ( n33211 , n4210 );
buf ( n33212 , n33211 );
not ( n4213 , n33212 );
not ( n4214 , n494 );
not ( n33215 , n2975 );
or ( n4216 , n4214 , n33215 );
nand ( n4217 , n2708 , n495 );
nand ( n4218 , n4216 , n4217 );
buf ( n33219 , n4218 );
not ( n4220 , n33219 );
or ( n4221 , n4213 , n4220 );
buf ( n33222 , n493 );
buf ( n33223 , n494 );
xor ( n4224 , n33222 , n33223 );
buf ( n33225 , n4224 );
buf ( n33226 , n33225 );
buf ( n33227 , n494 );
not ( n4228 , n33227 );
buf ( n33229 , n495 );
nand ( n4230 , n4228 , n33229 );
buf ( n33231 , n4230 );
buf ( n33232 , n33231 );
buf ( n33233 , n495 );
not ( n4234 , n33233 );
buf ( n33235 , n494 );
nand ( n33236 , n4234 , n33235 );
buf ( n33237 , n33236 );
buf ( n33238 , n33237 );
nand ( n4239 , n33226 , n33232 , n33238 );
buf ( n33240 , n4239 );
not ( n4241 , n33240 );
not ( n4242 , n4241 );
buf ( n33243 , n4242 );
xor ( n4244 , n493 , n519 );
buf ( n33245 , n4244 );
not ( n4249 , n33245 );
buf ( n33247 , n4249 );
buf ( n33248 , n33247 );
or ( n4252 , n33243 , n33248 );
nand ( n4253 , n4221 , n4252 );
buf ( n33251 , n4253 );
buf ( n33252 , n33251 );
and ( n4259 , n4207 , n33252 );
and ( n4260 , n33164 , n33206 );
or ( n33255 , n4259 , n4260 );
buf ( n33256 , n33255 );
buf ( n33257 , n33256 );
xor ( n4264 , n33147 , n33257 );
buf ( n33259 , n4264 );
buf ( n33260 , n33259 );
xor ( n4267 , n33107 , n33122 );
xor ( n4268 , n4267 , n33141 );
buf ( n33263 , n4268 );
buf ( n33264 , n33263 );
not ( n4271 , n4218 );
not ( n4272 , n4244 );
or ( n33267 , n4271 , n4272 );
xor ( n4274 , n520 , n493 );
nand ( n4275 , n4241 , n4274 );
nand ( n4276 , n33267 , n4275 );
buf ( n33271 , n4276 );
buf ( n33272 , n30912 );
buf ( n33273 , n514 );
buf ( n33274 , n499 );
xor ( n4281 , n33273 , n33274 );
buf ( n33276 , n4281 );
buf ( n33277 , n33276 );
not ( n4284 , n33277 );
buf ( n33279 , n4284 );
buf ( n33280 , n33279 );
or ( n33281 , n33272 , n33280 );
buf ( n33282 , n29543 );
buf ( n33283 , n513 );
buf ( n33284 , n499 );
xor ( n4291 , n33283 , n33284 );
buf ( n33286 , n4291 );
buf ( n33287 , n33286 );
nand ( n4294 , n33282 , n33287 );
buf ( n33289 , n4294 );
buf ( n33290 , n33289 );
nand ( n4297 , n33281 , n33290 );
buf ( n33292 , n4297 );
buf ( n33293 , n33292 );
xor ( n4300 , n33271 , n33293 );
buf ( n33295 , n520 );
buf ( n33296 , n494 );
or ( n33297 , n33295 , n33296 );
buf ( n33298 , n495 );
nand ( n4305 , n33297 , n33298 );
buf ( n33300 , n4305 );
buf ( n33301 , n33300 );
buf ( n33302 , n520 );
buf ( n33303 , n494 );
nand ( n4310 , n33302 , n33303 );
buf ( n33305 , n4310 );
buf ( n33306 , n33305 );
buf ( n33307 , n493 );
nand ( n4314 , n33301 , n33306 , n33307 );
buf ( n33309 , n4314 );
not ( n4316 , n33309 );
buf ( n33311 , n512 );
buf ( n33312 , n501 );
xor ( n4319 , n33311 , n33312 );
buf ( n33314 , n4319 );
not ( n4321 , n33314 );
not ( n4322 , n29640 );
or ( n4323 , n4321 , n4322 );
buf ( n33318 , n4118 );
buf ( n33319 , n29646 );
nand ( n4326 , n33318 , n33319 );
buf ( n33321 , n4326 );
nand ( n33322 , n4323 , n33321 );
not ( n33323 , n33322 );
or ( n33324 , n4316 , n33323 );
or ( n4331 , n33322 , n33309 );
nand ( n4332 , n33324 , n4331 );
buf ( n33327 , n4332 );
and ( n4334 , n4300 , n33327 );
and ( n4335 , n33271 , n33293 );
or ( n4336 , n4334 , n4335 );
buf ( n33331 , n4336 );
buf ( n33332 , n33331 );
xor ( n33333 , n33264 , n33332 );
xor ( n33334 , n33164 , n33206 );
xor ( n4344 , n33334 , n33252 );
buf ( n33336 , n4344 );
buf ( n33337 , n33336 );
and ( n4347 , n33333 , n33337 );
and ( n4348 , n33264 , n33332 );
or ( n4349 , n4347 , n4348 );
buf ( n33341 , n4349 );
buf ( n33342 , n33341 );
xor ( n33343 , n33260 , n33342 );
buf ( n33344 , n520 );
buf ( n33345 , n491 );
xor ( n4358 , n33344 , n33345 );
buf ( n33347 , n4358 );
buf ( n33348 , n33347 );
not ( n4361 , n33348 );
buf ( n33350 , n491 );
buf ( n33351 , n492 );
xnor ( n4364 , n33350 , n33351 );
buf ( n33353 , n4364 );
buf ( n33354 , n492 );
buf ( n33355 , n493 );
xor ( n33356 , n33354 , n33355 );
buf ( n33357 , n33356 );
nor ( n4370 , n33353 , n33357 );
buf ( n33359 , n4370 );
not ( n4372 , n33359 );
or ( n4373 , n4361 , n4372 );
buf ( n33362 , n33102 );
buf ( n33363 , n519 );
buf ( n33364 , n491 );
xor ( n4377 , n33363 , n33364 );
buf ( n33366 , n4377 );
buf ( n33367 , n33366 );
nand ( n4380 , n33362 , n33367 );
buf ( n33369 , n4380 );
buf ( n33370 , n33369 );
nand ( n4383 , n4373 , n33370 );
buf ( n33372 , n4383 );
buf ( n33373 , n33372 );
not ( n4386 , n33211 );
and ( n4387 , n33225 , n33237 , n33231 );
not ( n4388 , n4387 );
or ( n4389 , n4386 , n4388 );
buf ( n33378 , n494 );
buf ( n33379 , n495 );
xor ( n4392 , n33378 , n33379 );
buf ( n33381 , n4392 );
buf ( n33382 , n33381 );
buf ( n33383 , n517 );
buf ( n33384 , n493 );
xor ( n4397 , n33383 , n33384 );
buf ( n33386 , n4397 );
buf ( n33387 , n33386 );
nand ( n4400 , n33382 , n33387 );
buf ( n33389 , n4400 );
nand ( n4402 , n4389 , n33389 );
buf ( n33391 , n4402 );
xor ( n4404 , n33373 , n33391 );
buf ( n33393 , n512 );
buf ( n33394 , n499 );
xor ( n4407 , n33393 , n33394 );
buf ( n33396 , n4407 );
buf ( n33397 , n33396 );
not ( n4410 , n33397 );
buf ( n33399 , n30741 );
not ( n33400 , n33399 );
or ( n4413 , n4410 , n33400 );
buf ( n33402 , n511 );
buf ( n33403 , n499 );
xor ( n4416 , n33402 , n33403 );
buf ( n33405 , n4416 );
buf ( n33406 , n33405 );
buf ( n33407 , n29543 );
nand ( n4420 , n33406 , n33407 );
buf ( n33409 , n4420 );
buf ( n33410 , n33409 );
nand ( n4423 , n4413 , n33410 );
buf ( n33412 , n4423 );
buf ( n33413 , n33412 );
xor ( n4426 , n4404 , n33413 );
buf ( n33415 , n4426 );
buf ( n33416 , n33415 );
buf ( n33417 , n33134 );
not ( n4430 , n33417 );
buf ( n33419 , n29640 );
not ( n33420 , n33419 );
or ( n33421 , n4430 , n33420 );
buf ( n33422 , n29637 );
not ( n4435 , n33422 );
buf ( n33424 , n4435 );
buf ( n33425 , n33424 );
buf ( n33426 , n509 );
buf ( n33427 , n501 );
xor ( n4440 , n33426 , n33427 );
buf ( n33429 , n4440 );
buf ( n33430 , n33429 );
nand ( n33431 , n33425 , n33430 );
buf ( n33432 , n33431 );
buf ( n33433 , n33432 );
nand ( n4449 , n33421 , n33433 );
buf ( n33435 , n4449 );
buf ( n33436 , n33435 );
buf ( n33437 , n33172 );
not ( n4453 , n33437 );
buf ( n33439 , n33193 );
not ( n4458 , n33439 );
or ( n4459 , n4453 , n4458 );
xor ( n33442 , n515 , n495 );
nand ( n4461 , n30846 , n33442 );
buf ( n33444 , n4461 );
nand ( n4463 , n4459 , n33444 );
buf ( n33446 , n4463 );
buf ( n33447 , n33446 );
xor ( n4466 , n33436 , n33447 );
buf ( n33449 , n4109 );
not ( n4468 , n33449 );
buf ( n33451 , n30769 );
not ( n33452 , n33451 );
or ( n4471 , n4468 , n33452 );
buf ( n33454 , n1698 );
xor ( n4473 , n497 , n513 );
buf ( n33456 , n4473 );
nand ( n4475 , n33454 , n33456 );
buf ( n33458 , n4475 );
buf ( n33459 , n33458 );
nand ( n4478 , n4471 , n33459 );
buf ( n33461 , n4478 );
buf ( n33462 , n33461 );
xor ( n33463 , n4466 , n33462 );
buf ( n33464 , n33463 );
buf ( n33465 , n33464 );
xor ( n4484 , n33416 , n33465 );
buf ( n33467 , n33286 );
not ( n4486 , n33467 );
buf ( n33469 , n30741 );
not ( n4488 , n33469 );
or ( n4489 , n4486 , n4488 );
buf ( n33472 , n29543 );
buf ( n33473 , n33396 );
nand ( n4492 , n33472 , n33473 );
buf ( n33475 , n4492 );
buf ( n33476 , n33475 );
nand ( n33477 , n4489 , n33476 );
buf ( n33478 , n33477 );
buf ( n33479 , n33478 );
buf ( n33480 , n33322 );
buf ( n33481 , n33309 );
not ( n4500 , n33481 );
buf ( n33483 , n4500 );
buf ( n33484 , n33483 );
and ( n4503 , n33480 , n33484 );
buf ( n33486 , n4503 );
buf ( n33487 , n33486 );
xor ( n4506 , n33479 , n33487 );
buf ( n33489 , n510 );
buf ( n33490 , n503 );
xor ( n4509 , n33489 , n33490 );
buf ( n33492 , n4509 );
buf ( n33493 , n33492 );
not ( n4512 , n33493 );
buf ( n33495 , n29582 );
not ( n4514 , n33495 );
or ( n4515 , n4512 , n4514 );
buf ( n33498 , n33151 );
buf ( n33499 , n504 );
nand ( n4518 , n33498 , n33499 );
buf ( n33501 , n4518 );
buf ( n33502 , n33501 );
nand ( n4521 , n4515 , n33502 );
buf ( n33504 , n4521 );
buf ( n33505 , n33504 );
buf ( n33506 , n518 );
buf ( n33507 , n495 );
xor ( n4526 , n33506 , n33507 );
buf ( n33509 , n4526 );
buf ( n33510 , n33509 );
not ( n4529 , n33510 );
buf ( n33512 , n33193 );
not ( n4531 , n33512 );
or ( n4532 , n4529 , n4531 );
buf ( n33515 , n30846 );
buf ( n33516 , n33200 );
nand ( n4535 , n33515 , n33516 );
buf ( n33518 , n4535 );
buf ( n33519 , n33518 );
nand ( n4538 , n4532 , n33519 );
buf ( n33521 , n4538 );
buf ( n33522 , n33521 );
xor ( n4541 , n33505 , n33522 );
xor ( n4542 , n497 , n516 );
buf ( n33525 , n4542 );
not ( n4544 , n33525 );
buf ( n33527 , n30769 );
not ( n33528 , n33527 );
or ( n33529 , n4544 , n33528 );
buf ( n33530 , n1698 );
buf ( n33531 , n4102 );
nand ( n4550 , n33530 , n33531 );
buf ( n33533 , n4550 );
buf ( n33534 , n33533 );
nand ( n4553 , n33529 , n33534 );
buf ( n33536 , n4553 );
buf ( n33537 , n33536 );
and ( n4559 , n4541 , n33537 );
and ( n33539 , n33505 , n33522 );
or ( n4561 , n4559 , n33539 );
buf ( n33541 , n4561 );
buf ( n33542 , n33541 );
and ( n4564 , n4506 , n33542 );
and ( n4565 , n33479 , n33487 );
or ( n33545 , n4564 , n4565 );
buf ( n33546 , n33545 );
buf ( n33547 , n33546 );
xor ( n4572 , n4484 , n33547 );
buf ( n33549 , n4572 );
buf ( n33550 , n33549 );
xor ( n4575 , n33343 , n33550 );
buf ( n33552 , n4575 );
xor ( n4577 , n33479 , n33487 );
xor ( n4578 , n4577 , n33542 );
buf ( n33555 , n4578 );
buf ( n33556 , n33555 );
xor ( n4581 , n497 , n517 );
not ( n33558 , n4581 );
not ( n4583 , n30769 );
or ( n4584 , n33558 , n4583 );
buf ( n33561 , n1786 );
buf ( n33562 , n4542 );
nand ( n4587 , n33561 , n33562 );
buf ( n33564 , n4587 );
nand ( n4589 , n4584 , n33564 );
not ( n4590 , n4589 );
buf ( n33567 , n513 );
buf ( n33568 , n501 );
xor ( n4593 , n33567 , n33568 );
buf ( n33570 , n4593 );
not ( n4595 , n33570 );
not ( n4596 , n29640 );
or ( n4597 , n4595 , n4596 );
buf ( n33574 , n33314 );
buf ( n33575 , n33424 );
nand ( n4600 , n33574 , n33575 );
buf ( n33577 , n4600 );
nand ( n4602 , n4597 , n33577 );
not ( n4603 , n4602 );
buf ( n33580 , n33381 );
buf ( n33581 , n520 );
and ( n4606 , n33580 , n33581 );
buf ( n33583 , n4606 );
not ( n4608 , n33583 );
nand ( n4609 , n4603 , n4608 );
not ( n4610 , n4609 );
or ( n4611 , n4590 , n4610 );
nand ( n4612 , n33583 , n4602 );
nand ( n4613 , n4611 , n4612 );
not ( n4614 , n29734 );
and ( n4615 , n511 , n503 );
not ( n4616 , n511 );
and ( n4617 , n4616 , n956 );
nor ( n4618 , n4615 , n4617 );
not ( n4619 , n4618 );
or ( n4620 , n4614 , n4619 );
buf ( n33597 , n33492 );
buf ( n33598 , n504 );
nand ( n4623 , n33597 , n33598 );
buf ( n33600 , n4623 );
nand ( n4625 , n4620 , n33600 );
buf ( n33602 , n4625 );
buf ( n33603 , n519 );
buf ( n33604 , n495 );
xor ( n4629 , n33603 , n33604 );
buf ( n33606 , n4629 );
buf ( n33607 , n33606 );
not ( n4632 , n33607 );
buf ( n33609 , n33193 );
not ( n4634 , n33609 );
or ( n4635 , n4632 , n4634 );
buf ( n33612 , n30846 );
buf ( n33613 , n33509 );
nand ( n4638 , n33612 , n33613 );
buf ( n33615 , n4638 );
buf ( n33616 , n33615 );
nand ( n4641 , n4635 , n33616 );
buf ( n33618 , n4641 );
buf ( n33619 , n33618 );
xor ( n33620 , n33602 , n33619 );
buf ( n33621 , n30912 );
buf ( n33622 , n515 );
buf ( n33623 , n499 );
xor ( n4648 , n33622 , n33623 );
buf ( n33625 , n4648 );
buf ( n33626 , n33625 );
not ( n4651 , n33626 );
buf ( n33628 , n4651 );
buf ( n33629 , n33628 );
or ( n33630 , n33621 , n33629 );
buf ( n33631 , n29543 );
buf ( n33632 , n33276 );
nand ( n4657 , n33631 , n33632 );
buf ( n33634 , n4657 );
buf ( n33635 , n33634 );
nand ( n4660 , n33630 , n33635 );
buf ( n33637 , n4660 );
buf ( n33638 , n33637 );
and ( n4663 , n33620 , n33638 );
and ( n4664 , n33602 , n33619 );
or ( n4665 , n4663 , n4664 );
buf ( n33642 , n4665 );
xor ( n4667 , n4613 , n33642 );
xor ( n33644 , n33505 , n33522 );
xor ( n33645 , n33644 , n33537 );
buf ( n33646 , n33645 );
and ( n4671 , n4667 , n33646 );
and ( n4672 , n4613 , n33642 );
or ( n4673 , n4671 , n4672 );
buf ( n33650 , n4673 );
xor ( n4675 , n33556 , n33650 );
xor ( n4676 , n33264 , n33332 );
xor ( n33653 , n4676 , n33337 );
buf ( n33654 , n33653 );
buf ( n33655 , n33654 );
and ( n4683 , n4675 , n33655 );
and ( n4684 , n33556 , n33650 );
or ( n33658 , n4683 , n4684 );
buf ( n33659 , n33658 );
nor ( n4690 , n33552 , n33659 );
xor ( n4691 , n33556 , n33650 );
xor ( n4692 , n4691 , n33655 );
buf ( n33663 , n4692 );
xor ( n4694 , n33271 , n33293 );
xor ( n4695 , n4694 , n33327 );
buf ( n33666 , n4695 );
buf ( n33667 , n33666 );
xor ( n4698 , n4613 , n33642 );
xor ( n4699 , n4698 , n33646 );
buf ( n33670 , n4699 );
xor ( n4701 , n33667 , n33670 );
buf ( n33672 , n520 );
buf ( n33673 , n496 );
or ( n4704 , n33672 , n33673 );
buf ( n33675 , n497 );
nand ( n4706 , n4704 , n33675 );
buf ( n33677 , n4706 );
buf ( n33678 , n33677 );
buf ( n33679 , n520 );
buf ( n33680 , n496 );
nand ( n4711 , n33679 , n33680 );
buf ( n33682 , n4711 );
buf ( n33683 , n33682 );
buf ( n33684 , n495 );
and ( n4715 , n33678 , n33683 , n33684 );
buf ( n33686 , n4715 );
buf ( n33687 , n33686 );
buf ( n33688 , n30887 );
not ( n4719 , n33688 );
buf ( n33690 , n29640 );
not ( n4721 , n33690 );
or ( n33692 , n4719 , n4721 );
buf ( n33693 , n29649 );
buf ( n33694 , n33570 );
nand ( n4725 , n33693 , n33694 );
buf ( n33696 , n4725 );
buf ( n33697 , n33696 );
nand ( n4728 , n33692 , n33697 );
buf ( n33699 , n4728 );
buf ( n33700 , n33699 );
and ( n4731 , n33687 , n33700 );
buf ( n33702 , n4731 );
and ( n4733 , n33583 , n4602 );
not ( n4734 , n33583 );
and ( n4735 , n4734 , n4603 );
nor ( n4736 , n4733 , n4735 );
and ( n4737 , n4736 , n4589 );
not ( n4738 , n4736 );
not ( n4739 , n4589 );
and ( n33710 , n4738 , n4739 );
nor ( n4741 , n4737 , n33710 );
xor ( n4742 , n33702 , n4741 );
buf ( n33713 , n30834 );
not ( n4744 , n33713 );
buf ( n33715 , n29582 );
not ( n4746 , n33715 );
or ( n4747 , n4744 , n4746 );
buf ( n33718 , n4618 );
buf ( n33719 , n504 );
nand ( n4750 , n33718 , n33719 );
buf ( n33721 , n4750 );
buf ( n33722 , n33721 );
nand ( n4753 , n4747 , n33722 );
buf ( n33724 , n4753 );
buf ( n33725 , n33724 );
buf ( n33726 , n1788 );
not ( n4757 , n33726 );
buf ( n33728 , n30769 );
not ( n4759 , n33728 );
or ( n4760 , n4757 , n4759 );
buf ( n33731 , n1786 );
buf ( n33732 , n4581 );
nand ( n4763 , n33731 , n33732 );
buf ( n33734 , n4763 );
buf ( n33735 , n33734 );
nand ( n4766 , n4760 , n33735 );
buf ( n33737 , n4766 );
buf ( n33738 , n33737 );
xor ( n4769 , n33725 , n33738 );
buf ( n33740 , n495 );
buf ( n33741 , n520 );
and ( n4772 , n33740 , n33741 );
not ( n4773 , n33740 );
buf ( n33744 , n29690 );
and ( n33745 , n4773 , n33744 );
nor ( n4776 , n4772 , n33745 );
buf ( n33747 , n4776 );
buf ( n33748 , n33747 );
not ( n33749 , n33748 );
buf ( n33750 , n33178 );
buf ( n33751 , n33184 );
buf ( n33752 , n33190 );
and ( n4783 , n33750 , n33751 , n33752 );
buf ( n33754 , n4783 );
buf ( n33755 , n33754 );
buf ( n4786 , n33755 );
buf ( n33757 , n4786 );
buf ( n33758 , n33757 );
not ( n4789 , n33758 );
or ( n4790 , n33749 , n4789 );
buf ( n33761 , n33606 );
buf ( n33762 , n33167 );
nand ( n4793 , n33761 , n33762 );
buf ( n33764 , n4793 );
buf ( n33765 , n33764 );
nand ( n4796 , n4790 , n33765 );
buf ( n33767 , n4796 );
buf ( n33768 , n33767 );
and ( n33769 , n4769 , n33768 );
and ( n4800 , n33725 , n33738 );
or ( n4801 , n33769 , n4800 );
buf ( n33772 , n4801 );
and ( n4803 , n4742 , n33772 );
and ( n4804 , n33702 , n4741 );
or ( n4805 , n4803 , n4804 );
buf ( n33776 , n4805 );
and ( n4810 , n4701 , n33776 );
and ( n33778 , n33667 , n33670 );
or ( n4812 , n4810 , n33778 );
buf ( n33780 , n4812 );
nor ( n33781 , n33663 , n33780 );
nor ( n4818 , n4690 , n33781 );
not ( n4819 , n4818 );
xor ( n33784 , n33602 , n33619 );
xor ( n4821 , n33784 , n33638 );
buf ( n33786 , n4821 );
buf ( n33787 , n33786 );
buf ( n33788 , n30904 );
not ( n4825 , n33788 );
buf ( n33790 , n29535 );
not ( n4827 , n33790 );
or ( n4828 , n4825 , n4827 );
buf ( n33793 , n29543 );
buf ( n33794 , n33625 );
nand ( n4831 , n33793 , n33794 );
buf ( n33796 , n4831 );
buf ( n33797 , n33796 );
nand ( n4834 , n4828 , n33797 );
buf ( n33799 , n4834 );
buf ( n33800 , n33799 );
xor ( n4837 , n33687 , n33700 );
buf ( n33802 , n4837 );
buf ( n33803 , n33802 );
xor ( n4840 , n33800 , n33803 );
xor ( n4841 , n30842 , n30851 );
and ( n4842 , n4841 , n30867 );
and ( n4843 , n30842 , n30851 );
or ( n4844 , n4842 , n4843 );
buf ( n33809 , n4844 );
buf ( n33810 , n33809 );
and ( n4847 , n4840 , n33810 );
and ( n4848 , n33800 , n33803 );
or ( n4849 , n4847 , n4848 );
buf ( n33814 , n4849 );
buf ( n33815 , n33814 );
xor ( n4852 , n33787 , n33815 );
xor ( n4853 , n33702 , n4741 );
xor ( n4854 , n4853 , n33772 );
buf ( n33819 , n4854 );
xor ( n4856 , n4852 , n33819 );
buf ( n33821 , n4856 );
xor ( n4858 , n30894 , n30899 );
and ( n4859 , n4858 , n30918 );
and ( n4860 , n30894 , n30899 );
or ( n4861 , n4859 , n4860 );
buf ( n33826 , n4861 );
buf ( n33827 , n33826 );
xor ( n4864 , n33725 , n33738 );
xor ( n33829 , n4864 , n33768 );
buf ( n33830 , n33829 );
buf ( n33831 , n33830 );
xor ( n4868 , n33827 , n33831 );
xor ( n4869 , n33800 , n33803 );
xor ( n4870 , n4869 , n33810 );
buf ( n33835 , n4870 );
buf ( n33836 , n33835 );
and ( n4873 , n4868 , n33836 );
and ( n4874 , n33827 , n33831 );
or ( n4875 , n4873 , n4874 );
buf ( n33840 , n4875 );
nor ( n4877 , n33821 , n33840 );
not ( n4878 , n4877 );
xor ( n4879 , n33667 , n33670 );
xor ( n33844 , n4879 , n33776 );
buf ( n33845 , n33844 );
not ( n4882 , n33845 );
xor ( n4883 , n33787 , n33815 );
and ( n4884 , n4883 , n33819 );
and ( n33849 , n33787 , n33815 );
or ( n4886 , n4884 , n33849 );
buf ( n33851 , n4886 );
not ( n4888 , n33851 );
nand ( n4889 , n4882 , n4888 );
xor ( n33854 , n33827 , n33831 );
xor ( n4891 , n33854 , n33836 );
buf ( n33856 , n4891 );
not ( n4893 , n33856 );
xor ( n4894 , n30870 , n30876 );
and ( n4895 , n4894 , n30921 );
and ( n4896 , n30870 , n30876 );
or ( n4897 , n4895 , n4896 );
buf ( n33862 , n4897 );
not ( n4899 , n33862 );
nand ( n4900 , n4893 , n4899 );
not ( n4901 , n4900 );
nor ( n4902 , n4901 , n1857 );
nand ( n4903 , n4878 , n4889 , n1753 , n4902 );
nand ( n4904 , n33856 , n33862 );
nand ( n4905 , n4904 , n1859 );
nand ( n4906 , n4900 , n4905 );
nor ( n4907 , n4906 , n4877 );
nand ( n4908 , n33845 , n33851 );
nand ( n4909 , n33821 , n33840 );
nand ( n4910 , n4908 , n4909 );
or ( n4911 , n4907 , n4910 );
nand ( n4912 , n4911 , n4889 );
nand ( n4913 , n4903 , n4912 );
not ( n4914 , n4913 );
or ( n4915 , n4819 , n4914 );
nand ( n4916 , n33663 , n33780 );
or ( n4917 , n4690 , n4916 );
nand ( n4918 , n33552 , n33659 );
nand ( n4919 , n4917 , n4918 );
not ( n4920 , n4919 );
nand ( n4921 , n4915 , n4920 );
xor ( n4922 , n33416 , n33465 );
and ( n4923 , n4922 , n33547 );
and ( n4924 , n33416 , n33465 );
or ( n4925 , n4923 , n4924 );
buf ( n33890 , n4925 );
buf ( n33891 , n33890 );
xor ( n4928 , n490 , n491 );
and ( n4929 , n4928 , n520 );
not ( n4930 , n504 );
buf ( n33895 , n506 );
buf ( n33896 , n503 );
xor ( n4933 , n33895 , n33896 );
buf ( n33898 , n4933 );
not ( n4935 , n33898 );
or ( n33900 , n4930 , n4935 );
nand ( n33901 , n29734 , n4056 );
nand ( n33902 , n33900 , n33901 );
xor ( n4939 , n4929 , n33902 );
buf ( n33904 , n508 );
buf ( n33905 , n501 );
xor ( n4942 , n33904 , n33905 );
buf ( n33907 , n4942 );
not ( n4944 , n33907 );
not ( n33909 , n33424 );
or ( n4949 , n4944 , n33909 );
buf ( n33911 , n29637 );
buf ( n33912 , n29638 );
nand ( n4952 , n33911 , n33912 );
buf ( n33914 , n4952 );
not ( n4957 , n33914 );
nand ( n4958 , n4957 , n33429 );
nand ( n4959 , n4949 , n4958 );
xor ( n4960 , n4939 , n4959 );
buf ( n33919 , n4960 );
xor ( n4962 , n33373 , n33391 );
and ( n4963 , n4962 , n33413 );
and ( n4964 , n33373 , n33391 );
or ( n4965 , n4963 , n4964 );
buf ( n33924 , n4965 );
buf ( n33925 , n33924 );
xor ( n4968 , n33919 , n33925 );
xor ( n4969 , n33436 , n33447 );
and ( n4970 , n4969 , n33462 );
and ( n4971 , n33436 , n33447 );
or ( n4972 , n4970 , n4971 );
buf ( n33931 , n4972 );
buf ( n33932 , n33931 );
xor ( n4975 , n4968 , n33932 );
buf ( n33934 , n4975 );
buf ( n33935 , n33934 );
xor ( n4978 , n33891 , n33935 );
buf ( n33937 , n33069 );
buf ( n33938 , n33086 );
and ( n4981 , n33937 , n33938 );
buf ( n33940 , n4981 );
buf ( n33941 , n33940 );
buf ( n33942 , n33386 );
not ( n4985 , n33942 );
buf ( n33944 , n4241 );
not ( n4987 , n33944 );
or ( n4988 , n4985 , n4987 );
buf ( n33947 , n516 );
buf ( n33948 , n493 );
xor ( n4991 , n33947 , n33948 );
buf ( n33950 , n4991 );
buf ( n33951 , n33950 );
buf ( n33952 , n4218 );
nand ( n4995 , n33951 , n33952 );
buf ( n33954 , n4995 );
buf ( n33955 , n33954 );
nand ( n4998 , n4988 , n33955 );
buf ( n33957 , n4998 );
buf ( n33958 , n33957 );
xor ( n5001 , n33941 , n33958 );
buf ( n33960 , n33366 );
not ( n5003 , n33960 );
buf ( n33962 , n4370 );
not ( n5005 , n33962 );
buf ( n33964 , n5005 );
buf ( n33965 , n33964 );
not ( n5008 , n33965 );
buf ( n33967 , n5008 );
buf ( n33968 , n33967 );
not ( n5011 , n33968 );
or ( n5012 , n5003 , n5011 );
buf ( n33971 , n33102 );
buf ( n5014 , n33971 );
buf ( n33973 , n5014 );
buf ( n33974 , n33973 );
buf ( n33975 , n518 );
buf ( n33976 , n491 );
xor ( n5019 , n33975 , n33976 );
buf ( n33978 , n5019 );
buf ( n33979 , n33978 );
nand ( n5022 , n33974 , n33979 );
buf ( n33981 , n5022 );
buf ( n33982 , n33981 );
nand ( n33983 , n5012 , n33982 );
buf ( n33984 , n33983 );
buf ( n33985 , n33984 );
xor ( n5028 , n5001 , n33985 );
buf ( n33987 , n5028 );
buf ( n33988 , n33987 );
not ( n5031 , n4473 );
not ( n5032 , n30769 );
or ( n5033 , n5031 , n5032 );
buf ( n33992 , n29604 );
xor ( n5035 , n497 , n512 );
buf ( n33994 , n5035 );
nand ( n5037 , n33992 , n33994 );
buf ( n33996 , n5037 );
nand ( n5039 , n5033 , n33996 );
not ( n5040 , n5039 );
not ( n5041 , n33405 );
not ( n5042 , n29535 );
or ( n5043 , n5041 , n5042 );
buf ( n34002 , n29542 );
buf ( n34003 , n510 );
buf ( n34004 , n499 );
xor ( n5047 , n34003 , n34004 );
buf ( n34006 , n5047 );
buf ( n34007 , n34006 );
nand ( n5050 , n34002 , n34007 );
buf ( n34009 , n5050 );
nand ( n5052 , n5043 , n34009 );
not ( n5053 , n5052 );
and ( n5054 , n5040 , n5053 );
and ( n5055 , n5039 , n5052 );
nor ( n5056 , n5054 , n5055 );
nand ( n5057 , n33754 , n33442 );
not ( n5058 , n5057 );
not ( n5059 , n30846 );
buf ( n34018 , n514 );
buf ( n34019 , n495 );
xnor ( n5062 , n34018 , n34019 );
buf ( n34021 , n5062 );
nor ( n5064 , n5059 , n34021 );
nor ( n5065 , n5058 , n5064 );
buf ( n5066 , n5065 );
not ( n5067 , n5066 );
and ( n5068 , n5056 , n5067 );
not ( n5069 , n5056 );
and ( n5070 , n5069 , n5066 );
nor ( n5071 , n5068 , n5070 );
buf ( n34030 , n5071 );
xor ( n5073 , n33988 , n34030 );
xor ( n5074 , n33098 , n33146 );
and ( n5075 , n5074 , n33257 );
and ( n5076 , n33098 , n33146 );
or ( n5077 , n5075 , n5076 );
buf ( n34036 , n5077 );
buf ( n34037 , n34036 );
xor ( n5080 , n5073 , n34037 );
buf ( n34039 , n5080 );
buf ( n34040 , n34039 );
xor ( n5083 , n4978 , n34040 );
buf ( n34042 , n5083 );
xor ( n34043 , n33260 , n33342 );
and ( n34044 , n34043 , n33550 );
and ( n34045 , n33260 , n33342 );
or ( n5088 , n34044 , n34045 );
buf ( n34047 , n5088 );
nand ( n5090 , n34042 , n34047 );
not ( n5091 , n34042 );
not ( n5092 , n34047 );
nand ( n5093 , n5091 , n5092 );
nand ( n34052 , n5090 , n5093 );
and ( n5098 , n4921 , n34052 , n29519 );
nor ( n34054 , n4040 , n5098 );
not ( n5100 , n4038 );
nand ( n5101 , n5100 , n455 );
not ( n34057 , n5101 );
not ( n5106 , n3800 );
and ( n5107 , n34057 , n5106 );
not ( n5108 , n4921 );
nor ( n5109 , n34052 , n455 );
and ( n5110 , n5108 , n5109 );
nor ( n5111 , n5107 , n5110 );
buf ( n34064 , n541 );
not ( n5113 , n34064 );
buf ( n34066 , n5113 );
nand ( n5115 , n34054 , n5111 , n34066 );
buf ( n34068 , n5115 );
buf ( n5117 , n34068 );
buf ( n34070 , n5117 );
not ( n5119 , n4921 );
not ( n5120 , n5093 );
or ( n5121 , n5119 , n5120 );
nand ( n34074 , n5121 , n5090 );
not ( n5123 , n34074 );
buf ( n34076 , n5065 );
not ( n5125 , n34076 );
not ( n5126 , n5052 );
buf ( n34079 , n5126 );
not ( n5128 , n34079 );
or ( n5129 , n5125 , n5128 );
buf ( n34082 , n5039 );
nand ( n5131 , n5129 , n34082 );
buf ( n34084 , n5131 );
buf ( n34085 , n34084 );
buf ( n34086 , n5052 );
buf ( n34087 , n34021 );
not ( n5136 , n34087 );
buf ( n34089 , n30846 );
nand ( n5138 , n5136 , n34089 );
buf ( n34091 , n5138 );
nand ( n5140 , n34091 , n5057 );
buf ( n34093 , n5140 );
nand ( n5142 , n34086 , n34093 );
buf ( n34095 , n5142 );
buf ( n34096 , n34095 );
nand ( n5145 , n34085 , n34096 );
buf ( n34098 , n5145 );
buf ( n34099 , n34098 );
buf ( n34100 , n33907 );
not ( n5149 , n34100 );
buf ( n34102 , n33914 );
not ( n5151 , n34102 );
buf ( n34104 , n5151 );
buf ( n34105 , n34104 );
not ( n5154 , n34105 );
or ( n5155 , n5149 , n5154 );
buf ( n34108 , n33424 );
xor ( n5157 , n501 , n507 );
buf ( n34110 , n5157 );
nand ( n5159 , n34108 , n34110 );
buf ( n34112 , n5159 );
buf ( n34113 , n34112 );
nand ( n5162 , n5155 , n34113 );
buf ( n34115 , n5162 );
xor ( n5164 , n489 , n520 );
buf ( n34117 , n5164 );
not ( n5166 , n34117 );
not ( n5167 , n491 );
not ( n5168 , n490 );
nand ( n5169 , n5167 , n5168 , n489 );
not ( n5170 , n489 );
nand ( n5171 , n5170 , n491 , n490 );
nand ( n5172 , n5169 , n5171 );
buf ( n34125 , n5172 );
not ( n5174 , n34125 );
or ( n5175 , n5166 , n5174 );
and ( n5176 , n489 , n519 );
not ( n5177 , n489 );
not ( n5178 , n519 );
and ( n5179 , n5177 , n5178 );
nor ( n5180 , n5176 , n5179 );
nand ( n5181 , n4928 , n5180 );
buf ( n34134 , n5181 );
nand ( n5183 , n5175 , n34134 );
buf ( n34136 , n5183 );
xor ( n5185 , n34115 , n34136 );
buf ( n34138 , n5185 );
buf ( n34139 , n5035 );
not ( n5188 , n34139 );
buf ( n34141 , n1691 );
not ( n5190 , n34141 );
or ( n5191 , n5188 , n5190 );
buf ( n34144 , n29604 );
xor ( n5193 , n497 , n511 );
buf ( n34146 , n5193 );
nand ( n5195 , n34144 , n34146 );
buf ( n34148 , n5195 );
buf ( n34149 , n34148 );
nand ( n5198 , n5191 , n34149 );
buf ( n34151 , n5198 );
buf ( n34152 , n34151 );
and ( n5201 , n34138 , n34152 );
not ( n5202 , n34138 );
buf ( n34155 , n34151 );
not ( n5204 , n34155 );
buf ( n34157 , n5204 );
buf ( n34158 , n34157 );
and ( n5207 , n5202 , n34158 );
nor ( n5208 , n5201 , n5207 );
buf ( n34161 , n5208 );
buf ( n34162 , n34161 );
xor ( n5211 , n34099 , n34162 );
not ( n5212 , n33950 );
not ( n5213 , n4387 );
or ( n5214 , n5212 , n5213 );
buf ( n34167 , n515 );
buf ( n34168 , n493 );
xor ( n5217 , n34167 , n34168 );
buf ( n34170 , n5217 );
buf ( n34171 , n34170 );
buf ( n34172 , n33381 );
nand ( n5221 , n34171 , n34172 );
buf ( n34174 , n5221 );
nand ( n5223 , n5214 , n34174 );
buf ( n34176 , n5223 );
buf ( n34177 , n34006 );
not ( n5226 , n34177 );
buf ( n34179 , n30741 );
not ( n5228 , n34179 );
or ( n34181 , n5226 , n5228 );
buf ( n5230 , n29527 );
buf ( n34183 , n5230 );
xor ( n5232 , n499 , n509 );
buf ( n34185 , n5232 );
nand ( n5234 , n34183 , n34185 );
buf ( n34187 , n5234 );
buf ( n34188 , n34187 );
nand ( n5237 , n34181 , n34188 );
buf ( n34190 , n5237 );
buf ( n34191 , n34190 );
xor ( n5240 , n34176 , n34191 );
xor ( n5241 , n495 , n513 );
buf ( n34194 , n5241 );
not ( n5243 , n34194 );
buf ( n34196 , n33167 );
not ( n34197 , n34196 );
or ( n34198 , n5243 , n34197 );
buf ( n34199 , n33196 );
buf ( n34200 , n34021 );
or ( n5249 , n34199 , n34200 );
nand ( n5250 , n34198 , n5249 );
buf ( n34203 , n5250 );
buf ( n34204 , n34203 );
xor ( n34205 , n5240 , n34204 );
buf ( n34206 , n34205 );
buf ( n34207 , n34206 );
xor ( n5259 , n5211 , n34207 );
buf ( n34209 , n5259 );
buf ( n34210 , n34209 );
xor ( n5265 , n33988 , n34030 );
and ( n5266 , n5265 , n34037 );
and ( n5267 , n33988 , n34030 );
or ( n5268 , n5266 , n5267 );
buf ( n34215 , n5268 );
buf ( n34216 , n34215 );
xor ( n34217 , n34210 , n34216 );
xor ( n5272 , n33941 , n33958 );
and ( n5273 , n5272 , n33985 );
and ( n5274 , n33941 , n33958 );
or ( n5275 , n5273 , n5274 );
buf ( n34222 , n5275 );
buf ( n34223 , n34222 );
buf ( n34224 , n33978 );
not ( n5279 , n34224 );
buf ( n34226 , n33967 );
not ( n5281 , n34226 );
or ( n5282 , n5279 , n5281 );
buf ( n34229 , n33973 );
xor ( n5284 , n491 , n517 );
buf ( n34231 , n5284 );
nand ( n5286 , n34229 , n34231 );
buf ( n34233 , n5286 );
buf ( n34234 , n34233 );
nand ( n5289 , n5282 , n34234 );
buf ( n34236 , n5289 );
buf ( n34237 , n34236 );
buf ( n34238 , n520 );
buf ( n34239 , n490 );
or ( n5294 , n34238 , n34239 );
buf ( n34241 , n491 );
nand ( n5296 , n5294 , n34241 );
buf ( n34243 , n5296 );
buf ( n34244 , n34243 );
buf ( n34245 , n520 );
buf ( n34246 , n490 );
nand ( n5301 , n34245 , n34246 );
buf ( n34248 , n5301 );
buf ( n34249 , n34248 );
buf ( n34250 , n489 );
and ( n5305 , n34244 , n34249 , n34250 );
buf ( n34252 , n5305 );
buf ( n34253 , n34252 );
buf ( n34254 , n33898 );
not ( n5309 , n34254 );
buf ( n34256 , n29582 );
not ( n5311 , n34256 );
or ( n5312 , n5309 , n5311 );
xor ( n5313 , n503 , n505 );
buf ( n34260 , n5313 );
buf ( n34261 , n504 );
nand ( n5316 , n34260 , n34261 );
buf ( n34263 , n5316 );
buf ( n34264 , n34263 );
nand ( n5319 , n5312 , n34264 );
buf ( n34266 , n5319 );
buf ( n34267 , n34266 );
xor ( n5322 , n34253 , n34267 );
buf ( n34269 , n5322 );
buf ( n34270 , n34269 );
xor ( n5325 , n34237 , n34270 );
xor ( n5326 , n4929 , n33902 );
and ( n5327 , n5326 , n4959 );
and ( n5328 , n4929 , n33902 );
or ( n5329 , n5327 , n5328 );
buf ( n34276 , n5329 );
xor ( n5331 , n5325 , n34276 );
buf ( n34278 , n5331 );
buf ( n34279 , n34278 );
xor ( n5334 , n34223 , n34279 );
xor ( n5335 , n33919 , n33925 );
and ( n5336 , n5335 , n33932 );
and ( n5337 , n33919 , n33925 );
or ( n5338 , n5336 , n5337 );
buf ( n34285 , n5338 );
buf ( n34286 , n34285 );
xor ( n5341 , n5334 , n34286 );
buf ( n34288 , n5341 );
buf ( n34289 , n34288 );
xor ( n5344 , n34217 , n34289 );
buf ( n34291 , n5344 );
xor ( n34292 , n33891 , n33935 );
and ( n5347 , n34292 , n34040 );
and ( n5348 , n33891 , n33935 );
or ( n5349 , n5347 , n5348 );
buf ( n34296 , n5349 );
nor ( n5351 , n34291 , n34296 );
not ( n5352 , n5351 );
nand ( n5353 , n34291 , n34296 );
nand ( n5354 , n5352 , n5353 );
not ( n5355 , n5354 );
nand ( n5356 , n5355 , n29519 );
not ( n5357 , n5356 );
and ( n5358 , n5123 , n5357 );
not ( n5359 , n33042 );
not ( n5360 , n3800 );
or ( n5361 , n5359 , n5360 );
nand ( n34308 , n5361 , n4037 );
or ( n5363 , n3996 , n32985 );
nand ( n5364 , n5363 , n4010 );
nand ( n5365 , n32985 , n3996 );
nand ( n34312 , n5364 , n5365 );
buf ( n34313 , n34312 );
not ( n5368 , n3511 );
not ( n5369 , n3915 );
or ( n5370 , n5368 , n5369 );
nand ( n5371 , n882 , n493 );
not ( n5372 , n5371 );
nand ( n5373 , n2831 , n2704 );
not ( n5374 , n5373 );
or ( n5375 , n5372 , n5374 );
nand ( n5376 , n5375 , n3113 );
nand ( n5377 , n5370 , n5376 );
buf ( n34324 , n5377 );
not ( n5379 , n495 );
not ( n5380 , n3597 );
or ( n5381 , n5379 , n5380 );
buf ( n34328 , n1403 );
buf ( n34329 , n31784 );
nand ( n5384 , n34328 , n34329 );
buf ( n34331 , n5384 );
nand ( n5386 , n5381 , n34331 );
not ( n5387 , n5386 );
not ( n5388 , n2725 );
or ( n5389 , n5387 , n5388 );
nand ( n5390 , n3989 , n31812 );
nand ( n5391 , n5389 , n5390 );
buf ( n34338 , n5391 );
xor ( n5393 , n34324 , n34338 );
not ( n5394 , n799 );
not ( n5395 , n3971 );
or ( n5396 , n5394 , n5395 );
not ( n5397 , n499 );
not ( n5398 , n29492 );
or ( n5399 , n5397 , n5398 );
buf ( n34346 , n29493 );
buf ( n34347 , n29901 );
nand ( n5402 , n34346 , n34347 );
buf ( n34349 , n5402 );
nand ( n5404 , n5399 , n34349 );
nand ( n5405 , n5404 , n29884 );
nand ( n5406 , n5396 , n5405 );
buf ( n34353 , n5406 );
xor ( n5408 , n5393 , n34353 );
buf ( n34355 , n5408 );
buf ( n34356 , n34355 );
xor ( n5411 , n34313 , n34356 );
buf ( n34358 , n489 );
buf ( n34359 , n490 );
xnor ( n34360 , n34358 , n34359 );
buf ( n34361 , n34360 );
not ( n5416 , n34361 );
nand ( n5417 , n5416 , n3833 );
not ( n5418 , n5417 );
not ( n5419 , n5418 );
not ( n5420 , n489 );
not ( n5421 , n32849 );
or ( n34368 , n5420 , n5421 );
buf ( n34369 , n489 );
not ( n34370 , n34369 );
buf ( n34371 , n29939 );
nand ( n5429 , n34370 , n34371 );
buf ( n34373 , n5429 );
nand ( n5434 , n34368 , n34373 );
not ( n5435 , n5434 );
or ( n5436 , n5419 , n5435 );
not ( n5437 , n489 );
and ( n5438 , n29912 , n5437 );
not ( n5439 , n29912 );
and ( n5440 , n5439 , n489 );
nor ( n5441 , n5438 , n5440 );
nand ( n5442 , n5441 , n3832 );
nand ( n5443 , n5436 , n5442 );
buf ( n34384 , n5443 );
buf ( n34385 , n3072 );
not ( n5446 , n34385 );
and ( n5447 , n29501 , n497 );
not ( n5448 , n29501 );
and ( n5449 , n5448 , n30599 );
nor ( n5450 , n5447 , n5449 );
buf ( n34391 , n5450 );
not ( n5452 , n34391 );
or ( n5453 , n5446 , n5452 );
buf ( n34394 , n497 );
not ( n5455 , n34394 );
buf ( n34396 , n2678 );
not ( n5457 , n34396 );
or ( n5458 , n5455 , n5457 );
and ( n5459 , n456 , n463 );
not ( n5460 , n456 );
and ( n5461 , n5460 , n479 );
or ( n5462 , n5459 , n5461 );
buf ( n34403 , n5462 );
buf ( n34404 , n30599 );
nand ( n5465 , n34403 , n34404 );
buf ( n34406 , n5465 );
buf ( n34407 , n34406 );
nand ( n5468 , n5458 , n34407 );
buf ( n34409 , n5468 );
buf ( n34410 , n34409 );
buf ( n34411 , n910 );
nand ( n5472 , n34410 , n34411 );
buf ( n34413 , n5472 );
buf ( n34414 , n34413 );
nand ( n34415 , n5453 , n34414 );
buf ( n34416 , n34415 );
buf ( n34417 , n34416 );
xor ( n5478 , n34384 , n34417 );
buf ( n34419 , n30078 );
not ( n5480 , n34419 );
buf ( n34421 , n3873 );
not ( n5482 , n34421 );
or ( n5483 , n5480 , n5482 );
buf ( n34424 , n501 );
not ( n5485 , n34424 );
buf ( n34426 , n32467 );
not ( n5487 , n34426 );
or ( n5488 , n5485 , n5487 );
buf ( n34429 , n3434 );
buf ( n34430 , n984 );
nand ( n5491 , n34429 , n34430 );
buf ( n34432 , n5491 );
buf ( n34433 , n34432 );
nand ( n5494 , n5488 , n34433 );
buf ( n34435 , n5494 );
buf ( n34436 , n34435 );
buf ( n34437 , n1010 );
nand ( n5498 , n34436 , n34437 );
buf ( n34439 , n5498 );
buf ( n34440 , n34439 );
nand ( n34441 , n5483 , n34440 );
buf ( n34442 , n34441 );
buf ( n34443 , n34442 );
xor ( n5504 , n5478 , n34443 );
buf ( n34445 , n5504 );
buf ( n34446 , n34445 );
xor ( n5507 , n5411 , n34446 );
buf ( n34448 , n5507 );
buf ( n34449 , n34448 );
xor ( n5510 , n32970 , n4023 );
and ( n5511 , n5510 , n33035 );
and ( n5512 , n32970 , n4023 );
or ( n5513 , n5511 , n5512 );
buf ( n34454 , n5513 );
xor ( n5515 , n34449 , n34454 );
xor ( n5516 , n32935 , n32964 );
and ( n5517 , n5516 , n32968 );
and ( n5518 , n32935 , n32964 );
or ( n5519 , n5517 , n5518 );
buf ( n34460 , n5519 );
buf ( n34461 , n34460 );
not ( n5522 , n32949 );
buf ( n34463 , n3948 );
buf ( n5524 , n34463 );
buf ( n34465 , n5524 );
not ( n5526 , n34465 );
or ( n5527 , n5522 , n5526 );
and ( n5528 , n456 , n469 );
not ( n5529 , n456 );
and ( n5530 , n5529 , n485 );
nor ( n5531 , n5528 , n5530 );
and ( n5532 , n5531 , n5167 );
not ( n5533 , n5531 );
and ( n5534 , n5533 , n491 );
nor ( n5535 , n5532 , n5534 );
nand ( n5536 , n5535 , n3043 );
nand ( n5537 , n5527 , n5536 );
and ( n5538 , n29957 , n490 );
not ( n5539 , n489 );
nor ( n5540 , n5538 , n5539 );
not ( n5541 , n5168 );
not ( n5542 , n30592 );
or ( n5543 , n5541 , n5542 );
nand ( n5544 , n5543 , n491 );
nand ( n5545 , n5540 , n5544 );
not ( n5546 , n5545 );
buf ( n34487 , n504 );
not ( n5548 , n34487 );
buf ( n34489 , n503 );
not ( n5550 , n34489 );
and ( n5551 , n456 , n457 );
not ( n5552 , n456 );
and ( n5553 , n5552 , n473 );
nor ( n5554 , n5551 , n5553 );
buf ( n34495 , n5554 );
not ( n5556 , n34495 );
or ( n5557 , n5550 , n5556 );
and ( n5558 , n456 , n457 );
not ( n5559 , n456 );
and ( n5560 , n5559 , n473 );
nor ( n5561 , n5558 , n5560 );
not ( n5562 , n5561 );
buf ( n34503 , n5562 );
buf ( n34504 , n29987 );
nand ( n5565 , n34503 , n34504 );
buf ( n34506 , n5565 );
buf ( n34507 , n34506 );
nand ( n5568 , n5557 , n34507 );
buf ( n34509 , n5568 );
buf ( n34510 , n34509 );
not ( n5571 , n34510 );
or ( n5572 , n5548 , n5571 );
nand ( n5573 , n3857 , n29969 );
buf ( n34514 , n5573 );
nand ( n5575 , n5572 , n34514 );
buf ( n34516 , n5575 );
xor ( n5577 , n5546 , n34516 );
xor ( n5578 , n5537 , n5577 );
xor ( n5579 , n32853 , n32880 );
and ( n5580 , n5579 , n32899 );
and ( n5581 , n32853 , n32880 );
or ( n5582 , n5580 , n5581 );
buf ( n34523 , n5582 );
xor ( n34524 , n5578 , n34523 );
buf ( n34525 , n34524 );
xor ( n5586 , n34461 , n34525 );
buf ( n34527 , n32901 );
not ( n5588 , n34527 );
buf ( n34529 , n3820 );
not ( n34530 , n34529 );
buf ( n34531 , n34530 );
buf ( n34532 , n34531 );
not ( n5596 , n34532 );
or ( n5597 , n5588 , n5596 );
buf ( n34535 , n32901 );
not ( n5602 , n34535 );
buf ( n34537 , n5602 );
buf ( n34538 , n34537 );
not ( n5605 , n34538 );
buf ( n34540 , n3820 );
not ( n5607 , n34540 );
or ( n5608 , n5605 , n5607 );
buf ( n34543 , n3812 );
nand ( n5610 , n5608 , n34543 );
buf ( n34545 , n5610 );
buf ( n34546 , n34545 );
nand ( n5613 , n5597 , n34546 );
buf ( n34548 , n5613 );
buf ( n34549 , n34548 );
xor ( n5616 , n5586 , n34549 );
buf ( n34551 , n5616 );
buf ( n34552 , n34551 );
xor ( n5619 , n5515 , n34552 );
buf ( n34554 , n5619 );
xor ( n5621 , n3897 , n3901 );
and ( n5622 , n5621 , n4030 );
and ( n5623 , n3897 , n3901 );
or ( n5624 , n5622 , n5623 );
nor ( n5625 , n34554 , n5624 );
not ( n5626 , n5625 );
nand ( n5627 , n34554 , n5624 );
nand ( n34562 , n5626 , n5627 );
and ( n5629 , n34562 , n455 );
and ( n5630 , n34308 , n5629 );
nor ( n5631 , n5358 , n5630 );
not ( n5632 , n5631 );
not ( n5633 , n34308 );
not ( n5634 , n34562 );
nand ( n5635 , n5634 , n455 );
not ( n5636 , n5635 );
and ( n5637 , n5633 , n5636 );
not ( n5638 , n540 );
and ( n5639 , n5354 , n29519 );
nand ( n5640 , n34074 , n5639 );
nand ( n5641 , n5638 , n5640 );
nor ( n5642 , n5637 , n5641 );
not ( n5643 , n5642 );
or ( n5644 , n5632 , n5643 );
not ( n5645 , n5629 );
and ( n5646 , n5645 , n34308 );
not ( n5647 , n5635 );
nor ( n5648 , n34308 , n5647 );
nor ( n5649 , n5646 , n5648 );
not ( n5650 , n5356 );
not ( n5651 , n5650 );
not ( n5652 , n34074 );
not ( n34587 , n5652 );
or ( n5654 , n5651 , n34587 );
nand ( n5655 , n5654 , n5640 );
or ( n5656 , n5649 , n5655 );
nand ( n5657 , n5656 , n540 );
nand ( n5658 , n5644 , n5657 );
nand ( n5659 , n34070 , n5658 );
buf ( n5660 , n5659 );
nor ( n5661 , n5658 , n34070 );
not ( n5662 , n5661 );
nand ( n5663 , n5660 , n5662 );
nor ( n5664 , n5663 , n2618 );
not ( n34599 , n5664 );
buf ( n34600 , n545 );
not ( n5667 , n34600 );
not ( n5668 , n29519 );
not ( n5669 , n4877 );
buf ( n5670 , n4909 );
nand ( n5671 , n5669 , n5670 );
not ( n5672 , n5671 );
not ( n5673 , n4902 );
not ( n5674 , n1753 );
or ( n5675 , n5673 , n5674 );
nand ( n5676 , n5675 , n4906 );
not ( n5677 , n5676 );
or ( n5678 , n5672 , n5677 );
or ( n5679 , n5676 , n5671 );
nand ( n5680 , n5678 , n5679 );
not ( n5681 , n5680 );
or ( n5682 , n5668 , n5681 );
not ( n5683 , n3778 );
not ( n5684 , n1875 );
or ( n5685 , n5683 , n5684 );
buf ( n5686 , n3784 );
nand ( n5687 , n5685 , n5686 );
nand ( n5688 , n3761 , n3787 );
not ( n5689 , n5688 );
and ( n5690 , n5687 , n5689 );
not ( n5691 , n5687 );
and ( n5692 , n5691 , n5688 );
nor ( n5693 , n5690 , n5692 );
nand ( n5694 , n5693 , n455 );
nand ( n5695 , n5682 , n5694 );
buf ( n34630 , n5695 );
not ( n5697 , n34630 );
or ( n5698 , n5667 , n5697 );
buf ( n34633 , n5695 );
not ( n5700 , n34633 );
buf ( n34635 , n5700 );
buf ( n34636 , n34635 );
buf ( n34637 , n545 );
not ( n5704 , n34637 );
buf ( n34639 , n5704 );
buf ( n34640 , n34639 );
nand ( n5707 , n34636 , n34640 );
buf ( n34642 , n5707 );
buf ( n34643 , n34642 );
nand ( n5710 , n5698 , n34643 );
buf ( n34645 , n5710 );
buf ( n34646 , n34645 );
not ( n5713 , n2029 );
not ( n5714 , n5713 );
not ( n5715 , n1875 );
or ( n5716 , n5714 , n5715 );
buf ( n5717 , n2026 );
nand ( n5718 , n5716 , n5717 );
nand ( n5719 , n3780 , n3776 );
not ( n5720 , n5719 );
and ( n5721 , n5718 , n5720 );
not ( n5722 , n5718 );
and ( n5723 , n5722 , n5719 );
nor ( n5724 , n5721 , n5723 );
nand ( n5725 , n5724 , n455 );
not ( n5726 , n1858 );
not ( n5727 , n1753 );
or ( n5728 , n5726 , n5727 );
nand ( n5729 , n5728 , n1859 );
nand ( n5730 , n4900 , n4904 );
not ( n5731 , n5730 );
and ( n5732 , n5729 , n5731 );
not ( n5733 , n5729 );
and ( n5734 , n5733 , n5730 );
nor ( n5735 , n5732 , n5734 );
nand ( n5736 , n5735 , n29519 );
nand ( n5737 , n5725 , n5736 );
buf ( n34672 , n5737 );
not ( n5739 , n34672 );
buf ( n34674 , n546 );
not ( n5741 , n34674 );
buf ( n34676 , n5741 );
buf ( n34677 , n34676 );
nand ( n5744 , n5739 , n34677 );
buf ( n34679 , n5744 );
buf ( n34680 , n34679 );
or ( n5747 , n34646 , n34680 );
buf ( n34682 , n5747 );
buf ( n34683 , n34682 );
not ( n5753 , n546 );
not ( n34685 , n5737 );
or ( n5755 , n5753 , n34685 );
nand ( n5756 , n5725 , n5736 , n34676 );
nand ( n34688 , n5755 , n5756 );
buf ( n34689 , n34688 );
not ( n5762 , n2037 );
nand ( n5763 , n5762 , n30816 );
buf ( n34692 , n5763 );
and ( n5765 , n34689 , n34692 );
buf ( n34694 , n5765 );
buf ( n34695 , n34694 );
and ( n5768 , n34683 , n34695 );
buf ( n34697 , n34645 );
buf ( n34698 , n34679 );
and ( n5771 , n34697 , n34698 );
buf ( n34700 , n5771 );
buf ( n34701 , n34700 );
nor ( n5774 , n5768 , n34701 );
buf ( n34703 , n5774 );
buf ( n34704 , n34645 );
buf ( n34705 , n34679 );
or ( n5778 , n34704 , n34705 );
buf ( n34707 , n5778 );
buf ( n34708 , n34707 );
not ( n5781 , n30816 );
not ( n5782 , n31103 );
or ( n5783 , n5781 , n5782 );
nand ( n5784 , n5783 , n31109 );
not ( n5785 , n5784 );
not ( n5786 , n2053 );
not ( n5787 , n5786 );
or ( n5788 , n5785 , n5787 );
nand ( n5789 , n5788 , n2052 );
buf ( n34718 , n5789 );
not ( n5791 , n34688 );
not ( n5792 , n5763 );
nand ( n5793 , n5791 , n5792 );
buf ( n34722 , n5793 );
nand ( n5795 , n34708 , n34718 , n34722 );
buf ( n34724 , n5795 );
buf ( n34725 , n30813 );
buf ( n34726 , n2050 );
nor ( n5799 , n34725 , n34726 );
buf ( n34728 , n5799 );
nand ( n5801 , n34707 , n34728 , n5793 );
nand ( n5802 , n34703 , n34724 , n5801 );
not ( n5803 , n5802 );
not ( n5804 , n541 );
nand ( n5805 , n5111 , n34054 );
not ( n5806 , n5805 );
or ( n5807 , n5804 , n5806 );
nand ( n5808 , n5807 , n5115 );
buf ( n34737 , n5808 );
not ( n5810 , n34737 );
not ( n5811 , n3794 );
nand ( n5812 , n5811 , n3797 );
not ( n5813 , n5812 );
nand ( n5814 , n5813 , n455 );
not ( n5815 , n5814 );
or ( n5816 , n3288 , n3397 );
not ( n5817 , n5816 );
not ( n5818 , n3791 );
or ( n5819 , n5817 , n5818 );
nand ( n5820 , n5819 , n3795 );
not ( n5821 , n5820 );
nand ( n5822 , n5815 , n5821 );
not ( n5823 , n33781 );
not ( n5824 , n5823 );
not ( n5825 , n4913 );
or ( n5826 , n5824 , n5825 );
nand ( n5827 , n5826 , n4916 );
not ( n5828 , n4690 );
nand ( n5829 , n5828 , n4918 );
not ( n5830 , n5829 );
nand ( n5831 , n5830 , n29519 );
nor ( n5832 , n5827 , n5831 );
not ( n5833 , n5832 );
and ( n5834 , n5812 , n455 );
nand ( n5835 , n5820 , n5834 );
nand ( n5836 , n5827 , n5829 , n29519 );
nand ( n5837 , n5822 , n5833 , n5835 , n5836 );
buf ( n34766 , n5837 );
not ( n5839 , n34766 );
buf ( n34768 , n5839 );
buf ( n34769 , n34768 );
buf ( n34770 , n542 );
not ( n5843 , n34770 );
buf ( n34772 , n5843 );
buf ( n34773 , n34772 );
nand ( n5846 , n34769 , n34773 );
buf ( n34775 , n5846 );
buf ( n34776 , n34775 );
not ( n5849 , n34776 );
buf ( n34778 , n5849 );
buf ( n34779 , n34778 );
nand ( n5852 , n5810 , n34779 );
buf ( n34781 , n5852 );
buf ( n34782 , n34781 );
buf ( n34783 , n542 );
not ( n5856 , n34783 );
buf ( n34785 , n5837 );
not ( n5858 , n34785 );
or ( n5859 , n5856 , n5858 );
buf ( n34788 , n34768 );
buf ( n34789 , n34772 );
nand ( n5862 , n34788 , n34789 );
buf ( n34791 , n5862 );
buf ( n34792 , n34791 );
nand ( n5865 , n5859 , n34792 );
buf ( n34794 , n5865 );
buf ( n34795 , n34794 );
not ( n5868 , n29519 );
nand ( n5869 , n5823 , n4916 );
not ( n5870 , n5869 );
not ( n5871 , n4913 );
or ( n5872 , n5870 , n5871 );
or ( n5873 , n5869 , n4913 );
nand ( n5874 , n5872 , n5873 );
not ( n5875 , n5874 );
or ( n5876 , n5868 , n5875 );
nand ( n5877 , n5816 , n3795 );
not ( n5878 , n5877 );
not ( n5879 , n3791 );
or ( n5880 , n5878 , n5879 );
nand ( n5881 , n3779 , n3790 );
or ( n5882 , n5881 , n5877 );
nand ( n5883 , n5880 , n5882 );
nand ( n5884 , n5883 , n455 );
nand ( n5885 , n5876 , n5884 );
not ( n5886 , n5885 );
buf ( n34815 , n5886 );
buf ( n34816 , n543 );
not ( n5889 , n34816 );
buf ( n34818 , n5889 );
buf ( n34819 , n34818 );
nand ( n5892 , n34815 , n34819 );
buf ( n34821 , n5892 );
buf ( n34822 , n34821 );
or ( n5895 , n34795 , n34822 );
buf ( n34824 , n5895 );
buf ( n34825 , n34824 );
not ( n5898 , n34818 );
not ( n5899 , n5886 );
or ( n5900 , n5898 , n5899 );
buf ( n34829 , n34818 );
not ( n5902 , n34829 );
buf ( n34831 , n5885 );
nand ( n5904 , n5902 , n34831 );
buf ( n34833 , n5904 );
nand ( n5906 , n5900 , n34833 );
not ( n5907 , n3761 );
not ( n5908 , n5687 );
or ( n5909 , n5907 , n5908 );
nand ( n5910 , n5909 , n3787 );
or ( n5911 , n3674 , n32757 );
nand ( n5912 , n5911 , n3786 );
not ( n5913 , n5912 );
nand ( n5914 , n5913 , n455 );
nor ( n5915 , n5910 , n5914 );
not ( n5916 , n5915 );
nand ( n34845 , n5910 , n5912 , n455 );
not ( n34846 , n5669 );
not ( n5919 , n5676 );
or ( n5920 , n34846 , n5919 );
nand ( n34849 , n5920 , n5670 );
nand ( n5925 , n4889 , n4908 );
not ( n34851 , n5925 );
nand ( n5927 , n34851 , n29519 );
nor ( n5928 , n34849 , n5927 );
not ( n34854 , n5928 );
and ( n5933 , n5925 , n29519 );
nand ( n5934 , n34849 , n5933 );
nand ( n5935 , n5916 , n34845 , n34854 , n5934 );
buf ( n34858 , n5935 );
not ( n5937 , n34858 );
buf ( n34860 , n5937 );
buf ( n34861 , n544 );
not ( n5940 , n34861 );
buf ( n34863 , n5940 );
nand ( n5942 , n34860 , n34863 );
nor ( n5943 , n5906 , n5942 );
buf ( n34866 , n544 );
not ( n5945 , n34866 );
buf ( n34868 , n5935 );
not ( n5947 , n34868 );
or ( n34870 , n5945 , n5947 );
buf ( n34871 , n34860 );
buf ( n34872 , n34863 );
nand ( n5951 , n34871 , n34872 );
buf ( n34874 , n5951 );
buf ( n34875 , n34874 );
nand ( n5954 , n34870 , n34875 );
buf ( n34877 , n5954 );
buf ( n34878 , n34877 );
buf ( n34879 , n34642 );
buf ( n5958 , n34879 );
buf ( n34881 , n5958 );
buf ( n34882 , n34881 );
nor ( n5961 , n34878 , n34882 );
buf ( n34884 , n5961 );
nor ( n5963 , n5943 , n34884 );
buf ( n34886 , n5963 );
and ( n5965 , n34782 , n34825 , n34886 );
buf ( n34888 , n5965 );
not ( n5967 , n34888 );
or ( n5968 , n5803 , n5967 );
nand ( n5969 , n34824 , n34781 );
not ( n5970 , n5969 );
not ( n5971 , n5942 );
nand ( n5972 , n5886 , n34818 );
nand ( n5973 , n5971 , n34833 , n5972 );
not ( n5974 , n5973 );
buf ( n34897 , n34877 );
buf ( n34898 , n34881 );
and ( n5977 , n34897 , n34898 );
buf ( n34900 , n5977 );
not ( n5979 , n34900 );
or ( n5980 , n5974 , n5979 );
nand ( n5981 , n5906 , n5942 );
nand ( n5982 , n5980 , n5981 );
and ( n5983 , n5970 , n5982 );
buf ( n34906 , n34794 );
buf ( n34907 , n34821 );
nand ( n5986 , n34906 , n34907 );
buf ( n34909 , n5986 );
buf ( n34910 , n34909 );
not ( n5989 , n34910 );
buf ( n34912 , n5989 );
not ( n5991 , n34912 );
not ( n5992 , n34781 );
or ( n5993 , n5991 , n5992 );
buf ( n34916 , n5808 );
buf ( n5995 , n34916 );
buf ( n34918 , n5995 );
buf ( n34919 , n34918 );
buf ( n34920 , n34775 );
nand ( n5999 , n34919 , n34920 );
buf ( n34922 , n5999 );
nand ( n6001 , n5993 , n34922 );
nor ( n6002 , n5983 , n6001 );
nand ( n34925 , n5968 , n6002 );
buf ( n6004 , n34925 );
not ( n6005 , n6004 );
not ( n6006 , n6005 );
or ( n6007 , n34599 , n6006 );
not ( n6008 , n5663 );
nor ( n6009 , n6008 , n2618 );
and ( n6010 , n6009 , n6004 );
buf ( n34933 , n463 );
buf ( n34934 , n527 );
buf ( n34935 , n552 );
and ( n6014 , n34934 , n34935 );
buf ( n34937 , n6014 );
buf ( n34938 , n34937 );
xor ( n6017 , n34933 , n34938 );
buf ( n34940 , n6017 );
buf ( n34941 , n34940 );
buf ( n34942 , n464 );
buf ( n34943 , n528 );
buf ( n34944 , n552 );
and ( n6023 , n34943 , n34944 );
buf ( n34946 , n6023 );
buf ( n34947 , n34946 );
and ( n6026 , n34942 , n34947 );
buf ( n34949 , n6026 );
buf ( n34950 , n34949 );
xor ( n6029 , n34941 , n34950 );
buf ( n34952 , n531 );
buf ( n34953 , n549 );
and ( n6032 , n34952 , n34953 );
buf ( n34955 , n6032 );
buf ( n34956 , n34955 );
buf ( n34957 , n536 );
buf ( n34958 , n544 );
and ( n6037 , n34957 , n34958 );
buf ( n34960 , n6037 );
buf ( n34961 , n34960 );
xor ( n6040 , n34956 , n34961 );
buf ( n34963 , n529 );
buf ( n34964 , n551 );
and ( n6043 , n34963 , n34964 );
buf ( n34966 , n6043 );
buf ( n34967 , n34966 );
and ( n6046 , n6040 , n34967 );
and ( n6047 , n34956 , n34961 );
or ( n6048 , n6046 , n6047 );
buf ( n34971 , n6048 );
buf ( n34972 , n34971 );
and ( n6051 , n6029 , n34972 );
and ( n6052 , n34941 , n34950 );
or ( n6053 , n6051 , n6052 );
buf ( n34976 , n6053 );
buf ( n34977 , n34976 );
buf ( n34978 , n531 );
buf ( n34979 , n547 );
and ( n6058 , n34978 , n34979 );
buf ( n34981 , n6058 );
buf ( n34982 , n34981 );
buf ( n34983 , n462 );
buf ( n34984 , n526 );
buf ( n34985 , n552 );
and ( n6064 , n34984 , n34985 );
buf ( n34987 , n6064 );
buf ( n34988 , n34987 );
xor ( n6067 , n34983 , n34988 );
buf ( n34990 , n6067 );
buf ( n34991 , n34990 );
xor ( n6070 , n34982 , n34991 );
and ( n6071 , n34933 , n34938 );
buf ( n34994 , n6071 );
buf ( n34995 , n34994 );
xor ( n6074 , n6070 , n34995 );
buf ( n34997 , n6074 );
buf ( n34998 , n34997 );
xor ( n34999 , n34977 , n34998 );
buf ( n35000 , n528 );
buf ( n35001 , n551 );
and ( n6080 , n35000 , n35001 );
buf ( n35003 , n6080 );
buf ( n35004 , n35003 );
buf ( n35005 , n531 );
buf ( n35006 , n548 );
and ( n6088 , n35005 , n35006 );
buf ( n35008 , n6088 );
buf ( n35009 , n35008 );
xor ( n6094 , n35004 , n35009 );
buf ( n35011 , n532 );
buf ( n35012 , n547 );
and ( n6097 , n35011 , n35012 );
buf ( n35014 , n6097 );
buf ( n35015 , n35014 );
and ( n6100 , n6094 , n35015 );
and ( n6101 , n35004 , n35009 );
or ( n6102 , n6100 , n6101 );
buf ( n35019 , n6102 );
buf ( n35020 , n35019 );
buf ( n35021 , n529 );
buf ( n35022 , n550 );
and ( n6107 , n35021 , n35022 );
buf ( n35024 , n6107 );
buf ( n35025 , n35024 );
buf ( n35026 , n533 );
buf ( n35027 , n546 );
and ( n6112 , n35026 , n35027 );
buf ( n35029 , n6112 );
buf ( n35030 , n35029 );
xor ( n6115 , n35025 , n35030 );
buf ( n35032 , n534 );
buf ( n35033 , n545 );
and ( n6118 , n35032 , n35033 );
buf ( n35035 , n6118 );
buf ( n35036 , n35035 );
and ( n6121 , n6115 , n35036 );
and ( n6122 , n35025 , n35030 );
or ( n6123 , n6121 , n6122 );
buf ( n35040 , n6123 );
buf ( n35041 , n35040 );
xor ( n6126 , n35020 , n35041 );
buf ( n35043 , n530 );
buf ( n35044 , n549 );
and ( n6129 , n35043 , n35044 );
buf ( n35046 , n6129 );
buf ( n35047 , n35046 );
buf ( n35048 , n535 );
buf ( n35049 , n544 );
and ( n6134 , n35048 , n35049 );
buf ( n35051 , n6134 );
buf ( n35052 , n35051 );
xor ( n6137 , n35047 , n35052 );
buf ( n35054 , n536 );
buf ( n35055 , n543 );
and ( n6140 , n35054 , n35055 );
buf ( n35057 , n6140 );
buf ( n35058 , n35057 );
and ( n6143 , n6137 , n35058 );
and ( n35060 , n35047 , n35052 );
or ( n6145 , n6143 , n35060 );
buf ( n35062 , n6145 );
buf ( n35063 , n35062 );
xor ( n6148 , n6126 , n35063 );
buf ( n35065 , n6148 );
buf ( n35066 , n35065 );
xor ( n6151 , n34999 , n35066 );
buf ( n35068 , n6151 );
buf ( n35069 , n35068 );
and ( n6154 , n31601 , n31606 );
buf ( n35071 , n6154 );
buf ( n35072 , n35071 );
xor ( n6157 , n31545 , n31550 );
and ( n6158 , n6157 , n31556 );
and ( n6159 , n31545 , n31550 );
or ( n6160 , n6158 , n6159 );
buf ( n35077 , n6160 );
buf ( n35078 , n35077 );
xor ( n6163 , n35072 , n35078 );
xor ( n6164 , n31574 , n31579 );
and ( n6165 , n6164 , n31585 );
and ( n35082 , n31574 , n31579 );
or ( n6167 , n6165 , n35082 );
buf ( n35084 , n6167 );
buf ( n35085 , n35084 );
and ( n6170 , n6163 , n35085 );
and ( n6171 , n35072 , n35078 );
or ( n6172 , n6170 , n6171 );
buf ( n35089 , n6172 );
buf ( n35090 , n35089 );
buf ( n35091 , n530 );
buf ( n35092 , n550 );
and ( n6177 , n35091 , n35092 );
buf ( n35094 , n6177 );
buf ( n35095 , n35094 );
buf ( n35096 , n534 );
buf ( n35097 , n546 );
and ( n6182 , n35096 , n35097 );
buf ( n35099 , n6182 );
buf ( n35100 , n35099 );
xor ( n6185 , n35095 , n35100 );
buf ( n35102 , n535 );
buf ( n35103 , n545 );
and ( n6188 , n35102 , n35103 );
buf ( n35105 , n6188 );
buf ( n35106 , n35105 );
and ( n6191 , n6185 , n35106 );
and ( n6192 , n35095 , n35100 );
or ( n6193 , n6191 , n6192 );
buf ( n35110 , n6193 );
buf ( n35111 , n35110 );
xor ( n6196 , n35025 , n35030 );
xor ( n6197 , n6196 , n35036 );
buf ( n35114 , n6197 );
buf ( n35115 , n35114 );
xor ( n6200 , n35111 , n35115 );
xor ( n6201 , n35004 , n35009 );
xor ( n6202 , n6201 , n35015 );
buf ( n35119 , n6202 );
buf ( n35120 , n35119 );
xor ( n6205 , n6200 , n35120 );
buf ( n35122 , n6205 );
buf ( n35123 , n35122 );
xor ( n6208 , n35090 , n35123 );
xor ( n6209 , n35095 , n35100 );
xor ( n6210 , n6209 , n35106 );
buf ( n35127 , n6210 );
buf ( n35128 , n35127 );
xor ( n6213 , n34956 , n34961 );
xor ( n6214 , n6213 , n34967 );
buf ( n35131 , n6214 );
buf ( n35132 , n35131 );
xor ( n6217 , n35128 , n35132 );
xor ( n6218 , n31600 , n31609 );
and ( n6219 , n6218 , n31613 );
and ( n6220 , n31600 , n31609 );
or ( n6221 , n6219 , n6220 );
buf ( n35138 , n6221 );
buf ( n35139 , n35138 );
and ( n6224 , n6217 , n35139 );
and ( n6225 , n35128 , n35132 );
or ( n6226 , n6224 , n6225 );
buf ( n35143 , n6226 );
buf ( n35144 , n35143 );
and ( n6229 , n6208 , n35144 );
and ( n6230 , n35090 , n35123 );
or ( n6231 , n6229 , n6230 );
buf ( n35148 , n6231 );
buf ( n35149 , n35148 );
xor ( n6234 , n35069 , n35149 );
xor ( n6235 , n35111 , n35115 );
and ( n6236 , n6235 , n35120 );
and ( n6237 , n35111 , n35115 );
or ( n6238 , n6236 , n6237 );
buf ( n35155 , n6238 );
buf ( n35156 , n35155 );
buf ( n35157 , n527 );
buf ( n35158 , n551 );
and ( n35159 , n35157 , n35158 );
buf ( n35160 , n35159 );
buf ( n35161 , n35160 );
buf ( n35162 , n530 );
buf ( n35163 , n548 );
and ( n35164 , n35162 , n35163 );
buf ( n35165 , n35164 );
buf ( n35166 , n35165 );
xor ( n6257 , n35161 , n35166 );
buf ( n35168 , n536 );
buf ( n35169 , n542 );
and ( n6260 , n35168 , n35169 );
buf ( n35171 , n6260 );
buf ( n35172 , n35171 );
xor ( n6263 , n6257 , n35172 );
buf ( n35174 , n6263 );
buf ( n35175 , n35174 );
buf ( n35176 , n529 );
buf ( n35177 , n549 );
and ( n6268 , n35176 , n35177 );
buf ( n35179 , n6268 );
buf ( n35180 , n35179 );
buf ( n35181 , n534 );
buf ( n35182 , n544 );
and ( n6273 , n35181 , n35182 );
buf ( n35184 , n6273 );
buf ( n35185 , n35184 );
xor ( n6276 , n35180 , n35185 );
buf ( n35187 , n535 );
buf ( n35188 , n543 );
and ( n6279 , n35187 , n35188 );
buf ( n35190 , n6279 );
buf ( n35191 , n35190 );
xor ( n6282 , n6276 , n35191 );
buf ( n35193 , n6282 );
buf ( n35194 , n35193 );
xor ( n6285 , n35175 , n35194 );
buf ( n35196 , n528 );
buf ( n35197 , n550 );
and ( n6288 , n35196 , n35197 );
buf ( n35199 , n6288 );
buf ( n35200 , n35199 );
buf ( n35201 , n532 );
buf ( n35202 , n546 );
and ( n6293 , n35201 , n35202 );
buf ( n35204 , n6293 );
buf ( n35205 , n35204 );
xor ( n6296 , n35200 , n35205 );
buf ( n35207 , n533 );
buf ( n35208 , n545 );
and ( n6299 , n35207 , n35208 );
buf ( n35210 , n6299 );
buf ( n35211 , n35210 );
xor ( n6302 , n6296 , n35211 );
buf ( n35213 , n6302 );
buf ( n35214 , n35213 );
xor ( n6305 , n6285 , n35214 );
buf ( n35216 , n6305 );
buf ( n35217 , n35216 );
xor ( n6308 , n35156 , n35217 );
xor ( n6309 , n35047 , n35052 );
xor ( n6310 , n6309 , n35058 );
buf ( n35221 , n6310 );
buf ( n35222 , n35221 );
buf ( n35223 , n532 );
buf ( n35224 , n548 );
and ( n6315 , n35223 , n35224 );
buf ( n35226 , n6315 );
buf ( n35227 , n35226 );
buf ( n35228 , n533 );
buf ( n35229 , n547 );
and ( n6320 , n35228 , n35229 );
buf ( n35231 , n6320 );
buf ( n35232 , n35231 );
xor ( n6323 , n35227 , n35232 );
xor ( n6324 , n34942 , n34947 );
buf ( n35235 , n6324 );
buf ( n35236 , n35235 );
and ( n6327 , n6323 , n35236 );
and ( n6328 , n35227 , n35232 );
or ( n6329 , n6327 , n6328 );
buf ( n35240 , n6329 );
buf ( n35241 , n35240 );
xor ( n6332 , n35222 , n35241 );
xor ( n6333 , n34941 , n34950 );
xor ( n6334 , n6333 , n34972 );
buf ( n35245 , n6334 );
buf ( n35246 , n35245 );
and ( n6337 , n6332 , n35246 );
and ( n6338 , n35222 , n35241 );
or ( n6339 , n6337 , n6338 );
buf ( n35250 , n6339 );
buf ( n35251 , n35250 );
xor ( n6342 , n6308 , n35251 );
buf ( n35253 , n6342 );
buf ( n35254 , n35253 );
xor ( n6345 , n6234 , n35254 );
buf ( n35256 , n6345 );
xor ( n6347 , n35222 , n35241 );
xor ( n6348 , n6347 , n35246 );
buf ( n35259 , n6348 );
buf ( n35260 , n35259 );
xor ( n6351 , n35227 , n35232 );
xor ( n6352 , n6351 , n35236 );
buf ( n35263 , n6352 );
buf ( n35264 , n35263 );
xor ( n6355 , n35072 , n35078 );
xor ( n6356 , n6355 , n35085 );
buf ( n35267 , n6356 );
buf ( n35268 , n35267 );
xor ( n6359 , n35264 , n35268 );
xor ( n6360 , n31533 , n31539 );
and ( n6361 , n6360 , n31559 );
and ( n6362 , n31533 , n31539 );
or ( n6363 , n6361 , n6362 );
buf ( n35274 , n6363 );
buf ( n35275 , n35274 );
and ( n6366 , n6359 , n35275 );
and ( n6367 , n35264 , n35268 );
or ( n6368 , n6366 , n6367 );
buf ( n35279 , n6368 );
buf ( n35280 , n35279 );
xor ( n6371 , n35260 , n35280 );
xor ( n6372 , n35090 , n35123 );
xor ( n6373 , n6372 , n35144 );
buf ( n35284 , n6373 );
buf ( n35285 , n35284 );
and ( n6376 , n6371 , n35285 );
and ( n6377 , n35260 , n35280 );
or ( n6378 , n6376 , n6377 );
buf ( n35289 , n6378 );
or ( n6380 , n35256 , n35289 );
not ( n6381 , n6380 );
xor ( n6382 , n35069 , n35149 );
and ( n6383 , n6382 , n35254 );
and ( n6384 , n35069 , n35149 );
or ( n6385 , n6383 , n6384 );
buf ( n35296 , n6385 );
xor ( n6387 , n35020 , n35041 );
and ( n6388 , n6387 , n35063 );
and ( n6389 , n35020 , n35041 );
or ( n6390 , n6388 , n6389 );
buf ( n35301 , n6390 );
buf ( n35302 , n35301 );
xor ( n35303 , n35175 , n35194 );
and ( n6394 , n35303 , n35214 );
and ( n6395 , n35175 , n35194 );
or ( n35306 , n6394 , n6395 );
buf ( n35307 , n35306 );
buf ( n35308 , n35307 );
xor ( n6402 , n35302 , n35308 );
and ( n6403 , n34983 , n34988 );
buf ( n35311 , n6403 );
buf ( n35312 , n35311 );
xor ( n6409 , n35180 , n35185 );
and ( n6410 , n6409 , n35191 );
and ( n6411 , n35180 , n35185 );
or ( n6412 , n6410 , n6411 );
buf ( n35317 , n6412 );
buf ( n35318 , n35317 );
xor ( n6415 , n35312 , n35318 );
xor ( n6416 , n35161 , n35166 );
and ( n6417 , n6416 , n35172 );
and ( n6418 , n35161 , n35166 );
or ( n6419 , n6417 , n6418 );
buf ( n35324 , n6419 );
buf ( n35325 , n35324 );
xor ( n6422 , n6415 , n35325 );
buf ( n35327 , n6422 );
buf ( n35328 , n35327 );
xor ( n6425 , n6402 , n35328 );
buf ( n35330 , n6425 );
buf ( n35331 , n35330 );
xor ( n6428 , n35156 , n35217 );
and ( n6429 , n6428 , n35251 );
and ( n6430 , n35156 , n35217 );
or ( n6431 , n6429 , n6430 );
buf ( n35336 , n6431 );
buf ( n35337 , n35336 );
xor ( n6434 , n35331 , n35337 );
xor ( n6435 , n35200 , n35205 );
and ( n6436 , n6435 , n35211 );
and ( n6437 , n35200 , n35205 );
or ( n6438 , n6436 , n6437 );
buf ( n35343 , n6438 );
buf ( n35344 , n35343 );
buf ( n35345 , n526 );
buf ( n35346 , n551 );
and ( n6443 , n35345 , n35346 );
buf ( n35348 , n6443 );
buf ( n35349 , n35348 );
buf ( n35350 , n529 );
buf ( n35351 , n548 );
and ( n6448 , n35350 , n35351 );
buf ( n35353 , n6448 );
buf ( n35354 , n35353 );
xor ( n6451 , n35349 , n35354 );
buf ( n35356 , n535 );
buf ( n35357 , n542 );
and ( n6454 , n35356 , n35357 );
buf ( n35359 , n6454 );
buf ( n35360 , n35359 );
xor ( n6457 , n6451 , n35360 );
buf ( n35362 , n6457 );
buf ( n35363 , n35362 );
xor ( n6460 , n35344 , n35363 );
buf ( n35365 , n528 );
buf ( n35366 , n549 );
and ( n6463 , n35365 , n35366 );
buf ( n35368 , n6463 );
buf ( n35369 , n35368 );
buf ( n35370 , n533 );
buf ( n35371 , n544 );
and ( n6468 , n35370 , n35371 );
buf ( n35373 , n6468 );
buf ( n35374 , n35373 );
xor ( n6471 , n35369 , n35374 );
buf ( n35376 , n534 );
buf ( n35377 , n543 );
and ( n6474 , n35376 , n35377 );
buf ( n35379 , n6474 );
buf ( n35380 , n35379 );
xor ( n6477 , n6471 , n35380 );
buf ( n35382 , n6477 );
buf ( n35383 , n35382 );
xor ( n6480 , n6460 , n35383 );
buf ( n35385 , n6480 );
buf ( n35386 , n35385 );
buf ( n35387 , n527 );
buf ( n35388 , n550 );
and ( n6485 , n35387 , n35388 );
buf ( n35390 , n6485 );
buf ( n35391 , n35390 );
buf ( n35392 , n531 );
buf ( n35393 , n546 );
and ( n6490 , n35392 , n35393 );
buf ( n35395 , n6490 );
buf ( n35396 , n35395 );
xor ( n6493 , n35391 , n35396 );
buf ( n35398 , n532 );
buf ( n35399 , n545 );
and ( n6496 , n35398 , n35399 );
buf ( n35401 , n6496 );
buf ( n35402 , n35401 );
xor ( n6499 , n6493 , n35402 );
buf ( n35404 , n6499 );
buf ( n35405 , n35404 );
xor ( n6502 , n34982 , n34991 );
and ( n6503 , n6502 , n34995 );
and ( n6504 , n34982 , n34991 );
or ( n6505 , n6503 , n6504 );
buf ( n35410 , n6505 );
buf ( n35411 , n35410 );
xor ( n6508 , n35405 , n35411 );
buf ( n35413 , n536 );
buf ( n35414 , n541 );
and ( n6511 , n35413 , n35414 );
buf ( n35416 , n6511 );
buf ( n35417 , n35416 );
buf ( n35418 , n530 );
buf ( n35419 , n547 );
and ( n6516 , n35418 , n35419 );
buf ( n35421 , n6516 );
buf ( n35422 , n35421 );
xor ( n6519 , n35417 , n35422 );
buf ( n35424 , n461 );
buf ( n35425 , n525 );
buf ( n35426 , n552 );
and ( n6523 , n35425 , n35426 );
buf ( n35428 , n6523 );
buf ( n35429 , n35428 );
xor ( n6526 , n35424 , n35429 );
buf ( n35431 , n6526 );
buf ( n35432 , n35431 );
xor ( n6529 , n6519 , n35432 );
buf ( n35434 , n6529 );
buf ( n35435 , n35434 );
xor ( n6532 , n6508 , n35435 );
buf ( n35437 , n6532 );
buf ( n35438 , n35437 );
xor ( n6535 , n35386 , n35438 );
xor ( n6536 , n34977 , n34998 );
and ( n6537 , n6536 , n35066 );
and ( n35442 , n34977 , n34998 );
or ( n35443 , n6537 , n35442 );
buf ( n35444 , n35443 );
buf ( n35445 , n35444 );
xor ( n35446 , n6535 , n35445 );
buf ( n35447 , n35446 );
buf ( n35448 , n35447 );
xor ( n6548 , n6434 , n35448 );
buf ( n35450 , n6548 );
nor ( n35451 , n35296 , n35450 );
nor ( n6554 , n6381 , n35451 );
not ( n6555 , n6554 );
xor ( n6556 , n35260 , n35280 );
xor ( n6557 , n6556 , n35285 );
buf ( n35456 , n6557 );
buf ( n35457 , n35456 );
xor ( n6560 , n35128 , n35132 );
xor ( n6561 , n6560 , n35139 );
buf ( n35460 , n6561 );
buf ( n35461 , n35460 );
xor ( n6564 , n31588 , n31594 );
and ( n6565 , n6564 , n31616 );
and ( n6566 , n31588 , n31594 );
or ( n6567 , n6565 , n6566 );
buf ( n35466 , n6567 );
buf ( n35467 , n35466 );
xor ( n6570 , n35461 , n35467 );
xor ( n6571 , n35264 , n35268 );
xor ( n6572 , n6571 , n35275 );
buf ( n35471 , n6572 );
buf ( n35472 , n35471 );
and ( n6575 , n6570 , n35472 );
and ( n6576 , n35461 , n35467 );
or ( n6577 , n6575 , n6576 );
buf ( n35476 , n6577 );
buf ( n35477 , n35476 );
or ( n6580 , n35457 , n35477 );
buf ( n35479 , n6580 );
buf ( n35480 , n35479 );
not ( n6583 , n35480 );
xor ( n6584 , n35461 , n35467 );
xor ( n6585 , n6584 , n35472 );
buf ( n35484 , n6585 );
buf ( n35485 , n35484 );
xor ( n6588 , n31562 , n31568 );
and ( n6589 , n6588 , n31619 );
and ( n6590 , n31562 , n31568 );
or ( n6591 , n6589 , n6590 );
buf ( n35490 , n6591 );
buf ( n35491 , n35490 );
or ( n6594 , n35485 , n35491 );
buf ( n35493 , n6594 );
buf ( n35494 , n35493 );
not ( n6597 , n35494 );
buf ( n35496 , n31630 );
not ( n6599 , n35496 );
buf ( n35498 , n31656 );
not ( n6601 , n35498 );
or ( n6602 , n6599 , n6601 );
buf ( n35501 , n31635 );
nand ( n6604 , n6602 , n35501 );
buf ( n35503 , n6604 );
buf ( n35504 , n35503 );
not ( n6607 , n35504 );
or ( n6608 , n6597 , n6607 );
buf ( n35507 , n35484 );
buf ( n35508 , n35490 );
nand ( n6611 , n35507 , n35508 );
buf ( n35510 , n6611 );
buf ( n35511 , n35510 );
nand ( n6614 , n6608 , n35511 );
buf ( n35513 , n6614 );
buf ( n35514 , n35513 );
not ( n6617 , n35514 );
or ( n6618 , n6583 , n6617 );
buf ( n35517 , n35456 );
buf ( n35518 , n35476 );
nand ( n6621 , n35517 , n35518 );
buf ( n35520 , n6621 );
buf ( n35521 , n35520 );
nand ( n6624 , n6618 , n35521 );
buf ( n35523 , n6624 );
not ( n6626 , n35523 );
or ( n6627 , n6555 , n6626 );
not ( n6628 , n35451 );
buf ( n35527 , n35256 );
buf ( n35528 , n35289 );
nand ( n6631 , n35527 , n35528 );
buf ( n35530 , n6631 );
not ( n6633 , n35530 );
and ( n6634 , n6628 , n6633 );
buf ( n35533 , n35450 );
buf ( n35534 , n35296 );
and ( n6637 , n35533 , n35534 );
buf ( n35536 , n6637 );
nor ( n6639 , n6634 , n35536 );
nand ( n6640 , n6627 , n6639 );
buf ( n35539 , n6640 );
not ( n6642 , n35539 );
xor ( n6643 , n35344 , n35363 );
and ( n6644 , n6643 , n35383 );
and ( n6645 , n35344 , n35363 );
or ( n6646 , n6644 , n6645 );
buf ( n35545 , n6646 );
buf ( n35546 , n35545 );
xor ( n6649 , n35369 , n35374 );
and ( n6650 , n6649 , n35380 );
and ( n6651 , n35369 , n35374 );
or ( n6652 , n6650 , n6651 );
buf ( n35551 , n6652 );
buf ( n35552 , n35551 );
xor ( n6655 , n35349 , n35354 );
and ( n6656 , n6655 , n35360 );
and ( n6657 , n35349 , n35354 );
or ( n6658 , n6656 , n6657 );
buf ( n35557 , n6658 );
buf ( n35558 , n35557 );
xor ( n6661 , n35552 , n35558 );
buf ( n35560 , n535 );
buf ( n35561 , n541 );
and ( n6664 , n35560 , n35561 );
buf ( n35563 , n6664 );
buf ( n35564 , n35563 );
buf ( n35565 , n529 );
buf ( n35566 , n547 );
and ( n6669 , n35565 , n35566 );
buf ( n35568 , n6669 );
buf ( n35569 , n35568 );
xor ( n6672 , n35564 , n35569 );
buf ( n35571 , n536 );
buf ( n35572 , n540 );
and ( n6675 , n35571 , n35572 );
buf ( n35574 , n6675 );
buf ( n35575 , n35574 );
xor ( n6678 , n6672 , n35575 );
buf ( n35577 , n6678 );
buf ( n35578 , n35577 );
xor ( n6681 , n6661 , n35578 );
buf ( n35580 , n6681 );
buf ( n35581 , n35580 );
xor ( n6684 , n35546 , n35581 );
buf ( n35583 , n526 );
buf ( n35584 , n550 );
and ( n6690 , n35583 , n35584 );
buf ( n35586 , n6690 );
buf ( n35587 , n35586 );
buf ( n35588 , n530 );
buf ( n35589 , n546 );
and ( n6698 , n35588 , n35589 );
buf ( n35591 , n6698 );
buf ( n35592 , n35591 );
xor ( n6701 , n35587 , n35592 );
buf ( n35594 , n531 );
buf ( n35595 , n545 );
and ( n6704 , n35594 , n35595 );
buf ( n35597 , n6704 );
buf ( n35598 , n35597 );
xor ( n6707 , n6701 , n35598 );
buf ( n35600 , n6707 );
buf ( n35601 , n35600 );
buf ( n35602 , n527 );
buf ( n35603 , n549 );
and ( n6712 , n35602 , n35603 );
buf ( n35605 , n6712 );
buf ( n35606 , n35605 );
buf ( n35607 , n532 );
buf ( n35608 , n544 );
and ( n6717 , n35607 , n35608 );
buf ( n35610 , n6717 );
buf ( n35611 , n35610 );
xor ( n6720 , n35606 , n35611 );
buf ( n35613 , n533 );
buf ( n35614 , n543 );
and ( n6723 , n35613 , n35614 );
buf ( n35616 , n6723 );
buf ( n35617 , n35616 );
xor ( n6726 , n6720 , n35617 );
buf ( n35619 , n6726 );
buf ( n35620 , n35619 );
xor ( n6729 , n35601 , n35620 );
buf ( n35622 , n525 );
buf ( n35623 , n551 );
and ( n6732 , n35622 , n35623 );
buf ( n35625 , n6732 );
buf ( n35626 , n35625 );
buf ( n35627 , n528 );
buf ( n35628 , n548 );
and ( n6737 , n35627 , n35628 );
buf ( n35630 , n6737 );
buf ( n35631 , n35630 );
xor ( n6740 , n35626 , n35631 );
buf ( n35633 , n534 );
buf ( n35634 , n542 );
and ( n6743 , n35633 , n35634 );
buf ( n35636 , n6743 );
buf ( n35637 , n35636 );
xor ( n6746 , n6740 , n35637 );
buf ( n35639 , n6746 );
buf ( n35640 , n35639 );
xor ( n6749 , n6729 , n35640 );
buf ( n35642 , n6749 );
buf ( n35643 , n35642 );
xor ( n6752 , n6684 , n35643 );
buf ( n35645 , n6752 );
buf ( n35646 , n35645 );
xor ( n6755 , n35386 , n35438 );
and ( n6756 , n6755 , n35445 );
and ( n6757 , n35386 , n35438 );
or ( n6758 , n6756 , n6757 );
buf ( n35651 , n6758 );
buf ( n35652 , n35651 );
xor ( n6761 , n35646 , n35652 );
xor ( n6762 , n35405 , n35411 );
and ( n35655 , n6762 , n35435 );
and ( n6764 , n35405 , n35411 );
or ( n6765 , n35655 , n6764 );
buf ( n35658 , n6765 );
buf ( n35659 , n35658 );
xor ( n6768 , n35302 , n35308 );
and ( n6769 , n6768 , n35328 );
and ( n6770 , n35302 , n35308 );
or ( n6771 , n6769 , n6770 );
buf ( n35664 , n6771 );
buf ( n35665 , n35664 );
xor ( n6774 , n35659 , n35665 );
xor ( n6775 , n35417 , n35422 );
and ( n6776 , n6775 , n35432 );
and ( n6777 , n35417 , n35422 );
or ( n6778 , n6776 , n6777 );
buf ( n35671 , n6778 );
buf ( n35672 , n35671 );
xor ( n6781 , n35312 , n35318 );
and ( n6782 , n6781 , n35325 );
and ( n6783 , n35312 , n35318 );
or ( n6784 , n6782 , n6783 );
buf ( n35677 , n6784 );
buf ( n35678 , n35677 );
xor ( n6787 , n35672 , n35678 );
buf ( n35680 , n460 );
buf ( n35681 , n524 );
buf ( n35682 , n552 );
and ( n6791 , n35681 , n35682 );
buf ( n35684 , n6791 );
buf ( n35685 , n35684 );
xor ( n6794 , n35680 , n35685 );
buf ( n35687 , n6794 );
buf ( n35688 , n35687 );
and ( n6797 , n35424 , n35429 );
buf ( n35690 , n6797 );
buf ( n35691 , n35690 );
xor ( n6800 , n35688 , n35691 );
xor ( n6801 , n35391 , n35396 );
and ( n6802 , n6801 , n35402 );
and ( n6803 , n35391 , n35396 );
or ( n6804 , n6802 , n6803 );
buf ( n35697 , n6804 );
buf ( n35698 , n35697 );
xor ( n6807 , n6800 , n35698 );
buf ( n35700 , n6807 );
buf ( n35701 , n35700 );
xor ( n6810 , n6787 , n35701 );
buf ( n35703 , n6810 );
buf ( n35704 , n35703 );
xor ( n6813 , n6774 , n35704 );
buf ( n35706 , n6813 );
buf ( n35707 , n35706 );
xor ( n6816 , n6761 , n35707 );
buf ( n35709 , n6816 );
buf ( n35710 , n35709 );
xor ( n35711 , n35331 , n35337 );
and ( n35712 , n35711 , n35448 );
and ( n6821 , n35331 , n35337 );
or ( n6822 , n35712 , n6821 );
buf ( n35715 , n6822 );
buf ( n35716 , n35715 );
or ( n35717 , n35710 , n35716 );
buf ( n35718 , n35717 );
buf ( n35719 , n35718 );
buf ( n35720 , n35709 );
buf ( n35721 , n35715 );
nand ( n6836 , n35720 , n35721 );
buf ( n35723 , n6836 );
buf ( n35724 , n35723 );
nand ( n6839 , n35719 , n35724 );
buf ( n35726 , n6839 );
buf ( n35727 , n35726 );
not ( n6842 , n35727 );
or ( n6843 , n6642 , n6842 );
buf ( n35730 , n35726 );
buf ( n35731 , n6640 );
or ( n6846 , n35730 , n35731 );
nand ( n6847 , n6843 , n6846 );
buf ( n35734 , n6847 );
and ( n6849 , n35734 , n2356 );
nor ( n6850 , n6010 , n6849 );
nand ( n6851 , n6007 , n6850 );
not ( n6852 , n6851 );
not ( n6853 , n6852 );
buf ( n35740 , n35479 );
buf ( n35741 , n35520 );
nand ( n6856 , n35740 , n35741 );
buf ( n35743 , n6856 );
xnor ( n6858 , n35743 , n35513 );
not ( n6859 , n6858 );
not ( n6860 , n2356 );
or ( n6861 , n6859 , n6860 );
nand ( n6862 , n5981 , n5973 );
buf ( n35749 , n6862 );
not ( n6864 , n35749 );
buf ( n35751 , n6864 );
not ( n6866 , n35751 );
buf ( n35753 , n34884 );
not ( n6868 , n35753 );
buf ( n35755 , n6868 );
not ( n6870 , n35755 );
nand ( n6871 , n34703 , n5801 , n34724 );
not ( n6872 , n6871 );
or ( n6873 , n6870 , n6872 );
buf ( n35760 , n34900 );
not ( n6875 , n35760 );
buf ( n35762 , n6875 );
nand ( n6877 , n6873 , n35762 );
not ( n6878 , n6877 );
or ( n6879 , n6866 , n6878 );
nand ( n6880 , n6871 , n35755 );
and ( n6881 , n6880 , n6862 , n35762 );
nor ( n6882 , n6881 , n2618 );
nand ( n6883 , n6879 , n6882 );
nand ( n6884 , n6861 , n6883 );
not ( n6885 , n6884 );
not ( n6886 , n468 );
nand ( n6887 , n6885 , n6886 );
not ( n6888 , n2356 );
and ( n6889 , n35530 , n6380 );
xor ( n6890 , n6889 , n35523 );
not ( n6891 , n6890 );
or ( n6892 , n6888 , n6891 );
not ( n6893 , n5963 );
not ( n6894 , n6871 );
or ( n6895 , n6893 , n6894 );
not ( n35782 , n5982 );
nand ( n6897 , n6895 , n35782 );
not ( n6898 , n6897 );
buf ( n35785 , n34824 );
not ( n6900 , n35785 );
buf ( n35787 , n6900 );
buf ( n35788 , n35787 );
not ( n6903 , n35788 );
buf ( n35790 , n6903 );
buf ( n35791 , n35790 );
buf ( n35792 , n34909 );
nand ( n6907 , n35791 , n35792 );
buf ( n35794 , n6907 );
nand ( n6909 , n6898 , n35794 );
buf ( n35796 , n35794 );
not ( n6911 , n35796 );
buf ( n35798 , n6911 );
nand ( n6913 , n6897 , n35798 );
nand ( n6914 , n6909 , n6913 , n454 );
nand ( n6915 , n6892 , n6914 );
and ( n6916 , n6887 , n6915 );
not ( n6917 , n6916 );
not ( n6918 , n5963 );
nor ( n6919 , n6918 , n35787 );
buf ( n35806 , n6919 );
not ( n6921 , n35806 );
buf ( n6922 , n6871 );
buf ( n35809 , n6922 );
not ( n6924 , n35809 );
or ( n6925 , n6921 , n6924 );
and ( n6926 , n35790 , n5982 );
nor ( n6927 , n6926 , n34912 );
buf ( n35814 , n6927 );
nand ( n6929 , n6925 , n35814 );
buf ( n35816 , n6929 );
not ( n6931 , n35816 );
buf ( n35818 , n34781 );
buf ( n35819 , n34922 );
nand ( n6934 , n35818 , n35819 );
buf ( n35821 , n6934 );
nor ( n6936 , n35821 , n2618 );
and ( n6937 , n6931 , n6936 );
or ( n6938 , n35451 , n35536 );
buf ( n35825 , n6938 );
not ( n6940 , n35825 );
not ( n6941 , n6380 );
not ( n6942 , n35523 );
or ( n6943 , n6941 , n6942 );
nand ( n6944 , n6943 , n35530 );
buf ( n35831 , n6944 );
not ( n35832 , n35831 );
or ( n35833 , n6940 , n35832 );
buf ( n35834 , n6944 );
buf ( n35835 , n6938 );
or ( n35836 , n35834 , n35835 );
nand ( n6954 , n35833 , n35836 );
buf ( n35838 , n6954 );
and ( n6956 , n35838 , n2356 );
nor ( n6957 , n6937 , n6956 );
nand ( n35841 , n35816 , n35821 , n454 );
nand ( n6962 , n6957 , n35841 );
not ( n6963 , n6962 );
nor ( n6964 , n6917 , n6963 );
not ( n6965 , n6964 );
buf ( n35846 , n34694 );
not ( n6967 , n35846 );
buf ( n35848 , n6967 );
nand ( n6969 , n34728 , n5793 );
nand ( n6970 , n5793 , n5789 );
nand ( n6971 , n35848 , n6969 , n6970 );
not ( n6972 , n6971 );
not ( n6973 , n34700 );
nand ( n6974 , n6973 , n34682 );
nand ( n6975 , n6972 , n6974 );
not ( n6976 , n6974 );
nand ( n6977 , n6976 , n6971 );
nand ( n6978 , n6975 , n6977 , n454 );
nand ( n6979 , n6978 , n2617 );
nand ( n6980 , n6979 , n470 );
not ( n6981 , n6980 );
not ( n6982 , n5802 );
nand ( n6983 , n35755 , n35762 );
and ( n6984 , n6982 , n6983 );
not ( n6985 , n6982 );
not ( n6986 , n6983 );
and ( n6987 , n6985 , n6986 );
nor ( n6988 , n6984 , n6987 );
not ( n6989 , n6988 );
or ( n6990 , n6989 , n2356 );
buf ( n35871 , n35503 );
not ( n6992 , n35871 );
buf ( n35873 , n6992 );
not ( n6994 , n35873 );
buf ( n35875 , n35493 );
buf ( n35876 , n35510 );
and ( n6997 , n35875 , n35876 );
buf ( n35878 , n6997 );
not ( n6999 , n35878 );
or ( n7000 , n6994 , n6999 );
or ( n7001 , n35878 , n35873 );
nand ( n7002 , n7000 , n7001 );
nand ( n7003 , n7002 , n2356 );
not ( n7004 , n7003 );
nor ( n7005 , n7004 , n469 );
nand ( n7006 , n6990 , n7005 );
nand ( n7007 , n6981 , n7006 );
buf ( n35888 , n5793 );
buf ( n35889 , n35848 );
nand ( n7010 , n35888 , n35889 );
buf ( n35891 , n7010 );
not ( n7012 , n35891 );
buf ( n35893 , n5789 );
not ( n7014 , n35893 );
not ( n7015 , n34728 );
buf ( n35896 , n7015 );
nand ( n35897 , n7014 , n35896 );
buf ( n35898 , n35897 );
not ( n7019 , n35898 );
nand ( n7020 , n7012 , n7019 , n454 );
nand ( n7021 , n35891 , n35898 , n454 );
nand ( n7022 , n7020 , n7021 , n2476 );
not ( n7023 , n7022 );
not ( n7024 , n471 );
not ( n7025 , n472 );
not ( n7026 , n7025 );
nand ( n7027 , n7026 , n2358 );
nand ( n7028 , n7024 , n7027 );
not ( n7029 , n7028 );
or ( n7030 , n7023 , n7029 );
not ( n7031 , n7027 );
nand ( n7032 , n7031 , n471 );
nand ( n7033 , n7030 , n7032 );
not ( n7034 , n470 );
nand ( n7035 , n6975 , n454 , n6977 );
nand ( n7036 , n7034 , n7035 , n2617 );
nand ( n7037 , n7033 , n7006 , n7036 );
nand ( n7038 , n6988 , n454 );
nand ( n7039 , n7038 , n7003 );
nand ( n7040 , n7039 , n469 );
nand ( n7041 , n7007 , n7037 , n7040 );
buf ( n7042 , n7041 );
not ( n7043 , n7042 );
or ( n7044 , n6965 , n7043 );
buf ( n7045 , n6962 );
not ( n7046 , n6915 );
nand ( n7047 , n6884 , n468 );
nor ( n7048 , n7046 , n7047 );
nand ( n7049 , n7045 , n7048 );
nand ( n7050 , n7044 , n7049 );
not ( n7051 , n7050 );
or ( n7052 , n6853 , n7051 );
or ( n7053 , n6852 , n7050 );
nand ( n7054 , n7052 , n7053 );
not ( n7055 , n7054 );
or ( n7056 , n2630 , n7055 );
or ( n7057 , n2633 , n29502 );
nand ( n7058 , n7057 , n504 );
and ( n7059 , n456 , n465 );
not ( n7060 , n456 );
and ( n7061 , n7060 , n481 );
nor ( n7062 , n7059 , n7061 );
not ( n35943 , n7062 );
nand ( n35944 , n35943 , n29502 );
buf ( n7065 , n2678 );
not ( n7066 , n7065 );
and ( n35947 , n7058 , n35944 , n7066 );
buf ( n7071 , n29514 );
not ( n35949 , n7071 );
not ( n7073 , n497 );
buf ( n7074 , n973 );
not ( n35952 , n7074 );
not ( n7079 , n35952 );
or ( n7080 , n7073 , n7079 );
not ( n7081 , n497 );
nand ( n7082 , n7074 , n7081 );
nand ( n7083 , n7080 , n7082 );
not ( n7084 , n7083 );
or ( n7085 , n35949 , n7084 );
not ( n7086 , n498 );
not ( n7087 , n7074 );
not ( n7088 , n7087 );
or ( n7089 , n7086 , n7088 );
not ( n7090 , n7074 );
not ( n7091 , n7090 );
not ( n7092 , n498 );
nand ( n7093 , n7091 , n7092 );
nand ( n7094 , n7089 , n7093 );
not ( n7095 , n7094 );
not ( n7096 , n29514 );
and ( n7097 , n7074 , n7096 );
not ( n7098 , n7097 );
or ( n7099 , n7095 , n7098 );
nand ( n7100 , n7085 , n7099 );
xor ( n7101 , n35947 , n7100 );
not ( n7102 , n7062 );
not ( n7103 , n7102 );
and ( n7104 , n29502 , n7103 );
not ( n7105 , n29502 );
and ( n7106 , n7105 , n2633 );
nor ( n7107 , n7104 , n7106 );
not ( n7108 , n7107 );
and ( n7109 , n7108 , n504 );
not ( n7110 , n7071 );
not ( n7111 , n7094 );
or ( n7112 , n7110 , n7111 );
not ( n7113 , n499 );
not ( n7114 , n7087 );
or ( n7115 , n7113 , n7114 );
nand ( n7116 , n7074 , n1970 );
nand ( n7117 , n7115 , n7116 );
and ( n7118 , n7074 , n7096 );
nand ( n7119 , n7117 , n7118 );
nand ( n7120 , n7112 , n7119 );
xor ( n7121 , n7109 , n7120 );
not ( n7122 , n501 );
buf ( n7123 , n2831 );
not ( n7124 , n7123 );
and ( n7125 , n7122 , n7124 );
not ( n7126 , n7122 );
and ( n7127 , n7126 , n7123 );
nor ( n7128 , n7125 , n7127 );
not ( n7129 , n7128 );
xor ( n36004 , n29508 , n2831 );
not ( n7131 , n29508 );
not ( n7132 , n7090 );
and ( n7133 , n7131 , n7132 );
and ( n7134 , n35952 , n29508 );
nor ( n7135 , n7133 , n7134 );
and ( n7136 , n36004 , n7135 );
not ( n7137 , n7136 );
or ( n7138 , n7129 , n7137 );
xor ( n7139 , n7074 , n29508 );
not ( n7140 , n500 );
and ( n7141 , n7140 , n7124 );
not ( n7142 , n7140 );
and ( n7143 , n7142 , n2831 );
nor ( n7144 , n7141 , n7143 );
nand ( n7145 , n7139 , n7144 );
nand ( n7146 , n7138 , n7145 );
and ( n7147 , n7121 , n7146 );
and ( n7148 , n7109 , n7120 );
or ( n7149 , n7147 , n7148 );
xor ( n7150 , n7101 , n7149 );
not ( n7151 , n504 );
and ( n7152 , n7066 , n7151 );
and ( n7153 , n7065 , n504 );
nor ( n7154 , n7152 , n7153 );
not ( n7155 , n7154 );
not ( n7156 , n7155 );
not ( n7157 , n7065 );
and ( n7158 , n29502 , n7157 );
not ( n7159 , n29502 );
and ( n7160 , n7159 , n2671 );
nor ( n7161 , n7158 , n7160 );
and ( n7162 , n7161 , n7107 );
not ( n7163 , n7162 );
or ( n7164 , n7156 , n7163 );
not ( n7165 , n503 );
and ( n7166 , n7066 , n7165 );
and ( n7167 , n7065 , n503 );
nor ( n7168 , n7166 , n7167 );
or ( n7169 , n7168 , n7107 );
nand ( n36044 , n7164 , n7169 );
not ( n36045 , n7144 );
not ( n7172 , n7136 );
or ( n7173 , n36045 , n7172 );
not ( n36048 , n499 );
not ( n7178 , n2831 );
not ( n36050 , n7178 );
or ( n7180 , n36048 , n36050 );
nand ( n7181 , n7123 , n1970 );
nand ( n36053 , n7180 , n7181 );
nand ( n7186 , n7139 , n36053 );
nand ( n7187 , n7173 , n7186 );
xor ( n7188 , n36044 , n7187 );
buf ( n7189 , n933 );
not ( n7190 , n7189 );
and ( n7191 , n7190 , n2831 );
not ( n7192 , n7190 );
and ( n7193 , n7192 , n7178 );
nor ( n7194 , n7191 , n7193 );
not ( n7195 , n7194 );
not ( n7196 , n7195 );
and ( n7197 , n501 , n7103 );
not ( n7198 , n501 );
and ( n7199 , n7198 , n35943 );
nor ( n7200 , n7197 , n7199 );
not ( n7201 , n7200 );
not ( n7202 , n7201 );
or ( n7203 , n7196 , n7202 );
not ( n7204 , n502 );
and ( n7205 , n35943 , n7204 );
and ( n7206 , n7103 , n502 );
nor ( n7207 , n7205 , n7206 );
not ( n7208 , n7207 );
not ( n7209 , n2633 );
not ( n7210 , n7189 );
and ( n7211 , n7209 , n7210 );
and ( n7212 , n2633 , n7189 );
nor ( n7213 , n7211 , n7212 );
nand ( n7214 , n7194 , n7213 );
not ( n7215 , n7214 );
nand ( n7216 , n7208 , n7215 );
nand ( n7217 , n7203 , n7216 );
xor ( n7218 , n7188 , n7217 );
xor ( n7219 , n7150 , n7218 );
not ( n7220 , n7219 );
and ( n7221 , n503 , n7103 );
not ( n7222 , n503 );
and ( n7223 , n7222 , n2633 );
nor ( n7224 , n7221 , n7223 );
or ( n7225 , n7214 , n7224 );
not ( n7226 , n7195 );
or ( n7227 , n7226 , n7207 );
nand ( n7228 , n7225 , n7227 );
not ( n7229 , n7190 );
not ( n7230 , n7178 );
or ( n36099 , n7229 , n7230 );
nand ( n7232 , n36099 , n504 );
not ( n7233 , n7190 );
nand ( n7234 , n7233 , n7123 );
and ( n7235 , n7232 , n7234 , n35943 );
not ( n7236 , n7097 );
not ( n7237 , n500 );
not ( n7238 , n7087 );
or ( n7239 , n7237 , n7238 );
nand ( n7240 , n7074 , n7140 );
nand ( n7241 , n7239 , n7240 );
not ( n7242 , n7241 );
or ( n7243 , n7236 , n7242 );
nand ( n7244 , n7117 , n7071 );
nand ( n7245 , n7243 , n7244 );
and ( n7246 , n7235 , n7245 );
xor ( n7247 , n7228 , n7246 );
xor ( n7248 , n7109 , n7120 );
xor ( n7249 , n7248 , n7146 );
and ( n7250 , n7247 , n7249 );
and ( n7251 , n7228 , n7246 );
or ( n7252 , n7250 , n7251 );
not ( n7253 , n7252 );
nand ( n7254 , n7220 , n7253 );
nand ( n7255 , n7219 , n7252 );
nand ( n7256 , n7254 , n7255 );
not ( n7257 , n7256 );
xor ( n7258 , n7228 , n7246 );
xor ( n7259 , n7258 , n7249 );
not ( n7260 , n7259 );
and ( n7261 , n7204 , n7178 );
not ( n7262 , n7204 );
and ( n7263 , n7262 , n7123 );
nor ( n7264 , n7261 , n7263 );
not ( n7265 , n7264 );
not ( n7266 , n7136 );
or ( n36135 , n7265 , n7266 );
nand ( n36136 , n7139 , n7128 );
nand ( n7269 , n36135 , n36136 );
or ( n7270 , n7103 , n504 );
or ( n36139 , n35943 , n7151 );
nand ( n7275 , n7270 , n36139 );
not ( n36141 , n7275 );
not ( n7277 , n7215 );
or ( n7278 , n36141 , n7277 );
not ( n36144 , n7224 );
nand ( n7283 , n36144 , n7195 );
nand ( n7284 , n7278 , n7283 );
xor ( n7285 , n7269 , n7284 );
xor ( n7286 , n7235 , n7245 );
and ( n7287 , n7285 , n7286 );
and ( n7288 , n7269 , n7284 );
or ( n7289 , n7287 , n7288 );
not ( n7290 , n7289 );
nand ( n7291 , n7260 , n7290 );
not ( n7292 , n7291 );
xor ( n7293 , n7269 , n7284 );
xor ( n7294 , n7293 , n7286 );
not ( n7295 , n7294 );
and ( n7296 , n7195 , n504 );
xnor ( n7297 , n7123 , n7165 );
not ( n7298 , n7297 );
nand ( n7299 , n36004 , n7135 );
not ( n7300 , n7299 );
not ( n7301 , n7300 );
or ( n7302 , n7298 , n7301 );
nand ( n7303 , n7139 , n7264 );
nand ( n7304 , n7302 , n7303 );
xor ( n7305 , n7296 , n7304 );
not ( n7306 , n501 );
not ( n7307 , n35952 );
or ( n7308 , n7306 , n7307 );
nand ( n7309 , n7074 , n7122 );
nand ( n7310 , n7308 , n7309 );
not ( n7311 , n7310 );
or ( n7312 , n7311 , n7098 );
not ( n7313 , n7241 );
not ( n7314 , n7071 );
or ( n7315 , n7313 , n7314 );
nand ( n7316 , n7312 , n7315 );
and ( n7317 , n7305 , n7316 );
and ( n7318 , n7296 , n7304 );
or ( n7319 , n7317 , n7318 );
not ( n7320 , n7319 );
nand ( n7321 , n7295 , n7320 );
not ( n7322 , n7321 );
xor ( n7323 , n7296 , n7304 );
xor ( n36186 , n7323 , n7316 );
not ( n7325 , n7097 );
not ( n7326 , n502 );
not ( n7327 , n35952 );
or ( n7328 , n7326 , n7327 );
nand ( n7329 , n7091 , n7204 );
nand ( n7330 , n7328 , n7329 );
not ( n7331 , n7330 );
or ( n7332 , n7325 , n7331 );
nand ( n7333 , n7310 , n7071 );
nand ( n7334 , n7332 , n7333 );
not ( n7335 , n7334 );
and ( n7336 , n7091 , n29508 );
nor ( n7337 , n7336 , n7178 );
or ( n7338 , n7074 , n29508 );
nand ( n7339 , n7338 , n504 );
nand ( n7340 , n7337 , n7339 );
nor ( n7341 , n7335 , n7340 );
nor ( n7342 , n36186 , n7341 );
not ( n7343 , n7334 );
not ( n7344 , n7340 );
and ( n7345 , n7343 , n7344 );
and ( n7346 , n7334 , n7340 );
nor ( n7347 , n7345 , n7346 );
not ( n7348 , n7299 );
and ( n7349 , n7124 , n504 );
not ( n7350 , n7178 );
and ( n7351 , n7350 , n7151 );
nor ( n7352 , n7349 , n7351 );
not ( n7353 , n7352 );
and ( n36216 , n7348 , n7353 );
and ( n7355 , n7139 , n7297 );
nor ( n36218 , n36216 , n7355 );
and ( n7360 , n7347 , n36218 );
not ( n36220 , n7071 );
not ( n7362 , n7330 );
or ( n7363 , n36220 , n7362 );
not ( n36223 , n503 );
not ( n7368 , n7087 );
or ( n7369 , n36223 , n7368 );
nand ( n7370 , n7091 , n7165 );
nand ( n7371 , n7369 , n7370 );
nand ( n7372 , n7371 , n7118 );
nand ( n7373 , n7363 , n7372 );
and ( n7374 , n7139 , n504 );
nor ( n7375 , n7373 , n7374 );
nand ( n7376 , n7071 , n504 );
nand ( n7377 , n7091 , n7376 );
not ( n7378 , n7377 );
not ( n7379 , n7071 );
not ( n7380 , n7371 );
or ( n7381 , n7379 , n7380 );
nand ( n7382 , n29578 , n7097 );
nand ( n7383 , n7381 , n7382 );
nand ( n7384 , n7378 , n7383 );
or ( n7385 , n7375 , n7384 );
nand ( n7386 , n7373 , n7374 );
nand ( n7387 , n7385 , n7386 );
not ( n7388 , n7387 );
or ( n7389 , n7360 , n7388 );
or ( n7390 , n7347 , n36218 );
nand ( n7391 , n7389 , n7390 );
not ( n7392 , n7391 );
or ( n7393 , n7342 , n7392 );
nand ( n7394 , n36186 , n7341 );
nand ( n7395 , n7393 , n7394 );
not ( n7396 , n7395 );
or ( n7397 , n7322 , n7396 );
or ( n7398 , n7295 , n7320 );
nand ( n7399 , n7397 , n7398 );
not ( n7400 , n7399 );
or ( n7401 , n7292 , n7400 );
nand ( n7402 , n7259 , n7289 );
nand ( n36259 , n7401 , n7402 );
not ( n7404 , n36259 );
or ( n7405 , n7257 , n7404 );
or ( n7406 , n36259 , n7256 );
nand ( n7407 , n7405 , n7406 );
nand ( n7408 , n7407 , n2628 );
nand ( n7409 , n7056 , n7408 );
not ( n7410 , n2628 );
not ( n7411 , n7410 );
nand ( n7412 , n5642 , n5631 );
buf ( n36269 , n7412 );
not ( n7414 , n36269 );
buf ( n36271 , n539 );
not ( n7416 , n36271 );
not ( n7417 , n29519 );
and ( n7418 , n5352 , n5093 , n4818 );
not ( n7419 , n7418 );
not ( n7420 , n4913 );
or ( n7421 , n7419 , n7420 );
not ( n7422 , n34042 );
not ( n7423 , n34047 );
and ( n7424 , n7422 , n7423 );
nor ( n7425 , n7424 , n5351 );
and ( n7426 , n7425 , n4919 );
or ( n7427 , n5351 , n5090 );
nand ( n7428 , n7427 , n5353 );
nor ( n36285 , n7426 , n7428 );
nand ( n7433 , n7421 , n36285 );
not ( n36287 , n5180 );
not ( n7435 , n491 );
nand ( n7436 , n7435 , n5168 , n489 );
nand ( n36290 , n7436 , n5171 );
not ( n7441 , n36290 );
or ( n7442 , n36287 , n7441 );
buf ( n36293 , n4928 );
xor ( n7444 , n489 , n518 );
buf ( n36295 , n7444 );
nand ( n7446 , n36293 , n36295 );
buf ( n36297 , n7446 );
nand ( n7448 , n7442 , n36297 );
buf ( n36299 , n5193 );
not ( n7450 , n36299 );
buf ( n36301 , n497 );
buf ( n36302 , n498 );
xnor ( n7453 , n36301 , n36302 );
buf ( n36304 , n7453 );
nor ( n7455 , n36304 , n29602 );
buf ( n36306 , n7455 );
not ( n7457 , n36306 );
or ( n7458 , n7450 , n7457 );
buf ( n36309 , n29604 );
xor ( n7460 , n497 , n510 );
buf ( n36311 , n7460 );
nand ( n7462 , n36309 , n36311 );
buf ( n36313 , n7462 );
buf ( n36314 , n36313 );
nand ( n7465 , n7458 , n36314 );
buf ( n36316 , n7465 );
xor ( n7467 , n7448 , n36316 );
not ( n7468 , n5241 );
buf ( n36319 , n33190 );
buf ( n36320 , n33184 );
buf ( n36321 , n33178 );
and ( n36322 , n36319 , n36320 , n36321 );
buf ( n36323 , n36322 );
not ( n7474 , n36323 );
or ( n7475 , n7468 , n7474 );
buf ( n36326 , n30846 );
buf ( n36327 , n512 );
buf ( n36328 , n495 );
xor ( n7479 , n36327 , n36328 );
buf ( n36330 , n7479 );
buf ( n36331 , n36330 );
nand ( n7482 , n36326 , n36331 );
buf ( n36333 , n7482 );
nand ( n7484 , n7475 , n36333 );
xor ( n7485 , n7467 , n7484 );
not ( n7486 , n7485 );
buf ( n36337 , n520 );
buf ( n36338 , n489 );
and ( n7489 , n36337 , n36338 );
buf ( n36340 , n7489 );
buf ( n36341 , n36340 );
buf ( n36342 , n5313 );
not ( n7496 , n36342 );
buf ( n36344 , n29582 );
not ( n7498 , n36344 );
or ( n7499 , n7496 , n7498 );
buf ( n36347 , n503 );
buf ( n36348 , n504 );
nand ( n7505 , n36347 , n36348 );
buf ( n36350 , n7505 );
buf ( n36351 , n36350 );
nand ( n7508 , n7499 , n36351 );
buf ( n36353 , n7508 );
buf ( n36354 , n36353 );
xor ( n7511 , n36341 , n36354 );
buf ( n36356 , n5157 );
not ( n7513 , n36356 );
buf ( n36358 , n34104 );
not ( n7515 , n36358 );
or ( n7516 , n7513 , n7515 );
buf ( n36361 , n29646 );
buf ( n36362 , n506 );
buf ( n36363 , n501 );
xor ( n7520 , n36362 , n36363 );
buf ( n36365 , n7520 );
buf ( n36366 , n36365 );
nand ( n7523 , n36361 , n36366 );
buf ( n36368 , n7523 );
buf ( n36369 , n36368 );
nand ( n7526 , n7516 , n36369 );
buf ( n36371 , n7526 );
buf ( n36372 , n36371 );
xor ( n36373 , n7511 , n36372 );
buf ( n36374 , n36373 );
not ( n7531 , n36374 );
nand ( n7532 , n7486 , n7531 );
not ( n7533 , n7532 );
not ( n7534 , n5284 );
nor ( n7535 , n33357 , n33353 );
not ( n7536 , n7535 );
or ( n7537 , n7534 , n7536 );
buf ( n36382 , n33102 );
xor ( n7539 , n491 , n516 );
buf ( n36384 , n7539 );
nand ( n7541 , n36382 , n36384 );
buf ( n36386 , n7541 );
nand ( n36387 , n7537 , n36386 );
not ( n7547 , n4218 );
xor ( n36389 , n493 , n514 );
not ( n7549 , n36389 );
or ( n7550 , n7547 , n7549 );
nand ( n36392 , n4387 , n34170 );
nand ( n7555 , n7550 , n36392 );
xor ( n7556 , n36387 , n7555 );
buf ( n36395 , n5232 );
not ( n7558 , n36395 );
buf ( n36397 , n30741 );
not ( n7560 , n36397 );
or ( n7561 , n7558 , n7560 );
buf ( n36400 , n29543 );
xor ( n7563 , n499 , n508 );
buf ( n36402 , n7563 );
nand ( n7565 , n36400 , n36402 );
buf ( n36404 , n7565 );
buf ( n36405 , n36404 );
nand ( n7568 , n7561 , n36405 );
buf ( n36407 , n7568 );
xor ( n7570 , n7556 , n36407 );
buf ( n7571 , n7570 );
nand ( n7572 , n7533 , n7571 );
nand ( n7573 , n7485 , n36374 );
not ( n7574 , n7573 );
nand ( n7575 , n7574 , n7571 );
not ( n36414 , n7571 );
nor ( n7577 , n7486 , n36374 );
nand ( n7578 , n36414 , n7577 );
not ( n36417 , n36374 );
nor ( n7583 , n36417 , n7485 );
nand ( n7584 , n36414 , n7583 );
nand ( n7585 , n7572 , n7575 , n7578 , n7584 );
buf ( n36421 , n7585 );
xor ( n7587 , n34223 , n34279 );
and ( n7588 , n7587 , n34286 );
and ( n7589 , n34223 , n34279 );
or ( n7590 , n7588 , n7589 );
buf ( n36426 , n7590 );
buf ( n36427 , n36426 );
xor ( n7593 , n36421 , n36427 );
xor ( n7594 , n34237 , n34270 );
and ( n7595 , n7594 , n34276 );
and ( n7596 , n34237 , n34270 );
or ( n7597 , n7595 , n7596 );
buf ( n36433 , n7597 );
buf ( n36434 , n36433 );
and ( n7603 , n34253 , n34267 );
buf ( n36436 , n7603 );
buf ( n36437 , n36436 );
or ( n36438 , n34115 , n34151 );
nand ( n7610 , n36438 , n34136 );
buf ( n36440 , n34115 );
buf ( n36441 , n34151 );
nand ( n7613 , n36440 , n36441 );
buf ( n36443 , n7613 );
nand ( n36444 , n7610 , n36443 );
buf ( n36445 , n36444 );
xor ( n7620 , n36437 , n36445 );
xor ( n36447 , n34176 , n34191 );
and ( n7622 , n36447 , n34204 );
and ( n7623 , n34176 , n34191 );
or ( n36450 , n7622 , n7623 );
buf ( n36451 , n36450 );
buf ( n36452 , n36451 );
xor ( n36453 , n7620 , n36452 );
buf ( n36454 , n36453 );
buf ( n36455 , n36454 );
xor ( n36456 , n36434 , n36455 );
xor ( n7637 , n34099 , n34162 );
and ( n7638 , n7637 , n34207 );
and ( n36459 , n34099 , n34162 );
or ( n7640 , n7638 , n36459 );
buf ( n36461 , n7640 );
buf ( n36462 , n36461 );
xor ( n7646 , n36456 , n36462 );
buf ( n36464 , n7646 );
buf ( n36465 , n36464 );
xor ( n36466 , n7593 , n36465 );
buf ( n36467 , n36466 );
xor ( n36468 , n34210 , n34216 );
and ( n36469 , n36468 , n34289 );
and ( n36470 , n34210 , n34216 );
or ( n36471 , n36469 , n36470 );
buf ( n36472 , n36471 );
nor ( n36473 , n36467 , n36472 );
not ( n36474 , n36473 );
nand ( n36475 , n36467 , n36472 );
nand ( n36476 , n36474 , n36475 );
not ( n36477 , n36476 );
and ( n36478 , n7433 , n36477 );
not ( n36479 , n7433 );
and ( n36480 , n36479 , n36476 );
nor ( n36481 , n36478 , n36480 );
not ( n36482 , n36481 );
or ( n36483 , n7417 , n36482 );
not ( n36484 , n3072 );
not ( n36485 , n34409 );
or ( n36486 , n36484 , n36485 );
nand ( n36487 , n1492 , n1494 );
and ( n36488 , n36487 , n30599 );
and ( n36489 , n2803 , n36488 );
not ( n36490 , n2803 );
and ( n36491 , n36487 , n497 );
and ( n36492 , n36490 , n36491 );
nor ( n36493 , n36489 , n36492 );
nand ( n36494 , n36486 , n36493 );
not ( n36495 , n31812 );
not ( n36496 , n5386 );
or ( n36497 , n36495 , n36496 );
and ( n36498 , n29501 , n31784 );
not ( n36499 , n29501 );
and ( n36500 , n36499 , n495 );
or ( n36501 , n36498 , n36500 );
buf ( n36502 , n36501 );
buf ( n36503 , n1914 );
nand ( n36504 , n36502 , n36503 );
buf ( n36505 , n36504 );
nand ( n36506 , n36497 , n36505 );
xor ( n36507 , n36494 , n36506 );
buf ( n36508 , n3832 );
buf ( n36509 , n36508 );
not ( n36510 , n36509 );
xor ( n36511 , n489 , n29513 );
buf ( n36512 , n36511 );
not ( n36513 , n36512 );
or ( n36514 , n36510 , n36513 );
nand ( n36515 , n5441 , n5418 );
buf ( n36516 , n36515 );
nand ( n36517 , n36514 , n36516 );
buf ( n36518 , n36517 );
xor ( n36519 , n36507 , n36518 );
buf ( n36520 , n36519 );
not ( n36521 , n36520 );
buf ( n36522 , n29939 );
buf ( n36523 , n489 );
and ( n36524 , n36522 , n36523 );
buf ( n36525 , n36524 );
buf ( n36526 , n36525 );
buf ( n36527 , n29966 );
not ( n36528 , n36527 );
buf ( n36529 , n34509 );
not ( n36530 , n36529 );
or ( n36531 , n36528 , n36530 );
buf ( n36532 , n503 );
buf ( n36533 , n504 );
nand ( n36534 , n36532 , n36533 );
buf ( n36535 , n36534 );
buf ( n36536 , n36535 );
nand ( n36537 , n36531 , n36536 );
buf ( n36538 , n36537 );
buf ( n36539 , n36538 );
xor ( n36540 , n36526 , n36539 );
buf ( n36541 , n32034 );
not ( n36542 , n36541 );
buf ( n36543 , n34435 );
not ( n36544 , n36543 );
or ( n36545 , n36542 , n36544 );
or ( n36546 , n3855 , n743 );
nand ( n36547 , n3855 , n984 );
nand ( n36548 , n36546 , n36547 );
buf ( n36549 , n36548 );
buf ( n36550 , n1010 );
nand ( n36551 , n36549 , n36550 );
buf ( n36552 , n36551 );
buf ( n36553 , n36552 );
nand ( n36554 , n36545 , n36553 );
buf ( n36555 , n36554 );
buf ( n36556 , n36555 );
xor ( n36557 , n36540 , n36556 );
buf ( n36558 , n36557 );
not ( n36559 , n36558 );
buf ( n36560 , n798 );
not ( n36561 , n36560 );
buf ( n36562 , n36561 );
buf ( n36563 , n36562 );
not ( n36564 , n36563 );
buf ( n36565 , n5404 );
not ( n36566 , n36565 );
or ( n36567 , n36564 , n36566 );
buf ( n36568 , n499 );
not ( n36569 , n36568 );
buf ( n36570 , n3211 );
not ( n36571 , n36570 );
or ( n36572 , n36569 , n36571 );
not ( n36573 , n456 );
nand ( n36574 , n36573 , n3218 );
nand ( n36575 , n3215 , n456 );
nand ( n36576 , n36574 , n36575 , n29901 );
buf ( n36577 , n36576 );
nand ( n36578 , n36572 , n36577 );
buf ( n36579 , n36578 );
nand ( n36580 , n36579 , n745 );
buf ( n36581 , n36580 );
nand ( n36582 , n36567 , n36581 );
buf ( n36583 , n36582 );
not ( n36584 , n3045 );
buf ( n36585 , n491 );
not ( n36586 , n36585 );
buf ( n36587 , n854 );
not ( n36588 , n36587 );
or ( n36589 , n36586 , n36588 );
buf ( n36590 , n29507 );
buf ( n36591 , n3524 );
nand ( n36592 , n36590 , n36591 );
buf ( n36593 , n36592 );
buf ( n36594 , n36593 );
nand ( n36595 , n36589 , n36594 );
buf ( n36596 , n36595 );
not ( n36597 , n36596 );
or ( n36598 , n36584 , n36597 );
nand ( n36599 , n5535 , n3948 );
nand ( n36600 , n36598 , n36599 );
xor ( n36601 , n36583 , n36600 );
buf ( n36602 , n2978 );
not ( n36603 , n36602 );
not ( n36604 , n493 );
not ( n36605 , n929 );
or ( n36606 , n36604 , n36605 );
nand ( n36607 , n3063 , n2704 );
nand ( n36608 , n36606 , n36607 );
buf ( n36609 , n36608 );
not ( n36610 , n36609 );
or ( n36611 , n36603 , n36610 );
not ( n36612 , n5371 );
not ( n36613 , n5373 );
or ( n36614 , n36612 , n36613 );
nand ( n36615 , n36614 , n3511 );
buf ( n36616 , n36615 );
nand ( n36617 , n36611 , n36616 );
buf ( n36618 , n36617 );
xor ( n36619 , n36601 , n36618 );
nor ( n36620 , n36559 , n36619 );
nand ( n36621 , n36521 , n36620 );
not ( n36622 , n36558 );
and ( n36623 , n36619 , n36622 );
nand ( n36624 , n36521 , n36623 );
nand ( n36625 , n36619 , n36558 );
not ( n36626 , n36625 );
nand ( n36627 , n36626 , n36520 );
not ( n36628 , n36619 );
nand ( n36629 , n36628 , n36622 );
not ( n36630 , n36629 );
nand ( n36631 , n36630 , n36520 );
nand ( n36632 , n36621 , n36624 , n36627 , n36631 );
buf ( n36633 , n36632 );
xor ( n36634 , n34461 , n34525 );
and ( n36635 , n36634 , n34549 );
and ( n36636 , n34461 , n34525 );
or ( n36637 , n36635 , n36636 );
buf ( n36638 , n36637 );
buf ( n36639 , n36638 );
xor ( n36640 , n36633 , n36639 );
xor ( n36641 , n5537 , n5577 );
and ( n36642 , n36641 , n34523 );
and ( n36643 , n5537 , n5577 );
or ( n36644 , n36642 , n36643 );
buf ( n36645 , n36644 );
and ( n36646 , n5546 , n34516 );
buf ( n36647 , n36646 );
not ( n36648 , n34442 );
not ( n36649 , n5443 );
not ( n36650 , n3072 );
nor ( n36651 , n36650 , n4005 );
buf ( n36652 , n34409 );
not ( n36653 , n36652 );
buf ( n36654 , n33014 );
nor ( n36655 , n36653 , n36654 );
buf ( n36656 , n36655 );
nor ( n36657 , n36651 , n36656 );
nand ( n36658 , n36649 , n36657 );
not ( n36659 , n36658 );
or ( n36660 , n36648 , n36659 );
not ( n36661 , n5418 );
not ( n36662 , n5434 );
or ( n36663 , n36661 , n36662 );
nand ( n36664 , n36663 , n5442 );
nand ( n36665 , n36664 , n34416 );
nand ( n36666 , n36660 , n36665 );
buf ( n36667 , n36666 );
xor ( n36668 , n36647 , n36667 );
xor ( n36669 , n34324 , n34338 );
and ( n36670 , n36669 , n34353 );
and ( n36671 , n34324 , n34338 );
or ( n36672 , n36670 , n36671 );
buf ( n36673 , n36672 );
buf ( n36674 , n36673 );
xor ( n36675 , n36668 , n36674 );
buf ( n36676 , n36675 );
buf ( n36677 , n36676 );
xor ( n36678 , n36645 , n36677 );
xor ( n36679 , n34313 , n34356 );
and ( n36680 , n36679 , n34446 );
and ( n36681 , n34313 , n34356 );
or ( n36682 , n36680 , n36681 );
buf ( n36683 , n36682 );
buf ( n36684 , n36683 );
xor ( n36685 , n36678 , n36684 );
buf ( n36686 , n36685 );
buf ( n36687 , n36686 );
xor ( n36688 , n36640 , n36687 );
buf ( n36689 , n36688 );
xor ( n36690 , n34449 , n34454 );
and ( n36691 , n36690 , n34552 );
and ( n36692 , n34449 , n34454 );
or ( n36693 , n36691 , n36692 );
buf ( n36694 , n36693 );
nor ( n36695 , n36689 , n36694 );
not ( n36696 , n36695 );
nand ( n36697 , n36689 , n36694 );
buf ( n36698 , n36697 );
and ( n36699 , n36696 , n36698 );
not ( n36700 , n5881 );
nor ( n36701 , n33037 , n4035 );
not ( n36702 , n36701 );
nand ( n36703 , n5626 , n3671 , n36702 );
not ( n36704 , n36703 );
not ( n36705 , n36704 );
or ( n36706 , n36700 , n36705 );
nor ( n36707 , n5625 , n36701 );
and ( n36708 , n3798 , n36707 );
nor ( n36709 , n34554 , n5624 );
or ( n36710 , n36709 , n4037 );
nand ( n36711 , n36710 , n5627 );
nor ( n36712 , n36708 , n36711 );
nand ( n36713 , n36706 , n36712 );
xor ( n36714 , n36699 , n36713 );
nand ( n36715 , n36714 , n455 );
nand ( n36716 , n36483 , n36715 );
buf ( n36717 , n36716 );
not ( n36718 , n36717 );
or ( n36719 , n7416 , n36718 );
not ( n36720 , n29519 );
not ( n36721 , n36481 );
or ( n36722 , n36720 , n36721 );
and ( n36723 , n36714 , n455 );
nor ( n36724 , n36723 , n539 );
nand ( n36725 , n36722 , n36724 );
buf ( n36726 , n36725 );
nand ( n36727 , n36719 , n36726 );
buf ( n36728 , n36727 );
buf ( n36729 , n36728 );
not ( n36730 , n36729 );
or ( n36731 , n7414 , n36730 );
or ( n36732 , n36728 , n7412 );
buf ( n36733 , n36732 );
nand ( n36734 , n36731 , n36733 );
buf ( n36735 , n36734 );
buf ( n36736 , n36735 );
not ( n36737 , n36736 );
buf ( n36738 , n36737 );
not ( n36739 , n36738 );
not ( n36740 , n5982 );
not ( n36741 , n5970 );
or ( n36742 , n36740 , n36741 );
not ( n36743 , n6001 );
nand ( n36744 , n36742 , n36743 );
nand ( n36745 , n36744 , n5662 );
buf ( n36746 , n34888 );
nand ( n36747 , n6922 , n36746 , n5662 );
nand ( n36748 , n36745 , n5660 , n36747 );
not ( n36749 , n36748 );
or ( n36750 , n36739 , n36749 );
and ( n36751 , n36735 , n5660 );
and ( n36752 , n36751 , n36745 , n36747 );
nor ( n36753 , n36752 , n2618 );
nand ( n36754 , n36750 , n36753 );
xor ( n36755 , n35646 , n35652 );
and ( n36756 , n36755 , n35707 );
and ( n36757 , n35646 , n35652 );
or ( n36758 , n36756 , n36757 );
buf ( n36759 , n36758 );
buf ( n36760 , n36759 );
xor ( n36761 , n35587 , n35592 );
and ( n36762 , n36761 , n35598 );
and ( n36763 , n35587 , n35592 );
or ( n36764 , n36762 , n36763 );
buf ( n36765 , n36764 );
buf ( n36766 , n36765 );
xor ( n36767 , n35606 , n35611 );
and ( n36768 , n36767 , n35617 );
and ( n36769 , n35606 , n35611 );
or ( n36770 , n36768 , n36769 );
buf ( n36771 , n36770 );
buf ( n36772 , n36771 );
xor ( n36773 , n36766 , n36772 );
xor ( n36774 , n35564 , n35569 );
and ( n36775 , n36774 , n35575 );
and ( n36776 , n35564 , n35569 );
or ( n36777 , n36775 , n36776 );
buf ( n36778 , n36777 );
buf ( n36779 , n36778 );
xor ( n36780 , n36773 , n36779 );
buf ( n36781 , n36780 );
buf ( n36782 , n36781 );
xor ( n36783 , n35626 , n35631 );
and ( n36784 , n36783 , n35637 );
and ( n36785 , n35626 , n35631 );
or ( n36786 , n36784 , n36785 );
buf ( n36787 , n36786 );
buf ( n36788 , n36787 );
buf ( n36789 , n534 );
buf ( n36790 , n541 );
and ( n36791 , n36789 , n36790 );
buf ( n36792 , n36791 );
buf ( n36793 , n36792 );
buf ( n36794 , n528 );
buf ( n36795 , n547 );
and ( n36796 , n36794 , n36795 );
buf ( n36797 , n36796 );
buf ( n36798 , n36797 );
xor ( n36799 , n36793 , n36798 );
buf ( n36800 , n535 );
buf ( n36801 , n540 );
and ( n36802 , n36800 , n36801 );
buf ( n36803 , n36802 );
buf ( n36804 , n36803 );
xor ( n36805 , n36799 , n36804 );
buf ( n36806 , n36805 );
buf ( n36807 , n36806 );
xor ( n36808 , n36788 , n36807 );
buf ( n36809 , n525 );
buf ( n36810 , n550 );
and ( n36811 , n36809 , n36810 );
buf ( n36812 , n36811 );
buf ( n36813 , n36812 );
buf ( n36814 , n529 );
buf ( n36815 , n546 );
and ( n36816 , n36814 , n36815 );
buf ( n36817 , n36816 );
buf ( n36818 , n36817 );
xor ( n36819 , n36813 , n36818 );
buf ( n36820 , n530 );
buf ( n36821 , n545 );
and ( n36822 , n36820 , n36821 );
buf ( n36823 , n36822 );
buf ( n36824 , n36823 );
xor ( n36825 , n36819 , n36824 );
buf ( n36826 , n36825 );
buf ( n36827 , n36826 );
xor ( n36828 , n36808 , n36827 );
buf ( n36829 , n36828 );
buf ( n36830 , n36829 );
xor ( n36831 , n36782 , n36830 );
xor ( n36832 , n35672 , n35678 );
and ( n36833 , n36832 , n35701 );
and ( n36834 , n35672 , n35678 );
or ( n36835 , n36833 , n36834 );
buf ( n36836 , n36835 );
buf ( n36837 , n36836 );
xor ( n36838 , n36831 , n36837 );
buf ( n36839 , n36838 );
buf ( n36840 , n36839 );
xor ( n36841 , n35659 , n35665 );
and ( n36842 , n36841 , n35704 );
and ( n36843 , n35659 , n35665 );
or ( n36844 , n36842 , n36843 );
buf ( n36845 , n36844 );
buf ( n36846 , n36845 );
xor ( n36847 , n36840 , n36846 );
buf ( n36848 , n526 );
buf ( n36849 , n549 );
and ( n36850 , n36848 , n36849 );
buf ( n36851 , n36850 );
buf ( n36852 , n36851 );
buf ( n36853 , n531 );
buf ( n36854 , n544 );
and ( n36855 , n36853 , n36854 );
buf ( n36856 , n36855 );
buf ( n36857 , n36856 );
xor ( n36858 , n36852 , n36857 );
buf ( n36859 , n532 );
buf ( n36860 , n543 );
and ( n36861 , n36859 , n36860 );
buf ( n36862 , n36861 );
buf ( n36863 , n36862 );
xor ( n36864 , n36858 , n36863 );
buf ( n36865 , n36864 );
buf ( n36866 , n36865 );
buf ( n36867 , n524 );
buf ( n36868 , n551 );
and ( n36869 , n36867 , n36868 );
buf ( n36870 , n36869 );
buf ( n36871 , n36870 );
buf ( n36872 , n527 );
buf ( n36873 , n548 );
and ( n36874 , n36872 , n36873 );
buf ( n36875 , n36874 );
buf ( n36876 , n36875 );
xor ( n36877 , n36871 , n36876 );
buf ( n36878 , n533 );
buf ( n36879 , n542 );
and ( n36880 , n36878 , n36879 );
buf ( n36881 , n36880 );
buf ( n36882 , n36881 );
xor ( n36883 , n36877 , n36882 );
buf ( n36884 , n36883 );
buf ( n36885 , n36884 );
xor ( n36886 , n36866 , n36885 );
buf ( n36887 , n536 );
buf ( n36888 , n539 );
and ( n36889 , n36887 , n36888 );
buf ( n36890 , n36889 );
buf ( n36891 , n36890 );
buf ( n36892 , n459 );
buf ( n36893 , n523 );
buf ( n36894 , n552 );
and ( n36895 , n36893 , n36894 );
buf ( n36896 , n36895 );
buf ( n36897 , n36896 );
xor ( n36898 , n36892 , n36897 );
buf ( n36899 , n36898 );
buf ( n36900 , n36899 );
xor ( n36901 , n36891 , n36900 );
and ( n36902 , n35680 , n35685 );
buf ( n36903 , n36902 );
buf ( n36904 , n36903 );
xor ( n36905 , n36901 , n36904 );
buf ( n36906 , n36905 );
buf ( n36907 , n36906 );
xor ( n36908 , n36886 , n36907 );
buf ( n36909 , n36908 );
buf ( n36910 , n36909 );
xor ( n36911 , n35546 , n35581 );
and ( n36912 , n36911 , n35643 );
and ( n36913 , n35546 , n35581 );
or ( n36914 , n36912 , n36913 );
buf ( n36915 , n36914 );
buf ( n36916 , n36915 );
xor ( n36917 , n36910 , n36916 );
xor ( n36918 , n35688 , n35691 );
and ( n36919 , n36918 , n35698 );
and ( n36920 , n35688 , n35691 );
or ( n36921 , n36919 , n36920 );
buf ( n36922 , n36921 );
buf ( n36923 , n36922 );
xor ( n36924 , n35601 , n35620 );
and ( n36925 , n36924 , n35640 );
and ( n36926 , n35601 , n35620 );
or ( n36927 , n36925 , n36926 );
buf ( n36928 , n36927 );
buf ( n36929 , n36928 );
xor ( n36930 , n36923 , n36929 );
xor ( n36931 , n35552 , n35558 );
and ( n36932 , n36931 , n35578 );
and ( n36933 , n35552 , n35558 );
or ( n36934 , n36932 , n36933 );
buf ( n36935 , n36934 );
buf ( n36936 , n36935 );
xor ( n36937 , n36930 , n36936 );
buf ( n36938 , n36937 );
buf ( n36939 , n36938 );
xor ( n36940 , n36917 , n36939 );
buf ( n36941 , n36940 );
buf ( n36942 , n36941 );
xor ( n36943 , n36847 , n36942 );
buf ( n36944 , n36943 );
buf ( n36945 , n36944 );
xor ( n36946 , n36760 , n36945 );
buf ( n36947 , n35718 );
not ( n36948 , n36947 );
buf ( n36949 , n6640 );
not ( n36950 , n36949 );
or ( n36951 , n36948 , n36950 );
buf ( n36952 , n35723 );
nand ( n36953 , n36951 , n36952 );
buf ( n36954 , n36953 );
buf ( n36955 , n36954 );
xor ( n36956 , n36946 , n36955 );
buf ( n36957 , n36956 );
nand ( n36958 , n36957 , n2356 );
nand ( n36959 , n36754 , n36958 );
nand ( n36960 , n7041 , n6916 , n6851 , n6962 );
nor ( n36961 , n7046 , n7047 );
nand ( n36962 , n36961 , n6851 , n6962 );
nand ( n36963 , n36960 , n36962 );
buf ( n36964 , n36963 );
not ( n36965 , n36964 );
not ( n36966 , n36965 );
and ( n36967 , n36959 , n36966 );
not ( n36968 , n36959 );
and ( n36969 , n36968 , n36965 );
nor ( n36970 , n36967 , n36969 );
not ( n36971 , n36970 );
or ( n36972 , n7411 , n36971 );
xor ( n36973 , n36044 , n7187 );
and ( n36974 , n36973 , n7217 );
and ( n36975 , n36044 , n7187 );
or ( n36976 , n36974 , n36975 );
not ( n36977 , n2879 );
not ( n36978 , n36977 );
not ( n36979 , n32126 );
or ( n36980 , n36978 , n36979 );
nand ( n36981 , n2803 , n2879 );
nand ( n36982 , n36980 , n36981 );
nor ( n36983 , n36982 , n7151 );
not ( n36984 , n7071 );
not ( n36985 , n496 );
not ( n36986 , n7090 );
or ( n36987 , n36985 , n36986 );
not ( n36988 , n496 );
nand ( n36989 , n7074 , n36988 );
nand ( n36990 , n36987 , n36989 );
not ( n36991 , n36990 );
or ( n36992 , n36984 , n36991 );
nand ( n36993 , n7083 , n7118 );
nand ( n36994 , n36992 , n36993 );
xor ( n36995 , n36983 , n36994 );
and ( n36996 , n7204 , n7065 );
not ( n36997 , n7204 );
and ( n36998 , n36997 , n7066 );
nor ( n36999 , n36996 , n36998 );
not ( n37000 , n36999 );
not ( n37001 , n7108 );
or ( n37002 , n37000 , n37001 );
not ( n37003 , n7168 );
nand ( n37004 , n37003 , n7162 );
nand ( n37005 , n37002 , n37004 );
xor ( n37006 , n36995 , n37005 );
xor ( n37007 , n36976 , n37006 );
not ( n37008 , n7139 );
or ( n37009 , n7124 , n498 );
or ( n37010 , n7123 , n7092 );
nand ( n37011 , n37009 , n37010 );
not ( n37012 , n37011 );
or ( n37013 , n37008 , n37012 );
not ( n37014 , n36053 );
or ( n37015 , n37014 , n7299 );
nand ( n37016 , n37013 , n37015 );
or ( n37017 , n7214 , n7200 );
and ( n37018 , n35943 , n7140 );
and ( n37019 , n7062 , n500 );
nor ( n37020 , n37018 , n37019 );
or ( n37021 , n37020 , n7226 );
nand ( n37022 , n37017 , n37021 );
xor ( n37023 , n37016 , n37022 );
and ( n37024 , n35947 , n7100 );
xor ( n37025 , n37023 , n37024 );
xor ( n37026 , n37007 , n37025 );
xor ( n37027 , n7101 , n7149 );
and ( n37028 , n37027 , n7218 );
and ( n37029 , n7101 , n7149 );
or ( n37030 , n37028 , n37029 );
or ( n37031 , n37026 , n37030 );
nand ( n37032 , n37026 , n37030 );
nand ( n37033 , n37031 , n37032 );
not ( n37034 , n37033 );
not ( n37035 , n7254 );
not ( n37036 , n36259 );
or ( n37037 , n37035 , n37036 );
nand ( n37038 , n37037 , n7255 );
not ( n37039 , n37038 );
or ( n37040 , n37034 , n37039 );
or ( n37041 , n37038 , n37033 );
nand ( n37042 , n37040 , n37041 );
nand ( n37043 , n37042 , n2628 );
nand ( n37044 , n36972 , n37043 );
not ( n37045 , n7410 );
buf ( n37046 , n537 );
not ( n37047 , n37046 );
not ( n37048 , n29519 );
buf ( n37049 , n518 );
buf ( n37050 , n489 );
and ( n37051 , n37049 , n37050 );
buf ( n37052 , n37051 );
buf ( n37053 , n37052 );
buf ( n37054 , n511 );
buf ( n37055 , n495 );
xor ( n37056 , n37054 , n37055 );
buf ( n37057 , n37056 );
buf ( n37058 , n37057 );
not ( n37059 , n37058 );
buf ( n37060 , n36323 );
not ( n37061 , n37060 );
or ( n37062 , n37059 , n37061 );
buf ( n37063 , n30846 );
buf ( n37064 , n510 );
buf ( n37065 , n495 );
xor ( n37066 , n37064 , n37065 );
buf ( n37067 , n37066 );
buf ( n37068 , n37067 );
nand ( n37069 , n37063 , n37068 );
buf ( n37070 , n37069 );
buf ( n37071 , n37070 );
nand ( n37072 , n37062 , n37071 );
buf ( n37073 , n37072 );
buf ( n37074 , n37073 );
xor ( n37075 , n37053 , n37074 );
xor ( n37076 , n499 , n507 );
buf ( n37077 , n37076 );
not ( n37078 , n37077 );
buf ( n37079 , n30741 );
not ( n37080 , n37079 );
or ( n37081 , n37078 , n37080 );
buf ( n37082 , n5230 );
buf ( n37083 , n506 );
buf ( n37084 , n499 );
xor ( n37085 , n37083 , n37084 );
buf ( n37086 , n37085 );
buf ( n37087 , n37086 );
nand ( n37088 , n37082 , n37087 );
buf ( n37089 , n37088 );
buf ( n37090 , n37089 );
nand ( n37091 , n37081 , n37090 );
buf ( n37092 , n37091 );
buf ( n37093 , n37092 );
xor ( n37094 , n37075 , n37093 );
buf ( n37095 , n37094 );
buf ( n37096 , n37095 );
xor ( n37097 , n489 , n517 );
buf ( n37098 , n37097 );
not ( n37099 , n37098 );
buf ( n37100 , n5172 );
not ( n37101 , n37100 );
or ( n37102 , n37099 , n37101 );
buf ( n37103 , n4928 );
buf ( n37104 , n489 );
buf ( n37105 , n516 );
xor ( n37106 , n37104 , n37105 );
buf ( n37107 , n37106 );
buf ( n37108 , n37107 );
nand ( n37109 , n37103 , n37108 );
buf ( n37110 , n37109 );
buf ( n37111 , n37110 );
nand ( n37112 , n37102 , n37111 );
buf ( n37113 , n37112 );
buf ( n37114 , n37113 );
buf ( n37115 , n7460 );
not ( n37116 , n37115 );
buf ( n37117 , n1691 );
not ( n37118 , n37117 );
or ( n37119 , n37116 , n37118 );
buf ( n37120 , n1786 );
buf ( n37121 , n509 );
buf ( n37122 , n497 );
xor ( n37123 , n37121 , n37122 );
buf ( n37124 , n37123 );
buf ( n37125 , n37124 );
nand ( n37126 , n37120 , n37125 );
buf ( n37127 , n37126 );
buf ( n37128 , n37127 );
nand ( n37129 , n37119 , n37128 );
buf ( n37130 , n37129 );
buf ( n37131 , n37130 );
xor ( n37132 , n37114 , n37131 );
buf ( n37133 , n505 );
buf ( n37134 , n501 );
xor ( n37135 , n37133 , n37134 );
buf ( n37136 , n37135 );
buf ( n37137 , n37136 );
not ( n37138 , n37137 );
buf ( n37139 , n29640 );
not ( n37140 , n37139 );
or ( n37141 , n37138 , n37140 );
buf ( n37142 , n501 );
buf ( n37143 , n33424 );
nand ( n37144 , n37142 , n37143 );
buf ( n37145 , n37144 );
buf ( n37146 , n37145 );
nand ( n37147 , n37141 , n37146 );
buf ( n37148 , n37147 );
buf ( n37149 , n37148 );
not ( n37150 , n37149 );
buf ( n37151 , n37150 );
buf ( n37152 , n37151 );
xor ( n37153 , n37132 , n37152 );
buf ( n37154 , n37153 );
buf ( n37155 , n37154 );
xor ( n37156 , n37096 , n37155 );
xor ( n37157 , n36341 , n36354 );
and ( n37158 , n37157 , n36372 );
and ( n37159 , n36341 , n36354 );
or ( n37160 , n37158 , n37159 );
buf ( n37161 , n37160 );
buf ( n37162 , n37161 );
xor ( n37163 , n7448 , n36316 );
and ( n37164 , n37163 , n7484 );
and ( n37165 , n7448 , n36316 );
or ( n37166 , n37164 , n37165 );
buf ( n37167 , n37166 );
xor ( n37168 , n37162 , n37167 );
xor ( n37169 , n36387 , n7555 );
and ( n37170 , n37169 , n36407 );
and ( n37171 , n36387 , n7555 );
or ( n37172 , n37170 , n37171 );
buf ( n37173 , n37172 );
and ( n37174 , n37168 , n37173 );
and ( n37175 , n37162 , n37167 );
or ( n37176 , n37174 , n37175 );
buf ( n37177 , n37176 );
buf ( n37178 , n37177 );
xor ( n37179 , n37156 , n37178 );
buf ( n37180 , n37179 );
buf ( n37181 , n37180 );
buf ( n37182 , n37130 );
not ( n37183 , n37182 );
buf ( n37184 , n37183 );
buf ( n37185 , n37184 );
buf ( n37186 , n7539 );
not ( n37187 , n37186 );
buf ( n37188 , n33967 );
not ( n37189 , n37188 );
or ( n37190 , n37187 , n37189 );
buf ( n37191 , n33973 );
buf ( n37192 , n515 );
buf ( n37193 , n491 );
xor ( n37194 , n37192 , n37193 );
buf ( n37195 , n37194 );
buf ( n37196 , n37195 );
nand ( n37197 , n37191 , n37196 );
buf ( n37198 , n37197 );
buf ( n37199 , n37198 );
nand ( n37200 , n37190 , n37199 );
buf ( n37201 , n37200 );
buf ( n37202 , n37201 );
xor ( n37203 , n37185 , n37202 );
buf ( n37204 , n36389 );
not ( n37205 , n37204 );
buf ( n37206 , n4241 );
not ( n37207 , n37206 );
or ( n37208 , n37205 , n37207 );
buf ( n37209 , n4218 );
buf ( n37210 , n513 );
buf ( n37211 , n493 );
xor ( n37212 , n37210 , n37211 );
buf ( n37213 , n37212 );
buf ( n37214 , n37213 );
nand ( n37215 , n37209 , n37214 );
buf ( n37216 , n37215 );
buf ( n37217 , n37216 );
nand ( n37218 , n37208 , n37217 );
buf ( n37219 , n37218 );
buf ( n37220 , n37219 );
xor ( n37221 , n37203 , n37220 );
buf ( n37222 , n37221 );
not ( n37223 , n7532 );
not ( n37224 , n7570 );
or ( n37225 , n37223 , n37224 );
nand ( n37226 , n37225 , n7573 );
xor ( n37227 , n37222 , n37226 );
xor ( n37228 , n37162 , n37167 );
xor ( n37229 , n37228 , n37173 );
buf ( n37230 , n37229 );
and ( n37231 , n37227 , n37230 );
and ( n37232 , n37222 , n37226 );
or ( n37233 , n37231 , n37232 );
buf ( n37234 , n37233 );
xor ( n37235 , n37181 , n37234 );
xor ( n37236 , n37185 , n37202 );
and ( n37237 , n37236 , n37220 );
and ( n37238 , n37185 , n37202 );
or ( n37239 , n37237 , n37238 );
buf ( n37240 , n37239 );
buf ( n37241 , n37240 );
buf ( n37242 , n519 );
buf ( n37243 , n489 );
and ( n37244 , n37242 , n37243 );
buf ( n37245 , n37244 );
buf ( n37246 , n37245 );
buf ( n37247 , n7165 );
xor ( n37248 , n37246 , n37247 );
buf ( n37249 , n7444 );
not ( n37250 , n37249 );
buf ( n37251 , n36290 );
not ( n37252 , n37251 );
or ( n37253 , n37250 , n37252 );
xor ( n37254 , n490 , n491 );
not ( n37255 , n37254 );
buf ( n37256 , n37255 );
not ( n37257 , n37256 );
buf ( n37258 , n37097 );
nand ( n37259 , n37257 , n37258 );
buf ( n37260 , n37259 );
buf ( n37261 , n37260 );
nand ( n37262 , n37253 , n37261 );
buf ( n37263 , n37262 );
buf ( n37264 , n37263 );
and ( n37265 , n37248 , n37264 );
and ( n37266 , n37246 , n37247 );
or ( n37267 , n37265 , n37266 );
buf ( n37268 , n37267 );
buf ( n37269 , n37268 );
buf ( n37270 , n36330 );
not ( n37271 , n37270 );
buf ( n37272 , n36323 );
not ( n37273 , n37272 );
or ( n37274 , n37271 , n37273 );
buf ( n37275 , n30846 );
buf ( n37276 , n37057 );
nand ( n37277 , n37275 , n37276 );
buf ( n37278 , n37277 );
buf ( n37279 , n37278 );
nand ( n37280 , n37274 , n37279 );
buf ( n37281 , n37280 );
not ( n37282 , n37281 );
buf ( n37283 , n7563 );
not ( n37284 , n37283 );
buf ( n37285 , n30741 );
not ( n37286 , n37285 );
or ( n37287 , n37284 , n37286 );
buf ( n37288 , n5230 );
buf ( n37289 , n37076 );
nand ( n37290 , n37288 , n37289 );
buf ( n37291 , n37290 );
buf ( n37292 , n37291 );
nand ( n37293 , n37287 , n37292 );
buf ( n37294 , n37293 );
not ( n37295 , n37294 );
or ( n37296 , n37282 , n37295 );
buf ( n37297 , n37281 );
buf ( n37298 , n37294 );
nor ( n37299 , n37297 , n37298 );
buf ( n37300 , n37299 );
buf ( n37301 , n36365 );
not ( n37302 , n37301 );
buf ( n37303 , n29640 );
not ( n37304 , n37303 );
or ( n37305 , n37302 , n37304 );
buf ( n37306 , n33424 );
buf ( n37307 , n37136 );
nand ( n37308 , n37306 , n37307 );
buf ( n37309 , n37308 );
buf ( n37310 , n37309 );
nand ( n37311 , n37305 , n37310 );
buf ( n37312 , n37311 );
buf ( n37313 , n37312 );
not ( n37314 , n37313 );
buf ( n37315 , n37314 );
or ( n37316 , n37300 , n37315 );
nand ( n37317 , n37296 , n37316 );
buf ( n37318 , n37317 );
xor ( n37319 , n37269 , n37318 );
buf ( n37320 , n37124 );
not ( n37321 , n37320 );
buf ( n37322 , n7455 );
not ( n37323 , n37322 );
or ( n37324 , n37321 , n37323 );
buf ( n37325 , n1786 );
buf ( n37326 , n508 );
buf ( n37327 , n497 );
xor ( n37328 , n37326 , n37327 );
buf ( n37329 , n37328 );
buf ( n37330 , n37329 );
nand ( n37331 , n37325 , n37330 );
buf ( n37332 , n37331 );
buf ( n37333 , n37332 );
nand ( n37334 , n37324 , n37333 );
buf ( n37335 , n37334 );
buf ( n37336 , n37195 );
not ( n37337 , n37336 );
buf ( n37338 , n491 );
buf ( n37339 , n492 );
not ( n37340 , n37339 );
xor ( n37341 , n37338 , n37340 );
buf ( n37342 , n37341 );
buf ( n37343 , n37342 );
buf ( n37344 , n33357 );
nor ( n37345 , n37343 , n37344 );
buf ( n37346 , n37345 );
buf ( n37347 , n37346 );
not ( n37348 , n37347 );
or ( n37349 , n37337 , n37348 );
buf ( n37350 , n33102 );
xor ( n37351 , n491 , n514 );
buf ( n37352 , n37351 );
nand ( n37353 , n37350 , n37352 );
buf ( n37354 , n37353 );
buf ( n37355 , n37354 );
nand ( n37356 , n37349 , n37355 );
buf ( n37357 , n37356 );
xor ( n37358 , n37335 , n37357 );
not ( n37359 , n37213 );
not ( n37360 , n4387 );
or ( n37361 , n37359 , n37360 );
buf ( n37362 , n33381 );
buf ( n37363 , n512 );
buf ( n37364 , n493 );
xor ( n37365 , n37363 , n37364 );
buf ( n37366 , n37365 );
buf ( n37367 , n37366 );
nand ( n37368 , n37362 , n37367 );
buf ( n37369 , n37368 );
nand ( n37370 , n37361 , n37369 );
xor ( n37371 , n37358 , n37370 );
buf ( n37372 , n37371 );
xor ( n37373 , n37319 , n37372 );
buf ( n37374 , n37373 );
buf ( n37375 , n37374 );
xor ( n37376 , n37241 , n37375 );
xor ( n37377 , n37246 , n37247 );
xor ( n37378 , n37377 , n37264 );
buf ( n37379 , n37378 );
buf ( n37380 , n37379 );
xor ( n37381 , n37312 , n37281 );
xor ( n37382 , n37381 , n37294 );
buf ( n37383 , n37382 );
xor ( n37384 , n37380 , n37383 );
xor ( n37385 , n36437 , n36445 );
and ( n37386 , n37385 , n36452 );
and ( n37387 , n36437 , n36445 );
or ( n37388 , n37386 , n37387 );
buf ( n37389 , n37388 );
buf ( n37390 , n37389 );
and ( n37391 , n37384 , n37390 );
and ( n37392 , n37380 , n37383 );
or ( n37393 , n37391 , n37392 );
buf ( n37394 , n37393 );
buf ( n37395 , n37394 );
xor ( n37396 , n37376 , n37395 );
buf ( n37397 , n37396 );
buf ( n37398 , n37397 );
xor ( n37399 , n37235 , n37398 );
buf ( n37400 , n37399 );
not ( n37401 , n37400 );
xor ( n37402 , n37380 , n37383 );
xor ( n37403 , n37402 , n37390 );
buf ( n37404 , n37403 );
xor ( n37405 , n37222 , n37226 );
xor ( n37406 , n37405 , n37230 );
xor ( n37407 , n37404 , n37406 );
xor ( n37408 , n36434 , n36455 );
and ( n37409 , n37408 , n36462 );
and ( n37410 , n36434 , n36455 );
or ( n37411 , n37409 , n37410 );
buf ( n37412 , n37411 );
and ( n37413 , n37407 , n37412 );
and ( n37414 , n37404 , n37406 );
or ( n37415 , n37413 , n37414 );
not ( n37416 , n37415 );
nand ( n37417 , n37401 , n37416 );
nand ( n37418 , n37400 , n37415 );
nand ( n37419 , n37417 , n37418 );
buf ( n37420 , n37419 );
not ( n37421 , n37420 );
xor ( n37422 , n36421 , n36427 );
and ( n37423 , n37422 , n36465 );
and ( n37424 , n36421 , n36427 );
or ( n37425 , n37423 , n37424 );
buf ( n37426 , n37425 );
xor ( n37427 , n37404 , n37406 );
xor ( n37428 , n37427 , n37412 );
nor ( n37429 , n37426 , n37428 );
nor ( n37430 , n37429 , n36473 );
not ( n37431 , n37430 );
not ( n37432 , n7433 );
or ( n37433 , n37431 , n37432 );
nor ( n37434 , n37428 , n37426 );
or ( n37435 , n37434 , n36475 );
nand ( n37436 , n37428 , n37426 );
nand ( n37437 , n37435 , n37436 );
buf ( n37438 , n37437 );
not ( n37439 , n37438 );
nand ( n37440 , n37433 , n37439 );
not ( n37441 , n37440 );
or ( n37442 , n37421 , n37441 );
or ( n37443 , n37440 , n37420 );
nand ( n37444 , n37442 , n37443 );
not ( n37445 , n37444 );
or ( n37446 , n37048 , n37445 );
not ( n37447 , n36562 );
not ( n37448 , n499 );
not ( n37449 , n32467 );
or ( n37450 , n37448 , n37449 );
buf ( n37451 , n3434 );
buf ( n37452 , n29901 );
nand ( n37453 , n37451 , n37452 );
buf ( n37454 , n37453 );
nand ( n37455 , n37450 , n37454 );
not ( n37456 , n37455 );
or ( n37457 , n37447 , n37456 );
and ( n37458 , n456 , n458 );
not ( n37459 , n456 );
and ( n37460 , n37459 , n474 );
nor ( n37461 , n37458 , n37460 );
not ( n37462 , n37461 );
not ( n37463 , n37462 );
not ( n37464 , n29901 );
or ( n37465 , n37463 , n37464 );
nand ( n37466 , n499 , n37461 );
nand ( n37467 , n37465 , n37466 );
nand ( n37468 , n29884 , n37467 );
nand ( n37469 , n37457 , n37468 );
buf ( n37470 , n37469 );
buf ( n37471 , n29891 );
not ( n37472 , n37471 );
buf ( n37473 , n489 );
nand ( n37474 , n37472 , n37473 );
buf ( n37475 , n37474 );
buf ( n37476 , n37475 );
and ( n37477 , n37470 , n37476 );
not ( n37478 , n37470 );
buf ( n37479 , n37475 );
not ( n37480 , n37479 );
buf ( n37481 , n37480 );
buf ( n37482 , n37481 );
and ( n37483 , n37478 , n37482 );
nor ( n37484 , n37477 , n37483 );
buf ( n37485 , n37484 );
not ( n37486 , n1914 );
not ( n37487 , n495 );
not ( n37488 , n32975 );
or ( n37489 , n37487 , n37488 );
buf ( n37490 , n2803 );
buf ( n37491 , n31784 );
nand ( n37492 , n37490 , n37491 );
buf ( n37493 , n37492 );
nand ( n37494 , n37489 , n37493 );
not ( n37495 , n37494 );
or ( n37496 , n37486 , n37495 );
buf ( n37497 , n495 );
not ( n37498 , n37497 );
buf ( n37499 , n2678 );
not ( n37500 , n37499 );
or ( n37501 , n37498 , n37500 );
buf ( n37502 , n2879 );
buf ( n37503 , n31784 );
nand ( n37504 , n37502 , n37503 );
buf ( n37505 , n37504 );
buf ( n37506 , n37505 );
nand ( n37507 , n37501 , n37506 );
buf ( n37508 , n37507 );
nand ( n37509 , n37508 , n31812 );
nand ( n37510 , n37496 , n37509 );
not ( n37511 , n37510 );
and ( n37512 , n37485 , n37511 );
not ( n37513 , n37485 );
and ( n37514 , n37513 , n37510 );
nor ( n37515 , n37512 , n37514 );
buf ( n37516 , n37515 );
buf ( n37517 , n1010 );
not ( n37518 , n37517 );
buf ( n37519 , n984 );
nor ( n37520 , n37518 , n37519 );
buf ( n37521 , n37520 );
and ( n37522 , n984 , n5562 );
not ( n37523 , n984 );
and ( n37524 , n37523 , n5554 );
nor ( n37525 , n37522 , n37524 );
nor ( n37526 , n37525 , n2989 );
nor ( n37527 , n37521 , n37526 );
buf ( n37528 , n489 );
not ( n37529 , n37528 );
buf ( n37530 , n30090 );
not ( n37531 , n37530 );
or ( n37532 , n37529 , n37531 );
buf ( n37533 , n489 );
not ( n37534 , n37533 );
buf ( n37535 , n973 );
nand ( n37536 , n37534 , n37535 );
buf ( n37537 , n37536 );
buf ( n37538 , n37537 );
nand ( n37539 , n37532 , n37538 );
buf ( n37540 , n37539 );
not ( n37541 , n37540 );
not ( n37542 , n5417 );
not ( n37543 , n37542 );
or ( n37544 , n37541 , n37543 );
xor ( n37545 , n489 , n2845 );
not ( n37546 , n37545 );
nand ( n37547 , n37546 , n36508 );
nand ( n37548 , n37544 , n37547 );
xor ( n37549 , n37527 , n37548 );
not ( n37550 , n909 );
buf ( n37551 , n497 );
not ( n37552 , n37551 );
buf ( n37553 , n31829 );
not ( n37554 , n37553 );
or ( n37555 , n37552 , n37554 );
buf ( n37556 , n31826 );
buf ( n37557 , n30599 );
nand ( n37558 , n37556 , n37557 );
buf ( n37559 , n37558 );
buf ( n37560 , n37559 );
nand ( n37561 , n37555 , n37560 );
buf ( n37562 , n37561 );
not ( n37563 , n37562 );
or ( n37564 , n37550 , n37563 );
and ( n37565 , n2803 , n30599 );
not ( n37566 , n2803 );
and ( n37567 , n37566 , n497 );
or ( n37568 , n37565 , n37567 );
buf ( n37569 , n37568 );
buf ( n37570 , n30585 );
nand ( n37571 , n37569 , n37570 );
buf ( n37572 , n37571 );
nand ( n37573 , n37564 , n37572 );
xor ( n37574 , n37549 , n37573 );
buf ( n37575 , n37574 );
xor ( n37576 , n37516 , n37575 );
xor ( n37577 , n36526 , n36539 );
and ( n37578 , n37577 , n36556 );
and ( n37579 , n36526 , n36539 );
or ( n37580 , n37578 , n37579 );
buf ( n37581 , n37580 );
buf ( n37582 , n37581 );
xor ( n37583 , n36583 , n36600 );
and ( n37584 , n37583 , n36618 );
and ( n37585 , n36583 , n36600 );
or ( n37586 , n37584 , n37585 );
buf ( n37587 , n37586 );
xor ( n37588 , n37582 , n37587 );
xor ( n37589 , n36494 , n36506 );
and ( n37590 , n37589 , n36518 );
and ( n37591 , n36494 , n36506 );
or ( n37592 , n37590 , n37591 );
buf ( n37593 , n37592 );
and ( n37594 , n37588 , n37593 );
and ( n37595 , n37582 , n37587 );
or ( n37596 , n37594 , n37595 );
buf ( n37597 , n37596 );
buf ( n37598 , n37597 );
xor ( n37599 , n37576 , n37598 );
buf ( n37600 , n37599 );
buf ( n37601 , n37600 );
buf ( n37602 , n3146 );
not ( n37603 , n37602 );
buf ( n37604 , n36608 );
not ( n37605 , n37604 );
or ( n37606 , n37603 , n37605 );
not ( n37607 , n493 );
not ( n37608 , n3597 );
or ( n37609 , n37607 , n37608 );
or ( n37610 , n3597 , n493 );
nand ( n37611 , n37609 , n37610 );
nand ( n37612 , n2978 , n37611 );
buf ( n37613 , n37612 );
nand ( n37614 , n37606 , n37613 );
buf ( n37615 , n37614 );
buf ( n37616 , n37615 );
buf ( n37617 , n34465 );
not ( n37618 , n37617 );
buf ( n37619 , n36596 );
not ( n37620 , n37619 );
or ( n37621 , n37618 , n37620 );
buf ( n37622 , n491 );
not ( n37623 , n37622 );
buf ( n37624 , n882 );
not ( n37625 , n37624 );
or ( n37626 , n37623 , n37625 );
buf ( n37627 , n30008 );
buf ( n37628 , n3524 );
nand ( n37629 , n37627 , n37628 );
buf ( n37630 , n37629 );
buf ( n37631 , n37630 );
nand ( n37632 , n37626 , n37631 );
buf ( n37633 , n37632 );
buf ( n37634 , n37633 );
buf ( n37635 , n3045 );
nand ( n37636 , n37634 , n37635 );
buf ( n37637 , n37636 );
buf ( n37638 , n37637 );
nand ( n37639 , n37621 , n37638 );
buf ( n37640 , n37639 );
buf ( n37641 , n37640 );
xor ( n37642 , n37616 , n37641 );
buf ( n37643 , n37573 );
not ( n37644 , n37643 );
buf ( n37645 , n37644 );
buf ( n37646 , n37645 );
xor ( n37647 , n37642 , n37646 );
buf ( n37648 , n37647 );
not ( n37649 , n36519 );
not ( n37650 , n36629 );
or ( n37651 , n37649 , n37650 );
nand ( n37652 , n37651 , n36625 );
xor ( n37653 , n37648 , n37652 );
xor ( n37654 , n37582 , n37587 );
xor ( n37655 , n37654 , n37593 );
buf ( n37656 , n37655 );
and ( n37657 , n37653 , n37656 );
and ( n37658 , n37648 , n37652 );
or ( n37659 , n37657 , n37658 );
buf ( n37660 , n37659 );
xor ( n37661 , n37601 , n37660 );
xor ( n37662 , n37616 , n37641 );
and ( n37663 , n37662 , n37646 );
and ( n37664 , n37616 , n37641 );
or ( n37665 , n37663 , n37664 );
buf ( n37666 , n37665 );
buf ( n37667 , n37666 );
not ( n37668 , n29987 );
buf ( n37669 , n489 );
not ( n37670 , n37669 );
buf ( n37671 , n31951 );
nor ( n37672 , n37670 , n37671 );
buf ( n37673 , n37672 );
not ( n37674 , n37673 );
nand ( n37675 , n37668 , n37674 );
not ( n37676 , n37675 );
not ( n37677 , n5417 );
not ( n37678 , n37677 );
not ( n37679 , n36511 );
or ( n37680 , n37678 , n37679 );
buf ( n37681 , n37540 );
buf ( n37682 , n36508 );
nand ( n37683 , n37681 , n37682 );
buf ( n37684 , n37683 );
nand ( n37685 , n37680 , n37684 );
not ( n37686 , n37685 );
or ( n37687 , n37676 , n37686 );
nand ( n37688 , n37673 , n29987 );
nand ( n37689 , n37687 , n37688 );
not ( n37690 , n29884 );
not ( n37691 , n37455 );
or ( n37692 , n37690 , n37691 );
nand ( n37693 , n36579 , n799 );
nand ( n37694 , n37692 , n37693 );
not ( n37695 , n37694 );
buf ( n37696 , n31812 );
not ( n37697 , n37696 );
buf ( n37698 , n36501 );
not ( n37699 , n37698 );
or ( n37700 , n37697 , n37699 );
nand ( n37701 , n37508 , n2725 );
buf ( n37702 , n37701 );
nand ( n37703 , n37700 , n37702 );
buf ( n37704 , n37703 );
not ( n37705 , n37704 );
or ( n37706 , n37695 , n37705 );
buf ( n37707 , n37694 );
not ( n37708 , n31812 );
not ( n37709 , n36501 );
or ( n37710 , n37708 , n37709 );
nand ( n37711 , n37710 , n37701 );
buf ( n37712 , n37711 );
nor ( n37713 , n37707 , n37712 );
buf ( n37714 , n37713 );
not ( n37715 , n36548 );
not ( n37716 , n32034 );
or ( n37717 , n37715 , n37716 );
and ( n37718 , n503 , n953 );
not ( n37719 , n37718 );
not ( n37720 , n37719 );
not ( n37721 , n957 );
or ( n37722 , n37720 , n37721 );
not ( n37723 , n37525 );
nand ( n37724 , n37722 , n37723 );
nand ( n37725 , n37717 , n37724 );
buf ( n37726 , n37725 );
not ( n37727 , n37726 );
buf ( n37728 , n37727 );
or ( n37729 , n37714 , n37728 );
nand ( n37730 , n37706 , n37729 );
xor ( n37731 , n37689 , n37730 );
not ( n37732 , n3511 );
not ( n37733 , n37611 );
or ( n37734 , n37732 , n37733 );
buf ( n37735 , n493 );
not ( n37736 , n37735 );
buf ( n37737 , n1883 );
not ( n37738 , n37737 );
or ( n37739 , n37736 , n37738 );
buf ( n37740 , n29501 );
buf ( n37741 , n2704 );
nand ( n37742 , n37740 , n37741 );
buf ( n37743 , n37742 );
buf ( n37744 , n37743 );
nand ( n37745 , n37739 , n37744 );
buf ( n37746 , n37745 );
nand ( n37747 , n37746 , n2978 );
nand ( n37748 , n37734 , n37747 );
buf ( n37749 , n3948 );
not ( n37750 , n37749 );
buf ( n37751 , n37633 );
not ( n37752 , n37751 );
or ( n37753 , n37750 , n37752 );
not ( n37754 , n491 );
not ( n37755 , n933 );
or ( n37756 , n37754 , n37755 );
nand ( n37757 , n2944 , n3524 );
nand ( n37758 , n37756 , n37757 );
buf ( n37759 , n37758 );
not ( n37760 , n37759 );
buf ( n37761 , n3045 );
nand ( n37762 , n37760 , n37761 );
buf ( n37763 , n37762 );
buf ( n37764 , n37763 );
nand ( n37765 , n37753 , n37764 );
buf ( n37766 , n37765 );
xor ( n37767 , n37748 , n37766 );
buf ( n37768 , n910 );
not ( n37769 , n37768 );
buf ( n37770 , n497 );
not ( n37771 , n37770 );
buf ( n37772 , n3211 );
not ( n37773 , n37772 );
or ( n37774 , n37771 , n37773 );
buf ( n37775 , n3220 );
buf ( n37776 , n30599 );
nand ( n37777 , n37775 , n37776 );
buf ( n37778 , n37777 );
buf ( n37779 , n37778 );
nand ( n37780 , n37774 , n37779 );
buf ( n37781 , n37780 );
buf ( n37782 , n37781 );
not ( n37783 , n37782 );
or ( n37784 , n37769 , n37783 );
buf ( n37785 , n37562 );
buf ( n37786 , n30585 );
nand ( n37787 , n37785 , n37786 );
buf ( n37788 , n37787 );
buf ( n37789 , n37788 );
nand ( n37790 , n37784 , n37789 );
buf ( n37791 , n37790 );
xor ( n37792 , n37767 , n37791 );
xor ( n37793 , n37731 , n37792 );
buf ( n37794 , n37793 );
xor ( n37795 , n37667 , n37794 );
xor ( n37796 , n37674 , n29987 );
not ( n37797 , n37685 );
xor ( n37798 , n37796 , n37797 );
buf ( n37799 , n37798 );
not ( n37800 , n37711 );
not ( n37801 , n37800 );
not ( n37802 , n37725 );
not ( n37803 , n37694 );
not ( n37804 , n37803 );
or ( n37805 , n37802 , n37804 );
or ( n37806 , n37803 , n37725 );
nand ( n37807 , n37805 , n37806 );
not ( n37808 , n37807 );
or ( n37809 , n37801 , n37808 );
or ( n37810 , n37807 , n37800 );
nand ( n37811 , n37809 , n37810 );
buf ( n37812 , n37811 );
xor ( n37813 , n37799 , n37812 );
xor ( n37814 , n36647 , n36667 );
and ( n37815 , n37814 , n36674 );
and ( n37816 , n36647 , n36667 );
or ( n37817 , n37815 , n37816 );
buf ( n37818 , n37817 );
buf ( n37819 , n37818 );
and ( n37820 , n37813 , n37819 );
and ( n37821 , n37799 , n37812 );
or ( n37822 , n37820 , n37821 );
buf ( n37823 , n37822 );
buf ( n37824 , n37823 );
xor ( n37825 , n37795 , n37824 );
buf ( n37826 , n37825 );
buf ( n37827 , n37826 );
xor ( n37828 , n37661 , n37827 );
buf ( n37829 , n37828 );
not ( n37830 , n37829 );
xor ( n37831 , n37799 , n37812 );
xor ( n37832 , n37831 , n37819 );
buf ( n37833 , n37832 );
xor ( n37834 , n37648 , n37652 );
xor ( n37835 , n37834 , n37656 );
xor ( n37836 , n37833 , n37835 );
xor ( n37837 , n36645 , n36677 );
and ( n37838 , n37837 , n36684 );
and ( n37839 , n36645 , n36677 );
or ( n37840 , n37838 , n37839 );
buf ( n37841 , n37840 );
and ( n37842 , n37836 , n37841 );
and ( n37843 , n37833 , n37835 );
or ( n37844 , n37842 , n37843 );
not ( n37845 , n37844 );
nand ( n37846 , n37830 , n37845 );
not ( n37847 , n37846 );
not ( n37848 , n37847 );
nand ( n37849 , n37829 , n37844 );
nand ( n37850 , n37848 , n37849 );
not ( n37851 , n37850 );
not ( n37852 , n37851 );
xor ( n37853 , n37833 , n37835 );
xor ( n37854 , n37853 , n37841 );
xor ( n37855 , n36633 , n36639 );
and ( n37856 , n37855 , n36687 );
and ( n37857 , n36633 , n36639 );
or ( n37858 , n37856 , n37857 );
buf ( n37859 , n37858 );
nor ( n37860 , n37854 , n37859 );
or ( n37861 , n37860 , n36697 );
nand ( n37862 , n37854 , n37859 );
nand ( n37863 , n37861 , n37862 );
buf ( n37864 , n37863 );
not ( n37865 , n37864 );
nor ( n37866 , n37859 , n37854 );
nor ( n37867 , n37866 , n36695 );
buf ( n37868 , n37867 );
nand ( n37869 , n36713 , n37868 );
nand ( n37870 , n37865 , n37869 );
not ( n37871 , n37870 );
or ( n37872 , n37852 , n37871 );
and ( n37873 , n37869 , n37865 , n37850 );
not ( n37874 , n455 );
nor ( n37875 , n37873 , n37874 );
nand ( n37876 , n37872 , n37875 );
nand ( n37877 , n37446 , n37876 );
buf ( n37878 , n37877 );
not ( n37879 , n37878 );
or ( n37880 , n37047 , n37879 );
buf ( n37881 , n37877 );
not ( n37882 , n37881 );
buf ( n37883 , n537 );
not ( n37884 , n37883 );
buf ( n37885 , n37884 );
buf ( n37886 , n37885 );
nand ( n37887 , n37882 , n37886 );
buf ( n37888 , n37887 );
buf ( n37889 , n37888 );
nand ( n37890 , n37880 , n37889 );
buf ( n37891 , n37890 );
not ( n37892 , n36474 );
not ( n37893 , n7433 );
or ( n37894 , n37892 , n37893 );
buf ( n37895 , n36475 );
nand ( n37896 , n37894 , n37895 );
not ( n37897 , n37429 );
nand ( n37898 , n37897 , n37436 );
and ( n37899 , n37898 , n29519 );
and ( n37900 , n37896 , n37899 );
not ( n37901 , n37896 );
not ( n37902 , n29519 );
nor ( n37903 , n37902 , n37898 );
and ( n37904 , n37901 , n37903 );
nor ( n37905 , n37900 , n37904 );
not ( n37906 , n36696 );
not ( n37907 , n36713 );
or ( n37908 , n37906 , n37907 );
nand ( n37909 , n37908 , n36698 );
not ( n37910 , n37909 );
not ( n37911 , n37866 );
nand ( n37912 , n37911 , n37862 );
not ( n37913 , n37912 );
nand ( n37914 , n37913 , n455 );
not ( n37915 , n37914 );
nand ( n37916 , n37910 , n37915 );
and ( n37917 , n37912 , n455 );
nand ( n37918 , n37909 , n37917 );
buf ( n37919 , n538 );
not ( n37920 , n37919 );
buf ( n37921 , n37920 );
nand ( n37922 , n37905 , n37916 , n37918 , n37921 );
buf ( n37923 , n37922 );
buf ( n37924 , n37923 );
buf ( n37925 , n37924 );
nor ( n37926 , n37891 , n37925 );
not ( n37927 , n37926 );
not ( n37928 , n37927 );
not ( n37929 , n7412 );
not ( n37930 , n36728 );
or ( n37931 , n37929 , n37930 );
nand ( n37932 , n37931 , n5659 );
not ( n37933 , n538 );
nand ( n37934 , n37905 , n37916 , n37918 );
not ( n37935 , n37934 );
or ( n37936 , n37933 , n37935 );
nand ( n37937 , n37916 , n37905 , n37918 , n37921 );
nand ( n37938 , n37936 , n37937 );
not ( n37939 , n37938 );
buf ( n37940 , n36725 );
not ( n37941 , n37940 );
buf ( n37942 , n37941 );
nand ( n37943 , n37939 , n37942 );
or ( n37944 , n36728 , n7412 );
nand ( n37945 , n37932 , n37943 , n37944 );
buf ( n37946 , n37891 );
buf ( n37947 , n37925 );
nand ( n37948 , n37946 , n37947 );
buf ( n37949 , n37948 );
buf ( n37950 , n37938 );
buf ( n37951 , n37950 );
buf ( n37952 , n36725 );
nand ( n37953 , n37951 , n37952 );
buf ( n37954 , n37953 );
nand ( n37955 , n37945 , n37949 , n37954 );
not ( n37956 , n37955 );
or ( n37957 , n37928 , n37956 );
not ( n37958 , n5661 );
nand ( n37959 , n36732 , n37958 );
not ( n37960 , n37959 );
not ( n37961 , n37938 );
nand ( n37962 , n37961 , n37942 );
not ( n37963 , n37962 );
nor ( n37964 , n37926 , n37963 );
nand ( n37965 , n34925 , n37960 , n37964 );
nand ( n37966 , n37957 , n37965 );
buf ( n37967 , n37966 );
not ( n37968 , n37967 );
not ( n37969 , n29519 );
not ( n37970 , n7433 );
xor ( n37971 , n37114 , n37131 );
and ( n37972 , n37971 , n37152 );
and ( n37973 , n37114 , n37131 );
or ( n37974 , n37972 , n37973 );
buf ( n37975 , n37974 );
buf ( n37976 , n37975 );
buf ( n37977 , n517 );
buf ( n37978 , n489 );
and ( n37979 , n37977 , n37978 );
buf ( n37980 , n37979 );
buf ( n37981 , n37980 );
buf ( n37982 , n37329 );
not ( n37983 , n37982 );
buf ( n37984 , n7455 );
not ( n37985 , n37984 );
or ( n37986 , n37983 , n37985 );
buf ( n37987 , n1786 );
buf ( n37988 , n507 );
buf ( n37989 , n497 );
xor ( n37990 , n37988 , n37989 );
buf ( n37991 , n37990 );
buf ( n37992 , n37991 );
nand ( n37993 , n37987 , n37992 );
buf ( n37994 , n37993 );
buf ( n37995 , n37994 );
nand ( n37996 , n37986 , n37995 );
buf ( n37997 , n37996 );
buf ( n37998 , n37997 );
xor ( n37999 , n37981 , n37998 );
buf ( n38000 , n37366 );
not ( n38001 , n38000 );
buf ( n38002 , n4241 );
not ( n38003 , n38002 );
or ( n38004 , n38001 , n38003 );
buf ( n38005 , n4218 );
xor ( n38006 , n493 , n511 );
buf ( n38007 , n38006 );
nand ( n38008 , n38005 , n38007 );
buf ( n38009 , n38008 );
buf ( n38010 , n38009 );
nand ( n38011 , n38004 , n38010 );
buf ( n38012 , n38011 );
buf ( n38013 , n38012 );
xor ( n38014 , n37999 , n38013 );
buf ( n38015 , n38014 );
buf ( n38016 , n38015 );
xor ( n38017 , n37976 , n38016 );
buf ( n38018 , n37151 );
not ( n38019 , n38018 );
buf ( n38020 , n37107 );
not ( n38021 , n38020 );
buf ( n38022 , n36290 );
not ( n38023 , n38022 );
or ( n38024 , n38021 , n38023 );
buf ( n38025 , n4928 );
buf ( n38026 , n489 );
buf ( n38027 , n515 );
xor ( n38028 , n38026 , n38027 );
buf ( n38029 , n38028 );
buf ( n38030 , n38029 );
nand ( n38031 , n38025 , n38030 );
buf ( n38032 , n38031 );
buf ( n38033 , n38032 );
nand ( n38034 , n38024 , n38033 );
buf ( n38035 , n38034 );
buf ( n38036 , n37351 );
not ( n38037 , n38036 );
buf ( n38038 , n4370 );
not ( n38039 , n38038 );
or ( n38040 , n38037 , n38039 );
buf ( n38041 , n33102 );
buf ( n38042 , n513 );
buf ( n38043 , n491 );
xor ( n38044 , n38042 , n38043 );
buf ( n38045 , n38044 );
buf ( n38046 , n38045 );
nand ( n38047 , n38041 , n38046 );
buf ( n38048 , n38047 );
buf ( n38049 , n38048 );
nand ( n38050 , n38040 , n38049 );
buf ( n38051 , n38050 );
xor ( n38052 , n38035 , n38051 );
buf ( n38053 , n38052 );
not ( n38054 , n38053 );
or ( n38055 , n38019 , n38054 );
buf ( n38056 , n38052 );
buf ( n38057 , n37151 );
or ( n38058 , n38056 , n38057 );
nand ( n38059 , n38055 , n38058 );
buf ( n38060 , n38059 );
buf ( n38061 , n38060 );
xor ( n38062 , n38017 , n38061 );
buf ( n38063 , n38062 );
buf ( n38064 , n38063 );
xor ( n38065 , n37241 , n37375 );
and ( n38066 , n38065 , n37395 );
and ( n38067 , n37241 , n37375 );
or ( n38068 , n38066 , n38067 );
buf ( n38069 , n38068 );
buf ( n38070 , n38069 );
xor ( n38071 , n38064 , n38070 );
xor ( n38072 , n37269 , n37318 );
and ( n38073 , n38072 , n37372 );
and ( n38074 , n37269 , n37318 );
or ( n38075 , n38073 , n38074 );
buf ( n38076 , n38075 );
buf ( n38077 , n38076 );
buf ( n38078 , n37357 );
not ( n38079 , n38078 );
buf ( n38080 , n37370 );
not ( n38081 , n38080 );
or ( n38082 , n38079 , n38081 );
buf ( n38083 , n37370 );
buf ( n38084 , n37357 );
or ( n38085 , n38083 , n38084 );
buf ( n38086 , n37335 );
nand ( n38087 , n38085 , n38086 );
buf ( n38088 , n38087 );
buf ( n38089 , n38088 );
nand ( n38090 , n38082 , n38089 );
buf ( n38091 , n38090 );
buf ( n38092 , n38091 );
xor ( n38093 , n37053 , n37074 );
and ( n38094 , n38093 , n37093 );
and ( n38095 , n37053 , n37074 );
or ( n38096 , n38094 , n38095 );
buf ( n38097 , n38096 );
buf ( n38098 , n38097 );
xor ( n38099 , n38092 , n38098 );
buf ( n38100 , n29646 );
not ( n38101 , n38100 );
buf ( n38102 , n38101 );
buf ( n38103 , n38102 );
not ( n38104 , n38103 );
buf ( n38105 , n33914 );
not ( n38106 , n38105 );
or ( n38107 , n38104 , n38106 );
buf ( n38108 , n501 );
nand ( n38109 , n38107 , n38108 );
buf ( n38110 , n38109 );
buf ( n38111 , n38110 );
buf ( n38112 , n37067 );
not ( n38113 , n38112 );
buf ( n38114 , n36323 );
not ( n38115 , n38114 );
or ( n38116 , n38113 , n38115 );
buf ( n38117 , n30846 );
buf ( n38118 , n509 );
buf ( n38119 , n495 );
xor ( n38120 , n38118 , n38119 );
buf ( n38121 , n38120 );
buf ( n38122 , n38121 );
nand ( n38123 , n38117 , n38122 );
buf ( n38124 , n38123 );
buf ( n38125 , n38124 );
nand ( n38126 , n38116 , n38125 );
buf ( n38127 , n38126 );
buf ( n38128 , n38127 );
xor ( n38129 , n38111 , n38128 );
buf ( n38130 , n37086 );
not ( n38131 , n38130 );
buf ( n38132 , n29535 );
not ( n38133 , n38132 );
or ( n38134 , n38131 , n38133 );
buf ( n38135 , n5230 );
buf ( n38136 , n505 );
buf ( n38137 , n499 );
xor ( n38138 , n38136 , n38137 );
buf ( n38139 , n38138 );
buf ( n38140 , n38139 );
nand ( n38141 , n38135 , n38140 );
buf ( n38142 , n38141 );
buf ( n38143 , n38142 );
nand ( n38144 , n38134 , n38143 );
buf ( n38145 , n38144 );
buf ( n38146 , n38145 );
xor ( n38147 , n38129 , n38146 );
buf ( n38148 , n38147 );
buf ( n38149 , n38148 );
xor ( n38150 , n38099 , n38149 );
buf ( n38151 , n38150 );
buf ( n38152 , n38151 );
xor ( n38153 , n38077 , n38152 );
xor ( n38154 , n37096 , n37155 );
and ( n38155 , n38154 , n37178 );
and ( n38156 , n37096 , n37155 );
or ( n38157 , n38155 , n38156 );
buf ( n38158 , n38157 );
buf ( n38159 , n38158 );
xor ( n38160 , n38153 , n38159 );
buf ( n38161 , n38160 );
buf ( n38162 , n38161 );
xor ( n38163 , n38071 , n38162 );
buf ( n38164 , n38163 );
not ( n38165 , n38164 );
xor ( n38166 , n37181 , n37234 );
and ( n38167 , n38166 , n37398 );
and ( n38168 , n37181 , n37234 );
or ( n38169 , n38167 , n38168 );
buf ( n38170 , n38169 );
not ( n38171 , n38170 );
nand ( n38172 , n38165 , n38171 );
nand ( n38173 , n37430 , n38172 , n37417 );
not ( n38174 , n38173 );
not ( n38175 , n38174 );
or ( n38176 , n37970 , n38175 );
not ( n38177 , n37417 );
nor ( n38178 , n38164 , n38170 );
nor ( n38179 , n38177 , n38178 );
and ( n38180 , n37438 , n38179 );
not ( n38181 , n37418 );
not ( n38182 , n38181 );
not ( n38183 , n38172 );
or ( n38184 , n38182 , n38183 );
nand ( n38185 , n38164 , n38170 );
nand ( n38186 , n38184 , n38185 );
nor ( n38187 , n38180 , n38186 );
nand ( n38188 , n38176 , n38187 );
xor ( n38189 , n38064 , n38070 );
and ( n38190 , n38189 , n38162 );
and ( n38191 , n38064 , n38070 );
or ( n38192 , n38190 , n38191 );
buf ( n38193 , n38192 );
not ( n38194 , n38193 );
xor ( n38195 , n37976 , n38016 );
and ( n38196 , n38195 , n38061 );
and ( n38197 , n37976 , n38016 );
or ( n38198 , n38196 , n38197 );
buf ( n38199 , n38198 );
buf ( n38200 , n38199 );
xor ( n38201 , n38077 , n38152 );
and ( n38202 , n38201 , n38159 );
and ( n38203 , n38077 , n38152 );
or ( n38204 , n38202 , n38203 );
buf ( n38205 , n38204 );
buf ( n38206 , n38205 );
xor ( n38207 , n38200 , n38206 );
buf ( n38208 , n38139 );
not ( n38209 , n38208 );
buf ( n38210 , n30741 );
not ( n38211 , n38210 );
or ( n38212 , n38209 , n38211 );
buf ( n38213 , n499 );
buf ( n38214 , n5230 );
nand ( n38215 , n38213 , n38214 );
buf ( n38216 , n38215 );
buf ( n38217 , n38216 );
nand ( n38218 , n38212 , n38217 );
buf ( n38219 , n38218 );
not ( n38220 , n38219 );
buf ( n38221 , n38220 );
xor ( n38222 , n37981 , n37998 );
and ( n38223 , n38222 , n38013 );
and ( n38224 , n37981 , n37998 );
or ( n38225 , n38223 , n38224 );
buf ( n38226 , n38225 );
buf ( n38227 , n38226 );
xor ( n38228 , n38221 , n38227 );
xor ( n38229 , n38111 , n38128 );
and ( n38230 , n38229 , n38146 );
and ( n38231 , n38111 , n38128 );
or ( n38232 , n38230 , n38231 );
buf ( n38233 , n38232 );
buf ( n38234 , n38233 );
xor ( n38235 , n38228 , n38234 );
buf ( n38236 , n38235 );
buf ( n38237 , n38236 );
xor ( n38238 , n38092 , n38098 );
and ( n38239 , n38238 , n38149 );
and ( n38240 , n38092 , n38098 );
or ( n38241 , n38239 , n38240 );
buf ( n38242 , n38241 );
buf ( n38243 , n38242 );
xor ( n38244 , n38237 , n38243 );
buf ( n38245 , n38035 );
buf ( n38246 , n38051 );
or ( n38247 , n38245 , n38246 );
buf ( n38248 , n37148 );
nand ( n38249 , n38247 , n38248 );
buf ( n38250 , n38249 );
buf ( n38251 , n38250 );
buf ( n38252 , n38035 );
buf ( n38253 , n38051 );
nand ( n38254 , n38252 , n38253 );
buf ( n38255 , n38254 );
buf ( n38256 , n38255 );
nand ( n38257 , n38251 , n38256 );
buf ( n38258 , n38257 );
buf ( n38259 , n38258 );
not ( n38260 , n38045 );
not ( n38261 , n37346 );
or ( n38262 , n38260 , n38261 );
buf ( n38263 , n512 );
buf ( n38264 , n491 );
xor ( n38265 , n38263 , n38264 );
buf ( n38266 , n38265 );
nand ( n38267 , n38266 , n33102 );
nand ( n38268 , n38262 , n38267 );
buf ( n38269 , n38268 );
buf ( n38270 , n37991 );
not ( n38271 , n38270 );
buf ( n38272 , n7455 );
not ( n38273 , n38272 );
or ( n38274 , n38271 , n38273 );
buf ( n38275 , n1786 );
buf ( n38276 , n506 );
buf ( n38277 , n497 );
xor ( n38278 , n38276 , n38277 );
buf ( n38279 , n38278 );
buf ( n38280 , n38279 );
nand ( n38281 , n38275 , n38280 );
buf ( n38282 , n38281 );
buf ( n38283 , n38282 );
nand ( n38284 , n38274 , n38283 );
buf ( n38285 , n38284 );
buf ( n38286 , n38285 );
xor ( n38287 , n38269 , n38286 );
buf ( n38288 , n38006 );
not ( n38289 , n38288 );
buf ( n38290 , n4241 );
not ( n38291 , n38290 );
or ( n38292 , n38289 , n38291 );
buf ( n38293 , n4218 );
buf ( n38294 , n510 );
buf ( n38295 , n493 );
xor ( n38296 , n38294 , n38295 );
buf ( n38297 , n38296 );
buf ( n38298 , n38297 );
nand ( n38299 , n38293 , n38298 );
buf ( n38300 , n38299 );
buf ( n38301 , n38300 );
nand ( n38302 , n38292 , n38301 );
buf ( n38303 , n38302 );
buf ( n38304 , n38303 );
xor ( n38305 , n38287 , n38304 );
buf ( n38306 , n38305 );
buf ( n38307 , n38306 );
xor ( n38308 , n38259 , n38307 );
and ( n38309 , n37104 , n37105 );
buf ( n38310 , n38309 );
buf ( n38311 , n38310 );
buf ( n38312 , n38029 );
not ( n38313 , n38312 );
buf ( n38314 , n5172 );
not ( n38315 , n38314 );
or ( n38316 , n38313 , n38315 );
buf ( n38317 , n37254 );
buf ( n38318 , n489 );
buf ( n38319 , n514 );
xor ( n38320 , n38318 , n38319 );
buf ( n38321 , n38320 );
buf ( n38322 , n38321 );
nand ( n38323 , n38317 , n38322 );
buf ( n38324 , n38323 );
buf ( n38325 , n38324 );
nand ( n38326 , n38316 , n38325 );
buf ( n38327 , n38326 );
buf ( n38328 , n38327 );
xor ( n38329 , n38311 , n38328 );
buf ( n38330 , n38121 );
not ( n38331 , n38330 );
buf ( n38332 , n33757 );
not ( n38333 , n38332 );
or ( n38334 , n38331 , n38333 );
buf ( n38335 , n33167 );
buf ( n38336 , n508 );
buf ( n38337 , n495 );
xor ( n38338 , n38336 , n38337 );
buf ( n38339 , n38338 );
buf ( n38340 , n38339 );
nand ( n38341 , n38335 , n38340 );
buf ( n38342 , n38341 );
buf ( n38343 , n38342 );
nand ( n38344 , n38334 , n38343 );
buf ( n38345 , n38344 );
buf ( n38346 , n38345 );
xor ( n38347 , n38329 , n38346 );
buf ( n38348 , n38347 );
buf ( n38349 , n38348 );
xor ( n38350 , n38308 , n38349 );
buf ( n38351 , n38350 );
buf ( n38352 , n38351 );
xor ( n38353 , n38244 , n38352 );
buf ( n38354 , n38353 );
buf ( n38355 , n38354 );
xor ( n38356 , n38207 , n38355 );
buf ( n38357 , n38356 );
not ( n38358 , n38357 );
nand ( n38359 , n38194 , n38358 );
nand ( n38360 , n38357 , n38193 );
nand ( n38361 , n38359 , n38360 );
xnor ( n38362 , n38188 , n38361 );
not ( n38363 , n38362 );
or ( n38364 , n37969 , n38363 );
not ( n38365 , n5881 );
not ( n38366 , n36704 );
or ( n38367 , n38365 , n38366 );
nand ( n38368 , n38367 , n36712 );
not ( n38369 , n38368 );
xor ( n38370 , n37527 , n37548 );
and ( n38371 , n38370 , n37573 );
and ( n38372 , n37527 , n37548 );
or ( n38373 , n38371 , n38372 );
buf ( n38374 , n38373 );
buf ( n38375 , n30096 );
buf ( n38376 , n489 );
and ( n38377 , n38375 , n38376 );
buf ( n38378 , n38377 );
buf ( n38379 , n38378 );
not ( n38380 , n3146 );
not ( n38381 , n37746 );
or ( n38382 , n38380 , n38381 );
buf ( n38383 , n493 );
not ( n38384 , n38383 );
buf ( n38385 , n2678 );
not ( n38386 , n38385 );
or ( n38387 , n38384 , n38386 );
and ( n38388 , n456 , n463 );
not ( n38389 , n456 );
and ( n38390 , n38389 , n479 );
or ( n38391 , n38388 , n38390 );
nand ( n38392 , n38391 , n2704 );
buf ( n38393 , n38392 );
nand ( n38394 , n38387 , n38393 );
buf ( n38395 , n38394 );
nand ( n38396 , n38395 , n2978 );
nand ( n38397 , n38382 , n38396 );
buf ( n38398 , n38397 );
xor ( n38399 , n38379 , n38398 );
buf ( n38400 , n30585 );
not ( n38401 , n38400 );
buf ( n38402 , n37781 );
not ( n38403 , n38402 );
or ( n38404 , n38401 , n38403 );
buf ( n38405 , n497 );
not ( n38406 , n38405 );
and ( n38407 , n456 , n459 );
not ( n38408 , n456 );
and ( n38409 , n38408 , n475 );
nor ( n38410 , n38407 , n38409 );
buf ( n38411 , n38410 );
not ( n38412 , n38411 );
or ( n38413 , n38406 , n38412 );
not ( n38414 , n3433 );
buf ( n38415 , n38414 );
buf ( n38416 , n30599 );
nand ( n38417 , n38415 , n38416 );
buf ( n38418 , n38417 );
buf ( n38419 , n38418 );
nand ( n38420 , n38413 , n38419 );
buf ( n38421 , n38420 );
buf ( n38422 , n38421 );
buf ( n38423 , n910 );
nand ( n38424 , n38422 , n38423 );
buf ( n38425 , n38424 );
buf ( n38426 , n38425 );
nand ( n38427 , n38404 , n38426 );
buf ( n38428 , n38427 );
buf ( n38429 , n38428 );
xor ( n38430 , n38399 , n38429 );
buf ( n38431 , n38430 );
buf ( n38432 , n38431 );
xor ( n38433 , n38374 , n38432 );
buf ( n38434 , n37545 );
not ( n38435 , n38434 );
buf ( n38436 , n37677 );
not ( n38437 , n38436 );
buf ( n38438 , n38437 );
buf ( n38439 , n38438 );
not ( n38440 , n38439 );
and ( n38441 , n38435 , n38440 );
xor ( n38442 , n489 , n2831 );
buf ( n38443 , n38442 );
buf ( n38444 , n36508 );
and ( n38445 , n38443 , n38444 );
nor ( n38446 , n38441 , n38445 );
buf ( n38447 , n38446 );
buf ( n38448 , n38447 );
not ( n38449 , n38448 );
buf ( n38450 , n38449 );
not ( n38451 , n38450 );
not ( n38452 , n3045 );
buf ( n38453 , n491 );
not ( n38454 , n38453 );
buf ( n38455 , n30496 );
not ( n38456 , n38455 );
or ( n38457 , n38454 , n38456 );
buf ( n38458 , n1403 );
buf ( n38459 , n3524 );
nand ( n38460 , n38458 , n38459 );
buf ( n38461 , n38460 );
buf ( n38462 , n38461 );
nand ( n38463 , n38457 , n38462 );
buf ( n38464 , n38463 );
not ( n38465 , n38464 );
or ( n38466 , n38452 , n38465 );
not ( n38467 , n37758 );
not ( n38468 , n3554 );
nand ( n38469 , n38467 , n38468 );
nand ( n38470 , n38466 , n38469 );
not ( n38471 , n38470 );
not ( n38472 , n38471 );
or ( n38473 , n38451 , n38472 );
buf ( n38474 , n38447 );
buf ( n38475 , n38470 );
nand ( n38476 , n38474 , n38475 );
buf ( n38477 , n38476 );
nand ( n38478 , n38473 , n38477 );
buf ( n38479 , n38478 );
buf ( n38480 , n37527 );
not ( n38481 , n38480 );
buf ( n38482 , n38481 );
buf ( n38483 , n38482 );
xor ( n38484 , n38479 , n38483 );
buf ( n38485 , n38484 );
buf ( n38486 , n38485 );
xor ( n38487 , n38433 , n38486 );
buf ( n38488 , n38487 );
xor ( n38489 , n37667 , n37794 );
and ( n38490 , n38489 , n37824 );
and ( n38491 , n37667 , n37794 );
or ( n38492 , n38490 , n38491 );
buf ( n38493 , n38492 );
xor ( n38494 , n38488 , n38493 );
xor ( n38495 , n37689 , n37730 );
and ( n38496 , n38495 , n37792 );
and ( n38497 , n37689 , n37730 );
or ( n38498 , n38496 , n38497 );
buf ( n38499 , n38498 );
not ( n38500 , n37469 );
not ( n38501 , n37481 );
or ( n38502 , n38500 , n38501 );
or ( n38503 , n37481 , n37469 );
nand ( n38504 , n38503 , n37510 );
nand ( n38505 , n38502 , n38504 );
buf ( n38506 , n38505 );
not ( n38507 , n37719 );
not ( n38508 , n957 );
nor ( n38509 , n38508 , n960 );
not ( n38510 , n38509 );
or ( n38511 , n38507 , n38510 );
nand ( n38512 , n38511 , n501 );
buf ( n38513 , n38512 );
buf ( n38514 , n799 );
not ( n38515 , n38514 );
buf ( n38516 , n37467 );
not ( n38517 , n38516 );
or ( n38518 , n38515 , n38517 );
buf ( n38519 , n499 );
not ( n38520 , n38519 );
not ( n38521 , n5562 );
buf ( n38522 , n38521 );
not ( n38523 , n38522 );
or ( n38524 , n38520 , n38523 );
buf ( n38525 , n5562 );
buf ( n38526 , n29901 );
nand ( n38527 , n38525 , n38526 );
buf ( n38528 , n38527 );
buf ( n38529 , n38528 );
nand ( n38530 , n38524 , n38529 );
buf ( n38531 , n38530 );
buf ( n38532 , n38531 );
buf ( n38533 , n29884 );
nand ( n38534 , n38532 , n38533 );
buf ( n38535 , n38534 );
buf ( n38536 , n38535 );
nand ( n38537 , n38518 , n38536 );
buf ( n38538 , n38537 );
buf ( n38539 , n38538 );
xor ( n38540 , n38513 , n38539 );
buf ( n38541 , n3271 );
not ( n38542 , n38541 );
buf ( n38543 , n495 );
not ( n38544 , n38543 );
buf ( n38545 , n32660 );
not ( n38546 , n38545 );
or ( n38547 , n38544 , n38546 );
buf ( n38548 , n32660 );
not ( n38549 , n38548 );
buf ( n38550 , n31784 );
nand ( n38551 , n38549 , n38550 );
buf ( n38552 , n38551 );
buf ( n38553 , n38552 );
nand ( n38554 , n38547 , n38553 );
buf ( n38555 , n38554 );
buf ( n38556 , n38555 );
not ( n38557 , n38556 );
or ( n38558 , n38542 , n38557 );
nand ( n38559 , n37494 , n31812 );
buf ( n38560 , n38559 );
nand ( n38561 , n38558 , n38560 );
buf ( n38562 , n38561 );
buf ( n38563 , n38562 );
xor ( n38564 , n38540 , n38563 );
buf ( n38565 , n38564 );
buf ( n38566 , n38565 );
xor ( n38567 , n38506 , n38566 );
xor ( n38568 , n37748 , n37766 );
and ( n38569 , n38568 , n37791 );
and ( n38570 , n37748 , n37766 );
or ( n38571 , n38569 , n38570 );
buf ( n38572 , n38571 );
xor ( n38573 , n38567 , n38572 );
buf ( n38574 , n38573 );
buf ( n38575 , n38574 );
xor ( n38576 , n38499 , n38575 );
xor ( n38577 , n37516 , n37575 );
and ( n38578 , n38577 , n37598 );
and ( n38579 , n37516 , n37575 );
or ( n38580 , n38578 , n38579 );
buf ( n38581 , n38580 );
buf ( n38582 , n38581 );
xor ( n38583 , n38576 , n38582 );
buf ( n38584 , n38583 );
xor ( n38585 , n38494 , n38584 );
not ( n38586 , n38585 );
xor ( n38587 , n37601 , n37660 );
and ( n38588 , n38587 , n37827 );
and ( n38589 , n37601 , n37660 );
or ( n38590 , n38588 , n38589 );
buf ( n38591 , n38590 );
not ( n38592 , n38591 );
nand ( n38593 , n38586 , n38592 );
nand ( n38594 , n38593 , n37867 , n37846 );
not ( n38595 , n38594 );
not ( n38596 , n38595 );
or ( n38597 , n38369 , n38596 );
nor ( n38598 , n38591 , n38585 );
nor ( n38599 , n38598 , n37847 );
and ( n38600 , n37864 , n38599 );
not ( n38601 , n37849 );
not ( n38602 , n38601 );
not ( n38603 , n38593 );
or ( n38604 , n38602 , n38603 );
nand ( n38605 , n38591 , n38585 );
buf ( n38606 , n38605 );
nand ( n38607 , n38604 , n38606 );
nor ( n38608 , n38600 , n38607 );
nand ( n38609 , n38597 , n38608 );
xor ( n38610 , n38374 , n38432 );
and ( n38611 , n38610 , n38486 );
and ( n38612 , n38374 , n38432 );
or ( n38613 , n38611 , n38612 );
buf ( n38614 , n38613 );
buf ( n38615 , n38614 );
xor ( n38616 , n38499 , n38575 );
and ( n38617 , n38616 , n38582 );
and ( n38618 , n38499 , n38575 );
or ( n38619 , n38617 , n38618 );
buf ( n38620 , n38619 );
buf ( n38621 , n38620 );
xor ( n38622 , n38615 , n38621 );
buf ( n38623 , n799 );
not ( n38624 , n38623 );
buf ( n38625 , n38531 );
not ( n38626 , n38625 );
or ( n38627 , n38624 , n38626 );
buf ( n38628 , n29901 );
not ( n38629 , n38628 );
buf ( n38630 , n29884 );
nand ( n38631 , n38629 , n38630 );
buf ( n38632 , n38631 );
buf ( n38633 , n38632 );
nand ( n38634 , n38627 , n38633 );
buf ( n38635 , n38634 );
buf ( n38636 , n38635 );
not ( n38637 , n38636 );
buf ( n38638 , n38637 );
buf ( n38639 , n38638 );
xor ( n38640 , n38513 , n38539 );
and ( n38641 , n38640 , n38563 );
and ( n38642 , n38513 , n38539 );
or ( n38643 , n38641 , n38642 );
buf ( n38644 , n38643 );
buf ( n38645 , n38644 );
xor ( n38646 , n38639 , n38645 );
xor ( n38647 , n38379 , n38398 );
and ( n38648 , n38647 , n38429 );
and ( n38649 , n38379 , n38398 );
or ( n38650 , n38648 , n38649 );
buf ( n38651 , n38650 );
buf ( n38652 , n38651 );
xor ( n38653 , n38646 , n38652 );
buf ( n38654 , n38653 );
buf ( n38655 , n38654 );
xor ( n38656 , n38506 , n38566 );
and ( n38657 , n38656 , n38572 );
and ( n38658 , n38506 , n38566 );
or ( n38659 , n38657 , n38658 );
buf ( n38660 , n38659 );
buf ( n38661 , n38660 );
xor ( n38662 , n38655 , n38661 );
buf ( n38663 , n38470 );
not ( n38664 , n38663 );
buf ( n38665 , n38450 );
not ( n38666 , n38665 );
or ( n38667 , n38664 , n38666 );
not ( n38668 , n38447 );
not ( n38669 , n38471 );
or ( n38670 , n38668 , n38669 );
nand ( n38671 , n38670 , n38482 );
buf ( n38672 , n38671 );
nand ( n38673 , n38667 , n38672 );
buf ( n38674 , n38673 );
buf ( n38675 , n38674 );
buf ( n38676 , n29983 );
buf ( n38677 , n489 );
and ( n38678 , n38676 , n38677 );
buf ( n38679 , n38678 );
buf ( n38680 , n38679 );
buf ( n38681 , n37542 );
not ( n38682 , n38681 );
buf ( n38683 , n38442 );
not ( n38684 , n38683 );
or ( n38685 , n38682 , n38684 );
buf ( n38686 , n489 );
buf ( n38687 , n933 );
xor ( n38688 , n38686 , n38687 );
buf ( n38689 , n38688 );
buf ( n38690 , n38689 );
buf ( n38691 , n36508 );
nand ( n38692 , n38690 , n38691 );
buf ( n38693 , n38692 );
buf ( n38694 , n38693 );
nand ( n38695 , n38685 , n38694 );
buf ( n38696 , n38695 );
buf ( n38697 , n38696 );
xor ( n38698 , n38680 , n38697 );
buf ( n38699 , n2725 );
not ( n38700 , n38699 );
buf ( n38701 , n495 );
not ( n38702 , n38701 );
buf ( n38703 , n3211 );
not ( n38704 , n38703 );
or ( n38705 , n38702 , n38704 );
buf ( n38706 , n3220 );
buf ( n38707 , n31784 );
nand ( n38708 , n38706 , n38707 );
buf ( n38709 , n38708 );
buf ( n38710 , n38709 );
nand ( n38711 , n38705 , n38710 );
buf ( n38712 , n38711 );
buf ( n38713 , n38712 );
not ( n38714 , n38713 );
or ( n38715 , n38700 , n38714 );
buf ( n38716 , n38555 );
buf ( n38717 , n31812 );
nand ( n38718 , n38716 , n38717 );
buf ( n38719 , n38718 );
buf ( n38720 , n38719 );
nand ( n38721 , n38715 , n38720 );
buf ( n38722 , n38721 );
buf ( n38723 , n38722 );
xor ( n38724 , n38698 , n38723 );
buf ( n38725 , n38724 );
buf ( n38726 , n38725 );
xor ( n38727 , n38675 , n38726 );
buf ( n38728 , n30585 );
not ( n38729 , n38728 );
buf ( n38730 , n38421 );
not ( n38731 , n38730 );
or ( n38732 , n38729 , n38731 );
not ( n38733 , n497 );
not ( n38734 , n3848 );
or ( n38735 , n38733 , n38734 );
buf ( n38736 , n37462 );
buf ( n38737 , n30599 );
nand ( n38738 , n38736 , n38737 );
buf ( n38739 , n38738 );
nand ( n38740 , n38735 , n38739 );
buf ( n38741 , n38740 );
buf ( n38742 , n910 );
nand ( n38743 , n38741 , n38742 );
buf ( n38744 , n38743 );
buf ( n38745 , n38744 );
nand ( n38746 , n38732 , n38745 );
buf ( n38747 , n38746 );
buf ( n38748 , n3045 );
not ( n38749 , n38748 );
buf ( n38750 , n491 );
not ( n38751 , n38750 );
buf ( n38752 , n1883 );
not ( n38753 , n38752 );
or ( n38754 , n38751 , n38753 );
buf ( n38755 , n29501 );
buf ( n38756 , n3524 );
nand ( n38757 , n38755 , n38756 );
buf ( n38758 , n38757 );
buf ( n38759 , n38758 );
nand ( n38760 , n38754 , n38759 );
buf ( n38761 , n38760 );
buf ( n38762 , n38761 );
not ( n38763 , n38762 );
or ( n38764 , n38749 , n38763 );
buf ( n38765 , n38464 );
buf ( n38766 , n3948 );
nand ( n38767 , n38765 , n38766 );
buf ( n38768 , n38767 );
buf ( n38769 , n38768 );
nand ( n38770 , n38764 , n38769 );
buf ( n38771 , n38770 );
xor ( n38772 , n38747 , n38771 );
not ( n38773 , n3113 );
buf ( n38774 , n493 );
not ( n38775 , n38774 );
buf ( n38776 , n32975 );
not ( n38777 , n38776 );
or ( n38778 , n38775 , n38777 );
buf ( n38779 , n2803 );
buf ( n38780 , n2704 );
nand ( n38781 , n38779 , n38780 );
buf ( n38782 , n38781 );
buf ( n38783 , n38782 );
nand ( n38784 , n38778 , n38783 );
buf ( n38785 , n38784 );
not ( n38786 , n38785 );
or ( n38787 , n38773 , n38786 );
nand ( n38788 , n38395 , n3146 );
nand ( n38789 , n38787 , n38788 );
xor ( n38790 , n38772 , n38789 );
buf ( n38791 , n38790 );
xor ( n38792 , n38727 , n38791 );
buf ( n38793 , n38792 );
buf ( n38794 , n38793 );
xor ( n38795 , n38662 , n38794 );
buf ( n38796 , n38795 );
buf ( n38797 , n38796 );
xor ( n38798 , n38622 , n38797 );
buf ( n38799 , n38798 );
not ( n38800 , n38799 );
xor ( n38801 , n38488 , n38493 );
and ( n38802 , n38801 , n38584 );
and ( n38803 , n38488 , n38493 );
or ( n38804 , n38802 , n38803 );
not ( n38805 , n38804 );
nand ( n38806 , n38800 , n38805 );
not ( n38807 , n38799 );
not ( n38808 , n38807 );
nand ( n38809 , n38808 , n38804 );
nand ( n38810 , n38806 , n38809 );
not ( n38811 , n38810 );
and ( n38812 , n38609 , n38811 );
not ( n38813 , n38609 );
and ( n38814 , n38813 , n38810 );
nor ( n38815 , n38812 , n38814 );
nand ( n38816 , n38815 , n455 );
nand ( n38817 , n38364 , n38816 );
not ( n38818 , n38817 );
not ( n38819 , n37849 );
not ( n38820 , n37869 );
not ( n38821 , n37865 );
or ( n38822 , n38820 , n38821 );
buf ( n38823 , n37846 );
nand ( n38824 , n38822 , n38823 );
not ( n38825 , n38824 );
or ( n38826 , n38819 , n38825 );
buf ( n38827 , n38593 );
and ( n38828 , n38827 , n38606 );
nor ( n38829 , n38828 , n29519 );
nand ( n38830 , n38826 , n38829 );
not ( n38831 , n37418 );
nand ( n38832 , n37440 , n37417 );
not ( n38833 , n38832 );
or ( n38834 , n38831 , n38833 );
and ( n38835 , n38172 , n38185 );
nor ( n38836 , n38835 , n455 );
nand ( n38837 , n38834 , n38836 );
not ( n38838 , n455 );
not ( n38839 , n37844 );
not ( n38840 , n37829 );
or ( n38841 , n38839 , n38840 );
nand ( n38842 , n38841 , n38605 );
nor ( n38843 , n38838 , n38842 );
and ( n38844 , n38827 , n38843 );
nand ( n38845 , n38824 , n38844 );
and ( n38846 , n38185 , n37418 );
not ( n38847 , n38846 );
nor ( n38848 , n38847 , n38178 , n455 );
nand ( n38849 , n38832 , n38848 );
nand ( n38850 , n38830 , n38837 , n38845 , n38849 );
nor ( n38851 , n38818 , n38850 );
buf ( n38852 , n38851 );
nand ( n38853 , n38830 , n38837 , n38845 , n38849 );
not ( n38854 , n38853 );
buf ( n38855 , n37877 );
buf ( n38856 , n537 );
or ( n38857 , n38855 , n38856 );
buf ( n38858 , n38857 );
nor ( n38859 , n38854 , n38858 );
buf ( n38860 , n38859 );
nor ( n38861 , n38852 , n38860 );
buf ( n38862 , n38861 );
buf ( n38863 , n38862 );
buf ( n38864 , n38863 );
buf ( n38865 , n38864 );
not ( n38866 , n38359 );
not ( n38867 , n38188 );
or ( n38868 , n38866 , n38867 );
nand ( n38869 , n38868 , n38360 );
xor ( n38870 , n38311 , n38328 );
and ( n38871 , n38870 , n38346 );
and ( n38872 , n38311 , n38328 );
or ( n38873 , n38871 , n38872 );
buf ( n38874 , n38873 );
buf ( n38875 , n38874 );
not ( n38876 , n29534 );
not ( n38877 , n29542 );
not ( n38878 , n38877 );
or ( n38879 , n38876 , n38878 );
nand ( n38880 , n38879 , n499 );
buf ( n38881 , n38880 );
buf ( n38882 , n38279 );
not ( n38883 , n38882 );
buf ( n38884 , n30769 );
not ( n38885 , n38884 );
or ( n38886 , n38883 , n38885 );
buf ( n38887 , n1786 );
buf ( n38888 , n505 );
buf ( n38889 , n497 );
xor ( n38890 , n38888 , n38889 );
buf ( n38891 , n38890 );
buf ( n38892 , n38891 );
nand ( n38893 , n38887 , n38892 );
buf ( n38894 , n38893 );
buf ( n38895 , n38894 );
nand ( n38896 , n38886 , n38895 );
buf ( n38897 , n38896 );
buf ( n38898 , n38897 );
xor ( n38899 , n38881 , n38898 );
buf ( n38900 , n38297 );
not ( n38901 , n38900 );
buf ( n38902 , n4241 );
not ( n38903 , n38902 );
or ( n38904 , n38901 , n38903 );
buf ( n38905 , n4218 );
buf ( n38906 , n509 );
buf ( n38907 , n493 );
xor ( n38908 , n38906 , n38907 );
buf ( n38909 , n38908 );
buf ( n38910 , n38909 );
nand ( n38911 , n38905 , n38910 );
buf ( n38912 , n38911 );
buf ( n38913 , n38912 );
nand ( n38914 , n38904 , n38913 );
buf ( n38915 , n38914 );
buf ( n38916 , n38915 );
xor ( n38917 , n38899 , n38916 );
buf ( n38918 , n38917 );
buf ( n38919 , n38918 );
xor ( n38920 , n38875 , n38919 );
buf ( n38921 , n38321 );
not ( n38922 , n38921 );
buf ( n38923 , n36290 );
not ( n38924 , n38923 );
or ( n38925 , n38922 , n38924 );
buf ( n38926 , n37254 );
buf ( n38927 , n489 );
buf ( n38928 , n513 );
xor ( n38929 , n38927 , n38928 );
buf ( n38930 , n38929 );
buf ( n38931 , n38930 );
nand ( n38932 , n38926 , n38931 );
buf ( n38933 , n38932 );
buf ( n38934 , n38933 );
nand ( n38935 , n38925 , n38934 );
buf ( n38936 , n38935 );
buf ( n38937 , n38936 );
buf ( n38938 , n38266 );
not ( n38939 , n38938 );
buf ( n38940 , n33967 );
not ( n38941 , n38940 );
or ( n38942 , n38939 , n38941 );
buf ( n38943 , n33973 );
buf ( n38944 , n511 );
buf ( n38945 , n491 );
xor ( n38946 , n38944 , n38945 );
buf ( n38947 , n38946 );
buf ( n38948 , n38947 );
nand ( n38949 , n38943 , n38948 );
buf ( n38950 , n38949 );
buf ( n38951 , n38950 );
nand ( n38952 , n38942 , n38951 );
buf ( n38953 , n38952 );
buf ( n38954 , n38953 );
xor ( n38955 , n38937 , n38954 );
buf ( n38956 , n38339 );
not ( n38957 , n38956 );
buf ( n38958 , n33754 );
not ( n38959 , n38958 );
or ( n38960 , n38957 , n38959 );
buf ( n38961 , n507 );
buf ( n38962 , n495 );
xor ( n38963 , n38961 , n38962 );
buf ( n38964 , n38963 );
buf ( n38965 , n38964 );
buf ( n38966 , n33167 );
nand ( n38967 , n38965 , n38966 );
buf ( n38968 , n38967 );
buf ( n38969 , n38968 );
nand ( n38970 , n38960 , n38969 );
buf ( n38971 , n38970 );
buf ( n38972 , n38971 );
xor ( n38973 , n38955 , n38972 );
buf ( n38974 , n38973 );
buf ( n38975 , n38974 );
xor ( n38976 , n38920 , n38975 );
buf ( n38977 , n38976 );
and ( n38978 , n38026 , n38027 );
buf ( n38979 , n38978 );
xor ( n38980 , n38979 , n38219 );
xor ( n38981 , n38269 , n38286 );
and ( n38982 , n38981 , n38304 );
and ( n38983 , n38269 , n38286 );
or ( n38984 , n38982 , n38983 );
buf ( n38985 , n38984 );
xor ( n38986 , n38980 , n38985 );
buf ( n38987 , n38986 );
xor ( n38988 , n38221 , n38227 );
and ( n38989 , n38988 , n38234 );
and ( n38990 , n38221 , n38227 );
or ( n38991 , n38989 , n38990 );
buf ( n38992 , n38991 );
buf ( n38993 , n38992 );
xor ( n38994 , n38987 , n38993 );
xor ( n38995 , n38259 , n38307 );
and ( n38996 , n38995 , n38349 );
and ( n38997 , n38259 , n38307 );
or ( n38998 , n38996 , n38997 );
buf ( n38999 , n38998 );
buf ( n39000 , n38999 );
xor ( n39001 , n38994 , n39000 );
buf ( n39002 , n39001 );
xor ( n39003 , n38977 , n39002 );
xor ( n39004 , n38237 , n38243 );
and ( n39005 , n39004 , n38352 );
and ( n39006 , n38237 , n38243 );
or ( n39007 , n39005 , n39006 );
buf ( n39008 , n39007 );
xor ( n39009 , n39003 , n39008 );
not ( n39010 , n39009 );
xor ( n39011 , n38200 , n38206 );
and ( n39012 , n39011 , n38355 );
and ( n39013 , n38200 , n38206 );
or ( n39014 , n39012 , n39013 );
buf ( n39015 , n39014 );
not ( n39016 , n39015 );
nand ( n39017 , n39010 , n39016 );
nand ( n39018 , n39009 , n39015 );
nand ( n39019 , n39017 , n39018 );
xnor ( n39020 , n38869 , n39019 );
nand ( n39021 , n39020 , n29519 );
not ( n39022 , n39021 );
not ( n39023 , n38806 );
not ( n39024 , n38609 );
or ( n39025 , n39023 , n39024 );
buf ( n39026 , n38809 );
nand ( n39027 , n39025 , n39026 );
xor ( n39028 , n38680 , n38697 );
and ( n39029 , n39028 , n38723 );
and ( n39030 , n38680 , n38697 );
or ( n39031 , n39029 , n39030 );
buf ( n39032 , n39031 );
buf ( n39033 , n39032 );
not ( n39034 , n29884 );
buf ( n39035 , n39034 );
not ( n39036 , n39035 );
buf ( n39037 , n798 );
not ( n39038 , n39037 );
or ( n39039 , n39036 , n39038 );
buf ( n39040 , n499 );
nand ( n39041 , n39039 , n39040 );
buf ( n39042 , n39041 );
buf ( n39043 , n39042 );
buf ( n39044 , n909 );
not ( n39045 , n39044 );
buf ( n39046 , n497 );
not ( n39047 , n39046 );
buf ( n39048 , n38521 );
not ( n39049 , n39048 );
or ( n39050 , n39047 , n39049 );
buf ( n39051 , n5562 );
buf ( n39052 , n30599 );
nand ( n39053 , n39051 , n39052 );
buf ( n39054 , n39053 );
buf ( n39055 , n39054 );
nand ( n39056 , n39050 , n39055 );
buf ( n39057 , n39056 );
buf ( n39058 , n39057 );
not ( n39059 , n39058 );
or ( n39060 , n39045 , n39059 );
buf ( n39061 , n38740 );
buf ( n39062 , n30585 );
nand ( n39063 , n39061 , n39062 );
buf ( n39064 , n39063 );
buf ( n39065 , n39064 );
nand ( n39066 , n39060 , n39065 );
buf ( n39067 , n39066 );
buf ( n39068 , n39067 );
xor ( n39069 , n39043 , n39068 );
buf ( n39070 , n3113 );
not ( n39071 , n39070 );
buf ( n39072 , n493 );
not ( n39073 , n39072 );
buf ( n39074 , n31829 );
not ( n39075 , n39074 );
or ( n39076 , n39073 , n39075 );
buf ( n39077 , n31826 );
buf ( n39078 , n2704 );
nand ( n39079 , n39077 , n39078 );
buf ( n39080 , n39079 );
buf ( n39081 , n39080 );
nand ( n39082 , n39076 , n39081 );
buf ( n39083 , n39082 );
buf ( n39084 , n39083 );
not ( n39085 , n39084 );
or ( n39086 , n39071 , n39085 );
buf ( n39087 , n38785 );
buf ( n39088 , n3146 );
nand ( n39089 , n39087 , n39088 );
buf ( n39090 , n39089 );
buf ( n39091 , n39090 );
nand ( n39092 , n39086 , n39091 );
buf ( n39093 , n39092 );
buf ( n39094 , n39093 );
xor ( n39095 , n39069 , n39094 );
buf ( n39096 , n39095 );
buf ( n39097 , n39096 );
xor ( n39098 , n39033 , n39097 );
buf ( n39099 , n31812 );
not ( n39100 , n39099 );
buf ( n39101 , n38712 );
not ( n39102 , n39101 );
or ( n39103 , n39100 , n39102 );
buf ( n39104 , n495 );
not ( n39105 , n39104 );
buf ( n39106 , n38410 );
not ( n39107 , n39106 );
or ( n39108 , n39105 , n39107 );
buf ( n39109 , n38414 );
buf ( n39110 , n31784 );
nand ( n39111 , n39109 , n39110 );
buf ( n39112 , n39111 );
buf ( n39113 , n39112 );
nand ( n39114 , n39108 , n39113 );
buf ( n39115 , n39114 );
buf ( n39116 , n39115 );
buf ( n39117 , n3271 );
nand ( n39118 , n39116 , n39117 );
buf ( n39119 , n39118 );
buf ( n39120 , n39119 );
nand ( n39121 , n39103 , n39120 );
buf ( n39122 , n39121 );
buf ( n39123 , n39122 );
buf ( n39124 , n3045 );
not ( n39125 , n39124 );
buf ( n39126 , n491 );
not ( n39127 , n39126 );
buf ( n39128 , n2671 );
not ( n39129 , n39128 );
or ( n39130 , n39127 , n39129 );
nand ( n39131 , n38391 , n3524 );
buf ( n39132 , n39131 );
nand ( n39133 , n39130 , n39132 );
buf ( n39134 , n39133 );
buf ( n39135 , n39134 );
not ( n39136 , n39135 );
or ( n39137 , n39125 , n39136 );
buf ( n39138 , n38761 );
buf ( n39139 , n3948 );
nand ( n39140 , n39138 , n39139 );
buf ( n39141 , n39140 );
buf ( n39142 , n39141 );
nand ( n39143 , n39137 , n39142 );
buf ( n39144 , n39143 );
buf ( n39145 , n39144 );
xor ( n39146 , n39123 , n39145 );
buf ( n39147 , n37542 );
buf ( n39148 , n39147 );
buf ( n39149 , n39148 );
buf ( n39150 , n39149 );
not ( n39151 , n39150 );
buf ( n39152 , n38689 );
not ( n39153 , n39152 );
or ( n39154 , n39151 , n39153 );
buf ( n39155 , n489 );
buf ( n39156 , n2633 );
xor ( n39157 , n39155 , n39156 );
buf ( n39158 , n39157 );
buf ( n39159 , n39158 );
buf ( n39160 , n36508 );
nand ( n39161 , n39159 , n39160 );
buf ( n39162 , n39161 );
buf ( n39163 , n39162 );
nand ( n39164 , n39154 , n39163 );
buf ( n39165 , n39164 );
buf ( n39166 , n39165 );
xor ( n39167 , n39146 , n39166 );
buf ( n39168 , n39167 );
buf ( n39169 , n39168 );
xor ( n39170 , n39098 , n39169 );
buf ( n39171 , n39170 );
and ( n39172 , n489 , n2831 );
buf ( n39173 , n39172 );
buf ( n39174 , n38635 );
xor ( n39175 , n39173 , n39174 );
buf ( n39176 , n38789 );
not ( n39177 , n39176 );
buf ( n39178 , n38771 );
not ( n39179 , n39178 );
or ( n39180 , n39177 , n39179 );
buf ( n39181 , n38771 );
buf ( n39182 , n38789 );
or ( n39183 , n39181 , n39182 );
buf ( n39184 , n38747 );
nand ( n39185 , n39183 , n39184 );
buf ( n39186 , n39185 );
buf ( n39187 , n39186 );
nand ( n39188 , n39180 , n39187 );
buf ( n39189 , n39188 );
buf ( n39190 , n39189 );
xor ( n39191 , n39175 , n39190 );
buf ( n39192 , n39191 );
buf ( n39193 , n39192 );
xor ( n39194 , n38639 , n38645 );
and ( n39195 , n39194 , n38652 );
and ( n39196 , n38639 , n38645 );
or ( n39197 , n39195 , n39196 );
buf ( n39198 , n39197 );
buf ( n39199 , n39198 );
xor ( n39200 , n39193 , n39199 );
xor ( n39201 , n38675 , n38726 );
and ( n39202 , n39201 , n38791 );
and ( n39203 , n38675 , n38726 );
or ( n39204 , n39202 , n39203 );
buf ( n39205 , n39204 );
buf ( n39206 , n39205 );
xor ( n39207 , n39200 , n39206 );
buf ( n39208 , n39207 );
xor ( n39209 , n39171 , n39208 );
xor ( n39210 , n38655 , n38661 );
and ( n39211 , n39210 , n38794 );
and ( n39212 , n38655 , n38661 );
or ( n39213 , n39211 , n39212 );
buf ( n39214 , n39213 );
xor ( n39215 , n39209 , n39214 );
not ( n39216 , n39215 );
xor ( n39217 , n38615 , n38621 );
and ( n39218 , n39217 , n38797 );
and ( n39219 , n38615 , n38621 );
or ( n39220 , n39218 , n39219 );
buf ( n39221 , n39220 );
not ( n39222 , n39221 );
nand ( n39223 , n39216 , n39222 );
nand ( n39224 , n39221 , n39215 );
nand ( n39225 , n39223 , n39224 );
not ( n39226 , n39225 );
and ( n39227 , n39027 , n39226 );
not ( n39228 , n39027 );
and ( n39229 , n39228 , n39225 );
nor ( n39230 , n39227 , n39229 );
nand ( n39231 , n39230 , n455 );
not ( n39232 , n39231 );
or ( n39233 , n39022 , n39232 );
nand ( n39234 , n39233 , n38818 );
buf ( n39235 , n39234 );
buf ( n39236 , n39235 );
buf ( n39237 , n39236 );
and ( n39238 , n38865 , n39237 );
buf ( n39239 , n39238 );
not ( n39240 , n39239 );
or ( n39241 , n37968 , n39240 );
buf ( n39242 , n38858 );
not ( n39243 , n39242 );
buf ( n39244 , n39243 );
not ( n39245 , n39244 );
nor ( n39246 , n38817 , n38853 );
nand ( n39247 , n39245 , n39246 );
buf ( n39248 , n38818 );
nand ( n39249 , n39248 , n38853 );
nand ( n39250 , n39247 , n39249 );
buf ( n39251 , n39250 );
buf ( n39252 , n39237 );
and ( n39253 , n39251 , n39252 );
not ( n39254 , n29519 );
not ( n39255 , n39020 );
or ( n39256 , n39254 , n39255 );
nand ( n39257 , n39256 , n39231 );
not ( n39258 , n39257 );
not ( n39259 , n39258 );
nor ( n39260 , n39259 , n39248 );
buf ( n39261 , n39260 );
nor ( n39262 , n39253 , n39261 );
buf ( n39263 , n39262 );
buf ( n39264 , n39263 );
nand ( n39265 , n39241 , n39264 );
buf ( n39266 , n39265 );
not ( n39267 , n39259 );
xor ( n39268 , n39123 , n39145 );
and ( n39269 , n39268 , n39166 );
and ( n39270 , n39123 , n39145 );
or ( n39271 , n39269 , n39270 );
buf ( n39272 , n39271 );
buf ( n39273 , n39272 );
xor ( n39274 , n39043 , n39068 );
and ( n39275 , n39274 , n39094 );
and ( n39276 , n39043 , n39068 );
or ( n39277 , n39275 , n39276 );
buf ( n39278 , n39277 );
buf ( n39279 , n39278 );
xor ( n39280 , n39273 , n39279 );
not ( n39281 , n3948 );
not ( n39282 , n39134 );
or ( n39283 , n39281 , n39282 );
buf ( n39284 , n491 );
not ( n39285 , n39284 );
buf ( n39286 , n32126 );
not ( n39287 , n39286 );
or ( n39288 , n39285 , n39287 );
buf ( n39289 , n2803 );
buf ( n39290 , n3524 );
nand ( n39291 , n39289 , n39290 );
buf ( n39292 , n39291 );
buf ( n39293 , n39292 );
nand ( n39294 , n39288 , n39293 );
buf ( n39295 , n39294 );
buf ( n39296 , n39295 );
buf ( n39297 , n3045 );
nand ( n39298 , n39296 , n39297 );
buf ( n39299 , n39298 );
nand ( n39300 , n39283 , n39299 );
buf ( n39301 , n30585 );
not ( n39302 , n39301 );
buf ( n39303 , n39057 );
not ( n39304 , n39303 );
or ( n39305 , n39302 , n39304 );
buf ( n39306 , n30599 );
not ( n39307 , n39306 );
buf ( n39308 , n910 );
nand ( n39309 , n39307 , n39308 );
buf ( n39310 , n39309 );
buf ( n39311 , n39310 );
nand ( n39312 , n39305 , n39311 );
buf ( n39313 , n39312 );
xor ( n39314 , n39300 , n39313 );
buf ( n39315 , n39149 );
not ( n39316 , n39315 );
buf ( n39317 , n39158 );
not ( n39318 , n39317 );
or ( n39319 , n39316 , n39318 );
buf ( n39320 , n489 );
buf ( n39321 , n31693 );
not ( n39322 , n39321 );
buf ( n39323 , n39322 );
buf ( n39324 , n39323 );
xor ( n39325 , n39320 , n39324 );
buf ( n39326 , n39325 );
buf ( n39327 , n39326 );
buf ( n39328 , n36508 );
nand ( n39329 , n39327 , n39328 );
buf ( n39330 , n39329 );
buf ( n39331 , n39330 );
nand ( n39332 , n39319 , n39331 );
buf ( n39333 , n39332 );
xor ( n39334 , n39314 , n39333 );
buf ( n39335 , n39334 );
xor ( n39336 , n39280 , n39335 );
buf ( n39337 , n39336 );
buf ( n39338 , n39337 );
xor ( n39339 , n39193 , n39199 );
and ( n39340 , n39339 , n39206 );
and ( n39341 , n39193 , n39199 );
or ( n39342 , n39340 , n39341 );
buf ( n39343 , n39342 );
buf ( n39344 , n39343 );
xor ( n39345 , n39338 , n39344 );
and ( n39346 , n38686 , n38687 );
buf ( n39347 , n39346 );
buf ( n39348 , n39347 );
buf ( n39349 , n31812 );
not ( n39350 , n39349 );
buf ( n39351 , n39115 );
not ( n39352 , n39351 );
or ( n39353 , n39350 , n39352 );
not ( n39354 , n37462 );
not ( n39355 , n31784 );
or ( n39356 , n39354 , n39355 );
nand ( n39357 , n3854 , n495 );
nand ( n39358 , n39356 , n39357 );
buf ( n39359 , n39358 );
buf ( n39360 , n2725 );
nand ( n39361 , n39359 , n39360 );
buf ( n39362 , n39361 );
buf ( n39363 , n39362 );
nand ( n39364 , n39353 , n39363 );
buf ( n39365 , n39364 );
buf ( n39366 , n39365 );
not ( n39367 , n39366 );
buf ( n39368 , n39367 );
buf ( n39369 , n39368 );
xor ( n39370 , n39348 , n39369 );
buf ( n39371 , n3146 );
not ( n39372 , n39371 );
buf ( n39373 , n39083 );
not ( n39374 , n39373 );
or ( n39375 , n39372 , n39374 );
buf ( n39376 , n2704 );
not ( n39377 , n39376 );
buf ( n39378 , n3220 );
not ( n39379 , n39378 );
or ( n39380 , n39377 , n39379 );
buf ( n39381 , n3211 );
not ( n39382 , n39381 );
buf ( n39383 , n39382 );
buf ( n39384 , n39383 );
buf ( n39385 , n2704 );
or ( n39386 , n39384 , n39385 );
nand ( n39387 , n39380 , n39386 );
buf ( n39388 , n39387 );
buf ( n39389 , n39388 );
buf ( n39390 , n3113 );
nand ( n39391 , n39389 , n39390 );
buf ( n39392 , n39391 );
buf ( n39393 , n39392 );
nand ( n39394 , n39375 , n39393 );
buf ( n39395 , n39394 );
buf ( n39396 , n39395 );
xor ( n39397 , n39370 , n39396 );
buf ( n39398 , n39397 );
buf ( n39399 , n39398 );
xor ( n39400 , n39173 , n39174 );
and ( n39401 , n39400 , n39190 );
and ( n39402 , n39173 , n39174 );
or ( n39403 , n39401 , n39402 );
buf ( n39404 , n39403 );
buf ( n39405 , n39404 );
xor ( n39406 , n39399 , n39405 );
xor ( n39407 , n39033 , n39097 );
and ( n39408 , n39407 , n39169 );
and ( n39409 , n39033 , n39097 );
or ( n39410 , n39408 , n39409 );
buf ( n39411 , n39410 );
buf ( n39412 , n39411 );
xor ( n39413 , n39406 , n39412 );
buf ( n39414 , n39413 );
buf ( n39415 , n39414 );
xor ( n39416 , n39345 , n39415 );
buf ( n39417 , n39416 );
not ( n39418 , n39417 );
xor ( n39419 , n39171 , n39208 );
and ( n39420 , n39419 , n39214 );
and ( n39421 , n39171 , n39208 );
or ( n39422 , n39420 , n39421 );
not ( n39423 , n39422 );
nand ( n39424 , n39418 , n39423 );
not ( n39425 , n39424 );
not ( n39426 , n39425 );
nand ( n39427 , n39417 , n39422 );
buf ( n39428 , n39427 );
and ( n39429 , n39426 , n39428 );
nand ( n39430 , n39216 , n39222 );
not ( n39431 , n39430 );
not ( n39432 , n38806 );
nor ( n39433 , n39431 , n39432 );
not ( n39434 , n39433 );
not ( n39435 , n38609 );
or ( n39436 , n39434 , n39435 );
nor ( n39437 , n38807 , n38805 );
nand ( n39438 , n39223 , n39437 );
nand ( n39439 , n39221 , n39215 );
nand ( n39440 , n39438 , n39439 );
not ( n39441 , n39440 );
nand ( n39442 , n39436 , n39441 );
xor ( n39443 , n39429 , n39442 );
nand ( n39444 , n39443 , n455 );
and ( n39445 , n38359 , n39017 );
not ( n39446 , n39445 );
not ( n39447 , n38188 );
or ( n39448 , n39446 , n39447 );
not ( n39449 , n38360 );
nand ( n39450 , n39449 , n39017 );
nand ( n39451 , n39450 , n39018 );
not ( n39452 , n39451 );
nand ( n39453 , n39448 , n39452 );
buf ( n39454 , n38947 );
not ( n39455 , n39454 );
buf ( n39456 , n4370 );
not ( n39457 , n39456 );
or ( n39458 , n39455 , n39457 );
buf ( n39459 , n33102 );
buf ( n39460 , n510 );
buf ( n39461 , n491 );
xor ( n39462 , n39460 , n39461 );
buf ( n39463 , n39462 );
buf ( n39464 , n39463 );
nand ( n39465 , n39459 , n39464 );
buf ( n39466 , n39465 );
buf ( n39467 , n39466 );
nand ( n39468 , n39458 , n39467 );
buf ( n39469 , n39468 );
buf ( n39470 , n38891 );
not ( n39471 , n39470 );
buf ( n39472 , n1691 );
not ( n39473 , n39472 );
or ( n39474 , n39471 , n39473 );
buf ( n39475 , n29604 );
buf ( n39476 , n497 );
nand ( n39477 , n39475 , n39476 );
buf ( n39478 , n39477 );
buf ( n39479 , n39478 );
nand ( n39480 , n39474 , n39479 );
buf ( n39481 , n39480 );
xor ( n39482 , n39469 , n39481 );
buf ( n39483 , n38930 );
not ( n39484 , n39483 );
buf ( n39485 , n5172 );
not ( n39486 , n39485 );
or ( n39487 , n39484 , n39486 );
buf ( n39488 , n37254 );
buf ( n39489 , n489 );
buf ( n39490 , n512 );
xor ( n39491 , n39489 , n39490 );
buf ( n39492 , n39491 );
buf ( n39493 , n39492 );
nand ( n39494 , n39488 , n39493 );
buf ( n39495 , n39494 );
buf ( n39496 , n39495 );
nand ( n39497 , n39487 , n39496 );
buf ( n39498 , n39497 );
xor ( n39499 , n39482 , n39498 );
buf ( n39500 , n39499 );
xor ( n39501 , n38881 , n38898 );
and ( n39502 , n39501 , n38916 );
and ( n39503 , n38881 , n38898 );
or ( n39504 , n39502 , n39503 );
buf ( n39505 , n39504 );
buf ( n39506 , n39505 );
xor ( n39507 , n39500 , n39506 );
xor ( n39508 , n38937 , n38954 );
and ( n39509 , n39508 , n38972 );
and ( n39510 , n38937 , n38954 );
or ( n39511 , n39509 , n39510 );
buf ( n39512 , n39511 );
buf ( n39513 , n39512 );
xor ( n39514 , n39507 , n39513 );
buf ( n39515 , n39514 );
xor ( n39516 , n38987 , n38993 );
and ( n39517 , n39516 , n39000 );
and ( n39518 , n38987 , n38993 );
or ( n39519 , n39517 , n39518 );
buf ( n39520 , n39519 );
xor ( n39521 , n39515 , n39520 );
and ( n39522 , n38318 , n38319 );
buf ( n39523 , n39522 );
buf ( n39524 , n39523 );
buf ( n39525 , n38909 );
not ( n39526 , n39525 );
buf ( n39527 , n4241 );
not ( n39528 , n39527 );
or ( n39529 , n39526 , n39528 );
buf ( n39530 , n508 );
buf ( n39531 , n493 );
xor ( n39532 , n39530 , n39531 );
buf ( n39533 , n39532 );
buf ( n39534 , n39533 );
buf ( n39535 , n4218 );
nand ( n39536 , n39534 , n39535 );
buf ( n39537 , n39536 );
buf ( n39538 , n39537 );
nand ( n39539 , n39529 , n39538 );
buf ( n39540 , n39539 );
buf ( n39541 , n39540 );
xor ( n39542 , n39524 , n39541 );
buf ( n39543 , n38964 );
not ( n39544 , n39543 );
buf ( n39545 , n33754 );
not ( n39546 , n39545 );
or ( n39547 , n39544 , n39546 );
buf ( n39548 , n33167 );
buf ( n39549 , n495 );
buf ( n39550 , n506 );
xor ( n39551 , n39549 , n39550 );
buf ( n39552 , n39551 );
buf ( n39553 , n39552 );
nand ( n39554 , n39548 , n39553 );
buf ( n39555 , n39554 );
buf ( n39556 , n39555 );
nand ( n39557 , n39547 , n39556 );
buf ( n39558 , n39557 );
buf ( n39559 , n39558 );
not ( n39560 , n39559 );
buf ( n39561 , n39560 );
buf ( n39562 , n39561 );
xor ( n39563 , n39542 , n39562 );
buf ( n39564 , n39563 );
buf ( n39565 , n39564 );
nand ( n39566 , n38979 , n38219 );
nand ( n39567 , n38979 , n38985 );
nand ( n39568 , n38219 , n38985 );
nand ( n39569 , n39566 , n39567 , n39568 );
buf ( n39570 , n39569 );
xor ( n39571 , n39565 , n39570 );
xor ( n39572 , n38875 , n38919 );
and ( n39573 , n39572 , n38975 );
and ( n39574 , n38875 , n38919 );
or ( n39575 , n39573 , n39574 );
buf ( n39576 , n39575 );
buf ( n39577 , n39576 );
xor ( n39578 , n39571 , n39577 );
buf ( n39579 , n39578 );
xor ( n39580 , n39521 , n39579 );
not ( n39581 , n39580 );
xor ( n39582 , n38977 , n39002 );
and ( n39583 , n39582 , n39008 );
and ( n39584 , n38977 , n39002 );
or ( n39585 , n39583 , n39584 );
not ( n39586 , n39585 );
nand ( n39587 , n39581 , n39586 );
nand ( n39588 , n39580 , n39585 );
nand ( n39589 , n39587 , n39588 );
not ( n39590 , n39589 );
and ( n39591 , n39453 , n39590 );
not ( n39592 , n39453 );
and ( n39593 , n39592 , n39589 );
nor ( n39594 , n39591 , n39593 );
nand ( n39595 , n39594 , n29519 );
nand ( n39596 , n39444 , n39595 );
not ( n39597 , n39596 );
buf ( n39598 , n39597 );
not ( n39599 , n39598 );
or ( n39600 , n39267 , n39599 );
not ( n39601 , n39257 );
not ( n39602 , n455 );
not ( n39603 , n39443 );
or ( n39604 , n39602 , n39603 );
nand ( n39605 , n39604 , n39595 );
nand ( n39606 , n39601 , n39605 );
buf ( n39607 , n39606 );
nand ( n39608 , n39600 , n39607 );
and ( n39609 , n39608 , n454 );
and ( n39610 , n39266 , n39609 );
not ( n39611 , n39266 );
not ( n39612 , n454 );
nor ( n39613 , n39612 , n39608 );
and ( n39614 , n39611 , n39613 );
nor ( n39615 , n39610 , n39614 );
buf ( n39616 , n526 );
buf ( n39617 , n546 );
and ( n39618 , n39616 , n39617 );
buf ( n39619 , n39618 );
buf ( n39620 , n39619 );
buf ( n39621 , n532 );
buf ( n39622 , n540 );
and ( n39623 , n39621 , n39622 );
buf ( n39624 , n39623 );
buf ( n39625 , n39624 );
xor ( n39626 , n39620 , n39625 );
buf ( n39627 , n533 );
buf ( n39628 , n539 );
and ( n39629 , n39627 , n39628 );
buf ( n39630 , n39629 );
buf ( n39631 , n39630 );
xor ( n39632 , n39626 , n39631 );
buf ( n39633 , n39632 );
buf ( n39634 , n39633 );
buf ( n39635 , n530 );
buf ( n39636 , n542 );
and ( n39637 , n39635 , n39636 );
buf ( n39638 , n39637 );
buf ( n39639 , n39638 );
buf ( n39640 , n531 );
buf ( n39641 , n541 );
and ( n39642 , n39640 , n39641 );
buf ( n39643 , n39642 );
buf ( n39644 , n39643 );
xor ( n39645 , n39639 , n39644 );
buf ( n39646 , n523 );
buf ( n39647 , n549 );
and ( n39648 , n39646 , n39647 );
buf ( n39649 , n39648 );
buf ( n39650 , n39649 );
xor ( n39651 , n39645 , n39650 );
buf ( n39652 , n39651 );
buf ( n39653 , n39652 );
xor ( n39654 , n39634 , n39653 );
buf ( n39655 , n529 );
buf ( n39656 , n545 );
and ( n39657 , n39655 , n39656 );
buf ( n39658 , n39657 );
buf ( n39659 , n39658 );
buf ( n39660 , n525 );
buf ( n39661 , n549 );
and ( n39662 , n39660 , n39661 );
buf ( n39663 , n39662 );
buf ( n39664 , n39663 );
xor ( n39665 , n39659 , n39664 );
buf ( n39666 , n530 );
buf ( n39667 , n544 );
and ( n39668 , n39666 , n39667 );
buf ( n39669 , n39668 );
buf ( n39670 , n39669 );
and ( n39671 , n39665 , n39670 );
and ( n39672 , n39659 , n39664 );
or ( n39673 , n39671 , n39672 );
buf ( n39674 , n39673 );
buf ( n39675 , n39674 );
buf ( n39676 , n531 );
buf ( n39677 , n543 );
and ( n39678 , n39676 , n39677 );
buf ( n39679 , n39678 );
buf ( n39680 , n39679 );
buf ( n39681 , n523 );
buf ( n39682 , n551 );
and ( n39683 , n39681 , n39682 );
buf ( n39684 , n39683 );
buf ( n39685 , n39684 );
xor ( n39686 , n39680 , n39685 );
buf ( n39687 , n526 );
buf ( n39688 , n548 );
and ( n39689 , n39687 , n39688 );
buf ( n39690 , n39689 );
buf ( n39691 , n39690 );
and ( n39692 , n39686 , n39691 );
and ( n39693 , n39680 , n39685 );
or ( n39694 , n39692 , n39693 );
buf ( n39695 , n39694 );
buf ( n39696 , n39695 );
xor ( n39697 , n39675 , n39696 );
buf ( n39698 , n532 );
buf ( n39699 , n542 );
and ( n39700 , n39698 , n39699 );
buf ( n39701 , n39700 );
buf ( n39702 , n39701 );
buf ( n39703 , n533 );
buf ( n39704 , n541 );
and ( n39705 , n39703 , n39704 );
buf ( n39706 , n39705 );
buf ( n39707 , n39706 );
xor ( n39708 , n39702 , n39707 );
buf ( n39709 , n527 );
buf ( n39710 , n547 );
and ( n39711 , n39709 , n39710 );
buf ( n39712 , n39711 );
buf ( n39713 , n39712 );
and ( n39714 , n39708 , n39713 );
and ( n39715 , n39702 , n39707 );
or ( n39716 , n39714 , n39715 );
buf ( n39717 , n39716 );
buf ( n39718 , n39717 );
and ( n39719 , n39697 , n39718 );
and ( n39720 , n39675 , n39696 );
or ( n39721 , n39719 , n39720 );
buf ( n39722 , n39721 );
buf ( n39723 , n39722 );
xor ( n39724 , n39654 , n39723 );
buf ( n39725 , n39724 );
buf ( n39726 , n39725 );
buf ( n39727 , n457 );
buf ( n39728 , n521 );
buf ( n39729 , n552 );
and ( n39730 , n39728 , n39729 );
buf ( n39731 , n39730 );
buf ( n39732 , n39731 );
xor ( n39733 , n39727 , n39732 );
buf ( n39734 , n39733 );
buf ( n39735 , n39734 );
buf ( n39736 , n458 );
buf ( n39737 , n522 );
buf ( n39738 , n552 );
and ( n39739 , n39737 , n39738 );
buf ( n39740 , n39739 );
buf ( n39741 , n39740 );
and ( n39742 , n39736 , n39741 );
buf ( n39743 , n39742 );
buf ( n39744 , n39743 );
xor ( n39745 , n39735 , n39744 );
buf ( n39746 , n524 );
buf ( n39747 , n550 );
and ( n39748 , n39746 , n39747 );
buf ( n39749 , n39748 );
buf ( n39750 , n39749 );
buf ( n39751 , n528 );
buf ( n39752 , n546 );
and ( n39753 , n39751 , n39752 );
buf ( n39754 , n39753 );
buf ( n39755 , n39754 );
xor ( n39756 , n39750 , n39755 );
buf ( n39757 , n536 );
buf ( n39758 , n538 );
and ( n39759 , n39757 , n39758 );
buf ( n39760 , n39759 );
buf ( n39761 , n39760 );
and ( n39762 , n39756 , n39761 );
and ( n39763 , n39750 , n39755 );
or ( n39764 , n39762 , n39763 );
buf ( n39765 , n39764 );
buf ( n39766 , n39765 );
xor ( n39767 , n39745 , n39766 );
buf ( n39768 , n39767 );
buf ( n39769 , n39768 );
xor ( n39770 , n39736 , n39741 );
buf ( n39771 , n39770 );
buf ( n39772 , n39771 );
xor ( n39773 , n36852 , n36857 );
and ( n39774 , n39773 , n36863 );
and ( n39775 , n36852 , n36857 );
or ( n39776 , n39774 , n39775 );
buf ( n39777 , n39776 );
buf ( n39778 , n39777 );
xor ( n39779 , n39772 , n39778 );
xor ( n39780 , n36813 , n36818 );
and ( n39781 , n39780 , n36824 );
and ( n39782 , n36813 , n36818 );
or ( n39783 , n39781 , n39782 );
buf ( n39784 , n39783 );
buf ( n39785 , n39784 );
and ( n39786 , n39779 , n39785 );
and ( n39787 , n39772 , n39778 );
or ( n39788 , n39786 , n39787 );
buf ( n39789 , n39788 );
buf ( n39790 , n39789 );
xor ( n39791 , n39769 , n39790 );
xor ( n39792 , n39702 , n39707 );
xor ( n39793 , n39792 , n39713 );
buf ( n39794 , n39793 );
buf ( n39795 , n39794 );
xor ( n39796 , n39659 , n39664 );
xor ( n39797 , n39796 , n39670 );
buf ( n39798 , n39797 );
buf ( n39799 , n39798 );
xor ( n39800 , n39795 , n39799 );
xor ( n39801 , n39680 , n39685 );
xor ( n39802 , n39801 , n39691 );
buf ( n39803 , n39802 );
buf ( n39804 , n39803 );
and ( n39805 , n39800 , n39804 );
and ( n39806 , n39795 , n39799 );
or ( n39807 , n39805 , n39806 );
buf ( n39808 , n39807 );
buf ( n39809 , n39808 );
and ( n39810 , n39791 , n39809 );
and ( n39811 , n39769 , n39790 );
or ( n39812 , n39810 , n39811 );
buf ( n39813 , n39812 );
buf ( n39814 , n39813 );
xor ( n39815 , n39726 , n39814 );
xor ( n39816 , n39675 , n39696 );
xor ( n39817 , n39816 , n39718 );
buf ( n39818 , n39817 );
buf ( n39819 , n39818 );
xor ( n39820 , n36871 , n36876 );
and ( n39821 , n39820 , n36882 );
and ( n39822 , n36871 , n36876 );
or ( n39823 , n39821 , n39822 );
buf ( n39824 , n39823 );
buf ( n39825 , n39824 );
xor ( n39826 , n36793 , n36798 );
and ( n39827 , n39826 , n36804 );
and ( n39828 , n36793 , n36798 );
or ( n39829 , n39827 , n39828 );
buf ( n39830 , n39829 );
buf ( n39831 , n39830 );
xor ( n39832 , n39825 , n39831 );
xor ( n39833 , n39750 , n39755 );
xor ( n39834 , n39833 , n39761 );
buf ( n39835 , n39834 );
buf ( n39836 , n39835 );
and ( n39837 , n39832 , n39836 );
and ( n39838 , n39825 , n39831 );
or ( n39839 , n39837 , n39838 );
buf ( n39840 , n39839 );
buf ( n39841 , n39840 );
xor ( n39842 , n39819 , n39841 );
buf ( n39843 , n529 );
buf ( n39844 , n544 );
and ( n39845 , n39843 , n39844 );
buf ( n39846 , n39845 );
buf ( n39847 , n39846 );
buf ( n39848 , n530 );
buf ( n39849 , n543 );
and ( n39850 , n39848 , n39849 );
buf ( n39851 , n39850 );
buf ( n39852 , n39851 );
xor ( n39853 , n39847 , n39852 );
buf ( n39854 , n522 );
buf ( n39855 , n551 );
and ( n39856 , n39854 , n39855 );
buf ( n39857 , n39856 );
buf ( n39858 , n39857 );
xor ( n39859 , n39853 , n39858 );
buf ( n39860 , n39859 );
buf ( n39861 , n39860 );
buf ( n39862 , n525 );
buf ( n39863 , n548 );
and ( n39864 , n39862 , n39863 );
buf ( n39865 , n39864 );
buf ( n39866 , n39865 );
buf ( n39867 , n531 );
buf ( n39868 , n542 );
and ( n39869 , n39867 , n39868 );
buf ( n39870 , n39869 );
buf ( n39871 , n39870 );
xor ( n39872 , n39866 , n39871 );
buf ( n39873 , n532 );
buf ( n39874 , n541 );
and ( n39875 , n39873 , n39874 );
buf ( n39876 , n39875 );
buf ( n39877 , n39876 );
xor ( n39878 , n39872 , n39877 );
buf ( n39879 , n39878 );
buf ( n39880 , n39879 );
xor ( n39881 , n39861 , n39880 );
buf ( n39882 , n534 );
buf ( n39883 , n540 );
and ( n39884 , n39882 , n39883 );
buf ( n39885 , n39884 );
buf ( n39886 , n39885 );
buf ( n39887 , n535 );
buf ( n39888 , n539 );
and ( n39889 , n39887 , n39888 );
buf ( n39890 , n39889 );
buf ( n39891 , n39890 );
xor ( n39892 , n39886 , n39891 );
and ( n39893 , n36892 , n36897 );
buf ( n39894 , n39893 );
buf ( n39895 , n39894 );
and ( n39896 , n39892 , n39895 );
and ( n39897 , n39886 , n39891 );
or ( n39898 , n39896 , n39897 );
buf ( n39899 , n39898 );
buf ( n39900 , n39899 );
xor ( n39901 , n39881 , n39900 );
buf ( n39902 , n39901 );
buf ( n39903 , n39902 );
and ( n39904 , n39842 , n39903 );
and ( n39905 , n39819 , n39841 );
or ( n39906 , n39904 , n39905 );
buf ( n39907 , n39906 );
buf ( n39908 , n39907 );
xor ( n39909 , n39815 , n39908 );
buf ( n39910 , n39909 );
buf ( n39911 , n39910 );
xor ( n39912 , n39769 , n39790 );
xor ( n39913 , n39912 , n39809 );
buf ( n39914 , n39913 );
buf ( n39915 , n39914 );
xor ( n39916 , n39819 , n39841 );
xor ( n39917 , n39916 , n39903 );
buf ( n39918 , n39917 );
buf ( n39919 , n39918 );
xor ( n39920 , n39915 , n39919 );
xor ( n39921 , n39795 , n39799 );
xor ( n39922 , n39921 , n39804 );
buf ( n39923 , n39922 );
buf ( n39924 , n39923 );
xor ( n39925 , n36866 , n36885 );
and ( n39926 , n39925 , n36907 );
and ( n39927 , n36866 , n36885 );
or ( n39928 , n39926 , n39927 );
buf ( n39929 , n39928 );
buf ( n39930 , n39929 );
xor ( n39931 , n39924 , n39930 );
xor ( n39932 , n39886 , n39891 );
xor ( n39933 , n39932 , n39895 );
buf ( n39934 , n39933 );
buf ( n39935 , n39934 );
xor ( n39936 , n36891 , n36900 );
and ( n39937 , n39936 , n36904 );
and ( n39938 , n36891 , n36900 );
or ( n39939 , n39937 , n39938 );
buf ( n39940 , n39939 );
buf ( n39941 , n39940 );
xor ( n39942 , n39935 , n39941 );
xor ( n39943 , n36766 , n36772 );
and ( n39944 , n39943 , n36779 );
and ( n39945 , n36766 , n36772 );
or ( n39946 , n39944 , n39945 );
buf ( n39947 , n39946 );
buf ( n39948 , n39947 );
xor ( n39949 , n39942 , n39948 );
buf ( n39950 , n39949 );
buf ( n39951 , n39950 );
and ( n39952 , n39931 , n39951 );
and ( n39953 , n39924 , n39930 );
or ( n39954 , n39952 , n39953 );
buf ( n39955 , n39954 );
buf ( n39956 , n39955 );
and ( n39957 , n39920 , n39956 );
and ( n39958 , n39915 , n39919 );
or ( n39959 , n39957 , n39958 );
buf ( n39960 , n39959 );
buf ( n39961 , n39960 );
xor ( n39962 , n39911 , n39961 );
xor ( n39963 , n39735 , n39744 );
and ( n39964 , n39963 , n39766 );
and ( n39965 , n39735 , n39744 );
or ( n39966 , n39964 , n39965 );
buf ( n39967 , n39966 );
buf ( n39968 , n39967 );
xor ( n39969 , n39847 , n39852 );
and ( n39970 , n39969 , n39858 );
and ( n39971 , n39847 , n39852 );
or ( n39972 , n39970 , n39971 );
buf ( n39973 , n39972 );
buf ( n39974 , n39973 );
xor ( n39975 , n39866 , n39871 );
and ( n39976 , n39975 , n39877 );
and ( n39977 , n39866 , n39871 );
or ( n39978 , n39976 , n39977 );
buf ( n39979 , n39978 );
buf ( n39980 , n39979 );
xor ( n39981 , n39974 , n39980 );
buf ( n39982 , n526 );
buf ( n39983 , n547 );
and ( n39984 , n39982 , n39983 );
buf ( n39985 , n39984 );
buf ( n39986 , n39985 );
buf ( n39987 , n533 );
buf ( n39988 , n540 );
and ( n39989 , n39987 , n39988 );
buf ( n39990 , n39989 );
buf ( n39991 , n39990 );
xor ( n39992 , n39986 , n39991 );
buf ( n39993 , n534 );
buf ( n39994 , n539 );
and ( n39995 , n39993 , n39994 );
buf ( n39996 , n39995 );
buf ( n39997 , n39996 );
and ( n39998 , n39992 , n39997 );
and ( n39999 , n39986 , n39991 );
or ( n40000 , n39998 , n39999 );
buf ( n40001 , n40000 );
buf ( n40002 , n40001 );
xor ( n40003 , n39981 , n40002 );
buf ( n40004 , n40003 );
buf ( n40005 , n40004 );
xor ( n40006 , n39968 , n40005 );
and ( n40007 , n39727 , n39732 );
buf ( n40008 , n40007 );
buf ( n40009 , n40008 );
buf ( n40010 , n523 );
buf ( n40011 , n550 );
and ( n40012 , n40010 , n40011 );
buf ( n40013 , n40012 );
buf ( n40014 , n40013 );
buf ( n40015 , n527 );
buf ( n40016 , n546 );
and ( n40017 , n40015 , n40016 );
buf ( n40018 , n40017 );
buf ( n40019 , n40018 );
xor ( n40020 , n40014 , n40019 );
buf ( n40021 , n535 );
buf ( n40022 , n538 );
and ( n40023 , n40021 , n40022 );
buf ( n40024 , n40023 );
buf ( n40025 , n40024 );
and ( n40026 , n40020 , n40025 );
and ( n40027 , n40014 , n40019 );
or ( n40028 , n40026 , n40027 );
buf ( n40029 , n40028 );
buf ( n40030 , n40029 );
xor ( n40031 , n40009 , n40030 );
buf ( n40032 , n536 );
buf ( n40033 , n537 );
and ( n40034 , n40032 , n40033 );
buf ( n40035 , n40034 );
buf ( n40036 , n40035 );
buf ( n40037 , n528 );
buf ( n40038 , n545 );
and ( n40039 , n40037 , n40038 );
buf ( n40040 , n40039 );
buf ( n40041 , n40040 );
xor ( n40042 , n40036 , n40041 );
buf ( n40043 , n524 );
buf ( n40044 , n549 );
and ( n40045 , n40043 , n40044 );
buf ( n40046 , n40045 );
buf ( n40047 , n40046 );
and ( n40048 , n40042 , n40047 );
and ( n40049 , n40036 , n40041 );
or ( n40050 , n40048 , n40049 );
buf ( n40051 , n40050 );
buf ( n40052 , n40051 );
xor ( n40053 , n40031 , n40052 );
buf ( n40054 , n40053 );
buf ( n40055 , n40054 );
xor ( n40056 , n40006 , n40055 );
buf ( n40057 , n40056 );
buf ( n40058 , n40057 );
xor ( n40059 , n39986 , n39991 );
xor ( n40060 , n40059 , n39997 );
buf ( n40061 , n40060 );
buf ( n40062 , n40061 );
xor ( n40063 , n40014 , n40019 );
xor ( n40064 , n40063 , n40025 );
buf ( n40065 , n40064 );
buf ( n40066 , n40065 );
xor ( n40067 , n40062 , n40066 );
xor ( n40068 , n40036 , n40041 );
xor ( n40069 , n40068 , n40047 );
buf ( n40070 , n40069 );
buf ( n40071 , n40070 );
and ( n40072 , n40067 , n40071 );
and ( n40073 , n40062 , n40066 );
or ( n40074 , n40072 , n40073 );
buf ( n40075 , n40074 );
buf ( n40076 , n40075 );
xor ( n40077 , n39861 , n39880 );
and ( n40078 , n40077 , n39900 );
and ( n40079 , n39861 , n39880 );
or ( n40080 , n40078 , n40079 );
buf ( n40081 , n40080 );
buf ( n40082 , n40081 );
xor ( n40083 , n40076 , n40082 );
buf ( n40084 , n521 );
buf ( n40085 , n551 );
and ( n40086 , n40084 , n40085 );
buf ( n40087 , n40086 );
buf ( n40088 , n40087 );
buf ( n40089 , n522 );
buf ( n40090 , n550 );
and ( n40091 , n40089 , n40090 );
buf ( n40092 , n40091 );
buf ( n40093 , n40092 );
xor ( n40094 , n40088 , n40093 );
buf ( n40095 , n524 );
buf ( n40096 , n548 );
and ( n40097 , n40095 , n40096 );
buf ( n40098 , n40097 );
buf ( n40099 , n40098 );
xor ( n40100 , n40094 , n40099 );
buf ( n40101 , n40100 );
buf ( n40102 , n40101 );
buf ( n40103 , n528 );
buf ( n40104 , n544 );
and ( n40105 , n40103 , n40104 );
buf ( n40106 , n40105 );
buf ( n40107 , n40106 );
buf ( n40108 , n529 );
buf ( n40109 , n543 );
and ( n40110 , n40108 , n40109 );
buf ( n40111 , n40110 );
buf ( n40112 , n40111 );
xor ( n40113 , n40107 , n40112 );
buf ( n40114 , n525 );
buf ( n40115 , n547 );
and ( n40116 , n40114 , n40115 );
buf ( n40117 , n40116 );
buf ( n40118 , n40117 );
xor ( n40119 , n40113 , n40118 );
buf ( n40120 , n40119 );
buf ( n40121 , n40120 );
xor ( n40122 , n40102 , n40121 );
buf ( n40123 , n527 );
buf ( n40124 , n545 );
and ( n40125 , n40123 , n40124 );
buf ( n40126 , n40125 );
buf ( n40127 , n40126 );
buf ( n40128 , n534 );
buf ( n40129 , n538 );
and ( n40130 , n40128 , n40129 );
buf ( n40131 , n40130 );
buf ( n40132 , n40131 );
xor ( n40133 , n40127 , n40132 );
buf ( n40134 , n535 );
buf ( n40135 , n537 );
and ( n40136 , n40134 , n40135 );
buf ( n40137 , n40136 );
buf ( n40138 , n40137 );
xor ( n40139 , n40133 , n40138 );
buf ( n40140 , n40139 );
buf ( n40141 , n40140 );
xor ( n40142 , n40122 , n40141 );
buf ( n40143 , n40142 );
buf ( n40144 , n40143 );
xor ( n40145 , n40083 , n40144 );
buf ( n40146 , n40145 );
buf ( n40147 , n40146 );
xor ( n40148 , n40058 , n40147 );
xor ( n40149 , n40062 , n40066 );
xor ( n40150 , n40149 , n40071 );
buf ( n40151 , n40150 );
buf ( n40152 , n40151 );
xor ( n40153 , n39935 , n39941 );
and ( n40154 , n40153 , n39948 );
and ( n40155 , n39935 , n39941 );
or ( n40156 , n40154 , n40155 );
buf ( n40157 , n40156 );
buf ( n40158 , n40157 );
xor ( n40159 , n40152 , n40158 );
xor ( n40160 , n39772 , n39778 );
xor ( n40161 , n40160 , n39785 );
buf ( n40162 , n40161 );
buf ( n40163 , n40162 );
xor ( n40164 , n36788 , n36807 );
and ( n40165 , n40164 , n36827 );
and ( n40166 , n36788 , n36807 );
or ( n40167 , n40165 , n40166 );
buf ( n40168 , n40167 );
buf ( n40169 , n40168 );
xor ( n40170 , n40163 , n40169 );
xor ( n40171 , n39825 , n39831 );
xor ( n40172 , n40171 , n39836 );
buf ( n40173 , n40172 );
buf ( n40174 , n40173 );
and ( n40175 , n40170 , n40174 );
and ( n40176 , n40163 , n40169 );
or ( n40177 , n40175 , n40176 );
buf ( n40178 , n40177 );
buf ( n40179 , n40178 );
and ( n40180 , n40159 , n40179 );
and ( n40181 , n40152 , n40158 );
or ( n40182 , n40180 , n40181 );
buf ( n40183 , n40182 );
buf ( n40184 , n40183 );
xor ( n40185 , n40148 , n40184 );
buf ( n40186 , n40185 );
buf ( n40187 , n40186 );
xor ( n40188 , n39962 , n40187 );
buf ( n40189 , n40188 );
buf ( n40190 , n40189 );
xor ( n40191 , n40152 , n40158 );
xor ( n40192 , n40191 , n40179 );
buf ( n40193 , n40192 );
buf ( n40194 , n40193 );
xor ( n40195 , n39915 , n39919 );
xor ( n40196 , n40195 , n39956 );
buf ( n40197 , n40196 );
buf ( n40198 , n40197 );
xor ( n40199 , n40194 , n40198 );
xor ( n40200 , n36923 , n36929 );
and ( n40201 , n40200 , n36936 );
and ( n40202 , n36923 , n36929 );
or ( n40203 , n40201 , n40202 );
buf ( n40204 , n40203 );
buf ( n40205 , n40204 );
xor ( n40206 , n40163 , n40169 );
xor ( n40207 , n40206 , n40174 );
buf ( n40208 , n40207 );
buf ( n40209 , n40208 );
xor ( n40210 , n40205 , n40209 );
xor ( n40211 , n36782 , n36830 );
and ( n40212 , n40211 , n36837 );
and ( n40213 , n36782 , n36830 );
or ( n40214 , n40212 , n40213 );
buf ( n40215 , n40214 );
buf ( n40216 , n40215 );
and ( n40217 , n40210 , n40216 );
and ( n40218 , n40205 , n40209 );
or ( n40219 , n40217 , n40218 );
buf ( n40220 , n40219 );
buf ( n40221 , n40220 );
and ( n40222 , n40199 , n40221 );
and ( n40223 , n40194 , n40198 );
or ( n40224 , n40222 , n40223 );
buf ( n40225 , n40224 );
buf ( n40226 , n40225 );
or ( n40227 , n40190 , n40226 );
buf ( n40228 , n40227 );
not ( n40229 , n40228 );
xor ( n40230 , n39726 , n39814 );
and ( n40231 , n40230 , n39908 );
and ( n40232 , n39726 , n39814 );
or ( n40233 , n40231 , n40232 );
buf ( n40234 , n40233 );
buf ( n40235 , n40234 );
xor ( n40236 , n40058 , n40147 );
and ( n40237 , n40236 , n40184 );
and ( n40238 , n40058 , n40147 );
or ( n40239 , n40237 , n40238 );
buf ( n40240 , n40239 );
buf ( n40241 , n40240 );
xor ( n40242 , n40235 , n40241 );
xor ( n40243 , n40076 , n40082 );
and ( n40244 , n40243 , n40144 );
and ( n40245 , n40076 , n40082 );
or ( n40246 , n40244 , n40245 );
buf ( n40247 , n40246 );
buf ( n40248 , n40247 );
xor ( n40249 , n40102 , n40121 );
and ( n40250 , n40249 , n40141 );
and ( n40251 , n40102 , n40121 );
or ( n40252 , n40250 , n40251 );
buf ( n40253 , n40252 );
buf ( n40254 , n40253 );
xor ( n40255 , n40088 , n40093 );
and ( n40256 , n40255 , n40099 );
and ( n40257 , n40088 , n40093 );
or ( n40258 , n40256 , n40257 );
buf ( n40259 , n40258 );
buf ( n40260 , n40259 );
buf ( n40261 , n528 );
buf ( n40262 , n543 );
and ( n40263 , n40261 , n40262 );
buf ( n40264 , n40263 );
buf ( n40265 , n40264 );
buf ( n40266 , n529 );
buf ( n40267 , n542 );
and ( n40268 , n40266 , n40267 );
buf ( n40269 , n40268 );
buf ( n40270 , n40269 );
xor ( n40271 , n40265 , n40270 );
buf ( n40272 , n525 );
buf ( n40273 , n546 );
and ( n40274 , n40272 , n40273 );
buf ( n40275 , n40274 );
buf ( n40276 , n40275 );
xor ( n40277 , n40271 , n40276 );
buf ( n40278 , n40277 );
buf ( n40279 , n40278 );
xor ( n40280 , n40260 , n40279 );
buf ( n40281 , n521 );
buf ( n40282 , n550 );
and ( n40283 , n40281 , n40282 );
buf ( n40284 , n40283 );
buf ( n40285 , n40284 );
buf ( n40286 , n522 );
buf ( n40287 , n549 );
and ( n40288 , n40286 , n40287 );
buf ( n40289 , n40288 );
buf ( n40290 , n40289 );
xor ( n40291 , n40285 , n40290 );
buf ( n40292 , n524 );
buf ( n40293 , n547 );
and ( n40294 , n40292 , n40293 );
buf ( n40295 , n40294 );
buf ( n40296 , n40295 );
xor ( n40297 , n40291 , n40296 );
buf ( n40298 , n40297 );
buf ( n40299 , n40298 );
xor ( n40300 , n40280 , n40299 );
buf ( n40301 , n40300 );
buf ( n40302 , n40301 );
xor ( n40303 , n40254 , n40302 );
buf ( n40304 , n526 );
buf ( n40305 , n545 );
and ( n40306 , n40304 , n40305 );
buf ( n40307 , n40306 );
buf ( n40308 , n40307 );
buf ( n40309 , n532 );
buf ( n40310 , n539 );
and ( n40311 , n40309 , n40310 );
buf ( n40312 , n40311 );
buf ( n40313 , n40312 );
xor ( n40314 , n40308 , n40313 );
buf ( n40315 , n533 );
buf ( n40316 , n538 );
and ( n40317 , n40315 , n40316 );
buf ( n40318 , n40317 );
buf ( n40319 , n40318 );
xor ( n40320 , n40314 , n40319 );
buf ( n40321 , n40320 );
buf ( n40322 , n40321 );
buf ( n40323 , n530 );
buf ( n40324 , n541 );
and ( n40325 , n40323 , n40324 );
buf ( n40326 , n40325 );
buf ( n40327 , n40326 );
buf ( n40328 , n531 );
buf ( n40329 , n540 );
and ( n40330 , n40328 , n40329 );
buf ( n40331 , n40330 );
buf ( n40332 , n40331 );
xor ( n40333 , n40327 , n40332 );
buf ( n40334 , n523 );
buf ( n40335 , n548 );
and ( n40336 , n40334 , n40335 );
buf ( n40337 , n40336 );
buf ( n40338 , n40337 );
xor ( n40339 , n40333 , n40338 );
buf ( n40340 , n40339 );
buf ( n40341 , n40340 );
xor ( n40342 , n40322 , n40341 );
buf ( n40343 , n527 );
buf ( n40344 , n544 );
and ( n40345 , n40343 , n40344 );
buf ( n40346 , n40345 );
buf ( n40347 , n40346 );
buf ( n40348 , n534 );
buf ( n40349 , n537 );
and ( n40350 , n40348 , n40349 );
buf ( n40351 , n40350 );
buf ( n40352 , n40351 );
xor ( n40353 , n40347 , n40352 );
xor ( n40354 , n40127 , n40132 );
and ( n40355 , n40354 , n40138 );
and ( n40356 , n40127 , n40132 );
or ( n40357 , n40355 , n40356 );
buf ( n40358 , n40357 );
buf ( n40359 , n40358 );
xor ( n40360 , n40353 , n40359 );
buf ( n40361 , n40360 );
buf ( n40362 , n40361 );
xor ( n40363 , n40342 , n40362 );
buf ( n40364 , n40363 );
buf ( n40365 , n40364 );
xor ( n40366 , n40303 , n40365 );
buf ( n40367 , n40366 );
buf ( n40368 , n40367 );
xor ( n40369 , n40248 , n40368 );
xor ( n40370 , n39634 , n39653 );
and ( n40371 , n40370 , n39723 );
and ( n40372 , n39634 , n39653 );
or ( n40373 , n40371 , n40372 );
buf ( n40374 , n40373 );
buf ( n40375 , n40374 );
xor ( n40376 , n40009 , n40030 );
and ( n40377 , n40376 , n40052 );
and ( n40378 , n40009 , n40030 );
or ( n40379 , n40377 , n40378 );
buf ( n40380 , n40379 );
buf ( n40381 , n40380 );
xor ( n40382 , n39974 , n39980 );
and ( n40383 , n40382 , n40002 );
and ( n40384 , n39974 , n39980 );
or ( n40385 , n40383 , n40384 );
buf ( n40386 , n40385 );
buf ( n40387 , n40386 );
xor ( n40388 , n40381 , n40387 );
xor ( n40389 , n40107 , n40112 );
and ( n40390 , n40389 , n40118 );
and ( n40391 , n40107 , n40112 );
or ( n40392 , n40390 , n40391 );
buf ( n40393 , n40392 );
buf ( n40394 , n40393 );
xor ( n40395 , n39639 , n39644 );
and ( n40396 , n40395 , n39650 );
and ( n40397 , n39639 , n39644 );
or ( n40398 , n40396 , n40397 );
buf ( n40399 , n40398 );
buf ( n40400 , n40399 );
xor ( n40401 , n40394 , n40400 );
xor ( n40402 , n39620 , n39625 );
and ( n40403 , n40402 , n39631 );
and ( n40404 , n39620 , n39625 );
or ( n40405 , n40403 , n40404 );
buf ( n40406 , n40405 );
buf ( n40407 , n40406 );
xor ( n40408 , n40401 , n40407 );
buf ( n40409 , n40408 );
buf ( n40410 , n40409 );
xor ( n40411 , n40388 , n40410 );
buf ( n40412 , n40411 );
buf ( n40413 , n40412 );
xor ( n40414 , n40375 , n40413 );
xor ( n40415 , n39968 , n40005 );
and ( n40416 , n40415 , n40055 );
and ( n40417 , n39968 , n40005 );
or ( n40418 , n40416 , n40417 );
buf ( n40419 , n40418 );
buf ( n40420 , n40419 );
xor ( n40421 , n40414 , n40420 );
buf ( n40422 , n40421 );
buf ( n40423 , n40422 );
xor ( n40424 , n40369 , n40423 );
buf ( n40425 , n40424 );
buf ( n40426 , n40425 );
xor ( n40427 , n40242 , n40426 );
buf ( n40428 , n40427 );
not ( n40429 , n40428 );
xor ( n40430 , n39911 , n39961 );
and ( n40431 , n40430 , n40187 );
and ( n40432 , n39911 , n39961 );
or ( n40433 , n40431 , n40432 );
buf ( n40434 , n40433 );
not ( n40435 , n40434 );
nand ( n40436 , n40429 , n40435 );
not ( n40437 , n40436 );
nor ( n40438 , n40229 , n40437 );
not ( n40439 , n40438 );
xor ( n40440 , n40194 , n40198 );
xor ( n40441 , n40440 , n40221 );
buf ( n40442 , n40441 );
buf ( n40443 , n40442 );
xor ( n40444 , n39924 , n39930 );
xor ( n40445 , n40444 , n39951 );
buf ( n40446 , n40445 );
buf ( n40447 , n40446 );
xor ( n40448 , n36910 , n36916 );
and ( n40449 , n40448 , n36939 );
and ( n40450 , n36910 , n36916 );
or ( n40451 , n40449 , n40450 );
buf ( n40452 , n40451 );
buf ( n40453 , n40452 );
xor ( n40454 , n40447 , n40453 );
xor ( n40455 , n40205 , n40209 );
xor ( n40456 , n40455 , n40216 );
buf ( n40457 , n40456 );
buf ( n40458 , n40457 );
and ( n40459 , n40454 , n40458 );
and ( n40460 , n40447 , n40453 );
or ( n40461 , n40459 , n40460 );
buf ( n40462 , n40461 );
buf ( n40463 , n40462 );
nor ( n40464 , n40443 , n40463 );
buf ( n40465 , n40464 );
xor ( n40466 , n36840 , n36846 );
and ( n40467 , n40466 , n36942 );
and ( n40468 , n36840 , n36846 );
or ( n40469 , n40467 , n40468 );
buf ( n40470 , n40469 );
buf ( n40471 , n40470 );
xor ( n40472 , n40447 , n40453 );
xor ( n40473 , n40472 , n40458 );
buf ( n40474 , n40473 );
buf ( n40475 , n40474 );
nand ( n40476 , n40471 , n40475 );
buf ( n40477 , n40476 );
or ( n40478 , n40465 , n40477 );
buf ( n40479 , n40442 );
buf ( n40480 , n40462 );
nand ( n40481 , n40479 , n40480 );
buf ( n40482 , n40481 );
nand ( n40483 , n40478 , n40482 );
not ( n40484 , n40483 );
xor ( n40485 , n36760 , n36945 );
and ( n40486 , n40485 , n36955 );
and ( n40487 , n36760 , n36945 );
or ( n40488 , n40486 , n40487 );
buf ( n40489 , n40488 );
buf ( n40490 , n40489 );
buf ( n40491 , n40465 );
buf ( n40492 , n40470 );
buf ( n40493 , n40474 );
nor ( n40494 , n40492 , n40493 );
buf ( n40495 , n40494 );
buf ( n40496 , n40495 );
nor ( n40497 , n40491 , n40496 );
buf ( n40498 , n40497 );
buf ( n40499 , n40498 );
nand ( n40500 , n40490 , n40499 );
buf ( n40501 , n40500 );
nand ( n40502 , n40484 , n40501 );
not ( n40503 , n40502 );
or ( n40504 , n40439 , n40503 );
and ( n40505 , n40189 , n40225 );
not ( n40506 , n40505 );
not ( n40507 , n40436 );
or ( n40508 , n40506 , n40507 );
buf ( n40509 , n40428 );
buf ( n40510 , n40434 );
nand ( n40511 , n40509 , n40510 );
buf ( n40512 , n40511 );
nand ( n40513 , n40508 , n40512 );
buf ( n40514 , n40513 );
not ( n40515 , n40514 );
buf ( n40516 , n40515 );
nand ( n40517 , n40504 , n40516 );
not ( n40518 , n40517 );
buf ( n40519 , n530 );
buf ( n40520 , n540 );
and ( n40521 , n40519 , n40520 );
buf ( n40522 , n40521 );
buf ( n40523 , n40522 );
buf ( n40524 , n531 );
buf ( n40525 , n539 );
and ( n40526 , n40524 , n40525 );
buf ( n40527 , n40526 );
buf ( n40528 , n40527 );
xor ( n40529 , n40523 , n40528 );
buf ( n40530 , n523 );
buf ( n40531 , n547 );
and ( n40532 , n40530 , n40531 );
buf ( n40533 , n40532 );
buf ( n40534 , n40533 );
and ( n40535 , n40529 , n40534 );
and ( n40536 , n40523 , n40528 );
or ( n40537 , n40535 , n40536 );
buf ( n40538 , n40537 );
buf ( n40539 , n40538 );
buf ( n40540 , n530 );
buf ( n40541 , n539 );
and ( n40542 , n40540 , n40541 );
buf ( n40543 , n40542 );
buf ( n40544 , n40543 );
buf ( n40545 , n531 );
buf ( n40546 , n538 );
and ( n40547 , n40545 , n40546 );
buf ( n40548 , n40547 );
buf ( n40549 , n40548 );
xor ( n40550 , n40544 , n40549 );
buf ( n40551 , n523 );
buf ( n40552 , n546 );
and ( n40553 , n40551 , n40552 );
buf ( n40554 , n40553 );
buf ( n40555 , n40554 );
xor ( n40556 , n40550 , n40555 );
buf ( n40557 , n40556 );
buf ( n40558 , n40557 );
xor ( n40559 , n40539 , n40558 );
buf ( n40560 , n526 );
buf ( n40561 , n543 );
and ( n40562 , n40560 , n40561 );
buf ( n40563 , n40562 );
buf ( n40564 , n40563 );
buf ( n40565 , n532 );
buf ( n40566 , n537 );
and ( n40567 , n40565 , n40566 );
buf ( n40568 , n40567 );
buf ( n40569 , n40568 );
xor ( n40570 , n40564 , n40569 );
buf ( n40571 , n527 );
buf ( n40572 , n542 );
and ( n40573 , n40571 , n40572 );
buf ( n40574 , n40573 );
buf ( n40575 , n40574 );
xor ( n40576 , n40570 , n40575 );
buf ( n40577 , n40576 );
buf ( n40578 , n40577 );
xor ( n40579 , n40559 , n40578 );
buf ( n40580 , n40579 );
buf ( n40581 , n40580 );
buf ( n40582 , n521 );
buf ( n40583 , n548 );
and ( n40584 , n40582 , n40583 );
buf ( n40585 , n40584 );
buf ( n40586 , n40585 );
buf ( n40587 , n522 );
buf ( n40588 , n547 );
and ( n40589 , n40587 , n40588 );
buf ( n40590 , n40589 );
buf ( n40591 , n40590 );
xor ( n40592 , n40586 , n40591 );
buf ( n40593 , n524 );
buf ( n40594 , n545 );
and ( n40595 , n40593 , n40594 );
buf ( n40596 , n40595 );
buf ( n40597 , n40596 );
xor ( n40598 , n40592 , n40597 );
buf ( n40599 , n40598 );
buf ( n40600 , n40599 );
buf ( n40601 , n528 );
buf ( n40602 , n541 );
and ( n40603 , n40601 , n40602 );
buf ( n40604 , n40603 );
buf ( n40605 , n40604 );
buf ( n40606 , n529 );
buf ( n40607 , n540 );
and ( n40608 , n40606 , n40607 );
buf ( n40609 , n40608 );
buf ( n40610 , n40609 );
xor ( n40611 , n40605 , n40610 );
buf ( n40612 , n525 );
buf ( n40613 , n544 );
and ( n40614 , n40612 , n40613 );
buf ( n40615 , n40614 );
buf ( n40616 , n40615 );
xor ( n40617 , n40611 , n40616 );
buf ( n40618 , n40617 );
buf ( n40619 , n40618 );
xor ( n40620 , n40600 , n40619 );
buf ( n40621 , n527 );
buf ( n40622 , n543 );
and ( n40623 , n40621 , n40622 );
buf ( n40624 , n40623 );
buf ( n40625 , n40624 );
xor ( n40626 , n40327 , n40332 );
and ( n40627 , n40626 , n40338 );
and ( n40628 , n40327 , n40332 );
or ( n40629 , n40627 , n40628 );
buf ( n40630 , n40629 );
buf ( n40631 , n40630 );
xor ( n40632 , n40625 , n40631 );
xor ( n40633 , n40308 , n40313 );
and ( n40634 , n40633 , n40319 );
and ( n40635 , n40308 , n40313 );
or ( n40636 , n40634 , n40635 );
buf ( n40637 , n40636 );
buf ( n40638 , n40637 );
and ( n40639 , n40632 , n40638 );
and ( n40640 , n40625 , n40631 );
or ( n40641 , n40639 , n40640 );
buf ( n40642 , n40641 );
buf ( n40643 , n40642 );
xor ( n40644 , n40620 , n40643 );
buf ( n40645 , n40644 );
buf ( n40646 , n40645 );
xor ( n40647 , n40581 , n40646 );
xor ( n40648 , n40347 , n40352 );
and ( n40649 , n40648 , n40359 );
and ( n40650 , n40347 , n40352 );
or ( n40651 , n40649 , n40650 );
buf ( n40652 , n40651 );
buf ( n40653 , n40652 );
xor ( n40654 , n40394 , n40400 );
and ( n40655 , n40654 , n40407 );
and ( n40656 , n40394 , n40400 );
or ( n40657 , n40655 , n40656 );
buf ( n40658 , n40657 );
buf ( n40659 , n40658 );
xor ( n40660 , n40653 , n40659 );
xor ( n40661 , n40625 , n40631 );
xor ( n40662 , n40661 , n40638 );
buf ( n40663 , n40662 );
buf ( n40664 , n40663 );
and ( n40665 , n40660 , n40664 );
and ( n40666 , n40653 , n40659 );
or ( n40667 , n40665 , n40666 );
buf ( n40668 , n40667 );
buf ( n40669 , n40668 );
xor ( n40670 , n40647 , n40669 );
buf ( n40671 , n40670 );
buf ( n40672 , n40671 );
buf ( n40673 , n526 );
buf ( n40674 , n544 );
and ( n40675 , n40673 , n40674 );
buf ( n40676 , n40675 );
buf ( n40677 , n40676 );
buf ( n40678 , n532 );
buf ( n40679 , n538 );
and ( n40680 , n40678 , n40679 );
buf ( n40681 , n40680 );
buf ( n40682 , n40681 );
xor ( n40683 , n40677 , n40682 );
buf ( n40684 , n533 );
buf ( n40685 , n537 );
and ( n40686 , n40684 , n40685 );
buf ( n40687 , n40686 );
buf ( n40688 , n40687 );
and ( n40689 , n40683 , n40688 );
and ( n40690 , n40677 , n40682 );
or ( n40691 , n40689 , n40690 );
buf ( n40692 , n40691 );
buf ( n40693 , n40692 );
buf ( n40694 , n521 );
buf ( n40695 , n549 );
and ( n40696 , n40694 , n40695 );
buf ( n40697 , n40696 );
buf ( n40698 , n40697 );
buf ( n40699 , n522 );
buf ( n40700 , n548 );
and ( n40701 , n40699 , n40700 );
buf ( n40702 , n40701 );
buf ( n40703 , n40702 );
xor ( n40704 , n40698 , n40703 );
buf ( n40705 , n524 );
buf ( n40706 , n546 );
and ( n40707 , n40705 , n40706 );
buf ( n40708 , n40707 );
buf ( n40709 , n40708 );
and ( n40710 , n40704 , n40709 );
and ( n40711 , n40698 , n40703 );
or ( n40712 , n40710 , n40711 );
buf ( n40713 , n40712 );
buf ( n40714 , n40713 );
xor ( n40715 , n40693 , n40714 );
buf ( n40716 , n528 );
buf ( n40717 , n542 );
and ( n40718 , n40716 , n40717 );
buf ( n40719 , n40718 );
buf ( n40720 , n40719 );
buf ( n40721 , n529 );
buf ( n40722 , n541 );
and ( n40723 , n40721 , n40722 );
buf ( n40724 , n40723 );
buf ( n40725 , n40724 );
xor ( n40726 , n40720 , n40725 );
buf ( n40727 , n525 );
buf ( n40728 , n545 );
and ( n40729 , n40727 , n40728 );
buf ( n40730 , n40729 );
buf ( n40731 , n40730 );
and ( n40732 , n40726 , n40731 );
and ( n40733 , n40720 , n40725 );
or ( n40734 , n40732 , n40733 );
buf ( n40735 , n40734 );
buf ( n40736 , n40735 );
xor ( n40737 , n40715 , n40736 );
buf ( n40738 , n40737 );
buf ( n40739 , n40738 );
xor ( n40740 , n40698 , n40703 );
xor ( n40741 , n40740 , n40709 );
buf ( n40742 , n40741 );
buf ( n40743 , n40742 );
xor ( n40744 , n40523 , n40528 );
xor ( n40745 , n40744 , n40534 );
buf ( n40746 , n40745 );
buf ( n40747 , n40746 );
xor ( n40748 , n40743 , n40747 );
xor ( n40749 , n40720 , n40725 );
xor ( n40750 , n40749 , n40731 );
buf ( n40751 , n40750 );
buf ( n40752 , n40751 );
and ( n40753 , n40748 , n40752 );
and ( n40754 , n40743 , n40747 );
or ( n40755 , n40753 , n40754 );
buf ( n40756 , n40755 );
buf ( n40757 , n40756 );
xor ( n40758 , n40739 , n40757 );
xor ( n40759 , n40285 , n40290 );
and ( n40760 , n40759 , n40296 );
and ( n40761 , n40285 , n40290 );
or ( n40762 , n40760 , n40761 );
buf ( n40763 , n40762 );
buf ( n40764 , n40763 );
xor ( n40765 , n40265 , n40270 );
and ( n40766 , n40765 , n40276 );
and ( n40767 , n40265 , n40270 );
or ( n40768 , n40766 , n40767 );
buf ( n40769 , n40768 );
buf ( n40770 , n40769 );
xor ( n40771 , n40764 , n40770 );
xor ( n40772 , n40677 , n40682 );
xor ( n40773 , n40772 , n40688 );
buf ( n40774 , n40773 );
buf ( n40775 , n40774 );
and ( n40776 , n40771 , n40775 );
and ( n40777 , n40764 , n40770 );
or ( n40778 , n40776 , n40777 );
buf ( n40779 , n40778 );
buf ( n40780 , n40779 );
xor ( n40781 , n40758 , n40780 );
buf ( n40782 , n40781 );
buf ( n40783 , n40782 );
xor ( n40784 , n40260 , n40279 );
and ( n40785 , n40784 , n40299 );
and ( n40786 , n40260 , n40279 );
or ( n40787 , n40785 , n40786 );
buf ( n40788 , n40787 );
buf ( n40789 , n40788 );
xor ( n40790 , n40764 , n40770 );
xor ( n40791 , n40790 , n40775 );
buf ( n40792 , n40791 );
buf ( n40793 , n40792 );
xor ( n40794 , n40789 , n40793 );
xor ( n40795 , n40743 , n40747 );
xor ( n40796 , n40795 , n40752 );
buf ( n40797 , n40796 );
buf ( n40798 , n40797 );
and ( n40799 , n40794 , n40798 );
and ( n40800 , n40789 , n40793 );
or ( n40801 , n40799 , n40800 );
buf ( n40802 , n40801 );
buf ( n40803 , n40802 );
xor ( n40804 , n40783 , n40803 );
xor ( n40805 , n40322 , n40341 );
and ( n40806 , n40805 , n40362 );
and ( n40807 , n40322 , n40341 );
or ( n40808 , n40806 , n40807 );
buf ( n40809 , n40808 );
buf ( n40810 , n40809 );
xor ( n40811 , n40381 , n40387 );
and ( n40812 , n40811 , n40410 );
and ( n40813 , n40381 , n40387 );
or ( n40814 , n40812 , n40813 );
buf ( n40815 , n40814 );
buf ( n40816 , n40815 );
xor ( n40817 , n40810 , n40816 );
xor ( n40818 , n40653 , n40659 );
xor ( n40819 , n40818 , n40664 );
buf ( n40820 , n40819 );
buf ( n40821 , n40820 );
and ( n40822 , n40817 , n40821 );
and ( n40823 , n40810 , n40816 );
or ( n40824 , n40822 , n40823 );
buf ( n40825 , n40824 );
buf ( n40826 , n40825 );
xor ( n40827 , n40804 , n40826 );
buf ( n40828 , n40827 );
buf ( n40829 , n40828 );
xor ( n40830 , n40672 , n40829 );
xor ( n40831 , n40789 , n40793 );
xor ( n40832 , n40831 , n40798 );
buf ( n40833 , n40832 );
buf ( n40834 , n40833 );
xor ( n40835 , n40254 , n40302 );
and ( n40836 , n40835 , n40365 );
and ( n40837 , n40254 , n40302 );
or ( n40838 , n40836 , n40837 );
buf ( n40839 , n40838 );
buf ( n40840 , n40839 );
xor ( n40841 , n40834 , n40840 );
xor ( n40842 , n40375 , n40413 );
and ( n40843 , n40842 , n40420 );
and ( n40844 , n40375 , n40413 );
or ( n40845 , n40843 , n40844 );
buf ( n40846 , n40845 );
buf ( n40847 , n40846 );
and ( n40848 , n40841 , n40847 );
and ( n40849 , n40834 , n40840 );
or ( n40850 , n40848 , n40849 );
buf ( n40851 , n40850 );
buf ( n40852 , n40851 );
xor ( n40853 , n40830 , n40852 );
buf ( n40854 , n40853 );
buf ( n40855 , n40854 );
not ( n40856 , n40855 );
buf ( n40857 , n40856 );
buf ( n40858 , n40857 );
xor ( n40859 , n40810 , n40816 );
xor ( n40860 , n40859 , n40821 );
buf ( n40861 , n40860 );
buf ( n40862 , n40861 );
xor ( n40863 , n40834 , n40840 );
xor ( n40864 , n40863 , n40847 );
buf ( n40865 , n40864 );
buf ( n40866 , n40865 );
xor ( n40867 , n40862 , n40866 );
xor ( n40868 , n40248 , n40368 );
and ( n40869 , n40868 , n40423 );
and ( n40870 , n40248 , n40368 );
or ( n40871 , n40869 , n40870 );
buf ( n40872 , n40871 );
buf ( n40873 , n40872 );
and ( n40874 , n40867 , n40873 );
and ( n40875 , n40862 , n40866 );
or ( n40876 , n40874 , n40875 );
buf ( n40877 , n40876 );
buf ( n40878 , n40877 );
not ( n40879 , n40878 );
buf ( n40880 , n40879 );
buf ( n40881 , n40880 );
or ( n40882 , n40858 , n40881 );
buf ( n40883 , n40882 );
nand ( n40884 , n40857 , n40880 );
nand ( n40885 , n40883 , n40884 );
xor ( n40886 , n40862 , n40866 );
xor ( n40887 , n40886 , n40873 );
buf ( n40888 , n40887 );
buf ( n40889 , n40888 );
xor ( n40890 , n40235 , n40241 );
and ( n40891 , n40890 , n40426 );
and ( n40892 , n40235 , n40241 );
or ( n40893 , n40891 , n40892 );
buf ( n40894 , n40893 );
buf ( n40895 , n40894 );
nand ( n40896 , n40889 , n40895 );
buf ( n40897 , n40896 );
and ( n40898 , n40885 , n40897 );
nand ( n40899 , n40518 , n40898 );
or ( n40900 , n40894 , n40888 );
not ( n40901 , n40900 );
nor ( n40902 , n40901 , n40885 );
nand ( n40903 , n40517 , n40902 );
not ( n40904 , n40885 );
not ( n40905 , n40897 );
and ( n40906 , n40904 , n40905 );
not ( n40907 , n40900 );
nand ( n40908 , n40907 , n40885 , n40897 );
nand ( n40909 , n40908 , n2356 );
nor ( n40910 , n40906 , n40909 );
nand ( n40911 , n40899 , n40903 , n40910 );
nand ( n40912 , n39615 , n40911 );
not ( n40913 , n38865 );
not ( n40914 , n37966 );
or ( n40915 , n40913 , n40914 );
buf ( n40916 , n39250 );
not ( n40917 , n40916 );
buf ( n40918 , n40917 );
nand ( n40919 , n40915 , n40918 );
buf ( n40920 , n39260 );
not ( n40921 , n40920 );
buf ( n40922 , n39237 );
nand ( n40923 , n40921 , n40922 );
buf ( n40924 , n40923 );
and ( n40925 , n40924 , n454 );
and ( n40926 , n40919 , n40925 );
not ( n40927 , n40919 );
nor ( n40928 , n40924 , n2618 );
and ( n40929 , n40927 , n40928 );
nor ( n40930 , n40926 , n40929 );
buf ( n40931 , n40900 );
buf ( n40932 , n40897 );
nand ( n40933 , n40931 , n40932 );
buf ( n40934 , n40933 );
buf ( n40935 , n40934 );
not ( n40936 , n40935 );
buf ( n40937 , n40517 );
not ( n40938 , n40937 );
or ( n40939 , n40936 , n40938 );
buf ( n40940 , n40517 );
buf ( n40941 , n40934 );
or ( n40942 , n40940 , n40941 );
nand ( n40943 , n40939 , n40942 );
buf ( n40944 , n40943 );
nand ( n40945 , n2356 , n40944 );
nand ( n40946 , n40930 , n40945 );
nand ( n40947 , n36963 , n40912 , n40946 );
not ( n40948 , n40947 );
not ( n40949 , n37932 );
not ( n40950 , n40949 );
not ( n40951 , n37944 );
not ( n40952 , n40951 );
and ( n40953 , n40950 , n40952 );
and ( n40954 , n36744 , n37960 );
nor ( n40955 , n40953 , n40954 );
nand ( n40956 , n36746 , n37960 , n6922 );
nand ( n40957 , n40955 , n40956 );
nand ( n40958 , n37962 , n37954 );
not ( n40959 , n40958 );
and ( n40960 , n40957 , n40959 );
not ( n40961 , n40957 );
and ( n40962 , n40961 , n40958 );
nor ( n40963 , n40960 , n40962 );
nand ( n40964 , n40963 , n454 );
buf ( n40965 , n40489 );
buf ( n40966 , n40495 );
not ( n40967 , n40966 );
buf ( n40968 , n40477 );
nand ( n40969 , n40967 , n40968 );
buf ( n40970 , n40969 );
buf ( n40971 , n40970 );
xnor ( n40972 , n40965 , n40971 );
buf ( n40973 , n40972 );
nand ( n40974 , n40973 , n2356 );
nand ( n40975 , n40964 , n40974 );
nand ( n40976 , n40975 , n36959 );
not ( n40977 , n40976 );
buf ( n40978 , n38859 );
not ( n40979 , n40978 );
buf ( n40980 , n40979 );
not ( n40981 , n40980 );
not ( n40982 , n37966 );
or ( n40983 , n40981 , n40982 );
not ( n40984 , n38853 );
nand ( n40985 , n40984 , n38858 );
nand ( n40986 , n40983 , n40985 );
not ( n40987 , n40986 );
buf ( n40988 , n38851 );
not ( n40989 , n40988 );
buf ( n40990 , n39249 );
nand ( n40991 , n40989 , n40990 );
buf ( n40992 , n40991 );
not ( n40993 , n40992 );
and ( n40994 , n40993 , n454 );
nand ( n40995 , n40987 , n40994 );
not ( n40996 , n40993 );
nand ( n40997 , n40996 , n40986 , n454 );
not ( n40998 , n454 );
nand ( n40999 , n40512 , n40436 );
buf ( n41000 , n40999 );
not ( n41001 , n41000 );
not ( n41002 , n40228 );
not ( n41003 , n40502 );
or ( n41004 , n41002 , n41003 );
not ( n41005 , n40505 );
nand ( n41006 , n41004 , n41005 );
buf ( n41007 , n41006 );
not ( n41008 , n41007 );
or ( n41009 , n41001 , n41008 );
buf ( n41010 , n41006 );
buf ( n41011 , n40999 );
or ( n41012 , n41010 , n41011 );
nand ( n41013 , n41009 , n41012 );
buf ( n41014 , n41013 );
nand ( n41015 , n40998 , n41014 );
nand ( n41016 , n40995 , n40997 , n41015 );
nand ( n41017 , n41005 , n40228 );
xnor ( n41018 , n40502 , n41017 );
not ( n41019 , n41018 );
not ( n41020 , n2356 );
or ( n41021 , n41019 , n41020 );
not ( n41022 , n37927 );
not ( n41023 , n37955 );
or ( n41024 , n41022 , n41023 );
nand ( n41025 , n41024 , n37965 );
not ( n41026 , n41025 );
not ( n41027 , n41026 );
not ( n41028 , n41027 );
nand ( n41029 , n40985 , n40980 );
nand ( n41030 , n41028 , n41029 );
or ( n41031 , n41026 , n41029 );
nand ( n41032 , n41030 , n41031 , n454 );
nand ( n41033 , n41021 , n41032 );
buf ( n41034 , n37949 );
nand ( n41035 , n41034 , n37927 );
not ( n41036 , n41035 );
and ( n41037 , n37943 , n36732 , n37958 );
buf ( n41038 , n41037 );
buf ( n41039 , n36746 );
buf ( n41040 , n6922 );
nand ( n41041 , n41038 , n41039 , n41040 );
buf ( n41042 , n41041 );
buf ( n41043 , n37945 );
buf ( n41044 , n37954 );
and ( n41045 , n41043 , n41044 );
buf ( n41046 , n41045 );
nand ( n41047 , n41037 , n36744 );
nand ( n41048 , n41036 , n41042 , n41046 , n41047 );
not ( n41049 , n41048 );
nand ( n41050 , n41042 , n41046 , n41047 );
nand ( n41051 , n41050 , n41035 );
not ( n41052 , n41051 );
or ( n41053 , n41049 , n41052 );
nand ( n41054 , n41053 , n454 );
buf ( n41055 , n40465 );
not ( n41056 , n41055 );
buf ( n41057 , n40482 );
nand ( n41058 , n41056 , n41057 );
buf ( n41059 , n41058 );
buf ( n41060 , n41059 );
not ( n41061 , n41060 );
buf ( n41062 , n40489 );
not ( n41063 , n41062 );
buf ( n41064 , n41063 );
buf ( n41065 , n41064 );
buf ( n41066 , n40495 );
or ( n41067 , n41065 , n41066 );
buf ( n41068 , n40477 );
nand ( n41069 , n41067 , n41068 );
buf ( n41070 , n41069 );
buf ( n41071 , n41070 );
not ( n41072 , n41071 );
or ( n41073 , n41061 , n41072 );
buf ( n41074 , n41070 );
buf ( n41075 , n41059 );
or ( n41076 , n41074 , n41075 );
nand ( n41077 , n41073 , n41076 );
buf ( n41078 , n41077 );
nand ( n41079 , n2356 , n41078 );
nand ( n41080 , n41054 , n41079 );
nand ( n41081 , n40977 , n41016 , n41033 , n41080 );
not ( n41082 , n41081 );
and ( n41083 , n38862 , n39606 , n39234 );
not ( n41084 , n41083 );
not ( n41085 , n41025 );
or ( n41086 , n41084 , n41085 );
nand ( n41087 , n39258 , n39244 , n39246 );
nand ( n41088 , n41087 , n39598 );
not ( n41089 , n41088 );
not ( n41090 , n41089 );
nand ( n41091 , n41086 , n41090 );
xor ( n41092 , n39500 , n39506 );
and ( n41093 , n41092 , n39513 );
and ( n41094 , n39500 , n39506 );
or ( n41095 , n41093 , n41094 );
buf ( n41096 , n41095 );
buf ( n41097 , n41096 );
xor ( n41098 , n39524 , n39541 );
and ( n41099 , n41098 , n39562 );
and ( n41100 , n39524 , n39541 );
or ( n41101 , n41099 , n41100 );
buf ( n41102 , n41101 );
buf ( n41103 , n41102 );
buf ( n41104 , n39463 );
not ( n41105 , n41104 );
buf ( n41106 , n33967 );
not ( n41107 , n41106 );
or ( n41108 , n41105 , n41107 );
xnor ( n41109 , n491 , n509 );
buf ( n41110 , n41109 );
not ( n41111 , n41110 );
buf ( n41112 , n33973 );
nand ( n41113 , n41111 , n41112 );
buf ( n41114 , n41113 );
buf ( n41115 , n41114 );
nand ( n41116 , n41108 , n41115 );
buf ( n41117 , n41116 );
buf ( n41118 , n41117 );
buf ( n41119 , n1698 );
buf ( n41120 , n30769 );
or ( n41121 , n41119 , n41120 );
buf ( n41122 , n497 );
nand ( n41123 , n41121 , n41122 );
buf ( n41124 , n41123 );
buf ( n41125 , n41124 );
xor ( n41126 , n41118 , n41125 );
buf ( n41127 , n39552 );
not ( n41128 , n41127 );
buf ( n41129 , n33757 );
not ( n41130 , n41129 );
or ( n41131 , n41128 , n41130 );
buf ( n41132 , n495 );
buf ( n41133 , n505 );
xnor ( n41134 , n41132 , n41133 );
buf ( n41135 , n41134 );
buf ( n41136 , n41135 );
not ( n41137 , n41136 );
buf ( n41138 , n33167 );
nand ( n41139 , n41137 , n41138 );
buf ( n41140 , n41139 );
buf ( n41141 , n41140 );
nand ( n41142 , n41131 , n41141 );
buf ( n41143 , n41142 );
buf ( n41144 , n41143 );
xor ( n41145 , n41126 , n41144 );
buf ( n41146 , n41145 );
buf ( n41147 , n41146 );
xor ( n41148 , n41103 , n41147 );
buf ( n41149 , n39558 );
buf ( n41150 , n39469 );
not ( n41151 , n41150 );
buf ( n41152 , n39481 );
not ( n41153 , n41152 );
or ( n41154 , n41151 , n41153 );
buf ( n41155 , n39481 );
buf ( n41156 , n39469 );
or ( n41157 , n41155 , n41156 );
buf ( n41158 , n39498 );
nand ( n41159 , n41157 , n41158 );
buf ( n41160 , n41159 );
buf ( n41161 , n41160 );
nand ( n41162 , n41154 , n41161 );
buf ( n41163 , n41162 );
buf ( n41164 , n41163 );
xor ( n41165 , n41149 , n41164 );
and ( n41166 , n38927 , n38928 );
buf ( n41167 , n41166 );
buf ( n41168 , n41167 );
buf ( n41169 , n39533 );
not ( n41170 , n41169 );
buf ( n41171 , n4241 );
not ( n41172 , n41171 );
or ( n41173 , n41170 , n41172 );
buf ( n41174 , n4218 );
buf ( n41175 , n507 );
buf ( n41176 , n493 );
xor ( n41177 , n41175 , n41176 );
buf ( n41178 , n41177 );
buf ( n41179 , n41178 );
nand ( n41180 , n41174 , n41179 );
buf ( n41181 , n41180 );
buf ( n41182 , n41181 );
nand ( n41183 , n41173 , n41182 );
buf ( n41184 , n41183 );
buf ( n41185 , n41184 );
xor ( n41186 , n41168 , n41185 );
buf ( n41187 , n39492 );
not ( n41188 , n41187 );
buf ( n41189 , n36290 );
not ( n41190 , n41189 );
or ( n41191 , n41188 , n41190 );
buf ( n41192 , n37254 );
buf ( n41193 , n489 );
buf ( n41194 , n511 );
xor ( n41195 , n41193 , n41194 );
buf ( n41196 , n41195 );
buf ( n41197 , n41196 );
nand ( n41198 , n41192 , n41197 );
buf ( n41199 , n41198 );
buf ( n41200 , n41199 );
nand ( n41201 , n41191 , n41200 );
buf ( n41202 , n41201 );
buf ( n41203 , n41202 );
xor ( n41204 , n41186 , n41203 );
buf ( n41205 , n41204 );
buf ( n41206 , n41205 );
xor ( n41207 , n41165 , n41206 );
buf ( n41208 , n41207 );
buf ( n41209 , n41208 );
xor ( n41210 , n41148 , n41209 );
buf ( n41211 , n41210 );
buf ( n41212 , n41211 );
xor ( n41213 , n41097 , n41212 );
xor ( n41214 , n39565 , n39570 );
and ( n41215 , n41214 , n39577 );
and ( n41216 , n39565 , n39570 );
or ( n41217 , n41215 , n41216 );
buf ( n41218 , n41217 );
buf ( n41219 , n41218 );
xor ( n41220 , n41213 , n41219 );
buf ( n41221 , n41220 );
xor ( n41222 , n39515 , n39520 );
and ( n41223 , n41222 , n39579 );
and ( n41224 , n39515 , n39520 );
or ( n41225 , n41223 , n41224 );
nand ( n41226 , n41221 , n41225 );
not ( n41227 , n41221 );
not ( n41228 , n41225 );
nand ( n41229 , n41227 , n41228 );
and ( n41230 , n41226 , n41229 );
and ( n41231 , n38359 , n39587 , n39017 );
not ( n41232 , n41231 );
not ( n41233 , n38188 );
or ( n41234 , n41232 , n41233 );
not ( n41235 , n39587 );
not ( n41236 , n39451 );
or ( n41237 , n41235 , n41236 );
nand ( n41238 , n41237 , n39588 );
not ( n41239 , n41238 );
nand ( n41240 , n41234 , n41239 );
xor ( n41241 , n41230 , n41240 );
nand ( n41242 , n41241 , n29519 );
nand ( n41243 , n39430 , n38806 );
nor ( n41244 , n41243 , n39425 );
not ( n41245 , n41244 );
not ( n41246 , n38609 );
or ( n41247 , n41245 , n41246 );
not ( n41248 , n39426 );
not ( n41249 , n39440 );
or ( n41250 , n41248 , n41249 );
nand ( n41251 , n41250 , n39428 );
not ( n41252 , n41251 );
nand ( n41253 , n41247 , n41252 );
xor ( n41254 , n39273 , n39279 );
and ( n41255 , n41254 , n39335 );
and ( n41256 , n39273 , n39279 );
or ( n41257 , n41255 , n41256 );
buf ( n41258 , n41257 );
buf ( n41259 , n41258 );
xor ( n41260 , n39348 , n39369 );
and ( n41261 , n41260 , n39396 );
and ( n41262 , n39348 , n39369 );
or ( n41263 , n41261 , n41262 );
buf ( n41264 , n41263 );
buf ( n41265 , n41264 );
buf ( n41266 , n33014 );
not ( n41267 , n41266 );
buf ( n41268 , n30585 );
not ( n41269 , n41268 );
buf ( n41270 , n41269 );
buf ( n41271 , n41270 );
not ( n41272 , n41271 );
or ( n41273 , n41267 , n41272 );
buf ( n41274 , n497 );
nand ( n41275 , n41273 , n41274 );
buf ( n41276 , n41275 );
buf ( n41277 , n41276 );
buf ( n41278 , n34465 );
not ( n41279 , n41278 );
buf ( n41280 , n39295 );
not ( n41281 , n41280 );
or ( n41282 , n41279 , n41281 );
buf ( n41283 , n491 );
not ( n41284 , n41283 );
buf ( n41285 , n31829 );
not ( n41286 , n41285 );
or ( n41287 , n41284 , n41286 );
buf ( n41288 , n31826 );
buf ( n41289 , n3524 );
nand ( n41290 , n41288 , n41289 );
buf ( n41291 , n41290 );
buf ( n41292 , n41291 );
nand ( n41293 , n41287 , n41292 );
buf ( n41294 , n41293 );
buf ( n41295 , n41294 );
buf ( n41296 , n3045 );
nand ( n41297 , n41295 , n41296 );
buf ( n41298 , n41297 );
buf ( n41299 , n41298 );
nand ( n41300 , n41282 , n41299 );
buf ( n41301 , n41300 );
buf ( n41302 , n41301 );
xor ( n41303 , n41277 , n41302 );
buf ( n41304 , n31812 );
not ( n41305 , n41304 );
buf ( n41306 , n39358 );
not ( n41307 , n41306 );
or ( n41308 , n41305 , n41307 );
buf ( n41309 , n495 );
not ( n41310 , n41309 );
buf ( n41311 , n5561 );
buf ( n41312 , n41311 );
buf ( n41313 , n41312 );
not ( n41314 , n41313 );
or ( n41315 , n41310 , n41314 );
not ( n41316 , n41311 );
buf ( n41317 , n41316 );
buf ( n41318 , n31784 );
nand ( n41319 , n41317 , n41318 );
buf ( n41320 , n41319 );
buf ( n41321 , n41320 );
nand ( n41322 , n41315 , n41321 );
buf ( n41323 , n41322 );
buf ( n41324 , n41323 );
buf ( n41325 , n2725 );
nand ( n41326 , n41324 , n41325 );
buf ( n41327 , n41326 );
buf ( n41328 , n41327 );
nand ( n41329 , n41308 , n41328 );
buf ( n41330 , n41329 );
buf ( n41331 , n41330 );
xor ( n41332 , n41303 , n41331 );
buf ( n41333 , n41332 );
buf ( n41334 , n41333 );
xor ( n41335 , n41265 , n41334 );
buf ( n41336 , n39365 );
buf ( n41337 , n3948 );
not ( n41338 , n41337 );
buf ( n41339 , n39134 );
not ( n41340 , n41339 );
or ( n41341 , n41338 , n41340 );
buf ( n41342 , n39299 );
nand ( n41343 , n41341 , n41342 );
buf ( n41344 , n41343 );
buf ( n41345 , n41344 );
buf ( n41346 , n39313 );
or ( n41347 , n41345 , n41346 );
buf ( n41348 , n39333 );
nand ( n41349 , n41347 , n41348 );
buf ( n41350 , n41349 );
buf ( n41351 , n41350 );
buf ( n41352 , n41344 );
buf ( n41353 , n39313 );
nand ( n41354 , n41352 , n41353 );
buf ( n41355 , n41354 );
buf ( n41356 , n41355 );
nand ( n41357 , n41351 , n41356 );
buf ( n41358 , n41357 );
buf ( n41359 , n41358 );
xor ( n41360 , n41336 , n41359 );
and ( n41361 , n39155 , n39156 );
buf ( n41362 , n41361 );
buf ( n41363 , n41362 );
not ( n41364 , n2978 );
buf ( n41365 , n38414 );
buf ( n41366 , n2704 );
nand ( n41367 , n41365 , n41366 );
buf ( n41368 , n41367 );
nand ( n41369 , n38410 , n493 );
nand ( n41370 , n41368 , n41369 );
not ( n41371 , n41370 );
or ( n41372 , n41364 , n41371 );
buf ( n41373 , n39388 );
buf ( n41374 , n3146 );
nand ( n41375 , n41373 , n41374 );
buf ( n41376 , n41375 );
nand ( n41377 , n41372 , n41376 );
buf ( n41378 , n41377 );
xor ( n41379 , n41363 , n41378 );
buf ( n41380 , n36508 );
not ( n41381 , n41380 );
and ( n41382 , n489 , n38391 );
not ( n41383 , n489 );
and ( n41384 , n41383 , n2671 );
nor ( n41385 , n41382 , n41384 );
buf ( n41386 , n41385 );
not ( n41387 , n41386 );
or ( n41388 , n41381 , n41387 );
buf ( n41389 , n39326 );
buf ( n41390 , n37542 );
nand ( n41391 , n41389 , n41390 );
buf ( n41392 , n41391 );
buf ( n41393 , n41392 );
nand ( n41394 , n41388 , n41393 );
buf ( n41395 , n41394 );
buf ( n41396 , n41395 );
xor ( n41397 , n41379 , n41396 );
buf ( n41398 , n41397 );
buf ( n41399 , n41398 );
xor ( n41400 , n41360 , n41399 );
buf ( n41401 , n41400 );
buf ( n41402 , n41401 );
xor ( n41403 , n41335 , n41402 );
buf ( n41404 , n41403 );
buf ( n41405 , n41404 );
xor ( n41406 , n41259 , n41405 );
xor ( n41407 , n39399 , n39405 );
and ( n41408 , n41407 , n39412 );
and ( n41409 , n39399 , n39405 );
or ( n41410 , n41408 , n41409 );
buf ( n41411 , n41410 );
buf ( n41412 , n41411 );
xor ( n41413 , n41406 , n41412 );
buf ( n41414 , n41413 );
not ( n41415 , n41414 );
xor ( n41416 , n39338 , n39344 );
and ( n41417 , n41416 , n39415 );
and ( n41418 , n39338 , n39344 );
or ( n41419 , n41417 , n41418 );
buf ( n41420 , n41419 );
not ( n41421 , n41420 );
nand ( n41422 , n41415 , n41421 );
not ( n41423 , n41422 );
not ( n41424 , n41423 );
not ( n41425 , n41421 );
buf ( n41426 , n41414 );
nand ( n41427 , n41425 , n41426 );
nand ( n41428 , n41424 , n41427 );
not ( n41429 , n41428 );
and ( n41430 , n41253 , n41429 );
not ( n41431 , n41253 );
and ( n41432 , n41431 , n41428 );
nor ( n41433 , n41430 , n41432 );
nand ( n41434 , n41433 , n455 );
nand ( n41435 , n41242 , n41434 );
nand ( n41436 , n41435 , n39597 );
not ( n41437 , n41436 );
not ( n41438 , n29519 );
not ( n41439 , n41241 );
or ( n41440 , n41438 , n41439 );
nand ( n41441 , n41433 , n455 );
nand ( n41442 , n41440 , n41441 );
nor ( n41443 , n39597 , n41442 );
buf ( n41444 , n41443 );
or ( n41445 , n41437 , n41444 );
xnor ( n41446 , n41091 , n41445 );
not ( n41447 , n41446 );
not ( n41448 , n454 );
or ( n41449 , n41447 , n41448 );
xor ( n41450 , n40672 , n40829 );
and ( n41451 , n41450 , n40852 );
and ( n41452 , n40672 , n40829 );
or ( n41453 , n41451 , n41452 );
buf ( n41454 , n41453 );
buf ( n41455 , n41454 );
xor ( n41456 , n40581 , n40646 );
and ( n41457 , n41456 , n40669 );
and ( n41458 , n40581 , n40646 );
or ( n41459 , n41457 , n41458 );
buf ( n41460 , n41459 );
buf ( n41461 , n41460 );
xor ( n41462 , n40693 , n40714 );
and ( n41463 , n41462 , n40736 );
and ( n41464 , n40693 , n40714 );
or ( n41465 , n41463 , n41464 );
buf ( n41466 , n41465 );
buf ( n41467 , n41466 );
buf ( n41468 , n526 );
buf ( n41469 , n542 );
and ( n41470 , n41468 , n41469 );
buf ( n41471 , n41470 );
buf ( n41472 , n41471 );
buf ( n41473 , n527 );
buf ( n41474 , n541 );
and ( n41475 , n41473 , n41474 );
buf ( n41476 , n41475 );
buf ( n41477 , n41476 );
xor ( n41478 , n41472 , n41477 );
xor ( n41479 , n40564 , n40569 );
and ( n41480 , n41479 , n40575 );
and ( n41481 , n40564 , n40569 );
or ( n41482 , n41480 , n41481 );
buf ( n41483 , n41482 );
buf ( n41484 , n41483 );
xor ( n41485 , n41478 , n41484 );
buf ( n41486 , n41485 );
buf ( n41487 , n41486 );
xor ( n41488 , n41467 , n41487 );
xor ( n41489 , n40586 , n40591 );
and ( n41490 , n41489 , n40597 );
and ( n41491 , n40586 , n40591 );
or ( n41492 , n41490 , n41491 );
buf ( n41493 , n41492 );
buf ( n41494 , n41493 );
xor ( n41495 , n40605 , n40610 );
and ( n41496 , n41495 , n40616 );
and ( n41497 , n40605 , n40610 );
or ( n41498 , n41496 , n41497 );
buf ( n41499 , n41498 );
buf ( n41500 , n41499 );
xor ( n41501 , n41494 , n41500 );
xor ( n41502 , n40544 , n40549 );
and ( n41503 , n41502 , n40555 );
and ( n41504 , n40544 , n40549 );
or ( n41505 , n41503 , n41504 );
buf ( n41506 , n41505 );
buf ( n41507 , n41506 );
xor ( n41508 , n41501 , n41507 );
buf ( n41509 , n41508 );
buf ( n41510 , n41509 );
xor ( n41511 , n41488 , n41510 );
buf ( n41512 , n41511 );
buf ( n41513 , n41512 );
xor ( n41514 , n40739 , n40757 );
and ( n41515 , n41514 , n40780 );
and ( n41516 , n40739 , n40757 );
or ( n41517 , n41515 , n41516 );
buf ( n41518 , n41517 );
buf ( n41519 , n41518 );
xor ( n41520 , n41513 , n41519 );
xor ( n41521 , n40539 , n40558 );
and ( n41522 , n41521 , n40578 );
and ( n41523 , n40539 , n40558 );
or ( n41524 , n41522 , n41523 );
buf ( n41525 , n41524 );
buf ( n41526 , n41525 );
buf ( n41527 , n528 );
buf ( n41528 , n540 );
and ( n41529 , n41527 , n41528 );
buf ( n41530 , n41529 );
buf ( n41531 , n41530 );
buf ( n41532 , n529 );
buf ( n41533 , n539 );
and ( n41534 , n41532 , n41533 );
buf ( n41535 , n41534 );
buf ( n41536 , n41535 );
xor ( n41537 , n41531 , n41536 );
buf ( n41538 , n525 );
buf ( n41539 , n543 );
and ( n41540 , n41538 , n41539 );
buf ( n41541 , n41540 );
buf ( n41542 , n41541 );
xor ( n41543 , n41537 , n41542 );
buf ( n41544 , n41543 );
buf ( n41545 , n41544 );
buf ( n41546 , n530 );
buf ( n41547 , n538 );
and ( n41548 , n41546 , n41547 );
buf ( n41549 , n41548 );
buf ( n41550 , n41549 );
buf ( n41551 , n531 );
buf ( n41552 , n537 );
and ( n41553 , n41551 , n41552 );
buf ( n41554 , n41553 );
buf ( n41555 , n41554 );
xor ( n41556 , n41550 , n41555 );
buf ( n41557 , n523 );
buf ( n41558 , n545 );
and ( n41559 , n41557 , n41558 );
buf ( n41560 , n41559 );
buf ( n41561 , n41560 );
xor ( n41562 , n41556 , n41561 );
buf ( n41563 , n41562 );
buf ( n41564 , n41563 );
xor ( n41565 , n41545 , n41564 );
buf ( n41566 , n521 );
buf ( n41567 , n547 );
and ( n41568 , n41566 , n41567 );
buf ( n41569 , n41568 );
buf ( n41570 , n41569 );
buf ( n41571 , n522 );
buf ( n41572 , n546 );
and ( n41573 , n41571 , n41572 );
buf ( n41574 , n41573 );
buf ( n41575 , n41574 );
xor ( n41576 , n41570 , n41575 );
buf ( n41577 , n524 );
buf ( n41578 , n544 );
and ( n41579 , n41577 , n41578 );
buf ( n41580 , n41579 );
buf ( n41581 , n41580 );
xor ( n41582 , n41576 , n41581 );
buf ( n41583 , n41582 );
buf ( n41584 , n41583 );
xor ( n41585 , n41565 , n41584 );
buf ( n41586 , n41585 );
buf ( n41587 , n41586 );
xor ( n41588 , n41526 , n41587 );
xor ( n41589 , n40600 , n40619 );
and ( n41590 , n41589 , n40643 );
and ( n41591 , n40600 , n40619 );
or ( n41592 , n41590 , n41591 );
buf ( n41593 , n41592 );
buf ( n41594 , n41593 );
xor ( n41595 , n41588 , n41594 );
buf ( n41596 , n41595 );
buf ( n41597 , n41596 );
xor ( n41598 , n41520 , n41597 );
buf ( n41599 , n41598 );
buf ( n41600 , n41599 );
xor ( n41601 , n41461 , n41600 );
xor ( n41602 , n40783 , n40803 );
and ( n41603 , n41602 , n40826 );
and ( n41604 , n40783 , n40803 );
or ( n41605 , n41603 , n41604 );
buf ( n41606 , n41605 );
buf ( n41607 , n41606 );
xor ( n41608 , n41601 , n41607 );
buf ( n41609 , n41608 );
buf ( n41610 , n41609 );
or ( n41611 , n41455 , n41610 );
buf ( n41612 , n41611 );
buf ( n41613 , n41612 );
buf ( n41614 , n41609 );
buf ( n41615 , n41454 );
nand ( n41616 , n41614 , n41615 );
buf ( n41617 , n41616 );
buf ( n41618 , n41617 );
nand ( n41619 , n41613 , n41618 );
buf ( n41620 , n41619 );
buf ( n41621 , n41620 );
not ( n41622 , n41621 );
not ( n41623 , n40501 );
not ( n41624 , n40437 );
nand ( n41625 , n41624 , n40884 , n40228 , n40900 );
not ( n41626 , n41625 );
and ( n41627 , n41623 , n41626 );
buf ( n41628 , n40900 );
not ( n41629 , n41628 );
buf ( n41630 , n40513 );
not ( n41631 , n41630 );
or ( n41632 , n41629 , n41631 );
buf ( n41633 , n40897 );
nand ( n41634 , n41632 , n41633 );
buf ( n41635 , n41634 );
nand ( n41636 , n41635 , n40884 );
nand ( n41637 , n40438 , n40884 , n40483 , n40900 );
nand ( n41638 , n41636 , n41637 , n40883 );
nor ( n41639 , n41627 , n41638 );
not ( n41640 , n41639 );
buf ( n41641 , n41640 );
buf ( n41642 , n41641 );
not ( n41643 , n41642 );
or ( n41644 , n41622 , n41643 );
buf ( n41645 , n41641 );
buf ( n41646 , n41620 );
or ( n41647 , n41645 , n41646 );
nand ( n41648 , n41644 , n41647 );
buf ( n41649 , n41648 );
nand ( n41650 , n41649 , n2356 );
buf ( n41651 , n41650 );
nand ( n41652 , n41449 , n41651 );
nand ( n41653 , n40948 , n41082 , n41652 );
not ( n41654 , n41653 );
not ( n41655 , n454 );
buf ( n41656 , n37966 );
not ( n41657 , n41656 );
nand ( n41658 , n39606 , n38862 , n39234 );
nor ( n41659 , n41437 , n41658 );
buf ( n41660 , n41659 );
not ( n41661 , n41660 );
or ( n41662 , n41657 , n41661 );
and ( n41663 , n41087 , n39598 , n41436 );
nor ( n41664 , n41444 , n41663 );
buf ( n41665 , n41664 );
nand ( n41666 , n41662 , n41665 );
buf ( n41667 , n41666 );
not ( n41668 , n29519 );
not ( n41669 , n41229 );
nor ( n41670 , n38173 , n41669 );
nand ( n41671 , n41670 , n7433 , n41231 );
not ( n41672 , n37417 );
not ( n41673 , n37437 );
or ( n41674 , n41672 , n41673 );
nand ( n41675 , n41674 , n38846 );
not ( n41676 , n41228 );
not ( n41677 , n41221 );
not ( n41678 , n41677 );
or ( n41679 , n41676 , n41678 );
nand ( n41680 , n41679 , n39587 );
nor ( n41681 , n38178 , n41680 );
nand ( n41682 , n41675 , n41681 , n39445 );
not ( n41683 , n41682 );
not ( n41684 , n39450 );
and ( n41685 , n39018 , n39588 );
not ( n41686 , n41685 );
or ( n41687 , n41684 , n41686 );
not ( n41688 , n41680 );
nand ( n41689 , n41687 , n41688 );
nand ( n41690 , n41689 , n41226 );
nor ( n41691 , n41683 , n41690 );
nand ( n41692 , n41671 , n41691 );
xor ( n41693 , n41097 , n41212 );
and ( n41694 , n41693 , n41219 );
and ( n41695 , n41097 , n41212 );
or ( n41696 , n41694 , n41695 );
buf ( n41697 , n41696 );
xor ( n41698 , n41149 , n41164 );
and ( n41699 , n41698 , n41206 );
and ( n41700 , n41149 , n41164 );
or ( n41701 , n41699 , n41700 );
buf ( n41702 , n41701 );
buf ( n41703 , n41702 );
and ( n41704 , n39489 , n39490 );
buf ( n41705 , n41704 );
buf ( n41706 , n41705 );
buf ( n41707 , n489 );
buf ( n41708 , n510 );
xor ( n41709 , n41707 , n41708 );
buf ( n41710 , n41709 );
buf ( n41711 , n41710 );
not ( n41712 , n41711 );
buf ( n41713 , n37254 );
not ( n41714 , n41713 );
or ( n41715 , n41712 , n41714 );
buf ( n41716 , n5172 );
buf ( n41717 , n41716 );
buf ( n41718 , n41717 );
buf ( n41719 , n41718 );
buf ( n41720 , n41196 );
nand ( n41721 , n41719 , n41720 );
buf ( n41722 , n41721 );
buf ( n41723 , n41722 );
nand ( n41724 , n41715 , n41723 );
buf ( n41725 , n41724 );
buf ( n41726 , n41725 );
xor ( n41727 , n41706 , n41726 );
buf ( n41728 , n495 );
not ( n41729 , n41728 );
buf ( n41730 , n33167 );
not ( n41731 , n41730 );
or ( n41732 , n41729 , n41731 );
buf ( n41733 , n33757 );
not ( n41734 , n41733 );
buf ( n41735 , n41734 );
buf ( n41736 , n41735 );
buf ( n41737 , n41135 );
or ( n41738 , n41736 , n41737 );
nand ( n41739 , n41732 , n41738 );
buf ( n41740 , n41739 );
buf ( n41741 , n41740 );
xor ( n41742 , n41727 , n41741 );
buf ( n41743 , n41742 );
buf ( n41744 , n41743 );
xor ( n41745 , n41118 , n41125 );
and ( n41746 , n41745 , n41144 );
and ( n41747 , n41118 , n41125 );
or ( n41748 , n41746 , n41747 );
buf ( n41749 , n41748 );
buf ( n41750 , n41749 );
xor ( n41751 , n41744 , n41750 );
buf ( n41752 , n33964 );
buf ( n41753 , n41109 );
or ( n41754 , n41752 , n41753 );
buf ( n41755 , n33973 );
not ( n41756 , n41755 );
buf ( n41757 , n41756 );
buf ( n41758 , n41757 );
buf ( n41759 , n508 );
buf ( n41760 , n491 );
xor ( n41761 , n41759 , n41760 );
buf ( n41762 , n41761 );
buf ( n41763 , n41762 );
not ( n41764 , n41763 );
buf ( n41765 , n41764 );
buf ( n41766 , n41765 );
or ( n41767 , n41758 , n41766 );
nand ( n41768 , n41754 , n41767 );
buf ( n41769 , n41768 );
buf ( n41770 , n41769 );
buf ( n41771 , n41178 );
not ( n41772 , n41771 );
buf ( n41773 , n4241 );
not ( n41774 , n41773 );
or ( n41775 , n41772 , n41774 );
not ( n41776 , n4218 );
buf ( n41777 , n41776 );
buf ( n41778 , n506 );
buf ( n41779 , n493 );
xnor ( n41780 , n41778 , n41779 );
buf ( n41781 , n41780 );
buf ( n41782 , n41781 );
or ( n41783 , n41777 , n41782 );
buf ( n41784 , n41783 );
buf ( n41785 , n41784 );
nand ( n41786 , n41775 , n41785 );
buf ( n41787 , n41786 );
buf ( n41788 , n41787 );
not ( n41789 , n41788 );
buf ( n41790 , n41789 );
buf ( n41791 , n41790 );
xor ( n41792 , n41770 , n41791 );
xor ( n41793 , n41168 , n41185 );
and ( n41794 , n41793 , n41203 );
and ( n41795 , n41168 , n41185 );
or ( n41796 , n41794 , n41795 );
buf ( n41797 , n41796 );
buf ( n41798 , n41797 );
xor ( n41799 , n41792 , n41798 );
buf ( n41800 , n41799 );
buf ( n41801 , n41800 );
xor ( n41802 , n41751 , n41801 );
buf ( n41803 , n41802 );
buf ( n41804 , n41803 );
xor ( n41805 , n41703 , n41804 );
xor ( n41806 , n41103 , n41147 );
and ( n41807 , n41806 , n41209 );
and ( n41808 , n41103 , n41147 );
or ( n41809 , n41807 , n41808 );
buf ( n41810 , n41809 );
buf ( n41811 , n41810 );
xor ( n41812 , n41805 , n41811 );
buf ( n41813 , n41812 );
nor ( n41814 , n41697 , n41813 );
not ( n41815 , n41814 );
nand ( n41816 , n41813 , n41697 );
nand ( n41817 , n41815 , n41816 );
xnor ( n41818 , n41692 , n41817 );
not ( n41819 , n41818 );
or ( n41820 , n41668 , n41819 );
xor ( n41821 , n41336 , n41359 );
and ( n41822 , n41821 , n41399 );
and ( n41823 , n41336 , n41359 );
or ( n41824 , n41822 , n41823 );
buf ( n41825 , n41824 );
buf ( n41826 , n41825 );
and ( n41827 , n39320 , n39324 );
buf ( n41828 , n41827 );
buf ( n41829 , n41828 );
buf ( n41830 , n31812 );
not ( n41831 , n41830 );
buf ( n41832 , n41323 );
not ( n41833 , n41832 );
or ( n41834 , n41831 , n41833 );
buf ( n41835 , n2725 );
buf ( n41836 , n495 );
nand ( n41837 , n41835 , n41836 );
buf ( n41838 , n41837 );
buf ( n41839 , n41838 );
nand ( n41840 , n41834 , n41839 );
buf ( n41841 , n41840 );
buf ( n41842 , n41841 );
xor ( n41843 , n41829 , n41842 );
buf ( n41844 , n39149 );
not ( n41845 , n41844 );
buf ( n41846 , n41385 );
not ( n41847 , n41846 );
or ( n41848 , n41845 , n41847 );
buf ( n41849 , n489 );
buf ( n41850 , n2803 );
xor ( n41851 , n41849 , n41850 );
buf ( n41852 , n41851 );
buf ( n41853 , n41852 );
buf ( n41854 , n36508 );
nand ( n41855 , n41853 , n41854 );
buf ( n41856 , n41855 );
buf ( n41857 , n41856 );
nand ( n41858 , n41848 , n41857 );
buf ( n41859 , n41858 );
buf ( n41860 , n41859 );
xor ( n41861 , n41843 , n41860 );
buf ( n41862 , n41861 );
buf ( n41863 , n41862 );
xor ( n41864 , n41277 , n41302 );
and ( n41865 , n41864 , n41331 );
and ( n41866 , n41277 , n41302 );
or ( n41867 , n41865 , n41866 );
buf ( n41868 , n41867 );
buf ( n41869 , n41868 );
xor ( n41870 , n41863 , n41869 );
buf ( n41871 , n34465 );
not ( n41872 , n41871 );
buf ( n41873 , n41294 );
not ( n41874 , n41873 );
or ( n41875 , n41872 , n41874 );
buf ( n41876 , n491 );
not ( n41877 , n41876 );
buf ( n41878 , n3211 );
not ( n41879 , n41878 );
or ( n41880 , n41877 , n41879 );
buf ( n41881 , n39383 );
buf ( n41882 , n3524 );
nand ( n41883 , n41881 , n41882 );
buf ( n41884 , n41883 );
buf ( n41885 , n41884 );
nand ( n41886 , n41880 , n41885 );
buf ( n41887 , n41886 );
buf ( n41888 , n41887 );
buf ( n41889 , n3045 );
nand ( n41890 , n41888 , n41889 );
buf ( n41891 , n41890 );
buf ( n41892 , n41891 );
nand ( n41893 , n41875 , n41892 );
buf ( n41894 , n41893 );
buf ( n41895 , n41894 );
buf ( n41896 , n3146 );
not ( n41897 , n41896 );
buf ( n41898 , n41370 );
not ( n41899 , n41898 );
or ( n41900 , n41897 , n41899 );
buf ( n41901 , n2704 );
not ( n41902 , n37462 );
buf ( n41903 , n41902 );
and ( n41904 , n41901 , n41903 );
not ( n41905 , n41901 );
buf ( n41906 , n37462 );
and ( n41907 , n41905 , n41906 );
nor ( n41908 , n41904 , n41907 );
buf ( n41909 , n41908 );
buf ( n41910 , n41909 );
buf ( n41911 , n3113 );
nand ( n41912 , n41910 , n41911 );
buf ( n41913 , n41912 );
buf ( n41914 , n41913 );
nand ( n41915 , n41900 , n41914 );
buf ( n41916 , n41915 );
buf ( n41917 , n41916 );
not ( n41918 , n41917 );
buf ( n41919 , n41918 );
buf ( n41920 , n41919 );
xor ( n41921 , n41895 , n41920 );
xor ( n41922 , n41363 , n41378 );
and ( n41923 , n41922 , n41396 );
and ( n41924 , n41363 , n41378 );
or ( n41925 , n41923 , n41924 );
buf ( n41926 , n41925 );
buf ( n41927 , n41926 );
xor ( n41928 , n41921 , n41927 );
buf ( n41929 , n41928 );
buf ( n41930 , n41929 );
xor ( n41931 , n41870 , n41930 );
buf ( n41932 , n41931 );
buf ( n41933 , n41932 );
xor ( n41934 , n41826 , n41933 );
xor ( n41935 , n41265 , n41334 );
and ( n41936 , n41935 , n41402 );
and ( n41937 , n41265 , n41334 );
or ( n41938 , n41936 , n41937 );
buf ( n41939 , n41938 );
buf ( n41940 , n41939 );
xor ( n41941 , n41934 , n41940 );
buf ( n41942 , n41941 );
xor ( n41943 , n41259 , n41405 );
and ( n41944 , n41943 , n41412 );
and ( n41945 , n41259 , n41405 );
or ( n41946 , n41944 , n41945 );
buf ( n41947 , n41946 );
nand ( n41948 , n41942 , n41947 );
not ( n41949 , n41948 );
nor ( n41950 , n41942 , n41947 );
nor ( n41951 , n41949 , n41950 );
not ( n41952 , n37846 );
not ( n41953 , n37863 );
or ( n41954 , n41952 , n41953 );
not ( n41955 , n38842 );
nand ( n41956 , n41954 , n41955 );
not ( n41957 , n39430 );
nor ( n41958 , n41957 , n39432 );
nand ( n41959 , n41422 , n39424 );
nor ( n41960 , n38598 , n41959 );
nand ( n41961 , n41956 , n41958 , n41960 );
not ( n41962 , n41961 );
and ( n41963 , n39224 , n39427 );
not ( n41964 , n41963 );
not ( n41965 , n39438 );
or ( n41966 , n41964 , n41965 );
not ( n41967 , n41959 );
nand ( n41968 , n41966 , n41967 );
nand ( n41969 , n41968 , n41427 );
nor ( n41970 , n41962 , n41969 );
nor ( n41971 , n38594 , n41423 );
nand ( n41972 , n41971 , n41244 , n38368 );
nand ( n41973 , n41970 , n41972 );
xor ( n41974 , n41951 , n41973 );
nand ( n41975 , n41974 , n455 );
nand ( n41976 , n41820 , n41975 );
not ( n41977 , n29519 );
not ( n41978 , n41241 );
or ( n41979 , n41977 , n41978 );
nand ( n41980 , n41979 , n41434 );
buf ( n41981 , n41980 );
not ( n41982 , n41981 );
buf ( n41983 , n41982 );
nand ( n41984 , n41976 , n41983 );
not ( n41985 , n41976 );
buf ( n41986 , n41442 );
nand ( n41987 , n41985 , n41986 );
nand ( n41988 , n41984 , n41987 );
buf ( n41989 , n41988 );
not ( n41990 , n41989 );
buf ( n41991 , n41990 );
and ( n41992 , n41667 , n41991 );
not ( n41993 , n41667 );
and ( n41994 , n41993 , n41988 );
nor ( n41995 , n41992 , n41994 );
not ( n41996 , n41995 );
or ( n41997 , n41655 , n41996 );
xor ( n41998 , n41526 , n41587 );
and ( n41999 , n41998 , n41594 );
and ( n42000 , n41526 , n41587 );
or ( n42001 , n41999 , n42000 );
buf ( n42002 , n42001 );
buf ( n42003 , n42002 );
buf ( n42004 , n530 );
buf ( n42005 , n537 );
and ( n42006 , n42004 , n42005 );
buf ( n42007 , n42006 );
buf ( n42008 , n42007 );
buf ( n42009 , n523 );
buf ( n42010 , n544 );
and ( n42011 , n42009 , n42010 );
buf ( n42012 , n42011 );
buf ( n42013 , n42012 );
xor ( n42014 , n42008 , n42013 );
buf ( n42015 , n526 );
buf ( n42016 , n541 );
and ( n42017 , n42015 , n42016 );
buf ( n42018 , n42017 );
buf ( n42019 , n42018 );
xor ( n42020 , n42014 , n42019 );
buf ( n42021 , n42020 );
buf ( n42022 , n42021 );
xor ( n42023 , n41494 , n41500 );
and ( n42024 , n42023 , n41507 );
and ( n42025 , n41494 , n41500 );
or ( n42026 , n42024 , n42025 );
buf ( n42027 , n42026 );
buf ( n42028 , n42027 );
xor ( n42029 , n42022 , n42028 );
xor ( n42030 , n41472 , n41477 );
and ( n42031 , n42030 , n41484 );
and ( n42032 , n41472 , n41477 );
or ( n42033 , n42031 , n42032 );
buf ( n42034 , n42033 );
buf ( n42035 , n42034 );
xor ( n42036 , n42029 , n42035 );
buf ( n42037 , n42036 );
buf ( n42038 , n42037 );
xor ( n42039 , n41467 , n41487 );
and ( n42040 , n42039 , n41510 );
and ( n42041 , n41467 , n41487 );
or ( n42042 , n42040 , n42041 );
buf ( n42043 , n42042 );
buf ( n42044 , n42043 );
xor ( n42045 , n42038 , n42044 );
buf ( n42046 , n527 );
buf ( n42047 , n540 );
and ( n42048 , n42046 , n42047 );
buf ( n42049 , n42048 );
buf ( n42050 , n42049 );
xor ( n42051 , n41570 , n41575 );
and ( n42052 , n42051 , n41581 );
and ( n42053 , n41570 , n41575 );
or ( n42054 , n42052 , n42053 );
buf ( n42055 , n42054 );
buf ( n42056 , n42055 );
xor ( n42057 , n42050 , n42056 );
xor ( n42058 , n41531 , n41536 );
and ( n42059 , n42058 , n41542 );
and ( n42060 , n41531 , n41536 );
or ( n42061 , n42059 , n42060 );
buf ( n42062 , n42061 );
buf ( n42063 , n42062 );
xor ( n42064 , n42057 , n42063 );
buf ( n42065 , n42064 );
buf ( n42066 , n42065 );
xor ( n42067 , n41545 , n41564 );
and ( n42068 , n42067 , n41584 );
and ( n42069 , n41545 , n41564 );
or ( n42070 , n42068 , n42069 );
buf ( n42071 , n42070 );
buf ( n42072 , n42071 );
xor ( n42073 , n42066 , n42072 );
xor ( n42074 , n41550 , n41555 );
and ( n42075 , n42074 , n41561 );
and ( n42076 , n41550 , n41555 );
or ( n42077 , n42075 , n42076 );
buf ( n42078 , n42077 );
buf ( n42079 , n42078 );
buf ( n42080 , n521 );
buf ( n42081 , n546 );
and ( n42082 , n42080 , n42081 );
buf ( n42083 , n42082 );
buf ( n42084 , n42083 );
buf ( n42085 , n522 );
buf ( n42086 , n545 );
and ( n42087 , n42085 , n42086 );
buf ( n42088 , n42087 );
buf ( n42089 , n42088 );
xor ( n42090 , n42084 , n42089 );
buf ( n42091 , n524 );
buf ( n42092 , n543 );
and ( n42093 , n42091 , n42092 );
buf ( n42094 , n42093 );
buf ( n42095 , n42094 );
xor ( n42096 , n42090 , n42095 );
buf ( n42097 , n42096 );
buf ( n42098 , n42097 );
xor ( n42099 , n42079 , n42098 );
buf ( n42100 , n528 );
buf ( n42101 , n539 );
and ( n42102 , n42100 , n42101 );
buf ( n42103 , n42102 );
buf ( n42104 , n42103 );
buf ( n42105 , n529 );
buf ( n42106 , n538 );
and ( n42107 , n42105 , n42106 );
buf ( n42108 , n42107 );
buf ( n42109 , n42108 );
xor ( n42110 , n42104 , n42109 );
buf ( n42111 , n525 );
buf ( n42112 , n542 );
and ( n42113 , n42111 , n42112 );
buf ( n42114 , n42113 );
buf ( n42115 , n42114 );
xor ( n42116 , n42110 , n42115 );
buf ( n42117 , n42116 );
buf ( n42118 , n42117 );
xor ( n42119 , n42099 , n42118 );
buf ( n42120 , n42119 );
buf ( n42121 , n42120 );
xor ( n42122 , n42073 , n42121 );
buf ( n42123 , n42122 );
buf ( n42124 , n42123 );
xor ( n42125 , n42045 , n42124 );
buf ( n42126 , n42125 );
buf ( n42127 , n42126 );
xor ( n42128 , n42003 , n42127 );
xor ( n42129 , n41513 , n41519 );
and ( n42130 , n42129 , n41597 );
and ( n42131 , n41513 , n41519 );
or ( n42132 , n42130 , n42131 );
buf ( n42133 , n42132 );
buf ( n42134 , n42133 );
xor ( n42135 , n42128 , n42134 );
buf ( n42136 , n42135 );
xor ( n42137 , n41461 , n41600 );
and ( n42138 , n42137 , n41607 );
and ( n42139 , n41461 , n41600 );
or ( n42140 , n42138 , n42139 );
buf ( n42141 , n42140 );
nor ( n42142 , n42136 , n42141 );
buf ( n42143 , n42142 );
not ( n42144 , n42143 );
buf ( n42145 , n42141 );
buf ( n42146 , n42136 );
nand ( n42147 , n42145 , n42146 );
buf ( n42148 , n42147 );
buf ( n42149 , n42148 );
nand ( n42150 , n42144 , n42149 );
buf ( n42151 , n42150 );
buf ( n42152 , n42151 );
not ( n42153 , n42152 );
buf ( n42154 , n41612 );
not ( n42155 , n42154 );
buf ( n42156 , n41640 );
not ( n42157 , n42156 );
or ( n42158 , n42155 , n42157 );
buf ( n42159 , n41617 );
nand ( n42160 , n42158 , n42159 );
buf ( n42161 , n42160 );
buf ( n42162 , n42161 );
not ( n42163 , n42162 );
or ( n42164 , n42153 , n42163 );
buf ( n42165 , n42161 );
buf ( n42166 , n42151 );
or ( n42167 , n42165 , n42166 );
nand ( n42168 , n42164 , n42167 );
buf ( n42169 , n42168 );
nand ( n42170 , n42169 , n2356 );
nand ( n42171 , n41997 , n42170 );
xor ( n42172 , n41654 , n42171 );
not ( n42173 , n42172 );
or ( n42174 , n37045 , n42173 );
not ( n42175 , n7162 );
and ( n42176 , n7157 , n7081 );
and ( n42177 , n7065 , n497 );
nor ( n42178 , n42176 , n42177 );
or ( n42179 , n42175 , n42178 );
and ( n42180 , n7066 , n36988 );
and ( n42181 , n7065 , n496 );
nor ( n42182 , n42180 , n42181 );
not ( n42183 , n7108 );
or ( n42184 , n42182 , n42183 );
nand ( n42185 , n42179 , n42184 );
not ( n42186 , n29494 );
not ( n42187 , n42186 );
and ( n42188 , n42187 , n1970 );
not ( n42189 , n29494 );
and ( n42190 , n42189 , n499 );
nor ( n42191 , n42188 , n42190 );
not ( n42192 , n42191 );
not ( n42193 , n42192 );
buf ( n42194 , n2803 );
not ( n42195 , n42194 );
nand ( n42196 , n42195 , n29494 );
not ( n42197 , n29494 );
nand ( n42198 , n42197 , n42194 );
nand ( n42199 , n42196 , n42198 );
nand ( n42200 , n36982 , n42199 );
not ( n42201 , n42200 );
not ( n42202 , n42201 );
or ( n42203 , n42193 , n42202 );
not ( n42204 , n42189 );
and ( n42205 , n42204 , n7092 );
not ( n42206 , n29494 );
and ( n42207 , n42206 , n498 );
nor ( n42208 , n42205 , n42207 );
not ( n42209 , n42208 );
not ( n42210 , n36982 );
nand ( n42211 , n42209 , n42210 );
nand ( n42212 , n42203 , n42211 );
xor ( n42213 , n42185 , n42212 );
not ( n42214 , n495 );
and ( n42215 , n35943 , n42214 );
not ( n42216 , n35943 );
and ( n42217 , n42216 , n495 );
nor ( n42218 , n42215 , n42217 );
or ( n42219 , n7214 , n42218 );
buf ( n42220 , n7226 );
not ( n42221 , n494 );
and ( n42222 , n35943 , n42221 );
and ( n42223 , n42216 , n494 );
nor ( n42224 , n42222 , n42223 );
or ( n42225 , n42220 , n42224 );
nand ( n42226 , n42219 , n42225 );
and ( n42227 , n42213 , n42226 );
and ( n42228 , n42185 , n42212 );
or ( n42229 , n42227 , n42228 );
not ( n42230 , n42201 );
not ( n42231 , n42208 );
not ( n42232 , n42231 );
or ( n42233 , n42230 , n42232 );
and ( n42234 , n42187 , n7081 );
and ( n42235 , n42189 , n497 );
nor ( n42236 , n42234 , n42235 );
not ( n42237 , n42236 );
nand ( n42238 , n42237 , n42210 );
nand ( n42239 , n42233 , n42238 );
or ( n42240 , n7214 , n42224 );
not ( n42241 , n493 );
not ( n42242 , n35943 );
or ( n42243 , n42241 , n42242 );
or ( n42244 , n7102 , n493 );
nand ( n42245 , n42243 , n42244 );
or ( n42246 , n7226 , n42245 );
nand ( n42247 , n42240 , n42246 );
xor ( n42248 , n42239 , n42247 );
buf ( n42249 , n3220 );
and ( n42250 , n42249 , n29494 );
not ( n42251 , n42249 );
and ( n42252 , n42251 , n42186 );
or ( n42253 , n42250 , n42252 );
and ( n42254 , n42249 , n38414 );
not ( n42255 , n42249 );
buf ( n42256 , n3434 );
not ( n42257 , n42256 );
and ( n42258 , n42255 , n42257 );
nor ( n42259 , n42254 , n42258 );
nand ( n42260 , n42253 , n42259 );
buf ( n42261 , n42256 );
and ( n42262 , n42261 , n7140 );
not ( n42263 , n42261 );
and ( n42264 , n42263 , n500 );
nor ( n42265 , n42262 , n42264 );
or ( n42266 , n42260 , n42265 );
and ( n42267 , n42261 , n1970 );
not ( n42268 , n42261 );
and ( n42269 , n42268 , n499 );
nor ( n42270 , n42267 , n42269 );
buf ( n42271 , n42253 );
or ( n42272 , n42270 , n42271 );
nand ( n42273 , n42266 , n42272 );
xor ( n42274 , n42248 , n42273 );
xor ( n42275 , n42229 , n42274 );
not ( n42276 , n492 );
and ( n42277 , n7123 , n42276 );
and ( n42278 , n7178 , n492 );
nor ( n42279 , n42277 , n42278 );
or ( n42280 , n7299 , n42279 );
not ( n42281 , n7139 );
not ( n42282 , n491 );
and ( n42283 , n7123 , n42282 );
and ( n42284 , n7178 , n491 );
nor ( n42285 , n42283 , n42284 );
or ( n42286 , n42281 , n42285 );
nand ( n42287 , n42280 , n42286 );
nor ( n42288 , n41312 , n7165 );
xor ( n42289 , n42287 , n42288 );
not ( n42290 , n42175 );
not ( n42291 , n42290 );
or ( n42292 , n42291 , n42182 );
not ( n42293 , n7108 );
not ( n42294 , n7065 );
and ( n42295 , n42214 , n42294 );
not ( n42296 , n42214 );
and ( n42297 , n42296 , n7065 );
nor ( n42298 , n42295 , n42297 );
or ( n42299 , n42293 , n42298 );
nand ( n42300 , n42292 , n42299 );
xor ( n42301 , n42289 , n42300 );
xor ( n42302 , n42275 , n42301 );
xor ( n42303 , n42185 , n42212 );
xor ( n42304 , n42303 , n42226 );
not ( n42305 , n42260 );
not ( n42306 , n42305 );
and ( n42307 , n42261 , n7122 );
and ( n42308 , n42263 , n501 );
nor ( n42309 , n42307 , n42308 );
or ( n42310 , n42306 , n42309 );
or ( n42311 , n42265 , n42271 );
nand ( n42312 , n42310 , n42311 );
xor ( n42313 , n41902 , n42256 );
xnor ( n42314 , n41902 , n41316 );
nand ( n42315 , n42313 , n42314 );
not ( n42316 , n41312 );
and ( n42317 , n42316 , n7165 );
and ( n42318 , n41312 , n503 );
nor ( n42319 , n42317 , n42318 );
or ( n42320 , n42315 , n42319 );
buf ( n42321 , n42313 );
and ( n42322 , n42316 , n7204 );
and ( n42323 , n41312 , n502 );
nor ( n42324 , n42322 , n42323 );
or ( n42325 , n42321 , n42324 );
nand ( n42326 , n42320 , n42325 );
xor ( n42327 , n42312 , n42326 );
not ( n42328 , n41902 );
and ( n42329 , n42261 , n42328 );
and ( n42330 , n42263 , n41902 );
nor ( n42331 , n42330 , n7151 );
nor ( n42332 , n42329 , n42331 , n41312 );
not ( n42333 , n7071 );
and ( n42334 , n7074 , n42282 );
and ( n42335 , n7087 , n491 );
nor ( n42336 , n42334 , n42335 );
not ( n42337 , n42336 );
not ( n42338 , n42337 );
or ( n42339 , n42333 , n42338 );
and ( n42340 , n7074 , n42276 );
and ( n42341 , n7087 , n492 );
nor ( n42342 , n42340 , n42341 );
or ( n42343 , n42342 , n7098 );
nand ( n42344 , n42339 , n42343 );
and ( n42345 , n42332 , n42344 );
xor ( n42346 , n42327 , n42345 );
xor ( n42347 , n42304 , n42346 );
xor ( n42348 , n42332 , n42344 );
nor ( n42349 , n42321 , n7151 );
and ( n42350 , n7123 , n42214 );
and ( n42351 , n7178 , n495 );
nor ( n42352 , n42350 , n42351 );
or ( n42353 , n7299 , n42352 );
and ( n42354 , n7123 , n42221 );
and ( n42355 , n7178 , n494 );
nor ( n42356 , n42354 , n42355 );
or ( n42357 , n42281 , n42356 );
nand ( n42358 , n42353 , n42357 );
xor ( n42359 , n42349 , n42358 );
and ( n42360 , n7066 , n1970 );
and ( n42361 , n7065 , n499 );
nor ( n42362 , n42360 , n42361 );
or ( n42363 , n42291 , n42362 );
and ( n42364 , n7066 , n7092 );
and ( n42365 , n7065 , n498 );
nor ( n42366 , n42364 , n42365 );
or ( n42367 , n42366 , n42293 );
nand ( n42368 , n42363 , n42367 );
and ( n42369 , n42359 , n42368 );
and ( n42370 , n42349 , n42358 );
or ( n42371 , n42369 , n42370 );
xor ( n42372 , n42348 , n42371 );
and ( n42373 , n42187 , n7122 );
and ( n42374 , n42189 , n501 );
nor ( n42375 , n42373 , n42374 );
or ( n42376 , n42200 , n42375 );
and ( n42377 , n42187 , n7140 );
and ( n42378 , n42206 , n500 );
nor ( n42379 , n42377 , n42378 );
or ( n42380 , n42379 , n36982 );
nand ( n42381 , n42376 , n42380 );
not ( n42382 , n493 );
and ( n42383 , n7074 , n42382 );
and ( n42384 , n7087 , n493 );
nor ( n42385 , n42383 , n42384 );
or ( n42386 , n42385 , n7098 );
or ( n42387 , n42342 , n7314 );
nand ( n42388 , n42386 , n42387 );
xor ( n42389 , n42381 , n42388 );
and ( n42390 , n42261 , n7165 );
and ( n42391 , n42263 , n503 );
nor ( n42392 , n42390 , n42391 );
or ( n42393 , n42392 , n42260 );
and ( n42394 , n42261 , n7204 );
and ( n42395 , n42263 , n502 );
nor ( n42396 , n42394 , n42395 );
or ( n42397 , n42396 , n42271 );
nand ( n42398 , n42393 , n42397 );
and ( n42399 , n42389 , n42398 );
and ( n42400 , n42381 , n42388 );
or ( n42401 , n42399 , n42400 );
and ( n42402 , n42372 , n42401 );
and ( n42403 , n42348 , n42371 );
or ( n42404 , n42402 , n42403 );
and ( n42405 , n42347 , n42404 );
and ( n42406 , n42304 , n42346 );
or ( n42407 , n42405 , n42406 );
xor ( n42408 , n42302 , n42407 );
xor ( n42409 , n42312 , n42326 );
and ( n42410 , n42409 , n42345 );
and ( n42411 , n42312 , n42326 );
or ( n42412 , n42410 , n42411 );
or ( n42413 , n42315 , n42324 );
and ( n42414 , n42316 , n7122 );
and ( n42415 , n41312 , n501 );
nor ( n42416 , n42414 , n42415 );
or ( n42417 , n42416 , n42321 );
nand ( n42418 , n42413 , n42417 );
not ( n42419 , n490 );
and ( n42420 , n7074 , n42419 );
and ( n42421 , n7087 , n490 );
nor ( n42422 , n42420 , n42421 );
or ( n42423 , n42422 , n7098 );
and ( n42424 , n7074 , n5539 );
and ( n42425 , n7087 , n489 );
nor ( n42426 , n42424 , n42425 );
or ( n42427 , n42426 , n7314 );
nand ( n42428 , n42423 , n42427 );
xor ( n42429 , n42418 , n42428 );
nor ( n42430 , n41312 , n7151 );
or ( n42431 , n42336 , n7098 );
or ( n42432 , n42422 , n7314 );
nand ( n42433 , n42431 , n42432 );
xor ( n42434 , n42430 , n42433 );
and ( n42435 , n7350 , n42382 );
and ( n42436 , n7178 , n493 );
nor ( n42437 , n42435 , n42436 );
or ( n42438 , n7299 , n42437 );
or ( n42439 , n42281 , n42279 );
nand ( n42440 , n42438 , n42439 );
and ( n42441 , n42434 , n42440 );
and ( n42442 , n42430 , n42433 );
or ( n42443 , n42441 , n42442 );
xor ( n42444 , n42429 , n42443 );
xor ( n42445 , n42412 , n42444 );
or ( n42446 , n7299 , n42356 );
or ( n42447 , n42281 , n42437 );
nand ( n42448 , n42446 , n42447 );
or ( n42449 , n42291 , n42366 );
or ( n42450 , n42178 , n42293 );
nand ( n42451 , n42449 , n42450 );
xor ( n42452 , n42448 , n42451 );
not ( n42453 , n42198 );
not ( n42454 , n42196 );
or ( n42455 , n42453 , n42454 );
buf ( n42456 , n36982 );
nand ( n42457 , n42455 , n42456 );
or ( n42458 , n42457 , n42379 );
or ( n42459 , n42191 , n42456 );
nand ( n42460 , n42458 , n42459 );
and ( n42461 , n42452 , n42460 );
and ( n42462 , n42448 , n42451 );
or ( n42463 , n42461 , n42462 );
and ( n42464 , n35943 , n36988 );
and ( n42465 , n42216 , n496 );
nor ( n42466 , n42464 , n42465 );
or ( n42467 , n7214 , n42466 );
or ( n42468 , n42218 , n42220 );
nand ( n42469 , n42467 , n42468 );
or ( n42470 , n42260 , n42396 );
or ( n42471 , n42309 , n42271 );
nand ( n42472 , n42470 , n42471 );
xor ( n42473 , n42469 , n42472 );
and ( n42474 , n42316 , n7151 );
and ( n42475 , n41312 , n504 );
nor ( n42476 , n42474 , n42475 );
or ( n42477 , n42315 , n42476 );
or ( n42478 , n42321 , n42319 );
nand ( n42479 , n42477 , n42478 );
and ( n42480 , n42473 , n42479 );
and ( n42481 , n42469 , n42472 );
or ( n42482 , n42480 , n42481 );
xor ( n42483 , n42463 , n42482 );
xor ( n42484 , n42430 , n42433 );
xor ( n42485 , n42484 , n42440 );
and ( n42486 , n42483 , n42485 );
and ( n42487 , n42463 , n42482 );
or ( n42488 , n42486 , n42487 );
xor ( n42489 , n42445 , n42488 );
xor ( n42490 , n42408 , n42489 );
xor ( n42491 , n42463 , n42482 );
xor ( n42492 , n42491 , n42485 );
xor ( n42493 , n42304 , n42346 );
xor ( n42494 , n42493 , n42404 );
xor ( n42495 , n42492 , n42494 );
xor ( n42496 , n42469 , n42472 );
xor ( n42497 , n42496 , n42479 );
xor ( n42498 , n42448 , n42451 );
xor ( n42499 , n42498 , n42460 );
xor ( n42500 , n42497 , n42499 );
and ( n42501 , n35943 , n7081 );
and ( n42502 , n42216 , n497 );
nor ( n42503 , n42501 , n42502 );
or ( n42504 , n7214 , n42503 );
or ( n42505 , n42220 , n42466 );
nand ( n42506 , n42504 , n42505 );
or ( n42507 , n42187 , n42249 );
nand ( n42508 , n42507 , n504 );
nand ( n42509 , n42204 , n42249 );
and ( n42510 , n42508 , n42509 , n42261 );
xnor ( n42511 , n36988 , n7178 );
or ( n42512 , n7299 , n42511 );
or ( n42513 , n42281 , n42352 );
nand ( n42514 , n42512 , n42513 );
and ( n42515 , n42510 , n42514 );
xor ( n42516 , n42506 , n42515 );
and ( n42517 , n7066 , n7140 );
and ( n42518 , n7065 , n500 );
nor ( n42519 , n42517 , n42518 );
or ( n42520 , n42519 , n42175 );
or ( n42521 , n42362 , n42183 );
nand ( n42522 , n42520 , n42521 );
and ( n42523 , n42187 , n7204 );
and ( n42524 , n42186 , n502 );
nor ( n42525 , n42523 , n42524 );
not ( n42526 , n42525 );
not ( n42527 , n42526 );
not ( n42528 , n42201 );
or ( n42529 , n42527 , n42528 );
not ( n42530 , n42375 );
nand ( n42531 , n42530 , n42210 );
nand ( n42532 , n42529 , n42531 );
xor ( n42533 , n42522 , n42532 );
and ( n42534 , n494 , n35952 );
not ( n42535 , n494 );
and ( n42536 , n42535 , n7091 );
nor ( n42537 , n42534 , n42536 );
or ( n42538 , n42537 , n7098 );
or ( n42539 , n42385 , n7314 );
nand ( n42540 , n42538 , n42539 );
and ( n42541 , n42533 , n42540 );
and ( n42542 , n42522 , n42532 );
or ( n42543 , n42541 , n42542 );
and ( n42544 , n42516 , n42543 );
and ( n42545 , n42506 , n42515 );
or ( n42546 , n42544 , n42545 );
and ( n42547 , n42500 , n42546 );
and ( n42548 , n42497 , n42499 );
or ( n42549 , n42547 , n42548 );
and ( n42550 , n42495 , n42549 );
and ( n42551 , n42492 , n42494 );
or ( n42552 , n42550 , n42551 );
nand ( n42553 , n42490 , n42552 );
not ( n42554 , n42553 );
xor ( n42555 , n42492 , n42494 );
xor ( n42556 , n42555 , n42549 );
not ( n42557 , n42556 );
xor ( n42558 , n42348 , n42371 );
xor ( n42559 , n42558 , n42401 );
xor ( n42560 , n42381 , n42388 );
xor ( n42561 , n42560 , n42398 );
xor ( n42562 , n42349 , n42358 );
xor ( n42563 , n42562 , n42368 );
xor ( n42564 , n42561 , n42563 );
and ( n42565 , n42261 , n7151 );
and ( n42566 , n42263 , n504 );
nor ( n42567 , n42565 , n42566 );
or ( n42568 , n42306 , n42567 );
or ( n42569 , n42392 , n42271 );
nand ( n42570 , n42568 , n42569 );
and ( n42571 , n35943 , n7092 );
and ( n42572 , n7103 , n498 );
nor ( n42573 , n42571 , n42572 );
or ( n42574 , n7214 , n42573 );
or ( n42575 , n42503 , n42220 );
nand ( n42576 , n42574 , n42575 );
xor ( n42577 , n42570 , n42576 );
xor ( n42578 , n42510 , n42514 );
and ( n42579 , n42577 , n42578 );
and ( n42580 , n42570 , n42576 );
or ( n42581 , n42579 , n42580 );
and ( n42582 , n42564 , n42581 );
and ( n42583 , n42561 , n42563 );
or ( n42584 , n42582 , n42583 );
xor ( n42585 , n42559 , n42584 );
xor ( n42586 , n42497 , n42499 );
xor ( n42587 , n42586 , n42546 );
and ( n42588 , n42585 , n42587 );
and ( n42589 , n42559 , n42584 );
or ( n42590 , n42588 , n42589 );
not ( n42591 , n42590 );
nor ( n42592 , n42557 , n42591 );
nor ( n42593 , n42554 , n42592 );
not ( n42594 , n42490 );
not ( n42595 , n42552 );
nand ( n42596 , n42594 , n42595 );
not ( n42597 , n42596 );
or ( n42598 , n42593 , n42597 );
nand ( n42599 , n42557 , n42591 );
xor ( n42600 , n42506 , n42515 );
xor ( n42601 , n42600 , n42543 );
nor ( n42602 , n42253 , n7151 );
and ( n42603 , n497 , n7124 );
not ( n42604 , n497 );
and ( n42605 , n42604 , n7350 );
nor ( n42606 , n42603 , n42605 );
not ( n42607 , n42606 );
not ( n42608 , n42607 );
not ( n42609 , n7136 );
or ( n42610 , n42608 , n42609 );
not ( n42611 , n42511 );
nand ( n42612 , n42611 , n7139 );
nand ( n42613 , n42610 , n42612 );
xor ( n42614 , n42602 , n42613 );
and ( n42615 , n7066 , n7122 );
and ( n42616 , n7065 , n501 );
nor ( n42617 , n42615 , n42616 );
or ( n42618 , n42175 , n42617 );
or ( n42619 , n42519 , n42293 );
nand ( n42620 , n42618 , n42619 );
and ( n42621 , n42614 , n42620 );
and ( n42622 , n42602 , n42613 );
or ( n42623 , n42621 , n42622 );
not ( n42624 , n42210 );
not ( n42625 , n42526 );
or ( n42626 , n42624 , n42625 );
and ( n42627 , n503 , n42186 );
not ( n42628 , n503 );
and ( n42629 , n42628 , n29494 );
nor ( n42630 , n42627 , n42629 );
or ( n42631 , n42630 , n42200 );
nand ( n42632 , n42626 , n42631 );
and ( n42633 , n495 , n7090 );
not ( n42634 , n495 );
and ( n42635 , n42634 , n7074 );
nor ( n42636 , n42633 , n42635 );
or ( n42637 , n42636 , n7098 );
or ( n42638 , n42537 , n7314 );
nand ( n42639 , n42637 , n42638 );
xor ( n42640 , n42632 , n42639 );
and ( n42641 , n35943 , n1970 );
and ( n42642 , n7103 , n499 );
nor ( n42643 , n42641 , n42642 );
or ( n42644 , n7214 , n42643 );
or ( n42645 , n42573 , n7226 );
nand ( n42646 , n42644 , n42645 );
and ( n42647 , n42640 , n42646 );
and ( n42648 , n42632 , n42639 );
or ( n42649 , n42647 , n42648 );
xor ( n42650 , n42623 , n42649 );
xor ( n42651 , n42522 , n42532 );
xor ( n42652 , n42651 , n42540 );
and ( n42653 , n42650 , n42652 );
and ( n42654 , n42623 , n42649 );
or ( n42655 , n42653 , n42654 );
xor ( n42656 , n42601 , n42655 );
xor ( n42657 , n42561 , n42563 );
xor ( n42658 , n42657 , n42581 );
and ( n42659 , n42656 , n42658 );
and ( n42660 , n42601 , n42655 );
or ( n42661 , n42659 , n42660 );
xor ( n42662 , n42559 , n42584 );
xor ( n42663 , n42662 , n42587 );
xor ( n42664 , n42661 , n42663 );
xor ( n42665 , n42570 , n42576 );
xor ( n42666 , n42665 , n42578 );
xor ( n42667 , n42623 , n42649 );
xor ( n42668 , n42667 , n42652 );
xor ( n42669 , n42666 , n42668 );
or ( n42670 , n42294 , n42194 );
nand ( n42671 , n42670 , n504 );
nand ( n42672 , n7066 , n42194 );
and ( n42673 , n42671 , n42672 , n42187 );
not ( n42674 , n37011 );
not ( n42675 , n7136 );
or ( n42676 , n42674 , n42675 );
or ( n42677 , n42281 , n42606 );
nand ( n42678 , n42676 , n42677 );
and ( n42679 , n42673 , n42678 );
not ( n42680 , n36999 );
not ( n42681 , n7162 );
or ( n42682 , n42680 , n42681 );
not ( n42683 , n42617 );
nand ( n42684 , n42683 , n7108 );
nand ( n42685 , n42682 , n42684 );
and ( n42686 , n42187 , n7151 );
and ( n42687 , n42206 , n504 );
nor ( n42688 , n42686 , n42687 );
or ( n42689 , n42688 , n42200 );
or ( n42690 , n42630 , n36982 );
nand ( n42691 , n42689 , n42690 );
xor ( n42692 , n42685 , n42691 );
not ( n42693 , n7071 );
not ( n42694 , n42636 );
not ( n42695 , n42694 );
or ( n42696 , n42693 , n42695 );
not ( n42697 , n36990 );
or ( n42698 , n42697 , n7098 );
nand ( n42699 , n42696 , n42698 );
and ( n42700 , n42692 , n42699 );
and ( n42701 , n42685 , n42691 );
or ( n42702 , n42700 , n42701 );
xor ( n42703 , n42679 , n42702 );
xor ( n42704 , n42602 , n42613 );
xor ( n42705 , n42704 , n42620 );
and ( n42706 , n42703 , n42705 );
and ( n42707 , n42679 , n42702 );
or ( n42708 , n42706 , n42707 );
and ( n42709 , n42669 , n42708 );
and ( n42710 , n42666 , n42668 );
or ( n42711 , n42709 , n42710 );
xor ( n42712 , n42601 , n42655 );
xor ( n42713 , n42712 , n42658 );
xor ( n42714 , n42711 , n42713 );
xor ( n42715 , n42632 , n42639 );
xor ( n42716 , n42715 , n42646 );
or ( n42717 , n7214 , n37020 );
or ( n42718 , n42643 , n7226 );
nand ( n42719 , n42717 , n42718 );
xor ( n42720 , n42673 , n42678 );
xor ( n42721 , n42719 , n42720 );
xor ( n42722 , n36983 , n36994 );
and ( n42723 , n42722 , n37005 );
and ( n42724 , n36983 , n36994 );
or ( n42725 , n42723 , n42724 );
and ( n42726 , n42721 , n42725 );
and ( n42727 , n42719 , n42720 );
or ( n42728 , n42726 , n42727 );
xor ( n42729 , n42716 , n42728 );
xor ( n42730 , n42679 , n42702 );
xor ( n42731 , n42730 , n42705 );
and ( n42732 , n42729 , n42731 );
and ( n42733 , n42716 , n42728 );
or ( n42734 , n42732 , n42733 );
xor ( n42735 , n42666 , n42668 );
xor ( n42736 , n42735 , n42708 );
xor ( n42737 , n42734 , n42736 );
xor ( n42738 , n42685 , n42691 );
xor ( n42739 , n42738 , n42699 );
xor ( n42740 , n37016 , n37022 );
and ( n42741 , n42740 , n37024 );
and ( n42742 , n37016 , n37022 );
or ( n42743 , n42741 , n42742 );
xor ( n42744 , n42739 , n42743 );
xor ( n42745 , n42719 , n42720 );
xor ( n42746 , n42745 , n42725 );
and ( n42747 , n42744 , n42746 );
and ( n42748 , n42739 , n42743 );
or ( n42749 , n42747 , n42748 );
xor ( n42750 , n42716 , n42728 );
xor ( n42751 , n42750 , n42731 );
xor ( n42752 , n42749 , n42751 );
xor ( n42753 , n36976 , n37006 );
and ( n42754 , n42753 , n37025 );
and ( n42755 , n36976 , n37006 );
or ( n42756 , n42754 , n42755 );
xor ( n42757 , n42739 , n42743 );
xor ( n42758 , n42757 , n42746 );
xor ( n42759 , n42756 , n42758 );
not ( n42760 , n37031 );
not ( n42761 , n7254 );
not ( n42762 , n36259 );
or ( n42763 , n42761 , n42762 );
nand ( n42764 , n42763 , n7255 );
not ( n42765 , n42764 );
or ( n42766 , n42760 , n42765 );
nand ( n42767 , n42766 , n37032 );
and ( n42768 , n42759 , n42767 );
and ( n42769 , n42756 , n42758 );
or ( n42770 , n42768 , n42769 );
and ( n42771 , n42752 , n42770 );
and ( n42772 , n42749 , n42751 );
or ( n42773 , n42771 , n42772 );
and ( n42774 , n42737 , n42773 );
and ( n42775 , n42734 , n42736 );
or ( n42776 , n42774 , n42775 );
and ( n42777 , n42714 , n42776 );
and ( n42778 , n42711 , n42713 );
or ( n42779 , n42777 , n42778 );
and ( n42780 , n42664 , n42779 );
and ( n42781 , n42661 , n42663 );
or ( n42782 , n42780 , n42781 );
nand ( n42783 , n42599 , n42782 , n42596 );
nand ( n42784 , n42598 , n42783 );
buf ( n42785 , n42784 );
xor ( n42786 , n42239 , n42247 );
and ( n42787 , n42786 , n42273 );
and ( n42788 , n42239 , n42247 );
or ( n42789 , n42787 , n42788 );
or ( n42790 , n7214 , n42245 );
and ( n42791 , n35943 , n42276 );
and ( n42792 , n42216 , n492 );
nor ( n42793 , n42791 , n42792 );
or ( n42794 , n7226 , n42793 );
nand ( n42795 , n42790 , n42794 );
or ( n42796 , n42260 , n42270 );
and ( n42797 , n42261 , n7092 );
and ( n42798 , n42257 , n498 );
nor ( n42799 , n42797 , n42798 );
or ( n42800 , n42799 , n42253 );
nand ( n42801 , n42796 , n42800 );
xor ( n42802 , n42795 , n42801 );
or ( n42803 , n42315 , n42416 );
and ( n42804 , n42316 , n7140 );
and ( n42805 , n41312 , n500 );
nor ( n42806 , n42804 , n42805 );
or ( n42807 , n42806 , n42321 );
nand ( n42808 , n42803 , n42807 );
xor ( n42809 , n42802 , n42808 );
xor ( n42810 , n42789 , n42809 );
or ( n42811 , n42175 , n42298 );
and ( n42812 , n494 , n7065 );
not ( n42813 , n494 );
and ( n42814 , n42813 , n7066 );
nor ( n42815 , n42812 , n42814 );
or ( n42816 , n42183 , n42815 );
nand ( n42817 , n42811 , n42816 );
nor ( n42818 , n41312 , n7204 );
xor ( n42819 , n42817 , n42818 );
or ( n42820 , n42236 , n42200 );
and ( n42821 , n42187 , n36988 );
and ( n42822 , n42206 , n496 );
nor ( n42823 , n42821 , n42822 );
or ( n42824 , n42823 , n36982 );
nand ( n42825 , n42820 , n42824 );
xor ( n42826 , n42819 , n42825 );
xor ( n42827 , n42810 , n42826 );
or ( n42828 , n42426 , n7098 );
or ( n42829 , n7087 , n7314 );
nand ( n42830 , n42828 , n42829 );
or ( n42831 , n7299 , n42285 );
and ( n42832 , n7350 , n42419 );
and ( n42833 , n7124 , n490 );
nor ( n42834 , n42832 , n42833 );
or ( n42835 , n42281 , n42834 );
nand ( n42836 , n42831 , n42835 );
xor ( n42837 , n42830 , n42836 );
xor ( n42838 , n42287 , n42288 );
and ( n42839 , n42838 , n42300 );
and ( n42840 , n42287 , n42288 );
or ( n42841 , n42839 , n42840 );
xor ( n42842 , n42837 , n42841 );
xor ( n42843 , n42418 , n42428 );
and ( n42844 , n42843 , n42443 );
and ( n42845 , n42418 , n42428 );
or ( n42846 , n42844 , n42845 );
xor ( n42847 , n42842 , n42846 );
xor ( n42848 , n42229 , n42274 );
and ( n42849 , n42848 , n42301 );
and ( n42850 , n42229 , n42274 );
or ( n42851 , n42849 , n42850 );
xor ( n42852 , n42847 , n42851 );
xor ( n42853 , n42827 , n42852 );
xor ( n42854 , n42412 , n42444 );
and ( n42855 , n42854 , n42488 );
and ( n42856 , n42412 , n42444 );
or ( n42857 , n42855 , n42856 );
xor ( n42858 , n42853 , n42857 );
xor ( n42859 , n42302 , n42407 );
and ( n42860 , n42859 , n42489 );
and ( n42861 , n42302 , n42407 );
or ( n42862 , n42860 , n42861 );
or ( n42863 , n42858 , n42862 );
not ( n42864 , n42863 );
and ( n42865 , n42785 , n42864 );
nand ( n42866 , n42858 , n42862 );
not ( n42867 , n42866 );
and ( n42868 , n42785 , n42867 );
nor ( n42869 , n42865 , n42868 );
not ( n42870 , n42862 );
not ( n42871 , n42785 );
nand ( n42872 , n42870 , n42871 , n42858 );
not ( n42873 , n42858 );
nand ( n42874 , n42873 , n42871 , n42862 );
nand ( n42875 , n42869 , n42872 , n42874 );
nand ( n42876 , n42875 , n2628 );
nand ( n42877 , n42174 , n42876 );
not ( n42878 , n2629 );
buf ( n42879 , n40912 );
not ( n42880 , n42879 );
buf ( n42881 , n40946 );
and ( n42882 , n41016 , n42881 );
buf ( n42883 , n41033 );
nand ( n42884 , n42883 , n40977 , n41080 );
not ( n42885 , n42884 );
nand ( n42886 , n42882 , n36966 , n42885 );
not ( n42887 , n42886 );
or ( n42888 , n42880 , n42887 );
or ( n42889 , n42879 , n42886 );
nand ( n42890 , n42888 , n42889 );
not ( n42891 , n42890 );
or ( n42892 , n42878 , n42891 );
not ( n42893 , n42599 );
buf ( n42894 , n42782 );
and ( n42895 , n42893 , n42894 );
and ( n42896 , n42592 , n42894 );
nor ( n42897 , n42895 , n42896 );
not ( n42898 , n42590 );
not ( n42899 , n42894 );
nand ( n42900 , n42898 , n42899 , n42556 );
not ( n42901 , n42556 );
nand ( n42902 , n42901 , n42899 , n42590 );
nand ( n42903 , n42897 , n42900 , n42902 );
nand ( n42904 , n42903 , n2628 );
nand ( n42905 , n42892 , n42904 );
not ( n42906 , n2629 );
nand ( n42907 , n42885 , n36966 );
buf ( n42908 , n41016 );
not ( n42909 , n42908 );
and ( n42910 , n42907 , n42909 );
not ( n42911 , n42907 );
and ( n42912 , n42911 , n42908 );
nor ( n42913 , n42910 , n42912 );
not ( n42914 , n42913 );
or ( n42915 , n42906 , n42914 );
xor ( n42916 , n42711 , n42713 );
xor ( n42917 , n42916 , n42776 );
nand ( n42918 , n42917 , n2628 );
nand ( n42919 , n42915 , n42918 );
xor ( n42920 , n42734 , n42736 );
xor ( n42921 , n42920 , n42773 );
not ( n42922 , n42921 );
and ( n42923 , n2628 , n42922 );
not ( n42924 , n2628 );
not ( n42925 , n41080 );
buf ( n42926 , n40976 );
nor ( n42927 , n42925 , n42926 );
nand ( n42928 , n36966 , n42927 );
xor ( n42929 , n42928 , n42883 );
and ( n42930 , n42924 , n42929 );
nor ( n42931 , n42923 , n42930 );
and ( n42932 , n42261 , n36988 );
and ( n42933 , n42263 , n496 );
nor ( n42934 , n42932 , n42933 );
or ( n42935 , n42306 , n42934 );
and ( n42936 , n42261 , n42214 );
and ( n42937 , n42263 , n495 );
nor ( n42938 , n42936 , n42937 );
or ( n42939 , n42938 , n42271 );
nand ( n42940 , n42935 , n42939 );
and ( n42941 , n7066 , n42276 );
and ( n42942 , n7065 , n492 );
nor ( n42943 , n42941 , n42942 );
or ( n42944 , n42291 , n42943 );
and ( n42945 , n42294 , n42282 );
and ( n42946 , n7065 , n491 );
nor ( n42947 , n42945 , n42946 );
or ( n42948 , n42293 , n42947 );
nand ( n42949 , n42944 , n42948 );
xor ( n42950 , n42940 , n42949 );
and ( n42951 , n42316 , n7092 );
and ( n42952 , n41312 , n498 );
nor ( n42953 , n42951 , n42952 );
not ( n42954 , n42953 );
not ( n42955 , n42954 );
not ( n42956 , n42315 );
not ( n42957 , n42956 );
or ( n42958 , n42955 , n42957 );
and ( n42959 , n42316 , n7081 );
and ( n42960 , n41312 , n497 );
nor ( n42961 , n42959 , n42960 );
or ( n42962 , n42321 , n42961 );
nand ( n42963 , n42958 , n42962 );
and ( n42964 , n42950 , n42963 );
and ( n42965 , n42940 , n42949 );
or ( n42966 , n42964 , n42965 );
or ( n42967 , n7136 , n7139 );
nand ( n42968 , n42967 , n7350 );
and ( n42969 , n35943 , n42419 );
and ( n42970 , n42216 , n490 );
nor ( n42971 , n42969 , n42970 );
or ( n42972 , n7214 , n42971 );
and ( n42973 , n35943 , n5539 );
and ( n42974 , n42216 , n489 );
nor ( n42975 , n42973 , n42974 );
or ( n42976 , n42220 , n42975 );
nand ( n42977 , n42972 , n42976 );
xor ( n42978 , n42968 , n42977 );
not ( n42979 , n42210 );
and ( n42980 , n42204 , n42382 );
and ( n42981 , n42189 , n493 );
nor ( n42982 , n42980 , n42981 );
not ( n42983 , n42982 );
not ( n42984 , n42983 );
or ( n42985 , n42979 , n42984 );
and ( n42986 , n42204 , n42221 );
and ( n42987 , n42206 , n494 );
nor ( n42988 , n42986 , n42987 );
or ( n42989 , n42457 , n42988 );
nand ( n42990 , n42985 , n42989 );
and ( n42991 , n42978 , n42990 );
and ( n42992 , n42968 , n42977 );
or ( n42993 , n42991 , n42992 );
xor ( n42994 , n42966 , n42993 );
and ( n42995 , n42261 , n42221 );
and ( n42996 , n42263 , n494 );
nor ( n42997 , n42995 , n42996 );
or ( n42998 , n42997 , n42271 );
or ( n42999 , n42306 , n42938 );
nand ( n43000 , n42998 , n42999 );
or ( n43001 , n42315 , n42961 );
and ( n43002 , n42316 , n36988 );
and ( n43003 , n41312 , n496 );
nor ( n43004 , n43002 , n43003 );
or ( n43005 , n43004 , n42321 );
nand ( n43006 , n43001 , n43005 );
xor ( n43007 , n43000 , n43006 );
or ( n43008 , n7214 , n42975 );
or ( n43009 , n42220 , n42216 );
nand ( n43010 , n43008 , n43009 );
xor ( n43011 , n43007 , n43010 );
and ( n43012 , n42994 , n43011 );
and ( n43013 , n42966 , n42993 );
or ( n43014 , n43012 , n43013 );
not ( n43015 , n42220 );
or ( n43016 , n7215 , n43015 );
nand ( n43017 , n43016 , n35943 );
and ( n43018 , n42294 , n42419 );
and ( n43019 , n7065 , n490 );
nor ( n43020 , n43018 , n43019 );
or ( n43021 , n42291 , n43020 );
and ( n43022 , n42294 , n5539 );
and ( n43023 , n7065 , n489 );
nor ( n43024 , n43022 , n43023 );
or ( n43025 , n42293 , n43024 );
nand ( n43026 , n43021 , n43025 );
xor ( n43027 , n43017 , n43026 );
or ( n43028 , n42306 , n42997 );
and ( n43029 , n42261 , n42382 );
and ( n43030 , n42263 , n493 );
nor ( n43031 , n43029 , n43030 );
or ( n43032 , n42271 , n43031 );
nand ( n43033 , n43028 , n43032 );
xor ( n43034 , n43027 , n43033 );
buf ( n43035 , n42316 );
not ( n43036 , n43035 );
nor ( n43037 , n43036 , n7092 );
or ( n43038 , n42457 , n42982 );
and ( n43039 , n42204 , n42276 );
and ( n43040 , n42189 , n492 );
nor ( n43041 , n43039 , n43040 );
or ( n43042 , n42456 , n43041 );
nand ( n43043 , n43038 , n43042 );
xor ( n43044 , n43037 , n43043 );
or ( n43045 , n42291 , n42947 );
or ( n43046 , n42293 , n43020 );
nand ( n43047 , n43045 , n43046 );
not ( n43048 , n43047 );
and ( n43049 , n43044 , n43048 );
and ( n43050 , n43037 , n43043 );
or ( n43051 , n43049 , n43050 );
xor ( n43052 , n43034 , n43051 );
xor ( n43053 , n43000 , n43006 );
and ( n43054 , n43053 , n43010 );
and ( n43055 , n43000 , n43006 );
or ( n43056 , n43054 , n43055 );
xor ( n43057 , n43047 , n43056 );
or ( n43058 , n42315 , n43004 );
and ( n43059 , n43035 , n42214 );
and ( n43060 , n41312 , n495 );
nor ( n43061 , n43059 , n43060 );
or ( n43062 , n43061 , n42321 );
nand ( n43063 , n43058 , n43062 );
or ( n43064 , n42457 , n43041 );
and ( n43065 , n42204 , n42282 );
and ( n43066 , n42189 , n491 );
nor ( n43067 , n43065 , n43066 );
or ( n43068 , n42456 , n43067 );
nand ( n43069 , n43064 , n43068 );
xor ( n43070 , n43063 , n43069 );
nor ( n43071 , n41312 , n7081 );
xor ( n43072 , n43070 , n43071 );
xor ( n43073 , n43057 , n43072 );
xor ( n43074 , n43052 , n43073 );
xor ( n43075 , n43014 , n43074 );
xor ( n43076 , n43037 , n43043 );
xor ( n43077 , n43076 , n43048 );
nor ( n43078 , n43036 , n1970 );
and ( n43079 , n7350 , n5539 );
and ( n43080 , n7124 , n489 );
nor ( n43081 , n43079 , n43080 );
not ( n43082 , n43081 );
and ( n43083 , n7136 , n43082 );
and ( n43084 , n7139 , n7350 );
nor ( n43085 , n43083 , n43084 );
not ( n43086 , n43085 );
xor ( n43087 , n43078 , n43086 );
and ( n43088 , n35943 , n42282 );
and ( n43089 , n42216 , n491 );
nor ( n43090 , n43088 , n43089 );
or ( n43091 , n7214 , n43090 );
or ( n43092 , n42220 , n42971 );
nand ( n43093 , n43091 , n43092 );
and ( n43094 , n42186 , n495 );
and ( n43095 , n42204 , n42214 );
nor ( n43096 , n43094 , n43095 );
or ( n43097 , n42457 , n43096 );
or ( n43098 , n42988 , n36982 );
nand ( n43099 , n43097 , n43098 );
xor ( n43100 , n43093 , n43099 );
and ( n43101 , n42261 , n7081 );
and ( n43102 , n42263 , n497 );
nor ( n43103 , n43101 , n43102 );
or ( n43104 , n42306 , n43103 );
or ( n43105 , n42271 , n42934 );
nand ( n43106 , n43104 , n43105 );
and ( n43107 , n43100 , n43106 );
and ( n43108 , n43093 , n43099 );
or ( n43109 , n43107 , n43108 );
and ( n43110 , n43087 , n43109 );
and ( n43111 , n43078 , n43086 );
or ( n43112 , n43110 , n43111 );
xor ( n43113 , n43077 , n43112 );
or ( n43114 , n42943 , n42293 );
and ( n43115 , n7157 , n42382 );
and ( n43116 , n7065 , n493 );
nor ( n43117 , n43115 , n43116 );
not ( n43118 , n43117 );
nand ( n43119 , n43118 , n42290 );
nand ( n43120 , n43114 , n43119 );
and ( n43121 , n42316 , n1970 );
and ( n43122 , n41312 , n499 );
nor ( n43123 , n43121 , n43122 );
or ( n43124 , n42315 , n43123 );
or ( n43125 , n42953 , n42321 );
nand ( n43126 , n43124 , n43125 );
xor ( n43127 , n43120 , n43126 );
nor ( n43128 , n41312 , n7140 );
and ( n43129 , n43127 , n43128 );
and ( n43130 , n43120 , n43126 );
or ( n43131 , n43129 , n43130 );
xor ( n43132 , n42940 , n42949 );
xor ( n43133 , n43132 , n42963 );
xor ( n43134 , n43131 , n43133 );
xor ( n43135 , n42968 , n42977 );
xor ( n43136 , n43135 , n42990 );
and ( n43137 , n43134 , n43136 );
and ( n43138 , n43131 , n43133 );
or ( n43139 , n43137 , n43138 );
and ( n43140 , n43113 , n43139 );
and ( n43141 , n43077 , n43112 );
or ( n43142 , n43140 , n43141 );
and ( n43143 , n43075 , n43142 );
and ( n43144 , n43014 , n43074 );
or ( n43145 , n43143 , n43144 );
xor ( n43146 , n43047 , n43056 );
and ( n43147 , n43146 , n43072 );
and ( n43148 , n43047 , n43056 );
or ( n43149 , n43147 , n43148 );
xor ( n43150 , n43017 , n43026 );
and ( n43151 , n43150 , n43033 );
and ( n43152 , n43017 , n43026 );
or ( n43153 , n43151 , n43152 );
or ( n43154 , n42315 , n43061 );
and ( n43155 , n43035 , n42221 );
and ( n43156 , n41312 , n494 );
nor ( n43157 , n43155 , n43156 );
or ( n43158 , n43157 , n42321 );
nand ( n43159 , n43154 , n43158 );
nor ( n43160 , n43036 , n36988 );
xor ( n43161 , n43159 , n43160 );
or ( n43162 , n42291 , n43024 );
or ( n43163 , n42293 , n7065 );
nand ( n43164 , n43162 , n43163 );
xor ( n43165 , n43161 , n43164 );
xor ( n43166 , n43153 , n43165 );
or ( n43167 , n42306 , n43031 );
and ( n43168 , n42261 , n42276 );
and ( n43169 , n42263 , n492 );
nor ( n43170 , n43168 , n43169 );
or ( n43171 , n42271 , n43170 );
nand ( n43172 , n43167 , n43171 );
or ( n43173 , n42457 , n43067 );
and ( n43174 , n42204 , n42419 );
and ( n43175 , n42189 , n490 );
nor ( n43176 , n43174 , n43175 );
or ( n43177 , n42456 , n43176 );
nand ( n43178 , n43173 , n43177 );
not ( n43179 , n43178 );
xor ( n43180 , n43172 , n43179 );
xor ( n43181 , n43063 , n43069 );
and ( n43182 , n43181 , n43071 );
and ( n43183 , n43063 , n43069 );
or ( n43184 , n43182 , n43183 );
xor ( n43185 , n43180 , n43184 );
xor ( n43186 , n43166 , n43185 );
xor ( n43187 , n43149 , n43186 );
xor ( n43188 , n43034 , n43051 );
and ( n43189 , n43188 , n43073 );
and ( n43190 , n43034 , n43051 );
or ( n43191 , n43189 , n43190 );
xor ( n43192 , n43187 , n43191 );
or ( n43193 , n43145 , n43192 );
nand ( n43194 , n43145 , n43192 );
nand ( n43195 , n43193 , n43194 );
not ( n43196 , n43195 );
not ( n43197 , n42784 );
buf ( n43198 , n42866 );
nand ( n43199 , n43197 , n43198 );
xor ( n43200 , n43131 , n43133 );
xor ( n43201 , n43200 , n43136 );
xor ( n43202 , n43078 , n43086 );
xor ( n43203 , n43202 , n43109 );
or ( n43204 , n7299 , n42834 );
or ( n43205 , n42281 , n43081 );
nand ( n43206 , n43204 , n43205 );
or ( n43207 , n7118 , n7071 );
nand ( n43208 , n43207 , n7074 );
or ( n43209 , n43206 , n43208 );
xor ( n43210 , n43085 , n43209 );
nor ( n43211 , n41311 , n7122 );
or ( n43212 , n42175 , n42815 );
or ( n43213 , n43117 , n42293 );
nand ( n43214 , n43212 , n43213 );
xor ( n43215 , n43211 , n43214 );
not ( n43216 , n43096 );
not ( n43217 , n43216 );
not ( n43218 , n42456 );
not ( n43219 , n43218 );
or ( n43220 , n43217 , n43219 );
not ( n43221 , n42823 );
nand ( n43222 , n43221 , n42201 );
nand ( n43223 , n43220 , n43222 );
and ( n43224 , n43215 , n43223 );
and ( n43225 , n43211 , n43214 );
or ( n43226 , n43224 , n43225 );
and ( n43227 , n43210 , n43226 );
and ( n43228 , n43085 , n43209 );
or ( n43229 , n43227 , n43228 );
xor ( n43230 , n43203 , n43229 );
or ( n43231 , n7214 , n42793 );
or ( n43232 , n42220 , n43090 );
nand ( n43233 , n43231 , n43232 );
or ( n43234 , n42260 , n42799 );
or ( n43235 , n43103 , n42271 );
nand ( n43236 , n43234 , n43235 );
xor ( n43237 , n43233 , n43236 );
or ( n43238 , n42315 , n42806 );
or ( n43239 , n43123 , n42321 );
nand ( n43240 , n43238 , n43239 );
and ( n43241 , n43237 , n43240 );
and ( n43242 , n43233 , n43236 );
or ( n43243 , n43241 , n43242 );
xor ( n43244 , n43120 , n43126 );
xor ( n43245 , n43244 , n43128 );
xor ( n43246 , n43243 , n43245 );
xor ( n43247 , n43093 , n43099 );
xor ( n43248 , n43247 , n43106 );
and ( n43249 , n43246 , n43248 );
and ( n43250 , n43243 , n43245 );
or ( n43251 , n43249 , n43250 );
xor ( n43252 , n43230 , n43251 );
xor ( n43253 , n43201 , n43252 );
and ( n43254 , n42830 , n42836 );
xor ( n43255 , n42817 , n42818 );
and ( n43256 , n43255 , n42825 );
and ( n43257 , n42817 , n42818 );
or ( n43258 , n43256 , n43257 );
xor ( n43259 , n43254 , n43258 );
xor ( n43260 , n42795 , n42801 );
and ( n43261 , n43260 , n42808 );
and ( n43262 , n42795 , n42801 );
or ( n43263 , n43261 , n43262 );
and ( n43264 , n43259 , n43263 );
and ( n43265 , n43254 , n43258 );
or ( n43266 , n43264 , n43265 );
xor ( n43267 , n43085 , n43209 );
xor ( n43268 , n43267 , n43226 );
xor ( n43269 , n43266 , n43268 );
xor ( n43270 , n43233 , n43236 );
xor ( n43271 , n43270 , n43240 );
not ( n43272 , n43208 );
not ( n43273 , n43206 );
or ( n43274 , n43272 , n43273 );
nand ( n43275 , n43274 , n43209 );
xor ( n43276 , n43271 , n43275 );
xor ( n43277 , n43211 , n43214 );
xor ( n43278 , n43277 , n43223 );
and ( n43279 , n43276 , n43278 );
and ( n43280 , n43271 , n43275 );
or ( n43281 , n43279 , n43280 );
and ( n43282 , n43269 , n43281 );
and ( n43283 , n43266 , n43268 );
or ( n43284 , n43282 , n43283 );
xor ( n43285 , n43253 , n43284 );
xor ( n43286 , n43243 , n43245 );
xor ( n43287 , n43286 , n43248 );
and ( n43288 , n42837 , n42841 );
xor ( n43289 , n43254 , n43258 );
xor ( n43290 , n43289 , n43263 );
xor ( n43291 , n43288 , n43290 );
xor ( n43292 , n42789 , n42809 );
and ( n43293 , n43292 , n42826 );
and ( n43294 , n42789 , n42809 );
or ( n43295 , n43293 , n43294 );
and ( n43296 , n43291 , n43295 );
and ( n43297 , n43288 , n43290 );
or ( n43298 , n43296 , n43297 );
xor ( n43299 , n43287 , n43298 );
xor ( n43300 , n43266 , n43268 );
xor ( n43301 , n43300 , n43281 );
and ( n43302 , n43299 , n43301 );
and ( n43303 , n43287 , n43298 );
or ( n43304 , n43302 , n43303 );
nor ( n43305 , n43285 , n43304 );
not ( n43306 , n43305 );
xor ( n43307 , n43201 , n43252 );
and ( n43308 , n43307 , n43284 );
and ( n43309 , n43201 , n43252 );
or ( n43310 , n43308 , n43309 );
xor ( n43311 , n42966 , n42993 );
xor ( n43312 , n43311 , n43011 );
xor ( n43313 , n43077 , n43112 );
xor ( n43314 , n43313 , n43139 );
xor ( n43315 , n43312 , n43314 );
xor ( n43316 , n43203 , n43229 );
and ( n43317 , n43316 , n43251 );
and ( n43318 , n43203 , n43229 );
or ( n43319 , n43317 , n43318 );
xor ( n43320 , n43315 , n43319 );
or ( n43321 , n43310 , n43320 );
xor ( n43322 , n43271 , n43275 );
xor ( n43323 , n43322 , n43278 );
xor ( n43324 , n42842 , n42846 );
and ( n43325 , n43324 , n42851 );
and ( n43326 , n42842 , n42846 );
or ( n43327 , n43325 , n43326 );
xor ( n43328 , n43323 , n43327 );
xor ( n43329 , n43288 , n43290 );
xor ( n43330 , n43329 , n43295 );
xor ( n43331 , n43328 , n43330 );
xor ( n43332 , n42827 , n42852 );
and ( n43333 , n43332 , n42857 );
and ( n43334 , n42827 , n42852 );
or ( n43335 , n43333 , n43334 );
or ( n43336 , n43331 , n43335 );
not ( n43337 , n43336 );
xor ( n43338 , n43323 , n43327 );
and ( n43339 , n43338 , n43330 );
and ( n43340 , n43323 , n43327 );
or ( n43341 , n43339 , n43340 );
not ( n43342 , n43341 );
xor ( n43343 , n43287 , n43298 );
xor ( n43344 , n43343 , n43301 );
not ( n43345 , n43344 );
and ( n43346 , n43342 , n43345 );
buf ( n43347 , n43346 );
nor ( n43348 , n43337 , n43347 );
nand ( n43349 , n42864 , n42866 );
and ( n43350 , n43306 , n43321 , n43348 , n43349 );
and ( n43351 , n43199 , n43350 );
not ( n43352 , n43321 );
not ( n43353 , n43346 );
nand ( n43354 , n43335 , n43331 );
not ( n43355 , n43354 );
and ( n43356 , n43353 , n43355 );
nor ( n43357 , n43345 , n43342 );
nor ( n43358 , n43356 , n43357 );
or ( n43359 , n43358 , n43305 );
nand ( n43360 , n43285 , n43304 );
nand ( n43361 , n43359 , n43360 );
not ( n43362 , n43361 );
or ( n43363 , n43352 , n43362 );
nand ( n43364 , n43310 , n43320 );
nand ( n43365 , n43363 , n43364 );
nor ( n43366 , n43351 , n43365 );
xor ( n43367 , n43312 , n43314 );
and ( n43368 , n43367 , n43319 );
and ( n43369 , n43312 , n43314 );
or ( n43370 , n43368 , n43369 );
xor ( n43371 , n43014 , n43074 );
xor ( n43372 , n43371 , n43142 );
nor ( n43373 , n43370 , n43372 );
nor ( n43374 , n43366 , n43373 );
and ( n43375 , n43370 , n43372 );
or ( n43376 , n43374 , n43375 );
not ( n43377 , n43376 );
or ( n43378 , n43196 , n43377 );
or ( n43379 , n43376 , n43195 );
nand ( n43380 , n43378 , n43379 );
nand ( n43381 , n43380 , n2628 );
not ( n43382 , n43376 );
xor ( n43383 , n43149 , n43186 );
and ( n43384 , n43383 , n43191 );
and ( n43385 , n43149 , n43186 );
or ( n43386 , n43384 , n43385 );
not ( n43387 , n43386 );
xor ( n43388 , n43172 , n43179 );
and ( n43389 , n43388 , n43184 );
and ( n43390 , n43172 , n43179 );
or ( n43391 , n43389 , n43390 );
xor ( n43392 , n43159 , n43160 );
and ( n43393 , n43392 , n43164 );
and ( n43394 , n43159 , n43160 );
or ( n43395 , n43393 , n43394 );
or ( n43396 , n42290 , n7108 );
nand ( n43397 , n43396 , n42294 );
or ( n43398 , n42457 , n43176 );
and ( n43399 , n42204 , n5539 );
and ( n43400 , n42189 , n489 );
nor ( n43401 , n43399 , n43400 );
or ( n43402 , n42456 , n43401 );
nand ( n43403 , n43398 , n43402 );
xor ( n43404 , n43397 , n43403 );
or ( n43405 , n42315 , n43157 );
and ( n43406 , n43035 , n42382 );
and ( n43407 , n43036 , n493 );
nor ( n43408 , n43406 , n43407 );
or ( n43409 , n42321 , n43408 );
nand ( n43410 , n43405 , n43409 );
xor ( n43411 , n43404 , n43410 );
xor ( n43412 , n43395 , n43411 );
nor ( n43413 , n43036 , n42214 );
or ( n43414 , n42306 , n43170 );
and ( n43415 , n42261 , n42282 );
and ( n43416 , n42263 , n491 );
nor ( n43417 , n43415 , n43416 );
or ( n43418 , n42271 , n43417 );
nand ( n43419 , n43414 , n43418 );
xor ( n43420 , n43413 , n43419 );
xor ( n43421 , n43420 , n43178 );
xor ( n43422 , n43412 , n43421 );
xor ( n43423 , n43391 , n43422 );
xor ( n43424 , n43153 , n43165 );
and ( n43425 , n43424 , n43185 );
and ( n43426 , n43153 , n43165 );
or ( n43427 , n43425 , n43426 );
xor ( n43428 , n43423 , n43427 );
not ( n43429 , n43428 );
nand ( n43430 , n43387 , n43429 );
not ( n43431 , n43430 );
nor ( n43432 , n43387 , n43429 );
nor ( n43433 , n43431 , n43432 );
and ( n43434 , n43433 , n43194 );
nand ( n43435 , n43382 , n43434 );
not ( n43436 , n43193 );
nor ( n43437 , n43433 , n43436 );
nand ( n43438 , n43376 , n43437 );
and ( n43439 , n43433 , n43436 , n43194 );
nor ( n43440 , n43433 , n43194 );
nor ( n43441 , n43439 , n43440 );
nand ( n43442 , n43435 , n43438 , n43441 );
nand ( n43443 , n43442 , n2628 );
buf ( n43444 , n43366 );
nor ( n43445 , n43375 , n43373 );
xnor ( n43446 , n43444 , n43445 );
nand ( n43447 , n43446 , n2628 );
not ( n43448 , n36965 );
buf ( n43449 , n41082 );
nand ( n43450 , n43448 , n43449 );
not ( n43451 , n42881 );
and ( n43452 , n43450 , n43451 );
not ( n43453 , n43450 );
and ( n43454 , n43453 , n42881 );
nor ( n43455 , n43452 , n43454 );
nand ( n43456 , n43455 , n2629 );
buf ( n43457 , n2053 );
buf ( n43458 , n1735 );
nand ( n43459 , n43457 , n43458 );
buf ( n43460 , n43459 );
nand ( n43461 , n30476 , n454 );
or ( n43462 , n43460 , n43461 );
not ( n43463 , n31309 );
buf ( n43464 , n31315 );
not ( n43465 , n43464 );
buf ( n43466 , n31231 );
nor ( n43467 , n43465 , n43466 );
buf ( n43468 , n43467 );
not ( n43469 , n43468 );
or ( n43470 , n43463 , n43469 );
or ( n43471 , n43468 , n31309 );
nand ( n43472 , n43470 , n43471 );
or ( n43473 , n454 , n43472 );
not ( n43474 , n30476 );
nand ( n43475 , n43474 , n43460 , n454 );
nand ( n43476 , n43462 , n43473 , n43475 );
not ( n43477 , n43476 );
not ( n43478 , n7387 );
not ( n43479 , n7360 );
nand ( n43480 , n43479 , n7390 );
not ( n43481 , n43480 );
or ( n43482 , n43478 , n43481 );
or ( n43483 , n43480 , n7387 );
nand ( n43484 , n43482 , n43483 );
and ( n43485 , n2628 , n43484 );
not ( n43486 , n2628 );
not ( n43487 , n7036 );
not ( n43488 , n7033 );
or ( n43489 , n43487 , n43488 );
nand ( n43490 , n43489 , n6980 );
nand ( n43491 , n7006 , n7040 );
xnor ( n43492 , n43490 , n43491 );
and ( n43493 , n43486 , n43492 );
or ( n43494 , n43485 , n43493 );
not ( n43495 , n454 );
not ( n43496 , n41995 );
or ( n43497 , n43495 , n43496 );
nand ( n43498 , n43497 , n42170 );
not ( n43499 , n43498 );
not ( n43500 , n39597 );
not ( n43501 , n41442 );
not ( n43502 , n43501 );
or ( n43503 , n43500 , n43502 );
nand ( n43504 , n43503 , n41985 );
nand ( n43505 , C1 , n43504 );
buf ( n43506 , n43505 );
not ( n43507 , n41976 );
not ( n43508 , n41983 );
or ( n43509 , n43507 , n43508 );
not ( n43510 , n41242 );
not ( n43511 , n41434 );
or ( n43512 , n43510 , n43511 );
nand ( n43513 , n43512 , n39597 );
nand ( n43514 , n43509 , n43513 );
not ( n43515 , n43514 );
not ( n43516 , n43515 );
nor ( n43517 , n43516 , n41090 );
nor ( n43518 , n43506 , n43517 );
not ( n43519 , n43518 );
buf ( n43520 , n43514 );
nor ( n43521 , n43520 , n41658 );
nand ( n43522 , n43521 , n41025 );
not ( n43523 , n43522 );
or ( n43524 , n43519 , n43523 );
not ( n43525 , n41948 );
and ( n43526 , n41961 , n41427 );
buf ( n43527 , n41968 );
nand ( n43528 , n43526 , n41972 , n43527 );
not ( n43529 , n43528 );
not ( n43530 , n43529 );
or ( n43531 , n43525 , n43530 );
and ( n43532 , n41950 , n41948 );
xor ( n43533 , n41895 , n41920 );
and ( n43534 , n43533 , n41927 );
and ( n43535 , n41895 , n41920 );
or ( n43536 , n43534 , n43535 );
buf ( n43537 , n43536 );
buf ( n43538 , n43537 );
xor ( n43539 , n41829 , n41842 );
and ( n43540 , n43539 , n41860 );
and ( n43541 , n41829 , n41842 );
or ( n43542 , n43540 , n43541 );
buf ( n43543 , n43542 );
buf ( n43544 , n43543 );
not ( n43545 , n2724 );
not ( n43546 , n32280 );
or ( n43547 , n43545 , n43546 );
nand ( n43548 , n43547 , n495 );
buf ( n43549 , n43548 );
buf ( n43550 , n39149 );
not ( n43551 , n43550 );
buf ( n43552 , n41852 );
not ( n43553 , n43552 );
or ( n43554 , n43551 , n43553 );
buf ( n43555 , n489 );
buf ( n43556 , n31826 );
xor ( n43557 , n43555 , n43556 );
buf ( n43558 , n43557 );
buf ( n43559 , n43558 );
buf ( n43560 , n36508 );
nand ( n43561 , n43559 , n43560 );
buf ( n43562 , n43561 );
buf ( n43563 , n43562 );
nand ( n43564 , n43554 , n43563 );
buf ( n43565 , n43564 );
buf ( n43566 , n43565 );
xor ( n43567 , n43549 , n43566 );
buf ( n43568 , n3146 );
not ( n43569 , n43568 );
buf ( n43570 , n41909 );
not ( n43571 , n43570 );
or ( n43572 , n43569 , n43571 );
buf ( n43573 , n493 );
not ( n43574 , n43573 );
buf ( n43575 , n41312 );
not ( n43576 , n43575 );
or ( n43577 , n43574 , n43576 );
buf ( n43578 , n41316 );
buf ( n43579 , n2704 );
nand ( n43580 , n43578 , n43579 );
buf ( n43581 , n43580 );
buf ( n43582 , n43581 );
nand ( n43583 , n43577 , n43582 );
buf ( n43584 , n43583 );
buf ( n43585 , n43584 );
buf ( n43586 , n3113 );
nand ( n43587 , n43585 , n43586 );
buf ( n43588 , n43587 );
buf ( n43589 , n43588 );
nand ( n43590 , n43572 , n43589 );
buf ( n43591 , n43590 );
buf ( n43592 , n43591 );
xor ( n43593 , n43567 , n43592 );
buf ( n43594 , n43593 );
buf ( n43595 , n43594 );
xor ( n43596 , n43544 , n43595 );
and ( n43597 , n38391 , n489 );
buf ( n43598 , n43597 );
buf ( n43599 , n34465 );
not ( n43600 , n43599 );
buf ( n43601 , n41887 );
not ( n43602 , n43601 );
or ( n43603 , n43600 , n43602 );
buf ( n43604 , n491 );
not ( n43605 , n43604 );
buf ( n43606 , n38410 );
not ( n43607 , n43606 );
or ( n43608 , n43605 , n43607 );
buf ( n43609 , n38414 );
buf ( n43610 , n3524 );
nand ( n43611 , n43609 , n43610 );
buf ( n43612 , n43611 );
buf ( n43613 , n43612 );
nand ( n43614 , n43608 , n43613 );
buf ( n43615 , n43614 );
buf ( n43616 , n43615 );
buf ( n43617 , n3045 );
nand ( n43618 , n43616 , n43617 );
buf ( n43619 , n43618 );
buf ( n43620 , n43619 );
nand ( n43621 , n43603 , n43620 );
buf ( n43622 , n43621 );
buf ( n43623 , n43622 );
xor ( n43624 , n43598 , n43623 );
buf ( n43625 , n41916 );
xor ( n43626 , n43624 , n43625 );
buf ( n43627 , n43626 );
buf ( n43628 , n43627 );
xor ( n43629 , n43596 , n43628 );
buf ( n43630 , n43629 );
buf ( n43631 , n43630 );
xor ( n43632 , n43538 , n43631 );
xor ( n43633 , n41863 , n41869 );
and ( n43634 , n43633 , n41930 );
and ( n43635 , n41863 , n41869 );
or ( n43636 , n43634 , n43635 );
buf ( n43637 , n43636 );
buf ( n43638 , n43637 );
xor ( n43639 , n43632 , n43638 );
buf ( n43640 , n43639 );
xor ( n43641 , n41826 , n41933 );
and ( n43642 , n43641 , n41940 );
and ( n43643 , n41826 , n41933 );
or ( n43644 , n43642 , n43643 );
buf ( n43645 , n43644 );
nand ( n43646 , n43640 , n43645 );
not ( n43647 , n43646 );
nor ( n43648 , n43640 , n43645 );
nor ( n43649 , n43647 , n43648 );
nor ( n43650 , n43532 , n43649 , n29519 );
nand ( n43651 , n43531 , n43650 );
not ( n43652 , n41816 );
and ( n43653 , n41682 , n41226 );
nand ( n43654 , n43653 , n41671 , n41689 );
nand ( n43655 , n43654 , n41815 );
not ( n43656 , n43655 );
or ( n43657 , n43652 , n43656 );
xor ( n43658 , n41770 , n41791 );
and ( n43659 , n43658 , n41798 );
and ( n43660 , n41770 , n41791 );
or ( n43661 , n43659 , n43660 );
buf ( n43662 , n43661 );
buf ( n43663 , n43662 );
xor ( n43664 , n41706 , n41726 );
and ( n43665 , n43664 , n41741 );
and ( n43666 , n41706 , n41726 );
or ( n43667 , n43665 , n43666 );
buf ( n43668 , n43667 );
buf ( n43669 , n43668 );
and ( n43670 , n41193 , n41194 );
buf ( n43671 , n43670 );
not ( n43672 , n41762 );
not ( n43673 , n33967 );
or ( n43674 , n43672 , n43673 );
buf ( n43675 , n491 );
buf ( n43676 , n507 );
xnor ( n43677 , n43675 , n43676 );
buf ( n43678 , n43677 );
buf ( n43679 , n43678 );
not ( n43680 , n43679 );
buf ( n43681 , n33973 );
nand ( n43682 , n43680 , n43681 );
buf ( n43683 , n43682 );
nand ( n43684 , n43674 , n43683 );
xor ( n43685 , n43671 , n43684 );
xor ( n43686 , n43685 , n41787 );
buf ( n43687 , n43686 );
xor ( n43688 , n43669 , n43687 );
buf ( n43689 , n41710 );
not ( n43690 , n43689 );
buf ( n43691 , n41718 );
not ( n43692 , n43691 );
or ( n43693 , n43690 , n43692 );
buf ( n43694 , n37254 );
buf ( n43695 , n489 );
buf ( n43696 , n509 );
xor ( n43697 , n43695 , n43696 );
buf ( n43698 , n43697 );
buf ( n43699 , n43698 );
nand ( n43700 , n43694 , n43699 );
buf ( n43701 , n43700 );
buf ( n43702 , n43701 );
nand ( n43703 , n43693 , n43702 );
buf ( n43704 , n43703 );
buf ( n43705 , n43704 );
buf ( n43706 , n33167 );
not ( n43707 , n43706 );
buf ( n43708 , n43707 );
buf ( n43709 , n43708 );
not ( n43710 , n43709 );
buf ( n43711 , n41735 );
not ( n43712 , n43711 );
or ( n43713 , n43710 , n43712 );
buf ( n43714 , n495 );
nand ( n43715 , n43713 , n43714 );
buf ( n43716 , n43715 );
buf ( n43717 , n43716 );
xor ( n43718 , n43705 , n43717 );
buf ( n43719 , n493 );
buf ( n43720 , n505 );
and ( n43721 , n43719 , n43720 );
not ( n43722 , n43719 );
buf ( n43723 , n505 );
not ( n43724 , n43723 );
buf ( n43725 , n43724 );
buf ( n43726 , n43725 );
and ( n43727 , n43722 , n43726 );
nor ( n43728 , n43721 , n43727 );
buf ( n43729 , n43728 );
buf ( n43730 , n43729 );
not ( n43731 , n43730 );
not ( n43732 , n41776 );
buf ( n43733 , n43732 );
not ( n43734 , n43733 );
or ( n43735 , n43731 , n43734 );
buf ( n43736 , n4242 );
buf ( n43737 , n41781 );
or ( n43738 , n43736 , n43737 );
nand ( n43739 , n43735 , n43738 );
buf ( n43740 , n43739 );
buf ( n43741 , n43740 );
xor ( n43742 , n43718 , n43741 );
buf ( n43743 , n43742 );
buf ( n43744 , n43743 );
xor ( n43745 , n43688 , n43744 );
buf ( n43746 , n43745 );
buf ( n43747 , n43746 );
xor ( n43748 , n43663 , n43747 );
xor ( n43749 , n41744 , n41750 );
and ( n43750 , n43749 , n41801 );
and ( n43751 , n41744 , n41750 );
or ( n43752 , n43750 , n43751 );
buf ( n43753 , n43752 );
buf ( n43754 , n43753 );
xor ( n43755 , n43748 , n43754 );
buf ( n43756 , n43755 );
xor ( n43757 , n41703 , n41804 );
and ( n43758 , n43757 , n41811 );
and ( n43759 , n41703 , n41804 );
or ( n43760 , n43758 , n43759 );
buf ( n43761 , n43760 );
and ( n43762 , n43756 , n43761 );
nor ( n43763 , n43756 , n43761 );
nor ( n43764 , n43762 , n43763 );
nor ( n43765 , n43764 , n455 );
nand ( n43766 , n43657 , n43765 );
not ( n43767 , n41950 );
not ( n43768 , n43767 );
not ( n43769 , n43528 );
or ( n43770 , n43768 , n43769 );
and ( n43771 , n43649 , n41948 , n455 );
nand ( n43772 , n43770 , n43771 );
and ( n43773 , n43764 , n41816 , n29519 );
nand ( n43774 , n43655 , n43773 );
nand ( n43775 , n43651 , n43766 , n43772 , n43774 );
not ( n43776 , n43775 );
not ( n43777 , n43776 );
nor ( n43778 , n43777 , n41985 );
not ( n43779 , n43778 );
not ( n43780 , n29519 );
not ( n43781 , n41818 );
or ( n43782 , n43780 , n43781 );
nand ( n43783 , n43782 , n41975 );
not ( n43784 , n43783 );
nand ( n43785 , n43651 , n43766 , n43772 , n43774 );
nand ( n43786 , n43784 , n43785 );
buf ( n43787 , n43786 );
nand ( n43788 , n43779 , n43787 );
not ( n43789 , n43788 );
nor ( n43790 , n43789 , n2618 );
nand ( n43791 , n43524 , n43790 );
not ( n43792 , n454 );
nor ( n43793 , n43792 , n43788 );
nand ( n43794 , n43522 , n43793 , n43518 );
buf ( n43795 , n41639 );
buf ( n43796 , n42142 );
not ( n43797 , n43796 );
buf ( n43798 , n41612 );
nand ( n43799 , n43797 , n43798 );
buf ( n43800 , n43799 );
buf ( n43801 , n43800 );
nor ( n43802 , n43795 , n43801 );
buf ( n43803 , n43802 );
buf ( n43804 , n43803 );
or ( n43805 , n41617 , n42142 );
nand ( n43806 , n43805 , n42148 );
buf ( n43807 , n43806 );
or ( n43808 , n43804 , n43807 );
buf ( n43809 , n43808 );
xor ( n43810 , n42003 , n42127 );
and ( n43811 , n43810 , n42134 );
and ( n43812 , n42003 , n42127 );
or ( n43813 , n43811 , n43812 );
buf ( n43814 , n43813 );
buf ( n43815 , n43814 );
xor ( n43816 , n42050 , n42056 );
and ( n43817 , n43816 , n42063 );
and ( n43818 , n42050 , n42056 );
or ( n43819 , n43817 , n43818 );
buf ( n43820 , n43819 );
buf ( n43821 , n43820 );
xor ( n43822 , n42079 , n42098 );
and ( n43823 , n43822 , n42118 );
and ( n43824 , n42079 , n42098 );
or ( n43825 , n43823 , n43824 );
buf ( n43826 , n43825 );
buf ( n43827 , n43826 );
xor ( n43828 , n43821 , n43827 );
xor ( n43829 , n42084 , n42089 );
and ( n43830 , n43829 , n42095 );
and ( n43831 , n42084 , n42089 );
or ( n43832 , n43830 , n43831 );
buf ( n43833 , n43832 );
buf ( n43834 , n43833 );
xor ( n43835 , n42104 , n42109 );
and ( n43836 , n43835 , n42115 );
and ( n43837 , n42104 , n42109 );
or ( n43838 , n43836 , n43837 );
buf ( n43839 , n43838 );
buf ( n43840 , n43839 );
xor ( n43841 , n43834 , n43840 );
xor ( n43842 , n42008 , n42013 );
and ( n43843 , n43842 , n42019 );
and ( n43844 , n42008 , n42013 );
or ( n43845 , n43843 , n43844 );
buf ( n43846 , n43845 );
buf ( n43847 , n43846 );
xor ( n43848 , n43841 , n43847 );
buf ( n43849 , n43848 );
buf ( n43850 , n43849 );
xor ( n43851 , n43828 , n43850 );
buf ( n43852 , n43851 );
buf ( n43853 , n43852 );
buf ( n43854 , n521 );
buf ( n43855 , n545 );
and ( n43856 , n43854 , n43855 );
buf ( n43857 , n43856 );
buf ( n43858 , n43857 );
buf ( n43859 , n522 );
buf ( n43860 , n544 );
and ( n43861 , n43859 , n43860 );
buf ( n43862 , n43861 );
buf ( n43863 , n43862 );
xor ( n43864 , n43858 , n43863 );
buf ( n43865 , n524 );
buf ( n43866 , n542 );
and ( n43867 , n43865 , n43866 );
buf ( n43868 , n43867 );
buf ( n43869 , n43868 );
xor ( n43870 , n43864 , n43869 );
buf ( n43871 , n43870 );
buf ( n43872 , n43871 );
buf ( n43873 , n523 );
buf ( n43874 , n543 );
and ( n43875 , n43873 , n43874 );
buf ( n43876 , n43875 );
buf ( n43877 , n43876 );
buf ( n43878 , n526 );
buf ( n43879 , n540 );
and ( n43880 , n43878 , n43879 );
buf ( n43881 , n43880 );
buf ( n43882 , n43881 );
xor ( n43883 , n43877 , n43882 );
buf ( n43884 , n527 );
buf ( n43885 , n539 );
and ( n43886 , n43884 , n43885 );
buf ( n43887 , n43886 );
buf ( n43888 , n43887 );
xor ( n43889 , n43883 , n43888 );
buf ( n43890 , n43889 );
buf ( n43891 , n43890 );
xor ( n43892 , n43872 , n43891 );
buf ( n43893 , n528 );
buf ( n43894 , n538 );
and ( n43895 , n43893 , n43894 );
buf ( n43896 , n43895 );
buf ( n43897 , n43896 );
buf ( n43898 , n529 );
buf ( n43899 , n537 );
and ( n43900 , n43898 , n43899 );
buf ( n43901 , n43900 );
buf ( n43902 , n43901 );
xor ( n43903 , n43897 , n43902 );
buf ( n43904 , n525 );
buf ( n43905 , n541 );
and ( n43906 , n43904 , n43905 );
buf ( n43907 , n43906 );
buf ( n43908 , n43907 );
xor ( n43909 , n43903 , n43908 );
buf ( n43910 , n43909 );
buf ( n43911 , n43910 );
xor ( n43912 , n43892 , n43911 );
buf ( n43913 , n43912 );
buf ( n43914 , n43913 );
xor ( n43915 , n42022 , n42028 );
and ( n43916 , n43915 , n42035 );
and ( n43917 , n42022 , n42028 );
or ( n43918 , n43916 , n43917 );
buf ( n43919 , n43918 );
buf ( n43920 , n43919 );
xor ( n43921 , n43914 , n43920 );
xor ( n43922 , n42066 , n42072 );
and ( n43923 , n43922 , n42121 );
and ( n43924 , n42066 , n42072 );
or ( n43925 , n43923 , n43924 );
buf ( n43926 , n43925 );
buf ( n43927 , n43926 );
xor ( n43928 , n43921 , n43927 );
buf ( n43929 , n43928 );
buf ( n43930 , n43929 );
xor ( n43931 , n43853 , n43930 );
xor ( n43932 , n42038 , n42044 );
and ( n43933 , n43932 , n42124 );
and ( n43934 , n42038 , n42044 );
or ( n43935 , n43933 , n43934 );
buf ( n43936 , n43935 );
buf ( n43937 , n43936 );
xor ( n43938 , n43931 , n43937 );
buf ( n43939 , n43938 );
buf ( n43940 , n43939 );
or ( n43941 , n43815 , n43940 );
buf ( n43942 , n43941 );
buf ( n43943 , n43942 );
buf ( n43944 , n43814 );
buf ( n43945 , n43939 );
nand ( n43946 , n43944 , n43945 );
buf ( n43947 , n43946 );
buf ( n43948 , n43947 );
nand ( n43949 , n43943 , n43948 );
buf ( n43950 , n43949 );
not ( n43951 , n43950 );
and ( n43952 , n43809 , n43951 );
not ( n43953 , n43809 );
and ( n43954 , n43953 , n43950 );
nor ( n43955 , n43952 , n43954 );
nand ( n43956 , n43955 , n2356 );
and ( n43957 , n43791 , n43794 , n43956 );
nor ( n43958 , n43499 , n43957 );
not ( n43959 , n43776 );
nor ( n43960 , n41950 , n43648 );
not ( n43961 , n43960 );
nand ( n43962 , n41970 , n41972 );
not ( n43963 , n43962 );
or ( n43964 , n43961 , n43963 );
or ( n43965 , n41948 , n43648 );
nand ( n43966 , n43965 , n43646 );
not ( n43967 , n43966 );
nand ( n43968 , n43964 , n43967 );
not ( n43969 , n43968 );
not ( n43970 , n455 );
xor ( n43971 , n43538 , n43631 );
and ( n43972 , n43971 , n43638 );
and ( n43973 , n43538 , n43631 );
or ( n43974 , n43972 , n43973 );
buf ( n43975 , n43974 );
xor ( n43976 , n43598 , n43623 );
and ( n43977 , n43976 , n43625 );
and ( n43978 , n43598 , n43623 );
or ( n43979 , n43977 , n43978 );
buf ( n43980 , n43979 );
buf ( n43981 , n43980 );
buf ( n43982 , n43584 );
not ( n43983 , n43982 );
buf ( n43984 , n43983 );
or ( n43985 , n43984 , n3145 );
not ( n43986 , n2704 );
nand ( n43987 , n43986 , n2978 );
nand ( n43988 , n43985 , n43987 );
buf ( n43989 , n43988 );
not ( n43990 , n43989 );
buf ( n43991 , n43990 );
buf ( n43992 , n43991 );
xor ( n43993 , n43549 , n43566 );
and ( n43994 , n43993 , n43592 );
and ( n43995 , n43549 , n43566 );
or ( n43996 , n43994 , n43995 );
buf ( n43997 , n43996 );
buf ( n43998 , n43997 );
xor ( n43999 , n43992 , n43998 );
and ( n44000 , n41849 , n41850 );
buf ( n44001 , n44000 );
buf ( n44002 , n44001 );
buf ( n44003 , n39149 );
not ( n44004 , n44003 );
buf ( n44005 , n43558 );
not ( n44006 , n44005 );
or ( n44007 , n44004 , n44006 );
buf ( n44008 , n489 );
buf ( n44009 , n39383 );
xor ( n44010 , n44008 , n44009 );
buf ( n44011 , n44010 );
buf ( n44012 , n44011 );
buf ( n44013 , n36508 );
nand ( n44014 , n44012 , n44013 );
buf ( n44015 , n44014 );
buf ( n44016 , n44015 );
nand ( n44017 , n44007 , n44016 );
buf ( n44018 , n44017 );
buf ( n44019 , n44018 );
xor ( n44020 , n44002 , n44019 );
buf ( n44021 , n3045 );
not ( n44022 , n44021 );
buf ( n44023 , n491 );
buf ( n44024 , n37462 );
and ( n44025 , n44023 , n44024 );
not ( n44026 , n44023 );
buf ( n44027 , n41902 );
and ( n44028 , n44026 , n44027 );
nor ( n44029 , n44025 , n44028 );
buf ( n44030 , n44029 );
buf ( n44031 , n44030 );
not ( n44032 , n44031 );
or ( n44033 , n44022 , n44032 );
buf ( n44034 , n43615 );
buf ( n44035 , n34465 );
nand ( n44036 , n44034 , n44035 );
buf ( n44037 , n44036 );
buf ( n44038 , n44037 );
nand ( n44039 , n44033 , n44038 );
buf ( n44040 , n44039 );
buf ( n44041 , n44040 );
xor ( n44042 , n44020 , n44041 );
buf ( n44043 , n44042 );
buf ( n44044 , n44043 );
xor ( n44045 , n43999 , n44044 );
buf ( n44046 , n44045 );
buf ( n44047 , n44046 );
xor ( n44048 , n43981 , n44047 );
xor ( n44049 , n43544 , n43595 );
and ( n44050 , n44049 , n43628 );
and ( n44051 , n43544 , n43595 );
or ( n44052 , n44050 , n44051 );
buf ( n44053 , n44052 );
buf ( n44054 , n44053 );
xor ( n44055 , n44048 , n44054 );
buf ( n44056 , n44055 );
or ( n44057 , n43975 , n44056 );
nand ( n44058 , n43975 , n44056 );
nand ( n44059 , n44057 , n44058 );
nor ( n44060 , n43970 , n44059 );
nand ( n44061 , n43969 , n44060 );
nand ( n44062 , n43968 , n44059 , n455 );
nor ( n44063 , n41814 , n43763 );
not ( n44064 , n44063 );
not ( n44065 , n41692 );
or ( n44066 , n44064 , n44065 );
not ( n44067 , n43756 );
not ( n44068 , n43761 );
or ( n44069 , n44067 , n44068 );
or ( n44070 , n41816 , n43763 );
nand ( n44071 , n44069 , n44070 );
not ( n44072 , n44071 );
nand ( n44073 , n44066 , n44072 );
xor ( n44074 , n43663 , n43747 );
and ( n44075 , n44074 , n43754 );
and ( n44076 , n43663 , n43747 );
or ( n44077 , n44075 , n44076 );
buf ( n44078 , n44077 );
xor ( n44079 , n43671 , n43684 );
and ( n44080 , n44079 , n41787 );
and ( n44081 , n43671 , n43684 );
or ( n44082 , n44080 , n44081 );
buf ( n44083 , n44082 );
buf ( n44084 , n4241 );
buf ( n44085 , n43729 );
and ( n44086 , n44084 , n44085 );
buf ( n44087 , n43732 );
buf ( n44088 , n493 );
and ( n44089 , n44087 , n44088 );
nor ( n44090 , n44086 , n44089 );
buf ( n44091 , n44090 );
buf ( n44092 , n44091 );
and ( n44093 , n41707 , n41708 );
buf ( n44094 , n44093 );
buf ( n44095 , n44094 );
buf ( n44096 , n43698 );
not ( n44097 , n44096 );
buf ( n44098 , n41718 );
not ( n44099 , n44098 );
or ( n44100 , n44097 , n44099 );
buf ( n44101 , n508 );
buf ( n44102 , n489 );
xnor ( n44103 , n44101 , n44102 );
buf ( n44104 , n44103 );
buf ( n44105 , n44104 );
not ( n44106 , n44105 );
buf ( n44107 , n37254 );
nand ( n44108 , n44106 , n44107 );
buf ( n44109 , n44108 );
buf ( n44110 , n44109 );
nand ( n44111 , n44100 , n44110 );
buf ( n44112 , n44111 );
buf ( n44113 , n44112 );
xor ( n44114 , n44095 , n44113 );
buf ( n44115 , n33964 );
buf ( n44116 , n43678 );
or ( n44117 , n44115 , n44116 );
buf ( n44118 , n41757 );
buf ( n44119 , n5167 );
buf ( n44120 , n506 );
and ( n44121 , n44119 , n44120 );
buf ( n44122 , n506 );
not ( n44123 , n44122 );
buf ( n44124 , n44123 );
buf ( n44125 , n44124 );
buf ( n44126 , n491 );
and ( n44127 , n44125 , n44126 );
nor ( n44128 , n44121 , n44127 );
buf ( n44129 , n44128 );
buf ( n44130 , n44129 );
or ( n44131 , n44118 , n44130 );
nand ( n44132 , n44117 , n44131 );
buf ( n44133 , n44132 );
buf ( n44134 , n44133 );
xor ( n44135 , n44114 , n44134 );
buf ( n44136 , n44135 );
buf ( n44137 , n44136 );
xor ( n44138 , n44092 , n44137 );
xor ( n44139 , n43705 , n43717 );
and ( n44140 , n44139 , n43741 );
and ( n44141 , n43705 , n43717 );
or ( n44142 , n44140 , n44141 );
buf ( n44143 , n44142 );
buf ( n44144 , n44143 );
xor ( n44145 , n44138 , n44144 );
buf ( n44146 , n44145 );
buf ( n44147 , n44146 );
xor ( n44148 , n44083 , n44147 );
xor ( n44149 , n43669 , n43687 );
and ( n44150 , n44149 , n43744 );
and ( n44151 , n43669 , n43687 );
or ( n44152 , n44150 , n44151 );
buf ( n44153 , n44152 );
buf ( n44154 , n44153 );
xor ( n44155 , n44148 , n44154 );
buf ( n44156 , n44155 );
or ( n44157 , n44078 , n44156 );
nand ( n44158 , n44078 , n44156 );
nand ( n44159 , n44157 , n44158 );
not ( n44160 , n44159 );
nor ( n44161 , n44160 , n455 );
and ( n44162 , n44073 , n44161 );
not ( n44163 , n44073 );
nor ( n44164 , n44159 , n455 );
and ( n44165 , n44163 , n44164 );
nor ( n44166 , n44162 , n44165 );
nand ( n44167 , n44061 , n44062 , n44166 );
not ( n44168 , n44167 );
or ( n44169 , n43959 , n44168 );
nand ( n44170 , n44169 , n43786 );
nor ( n44171 , n43514 , n44170 );
nand ( n44172 , n41083 , n44171 );
not ( n44173 , n44172 );
not ( n44174 , n44173 );
not ( n44175 , n41027 );
or ( n44176 , n44174 , n44175 );
not ( n44177 , n44171 );
not ( n44178 , n41089 );
or ( n44179 , n44177 , n44178 );
buf ( n44180 , n44170 );
not ( n44181 , n44180 );
buf ( n44182 , n44181 );
and ( n44183 , n44182 , n43505 );
nand ( n44184 , n44167 , n43776 );
not ( n44185 , n44184 );
nor ( n44186 , n43777 , n41985 );
not ( n44187 , n44186 );
or ( n44188 , n44185 , n44187 );
not ( n44189 , n44167 );
nand ( n44190 , n44189 , n43777 );
nand ( n44191 , n44188 , n44190 );
nor ( n44192 , n44183 , n44191 );
nand ( n44193 , n44179 , n44192 );
buf ( n44194 , n44193 );
not ( n44195 , n44194 );
buf ( n44196 , n44195 );
nand ( n44197 , n44176 , n44196 );
not ( n44198 , n44197 );
nand ( n44199 , n43960 , n44057 );
not ( n44200 , n44199 );
not ( n44201 , n44200 );
not ( n44202 , n43962 );
or ( n44203 , n44201 , n44202 );
not ( n44204 , n44057 );
not ( n44205 , n43966 );
or ( n44206 , n44204 , n44205 );
nand ( n44207 , n44206 , n44058 );
not ( n44208 , n44207 );
nand ( n44209 , n44203 , n44208 );
xor ( n44210 , n43981 , n44047 );
and ( n44211 , n44210 , n44054 );
and ( n44212 , n43981 , n44047 );
or ( n44213 , n44211 , n44212 );
buf ( n44214 , n44213 );
buf ( n44215 , n3146 );
buf ( n44216 , n3113 );
or ( n44217 , n44215 , n44216 );
buf ( n44218 , n493 );
nand ( n44219 , n44217 , n44218 );
buf ( n44220 , n44219 );
buf ( n44221 , n44220 );
and ( n44222 , n43555 , n43556 );
buf ( n44223 , n44222 );
buf ( n44224 , n44223 );
xor ( n44225 , n44221 , n44224 );
buf ( n44226 , n34465 );
not ( n44227 , n44226 );
buf ( n44228 , n44030 );
not ( n44229 , n44228 );
or ( n44230 , n44227 , n44229 );
buf ( n44231 , n491 );
buf ( n44232 , n41312 );
and ( n44233 , n44231 , n44232 );
not ( n44234 , n44231 );
buf ( n44235 , n42316 );
and ( n44236 , n44234 , n44235 );
nor ( n44237 , n44233 , n44236 );
buf ( n44238 , n44237 );
buf ( n44239 , n44238 );
buf ( n44240 , n3044 );
or ( n44241 , n44239 , n44240 );
nand ( n44242 , n44230 , n44241 );
buf ( n44243 , n44242 );
buf ( n44244 , n44243 );
xor ( n44245 , n44225 , n44244 );
buf ( n44246 , n44245 );
buf ( n44247 , n44246 );
buf ( n44248 , n36508 );
not ( n44249 , n44248 );
buf ( n44250 , n489 );
buf ( n44251 , n38414 );
xor ( n44252 , n44250 , n44251 );
buf ( n44253 , n44252 );
buf ( n44254 , n44253 );
not ( n44255 , n44254 );
or ( n44256 , n44249 , n44255 );
buf ( n44257 , n44011 );
not ( n44258 , n44257 );
buf ( n44259 , n44258 );
buf ( n44260 , n44259 );
buf ( n44261 , n39149 );
not ( n44262 , n44261 );
buf ( n44263 , n44262 );
buf ( n44264 , n44263 );
or ( n44265 , n44260 , n44264 );
nand ( n44266 , n44256 , n44265 );
buf ( n44267 , n44266 );
buf ( n44268 , n44267 );
buf ( n44269 , n43988 );
xor ( n44270 , n44268 , n44269 );
xor ( n44271 , n44002 , n44019 );
and ( n44272 , n44271 , n44041 );
and ( n44273 , n44002 , n44019 );
or ( n44274 , n44272 , n44273 );
buf ( n44275 , n44274 );
buf ( n44276 , n44275 );
xor ( n44277 , n44270 , n44276 );
buf ( n44278 , n44277 );
buf ( n44279 , n44278 );
xor ( n44280 , n44247 , n44279 );
xor ( n44281 , n43992 , n43998 );
and ( n44282 , n44281 , n44044 );
and ( n44283 , n43992 , n43998 );
or ( n44284 , n44282 , n44283 );
buf ( n44285 , n44284 );
buf ( n44286 , n44285 );
xor ( n44287 , n44280 , n44286 );
buf ( n44288 , n44287 );
or ( n44289 , n44214 , n44288 );
nand ( n44290 , n44214 , n44288 );
and ( n44291 , n44289 , n44290 );
nand ( n44292 , n44209 , n44291 );
not ( n44293 , n44292 );
nor ( n44294 , n44209 , n44291 );
nor ( n44295 , n44294 , n37874 );
not ( n44296 , n44295 );
or ( n44297 , n44293 , n44296 );
not ( n44298 , n41671 );
not ( n44299 , n41691 );
or ( n44300 , n44298 , n44299 );
nand ( n44301 , n44063 , n44157 );
not ( n44302 , n44301 );
nand ( n44303 , n44300 , n44302 );
not ( n44304 , n44303 );
xor ( n44305 , n44083 , n44147 );
and ( n44306 , n44305 , n44154 );
and ( n44307 , n44083 , n44147 );
or ( n44308 , n44306 , n44307 );
buf ( n44309 , n44308 );
buf ( n44310 , n33964 );
buf ( n44311 , n44129 );
or ( n44312 , n44310 , n44311 );
buf ( n44313 , n41757 );
buf ( n44314 , n5167 );
buf ( n44315 , n505 );
and ( n44316 , n44314 , n44315 );
buf ( n44317 , n43725 );
buf ( n44318 , n491 );
and ( n44319 , n44317 , n44318 );
nor ( n44320 , n44316 , n44319 );
buf ( n44321 , n44320 );
buf ( n44322 , n44321 );
or ( n44323 , n44313 , n44322 );
nand ( n44324 , n44312 , n44323 );
buf ( n44325 , n44324 );
buf ( n44326 , n44325 );
and ( n44327 , n43695 , n43696 );
buf ( n44328 , n44327 );
buf ( n44329 , n44328 );
xor ( n44330 , n44326 , n44329 );
buf ( n44331 , n41776 );
not ( n44332 , n44331 );
buf ( n44333 , n4242 );
not ( n44334 , n44333 );
or ( n44335 , n44332 , n44334 );
buf ( n44336 , n493 );
nand ( n44337 , n44335 , n44336 );
buf ( n44338 , n44337 );
buf ( n44339 , n44338 );
xor ( n44340 , n44330 , n44339 );
buf ( n44341 , n44340 );
buf ( n44342 , n44341 );
buf ( n44343 , n44091 );
not ( n44344 , n44343 );
buf ( n44345 , n44344 );
buf ( n44346 , n44345 );
buf ( n44347 , n41718 );
not ( n44348 , n44347 );
buf ( n44349 , n44348 );
or ( n44350 , n44349 , n44104 );
buf ( n44351 , n5539 );
buf ( n44352 , n507 );
and ( n44353 , n44351 , n44352 );
buf ( n44354 , n507 );
not ( n44355 , n44354 );
buf ( n44356 , n44355 );
buf ( n44357 , n44356 );
buf ( n44358 , n489 );
and ( n44359 , n44357 , n44358 );
nor ( n44360 , n44353 , n44359 );
buf ( n44361 , n44360 );
or ( n44362 , n37255 , n44361 );
nand ( n44363 , n44350 , n44362 );
buf ( n44364 , n44363 );
xor ( n44365 , n44346 , n44364 );
xor ( n44366 , n44095 , n44113 );
and ( n44367 , n44366 , n44134 );
and ( n44368 , n44095 , n44113 );
or ( n44369 , n44367 , n44368 );
buf ( n44370 , n44369 );
buf ( n44371 , n44370 );
xor ( n44372 , n44365 , n44371 );
buf ( n44373 , n44372 );
buf ( n44374 , n44373 );
xor ( n44375 , n44342 , n44374 );
xor ( n44376 , n44092 , n44137 );
and ( n44377 , n44376 , n44144 );
and ( n44378 , n44092 , n44137 );
or ( n44379 , n44377 , n44378 );
buf ( n44380 , n44379 );
buf ( n44381 , n44380 );
xor ( n44382 , n44375 , n44381 );
buf ( n44383 , n44382 );
or ( n44384 , n44309 , n44383 );
nand ( n44385 , n44309 , n44383 );
and ( n44386 , n44384 , n44385 );
not ( n44387 , n44386 );
not ( n44388 , n44157 );
not ( n44389 , n44071 );
or ( n44390 , n44388 , n44389 );
nand ( n44391 , n44390 , n44158 );
buf ( n44392 , n44391 );
nor ( n44393 , n44387 , n44392 );
nor ( n44394 , n44393 , n44392 );
not ( n44395 , n44394 );
or ( n44396 , n44304 , n44395 );
not ( n44397 , n44386 );
or ( n44398 , n44393 , n44397 );
nand ( n44399 , n44398 , n29519 );
nor ( n44400 , n44303 , n44397 );
nor ( n44401 , n44399 , n44400 );
nand ( n44402 , n44396 , n44401 );
nand ( n44403 , n44297 , n44402 );
nand ( n44404 , n44403 , n44189 );
nor ( n44405 , n44403 , n44189 );
buf ( n44406 , n44405 );
not ( n44407 , n44406 );
buf ( n44408 , n44407 );
and ( n44409 , n44404 , n44408 );
and ( n44410 , n44409 , n454 );
nand ( n44411 , n44198 , n44410 );
nor ( n44412 , n2618 , n44409 );
nand ( n44413 , n44197 , n44412 );
not ( n44414 , n454 );
buf ( n44415 , n528 );
buf ( n44416 , n537 );
and ( n44417 , n44415 , n44416 );
buf ( n44418 , n44417 );
buf ( n44419 , n44418 );
buf ( n44420 , n525 );
buf ( n44421 , n540 );
and ( n44422 , n44420 , n44421 );
buf ( n44423 , n44422 );
buf ( n44424 , n44423 );
xor ( n44425 , n44419 , n44424 );
buf ( n44426 , n523 );
buf ( n44427 , n542 );
and ( n44428 , n44426 , n44427 );
buf ( n44429 , n44428 );
buf ( n44430 , n44429 );
xor ( n44431 , n44425 , n44430 );
buf ( n44432 , n44431 );
buf ( n44433 , n44432 );
buf ( n44434 , n526 );
buf ( n44435 , n539 );
and ( n44436 , n44434 , n44435 );
buf ( n44437 , n44436 );
buf ( n44438 , n44437 );
buf ( n44439 , n527 );
buf ( n44440 , n538 );
and ( n44441 , n44439 , n44440 );
buf ( n44442 , n44441 );
buf ( n44443 , n44442 );
xor ( n44444 , n44438 , n44443 );
xor ( n44445 , n43877 , n43882 );
and ( n44446 , n44445 , n43888 );
and ( n44447 , n43877 , n43882 );
or ( n44448 , n44446 , n44447 );
buf ( n44449 , n44448 );
buf ( n44450 , n44449 );
xor ( n44451 , n44444 , n44450 );
buf ( n44452 , n44451 );
buf ( n44453 , n44452 );
xor ( n44454 , n44433 , n44453 );
xor ( n44455 , n43834 , n43840 );
and ( n44456 , n44455 , n43847 );
and ( n44457 , n43834 , n43840 );
or ( n44458 , n44456 , n44457 );
buf ( n44459 , n44458 );
buf ( n44460 , n44459 );
xor ( n44461 , n44454 , n44460 );
buf ( n44462 , n44461 );
buf ( n44463 , n44462 );
xor ( n44464 , n43858 , n43863 );
and ( n44465 , n44464 , n43869 );
and ( n44466 , n43858 , n43863 );
or ( n44467 , n44465 , n44466 );
buf ( n44468 , n44467 );
buf ( n44469 , n44468 );
xor ( n44470 , n43897 , n43902 );
and ( n44471 , n44470 , n43908 );
and ( n44472 , n43897 , n43902 );
or ( n44473 , n44471 , n44472 );
buf ( n44474 , n44473 );
buf ( n44475 , n44474 );
xor ( n44476 , n44469 , n44475 );
buf ( n44477 , n521 );
buf ( n44478 , n544 );
and ( n44479 , n44477 , n44478 );
buf ( n44480 , n44479 );
buf ( n44481 , n44480 );
buf ( n44482 , n522 );
buf ( n44483 , n543 );
and ( n44484 , n44482 , n44483 );
buf ( n44485 , n44484 );
buf ( n44486 , n44485 );
xor ( n44487 , n44481 , n44486 );
buf ( n44488 , n524 );
buf ( n44489 , n541 );
and ( n44490 , n44488 , n44489 );
buf ( n44491 , n44490 );
buf ( n44492 , n44491 );
xor ( n44493 , n44487 , n44492 );
buf ( n44494 , n44493 );
buf ( n44495 , n44494 );
xor ( n44496 , n44476 , n44495 );
buf ( n44497 , n44496 );
buf ( n44498 , n44497 );
xor ( n44499 , n43872 , n43891 );
and ( n44500 , n44499 , n43911 );
and ( n44501 , n43872 , n43891 );
or ( n44502 , n44500 , n44501 );
buf ( n44503 , n44502 );
buf ( n44504 , n44503 );
xor ( n44505 , n44498 , n44504 );
xor ( n44506 , n43821 , n43827 );
and ( n44507 , n44506 , n43850 );
and ( n44508 , n43821 , n43827 );
or ( n44509 , n44507 , n44508 );
buf ( n44510 , n44509 );
buf ( n44511 , n44510 );
xor ( n44512 , n44505 , n44511 );
buf ( n44513 , n44512 );
buf ( n44514 , n44513 );
xor ( n44515 , n44463 , n44514 );
xor ( n44516 , n43914 , n43920 );
and ( n44517 , n44516 , n43927 );
and ( n44518 , n43914 , n43920 );
or ( n44519 , n44517 , n44518 );
buf ( n44520 , n44519 );
buf ( n44521 , n44520 );
and ( n44522 , n44515 , n44521 );
and ( n44523 , n44463 , n44514 );
or ( n44524 , n44522 , n44523 );
buf ( n44525 , n44524 );
buf ( n44526 , n44525 );
buf ( n44527 , n525 );
buf ( n44528 , n539 );
and ( n44529 , n44527 , n44528 );
buf ( n44530 , n44529 );
buf ( n44531 , n44530 );
buf ( n44532 , n523 );
buf ( n44533 , n541 );
and ( n44534 , n44532 , n44533 );
buf ( n44535 , n44534 );
buf ( n44536 , n44535 );
xor ( n44537 , n44531 , n44536 );
buf ( n44538 , n526 );
buf ( n44539 , n538 );
and ( n44540 , n44538 , n44539 );
buf ( n44541 , n44540 );
buf ( n44542 , n44541 );
xor ( n44543 , n44537 , n44542 );
buf ( n44544 , n44543 );
buf ( n44545 , n44544 );
buf ( n44546 , n521 );
buf ( n44547 , n543 );
and ( n44548 , n44546 , n44547 );
buf ( n44549 , n44548 );
buf ( n44550 , n44549 );
buf ( n44551 , n522 );
buf ( n44552 , n542 );
and ( n44553 , n44551 , n44552 );
buf ( n44554 , n44553 );
buf ( n44555 , n44554 );
xor ( n44556 , n44550 , n44555 );
buf ( n44557 , n524 );
buf ( n44558 , n540 );
and ( n44559 , n44557 , n44558 );
buf ( n44560 , n44559 );
buf ( n44561 , n44560 );
xor ( n44562 , n44556 , n44561 );
buf ( n44563 , n44562 );
buf ( n44564 , n44563 );
xor ( n44565 , n44545 , n44564 );
xor ( n44566 , n44438 , n44443 );
and ( n44567 , n44566 , n44450 );
and ( n44568 , n44438 , n44443 );
or ( n44569 , n44567 , n44568 );
buf ( n44570 , n44569 );
buf ( n44571 , n44570 );
xor ( n44572 , n44565 , n44571 );
buf ( n44573 , n44572 );
buf ( n44574 , n44573 );
buf ( n44575 , n527 );
buf ( n44576 , n537 );
and ( n44577 , n44575 , n44576 );
buf ( n44578 , n44577 );
buf ( n44579 , n44578 );
xor ( n44580 , n44481 , n44486 );
and ( n44581 , n44580 , n44492 );
and ( n44582 , n44481 , n44486 );
or ( n44583 , n44581 , n44582 );
buf ( n44584 , n44583 );
buf ( n44585 , n44584 );
xor ( n44586 , n44579 , n44585 );
xor ( n44587 , n44419 , n44424 );
and ( n44588 , n44587 , n44430 );
and ( n44589 , n44419 , n44424 );
or ( n44590 , n44588 , n44589 );
buf ( n44591 , n44590 );
buf ( n44592 , n44591 );
xor ( n44593 , n44586 , n44592 );
buf ( n44594 , n44593 );
buf ( n44595 , n44594 );
xor ( n44596 , n44469 , n44475 );
and ( n44597 , n44596 , n44495 );
and ( n44598 , n44469 , n44475 );
or ( n44599 , n44597 , n44598 );
buf ( n44600 , n44599 );
buf ( n44601 , n44600 );
xor ( n44602 , n44595 , n44601 );
xor ( n44603 , n44433 , n44453 );
and ( n44604 , n44603 , n44460 );
and ( n44605 , n44433 , n44453 );
or ( n44606 , n44604 , n44605 );
buf ( n44607 , n44606 );
buf ( n44608 , n44607 );
xor ( n44609 , n44602 , n44608 );
buf ( n44610 , n44609 );
buf ( n44611 , n44610 );
xor ( n44612 , n44574 , n44611 );
xor ( n44613 , n44498 , n44504 );
and ( n44614 , n44613 , n44511 );
and ( n44615 , n44498 , n44504 );
or ( n44616 , n44614 , n44615 );
buf ( n44617 , n44616 );
buf ( n44618 , n44617 );
xor ( n44619 , n44612 , n44618 );
buf ( n44620 , n44619 );
buf ( n44621 , n44620 );
and ( n44622 , n44526 , n44621 );
buf ( n44623 , n44622 );
buf ( n44624 , n44623 );
not ( n44625 , n44624 );
buf ( n44626 , n44625 );
buf ( n44627 , n44626 );
buf ( n44628 , n44525 );
buf ( n44629 , n44620 );
or ( n44630 , n44628 , n44629 );
buf ( n44631 , n44630 );
buf ( n44632 , n44631 );
nand ( n44633 , n44627 , n44632 );
buf ( n44634 , n44633 );
buf ( n44635 , n44634 );
not ( n44636 , n44635 );
buf ( n44637 , n43800 );
buf ( n44638 , n43942 );
xor ( n44639 , n43853 , n43930 );
and ( n44640 , n44639 , n43937 );
and ( n44641 , n43853 , n43930 );
or ( n44642 , n44640 , n44641 );
buf ( n44643 , n44642 );
buf ( n44644 , n44643 );
xor ( n44645 , n44463 , n44514 );
xor ( n44646 , n44645 , n44521 );
buf ( n44647 , n44646 );
buf ( n44648 , n44647 );
or ( n44649 , n44644 , n44648 );
buf ( n44650 , n44649 );
buf ( n44651 , n44650 );
nand ( n44652 , n44638 , n44651 );
buf ( n44653 , n44652 );
buf ( n44654 , n44653 );
nor ( n44655 , n44637 , n44654 );
buf ( n44656 , n44655 );
not ( n44657 , n44656 );
not ( n44658 , n41640 );
or ( n44659 , n44657 , n44658 );
or ( n44660 , n44643 , n44647 );
not ( n44661 , n43942 );
not ( n44662 , n43806 );
or ( n44663 , n44661 , n44662 );
nand ( n44664 , n44663 , n43947 );
nand ( n44665 , n44660 , n44664 );
nand ( n44666 , n44647 , n44643 );
nand ( n44667 , n44665 , n44666 );
not ( n44668 , n44667 );
nand ( n44669 , n44659 , n44668 );
buf ( n44670 , n44669 );
not ( n44671 , n44670 );
or ( n44672 , n44636 , n44671 );
buf ( n44673 , n44634 );
buf ( n44674 , n44669 );
or ( n44675 , n44673 , n44674 );
nand ( n44676 , n44672 , n44675 );
buf ( n44677 , n44676 );
nand ( n44678 , n44414 , n44677 );
nand ( n44679 , n44411 , n44413 , n44678 );
not ( n44680 , n2356 );
buf ( n44681 , n43942 );
not ( n44682 , n44681 );
buf ( n44683 , n43803 );
not ( n44684 , n44683 );
or ( n44685 , n44682 , n44684 );
buf ( n44686 , n43942 );
not ( n44687 , n44686 );
buf ( n44688 , n43806 );
not ( n44689 , n44688 );
or ( n44690 , n44687 , n44689 );
buf ( n44691 , n43947 );
nand ( n44692 , n44690 , n44691 );
buf ( n44693 , n44692 );
buf ( n44694 , n44693 );
not ( n44695 , n44694 );
buf ( n44696 , n44695 );
buf ( n44697 , n44696 );
nand ( n44698 , n44685 , n44697 );
buf ( n44699 , n44698 );
buf ( n44700 , n44699 );
buf ( n44701 , n44650 );
buf ( n44702 , n44666 );
nand ( n44703 , n44701 , n44702 );
buf ( n44704 , n44703 );
buf ( n44705 , n44704 );
xnor ( n44706 , n44700 , n44705 );
buf ( n44707 , n44706 );
not ( n44708 , n44707 );
or ( n44709 , n44680 , n44708 );
nand ( n44710 , n43515 , n43787 );
nor ( n44711 , n44710 , n41658 );
not ( n44712 , n44711 );
not ( n44713 , n37966 );
or ( n44714 , n44712 , n44713 );
not ( n44715 , n44710 );
not ( n44716 , n41090 );
and ( n44717 , n44715 , n44716 );
not ( n44718 , n43787 );
not ( n44719 , n43505 );
or ( n44720 , n44718 , n44719 );
not ( n44721 , n43778 );
nand ( n44722 , n44720 , n44721 );
nor ( n44723 , n44717 , n44722 );
nand ( n44724 , n44714 , n44723 );
not ( n44725 , n44724 );
buf ( n44726 , n44190 );
buf ( n44727 , n44726 );
buf ( n44728 , n44727 );
buf ( n44729 , n44184 );
nand ( n44730 , n44728 , n44729 );
not ( n44731 , n44730 );
nand ( n44732 , n44731 , n454 );
not ( n44733 , n44732 );
and ( n44734 , n44725 , n44733 );
nor ( n44735 , n44731 , n2618 );
and ( n44736 , n44724 , n44735 );
nor ( n44737 , n44734 , n44736 );
nand ( n44738 , n44709 , n44737 );
nand ( n44739 , n43958 , n44679 , n44738 );
not ( n44740 , n44739 );
nand ( n44741 , n44740 , n41654 );
buf ( n44742 , n6887 );
not ( n44743 , n44742 );
not ( n44744 , n7042 );
or ( n44745 , n44743 , n44744 );
nand ( n44746 , n44745 , n7047 );
buf ( n44747 , n6915 );
and ( n44748 , n44746 , n44747 );
not ( n44749 , n44746 );
and ( n44750 , n44749 , n7046 );
nor ( n44751 , n44748 , n44750 );
nand ( n44752 , n7036 , n6980 );
not ( n44753 , n7033 );
and ( n44754 , n44752 , n44753 );
not ( n44755 , n44752 );
and ( n44756 , n44755 , n7033 );
nor ( n44757 , n44754 , n44756 );
and ( n44758 , n2358 , n472 );
not ( n44759 , n2358 );
and ( n44760 , n44759 , n7025 );
nor ( n44761 , n44758 , n44760 );
xor ( n44762 , n44247 , n44279 );
and ( n44763 , n44762 , n44286 );
and ( n44764 , n44247 , n44279 );
or ( n44765 , n44763 , n44764 );
buf ( n44766 , n44765 );
xor ( n44767 , n44221 , n44224 );
and ( n44768 , n44767 , n44244 );
and ( n44769 , n44221 , n44224 );
or ( n44770 , n44768 , n44769 );
buf ( n44771 , n44770 );
buf ( n44772 , n44771 );
buf ( n44773 , n44238 );
not ( n44774 , n44773 );
buf ( n44775 , n44774 );
buf ( n44776 , n44775 );
buf ( n44777 , n34465 );
and ( n44778 , n44776 , n44777 );
buf ( n44779 , n3045 );
buf ( n44780 , n491 );
and ( n44781 , n44779 , n44780 );
nor ( n44782 , n44778 , n44781 );
buf ( n44783 , n44782 );
buf ( n44784 , n44783 );
and ( n44785 , n44008 , n44009 );
buf ( n44786 , n44785 );
buf ( n44787 , n44786 );
xor ( n44788 , n44784 , n44787 );
buf ( n44789 , n39149 );
not ( n44790 , n44789 );
buf ( n44791 , n44253 );
not ( n44792 , n44791 );
or ( n44793 , n44790 , n44792 );
buf ( n44794 , n37462 );
buf ( n44795 , n489 );
xnor ( n44796 , n44794 , n44795 );
buf ( n44797 , n44796 );
buf ( n44798 , n44797 );
buf ( n44799 , n36508 );
not ( n44800 , n44799 );
buf ( n44801 , n44800 );
buf ( n44802 , n44801 );
or ( n44803 , n44798 , n44802 );
nand ( n44804 , n44793 , n44803 );
buf ( n44805 , n44804 );
buf ( n44806 , n44805 );
xor ( n44807 , n44788 , n44806 );
buf ( n44808 , n44807 );
buf ( n44809 , n44808 );
xor ( n44810 , n44268 , n44269 );
and ( n44811 , n44810 , n44276 );
and ( n44812 , n44268 , n44269 );
or ( n44813 , n44811 , n44812 );
buf ( n44814 , n44813 );
buf ( n44815 , n44814 );
xor ( n44816 , n44772 , n44809 );
xor ( n44817 , n44816 , n44815 );
buf ( n44818 , n44817 );
xor ( n44819 , n44772 , n44809 );
and ( n44820 , n44819 , n44815 );
and ( n44821 , n44772 , n44809 );
or ( n44822 , n44820 , n44821 );
buf ( n44823 , n44822 );
buf ( n44824 , n44783 );
not ( n44825 , n44824 );
buf ( n44826 , n44825 );
buf ( n44827 , n44826 );
xor ( n44828 , n44784 , n44787 );
and ( n44829 , n44828 , n44806 );
and ( n44830 , n44784 , n44787 );
or ( n44831 , n44829 , n44830 );
buf ( n44832 , n44831 );
buf ( n44833 , n44832 );
buf ( n44834 , n34465 );
buf ( n44835 , n3045 );
or ( n44836 , n44834 , n44835 );
buf ( n44837 , n491 );
nand ( n44838 , n44836 , n44837 );
buf ( n44839 , n44838 );
buf ( n44840 , n44839 );
and ( n44841 , n44250 , n44251 );
buf ( n44842 , n44841 );
buf ( n44843 , n44842 );
xor ( n44844 , n44840 , n44843 );
buf ( n44845 , n36508 );
not ( n44846 , n44845 );
buf ( n44847 , n489 );
buf ( n44848 , n41311 );
and ( n44849 , n44847 , n44848 );
not ( n44850 , n44847 );
buf ( n44851 , n42316 );
and ( n44852 , n44850 , n44851 );
nor ( n44853 , n44849 , n44852 );
buf ( n44854 , n44853 );
buf ( n44855 , n44854 );
not ( n44856 , n44855 );
buf ( n44857 , n44856 );
buf ( n44858 , n44857 );
not ( n44859 , n44858 );
or ( n44860 , n44846 , n44859 );
buf ( n44861 , n44797 );
buf ( n44862 , n44263 );
or ( n44863 , n44861 , n44862 );
nand ( n44864 , n44860 , n44863 );
buf ( n44865 , n44864 );
buf ( n44866 , n44865 );
xor ( n44867 , n44844 , n44866 );
buf ( n44868 , n44867 );
buf ( n44869 , n44868 );
xor ( n44870 , n44827 , n44833 );
xor ( n44871 , n44870 , n44869 );
buf ( n44872 , n44871 );
xor ( n44873 , n44827 , n44833 );
and ( n44874 , n44873 , n44869 );
and ( n44875 , n44827 , n44833 );
or ( n44876 , n44874 , n44875 );
buf ( n44877 , n44876 );
buf ( n44878 , n44854 );
buf ( n44879 , n44263 );
or ( n44880 , n44878 , n44879 );
buf ( n44881 , n44801 );
buf ( n44882 , n5437 );
or ( n44883 , n44881 , n44882 );
nand ( n44884 , n44880 , n44883 );
buf ( n44885 , n44884 );
buf ( n44886 , n44885 );
buf ( n44887 , n42328 );
buf ( n44888 , n489 );
nand ( n44889 , n44887 , n44888 );
buf ( n44890 , n44889 );
buf ( n44891 , n44890 );
xor ( n44892 , n44840 , n44843 );
and ( n44893 , n44892 , n44866 );
and ( n44894 , n44840 , n44843 );
or ( n44895 , n44893 , n44894 );
buf ( n44896 , n44895 );
buf ( n44897 , n44896 );
xor ( n44898 , n44886 , n44891 );
xor ( n44899 , n44898 , n44897 );
buf ( n44900 , n44899 );
xor ( n44901 , n44886 , n44891 );
and ( n44902 , n44901 , n44897 );
and ( n44903 , n44886 , n44891 );
or ( n44904 , n44902 , n44903 );
buf ( n44905 , n44904 );
buf ( n44906 , n44890 );
buf ( n44907 , n43035 );
buf ( n44908 , n489 );
nand ( n44909 , n44907 , n44908 );
buf ( n44910 , n44909 );
buf ( n44911 , n44910 );
not ( n44912 , n44911 );
buf ( n44913 , n39149 );
buf ( n44914 , n36508 );
or ( n44915 , n44913 , n44914 );
buf ( n44916 , n489 );
nand ( n44917 , n44915 , n44916 );
buf ( n44918 , n44917 );
buf ( n44919 , n44918 );
not ( n44920 , n44919 );
or ( n44921 , n44912 , n44920 );
buf ( n44922 , n44918 );
buf ( n44923 , n44910 );
or ( n44924 , n44922 , n44923 );
nand ( n44925 , n44921 , n44924 );
buf ( n44926 , n44925 );
buf ( n44927 , n44926 );
buf ( n44928 , n44926 );
buf ( n44929 , n44890 );
not ( n44930 , n44906 );
not ( n44931 , n44927 );
or ( n44932 , n44930 , n44931 );
or ( n44933 , n44928 , n44929 );
nand ( n44934 , n44932 , n44933 );
buf ( n44935 , n44934 );
xor ( n44936 , n44342 , n44374 );
and ( n44937 , n44936 , n44381 );
and ( n44938 , n44342 , n44374 );
or ( n44939 , n44937 , n44938 );
buf ( n44940 , n44939 );
xor ( n44941 , n44326 , n44329 );
and ( n44942 , n44941 , n44339 );
and ( n44943 , n44326 , n44329 );
or ( n44944 , n44942 , n44943 );
buf ( n44945 , n44944 );
buf ( n44946 , n44945 );
buf ( n44947 , n44349 );
buf ( n44948 , n44361 );
or ( n44949 , n44947 , n44948 );
buf ( n44950 , n37255 );
buf ( n44951 , n5539 );
buf ( n44952 , n506 );
and ( n44953 , n44951 , n44952 );
buf ( n44954 , n44124 );
buf ( n44955 , n489 );
and ( n44956 , n44954 , n44955 );
nor ( n44957 , n44953 , n44956 );
buf ( n44958 , n44957 );
buf ( n44959 , n44958 );
or ( n44960 , n44950 , n44959 );
nand ( n44961 , n44949 , n44960 );
buf ( n44962 , n44961 );
buf ( n44963 , n44962 );
buf ( n44964 , n5539 );
buf ( n44965 , n33049 );
nor ( n44966 , n44964 , n44965 );
buf ( n44967 , n44966 );
buf ( n44968 , n44967 );
xor ( n44969 , n44963 , n44968 );
buf ( n44970 , n33964 );
not ( n44971 , n44970 );
buf ( n44972 , n44321 );
not ( n44973 , n44972 );
and ( n44974 , n44971 , n44973 );
buf ( n44975 , n33973 );
buf ( n44976 , n491 );
and ( n44977 , n44975 , n44976 );
nor ( n44978 , n44974 , n44977 );
buf ( n44979 , n44978 );
buf ( n44980 , n44979 );
xor ( n44981 , n44969 , n44980 );
buf ( n44982 , n44981 );
buf ( n44983 , n44982 );
xor ( n44984 , n44346 , n44364 );
and ( n44985 , n44984 , n44371 );
and ( n44986 , n44346 , n44364 );
or ( n44987 , n44985 , n44986 );
buf ( n44988 , n44987 );
buf ( n44989 , n44988 );
xor ( n44990 , n44946 , n44983 );
xor ( n44991 , n44990 , n44989 );
buf ( n44992 , n44991 );
xor ( n44993 , n44946 , n44983 );
and ( n44994 , n44993 , n44989 );
and ( n44995 , n44946 , n44983 );
or ( n44996 , n44994 , n44995 );
buf ( n44997 , n44996 );
xor ( n44998 , n44963 , n44968 );
and ( n44999 , n44998 , n44980 );
and ( n45000 , n44963 , n44968 );
or ( n45001 , n44999 , n45000 );
buf ( n45002 , n45001 );
buf ( n45003 , n45002 );
buf ( n45004 , n44979 );
not ( n45005 , n45004 );
buf ( n45006 , n45005 );
buf ( n45007 , n45006 );
buf ( n45008 , n33967 );
buf ( n45009 , n33973 );
or ( n45010 , n45008 , n45009 );
buf ( n45011 , n491 );
nand ( n45012 , n45010 , n45011 );
buf ( n45013 , n45012 );
buf ( n45014 , n45013 );
buf ( n45015 , n5539 );
buf ( n45016 , n44356 );
nor ( n45017 , n45015 , n45016 );
buf ( n45018 , n45017 );
buf ( n45019 , n45018 );
xor ( n45020 , n45014 , n45019 );
buf ( n45021 , n44349 );
buf ( n45022 , n44958 );
or ( n45023 , n45021 , n45022 );
buf ( n45024 , n37255 );
buf ( n45025 , n5539 );
buf ( n45026 , n505 );
and ( n45027 , n45025 , n45026 );
buf ( n45028 , n43725 );
buf ( n45029 , n489 );
and ( n45030 , n45028 , n45029 );
nor ( n45031 , n45027 , n45030 );
buf ( n45032 , n45031 );
buf ( n45033 , n45032 );
or ( n45034 , n45024 , n45033 );
nand ( n45035 , n45023 , n45034 );
buf ( n45036 , n45035 );
buf ( n45037 , n45036 );
xor ( n45038 , n45020 , n45037 );
buf ( n45039 , n45038 );
buf ( n45040 , n45039 );
xor ( n45041 , n45003 , n45007 );
xor ( n45042 , n45041 , n45040 );
buf ( n45043 , n45042 );
xor ( n45044 , n45003 , n45007 );
and ( n45045 , n45044 , n45040 );
and ( n45046 , n45003 , n45007 );
or ( n45047 , n45045 , n45046 );
buf ( n45048 , n45047 );
buf ( n45049 , n44349 );
buf ( n45050 , n45032 );
or ( n45051 , n45049 , n45050 );
buf ( n45052 , n37255 );
buf ( n45053 , n5539 );
or ( n45054 , n45052 , n45053 );
nand ( n45055 , n45051 , n45054 );
buf ( n45056 , n45055 );
buf ( n45057 , n45056 );
buf ( n45058 , n506 );
buf ( n45059 , n489 );
nand ( n45060 , n45058 , n45059 );
buf ( n45061 , n45060 );
buf ( n45062 , n45061 );
xor ( n45063 , n45014 , n45019 );
and ( n45064 , n45063 , n45037 );
and ( n45065 , n45014 , n45019 );
or ( n45066 , n45064 , n45065 );
buf ( n45067 , n45066 );
buf ( n45068 , n45067 );
xor ( n45069 , n45057 , n45062 );
xor ( n45070 , n45069 , n45068 );
buf ( n45071 , n45070 );
xor ( n45072 , n45057 , n45062 );
and ( n45073 , n45072 , n45068 );
and ( n45074 , n45057 , n45062 );
or ( n45075 , n45073 , n45074 );
buf ( n45076 , n45075 );
buf ( n45077 , n45061 );
buf ( n45078 , n505 );
buf ( n45079 , n489 );
nand ( n45080 , n45078 , n45079 );
buf ( n45081 , n45080 );
buf ( n45082 , n45081 );
not ( n45083 , n45082 );
buf ( n45084 , n41718 );
buf ( n45085 , n37254 );
or ( n45086 , n45084 , n45085 );
buf ( n45087 , n489 );
nand ( n45088 , n45086 , n45087 );
buf ( n45089 , n45088 );
buf ( n45090 , n45089 );
not ( n45091 , n45090 );
or ( n45092 , n45083 , n45091 );
buf ( n45093 , n45089 );
buf ( n45094 , n45081 );
or ( n45095 , n45093 , n45094 );
nand ( n45096 , n45092 , n45095 );
buf ( n45097 , n45096 );
buf ( n45098 , n45097 );
buf ( n45099 , n45097 );
buf ( n45100 , n45061 );
not ( n45101 , n45077 );
not ( n45102 , n45098 );
or ( n45103 , n45101 , n45102 );
or ( n45104 , n45099 , n45100 );
nand ( n45105 , n45103 , n45104 );
buf ( n45106 , n45105 );
xor ( n45107 , n44550 , n44555 );
and ( n45108 , n45107 , n44561 );
and ( n45109 , n44550 , n44555 );
or ( n45110 , n45108 , n45109 );
buf ( n45111 , n45110 );
xor ( n45112 , n44531 , n44536 );
and ( n45113 , n45112 , n44542 );
and ( n45114 , n44531 , n44536 );
or ( n45115 , n45113 , n45114 );
buf ( n45116 , n45115 );
xor ( n45117 , n44579 , n44585 );
and ( n45118 , n45117 , n44592 );
and ( n45119 , n44579 , n44585 );
or ( n45120 , n45118 , n45119 );
buf ( n45121 , n45120 );
xor ( n45122 , n44545 , n44564 );
and ( n45123 , n45122 , n44571 );
and ( n45124 , n44545 , n44564 );
or ( n45125 , n45123 , n45124 );
buf ( n45126 , n45125 );
xor ( n45127 , n44595 , n44601 );
and ( n45128 , n45127 , n44608 );
and ( n45129 , n44595 , n44601 );
or ( n45130 , n45128 , n45129 );
buf ( n45131 , n45130 );
xor ( n45132 , n44574 , n44611 );
and ( n45133 , n45132 , n44618 );
and ( n45134 , n44574 , n44611 );
or ( n45135 , n45133 , n45134 );
buf ( n45136 , n45135 );
buf ( n45137 , n521 );
buf ( n45138 , n542 );
and ( n45139 , n45137 , n45138 );
buf ( n45140 , n45139 );
buf ( n45141 , n45140 );
buf ( n45142 , n522 );
buf ( n45143 , n541 );
and ( n45144 , n45142 , n45143 );
buf ( n45145 , n45144 );
buf ( n45146 , n45145 );
buf ( n45147 , n524 );
buf ( n45148 , n539 );
and ( n45149 , n45147 , n45148 );
buf ( n45150 , n45149 );
buf ( n45151 , n45150 );
xor ( n45152 , n45141 , n45146 );
xor ( n45153 , n45152 , n45151 );
buf ( n45154 , n45153 );
xor ( n45155 , n45141 , n45146 );
and ( n45156 , n45155 , n45151 );
and ( n45157 , n45141 , n45146 );
or ( n45158 , n45156 , n45157 );
buf ( n45159 , n45158 );
buf ( n45160 , n525 );
buf ( n45161 , n538 );
and ( n45162 , n45160 , n45161 );
buf ( n45163 , n45162 );
buf ( n45164 , n45163 );
buf ( n45165 , n523 );
buf ( n45166 , n540 );
and ( n45167 , n45165 , n45166 );
buf ( n45168 , n45167 );
buf ( n45169 , n45168 );
buf ( n45170 , n526 );
buf ( n45171 , n537 );
and ( n45172 , n45170 , n45171 );
buf ( n45173 , n45172 );
buf ( n45174 , n45173 );
xor ( n45175 , n45164 , n45169 );
xor ( n45176 , n45175 , n45174 );
buf ( n45177 , n45176 );
xor ( n45178 , n45164 , n45169 );
and ( n45179 , n45178 , n45174 );
and ( n45180 , n45164 , n45169 );
or ( n45181 , n45179 , n45180 );
buf ( n45182 , n45181 );
buf ( n45183 , n45116 );
buf ( n45184 , n45111 );
buf ( n45185 , n45154 );
xor ( n45186 , n45183 , n45184 );
xor ( n45187 , n45186 , n45185 );
buf ( n45188 , n45187 );
xor ( n45189 , n45183 , n45184 );
and ( n45190 , n45189 , n45185 );
and ( n45191 , n45183 , n45184 );
or ( n45192 , n45190 , n45191 );
buf ( n45193 , n45192 );
buf ( n45194 , n45177 );
buf ( n45195 , n45121 );
buf ( n45196 , n45188 );
xor ( n45197 , n45194 , n45195 );
xor ( n45198 , n45197 , n45196 );
buf ( n45199 , n45198 );
xor ( n45200 , n45194 , n45195 );
and ( n45201 , n45200 , n45196 );
and ( n45202 , n45194 , n45195 );
or ( n45203 , n45201 , n45202 );
buf ( n45204 , n45203 );
buf ( n45205 , n45126 );
buf ( n45206 , n45199 );
buf ( n45207 , n45131 );
xor ( n45208 , n45205 , n45206 );
xor ( n45209 , n45208 , n45207 );
buf ( n45210 , n45209 );
xor ( n45211 , n45205 , n45206 );
and ( n45212 , n45211 , n45207 );
and ( n45213 , n45205 , n45206 );
or ( n45214 , n45212 , n45213 );
buf ( n45215 , n45214 );
buf ( n45216 , n521 );
buf ( n45217 , n541 );
and ( n45218 , n45216 , n45217 );
buf ( n45219 , n45218 );
buf ( n45220 , n45219 );
buf ( n45221 , n522 );
buf ( n45222 , n540 );
and ( n45223 , n45221 , n45222 );
buf ( n45224 , n45223 );
buf ( n45225 , n45224 );
buf ( n45226 , n524 );
buf ( n45227 , n538 );
and ( n45228 , n45226 , n45227 );
buf ( n45229 , n45228 );
buf ( n45230 , n45229 );
xor ( n45231 , n45220 , n45225 );
xor ( n45232 , n45231 , n45230 );
buf ( n45233 , n45232 );
xor ( n45234 , n45220 , n45225 );
and ( n45235 , n45234 , n45230 );
and ( n45236 , n45220 , n45225 );
or ( n45237 , n45235 , n45236 );
buf ( n45238 , n45237 );
buf ( n45239 , n525 );
buf ( n45240 , n537 );
and ( n45241 , n45239 , n45240 );
buf ( n45242 , n45241 );
buf ( n45243 , n45242 );
buf ( n45244 , n523 );
buf ( n45245 , n539 );
and ( n45246 , n45244 , n45245 );
buf ( n45247 , n45246 );
buf ( n45248 , n45247 );
buf ( n45249 , n45182 );
xor ( n45250 , n45243 , n45248 );
xor ( n45251 , n45250 , n45249 );
buf ( n45252 , n45251 );
xor ( n45253 , n45243 , n45248 );
and ( n45254 , n45253 , n45249 );
and ( n45255 , n45243 , n45248 );
or ( n45256 , n45254 , n45255 );
buf ( n45257 , n45256 );
buf ( n45258 , n45159 );
buf ( n45259 , n45233 );
buf ( n45260 , n45252 );
xor ( n45261 , n45258 , n45259 );
xor ( n45262 , n45261 , n45260 );
buf ( n45263 , n45262 );
xor ( n45264 , n45258 , n45259 );
and ( n45265 , n45264 , n45260 );
and ( n45266 , n45258 , n45259 );
or ( n45267 , n45265 , n45266 );
buf ( n45268 , n45267 );
buf ( n45269 , n45193 );
buf ( n45270 , n45263 );
buf ( n45271 , n45204 );
xor ( n45272 , n45269 , n45270 );
xor ( n45273 , n45272 , n45271 );
buf ( n45274 , n45273 );
xor ( n45275 , n45269 , n45270 );
and ( n45276 , n45275 , n45271 );
and ( n45277 , n45269 , n45270 );
or ( n45278 , n45276 , n45277 );
buf ( n45279 , n45278 );
buf ( n45280 , n521 );
buf ( n45281 , n540 );
and ( n45282 , n45280 , n45281 );
buf ( n45283 , n45282 );
buf ( n45284 , n45283 );
buf ( n45285 , n522 );
buf ( n45286 , n539 );
and ( n45287 , n45285 , n45286 );
buf ( n45288 , n45287 );
buf ( n45289 , n45288 );
buf ( n45290 , n524 );
not ( n45291 , n45290 );
buf ( n45292 , n537 );
not ( n45293 , n45292 );
buf ( n45294 , n45293 );
buf ( n45295 , n45294 );
nor ( n45296 , n45291 , n45295 );
buf ( n45297 , n45296 );
buf ( n45298 , n45297 );
xor ( n45299 , n45284 , n45289 );
xor ( n45300 , n45299 , n45298 );
buf ( n45301 , n45300 );
xor ( n45302 , n45284 , n45289 );
and ( n45303 , n45302 , n45298 );
and ( n45304 , n45284 , n45289 );
or ( n45305 , n45303 , n45304 );
buf ( n45306 , n45305 );
buf ( n45307 , n523 );
not ( n45308 , n45307 );
buf ( n45309 , n45308 );
buf ( n45310 , n45309 );
buf ( n45311 , n37921 );
nor ( n45312 , n45310 , n45311 );
buf ( n45313 , n45312 );
buf ( n45314 , n45313 );
buf ( n45315 , n45238 );
buf ( n45316 , n45301 );
xor ( n45317 , n45314 , n45315 );
xor ( n45318 , n45317 , n45316 );
buf ( n45319 , n45318 );
xor ( n45320 , n45314 , n45315 );
and ( n45321 , n45320 , n45316 );
and ( n45322 , n45314 , n45315 );
or ( n45323 , n45321 , n45322 );
buf ( n45324 , n45323 );
buf ( n45325 , n45257 );
buf ( n45326 , n45319 );
buf ( n45327 , n45268 );
xor ( n45328 , n45325 , n45326 );
xor ( n45329 , n45328 , n45327 );
buf ( n45330 , n45329 );
xor ( n45331 , n45325 , n45326 );
and ( n45332 , n45331 , n45327 );
and ( n45333 , n45325 , n45326 );
or ( n45334 , n45332 , n45333 );
buf ( n45335 , n45334 );
buf ( n45336 , n539 );
not ( n45337 , n45336 );
buf ( n45338 , n521 );
not ( n45339 , n45338 );
buf ( n45340 , n45339 );
buf ( n45341 , n45340 );
nor ( n45342 , n45337 , n45341 );
buf ( n45343 , n45342 );
buf ( n45344 , n45343 );
buf ( n45345 , n522 );
not ( n45346 , n45345 );
buf ( n45347 , n45346 );
buf ( n45348 , n45347 );
buf ( n45349 , n37921 );
nor ( n45350 , n45348 , n45349 );
buf ( n45351 , n45350 );
buf ( n45352 , n45351 );
buf ( n45353 , n45309 );
buf ( n45354 , n45294 );
nor ( n45355 , n45353 , n45354 );
buf ( n45356 , n45355 );
buf ( n45357 , n45356 );
xor ( n45358 , n45344 , n45352 );
xor ( n45359 , n45358 , n45357 );
buf ( n45360 , n45359 );
xor ( n45361 , n45344 , n45352 );
and ( n45362 , n45361 , n45357 );
and ( n45363 , n45344 , n45352 );
or ( n45364 , n45362 , n45363 );
buf ( n45365 , n45364 );
buf ( n45366 , n45306 );
buf ( n45367 , n45360 );
buf ( n45368 , n45324 );
xor ( n45369 , n45366 , n45367 );
xor ( n45370 , n45369 , n45368 );
buf ( n45371 , n45370 );
xor ( n45372 , n45366 , n45367 );
and ( n45373 , n45372 , n45368 );
and ( n45374 , n45366 , n45367 );
or ( n45375 , n45373 , n45374 );
buf ( n45376 , n45375 );
buf ( n45377 , n45340 );
buf ( n45378 , n37921 );
nor ( n45379 , n45377 , n45378 );
buf ( n45380 , n45379 );
buf ( n45381 , n45380 );
buf ( n45382 , n45347 );
buf ( n45383 , n45294 );
nor ( n45384 , n45382 , n45383 );
buf ( n45385 , n45384 );
buf ( n45386 , n45385 );
buf ( n45387 , n45365 );
xor ( n45388 , n45381 , n45386 );
xor ( n45389 , n45388 , n45387 );
buf ( n45390 , n45389 );
xor ( n45391 , n45381 , n45386 );
and ( n45392 , n45391 , n45387 );
and ( n45393 , n45381 , n45386 );
or ( n45394 , n45392 , n45393 );
buf ( n45395 , n45394 );
or ( n45396 , n45136 , n45210 );
and ( n45397 , n44631 , n45396 );
buf ( n45398 , n45397 );
buf ( n45399 , n44669 );
and ( n45400 , n44623 , n45396 );
and ( n45401 , n45136 , n45210 );
nor ( n45402 , n45400 , n45401 );
buf ( n45403 , n45402 );
not ( n45404 , n45398 );
not ( n45405 , n45399 );
or ( n45406 , n45404 , n45405 );
nand ( n45407 , n45406 , n45403 );
buf ( n45408 , n45407 );
buf ( n45409 , n44631 );
buf ( n45410 , n44669 );
buf ( n45411 , n44626 );
not ( n45412 , n45409 );
not ( n45413 , n45410 );
or ( n45414 , n45412 , n45413 );
nand ( n45415 , n45414 , n45411 );
buf ( n45416 , n45415 );
buf ( n45417 , n45215 );
not ( n45418 , n45417 );
buf ( n45419 , n45418 );
buf ( n45420 , n45419 );
buf ( n45421 , n45274 );
not ( n45422 , n45421 );
buf ( n45423 , n45422 );
buf ( n45424 , n45423 );
nand ( n45425 , n45420 , n45424 );
buf ( n45426 , n45425 );
and ( n45427 , n45396 , n45426 );
buf ( n45428 , n45427 );
buf ( n45429 , n45279 );
buf ( n45430 , n45330 );
or ( n45431 , n45429 , n45430 );
buf ( n45432 , n45431 );
buf ( n45433 , n45432 );
and ( n45434 , n45428 , n45433 );
buf ( n45435 , n45434 );
buf ( n45436 , n45435 );
buf ( n45437 , n44631 );
and ( n45438 , n45436 , n45437 );
buf ( n45439 , n45438 );
buf ( n45440 , n45439 );
buf ( n45441 , n44669 );
buf ( n45442 , n45435 );
buf ( n45443 , n44623 );
and ( n45444 , n45442 , n45443 );
not ( n45445 , n45426 );
buf ( n45446 , n45432 );
not ( n45447 , n45446 );
buf ( n45448 , n45447 );
nor ( n45449 , n45445 , n45448 );
not ( n45450 , n45449 );
not ( n45451 , n45401 );
or ( n45452 , n45450 , n45451 );
buf ( n45453 , n45419 );
buf ( n45454 , n45423 );
nor ( n45455 , n45453 , n45454 );
buf ( n45456 , n45455 );
not ( n45457 , n45456 );
not ( n45458 , n45457 );
not ( n45459 , n45448 );
and ( n45460 , n45458 , n45459 );
buf ( n45461 , n45279 );
buf ( n45462 , n45330 );
nand ( n45463 , n45461 , n45462 );
buf ( n45464 , n45463 );
not ( n45465 , n45464 );
nor ( n45466 , n45460 , n45465 );
nand ( n45467 , n45452 , n45466 );
buf ( n45468 , n45467 );
nor ( n45469 , n45444 , n45468 );
buf ( n45470 , n45469 );
buf ( n45471 , n45470 );
not ( n45472 , n45440 );
not ( n45473 , n45441 );
or ( n45474 , n45472 , n45473 );
nand ( n45475 , n45474 , n45471 );
buf ( n45476 , n45475 );
buf ( n45477 , n45335 );
buf ( n45478 , n45371 );
or ( n45479 , n45477 , n45478 );
buf ( n45480 , n45479 );
buf ( n45481 , n45480 );
buf ( n45482 , n44667 );
buf ( n45483 , n45439 );
nand ( n45484 , n45482 , n45483 );
buf ( n45485 , n45484 );
buf ( n45486 , n45485 );
buf ( n45487 , n45470 );
nand ( n45488 , n45486 , n45487 );
buf ( n45489 , n45488 );
buf ( n45490 , n45489 );
buf ( n45491 , n45335 );
buf ( n45492 , n45371 );
nand ( n45493 , n45491 , n45492 );
buf ( n45494 , n45493 );
buf ( n45495 , n45494 );
not ( n45496 , n45481 );
not ( n45497 , n45490 );
or ( n45498 , n45496 , n45497 );
nand ( n45499 , n45498 , n45495 );
buf ( n45500 , n45499 );
buf ( n45501 , n45467 );
buf ( n45502 , n45480 );
not ( n45503 , n45502 );
buf ( n45504 , n45376 );
buf ( n45505 , n45390 );
nor ( n45506 , n45504 , n45505 );
buf ( n45507 , n45506 );
buf ( n45508 , n45507 );
nor ( n45509 , n45503 , n45508 );
buf ( n45510 , n45509 );
buf ( n45511 , n45510 );
and ( n45512 , n45501 , n45511 );
buf ( n45513 , n45494 );
buf ( n45514 , n45507 );
or ( n45515 , n45513 , n45514 );
buf ( n45516 , n45376 );
buf ( n45517 , n45390 );
nand ( n45518 , n45516 , n45517 );
buf ( n45519 , n45518 );
buf ( n45520 , n45519 );
nand ( n45521 , n45515 , n45520 );
buf ( n45522 , n45521 );
buf ( n45523 , n45522 );
nor ( n45524 , n45512 , n45523 );
buf ( n45525 , n45524 );
buf ( n45526 , n45525 );
not ( n45527 , n45526 );
buf ( n45528 , n45527 );
buf ( n45529 , n45528 );
buf ( n45530 , n45395 );
not ( n45531 , n45530 );
buf ( n45532 , n45531 );
buf ( n45533 , n45532 );
buf ( n45534 , n521 );
buf ( n45535 , n537 );
nand ( n45536 , n45534 , n45535 );
buf ( n45537 , n45536 );
buf ( n45538 , n45537 );
nand ( n45539 , n45533 , n45538 );
buf ( n45540 , n45539 );
buf ( n45541 , n45540 );
buf ( n45542 , n45532 );
buf ( n45543 , n45537 );
nor ( n45544 , n45542 , n45543 );
buf ( n45545 , n45544 );
buf ( n45546 , n45545 );
and ( n45547 , n45529 , n45541 );
nor ( n45548 , n45547 , n45546 );
buf ( n45549 , n45548 );
and ( n45550 , n44623 , n45427 );
and ( n45551 , n45401 , n45426 );
nor ( n45552 , n45550 , n45551 , n45456 );
buf ( n45553 , n45552 );
buf ( n45554 , n45448 );
or ( n45555 , n45553 , n45554 );
buf ( n45556 , n45464 );
nand ( n45557 , n45555 , n45556 );
buf ( n45558 , n45557 );
buf ( n45559 , n45558 );
buf ( n45560 , n45510 );
buf ( n45561 , n45522 );
and ( n45562 , n45559 , n45560 );
nor ( n45563 , n45562 , n45561 );
buf ( n45564 , n45563 );
buf ( n45565 , n45439 );
buf ( n45566 , n45480 );
nand ( n45567 , n45565 , n45566 );
buf ( n45568 , n45567 );
buf ( n45569 , n45435 );
buf ( n45570 , n45510 );
buf ( n45571 , n45540 );
and ( n45572 , n45569 , n45570 , n45571 );
buf ( n45573 , n45572 );
buf ( n45574 , n44631 );
buf ( n45575 , n45427 );
and ( n45576 , n45574 , n45575 );
buf ( n45577 , n45576 );
buf ( n45578 , n45577 );
buf ( n45579 , n45432 );
buf ( n45580 , n45510 );
and ( n45581 , n45578 , n45579 , n45580 );
buf ( n45582 , n45581 );
buf ( n45583 , n45456 );
buf ( n45584 , n45426 );
not ( n45585 , n45583 );
nand ( n45586 , n45585 , n45584 );
buf ( n45587 , n45586 );
buf ( n45588 , n45480 );
buf ( n45589 , n45494 );
nand ( n45590 , n45588 , n45589 );
buf ( n45591 , n45590 );
buf ( n45592 , n31300 );
buf ( n45593 , n31306 );
not ( n45594 , n45593 );
buf ( n45595 , n31257 );
nand ( n45596 , n45594 , n45595 );
buf ( n45597 , n45596 );
buf ( n45598 , n45597 );
buf ( n45599 , n45597 );
buf ( n45600 , n31300 );
not ( n45601 , n45592 );
not ( n45602 , n45598 );
or ( n45603 , n45601 , n45602 );
or ( n45604 , n45599 , n45600 );
nand ( n45605 , n45603 , n45604 );
buf ( n45606 , n45605 );
buf ( n45607 , n45545 );
buf ( n45608 , n45540 );
not ( n45609 , n45607 );
nand ( n45610 , n45609 , n45608 );
buf ( n45611 , n45610 );
xor ( n45612 , n31267 , n31291 );
xor ( n45613 , n45612 , n31296 );
buf ( n45614 , n45613 );
xor ( n45615 , n31272 , n31282 );
xor ( n45616 , n45615 , n31286 );
buf ( n45617 , n45616 );
buf ( n45618 , n472 );
buf ( n45619 , n31278 );
buf ( n45620 , n31278 );
buf ( n45621 , n472 );
not ( n45622 , n45618 );
not ( n45623 , n45619 );
or ( n45624 , n45622 , n45623 );
or ( n45625 , n45620 , n45621 );
nand ( n45626 , n45624 , n45625 );
buf ( n45627 , n45626 );
not ( n45628 , n45582 );
not ( n45629 , n44669 );
or ( n45630 , n45628 , n45629 );
nand ( n45631 , n45630 , n45564 );
buf ( n45632 , n45631 );
buf ( n45633 , n45611 );
xnor ( n45634 , n45632 , n45633 );
buf ( n45635 , n45634 );
buf ( n45636 , n30470 );
not ( n45637 , n45636 );
buf ( n45638 , n30393 );
nand ( n45639 , n45637 , n45638 );
buf ( n45640 , n45639 );
buf ( n45641 , n45640 );
buf ( n45642 , n30453 );
not ( n45643 , n45642 );
buf ( n45644 , n30461 );
nand ( n45645 , n45643 , n45644 );
buf ( n45646 , n45645 );
buf ( n45647 , n45646 );
buf ( n45648 , n45646 );
buf ( n45649 , n45640 );
not ( n45650 , n45641 );
not ( n45651 , n45647 );
or ( n45652 , n45650 , n45651 );
or ( n45653 , n45648 , n45649 );
nand ( n45654 , n45652 , n45653 );
buf ( n45655 , n45654 );
buf ( n45656 , n30436 );
buf ( n45657 , n30450 );
buf ( n45658 , n30461 );
nand ( n45659 , n45657 , n45658 );
buf ( n45660 , n45659 );
buf ( n45661 , n45660 );
buf ( n45662 , n45660 );
buf ( n45663 , n30436 );
not ( n45664 , n45656 );
not ( n45665 , n45661 );
or ( n45666 , n45664 , n45665 );
or ( n45667 , n45662 , n45663 );
nand ( n45668 , n45666 , n45667 );
buf ( n45669 , n45668 );
buf ( n45670 , n44193 );
not ( n45671 , n29519 );
not ( n45672 , n44384 );
or ( n45673 , n44303 , n45672 );
not ( n45674 , n44391 );
not ( n45675 , n44384 );
or ( n45676 , n45674 , n45675 );
nand ( n45677 , n45676 , n44385 );
not ( n45678 , n45677 );
nand ( n45679 , n45673 , n45678 );
and ( n45680 , n44940 , n44992 );
not ( n45681 , n45680 );
or ( n45682 , n44940 , n44992 );
nand ( n45683 , n45681 , n45682 );
not ( n45684 , n45683 );
and ( n45685 , n45679 , n45684 );
not ( n45686 , n45679 );
and ( n45687 , n45686 , n45683 );
nor ( n45688 , n45685 , n45687 );
not ( n45689 , n45688 );
or ( n45690 , n45671 , n45689 );
not ( n45691 , n44289 );
nor ( n45692 , n45691 , n44199 );
not ( n45693 , n45692 );
not ( n45694 , n41973 );
or ( n45695 , n45693 , n45694 );
not ( n45696 , n44289 );
not ( n45697 , n44207 );
or ( n45698 , n45696 , n45697 );
nand ( n45699 , n45698 , n44290 );
not ( n45700 , n45699 );
nand ( n45701 , n45695 , n45700 );
and ( n45702 , n44766 , n44818 );
not ( n45703 , n45702 );
or ( n45704 , n44766 , n44818 );
nand ( n45705 , n45703 , n45704 );
not ( n45706 , n45705 );
and ( n45707 , n45701 , n45706 );
not ( n45708 , n45701 );
and ( n45709 , n45708 , n45705 );
nor ( n45710 , n45707 , n45709 );
nand ( n45711 , n45710 , n455 );
nand ( n45712 , n45690 , n45711 );
not ( n45713 , n45712 );
not ( n45714 , n44292 );
not ( n45715 , n44295 );
or ( n45716 , n45714 , n45715 );
nand ( n45717 , n45716 , n44402 );
not ( n45718 , n45717 );
not ( n45719 , n45718 );
or ( n45720 , n45713 , n45719 );
nand ( n45721 , n45720 , n44404 );
not ( n45722 , n45721 );
buf ( n45723 , n45722 );
nand ( n45724 , n45670 , n45723 );
buf ( n45725 , n45724 );
buf ( n45726 , n44404 );
buf ( n45727 , n44193 );
nand ( n45728 , n45726 , n45727 );
buf ( n45729 , n45728 );
xor ( n45730 , n30396 , n30411 );
xor ( n45731 , n45730 , n30432 );
buf ( n45732 , n45731 );
xor ( n45733 , n30413 , n30429 );
buf ( n45734 , n45733 );
not ( n45735 , n29519 );
not ( n45736 , n45688 );
or ( n45737 , n45735 , n45736 );
nand ( n45738 , n45737 , n45711 );
not ( n45739 , n45738 );
not ( n45740 , n29519 );
nand ( n45741 , n44384 , n45682 );
nor ( n45742 , n44301 , n45741 );
not ( n45743 , n45742 );
not ( n45744 , n41692 );
or ( n45745 , n45743 , n45744 );
and ( n45746 , n45677 , n45682 );
nor ( n45747 , n45746 , n45680 );
nand ( n45748 , n45745 , n45747 );
or ( n45749 , n44997 , n45043 );
nand ( n45750 , n44997 , n45043 );
nand ( n45751 , n45749 , n45750 );
xnor ( n45752 , n45748 , n45751 );
not ( n45753 , n45752 );
or ( n45754 , n45740 , n45753 );
nand ( n45755 , n44289 , n45704 );
nor ( n45756 , n44199 , n45755 );
not ( n45757 , n45756 );
not ( n45758 , n41973 );
or ( n45759 , n45757 , n45758 );
and ( n45760 , n45699 , n45704 );
nor ( n45761 , n45760 , n45702 );
nand ( n45762 , n45759 , n45761 );
or ( n45763 , n44823 , n44872 );
nand ( n45764 , n44823 , n44872 );
nand ( n45765 , n45763 , n45764 );
not ( n45766 , n45765 );
and ( n45767 , n45762 , n45766 );
not ( n45768 , n45762 );
and ( n45769 , n45768 , n45765 );
nor ( n45770 , n45767 , n45769 );
nand ( n45771 , n45770 , n455 );
nand ( n45772 , n45754 , n45771 );
nor ( n45773 , n45739 , n45772 );
buf ( n45774 , n45773 );
buf ( n45775 , n45774 );
buf ( n45776 , n45775 );
xor ( n45777 , n43397 , n43403 );
and ( n45778 , n45777 , n43410 );
and ( n45779 , n43397 , n43403 );
or ( n45780 , n45778 , n45779 );
xor ( n45781 , n43413 , n43419 );
and ( n45782 , n45781 , n43178 );
and ( n45783 , n43413 , n43419 );
or ( n45784 , n45782 , n45783 );
xor ( n45785 , n43395 , n43411 );
and ( n45786 , n45785 , n43421 );
and ( n45787 , n43395 , n43411 );
or ( n45788 , n45786 , n45787 );
xor ( n45789 , n43391 , n43422 );
and ( n45790 , n45789 , n43427 );
and ( n45791 , n43391 , n43422 );
or ( n45792 , n45790 , n45791 );
nor ( n45793 , n43036 , n42221 );
or ( n45794 , n42306 , n43417 );
and ( n45795 , n42261 , n42419 );
and ( n45796 , n42263 , n490 );
nor ( n45797 , n45795 , n45796 );
or ( n45798 , n42271 , n45797 );
nand ( n45799 , n45794 , n45798 );
xor ( n45800 , n45793 , n45799 );
or ( n45801 , n42315 , n43408 );
and ( n45802 , n43035 , n42276 );
and ( n45803 , n43036 , n492 );
nor ( n45804 , n45802 , n45803 );
or ( n45805 , n42321 , n45804 );
nand ( n45806 , n45801 , n45805 );
xor ( n45807 , n45800 , n45806 );
xor ( n45808 , n45793 , n45799 );
and ( n45809 , n45808 , n45806 );
and ( n45810 , n45793 , n45799 );
or ( n45811 , n45809 , n45810 );
or ( n45812 , n42457 , n43401 );
or ( n45813 , n42456 , n42189 );
nand ( n45814 , n45812 , n45813 );
not ( n45815 , n45814 );
xor ( n45816 , n45815 , n45780 );
xor ( n45817 , n45816 , n45807 );
xor ( n45818 , n45815 , n45780 );
and ( n45819 , n45818 , n45807 );
and ( n45820 , n45815 , n45780 );
or ( n45821 , n45819 , n45820 );
xor ( n45822 , n45784 , n45817 );
xor ( n45823 , n45822 , n45788 );
xor ( n45824 , n45784 , n45817 );
and ( n45825 , n45824 , n45788 );
and ( n45826 , n45784 , n45817 );
or ( n45827 , n45825 , n45826 );
not ( n45828 , n42457 );
or ( n45829 , n45828 , n43218 );
nand ( n45830 , n45829 , n42204 );
or ( n45831 , n42306 , n45797 );
and ( n45832 , n42261 , n5539 );
and ( n45833 , n42263 , n489 );
nor ( n45834 , n45832 , n45833 );
or ( n45835 , n42271 , n45834 );
nand ( n45836 , n45831 , n45835 );
xor ( n45837 , n45830 , n45836 );
nor ( n45838 , n43036 , n42382 );
xor ( n45839 , n45837 , n45838 );
xor ( n45840 , n45830 , n45836 );
and ( n45841 , n45840 , n45838 );
and ( n45842 , n45830 , n45836 );
or ( n45843 , n45841 , n45842 );
or ( n45844 , n42315 , n45804 );
and ( n45845 , n43035 , n42282 );
and ( n45846 , n43036 , n491 );
nor ( n45847 , n45845 , n45846 );
or ( n45848 , n42321 , n45847 );
nand ( n45849 , n45844 , n45848 );
xor ( n45850 , n45849 , n45814 );
xor ( n45851 , n45850 , n45811 );
xor ( n45852 , n45849 , n45814 );
and ( n45853 , n45852 , n45811 );
and ( n45854 , n45849 , n45814 );
or ( n45855 , n45853 , n45854 );
xor ( n45856 , n45839 , n45851 );
xor ( n45857 , n45856 , n45821 );
xor ( n45858 , n45839 , n45851 );
and ( n45859 , n45858 , n45821 );
and ( n45860 , n45839 , n45851 );
or ( n45861 , n45859 , n45860 );
or ( n45862 , n42315 , n45847 );
and ( n45863 , n43035 , n42419 );
and ( n45864 , n41312 , n490 );
nor ( n45865 , n45863 , n45864 );
or ( n45866 , n42321 , n45865 );
nand ( n45867 , n45862 , n45866 );
nor ( n45868 , n43036 , n42276 );
xor ( n45869 , n45867 , n45868 );
not ( n45870 , n45834 );
and ( n45871 , n42305 , n45870 );
not ( n45872 , n42271 );
and ( n45873 , n45872 , n42261 );
nor ( n45874 , n45871 , n45873 );
xor ( n45875 , n45869 , n45874 );
xor ( n45876 , n45867 , n45868 );
and ( n45877 , n45876 , n45874 );
and ( n45878 , n45867 , n45868 );
or ( n45879 , n45877 , n45878 );
xor ( n45880 , n45843 , n45875 );
xor ( n45881 , n45880 , n45855 );
xor ( n45882 , n45843 , n45875 );
and ( n45883 , n45882 , n45855 );
and ( n45884 , n45843 , n45875 );
or ( n45885 , n45883 , n45884 );
or ( n45886 , n42305 , n45872 );
nand ( n45887 , n45886 , n42261 );
or ( n45888 , n42315 , n45865 );
and ( n45889 , n43035 , n5539 );
and ( n45890 , n43036 , n489 );
nor ( n45891 , n45889 , n45890 );
or ( n45892 , n42321 , n45891 );
nand ( n45893 , n45888 , n45892 );
xor ( n45894 , n45887 , n45893 );
nor ( n45895 , n43036 , n42282 );
xor ( n45896 , n45894 , n45895 );
xor ( n45897 , n45887 , n45893 );
and ( n45898 , n45897 , n45895 );
and ( n45899 , n45887 , n45893 );
or ( n45900 , n45898 , n45899 );
not ( n45901 , n45874 );
xor ( n45902 , n45901 , n45896 );
xor ( n45903 , n45902 , n45879 );
xor ( n45904 , n45901 , n45896 );
and ( n45905 , n45904 , n45879 );
and ( n45906 , n45901 , n45896 );
or ( n45907 , n45905 , n45906 );
or ( n45908 , n42315 , n45891 );
or ( n45909 , n42321 , n43036 );
nand ( n45910 , n45908 , n45909 );
nand ( n45911 , n43035 , n490 );
xor ( n45912 , n45910 , n45911 );
xor ( n45913 , n45912 , n45900 );
xor ( n45914 , n45910 , n45911 );
and ( n45915 , n45914 , n45900 );
and ( n45916 , n45910 , n45911 );
or ( n45917 , n45915 , n45916 );
or ( n45918 , n45792 , n45823 );
not ( n45919 , n45918 );
and ( n45920 , n43193 , n43430 );
not ( n45921 , n45920 );
not ( n45922 , n43374 );
or ( n45923 , n45921 , n45922 );
not ( n45924 , n43375 );
not ( n45925 , n43193 );
or ( n45926 , n45924 , n45925 );
nand ( n45927 , n45926 , n43194 );
and ( n45928 , n45927 , n43430 );
nor ( n45929 , n45928 , n43432 );
nand ( n45930 , n45923 , n45929 );
not ( n45931 , n45930 );
or ( n45932 , n45919 , n45931 );
nand ( n45933 , n45792 , n45823 );
nand ( n45934 , n45932 , n45933 );
or ( n45935 , n43357 , n43347 );
not ( n45936 , n45935 );
not ( n45937 , n43336 );
not ( n45938 , n42863 );
not ( n45939 , n42784 );
or ( n45940 , n45938 , n45939 );
nand ( n45941 , n45940 , n43198 );
not ( n45942 , n45941 );
or ( n45943 , n45937 , n45942 );
nand ( n45944 , n45943 , n43354 );
not ( n45945 , n45944 );
or ( n45946 , n45936 , n45945 );
or ( n45947 , n45944 , n45935 );
nand ( n45948 , n45946 , n45947 );
nand ( n45949 , n43336 , n43354 );
not ( n45950 , n45949 );
not ( n45951 , n45941 );
or ( n45952 , n45950 , n45951 );
or ( n45953 , n45941 , n45949 );
nand ( n45954 , n45952 , n45953 );
xor ( n45955 , n42661 , n42663 );
xor ( n45956 , n45955 , n42779 );
nor ( n45957 , n45827 , n45857 );
not ( n45958 , n45957 );
not ( n45959 , n45933 );
and ( n45960 , n45958 , n45959 );
and ( n45961 , n45827 , n45857 );
nor ( n45962 , n45960 , n45961 );
or ( n45963 , n45861 , n45881 );
not ( n45964 , n45963 );
nor ( n45965 , n45885 , n45903 );
nor ( n45966 , n45964 , n45965 );
not ( n45967 , n45966 );
or ( n45968 , n45962 , n45967 );
nand ( n45969 , n45861 , n45881 );
not ( n45970 , n45969 );
not ( n45971 , n45965 );
and ( n45972 , n45970 , n45971 );
and ( n45973 , n45903 , n45885 );
nor ( n45974 , n45972 , n45973 );
nand ( n45975 , n45968 , n45974 );
not ( n45976 , n45907 );
not ( n45977 , n45913 );
nand ( n45978 , n45976 , n45977 );
and ( n45979 , n45975 , n45978 );
nor ( n45980 , n45976 , n45977 );
nor ( n45981 , n45979 , n45980 );
nand ( n45982 , n43306 , n43360 );
not ( n45983 , n45918 );
nor ( n45984 , n45983 , n45957 );
and ( n45985 , n45984 , n45966 , n45978 );
xor ( n45986 , n42756 , n42758 );
xor ( n45987 , n45986 , n42767 );
nand ( n45988 , n45918 , n45933 );
or ( n45989 , n45961 , n45957 );
nand ( n45990 , n45963 , n45969 );
or ( n45991 , n45965 , n45973 );
not ( n45992 , n7399 );
nand ( n45993 , n7291 , n7402 );
not ( n45994 , n45993 );
or ( n45995 , n45992 , n45994 );
or ( n45996 , n45993 , n7399 );
nand ( n45997 , n45995 , n45996 );
not ( n45998 , n45980 );
nand ( n45999 , n45998 , n45978 );
not ( n46000 , n45917 );
not ( n46001 , n42321 );
or ( n46002 , n42956 , n46001 );
nand ( n46003 , n46002 , n43035 );
nor ( n46004 , n43036 , n5539 );
xor ( n46005 , n46003 , n46004 );
not ( n46006 , n45911 );
xor ( n46007 , n46005 , n46006 );
not ( n46008 , n46007 );
and ( n46009 , n46000 , n46008 );
and ( n46010 , n45917 , n46007 );
nor ( n46011 , n46009 , n46010 );
not ( n46012 , n7391 );
not ( n46013 , n7342 );
nand ( n46014 , n46013 , n7394 );
not ( n46015 , n46014 );
or ( n46016 , n46012 , n46015 );
or ( n46017 , n46014 , n7391 );
nand ( n46018 , n46016 , n46017 );
and ( n46019 , n7295 , n7320 );
not ( n46020 , n7398 );
nor ( n46021 , n46019 , n46020 );
not ( n46022 , n7384 );
not ( n46023 , n7386 );
nor ( n46024 , n46023 , n7375 );
not ( n46025 , n46024 );
or ( n46026 , n46022 , n46025 );
or ( n46027 , n46024 , n7384 );
nand ( n46028 , n46026 , n46027 );
not ( n46029 , n7383 );
and ( n46030 , n46029 , n7377 );
not ( n46031 , n7384 );
nor ( n46032 , n46030 , n46031 );
not ( n46033 , n7376 );
not ( n46034 , n44905 );
not ( n46035 , n44935 );
and ( n46036 , n46034 , n46035 );
and ( n46037 , n44905 , n44935 );
nor ( n46038 , n46036 , n46037 );
nor ( n46039 , n46038 , n29519 );
nand ( n46040 , n46038 , n455 );
or ( n46041 , n44877 , n44900 );
nand ( n46042 , n44877 , n44900 );
nand ( n46043 , n46041 , n46042 );
not ( n46044 , n45076 );
not ( n46045 , n45106 );
and ( n46046 , n46044 , n46045 );
and ( n46047 , n45076 , n45106 );
nor ( n46048 , n46046 , n46047 );
nand ( n46049 , n45048 , n45071 );
or ( n46050 , n45048 , n45071 );
xor ( n46051 , n7395 , n46021 );
not ( n46052 , n45763 );
not ( n46053 , n45762 );
or ( n46054 , n46052 , n46053 );
nand ( n46055 , n46054 , n45764 );
not ( n46056 , n46043 );
and ( n46057 , n46055 , n46056 );
nor ( n46058 , n46057 , n37874 );
not ( n46059 , n46058 );
or ( n46060 , n44823 , n44872 );
nand ( n46061 , n46060 , n45762 );
nand ( n46062 , n46061 , n45764 , n46043 );
not ( n46063 , n46062 );
or ( n46064 , n46059 , n46063 );
nand ( n46065 , n46050 , n46049 );
not ( n46066 , n46065 );
not ( n46067 , n45749 );
not ( n46068 , n45748 );
or ( n46069 , n46067 , n46068 );
buf ( n46070 , n45750 );
nand ( n46071 , n46069 , n46070 );
not ( n46072 , n46071 );
or ( n46073 , n46066 , n46072 );
or ( n46074 , n46065 , n46071 );
nand ( n46075 , n46073 , n46074 );
nand ( n46076 , n46075 , n29519 );
nand ( n46077 , n46064 , n46076 );
not ( n46078 , n46077 );
not ( n46079 , n45772 );
not ( n46080 , n46079 );
or ( n46081 , n46078 , n46080 );
nand ( n46082 , n45739 , n45772 );
nand ( n46083 , n46081 , n46082 );
not ( n46084 , n46083 );
buf ( n46085 , n44405 );
not ( n46086 , n46085 );
buf ( n46087 , n45718 );
buf ( n46088 , n45712 );
nand ( n46089 , n46087 , n46088 );
buf ( n46090 , n46089 );
buf ( n46091 , n46090 );
not ( n46092 , n46091 );
or ( n46093 , n46086 , n46092 );
not ( n46094 , n45718 );
nand ( n46095 , n46094 , n45739 );
buf ( n46096 , n46095 );
nand ( n46097 , n46093 , n46096 );
buf ( n46098 , n46097 );
and ( n46099 , n46084 , n46098 );
buf ( n46100 , n45773 );
not ( n46101 , n46100 );
nand ( n46102 , n46077 , n46079 );
buf ( n46103 , n46102 );
not ( n46104 , n46103 );
or ( n46105 , n46101 , n46104 );
not ( n46106 , n46058 );
not ( n46107 , n46062 );
or ( n46108 , n46106 , n46107 );
nand ( n46109 , n46075 , n29519 );
nand ( n46110 , n46108 , n46109 );
or ( n46111 , n46110 , n46079 );
buf ( n46112 , n46111 );
nand ( n46113 , n46105 , n46112 );
buf ( n46114 , n46113 );
nor ( n46115 , n46099 , n46114 );
buf ( n46116 , n46110 );
not ( n46117 , n46116 );
buf ( n46118 , n46117 );
not ( n46119 , n46118 );
not ( n46120 , n46041 );
not ( n46121 , n46055 );
or ( n46122 , n46120 , n46121 );
nand ( n46123 , n46122 , n46042 );
nor ( n46124 , n46123 , n46040 );
not ( n46125 , n46124 );
not ( n46126 , n46050 );
not ( n46127 , n46071 );
or ( n46128 , n46126 , n46127 );
nand ( n46129 , n46128 , n46049 );
nor ( n46130 , n46048 , n455 );
and ( n46131 , n46129 , n46130 );
not ( n46132 , n46129 );
and ( n46133 , n46048 , n29519 );
and ( n46134 , n46132 , n46133 );
nor ( n46135 , n46131 , n46134 );
nand ( n46136 , n46123 , n46039 );
nand ( n46137 , n46125 , n46135 , n46136 );
nor ( n46138 , n46119 , n46137 );
nand ( n46139 , n44196 , n46115 , n46138 );
not ( n46140 , n46139 );
nand ( n46141 , n46084 , n45722 );
not ( n46142 , n46141 );
nand ( n46143 , n46137 , n46118 );
not ( n46144 , n46143 );
not ( n46145 , n46144 );
not ( n46146 , n41026 );
not ( n46147 , n44172 );
nand ( n46148 , n46142 , n46145 , n46146 , n46147 );
nand ( n46149 , n46140 , n46148 );
buf ( n46150 , n46149 );
not ( n46151 , n46150 );
buf ( n46152 , n46151 );
buf ( n46153 , n45930 );
nand ( n46154 , n44742 , n7047 );
not ( n46155 , n2356 );
not ( n46156 , n45591 );
and ( n46157 , n45476 , n46156 );
not ( n46158 , n45476 );
and ( n46159 , n46158 , n45591 );
nor ( n46160 , n46157 , n46159 );
not ( n46161 , n46160 );
or ( n46162 , n46155 , n46161 );
nand ( n46163 , n46084 , n45722 );
not ( n46164 , n46163 );
nand ( n46165 , n46164 , n44193 );
nand ( n46166 , n46164 , n46146 , n46147 );
nand ( n46167 , n46165 , n46166 , n46115 );
not ( n46168 , n46167 );
not ( n46169 , n46118 );
not ( n46170 , n46137 );
and ( n46171 , n46169 , n46170 );
nor ( n46172 , n46171 , n46144 );
not ( n46173 , n46172 );
nand ( n46174 , n46168 , n46173 );
nand ( n46175 , n46167 , n46172 );
nand ( n46176 , n46174 , n46175 , n454 );
nand ( n46177 , n46162 , n46176 );
buf ( n46178 , n46177 );
not ( n46179 , n2356 );
not ( n46180 , n45401 );
nand ( n46181 , n46180 , n45396 );
xnor ( n46182 , n45416 , n46181 );
not ( n46183 , n46182 );
or ( n46184 , n46179 , n46183 );
not ( n46185 , n45729 );
and ( n46186 , n46090 , n46095 );
buf ( n46187 , n46186 );
nand ( n46188 , n46185 , n46187 );
not ( n46189 , n46186 );
buf ( n46190 , n46146 );
buf ( n46191 , n44173 );
buf ( n46192 , n44404 );
nand ( n46193 , n46190 , n46191 , n46192 );
buf ( n46194 , n46193 );
nor ( n46195 , n46189 , n46194 );
not ( n46196 , n46186 );
not ( n46197 , n44408 );
not ( n46198 , n46197 );
or ( n46199 , n46196 , n46198 );
nand ( n46200 , n46199 , n454 );
nor ( n46201 , n46195 , n46200 );
nor ( n46202 , n46197 , n46186 );
nand ( n46203 , n45729 , n46202 , n46194 );
nand ( n46204 , n46188 , n46201 , n46203 );
nand ( n46205 , n46184 , n46204 );
nand ( n46206 , n46177 , n46205 );
buf ( n46207 , n46111 );
buf ( n46208 , n46102 );
nand ( n46209 , n46207 , n46208 );
buf ( n46210 , n46209 );
and ( n46211 , n46210 , n454 );
not ( n46212 , n46211 );
buf ( n46213 , n46146 );
not ( n46214 , n46082 );
nor ( n46215 , n46214 , n45721 );
buf ( n46216 , n46215 );
buf ( n46217 , n44173 );
nand ( n46218 , n46213 , n46216 , n46217 );
buf ( n46219 , n46218 );
buf ( n46220 , n44193 );
buf ( n46221 , n46215 );
nand ( n46222 , n46220 , n46221 );
buf ( n46223 , n46222 );
buf ( n46224 , n46082 );
buf ( n46225 , n46224 );
buf ( n46226 , n46098 );
and ( n46227 , n46225 , n46226 );
buf ( n46228 , n45776 );
nor ( n46229 , n46227 , n46228 );
buf ( n46230 , n46229 );
nand ( n46231 , n46219 , n46223 , n46230 );
not ( n46232 , n46231 );
or ( n46233 , n46212 , n46232 );
not ( n46234 , n45577 );
not ( n46235 , n44669 );
or ( n46236 , n46234 , n46235 );
nand ( n46237 , n46236 , n45552 );
buf ( n46238 , n45432 );
buf ( n46239 , n45464 );
nand ( n46240 , n46238 , n46239 );
buf ( n46241 , n46240 );
not ( n46242 , n46241 );
and ( n46243 , n46237 , n46242 );
not ( n46244 , n46237 );
and ( n46245 , n46244 , n46241 );
nor ( n46246 , n46243 , n46245 );
nand ( n46247 , n46246 , n2356 );
nand ( n46248 , n46233 , n46247 );
buf ( n46249 , n46223 );
buf ( n46250 , n46219 );
buf ( n46251 , n46230 );
nand ( n46252 , n46249 , n46250 , n46251 );
buf ( n46253 , n46252 );
not ( n46254 , n46210 );
nand ( n46255 , n46254 , n454 );
nor ( n46256 , n46253 , n46255 );
nor ( n46257 , n46248 , n46256 );
not ( n46258 , n46257 );
not ( n46259 , n2356 );
buf ( n46260 , n45408 );
buf ( n46261 , n45587 );
xnor ( n46262 , n46260 , n46261 );
buf ( n46263 , n46262 );
not ( n46264 , n46263 );
or ( n46265 , n46259 , n46264 );
nand ( n46266 , n46146 , n45722 , n44173 );
and ( n46267 , n46266 , n45725 );
not ( n46268 , n45776 );
not ( n46269 , n46098 );
and ( n46270 , n46224 , n46268 , n46269 , n454 );
and ( n46271 , n46267 , n46270 );
nand ( n46272 , n46266 , n45725 , n46269 );
and ( n46273 , n46224 , n46268 );
nor ( n46274 , n46273 , n2618 );
and ( n46275 , n46272 , n46274 );
nor ( n46276 , n46271 , n46275 );
nand ( n46277 , n46265 , n46276 );
nand ( n46278 , n46258 , n46277 );
nor ( n46279 , n46206 , n46278 );
not ( n46280 , n2356 );
not ( n46281 , n45500 );
nand ( n46282 , n44656 , n41640 );
or ( n46283 , n46282 , n45568 );
nand ( n46284 , n46281 , n46283 );
not ( n46285 , n45519 );
nor ( n46286 , n46285 , n45507 );
xor ( n46287 , n46284 , n46286 );
not ( n46288 , n46287 );
or ( n46289 , n46280 , n46288 );
not ( n46290 , n46149 );
not ( n46291 , n46148 );
not ( n46292 , n46137 );
not ( n46293 , n46292 );
nand ( n46294 , n46291 , n46293 );
not ( n46295 , n46294 );
or ( n46296 , n46290 , n46295 );
nand ( n46297 , n46296 , n454 );
nand ( n46298 , n46289 , n46297 );
nand ( n46299 , n43794 , n43791 , n43956 );
and ( n46300 , n43498 , n46299 );
not ( n46301 , n454 );
not ( n46302 , n46152 );
or ( n46303 , n46301 , n46302 );
not ( n46304 , n45416 );
not ( n46305 , n45573 );
or ( n46306 , n46304 , n46305 );
nand ( n46307 , n46306 , n45549 );
nand ( n46308 , n46307 , n2356 );
nand ( n46309 , n46303 , n46308 );
nand ( n46310 , n46298 , n46300 , n46309 );
not ( n46311 , n2356 );
not ( n46312 , n45635 );
or ( n46313 , n46311 , n46312 );
nand ( n46314 , n46152 , n454 );
nand ( n46315 , n46313 , n46314 );
nand ( n46316 , n44679 , n44738 );
not ( n46317 , n46316 );
nand ( n46318 , n46315 , n46317 );
nor ( n46319 , n46310 , n46318 );
not ( n46320 , n40947 );
nand ( n46321 , n46320 , n41082 , n41652 );
not ( n46322 , n46321 );
nand ( n46323 , n46279 , n46319 , n46322 );
not ( n46324 , n46314 );
buf ( n46325 , n46324 );
not ( n46326 , n45984 );
not ( n46327 , n45930 );
or ( n46328 , n46326 , n46327 );
nand ( n46329 , n46328 , n45962 );
xor ( n46330 , n45990 , n46329 );
not ( n46331 , n45963 );
not ( n46332 , n45984 );
not ( n46333 , n45930 );
or ( n46334 , n46332 , n46333 );
nand ( n46335 , n46334 , n45962 );
not ( n46336 , n46335 );
or ( n46337 , n46331 , n46336 );
nand ( n46338 , n46337 , n45969 );
not ( n46339 , n6916 );
not ( n46340 , n7041 );
or ( n46341 , n46339 , n46340 );
not ( n46342 , n7048 );
nand ( n46343 , n46341 , n46342 );
and ( n46344 , n46343 , n7045 );
not ( n46345 , n46343 );
and ( n46346 , n46345 , n6963 );
nor ( n46347 , n46344 , n46346 );
buf ( n46348 , n46277 );
not ( n46349 , n44741 );
or ( n46350 , n46330 , n2629 );
and ( n46351 , n42171 , n46299 );
not ( n46352 , n454 );
not ( n46353 , n44724 );
and ( n46354 , n44730 , n46353 );
not ( n46355 , n44730 );
and ( n46356 , n46355 , n44724 );
nor ( n46357 , n46354 , n46356 );
not ( n46358 , n46357 );
or ( n46359 , n46352 , n46358 );
nand ( n46360 , n44707 , n2356 );
nand ( n46361 , n46359 , n46360 );
nand ( n46362 , n46315 , n46351 , n46361 );
not ( n46363 , n2356 );
not ( n46364 , n46287 );
or ( n46365 , n46363 , n46364 );
nand ( n46366 , n46365 , n46297 );
or ( n46367 , n44410 , n44197 );
or ( n46368 , n44198 , n44412 );
nand ( n46369 , n46367 , n46368 );
nand ( n46370 , n46369 , n44678 );
nand ( n46371 , n46366 , n46370 );
nor ( n46372 , n46362 , n46371 );
nand ( n46373 , n46372 , n46279 , n46322 );
not ( n46374 , n46309 );
nand ( n46375 , n46374 , n7410 );
or ( n46376 , n46373 , n46375 );
nor ( n46377 , n46374 , n2628 );
nand ( n46378 , n46373 , n46377 );
nand ( n46379 , n46350 , n46376 , n46378 );
not ( n46380 , n46178 );
nand ( n46381 , n46277 , n46205 );
not ( n46382 , n46381 );
nand ( n46383 , n44740 , n46382 , n41654 , n46258 );
not ( n46384 , n46383 );
nand ( n46385 , n46380 , n46384 , n7410 );
and ( n46386 , n46366 , n7410 );
nor ( n46387 , n46348 , n2628 );
buf ( n46388 , n46205 );
nand ( n46389 , n46388 , n41654 , n44740 );
or ( n46390 , n46387 , n46389 );
not ( n46391 , n7410 );
not ( n46392 , n46348 );
or ( n46393 , n46391 , n46392 );
nand ( n46394 , n46393 , n46389 );
nand ( n46395 , n46390 , n46394 );
nand ( n46396 , n46395 , n43447 );
and ( n46397 , n46325 , n2627 );
not ( n46398 , n46258 );
nand ( n46399 , n44740 , n46382 , n41654 );
not ( n46400 , n46399 );
nand ( n46401 , n46400 , n46398 , n7410 );
not ( n46402 , n7410 );
nor ( n46403 , n46402 , n46398 );
nand ( n46404 , n46403 , n46399 );
nand ( n46405 , n46401 , n43381 , n46404 );
buf ( n46406 , n43358 );
nand ( n46407 , n46351 , n46361 );
and ( n46408 , n41654 , n44740 );
not ( n46409 , n43348 );
not ( n46410 , n45941 );
or ( n46411 , n46409 , n46410 );
nand ( n46412 , n46411 , n46406 );
not ( n46413 , n43306 );
nand ( n46414 , n43321 , n43364 );
nor ( n46415 , n46413 , n46414 );
nand ( n46416 , n46412 , n46415 );
not ( n46417 , n46414 );
not ( n46418 , n43360 );
and ( n46419 , n46417 , n46418 );
not ( n46420 , n43306 );
nand ( n46421 , n46420 , n46414 , n43360 );
nand ( n46422 , n46421 , n2628 );
nor ( n46423 , n46419 , n46422 );
not ( n46424 , n46278 );
buf ( n46425 , n42171 );
not ( n46426 , n43957 );
not ( n46427 , n454 );
not ( n46428 , n41446 );
or ( n46429 , n46427 , n46428 );
nand ( n46430 , n46429 , n41651 );
nand ( n46431 , n46425 , n46426 , n46430 );
nand ( n46432 , n42881 , n42879 );
nor ( n46433 , n46431 , n46432 );
xor ( n46434 , n45982 , n46412 );
or ( n46435 , n46434 , n2629 );
not ( n46436 , n46407 );
not ( n46437 , n46436 );
not ( n46438 , n46322 );
or ( n46439 , n46437 , n46438 );
nand ( n46440 , n44411 , n44413 , n44678 );
and ( n46441 , n46440 , n2629 );
nand ( n46442 , n46439 , n46441 );
not ( n46443 , n46440 );
nand ( n46444 , n46443 , n46322 , n2629 , n46436 );
nand ( n46445 , n46435 , n46442 , n46444 );
not ( n46446 , n46412 );
nand ( n46447 , n46446 , n46414 , n43360 );
nand ( n46448 , n46447 , n46423 , n46416 );
not ( n46449 , n46206 );
nor ( n46450 , n7027 , n471 );
nand ( n46451 , n46349 , n46388 );
not ( n46452 , n46388 );
nand ( n46453 , n46452 , n44741 );
nand ( n46454 , n46451 , n46453 , n7410 );
nand ( n46455 , n46454 , n46448 );
and ( n46456 , n46152 , n454 );
and ( n46457 , n46456 , n7410 );
not ( n46458 , n46457 );
and ( n46459 , n41082 , n40948 , n41652 );
and ( n46460 , n43498 , n46299 );
and ( n46461 , n46317 , n46460 );
nand ( n46462 , n46449 , n46424 , n46459 , n46461 );
not ( n46463 , n46462 );
or ( n46464 , n46458 , n46463 );
nand ( n46465 , n45999 , n45966 );
not ( n46466 , n46465 );
nand ( n46467 , n46466 , n45984 );
not ( n46468 , n46467 );
and ( n46469 , n45920 , n46468 , n43374 );
or ( n46470 , n45929 , n46467 );
not ( n46471 , n45962 );
not ( n46472 , n46465 );
and ( n46473 , n46471 , n46472 );
not ( n46474 , n45999 );
nor ( n46475 , n46474 , n45974 );
nor ( n46476 , n46473 , n46475 );
nand ( n46477 , n46470 , n46476 );
nor ( n46478 , n46469 , n46477 );
not ( n46479 , n46478 );
not ( n46480 , n45966 );
not ( n46481 , n46335 );
or ( n46482 , n46480 , n46481 );
not ( n46483 , n45974 );
nor ( n46484 , n46483 , n45999 );
nand ( n46485 , n46482 , n46484 );
not ( n46486 , n46485 );
or ( n46487 , n46479 , n46486 );
nand ( n46488 , n46487 , n2628 );
nand ( n46489 , n46464 , n46488 );
nand ( n46490 , n46315 , n2627 );
not ( n46491 , n46490 );
not ( n46492 , n46490 );
nor ( n46493 , n46492 , n46459 );
nor ( n46494 , n46491 , n46382 );
and ( n46495 , n46324 , n46258 , n46277 );
and ( n46496 , n42881 , n46430 , n42879 , n42908 );
nand ( n46497 , n46495 , n46449 , n46496 );
not ( n46498 , n46491 );
nand ( n46499 , n46160 , n2356 );
nand ( n46500 , n46499 , n46176 );
and ( n46501 , n46258 , n46500 );
nand ( n46502 , n46298 , n46440 );
nor ( n46503 , n46502 , n46407 );
nand ( n46504 , n46501 , n46503 );
nand ( n46505 , n46498 , n46504 );
not ( n46506 , n46315 );
not ( n46507 , n2627 );
not ( n46508 , n46507 );
and ( n46509 , n46506 , n46508 );
nor ( n46510 , n46509 , n46381 );
nand ( n46511 , n46501 , n46510 , n46503 , n46459 );
nor ( n46512 , n46493 , n46494 );
nand ( n46513 , n46505 , n46511 , n46512 );
not ( n46514 , n45989 );
not ( n46515 , n45934 );
or ( n46516 , n46514 , n46515 );
or ( n46517 , n45934 , n45989 );
nand ( n46518 , n46516 , n46517 );
nand ( n46519 , n46518 , n2628 );
nand ( n46520 , n46513 , n46519 );
and ( n46521 , n7028 , n7022 );
and ( n46522 , n7027 , n471 );
nor ( n46523 , n46522 , n7022 );
nor ( n46524 , n46521 , n46523 );
not ( n46525 , n46524 );
not ( n46526 , n7032 );
and ( n46527 , n7022 , n46526 );
not ( n46528 , n7022 );
and ( n46529 , n46528 , n46450 );
nor ( n46530 , n46527 , n46529 );
nand ( n46531 , n46525 , n46530 );
and ( n46532 , n46531 , n2627 );
and ( n46533 , n46032 , n2628 );
nor ( n46534 , n46532 , n46533 );
and ( n46535 , n44761 , n2627 );
and ( n46536 , n2628 , n46033 );
nor ( n46537 , n46535 , n46536 );
not ( n46538 , n46537 );
and ( n46539 , n46323 , n46397 );
nor ( n46540 , n46539 , C0 );
and ( n46541 , n45991 , n2628 );
and ( n46542 , n46338 , n46541 );
not ( n46543 , n46338 );
nor ( n46544 , n45991 , n2627 );
and ( n46545 , n46543 , n46544 );
nor ( n46546 , n46542 , n46545 );
nand ( n46547 , n46540 , n46546 );
nand ( n46548 , n46462 , n46457 );
not ( n46549 , n46548 );
buf ( n46550 , n44738 );
not ( n46551 , n46550 );
nand ( n46552 , n46551 , n43450 );
not ( n46553 , n43450 );
nand ( n46554 , n46553 , n46433 , n46550 );
not ( n46555 , n46433 );
and ( n46556 , n46555 , n46551 );
nor ( n46557 , n46556 , n2628 );
nand ( n46558 , n46552 , n46554 , n46557 );
nand ( n46559 , n45948 , n2628 );
nand ( n46560 , n46558 , n46559 );
nand ( n46561 , n46178 , n46383 , n7410 );
nand ( n46562 , n46385 , n46561 , n43443 );
nand ( n46563 , n41054 , n41079 );
not ( n46564 , n46366 );
nand ( n46565 , n46564 , n7410 );
nand ( n46566 , n46408 , n46279 );
or ( n46567 , n46565 , n46566 );
xor ( n46568 , n45988 , n46153 );
or ( n46569 , n46568 , n7410 );
nand ( n46570 , n46566 , n46386 );
nand ( n46571 , n46567 , n46569 , n46570 );
and ( n46572 , n46317 , n46300 );
buf ( n46573 , n46456 );
nor ( n46574 , n2628 , n46430 );
and ( n46575 , n36964 , n42908 , n42881 );
not ( n46576 , n42879 );
nor ( n46577 , n46576 , n42884 );
nand ( n46578 , n46574 , n46575 , n46577 );
not ( n46579 , n46577 );
not ( n46580 , n46575 );
or ( n46581 , n46579 , n46580 );
not ( n46582 , n46430 );
nor ( n46583 , n46582 , n2628 );
nand ( n46584 , n46581 , n46583 );
not ( n46585 , n42599 );
not ( n46586 , n42894 );
or ( n46587 , n46585 , n46586 );
not ( n46588 , n42592 );
nand ( n46589 , n46587 , n46588 );
not ( n46590 , n46589 );
nor ( n46591 , n42595 , n42490 );
and ( n46592 , n46590 , n46591 );
nor ( n46593 , n42594 , n42552 );
and ( n46594 , n46590 , n46593 );
nor ( n46595 , n46592 , n46594 );
and ( n46596 , n46589 , n42597 );
not ( n46597 , n42553 );
and ( n46598 , n46589 , n46597 );
nor ( n46599 , n46596 , n46598 );
nand ( n46600 , n46595 , n46599 );
nand ( n46601 , n46600 , n2628 );
nand ( n46602 , n46578 , n46584 , n46601 );
not ( n46603 , n46425 );
not ( n46604 , n46322 );
or ( n46605 , n46603 , n46604 );
not ( n46606 , n46426 );
nor ( n46607 , n46606 , n2628 );
nand ( n46608 , n46605 , n46607 );
and ( n46609 , n42171 , n7410 );
and ( n46610 , n46609 , n46322 , n43957 );
and ( n46611 , n2628 , n45954 );
nor ( n46612 , n46610 , n46611 );
nand ( n46613 , n46608 , n46612 );
not ( n46614 , n2627 );
not ( n46615 , n44757 );
or ( n46616 , n46614 , n46615 );
nand ( n46617 , n46028 , n2628 );
nand ( n46618 , n46616 , n46617 );
not ( n46619 , n2629 );
not ( n46620 , n40975 );
nand ( n46621 , n36964 , n36959 );
not ( n46622 , n46621 );
or ( n46623 , n46620 , n46622 );
or ( n46624 , n40975 , n46621 );
nand ( n46625 , n46623 , n46624 );
not ( n46626 , n46625 );
or ( n46627 , n46619 , n46626 );
nand ( n46628 , n45987 , n2628 );
nand ( n46629 , n46627 , n46628 );
not ( n46630 , n2629 );
not ( n46631 , n44751 );
or ( n46632 , n46630 , n46631 );
nand ( n46633 , n46051 , n2628 );
nand ( n46634 , n46632 , n46633 );
not ( n46635 , n2629 );
not ( n46636 , n46347 );
or ( n46637 , n46635 , n46636 );
nand ( n46638 , n45997 , n2628 );
nand ( n46639 , n46637 , n46638 );
not ( n46640 , n454 );
not ( n46641 , n45655 );
or ( n46642 , n46640 , n46641 );
nand ( n46643 , n45606 , n2618 );
nand ( n46644 , n46642 , n46643 );
not ( n46645 , n454 );
not ( n46646 , n45669 );
or ( n46647 , n46645 , n46646 );
nand ( n46648 , n45614 , n2618 );
nand ( n46649 , n46647 , n46648 );
not ( n46650 , n42907 );
nand ( n46651 , n46650 , n46572 );
nor ( n46652 , n46651 , n46497 , n2628 );
not ( n46653 , n46534 );
not ( n46654 , n2618 );
not ( n46655 , n45627 );
or ( n46656 , n46654 , n46655 );
nand ( n46657 , n45734 , n454 );
nand ( n46658 , n46656 , n46657 );
not ( n46659 , n454 );
not ( n46660 , n45732 );
or ( n46661 , n46659 , n46660 );
nand ( n46662 , n45617 , n2618 );
nand ( n46663 , n46661 , n46662 );
not ( n46664 , n46457 );
not ( n46665 , n46462 );
or ( n46666 , n46664 , n46665 );
not ( n46667 , n45930 );
not ( n46668 , n45985 );
or ( n46669 , n46667 , n46668 );
nand ( n46670 , n46669 , n45981 );
and ( n46671 , n46670 , n46011 );
not ( n46672 , n46670 );
not ( n46673 , n46011 );
and ( n46674 , n46672 , n46673 );
nor ( n46675 , n46671 , n46674 );
nand ( n46676 , n46675 , n2628 );
nand ( n46677 , n46666 , n46676 );
not ( n46678 , n42926 );
nor ( n46679 , n42926 , n46563 );
nand ( n46680 , n36966 , n46678 );
nand ( n46681 , n36966 , n46679 );
not ( n46682 , n46154 );
not ( n46683 , n7042 );
or ( n46684 , n46682 , n46683 );
or ( n46685 , n46154 , n7042 );
nand ( n46686 , n46684 , n46685 );
not ( n46687 , n45956 );
not ( n46688 , n2628 );
or ( n46689 , n46687 , n46688 );
nand ( n46690 , n46689 , n43456 );
and ( n46691 , n2627 , n46686 );
not ( n46692 , n2627 );
and ( n46693 , n46692 , n46018 );
or ( n46694 , n46691 , n46693 );
xor ( n46695 , n42749 , n42751 );
xor ( n46696 , n46695 , n42770 );
or ( n46697 , n46681 , n2628 );
and ( n46698 , n41080 , n7410 );
nand ( n46699 , n46680 , n46698 );
nand ( n46700 , n46696 , n2628 );
nand ( n46701 , n46697 , n46699 , n46700 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
not ( C1n , n0 );
or ( C1 , C1n , n0 );
endmodule
