module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 ;
output g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
     n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
     n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
     n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
     n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
     n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
     n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
     n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
     n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
     n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
     n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
     n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
     n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
     n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
     n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
     n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
     n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
     n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
     n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
     n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
     n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
     n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
     n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
     n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
     n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , 
     n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , 
     n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , 
     n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , 
     n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
     n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , 
     n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
     n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
     n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
     n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
     n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
     n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
     n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
     n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
     n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , 
     n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , 
     n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
     n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
     n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
     n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
     n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , 
     n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , 
     n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , 
     n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
     n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
     n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
     n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
     n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
     n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
     n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , 
     n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , 
     n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , 
     n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , 
     n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , 
     n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
     n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
     n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
     n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
     n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , 
     n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , 
     n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , 
     n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , 
     n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , 
     n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
     n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , 
     n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , 
     n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , 
     n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , 
     n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , 
     n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , 
     n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , 
     n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , 
     n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , 
     n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , 
     n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , 
     n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , 
     n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , 
     n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , 
     n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , 
     n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , 
     n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
     n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , 
     n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , 
     n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , 
     n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , 
     n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , 
     n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , 
     n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , 
     n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , 
     n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , 
     n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , 
     n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , 
     n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , 
     n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , 
     n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , 
     n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , 
     n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , 
     n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , 
     n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , 
     n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , 
     n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , 
     n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , 
     n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , 
     n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , 
     n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , 
     n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , 
     n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , 
     n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , 
     n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , 
     n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , 
     n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , 
     n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , 
     n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , 
     n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , 
     n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , 
     n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , 
     n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , 
     n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , 
     n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , 
     n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , 
     n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , 
     n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , 
     n3270 , n3271 , n3272 , n3273 , n3274 , n3275 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( n18 , g17 );
buf ( n19 , g18 );
buf ( n20 , g19 );
buf ( n21 , g20 );
buf ( n22 , g21 );
buf ( n23 , g22 );
buf ( n24 , g23 );
buf ( n25 , g24 );
buf ( n26 , g25 );
buf ( n27 , g26 );
buf ( n28 , g27 );
buf ( n29 , g28 );
buf ( n30 , g29 );
buf ( n31 , g30 );
buf ( n32 , g31 );
buf ( n33 , g32 );
buf ( n34 , g33 );
buf ( n35 , g34 );
buf ( n36 , g35 );
buf ( n37 , g36 );
buf ( n38 , g37 );
buf ( n39 , g38 );
buf ( n40 , g39 );
buf ( n41 , g40 );
buf ( n42 , g41 );
buf ( n43 , g42 );
buf ( n44 , g43 );
buf ( n45 , g44 );
buf ( n46 , g45 );
buf ( n47 , g46 );
buf ( n48 , g47 );
buf ( n49 , g48 );
buf ( n50 , g49 );
buf ( n51 , g50 );
buf ( n52 , g51 );
buf ( n53 , g52 );
buf ( n54 , g53 );
buf ( n55 , g54 );
buf ( n56 , g55 );
buf ( n57 , g56 );
buf ( n58 , g57 );
buf ( n59 , g58 );
buf ( n60 , g59 );
buf ( n61 , g60 );
buf ( n62 , g61 );
buf ( n63 , g62 );
buf ( n64 , g63 );
buf ( n65 , g64 );
buf ( n66 , g65 );
buf ( n67 , g66 );
buf ( n68 , g67 );
buf ( n69 , g68 );
buf ( n70 , g69 );
buf ( n71 , g70 );
buf ( n72 , g71 );
buf ( n73 , g72 );
buf ( n74 , g73 );
buf ( n75 , g74 );
buf ( n76 , g75 );
buf ( n77 , g76 );
buf ( n78 , g77 );
buf ( n79 , g78 );
buf ( n80 , g79 );
buf ( n81 , g80 );
buf ( n82 , g81 );
buf ( n83 , g82 );
buf ( n84 , g83 );
buf ( n85 , g84 );
buf ( n86 , g85 );
buf ( n87 , g86 );
buf ( n88 , g87 );
buf ( n89 , g88 );
buf ( n90 , g89 );
buf ( n91 , g90 );
buf ( n92 , g91 );
buf ( n93 , g92 );
buf ( n94 , g93 );
buf ( n95 , g94 );
buf ( n96 , g95 );
buf ( n97 , g96 );
buf ( n98 , g97 );
buf ( n99 , g98 );
buf ( n100 , g99 );
buf ( n101 , g100 );
buf ( n102 , g101 );
buf ( n103 , g102 );
buf ( n104 , g103 );
buf ( n105 , g104 );
buf ( n106 , g105 );
buf ( n107 , g106 );
buf ( n108 , g107 );
buf ( n109 , g108 );
buf ( n110 , g109 );
buf ( n111 , g110 );
buf ( n112 , g111 );
buf ( n113 , g112 );
buf ( n114 , g113 );
buf ( n115 , g114 );
buf ( n116 , g115 );
buf ( n117 , g116 );
buf ( n118 , g117 );
buf ( n119 , g118 );
buf ( n120 , g119 );
buf ( n121 , g120 );
buf ( n122 , g121 );
buf ( n123 , g122 );
buf ( n124 , g123 );
buf ( n125 , g124 );
buf ( n126 , g125 );
buf ( n127 , g126 );
buf ( n128 , g127 );
buf ( n129 , g128 );
buf ( n130 , g129 );
buf ( n131 , g130 );
buf ( n132 , g131 );
buf ( n133 , g132 );
buf ( n134 , g133 );
buf ( n135 , g134 );
buf ( n136 , g135 );
buf ( n137 , g136 );
buf ( n138 , g137 );
buf ( n139 , g138 );
buf ( n140 , g139 );
buf ( n141 , g140 );
buf ( n142 , g141 );
buf ( n143 , g142 );
buf ( n144 , g143 );
buf ( n145 , g144 );
buf ( n146 , g145 );
buf ( n147 , g146 );
buf ( n148 , g147 );
buf ( n149 , g148 );
buf ( n150 , g149 );
buf ( n151 , g150 );
buf ( n152 , g151 );
buf ( n153 , g152 );
buf ( n154 , g153 );
buf ( n155 , g154 );
buf ( n156 , g155 );
buf ( n157 , g156 );
buf ( n158 , g157 );
buf ( n159 , g158 );
buf ( n160 , g159 );
buf ( n161 , g160 );
buf ( n162 , g161 );
buf ( n163 , g162 );
buf ( n164 , g163 );
buf ( n165 , g164 );
buf ( n166 , g165 );
buf ( n167 , g166 );
buf ( n168 , g167 );
buf ( n169 , g168 );
buf ( n170 , g169 );
buf ( n171 , g170 );
buf ( n172 , g171 );
buf ( n173 , g172 );
buf ( n174 , g173 );
buf ( n175 , g174 );
buf ( n176 , g175 );
buf ( n177 , g176 );
buf ( n178 , g177 );
buf ( n179 , g178 );
buf ( g179 , n180 );
buf ( g180 , n181 );
buf ( g181 , n182 );
buf ( g182 , n183 );
buf ( g183 , n184 );
buf ( g184 , n185 );
buf ( g185 , n186 );
buf ( g186 , n187 );
buf ( g187 , n188 );
buf ( g188 , n189 );
buf ( g189 , n190 );
buf ( g190 , n191 );
buf ( g191 , n192 );
buf ( g192 , n193 );
buf ( g193 , n194 );
buf ( g194 , n195 );
buf ( g195 , n196 );
buf ( g196 , n197 );
buf ( g197 , n198 );
buf ( g198 , n199 );
buf ( g199 , n200 );
buf ( g200 , n201 );
buf ( g201 , n202 );
buf ( g202 , n203 );
buf ( g203 , n204 );
buf ( g204 , n205 );
buf ( g205 , n206 );
buf ( g206 , n207 );
buf ( g207 , n208 );
buf ( g208 , n209 );
buf ( g209 , n210 );
buf ( g210 , n211 );
buf ( g211 , n212 );
buf ( g212 , n213 );
buf ( g213 , n214 );
buf ( g214 , n215 );
buf ( g215 , n216 );
buf ( g216 , n217 );
buf ( g217 , n218 );
buf ( g218 , n219 );
buf ( g219 , n220 );
buf ( g220 , n221 );
buf ( g221 , n222 );
buf ( g222 , n223 );
buf ( g223 , n224 );
buf ( g224 , n225 );
buf ( g225 , n226 );
buf ( g226 , n227 );
buf ( g227 , n228 );
buf ( g228 , n229 );
buf ( g229 , n230 );
buf ( g230 , n231 );
buf ( g231 , n232 );
buf ( g232 , n233 );
buf ( g233 , n234 );
buf ( g234 , n235 );
buf ( g235 , n236 );
buf ( g236 , n237 );
buf ( g237 , n238 );
buf ( g238 , n239 );
buf ( g239 , n240 );
buf ( g240 , n241 );
buf ( g241 , n242 );
buf ( g242 , n243 );
buf ( n180 , n2610 );
buf ( n181 , n2627 );
buf ( n182 , n2719 );
buf ( n183 , n2733 );
buf ( n184 , n3137 );
buf ( n185 , n2846 );
buf ( n186 , n3154 );
buf ( n187 , n1883 );
buf ( n188 , n1951 );
buf ( n189 , n2084 );
buf ( n190 , n2015 );
buf ( n191 , n2215 );
buf ( n192 , n2266 );
buf ( n193 , n2144 );
buf ( n194 , n2469 );
buf ( n195 , n2533 );
buf ( n196 , n2895 );
buf ( n197 , n1893 );
buf ( n198 , n2021 );
buf ( n199 , n2149 );
buf ( n200 , n2024 );
buf ( n201 , n2220 );
buf ( n202 , n2271 );
buf ( n203 , n2152 );
buf ( n204 , n2557 );
buf ( n205 , n2553 );
buf ( n206 , n2899 );
buf ( n207 , n2973 );
buf ( n208 , n2421 );
buf ( n209 , n2706 );
buf ( n210 , n3086 );
buf ( n211 , n2365 );
buf ( n212 , n2344 );
buf ( n213 , n2549 );
buf ( n214 , n2573 );
buf ( n215 , n2640 );
buf ( n216 , n2657 );
buf ( n217 , n2831 );
buf ( n218 , n3049 );
buf ( n219 , n2923 );
buf ( n220 , n2992 );
buf ( n221 , n2912 );
buf ( n222 , n3105 );
buf ( n223 , n3246 );
buf ( n224 , n2800 );
buf ( n225 , n2997 );
buf ( n226 , n3192 );
buf ( n227 , n2797 );
buf ( n228 , n3197 );
buf ( n229 , n3012 );
buf ( n230 , n3171 );
buf ( n231 , n3236 );
buf ( n232 , n2939 );
buf ( n233 , n3121 );
buf ( n234 , n3214 );
buf ( n235 , n2426 );
buf ( n236 , n2804 );
buf ( n237 , n3125 );
buf ( n238 , n2816 );
buf ( n239 , n3026 );
buf ( n240 , n3226 );
buf ( n241 , n3275 );
buf ( n242 , n3253 );
buf ( n243 , n3270 );
not ( n246 , n80 );
not ( n247 , n1 );
not ( n248 , n22 );
and ( n249 , n247 , n248 );
not ( n250 , n247 );
nor ( n251 , n29 , n30 );
nor ( n252 , n19 , n28 );
nor ( n253 , n18 , n31 );
nor ( n254 , n20 , n32 );
nand ( n255 , n251 , n252 , n253 , n254 );
not ( n256 , n255 );
nor ( n257 , n6 , n7 );
nor ( n258 , n4 , n12 );
nor ( n259 , n5 , n13 );
and ( n260 , n257 , n258 , n259 );
nor ( n261 , n2 , n11 );
nor ( n262 , n8 , n14 );
nor ( n263 , n9 , n16 );
nand ( n264 , n262 , n263 );
not ( n265 , n264 );
nor ( n266 , n3 , n10 );
nor ( n267 , n15 , n17 );
nand ( n268 , n266 , n267 );
not ( n269 , n268 );
nand ( n270 , n260 , n261 , n265 , n269 );
not ( n271 , n270 );
nand ( n272 , n256 , n271 );
and ( n273 , n272 , n248 );
not ( n274 , n272 );
and ( n275 , n274 , n22 );
nor ( n276 , n273 , n275 );
and ( n277 , n250 , n276 );
or ( n278 , n249 , n277 );
not ( n279 , n27 );
not ( n280 , n26 );
not ( n281 , n25 );
not ( n282 , n24 );
not ( n283 , n23 );
nor ( n284 , n21 , n22 );
nand ( n285 , n282 , n283 , n284 );
nor ( n286 , n285 , n255 );
nand ( n287 , n280 , n281 , n286 , n271 );
not ( n288 , n287 );
and ( n289 , n1 , n279 , n288 );
not ( n290 , n289 );
not ( n291 , n290 );
not ( n292 , n291 );
not ( n293 , n1 );
and ( n294 , n293 , n31 );
not ( n295 , n293 );
not ( n296 , n270 );
nor ( n297 , n20 , n29 );
nor ( n298 , n18 , n19 );
nand ( n299 , n296 , n297 , n298 );
not ( n300 , n299 );
not ( n301 , n30 );
not ( n302 , n28 );
not ( n303 , n32 );
and ( n304 , n302 , n303 );
nand ( n305 , n300 , n301 , n304 );
not ( n306 , n31 );
and ( n307 , n305 , n306 );
not ( n308 , n305 );
and ( n309 , n308 , n31 );
nor ( n310 , n307 , n309 );
not ( n311 , n310 );
and ( n312 , n295 , n311 );
nor ( n313 , n294 , n312 );
buf ( n314 , n313 );
nor ( n315 , n292 , n314 );
not ( n316 , n292 );
not ( n317 , n316 );
not ( n318 , n1 );
and ( n319 , n318 , n30 );
not ( n320 , n318 );
nor ( n321 , n264 , n268 );
nand ( n322 , n260 , n261 , n321 );
not ( n323 , n322 );
nand ( n324 , n323 , n298 , n297 );
not ( n325 , n324 );
nand ( n326 , n304 , n325 );
xnor ( n327 , n326 , n30 );
not ( n328 , n327 );
and ( n329 , n320 , n328 );
nor ( n330 , n319 , n329 );
not ( n331 , n1 );
and ( n332 , n331 , n28 );
not ( n333 , n331 );
not ( n334 , n324 );
nand ( n335 , n334 , n303 );
and ( n336 , n335 , n302 );
not ( n337 , n335 );
and ( n338 , n337 , n28 );
nor ( n339 , n336 , n338 );
not ( n340 , n339 );
and ( n341 , n333 , n340 );
nor ( n342 , n332 , n341 );
not ( n343 , n29 );
not ( n344 , n1 );
not ( n345 , n344 );
or ( n346 , n343 , n345 );
not ( n347 , n20 );
not ( n348 , n347 );
not ( n349 , n322 );
nand ( n350 , n349 , n298 );
not ( n351 , n350 );
not ( n352 , n351 );
or ( n353 , n348 , n352 );
nand ( n354 , n353 , n29 );
not ( n355 , n29 );
nor ( n356 , n20 , n350 );
and ( n357 , n355 , n356 );
not ( n358 , n1 );
nor ( n359 , n357 , n358 );
nand ( n360 , n354 , n359 );
nand ( n361 , n346 , n360 );
not ( n362 , n299 );
not ( n363 , n362 );
not ( n364 , n32 );
and ( n365 , n363 , n364 );
and ( n366 , n32 , n362 );
nor ( n367 , n365 , n366 );
not ( n368 , n1 );
or ( n369 , n367 , n368 );
or ( n370 , n303 , n1 );
nand ( n371 , n369 , n370 );
nor ( n372 , n361 , n371 );
nand ( n373 , n330 , n342 , n372 );
not ( n374 , n373 );
or ( n375 , n317 , n374 );
not ( n376 , n9 );
not ( n377 , n8 );
nor ( n378 , n6 , n7 );
nand ( n379 , n376 , n377 , n378 );
nand ( n380 , n379 , n1 );
xor ( n381 , n380 , n2 );
not ( n382 , n381 );
not ( n383 , n382 );
not ( n384 , n6 );
nand ( n385 , n377 , n378 );
nand ( n386 , n1 , n385 );
and ( n387 , n386 , n376 );
not ( n388 , n386 );
and ( n389 , n388 , n9 );
or ( n390 , n387 , n389 );
and ( n391 , n384 , n390 );
not ( n392 , n10 );
not ( n393 , n2 );
not ( n394 , n3 );
nand ( n395 , n393 , n394 );
nand ( n396 , n376 , n377 , n257 );
nor ( n397 , n395 , n396 );
nor ( n398 , n4 , n5 );
nand ( n399 , n397 , n398 );
nor ( n400 , n11 , n399 );
not ( n401 , n400 );
or ( n402 , n392 , n401 );
not ( n403 , n379 );
not ( n404 , n395 );
nand ( n405 , n403 , n398 , n404 );
not ( n406 , n405 );
not ( n407 , n406 );
nor ( n408 , n407 , n11 );
or ( n409 , n10 , n408 );
nand ( n410 , n402 , n409 );
and ( n411 , n1 , n410 );
not ( n412 , n1 );
and ( n413 , n412 , n10 );
nor ( n414 , n411 , n413 );
nand ( n415 , n383 , n391 , n414 );
not ( n416 , n415 );
not ( n417 , n1 );
and ( n418 , n417 , n12 );
not ( n419 , n417 );
not ( n420 , n405 );
nor ( n421 , n10 , n11 );
not ( n422 , n13 );
nand ( n423 , n420 , n421 , n422 );
xor ( n424 , n423 , n12 );
and ( n425 , n419 , n424 );
nor ( n426 , n418 , n425 );
not ( n427 , n1 );
and ( n428 , n427 , n13 );
not ( n429 , n427 );
not ( n430 , n422 );
not ( n431 , n399 );
nand ( n432 , n421 , n431 );
not ( n433 , n432 );
and ( n434 , n430 , n433 );
and ( n435 , n422 , n432 );
nor ( n436 , n434 , n435 );
not ( n437 , n436 );
and ( n438 , n429 , n437 );
nor ( n439 , n428 , n438 );
not ( n440 , n1 );
not ( n441 , n6 );
not ( n442 , n7 );
or ( n443 , n441 , n442 );
nor ( n444 , n6 , n7 );
not ( n445 , n444 );
nand ( n446 , n443 , n445 );
or ( n447 , n440 , n446 );
not ( n448 , n1 );
nand ( n449 , n448 , n7 );
nand ( n450 , n447 , n449 );
not ( n451 , n450 );
not ( n452 , n1 );
nor ( n453 , n377 , n378 );
not ( n454 , n453 );
nand ( n455 , n454 , n385 );
or ( n456 , n452 , n455 );
not ( n457 , n1 );
nand ( n458 , n457 , n8 );
nand ( n459 , n456 , n458 );
not ( n460 , n459 );
and ( n461 , n451 , n460 );
nand ( n462 , n376 , n377 , n444 );
nor ( n463 , n395 , n462 );
not ( n464 , n463 );
nand ( n465 , n464 , n1 );
not ( n466 , n5 );
xor ( n467 , n465 , n466 );
not ( n468 , n467 );
not ( n469 , n4 );
not ( n470 , n1 );
not ( n471 , n470 );
or ( n472 , n469 , n471 );
not ( n473 , n4 );
and ( n474 , n466 , n463 );
not ( n475 , n474 );
not ( n476 , n475 );
or ( n477 , n473 , n476 );
not ( n478 , n4 );
and ( n479 , n478 , n474 );
not ( n480 , n1 );
nor ( n481 , n479 , n480 );
nand ( n482 , n477 , n481 );
nand ( n483 , n472 , n482 );
not ( n484 , n483 );
nand ( n485 , n461 , n468 , n484 );
not ( n486 , n445 );
nand ( n487 , n376 , n377 , n486 );
nor ( n488 , n2 , n487 );
not ( n489 , n488 );
nand ( n490 , n3 , n489 );
and ( n491 , n394 , n488 );
not ( n492 , n1 );
nor ( n493 , n491 , n492 );
and ( n494 , n490 , n493 );
nor ( n495 , n394 , n1 );
nor ( n496 , n494 , n495 );
not ( n497 , n496 );
not ( n498 , n11 );
not ( n499 , n1 );
not ( n500 , n499 );
or ( n501 , n498 , n500 );
not ( n502 , n408 );
nand ( n503 , n11 , n399 );
nand ( n504 , n502 , n503 , n1 );
not ( n505 , n504 );
not ( n506 , n505 );
nand ( n507 , n501 , n506 );
nor ( n508 , n485 , n497 , n507 );
nand ( n509 , n416 , n426 , n439 , n508 );
not ( n510 , n1 );
and ( n511 , n510 , n14 );
not ( n512 , n510 );
not ( n513 , n14 );
not ( n514 , n513 );
nor ( n515 , n10 , n11 );
not ( n516 , n12 );
nand ( n517 , n515 , n516 , n422 );
not ( n518 , n517 );
nand ( n519 , n518 , n431 );
not ( n520 , n519 );
and ( n521 , n514 , n520 );
and ( n522 , n513 , n519 );
nor ( n523 , n521 , n522 );
not ( n524 , n523 );
and ( n525 , n512 , n524 );
nor ( n526 , n511 , n525 );
not ( n527 , n1 );
and ( n528 , n527 , n16 );
not ( n529 , n527 );
not ( n530 , n399 );
nand ( n531 , n530 , n513 , n518 );
and ( n532 , n531 , n16 );
not ( n533 , n531 );
not ( n534 , n16 );
and ( n535 , n533 , n534 );
nor ( n536 , n532 , n535 );
and ( n537 , n529 , n536 );
nor ( n538 , n528 , n537 );
not ( n539 , n1 );
and ( n540 , n539 , n17 );
not ( n541 , n539 );
not ( n542 , n399 );
nand ( n543 , n513 , n534 );
nor ( n544 , n543 , n517 );
nand ( n545 , n542 , n544 );
and ( n546 , n545 , n17 );
not ( n547 , n545 );
not ( n548 , n17 );
and ( n549 , n547 , n548 );
nor ( n550 , n546 , n549 );
and ( n551 , n541 , n550 );
nor ( n552 , n540 , n551 );
nand ( n553 , n526 , n538 , n552 );
not ( n554 , n553 );
not ( n555 , n1 );
not ( n556 , n351 );
and ( n557 , n556 , n347 );
not ( n558 , n556 );
and ( n559 , n558 , n20 );
nor ( n560 , n557 , n559 );
nor ( n561 , n555 , n560 );
not ( n562 , n18 );
not ( n563 , n562 );
not ( n564 , n19 );
nand ( n565 , n564 , n271 );
not ( n566 , n565 );
or ( n567 , n563 , n566 );
and ( n568 , n261 , n376 , n534 );
not ( n569 , n10 );
not ( n570 , n15 );
and ( n571 , n394 , n569 , n570 , n548 );
nor ( n572 , n562 , n19 );
nor ( n573 , n8 , n14 );
and ( n574 , n258 , n259 );
and ( n575 , n573 , n486 , n574 );
nand ( n576 , n568 , n571 , n572 , n575 );
nand ( n577 , n567 , n576 );
not ( n578 , n577 );
and ( n579 , n1 , n578 );
not ( n580 , n1 );
and ( n581 , n347 , n580 , n562 );
nor ( n582 , n579 , n581 );
nor ( n583 , n561 , n582 );
not ( n584 , n1 );
not ( n585 , n399 );
nor ( n586 , n543 , n517 );
nand ( n587 , n585 , n586 , n548 );
and ( n588 , n587 , n15 );
not ( n589 , n587 );
and ( n590 , n589 , n570 );
nor ( n591 , n588 , n590 );
not ( n592 , n591 );
or ( n593 , n584 , n592 );
or ( n594 , n570 , n1 );
nand ( n595 , n593 , n594 );
nor ( n596 , n271 , n564 );
not ( n597 , n596 );
nand ( n598 , n597 , n1 , n565 );
not ( n599 , n598 );
nor ( n600 , n595 , n599 );
not ( n601 , n1 );
nand ( n602 , n19 , n601 );
nand ( n603 , n554 , n583 , n600 , n602 );
nor ( n604 , n509 , n603 );
nor ( n605 , n604 , n290 );
not ( n606 , n605 );
nand ( n607 , n375 , n606 );
nor ( n608 , n315 , n607 );
nor ( n609 , n278 , n608 );
not ( n610 , n609 );
nand ( n611 , n278 , n608 );
nand ( n612 , n610 , n611 );
not ( n613 , n612 );
not ( n614 , n613 );
not ( n615 , n159 );
not ( n616 , n615 );
not ( n617 , n1 );
and ( n618 , n617 , n21 );
not ( n619 , n617 );
not ( n620 , n21 );
nand ( n621 , n271 , n256 );
nor ( n622 , n22 , n621 );
not ( n623 , n622 );
or ( n624 , n620 , n623 );
nor ( n625 , n272 , n22 );
or ( n626 , n21 , n625 );
nand ( n627 , n624 , n626 );
and ( n628 , n619 , n627 );
nor ( n629 , n618 , n628 );
not ( n630 , n629 );
and ( n631 , n630 , n609 );
not ( n632 , n631 );
not ( n633 , n609 );
nand ( n634 , n629 , n633 );
nand ( n635 , n632 , n634 );
not ( n636 , n635 );
or ( n637 , n616 , n636 );
not ( n638 , n1 );
and ( n639 , n638 , n23 );
not ( n640 , n638 );
not ( n641 , n270 );
not ( n642 , n284 );
nor ( n643 , n29 , n30 );
nor ( n644 , n19 , n28 );
nor ( n645 , n18 , n31 );
nor ( n646 , n20 , n32 );
nand ( n647 , n643 , n644 , n645 , n646 );
nor ( n648 , n642 , n647 );
nand ( n649 , n641 , n648 );
not ( n650 , n649 );
not ( n651 , n650 );
not ( n652 , n23 );
and ( n653 , n651 , n652 );
not ( n654 , n651 );
and ( n655 , n654 , n23 );
nor ( n656 , n653 , n655 );
not ( n657 , n656 );
and ( n658 , n640 , n657 );
nor ( n659 , n639 , n658 );
and ( n660 , n631 , n659 );
not ( n661 , n631 );
not ( n662 , n659 );
and ( n663 , n661 , n662 );
nor ( n664 , n660 , n663 );
not ( n665 , n664 );
nand ( n666 , n637 , n665 );
not ( n667 , n666 );
or ( n668 , n614 , n667 );
not ( n669 , n664 );
nand ( n670 , n159 , n612 );
not ( n671 , n670 );
not ( n672 , n671 );
not ( n673 , n635 );
or ( n674 , n672 , n673 );
not ( n675 , n160 );
nand ( n676 , n674 , n675 );
nand ( n677 , n669 , n676 );
nand ( n678 , n668 , n677 );
not ( n679 , n678 );
not ( n680 , n669 );
not ( n681 , n635 );
not ( n682 , n615 );
not ( n683 , n613 );
or ( n684 , n682 , n683 );
nand ( n685 , n684 , n670 );
not ( n686 , n685 );
or ( n687 , n681 , n686 );
not ( n688 , n161 );
nand ( n689 , n687 , n688 );
not ( n690 , n689 );
or ( n691 , n680 , n690 );
not ( n692 , n635 );
nand ( n693 , n692 , n664 );
nand ( n694 , n691 , n693 );
not ( n695 , n694 );
nand ( n696 , n679 , n695 );
buf ( n697 , n314 );
not ( n698 , n607 );
xnor ( n699 , n697 , n698 );
not ( n700 , n699 );
not ( n701 , n664 );
nand ( n702 , n701 , n692 , n613 );
nand ( n703 , n158 , n702 );
nor ( n704 , n700 , n703 );
buf ( n705 , n704 );
not ( n706 , n705 );
not ( n707 , n361 );
nor ( n708 , n707 , n606 );
not ( n709 , n371 );
xnor ( n710 , n708 , n709 );
not ( n711 , n342 );
not ( n712 , n709 );
nand ( n713 , n712 , n708 );
not ( n714 , n713 );
nand ( n715 , n711 , n714 );
buf ( n716 , n330 );
not ( n717 , n716 );
and ( n718 , n715 , n717 );
not ( n719 , n715 );
and ( n720 , n719 , n716 );
nor ( n721 , n718 , n720 );
nand ( n722 , n710 , n721 );
not ( n723 , n707 );
not ( n724 , n723 );
not ( n725 , n606 );
not ( n726 , n725 );
and ( n727 , n724 , n726 );
nor ( n728 , n727 , n708 );
nor ( n729 , n728 , n710 );
not ( n730 , n729 );
and ( n731 , n713 , n711 );
not ( n732 , n713 );
not ( n733 , n711 );
and ( n734 , n732 , n733 );
nor ( n735 , n731 , n734 );
nand ( n736 , n735 , n721 );
not ( n737 , n736 );
not ( n738 , n737 );
not ( n739 , n735 );
not ( n740 , n721 );
nand ( n741 , n739 , n740 );
nand ( n742 , n738 , n741 );
and ( n743 , n722 , n730 , n742 );
or ( n744 , n696 , n706 , n743 );
not ( n745 , n744 );
nor ( n746 , n246 , n745 );
not ( n747 , n746 );
not ( n748 , n280 );
not ( n749 , n1 );
and ( n750 , n748 , n749 );
not ( n751 , n286 );
not ( n752 , n271 );
or ( n753 , n751 , n752 );
nand ( n754 , n753 , n26 );
not ( n755 , n24 );
not ( n756 , n23 );
nor ( n757 , n21 , n22 );
nand ( n758 , n755 , n756 , n757 );
nor ( n759 , n758 , n647 );
and ( n760 , n759 , n323 );
and ( n761 , n280 , n760 );
not ( n762 , n1 );
nor ( n763 , n761 , n762 );
and ( n764 , n754 , n763 );
nor ( n765 , n750 , n764 );
not ( n766 , n1 );
nand ( n767 , n24 , n766 );
not ( n768 , n23 );
not ( n769 , n768 );
not ( n770 , n650 );
or ( n771 , n769 , n770 );
nand ( n772 , n771 , n24 );
not ( n773 , n24 );
nor ( n774 , n23 , n649 );
and ( n775 , n773 , n774 );
not ( n776 , n1 );
nor ( n777 , n775 , n776 );
nand ( n778 , n772 , n777 );
and ( n779 , n767 , n778 );
not ( n780 , n373 );
and ( n781 , n313 , n659 );
nand ( n782 , n780 , n781 , n629 , n278 );
and ( n783 , n782 , n291 );
nor ( n784 , n783 , n605 );
nor ( n785 , n779 , n784 );
xnor ( n786 , n765 , n785 );
not ( n787 , n786 );
not ( n788 , n787 );
not ( n789 , n788 );
not ( n790 , n789 );
not ( n791 , n790 );
not ( n792 , n483 );
nand ( n793 , n792 , n598 );
not ( n794 , n793 );
nor ( n795 , n505 , n627 );
nor ( n796 , n467 , n591 );
nand ( n797 , n794 , n795 , n796 , n496 );
nand ( n798 , n384 , n436 , n523 );
not ( n799 , n798 );
nand ( n800 , n799 , n310 , n656 );
nor ( n801 , n797 , n800 );
not ( n802 , n550 );
nand ( n803 , n802 , n327 );
not ( n804 , n803 );
nand ( n805 , n339 , n778 );
nand ( n806 , n560 , n367 );
nand ( n807 , n276 , n765 );
nor ( n808 , n805 , n806 , n807 );
not ( n809 , n424 );
nor ( n810 , n450 , n459 );
nand ( n811 , n810 , n390 , n381 );
nor ( n812 , n410 , n811 );
nand ( n813 , n809 , n812 , n360 );
nor ( n814 , n813 , n536 , n577 );
nand ( n815 , n804 , n808 , n814 );
not ( n816 , n815 );
and ( n817 , n801 , n816 );
not ( n818 , n621 );
not ( n819 , n285 );
nand ( n820 , n818 , n280 , n819 );
not ( n821 , n820 );
and ( n822 , n281 , n821 );
not ( n823 , n1 );
nor ( n824 , n822 , n823 );
nand ( n825 , n25 , n820 );
and ( n826 , n824 , n825 );
not ( n827 , n1 );
and ( n828 , n25 , n827 );
nor ( n829 , n826 , n828 );
not ( n830 , n829 );
nand ( n831 , n289 , n830 );
nor ( n832 , n817 , n831 );
not ( n833 , n287 );
xor ( n834 , n279 , n833 );
and ( n835 , n1 , n834 );
not ( n836 , n1 );
and ( n837 , n836 , n27 );
or ( n838 , n835 , n837 );
and ( n839 , n832 , n838 );
not ( n840 , n832 );
not ( n841 , n838 );
and ( n842 , n840 , n841 );
nor ( n843 , n839 , n842 );
buf ( n844 , n843 );
and ( n845 , n801 , n816 );
nor ( n846 , n845 , n290 );
not ( n847 , n830 );
and ( n848 , n846 , n847 );
not ( n849 , n846 );
and ( n850 , n849 , n830 );
nor ( n851 , n848 , n850 );
not ( n852 , n851 );
nor ( n853 , n844 , n852 );
buf ( n854 , n853 );
not ( n855 , n854 );
not ( n856 , n855 );
not ( n857 , n84 );
not ( n858 , n857 );
and ( n859 , n856 , n858 );
not ( n860 , n851 );
nand ( n861 , n860 , n844 );
buf ( n862 , n861 );
not ( n863 , n862 );
and ( n864 , n83 , n863 );
nor ( n865 , n859 , n864 );
nand ( n866 , n844 , n851 );
not ( n867 , n866 );
not ( n868 , n867 );
not ( n869 , n868 );
and ( n870 , n81 , n869 );
not ( n871 , n844 );
nand ( n872 , n871 , n852 );
not ( n873 , n872 );
not ( n874 , n873 );
not ( n875 , n82 );
nor ( n876 , n874 , n875 );
nor ( n877 , n870 , n876 );
nand ( n878 , n865 , n877 );
not ( n879 , n878 );
not ( n880 , n879 );
not ( n881 , n861 );
and ( n882 , n47 , n881 );
not ( n883 , n844 );
nand ( n884 , n883 , n860 );
not ( n885 , n884 );
not ( n886 , n885 );
not ( n887 , n46 );
nor ( n888 , n886 , n887 );
nor ( n889 , n882 , n888 );
not ( n890 , n866 );
not ( n891 , n890 );
not ( n892 , n891 );
and ( n893 , n892 , n48 );
nor ( n894 , n860 , n844 );
not ( n895 , n894 );
not ( n896 , n45 );
nor ( n897 , n895 , n896 );
nor ( n898 , n893 , n897 );
nand ( n899 , n889 , n898 );
nand ( n900 , n860 , n844 );
not ( n901 , n900 );
and ( n902 , n51 , n901 );
not ( n903 , n885 );
not ( n904 , n50 );
nor ( n905 , n903 , n904 );
nor ( n906 , n902 , n905 );
not ( n907 , n891 );
and ( n908 , n907 , n49 );
not ( n909 , n894 );
not ( n910 , n52 );
nor ( n911 , n909 , n910 );
nor ( n912 , n908 , n911 );
nand ( n913 , n906 , n912 );
nand ( n914 , n899 , n913 );
not ( n915 , n914 );
buf ( n916 , n853 );
not ( n917 , n916 );
not ( n918 , n917 );
nand ( n919 , n918 , n36 );
not ( n920 , n868 );
nand ( n921 , n33 , n920 );
not ( n922 , n862 );
nand ( n923 , n35 , n922 );
buf ( n924 , n872 );
not ( n925 , n924 );
nand ( n926 , n925 , n34 );
nand ( n927 , n919 , n921 , n923 , n926 );
not ( n928 , n44 );
nor ( n929 , n855 , n928 );
not ( n930 , n42 );
not ( n931 , n867 );
nor ( n932 , n930 , n931 );
nor ( n933 , n929 , n932 );
not ( n934 , n43 );
not ( n935 , n934 );
buf ( n936 , n861 );
not ( n937 , n936 );
and ( n938 , n935 , n937 );
not ( n939 , n41 );
nor ( n940 , n924 , n939 );
nor ( n941 , n938 , n940 );
nand ( n942 , n933 , n941 );
nand ( n943 , n927 , n942 );
not ( n944 , n943 );
not ( n945 , n40 );
not ( n946 , n894 );
or ( n947 , n945 , n946 );
nand ( n948 , n890 , n37 );
nand ( n949 , n947 , n948 );
not ( n950 , n39 );
not ( n951 , n900 );
not ( n952 , n951 );
or ( n953 , n950 , n952 );
nand ( n954 , n885 , n38 );
nand ( n955 , n953 , n954 );
nor ( n956 , n949 , n955 );
not ( n957 , n956 );
not ( n958 , n936 );
not ( n959 , n958 );
not ( n960 , n959 );
nand ( n961 , n957 , n960 );
not ( n962 , n961 );
nand ( n963 , n915 , n944 , n962 );
not ( n964 , n963 );
not ( n965 , n916 );
not ( n966 , n68 );
nor ( n967 , n965 , n966 );
not ( n968 , n872 );
not ( n969 , n968 );
not ( n970 , n66 );
nor ( n971 , n969 , n970 );
nor ( n972 , n967 , n971 );
not ( n973 , n65 );
not ( n974 , n867 );
nor ( n975 , n973 , n974 );
not ( n976 , n67 );
nor ( n977 , n976 , n936 );
nor ( n978 , n975 , n977 );
nand ( n979 , n972 , n978 );
buf ( n980 , n979 );
not ( n981 , n980 );
and ( n982 , n61 , n869 );
not ( n983 , n916 );
not ( n984 , n64 );
nor ( n985 , n983 , n984 );
nor ( n986 , n982 , n985 );
and ( n987 , n63 , n958 );
not ( n988 , n873 );
not ( n989 , n62 );
nor ( n990 , n988 , n989 );
nor ( n991 , n987 , n990 );
nand ( n992 , n986 , n991 );
buf ( n993 , n992 );
not ( n994 , n993 );
nor ( n995 , n981 , n994 );
not ( n996 , n55 );
not ( n997 , n996 );
not ( n998 , n881 );
not ( n999 , n998 );
and ( n1000 , n997 , n999 );
not ( n1001 , n855 );
and ( n1002 , n56 , n1001 );
nor ( n1003 , n1000 , n1002 );
not ( n1004 , n54 );
not ( n1005 , n873 );
nor ( n1006 , n1004 , n1005 );
not ( n1007 , n53 );
nor ( n1008 , n1007 , n931 );
nor ( n1009 , n1006 , n1008 );
nand ( n1010 , n1003 , n1009 );
not ( n1011 , n60 );
nor ( n1012 , n1011 , n917 );
not ( n1013 , n57 );
nor ( n1014 , n1013 , n936 );
nor ( n1015 , n1012 , n1014 );
not ( n1016 , n59 );
not ( n1017 , n873 );
nor ( n1018 , n1016 , n1017 );
not ( n1019 , n58 );
nor ( n1020 , n974 , n1019 );
nor ( n1021 , n1018 , n1020 );
nand ( n1022 , n1015 , n1021 );
nand ( n1023 , n1010 , n1022 );
not ( n1024 , n1023 );
nand ( n1025 , n964 , n995 , n1024 );
not ( n1026 , n1025 );
not ( n1027 , n1026 );
not ( n1028 , n998 );
and ( n1029 , n71 , n1028 );
not ( n1030 , n72 );
nor ( n1031 , n1030 , n855 );
nor ( n1032 , n1029 , n1031 );
not ( n1033 , n931 );
and ( n1034 , n1033 , n69 );
not ( n1035 , n70 );
nor ( n1036 , n1005 , n1035 );
nor ( n1037 , n1034 , n1036 );
nand ( n1038 , n1032 , n1037 );
not ( n1039 , n924 );
nand ( n1040 , n1039 , n74 );
nand ( n1041 , n918 , n76 );
not ( n1042 , n868 );
nand ( n1043 , n1042 , n73 );
not ( n1044 , n862 );
nand ( n1045 , n75 , n1044 );
nand ( n1046 , n1040 , n1041 , n1043 , n1045 );
nand ( n1047 , n1038 , n1046 );
nor ( n1048 , n1027 , n1047 );
not ( n1049 , n1048 );
and ( n1050 , n880 , n1049 );
and ( n1051 , n879 , n1048 );
nor ( n1052 , n1050 , n1051 );
not ( n1053 , n1052 );
not ( n1054 , n1053 );
or ( n1055 , n791 , n1054 );
nor ( n1056 , n1023 , n1047 );
nand ( n1057 , n865 , n877 );
not ( n1058 , n80 );
not ( n1059 , n854 );
nor ( n1060 , n1058 , n1059 );
not ( n1061 , n78 );
nor ( n1062 , n1061 , n931 );
nor ( n1063 , n1060 , n1062 );
nand ( n1064 , n79 , n968 );
nand ( n1065 , n77 , n901 );
and ( n1066 , n1064 , n1065 );
nand ( n1067 , n1063 , n1066 );
nand ( n1068 , n1057 , n1067 );
nand ( n1069 , n992 , n913 , n979 , n899 );
nor ( n1070 , n1068 , n1069 );
nor ( n1071 , n961 , n943 );
and ( n1072 , n1056 , n1070 , n1071 );
buf ( n1073 , n1072 );
not ( n1074 , n120 );
buf ( n1075 , n916 );
not ( n1076 , n1075 );
or ( n1077 , n1074 , n1076 );
nand ( n1078 , n122 , n1039 );
nand ( n1079 , n1077 , n1078 );
not ( n1080 , n121 );
not ( n1081 , n868 );
not ( n1082 , n1081 );
or ( n1083 , n1080 , n1082 );
nand ( n1084 , n123 , n1044 );
nand ( n1085 , n1083 , n1084 );
nor ( n1086 , n1079 , n1085 );
not ( n1087 , n1086 );
xnor ( n1088 , n1073 , n1087 );
not ( n1089 , n1088 );
not ( n1090 , n1089 );
not ( n1091 , n1059 );
nand ( n1092 , n114 , n1091 );
not ( n1093 , n936 );
nand ( n1094 , n115 , n1093 );
not ( n1095 , n1017 );
nand ( n1096 , n113 , n1095 );
nand ( n1097 , n112 , n869 );
nand ( n1098 , n1092 , n1094 , n1096 , n1097 );
nand ( n1099 , n108 , n1091 );
nand ( n1100 , n111 , n1093 );
not ( n1101 , n1017 );
nand ( n1102 , n110 , n1101 );
nand ( n1103 , n109 , n1033 );
nand ( n1104 , n1099 , n1100 , n1102 , n1103 );
nand ( n1105 , n1098 , n1104 );
not ( n1106 , n87 );
not ( n1107 , n1106 );
not ( n1108 , n998 );
and ( n1109 , n1107 , n1108 );
not ( n1110 , n1059 );
and ( n1111 , n88 , n1110 );
nor ( n1112 , n1109 , n1111 );
not ( n1113 , n1112 );
not ( n1114 , n86 );
not ( n1115 , n1114 );
not ( n1116 , n931 );
and ( n1117 , n1115 , n1116 );
and ( n1118 , n85 , n1101 );
nor ( n1119 , n1117 , n1118 );
not ( n1120 , n1119 );
or ( n1121 , n1113 , n1120 );
nand ( n1122 , n91 , n1075 );
nand ( n1123 , n90 , n1101 );
not ( n1124 , n931 );
nand ( n1125 , n89 , n1124 );
nand ( n1126 , n92 , n1093 );
nand ( n1127 , n1122 , n1123 , n1125 , n1126 );
nand ( n1128 , n1121 , n1127 );
nor ( n1129 , n1105 , n1128 );
nand ( n1130 , n93 , n1124 );
nand ( n1131 , n94 , n1095 );
nand ( n1132 , n96 , n1001 );
nand ( n1133 , n95 , n863 );
nand ( n1134 , n1130 , n1131 , n1132 , n1133 );
not ( n1135 , n1134 );
not ( n1136 , n103 );
not ( n1137 , n1136 );
not ( n1138 , n998 );
and ( n1139 , n1137 , n1138 );
and ( n1140 , n102 , n1110 );
nor ( n1141 , n1139 , n1140 );
not ( n1142 , n1141 );
not ( n1143 , n100 );
not ( n1144 , n1143 );
not ( n1145 , n931 );
and ( n1146 , n1144 , n1145 );
and ( n1147 , n101 , n1095 );
nor ( n1148 , n1146 , n1147 );
not ( n1149 , n1148 );
or ( n1150 , n1142 , n1149 );
nand ( n1151 , n107 , n1075 );
nand ( n1152 , n1124 , n106 );
nand ( n1153 , n105 , n1039 );
nand ( n1154 , n104 , n863 );
nand ( n1155 , n1151 , n1152 , n1153 , n1154 );
nand ( n1156 , n1150 , n1155 );
nor ( n1157 , n1135 , n1156 );
nand ( n1158 , n138 , n918 );
not ( n1159 , n1158 );
not ( n1160 , n136 );
nor ( n1161 , n1160 , n1005 );
not ( n1162 , n137 );
nor ( n1163 , n1162 , n974 );
nor ( n1164 , n1161 , n1163 );
not ( n1165 , n1164 );
or ( n1166 , n1159 , n1165 );
buf ( n1167 , n854 );
nand ( n1168 , n141 , n1167 );
nand ( n1169 , n139 , n925 );
not ( n1170 , n868 );
nand ( n1171 , n1170 , n140 );
nand ( n1172 , n142 , n881 );
nand ( n1173 , n1168 , n1169 , n1171 , n1172 );
nand ( n1174 , n1166 , n1173 );
nand ( n1175 , n98 , n885 );
nand ( n1176 , n97 , n894 );
nand ( n1177 , n99 , n867 );
and ( n1178 , n1175 , n1176 , n1177 );
not ( n1179 , n1178 );
nand ( n1180 , n925 , n133 );
nand ( n1181 , n135 , n1167 );
nand ( n1182 , n1081 , n132 );
not ( n1183 , n862 );
nand ( n1184 , n134 , n1183 );
nand ( n1185 , n1180 , n1181 , n1182 , n1184 );
nand ( n1186 , n1179 , n1185 );
nand ( n1187 , n131 , n1167 );
nand ( n1188 , n1081 , n130 );
not ( n1189 , n924 );
nand ( n1190 , n1189 , n129 );
nand ( n1191 , n128 , n901 );
nand ( n1192 , n1187 , n1188 , n1190 , n1191 );
nand ( n1193 , n1042 , n124 );
not ( n1194 , n924 );
nand ( n1195 , n125 , n1194 );
nand ( n1196 , n126 , n1167 );
not ( n1197 , n862 );
nand ( n1198 , n127 , n1197 );
nand ( n1199 , n1193 , n1195 , n1196 , n1198 );
nand ( n1200 , n1192 , n1199 );
nor ( n1201 , n1174 , n1186 , n1200 );
not ( n1202 , n119 );
not ( n1203 , n1093 );
or ( n1204 , n1202 , n1203 );
nand ( n1205 , n116 , n1001 );
nand ( n1206 , n1204 , n1205 );
not ( n1207 , n118 );
not ( n1208 , n1033 );
or ( n1209 , n1207 , n1208 );
nand ( n1210 , n117 , n1095 );
nand ( n1211 , n1209 , n1210 );
nor ( n1212 , n1206 , n1211 );
nor ( n1213 , n1086 , n1212 );
and ( n1214 , n1129 , n1157 , n1201 , n1213 );
nand ( n1215 , n1214 , n1072 );
nand ( n1216 , n143 , n1101 );
and ( n1217 , n145 , n1124 );
and ( n1218 , n144 , n1091 );
nor ( n1219 , n1217 , n1218 );
and ( n1220 , n1216 , n1219 );
and ( n1221 , n1215 , n1220 );
not ( n1222 , n1215 );
not ( n1223 , n1220 );
and ( n1224 , n1222 , n1223 );
nor ( n1225 , n1221 , n1224 );
nand ( n1226 , n1075 , n149 );
nand ( n1227 , n1194 , n148 );
not ( n1228 , n862 );
nand ( n1229 , n1228 , n146 );
nand ( n1230 , n147 , n892 );
nand ( n1231 , n1226 , n1227 , n1229 , n1230 );
not ( n1232 , n1231 );
not ( n1233 , n1232 );
nand ( n1234 , n1225 , n1233 );
not ( n1235 , n1234 );
not ( n1236 , n914 );
not ( n1237 , n956 );
nand ( n1238 , n1237 , n960 );
not ( n1239 , n1238 );
nand ( n1240 , n1236 , n1239 );
not ( n1241 , n1240 );
buf ( n1242 , n927 );
nand ( n1243 , n1241 , n1242 );
buf ( n1244 , n942 );
not ( n1245 , n1244 );
not ( n1246 , n1245 );
and ( n1247 , n1243 , n1246 );
not ( n1248 , n1243 );
and ( n1249 , n1248 , n1245 );
nor ( n1250 , n1247 , n1249 );
not ( n1251 , n963 );
not ( n1252 , n980 );
not ( n1253 , n1252 );
and ( n1254 , n1251 , n1253 );
not ( n1255 , n1251 );
and ( n1256 , n1255 , n1252 );
or ( n1257 , n1254 , n1256 );
nor ( n1258 , n1250 , n1257 );
not ( n1259 , n151 );
not ( n1260 , n916 );
or ( n1261 , n1259 , n1260 );
nand ( n1262 , n150 , n951 );
nand ( n1263 , n1261 , n1262 );
not ( n1264 , n152 );
not ( n1265 , n885 );
or ( n1266 , n1264 , n1265 );
nand ( n1267 , n867 , n153 );
nand ( n1268 , n1266 , n1267 );
nor ( n1269 , n1263 , n1268 );
buf ( n1270 , n1269 );
not ( n1271 , n1270 );
nand ( n1272 , n157 , n968 );
nand ( n1273 , n156 , n894 );
nand ( n1274 , n154 , n951 );
nand ( n1275 , n155 , n867 );
nand ( n1276 , n1272 , n1273 , n1274 , n1275 );
not ( n1277 , n1276 );
not ( n1278 , n1277 );
nand ( n1279 , n1271 , n1278 );
not ( n1280 , n1279 );
nand ( n1281 , n898 , n889 );
and ( n1282 , n1239 , n1281 );
not ( n1283 , n1239 );
not ( n1284 , n1281 );
and ( n1285 , n1283 , n1284 );
nor ( n1286 , n1282 , n1285 );
not ( n1287 , n1239 );
not ( n1288 , n1287 );
not ( n1289 , n960 );
nand ( n1290 , n1289 , n956 );
not ( n1291 , n1290 );
nor ( n1292 , n1288 , n1291 );
nand ( n1293 , n1280 , n1286 , n1292 );
not ( n1294 , n1293 );
not ( n1295 , n1240 );
not ( n1296 , n1295 );
not ( n1297 , n1242 );
not ( n1298 , n1297 );
or ( n1299 , n1296 , n1298 );
or ( n1300 , n1297 , n1295 );
nand ( n1301 , n1299 , n1300 );
nand ( n1302 , n906 , n912 );
not ( n1303 , n1302 );
nand ( n1304 , n1281 , n1239 );
not ( n1305 , n1304 );
or ( n1306 , n1303 , n1305 );
or ( n1307 , n1302 , n1304 );
nand ( n1308 , n1306 , n1307 );
nand ( n1309 , n1294 , n1301 , n1308 );
not ( n1310 , n1309 );
nand ( n1311 , n1258 , n1310 );
not ( n1312 , n1311 );
not ( n1313 , n1026 );
not ( n1314 , n1038 );
not ( n1315 , n1314 );
not ( n1316 , n1315 );
not ( n1317 , n1316 );
not ( n1318 , n1317 );
not ( n1319 , n1318 );
and ( n1320 , n1313 , n1319 );
not ( n1321 , n1317 );
not ( n1322 , n1025 );
and ( n1323 , n1321 , n1322 );
nor ( n1324 , n1320 , n1323 );
buf ( n1325 , n1022 );
not ( n1326 , n1325 );
not ( n1327 , n1326 );
and ( n1328 , n1251 , n1327 , n995 );
nand ( n1329 , n1003 , n1009 );
not ( n1330 , n1329 );
xor ( n1331 , n1328 , n1330 );
nor ( n1332 , n1324 , n1331 );
nand ( n1333 , n1235 , n1312 , n1332 );
not ( n1334 , n1333 );
not ( n1335 , n1321 );
nand ( n1336 , n1335 , n1322 );
buf ( n1337 , n1046 );
not ( n1338 , n1337 );
buf ( n1339 , n1338 );
not ( n1340 , n1339 );
and ( n1341 , n1336 , n1340 );
not ( n1342 , n1336 );
and ( n1343 , n1342 , n1339 );
nor ( n1344 , n1341 , n1343 );
nand ( n1345 , n1251 , n995 );
buf ( n1346 , n1326 );
and ( n1347 , n1345 , n1346 );
not ( n1348 , n1345 );
not ( n1349 , n1346 );
and ( n1350 , n1348 , n1349 );
nor ( n1351 , n1347 , n1350 );
nand ( n1352 , n1253 , n1251 );
not ( n1353 , n994 );
not ( n1354 , n1353 );
and ( n1355 , n1352 , n1354 );
not ( n1356 , n1352 );
and ( n1357 , n1356 , n1353 );
nor ( n1358 , n1355 , n1357 );
nand ( n1359 , n1351 , n1358 );
nor ( n1360 , n1344 , n1359 );
nand ( n1361 , n1334 , n1360 );
nor ( n1362 , n1361 , n1052 );
nand ( n1363 , n878 , n1048 );
buf ( n1364 , n1067 );
not ( n1365 , n1364 );
xor ( n1366 , n1363 , n1365 );
nand ( n1367 , n1362 , n1366 );
not ( n1368 , n1367 );
not ( n1369 , n1368 );
or ( n1370 , n1090 , n1369 );
and ( n1371 , n1088 , n1367 );
buf ( n1372 , n786 );
not ( n1373 , n1372 );
not ( n1374 , n1373 );
nor ( n1375 , n1371 , n1374 );
nand ( n1376 , n1370 , n1375 );
nand ( n1377 , n1055 , n1376 );
not ( n1378 , n741 );
and ( n1379 , n1377 , n1378 );
not ( n1380 , n784 );
not ( n1381 , n779 );
not ( n1382 , n1381 );
and ( n1383 , n1380 , n1382 );
and ( n1384 , n1381 , n784 );
nor ( n1385 , n1383 , n1384 );
and ( n1386 , n765 , n1381 );
not ( n1387 , n765 );
and ( n1388 , n1387 , n779 );
nor ( n1389 , n1386 , n1388 );
nand ( n1390 , n1385 , n1389 );
buf ( n1391 , n1390 );
not ( n1392 , n1391 );
not ( n1393 , n1392 );
not ( n1394 , n1393 );
not ( n1395 , n1394 );
and ( n1396 , n1395 , n175 );
not ( n1397 , n1395 );
and ( n1398 , n1397 , n595 );
nor ( n1399 , n1396 , n1398 );
or ( n1400 , n552 , n1395 );
buf ( n1401 , n1391 );
not ( n1402 , n1401 );
not ( n1403 , n1402 );
nand ( n1404 , n176 , n1403 );
nand ( n1405 , n1400 , n1404 );
not ( n1406 , n1405 );
buf ( n1407 , n1406 );
not ( n1408 , n526 );
or ( n1409 , n1408 , n1395 );
not ( n1410 , n162 );
nand ( n1411 , n1410 , n1403 );
nand ( n1412 , n1409 , n1411 );
not ( n1413 , n1412 );
not ( n1414 , n1413 );
not ( n1415 , n538 );
not ( n1416 , n1394 );
or ( n1417 , n1415 , n1416 );
not ( n1418 , n177 );
not ( n1419 , n1392 );
nand ( n1420 , n1418 , n1419 );
nand ( n1421 , n1417 , n1420 );
nand ( n1422 , n1414 , n1421 );
not ( n1423 , n507 );
or ( n1424 , n1403 , n1423 );
nand ( n1425 , n165 , n1419 );
nand ( n1426 , n1424 , n1425 );
buf ( n1427 , n1426 );
not ( n1428 , n1427 );
not ( n1429 , n414 );
not ( n1430 , n1429 );
not ( n1431 , n1401 );
not ( n1432 , n1431 );
or ( n1433 , n1430 , n1432 );
buf ( n1434 , n1391 );
nand ( n1435 , n164 , n1434 );
nand ( n1436 , n1433 , n1435 );
not ( n1437 , n1436 );
nand ( n1438 , n1428 , n1437 );
not ( n1439 , n1438 );
not ( n1440 , n439 );
not ( n1441 , n1402 );
or ( n1442 , n1440 , n1441 );
not ( n1443 , n167 );
nand ( n1444 , n1443 , n1419 );
nand ( n1445 , n1442 , n1444 );
not ( n1446 , n426 );
not ( n1447 , n1394 );
or ( n1448 , n1446 , n1447 );
not ( n1449 , n163 );
nand ( n1450 , n1449 , n1419 );
nand ( n1451 , n1448 , n1450 );
not ( n1452 , n1451 );
buf ( n1453 , n1452 );
not ( n1454 , n1453 );
and ( n1455 , n1445 , n1454 );
or ( n1456 , n484 , n1401 );
nand ( n1457 , n166 , n1434 );
nand ( n1458 , n1456 , n1457 );
not ( n1459 , n1458 );
buf ( n1460 , n1459 );
not ( n1461 , n468 );
or ( n1462 , n1461 , n1401 );
not ( n1463 , n171 );
nand ( n1464 , n1463 , n1393 );
nand ( n1465 , n1462 , n1464 );
not ( n1466 , n1465 );
not ( n1467 , n1466 );
not ( n1468 , n1467 );
not ( n1469 , n170 );
not ( n1470 , n1391 );
or ( n1471 , n1469 , n1470 );
not ( n1472 , n390 );
nand ( n1473 , n1472 , n1392 );
nand ( n1474 , n1471 , n1473 );
not ( n1475 , n1474 );
not ( n1476 , n172 );
not ( n1477 , n1476 );
not ( n1478 , n1391 );
or ( n1479 , n1477 , n1478 );
nand ( n1480 , n1389 , n1385 );
not ( n1481 , n1480 );
nand ( n1482 , n460 , n1481 );
nand ( n1483 , n1479 , n1482 );
not ( n1484 , n1483 );
not ( n1485 , n174 );
not ( n1486 , n1480 );
or ( n1487 , n1485 , n1486 );
nand ( n1488 , n6 , n1481 );
nand ( n1489 , n1487 , n1488 );
not ( n1490 , n1489 );
not ( n1491 , n173 );
not ( n1492 , n1491 );
not ( n1493 , n1480 );
or ( n1494 , n1492 , n1493 );
nand ( n1495 , n451 , n1481 );
nand ( n1496 , n1494 , n1495 );
nand ( n1497 , n1490 , n1496 );
nor ( n1498 , n1484 , n1497 );
and ( n1499 , n1475 , n1498 );
not ( n1500 , n168 );
not ( n1501 , n1391 );
or ( n1502 , n1500 , n1501 );
not ( n1503 , n496 );
not ( n1504 , n1391 );
nand ( n1505 , n1503 , n1504 );
nand ( n1506 , n1502 , n1505 );
not ( n1507 , n1506 );
or ( n1508 , n382 , n1401 );
not ( n1509 , n169 );
nand ( n1510 , n1509 , n1434 );
nand ( n1511 , n1508 , n1510 );
not ( n1512 , n1511 );
not ( n1513 , n1512 );
nand ( n1514 , n1499 , n1507 , n1513 );
nor ( n1515 , n1468 , n1514 );
and ( n1516 , n1460 , n1515 );
nand ( n1517 , n1439 , n1455 , n1516 );
nor ( n1518 , n1422 , n1517 );
nand ( n1519 , n1407 , n1518 );
xnor ( n1520 , n1399 , n1519 );
not ( n1521 , n1520 );
and ( n1522 , n729 , n737 );
not ( n1523 , n1522 );
or ( n1524 , n1521 , n1523 );
not ( n1525 , n722 );
and ( n1526 , n735 , n1525 );
not ( n1527 , n1399 );
nand ( n1528 , n1526 , n1527 );
nand ( n1529 , n1524 , n1528 );
nor ( n1530 , n1379 , n1529 );
and ( n1531 , n1452 , n1329 );
not ( n1532 , n1413 );
not ( n1533 , n1316 );
or ( n1534 , n1532 , n1533 );
nand ( n1535 , n1412 , n1315 );
nand ( n1536 , n1534 , n1535 );
nand ( n1537 , n1531 , n1536 );
not ( n1538 , n1537 );
nand ( n1539 , n1413 , n1315 );
not ( n1540 , n1539 );
not ( n1541 , n1421 );
not ( n1542 , n1541 );
not ( n1543 , n1338 );
or ( n1544 , n1542 , n1543 );
nand ( n1545 , n1421 , n1337 );
nand ( n1546 , n1544 , n1545 );
or ( n1547 , n1540 , n1546 );
nand ( n1548 , n1538 , n1547 );
nand ( n1549 , n1540 , n1546 );
and ( n1550 , n1548 , n1549 );
not ( n1551 , n1550 );
nand ( n1552 , n1541 , n1337 );
not ( n1553 , n1552 );
or ( n1554 , n1406 , n878 );
nand ( n1555 , n1406 , n878 );
nand ( n1556 , n1554 , n1555 );
nor ( n1557 , n1553 , n1556 );
not ( n1558 , n1557 );
and ( n1559 , n1551 , n1558 );
nand ( n1560 , n1458 , n1244 );
not ( n1561 , n1560 );
not ( n1562 , n980 );
nor ( n1563 , n1427 , n1562 );
not ( n1564 , n1563 );
nand ( n1565 , n1427 , n1252 );
nand ( n1566 , n1564 , n1565 );
nand ( n1567 , n1561 , n1566 );
nand ( n1568 , n1426 , n980 );
not ( n1569 , n1568 );
nor ( n1570 , n1436 , n994 );
not ( n1571 , n1570 );
nand ( n1572 , n1436 , n994 );
nand ( n1573 , n1571 , n1572 );
nor ( n1574 , n1569 , n1573 );
nor ( n1575 , n1567 , n1574 );
not ( n1576 , n1573 );
not ( n1577 , n1569 );
nor ( n1578 , n1576 , n1577 );
nor ( n1579 , n1575 , n1578 );
not ( n1580 , n1445 );
nand ( n1581 , n1580 , n1326 );
not ( n1582 , n1581 );
and ( n1583 , n1445 , n1325 );
nor ( n1584 , n1582 , n1583 );
not ( n1585 , n1584 );
nand ( n1586 , n1436 , n993 );
not ( n1587 , n1586 );
nand ( n1588 , n1585 , n1587 );
and ( n1589 , n1579 , n1588 );
nand ( n1590 , n1584 , n1586 );
not ( n1591 , n1325 );
nor ( n1592 , n1591 , n1445 );
not ( n1593 , n1592 );
and ( n1594 , n1453 , n1330 );
and ( n1595 , n1451 , n1329 );
nor ( n1596 , n1594 , n1595 );
nand ( n1597 , n1593 , n1596 );
nand ( n1598 , n1590 , n1597 );
nor ( n1599 , n1589 , n1598 );
not ( n1600 , n1593 );
not ( n1601 , n1596 );
and ( n1602 , n1600 , n1601 );
nor ( n1603 , n1599 , n1602 );
not ( n1604 , n1603 );
or ( n1605 , n1531 , n1536 );
nand ( n1606 , n1605 , n1547 );
nor ( n1607 , n1557 , n1606 );
and ( n1608 , n1604 , n1607 );
nor ( n1609 , n1559 , n1608 );
or ( n1610 , n1566 , n1561 );
not ( n1611 , n1574 );
nand ( n1612 , n1610 , n1611 );
nor ( n1613 , n1612 , n1598 );
not ( n1614 , n1277 );
nand ( n1615 , n1614 , n1484 );
nand ( n1616 , n39 , n901 );
nand ( n1617 , n40 , n916 );
nand ( n1618 , n954 , n1616 , n1617 , n948 );
not ( n1619 , n959 );
and ( n1620 , n1618 , n1619 );
not ( n1621 , n1618 );
and ( n1622 , n1621 , n959 );
nor ( n1623 , n1620 , n1622 );
xor ( n1624 , n1475 , n1623 );
nand ( n1625 , n1615 , n1624 );
and ( n1626 , n1489 , n1231 );
not ( n1627 , n1496 );
not ( n1628 , n1627 );
not ( n1629 , n1270 );
or ( n1630 , n1628 , n1629 );
not ( n1631 , n1496 );
or ( n1632 , n1631 , n1270 );
nand ( n1633 , n1630 , n1632 );
nand ( n1634 , n1626 , n1633 );
nor ( n1635 , n1483 , n1276 );
not ( n1636 , n1635 );
not ( n1637 , n1276 );
not ( n1638 , n1637 );
nand ( n1639 , n1638 , n1483 );
nand ( n1640 , n1636 , n1639 );
not ( n1641 , n1631 );
nor ( n1642 , n1641 , n1270 );
nor ( n1643 , n1640 , n1642 );
or ( n1644 , n1634 , n1643 );
nand ( n1645 , n1642 , n1640 );
nand ( n1646 , n1644 , n1645 );
nand ( n1647 , n1625 , n1646 );
not ( n1648 , n1624 );
not ( n1649 , n1615 );
nand ( n1650 , n1648 , n1649 );
nand ( n1651 , n1647 , n1650 );
not ( n1652 , n1239 );
nand ( n1653 , n1474 , n1623 );
nand ( n1654 , n1652 , n1653 );
nor ( n1655 , n1511 , n1281 );
not ( n1656 , n1655 );
nand ( n1657 , n1511 , n1281 );
nand ( n1658 , n1656 , n1657 );
nor ( n1659 , n1654 , n1658 );
nand ( n1660 , n1512 , n1281 );
not ( n1661 , n1660 );
nor ( n1662 , n1507 , n1302 );
not ( n1663 , n1662 );
nand ( n1664 , n1507 , n1302 );
nand ( n1665 , n1663 , n1664 );
nor ( n1666 , n1661 , n1665 );
nor ( n1667 , n1659 , n1666 );
and ( n1668 , n1651 , n1667 );
nand ( n1669 , n1466 , n1242 );
not ( n1670 , n1669 );
not ( n1671 , n1244 );
nor ( n1672 , n1671 , n1458 );
not ( n1673 , n1672 );
not ( n1674 , n1459 );
nand ( n1675 , n1674 , n1245 );
nand ( n1676 , n1673 , n1675 );
nor ( n1677 , n1670 , n1676 );
nand ( n1678 , n1506 , n1302 );
not ( n1679 , n1678 );
nor ( n1680 , n1467 , n1242 );
not ( n1681 , n1680 );
nand ( n1682 , n1242 , n1465 );
nand ( n1683 , n1681 , n1682 );
nor ( n1684 , n1679 , n1683 );
nor ( n1685 , n1677 , n1684 );
nand ( n1686 , n1668 , n1685 );
nand ( n1687 , n1654 , n1658 );
or ( n1688 , n1687 , n1666 );
nand ( n1689 , n1661 , n1665 );
nand ( n1690 , n1688 , n1689 );
and ( n1691 , n1690 , n1685 );
nand ( n1692 , n1679 , n1683 );
nor ( n1693 , n1677 , n1692 );
nor ( n1694 , n1691 , n1693 );
nand ( n1695 , n1670 , n1676 );
not ( n1696 , n1695 );
not ( n1697 , n1696 );
nand ( n1698 , n1686 , n1694 , n1697 );
nand ( n1699 , n1613 , n1698 );
not ( n1700 , n1699 );
nand ( n1701 , n1700 , n1607 );
nand ( n1702 , n1553 , n1556 );
nand ( n1703 , n1609 , n1701 , n1702 );
nand ( n1704 , n1405 , n878 );
not ( n1705 , n1704 );
and ( n1706 , n1399 , n1364 );
not ( n1707 , n1399 );
not ( n1708 , n1364 );
and ( n1709 , n1707 , n1708 );
nor ( n1710 , n1706 , n1709 );
not ( n1711 , n1710 );
and ( n1712 , n1705 , n1711 );
and ( n1713 , n1704 , n1710 );
nor ( n1714 , n1712 , n1713 );
and ( n1715 , n1703 , n1714 );
not ( n1716 , n1703 );
not ( n1717 , n1714 );
and ( n1718 , n1716 , n1717 );
nor ( n1719 , n1715 , n1718 );
and ( n1720 , n740 , n728 );
not ( n1721 , n740 );
and ( n1722 , n1721 , n710 );
nor ( n1723 , n1720 , n1722 );
not ( n1724 , n1723 );
nor ( n1725 , n1724 , n742 );
buf ( n1726 , n1725 );
buf ( n1727 , n1726 );
buf ( n1728 , n1727 );
buf ( n1729 , n1728 );
nand ( n1730 , n1719 , n1729 );
not ( n1731 , n1535 );
not ( n1732 , n1421 );
not ( n1733 , n1338 );
or ( n1734 , n1732 , n1733 );
nand ( n1735 , n1734 , n1552 );
nor ( n1736 , n1731 , n1735 );
and ( n1737 , n1412 , n1314 );
not ( n1738 , n1737 );
nand ( n1739 , n1738 , n1539 );
nand ( n1740 , n1595 , n1739 );
nor ( n1741 , n1736 , n1740 );
and ( n1742 , n1731 , n1735 );
nor ( n1743 , n1741 , n1742 );
not ( n1744 , n1743 );
not ( n1745 , n1545 );
not ( n1746 , n1406 );
or ( n1747 , n1746 , n878 );
nand ( n1748 , n1747 , n1704 );
nor ( n1749 , n1745 , n1748 );
not ( n1750 , n1749 );
and ( n1751 , n1744 , n1750 );
not ( n1752 , n1563 );
not ( n1753 , n1752 );
not ( n1754 , n1586 );
nor ( n1755 , n1436 , n993 );
nor ( n1756 , n1754 , n1755 );
not ( n1757 , n1756 );
nand ( n1758 , n1753 , n1757 );
nor ( n1759 , n1426 , n980 );
not ( n1760 , n1759 );
nand ( n1761 , n1760 , n1568 );
and ( n1762 , n1672 , n1761 );
nand ( n1763 , n1752 , n1756 );
nand ( n1764 , n1762 , n1763 );
nand ( n1765 , n1758 , n1764 );
not ( n1766 , n1570 );
not ( n1767 , n1325 );
nand ( n1768 , n1445 , n1767 );
not ( n1769 , n1768 );
nor ( n1770 , n1769 , n1592 );
nand ( n1771 , n1766 , n1770 );
and ( n1772 , n1765 , n1771 );
not ( n1773 , n1770 );
and ( n1774 , n1570 , n1773 );
nor ( n1775 , n1772 , n1774 );
not ( n1776 , n1583 );
not ( n1777 , n1453 );
not ( n1778 , n1329 );
and ( n1779 , n1777 , n1778 );
nor ( n1780 , n1779 , n1531 );
nand ( n1781 , n1776 , n1780 );
not ( n1782 , n1781 );
or ( n1783 , n1775 , n1782 );
not ( n1784 , n1780 );
nand ( n1785 , n1583 , n1784 );
nand ( n1786 , n1783 , n1785 );
not ( n1787 , n1749 );
nor ( n1788 , n1595 , n1739 );
nor ( n1789 , n1788 , n1736 );
nand ( n1790 , n1787 , n1789 );
not ( n1791 , n1790 );
and ( n1792 , n1786 , n1791 );
nor ( n1793 , n1751 , n1792 );
not ( n1794 , n1763 );
nor ( n1795 , n1672 , n1761 );
nor ( n1796 , n1794 , n1795 );
nand ( n1797 , n1771 , n1796 , n1781 );
nor ( n1798 , n1797 , n1790 );
not ( n1799 , n1511 );
nor ( n1800 , n1799 , n1281 );
not ( n1801 , n1800 );
nand ( n1802 , n1801 , n1660 );
nand ( n1803 , n1475 , n1290 );
nand ( n1804 , n1652 , n1803 );
nand ( n1805 , n1802 , n1804 );
not ( n1806 , n1657 );
nor ( n1807 , n1506 , n1302 );
not ( n1808 , n1807 );
nand ( n1809 , n1808 , n1678 );
nor ( n1810 , n1806 , n1809 );
or ( n1811 , n1805 , n1810 );
nand ( n1812 , n1806 , n1809 );
nand ( n1813 , n1811 , n1812 );
nor ( n1814 , n1466 , n1242 );
not ( n1815 , n1814 );
nand ( n1816 , n1815 , n1669 );
not ( n1817 , n1664 );
nor ( n1818 , n1816 , n1817 );
not ( n1819 , n1682 );
nor ( n1820 , n1458 , n1244 );
not ( n1821 , n1820 );
nand ( n1822 , n1821 , n1560 );
nor ( n1823 , n1819 , n1822 );
nor ( n1824 , n1818 , n1823 );
and ( n1825 , n1813 , n1824 );
nand ( n1826 , n1817 , n1816 );
nor ( n1827 , n1826 , n1823 );
nor ( n1828 , n1825 , n1827 );
nor ( n1829 , n1802 , n1804 );
nor ( n1830 , n1829 , n1810 );
and ( n1831 , n1830 , n1824 );
not ( n1832 , n1623 );
nand ( n1833 , n1475 , n1832 );
and ( n1834 , n1653 , n1833 );
nand ( n1835 , n1639 , n1834 );
nor ( n1836 , n1231 , n1489 );
not ( n1837 , n1836 );
not ( n1838 , n1496 );
nor ( n1839 , n1263 , n1268 );
not ( n1840 , n1839 );
or ( n1841 , n1838 , n1840 );
or ( n1842 , n1496 , n1839 );
nand ( n1843 , n1841 , n1842 );
nand ( n1844 , n1231 , n1843 );
nand ( n1845 , n1837 , n1844 );
not ( n1846 , n1843 );
nand ( n1847 , n1232 , n1846 );
nand ( n1848 , n1845 , n1847 );
not ( n1849 , n1270 );
not ( n1850 , n1631 );
and ( n1851 , n1849 , n1850 );
not ( n1852 , n1277 );
nor ( n1853 , n1484 , n1852 );
not ( n1854 , n1853 );
nand ( n1855 , n1854 , n1615 );
nor ( n1856 , n1851 , n1855 );
or ( n1857 , n1848 , n1856 );
nand ( n1858 , n1851 , n1855 );
nand ( n1859 , n1857 , n1858 );
nand ( n1860 , n1835 , n1859 );
not ( n1861 , n1834 );
not ( n1862 , n1639 );
nand ( n1863 , n1861 , n1862 );
nand ( n1864 , n1860 , n1863 );
and ( n1865 , n1831 , n1864 );
and ( n1866 , n1819 , n1822 );
nor ( n1867 , n1865 , n1866 );
nand ( n1868 , n1828 , n1867 );
nand ( n1869 , n1798 , n1868 );
nand ( n1870 , n1745 , n1748 );
nand ( n1871 , n1793 , n1869 , n1870 );
xnor ( n1872 , n1555 , n1710 );
xor ( n1873 , n1871 , n1872 );
not ( n1874 , n728 );
not ( n1875 , n740 );
or ( n1876 , n1874 , n1875 );
not ( n1877 , n722 );
nand ( n1878 , n1877 , n736 );
nand ( n1879 , n1876 , n1878 );
nand ( n1880 , n1873 , n1879 );
nand ( n1881 , n1530 , n1730 , n1880 );
nand ( n1882 , n1881 , n745 );
nand ( n1883 , n747 , n1882 );
not ( n1884 , n743 );
nand ( n1885 , n1884 , n678 );
nor ( n1886 , n706 , n1885 );
nand ( n1887 , n695 , n1886 );
not ( n1888 , n79 );
and ( n1889 , n1887 , n1888 );
not ( n1890 , n1887 );
not ( n1891 , n1881 );
and ( n1892 , n1890 , n1891 );
nor ( n1893 , n1889 , n1892 );
not ( n1894 , n745 );
nor ( n1895 , n1373 , n1344 );
not ( n1896 , n1895 );
not ( n1897 , n1368 );
buf ( n1898 , n1362 );
not ( n1899 , n1898 );
not ( n1900 , n1366 );
nand ( n1901 , n1899 , n1900 );
nand ( n1902 , n1897 , n1901 , n789 );
nand ( n1903 , n1896 , n1902 );
nand ( n1904 , n1903 , n1378 );
not ( n1905 , n1603 );
not ( n1906 , n1699 );
or ( n1907 , n1905 , n1906 );
not ( n1908 , n1606 );
nand ( n1909 , n1907 , n1908 );
nand ( n1910 , n1909 , n1550 );
not ( n1911 , n1557 );
nand ( n1912 , n1911 , n1702 );
not ( n1913 , n1912 );
and ( n1914 , n1910 , n1913 );
not ( n1915 , n1910 );
and ( n1916 , n1915 , n1912 );
nor ( n1917 , n1914 , n1916 );
and ( n1918 , n1917 , n1729 );
not ( n1919 , n1518 );
and ( n1920 , n1919 , n1407 );
not ( n1921 , n1919 );
not ( n1922 , n1407 );
and ( n1923 , n1921 , n1922 );
nor ( n1924 , n1920 , n1923 );
or ( n1925 , n1924 , n1523 );
nand ( n1926 , n1526 , n1922 );
nand ( n1927 , n1925 , n1926 );
nor ( n1928 , n1918 , n1927 );
not ( n1929 , n1749 );
nand ( n1930 , n1929 , n1870 );
not ( n1931 , n1930 );
not ( n1932 , n1789 );
not ( n1933 , n1868 );
not ( n1934 , n1797 );
not ( n1935 , n1934 );
or ( n1936 , n1933 , n1935 );
not ( n1937 , n1786 );
nand ( n1938 , n1936 , n1937 );
not ( n1939 , n1938 );
or ( n1940 , n1932 , n1939 );
nand ( n1941 , n1940 , n1743 );
not ( n1942 , n1941 );
or ( n1943 , n1931 , n1942 );
or ( n1944 , n1941 , n1930 );
nand ( n1945 , n1943 , n1944 );
nand ( n1946 , n1879 , n1945 );
nand ( n1947 , n1904 , n1928 , n1946 );
not ( n1948 , n1947 );
or ( n1949 , n1894 , n1948 );
nand ( n1950 , n84 , n744 );
nand ( n1951 , n1949 , n1950 );
not ( n1952 , n1374 );
buf ( n1953 , n1331 );
not ( n1954 , n1953 );
not ( n1955 , n1954 );
or ( n1956 , n1952 , n1955 );
not ( n1957 , n1344 );
not ( n1958 , n1957 );
nor ( n1959 , n1234 , n1311 );
not ( n1960 , n1359 );
nand ( n1961 , n1959 , n1960 );
not ( n1962 , n1961 );
buf ( n1963 , n1332 );
nand ( n1964 , n1962 , n1963 );
not ( n1965 , n1964 );
not ( n1966 , n1965 );
or ( n1967 , n1958 , n1966 );
and ( n1968 , n1344 , n1964 );
nor ( n1969 , n1968 , n1372 );
nand ( n1970 , n1967 , n1969 );
nand ( n1971 , n1956 , n1970 );
nand ( n1972 , n1971 , n1378 );
buf ( n1973 , n1868 );
not ( n1974 , n1973 );
not ( n1975 , n1934 );
or ( n1976 , n1974 , n1975 );
nand ( n1977 , n1976 , n1937 );
not ( n1978 , n1788 );
nand ( n1979 , n1740 , n1978 );
not ( n1980 , n1979 );
and ( n1981 , n1977 , n1980 );
not ( n1982 , n1977 );
and ( n1983 , n1982 , n1979 );
nor ( n1984 , n1981 , n1983 );
nand ( n1985 , n1879 , n1984 );
not ( n1986 , n1414 );
not ( n1987 , n1986 );
not ( n1988 , n1987 );
not ( n1989 , n1517 );
or ( n1990 , n1988 , n1989 );
or ( n1991 , n1987 , n1517 );
nand ( n1992 , n1990 , n1991 );
and ( n1993 , n1522 , n1992 );
not ( n1994 , n1526 );
not ( n1995 , n1987 );
not ( n1996 , n1995 );
nor ( n1997 , n1994 , n1996 );
nor ( n1998 , n1993 , n1997 );
nand ( n1999 , n1972 , n1985 , n1998 );
or ( n2000 , n1724 , n742 );
buf ( n2001 , n2000 );
nand ( n2002 , n1603 , n1699 );
buf ( n2003 , n1537 );
nand ( n2004 , n2003 , n1605 );
not ( n2005 , n2004 );
and ( n2006 , n2002 , n2005 );
not ( n2007 , n2002 );
and ( n2008 , n2007 , n2004 );
nor ( n2009 , n2006 , n2008 );
not ( n2010 , n2009 );
nor ( n2011 , n2001 , n2010 );
nor ( n2012 , n1999 , n2011 );
or ( n2013 , n2012 , n744 );
or ( n2014 , n1030 , n745 );
nand ( n2015 , n2013 , n2014 );
not ( n2016 , n1887 );
not ( n2017 , n2016 );
not ( n2018 , n1947 );
or ( n2019 , n2017 , n2018 );
nand ( n2020 , n82 , n1887 );
nand ( n2021 , n2019 , n2020 );
or ( n2022 , n2012 , n1887 );
or ( n2023 , n1035 , n2016 );
nand ( n2024 , n2022 , n2023 );
not ( n2025 , n76 );
not ( n2026 , n744 );
or ( n2027 , n2025 , n2026 );
not ( n2028 , n2002 );
not ( n2029 , n1605 );
or ( n2030 , n2028 , n2029 );
buf ( n2031 , n2003 );
nand ( n2032 , n2030 , n2031 );
nand ( n2033 , n1549 , n1547 );
not ( n2034 , n2033 );
and ( n2035 , n2032 , n2034 );
not ( n2036 , n2032 );
and ( n2037 , n2036 , n2033 );
nor ( n2038 , n2035 , n2037 );
and ( n2039 , n1729 , n2038 );
not ( n2040 , n1879 );
not ( n2041 , n1868 );
not ( n2042 , n1934 );
or ( n2043 , n2041 , n2042 );
nand ( n2044 , n2043 , n1937 );
not ( n2045 , n2044 );
not ( n2046 , n1978 );
or ( n2047 , n2045 , n2046 );
nand ( n2048 , n2047 , n1740 );
nor ( n2049 , n1742 , n1736 );
and ( n2050 , n2048 , n2049 );
not ( n2051 , n2048 );
not ( n2052 , n2049 );
and ( n2053 , n2051 , n2052 );
nor ( n2054 , n2050 , n2053 );
not ( n2055 , n2054 );
or ( n2056 , n2040 , n2055 );
and ( n2057 , n1052 , n1361 );
nor ( n2058 , n2057 , n1372 );
not ( n2059 , n2058 );
not ( n2060 , n1898 );
not ( n2061 , n2060 );
or ( n2062 , n2059 , n2061 );
not ( n2063 , n786 );
not ( n2064 , n2063 );
buf ( n2065 , n1324 );
not ( n2066 , n2065 );
nand ( n2067 , n2064 , n2066 );
nand ( n2068 , n2062 , n2067 );
and ( n2069 , n1378 , n2068 );
not ( n2070 , n1517 );
not ( n2071 , n1986 );
nand ( n2072 , n2070 , n2071 );
and ( n2073 , n2072 , n1421 );
not ( n2074 , n2072 );
and ( n2075 , n2074 , n1541 );
nor ( n2076 , n2073 , n2075 );
or ( n2077 , n1523 , n2076 );
or ( n2078 , n1994 , n1421 );
nand ( n2079 , n2077 , n2078 );
nor ( n2080 , n2069 , n2079 );
nand ( n2081 , n2056 , n2080 );
nor ( n2082 , n2039 , n2081 );
or ( n2083 , n2082 , n744 );
nand ( n2084 , n2027 , n2083 );
not ( n2085 , n1973 );
not ( n2086 , n1795 );
not ( n2087 , n2086 );
or ( n2088 , n2085 , n2087 );
not ( n2089 , n1762 );
nand ( n2090 , n2088 , n2089 );
nand ( n2091 , n1758 , n1763 );
not ( n2092 , n2091 );
and ( n2093 , n2090 , n2092 );
not ( n2094 , n2090 );
and ( n2095 , n2094 , n2091 );
nor ( n2096 , n2093 , n2095 );
nand ( n2097 , n1879 , n2096 );
not ( n2098 , n788 );
buf ( n2099 , n1257 );
not ( n2100 , n2099 );
not ( n2101 , n2100 );
or ( n2102 , n2098 , n2101 );
not ( n2103 , n1351 );
not ( n2104 , n2103 );
buf ( n2105 , n1358 );
nand ( n2106 , n1959 , n2105 );
not ( n2107 , n2106 );
not ( n2108 , n2107 );
not ( n2109 , n2108 );
or ( n2110 , n2104 , n2109 );
and ( n2111 , n1351 , n2107 );
nor ( n2112 , n2111 , n1372 );
nand ( n2113 , n2110 , n2112 );
nand ( n2114 , n2102 , n2113 );
nand ( n2115 , n1378 , n2114 );
buf ( n2116 , n1428 );
nand ( n2117 , n2116 , n1516 );
and ( n2118 , n2117 , n1436 );
not ( n2119 , n2117 );
and ( n2120 , n2119 , n1437 );
nor ( n2121 , n2118 , n2120 );
and ( n2122 , n1522 , n2121 );
nor ( n2123 , n1994 , n1437 );
nor ( n2124 , n2122 , n2123 );
nand ( n2125 , n2097 , n2115 , n2124 );
and ( n2126 , n1668 , n1685 );
nor ( n2127 , n2126 , n1696 );
nand ( n2128 , n2127 , n1694 );
and ( n2129 , n1610 , n2128 );
not ( n2130 , n1567 );
nor ( n2131 , n2129 , n2130 );
not ( n2132 , n2131 );
not ( n2133 , n1611 );
nor ( n2134 , n1578 , n2133 );
not ( n2135 , n2134 );
or ( n2136 , n2132 , n2135 );
or ( n2137 , n2131 , n2134 );
nand ( n2138 , n2136 , n2137 );
not ( n2139 , n2138 );
nor ( n2140 , n2001 , n2139 );
nor ( n2141 , n2125 , n2140 );
or ( n2142 , n2141 , n744 );
or ( n2143 , n984 , n745 );
nand ( n2144 , n2142 , n2143 );
not ( n2145 , n74 );
not ( n2146 , n1887 );
or ( n2147 , n2145 , n2146 );
or ( n2148 , n2082 , n1887 );
nand ( n2149 , n2147 , n2148 );
or ( n2150 , n2141 , n1887 );
or ( n2151 , n989 , n2016 );
nand ( n2152 , n2150 , n2151 );
not ( n2153 , n745 );
nand ( n2154 , n1372 , n1351 );
not ( n2155 , n2065 );
nor ( n2156 , n1961 , n1953 );
not ( n2157 , n2156 );
not ( n2158 , n2157 );
or ( n2159 , n2155 , n2158 );
not ( n2160 , n2065 );
and ( n2161 , n2160 , n2156 );
nor ( n2162 , n2161 , n1372 );
nand ( n2163 , n2159 , n2162 );
nand ( n2164 , n2154 , n2163 );
and ( n2165 , n1378 , n2164 );
not ( n2166 , n1879 );
not ( n2167 , n1973 );
and ( n2168 , n1796 , n1771 );
not ( n2169 , n2168 );
or ( n2170 , n2167 , n2169 );
buf ( n2171 , n1775 );
nand ( n2172 , n2170 , n2171 );
nand ( n2173 , n1785 , n1781 );
and ( n2174 , n2172 , n2173 );
not ( n2175 , n2172 );
not ( n2176 , n2173 );
and ( n2177 , n2175 , n2176 );
nor ( n2178 , n2174 , n2177 );
nor ( n2179 , n2166 , n2178 );
nor ( n2180 , n2165 , n2179 );
not ( n2181 , n1579 );
not ( n2182 , n1612 );
nand ( n2183 , n2128 , n2182 );
not ( n2184 , n2183 );
or ( n2185 , n2181 , n2184 );
nand ( n2186 , n2185 , n1590 );
nand ( n2187 , n2186 , n1588 );
not ( n2188 , n1597 );
nor ( n2189 , n1602 , n2188 );
and ( n2190 , n2187 , n2189 );
not ( n2191 , n2187 );
not ( n2192 , n2189 );
and ( n2193 , n2191 , n2192 );
nor ( n2194 , n2190 , n2193 );
and ( n2195 , n2194 , n1729 );
not ( n2196 , n1516 );
nor ( n2197 , n2196 , n1438 );
nand ( n2198 , n1445 , n2197 );
buf ( n2199 , n1454 );
not ( n2200 , n2199 );
and ( n2201 , n2198 , n2200 );
not ( n2202 , n2198 );
and ( n2203 , n2202 , n2199 );
nor ( n2204 , n2201 , n2203 );
not ( n2205 , n2204 );
or ( n2206 , n2205 , n1523 );
buf ( n2207 , n2199 );
or ( n2208 , n1994 , n2207 );
nand ( n2209 , n2206 , n2208 );
nor ( n2210 , n2195 , n2209 );
nand ( n2211 , n2180 , n2210 );
not ( n2212 , n2211 );
or ( n2213 , n2153 , n2212 );
nand ( n2214 , n56 , n744 );
nand ( n2215 , n2213 , n2214 );
not ( n2216 , n2016 );
not ( n2217 , n2211 );
or ( n2218 , n2216 , n2217 );
nand ( n2219 , n54 , n1887 );
nand ( n2220 , n2218 , n2219 );
not ( n2221 , n60 );
not ( n2222 , n744 );
or ( n2223 , n2221 , n2222 );
not ( n2224 , n1973 );
not ( n2225 , n1796 );
or ( n2226 , n2224 , n2225 );
not ( n2227 , n1765 );
nand ( n2228 , n2226 , n2227 );
not ( n2229 , n1774 );
nand ( n2230 , n2229 , n1771 );
not ( n2231 , n2230 );
and ( n2232 , n2228 , n2231 );
not ( n2233 , n2228 );
and ( n2234 , n2233 , n2230 );
nor ( n2235 , n2232 , n2234 );
nand ( n2236 , n1879 , n2235 );
not ( n2237 , n2157 );
and ( n2238 , n1961 , n1953 );
nor ( n2239 , n2238 , n1372 );
not ( n2240 , n2239 );
or ( n2241 , n2237 , n2240 );
buf ( n2242 , n2105 );
nand ( n2243 , n2064 , n2242 );
nand ( n2244 , n2241 , n2243 );
nand ( n2245 , n1378 , n2244 );
not ( n2246 , n1580 );
not ( n2247 , n2197 );
or ( n2248 , n2246 , n2247 );
or ( n2249 , n1580 , n2197 );
nand ( n2250 , n2248 , n2249 );
and ( n2251 , n1522 , n2250 );
nor ( n2252 , n1994 , n1445 );
nor ( n2253 , n2251 , n2252 );
nand ( n2254 , n2236 , n2245 , n2253 );
nand ( n2255 , n1579 , n2183 );
nand ( n2256 , n1588 , n1590 );
not ( n2257 , n2256 );
and ( n2258 , n2255 , n2257 );
not ( n2259 , n2255 );
and ( n2260 , n2259 , n2256 );
nor ( n2261 , n2258 , n2260 );
not ( n2262 , n2261 );
nor ( n2263 , n2001 , n2262 );
nor ( n2264 , n2254 , n2263 );
or ( n2265 , n2264 , n744 );
nand ( n2266 , n2223 , n2265 );
not ( n2267 , n59 );
not ( n2268 , n1887 );
or ( n2269 , n2267 , n2268 );
or ( n2270 , n2264 , n1887 );
nand ( n2271 , n2269 , n2270 );
nand ( n2272 , n699 , n678 , n694 );
not ( n2273 , n2272 );
nand ( n2274 , n158 , n729 );
not ( n2275 , n702 );
nor ( n2276 , n2274 , n2275 );
nand ( n2277 , n2273 , n2276 , n1378 );
not ( n2278 , n2277 );
not ( n2279 , n2278 );
not ( n2280 , n2279 );
not ( n2281 , n2280 );
not ( n2282 , n2281 );
nand ( n2283 , n1903 , n2282 );
nor ( n2284 , n1723 , n742 );
buf ( n2285 , n2284 );
nor ( n2286 , n703 , n2272 );
nand ( n2287 , n2285 , n2286 );
not ( n2288 , n2287 );
and ( n2289 , n1945 , n2288 );
not ( n2290 , n1526 );
not ( n2291 , n2286 );
or ( n2292 , n2290 , n2291 );
not ( n2293 , n710 );
nand ( n2294 , n728 , n2293 , n737 );
not ( n2295 , n2294 );
nand ( n2296 , n2295 , n704 );
nand ( n2297 , n2292 , n2296 );
not ( n2298 , n2297 );
not ( n2299 , n2298 );
and ( n2300 , n1922 , n2299 );
not ( n2301 , n158 );
and ( n2302 , n83 , n2301 );
nor ( n2303 , n2300 , n2302 );
not ( n2304 , n2272 );
nor ( n2305 , n2274 , n2275 );
nand ( n2306 , n2304 , n2305 , n737 );
not ( n2307 , n2306 );
not ( n2308 , n2307 );
buf ( n2309 , n2308 );
not ( n2310 , n2309 );
not ( n2311 , n1924 );
nand ( n2312 , n2310 , n2311 );
not ( n2313 , n75 );
nand ( n2314 , n39 , n47 );
not ( n2315 , n2314 );
and ( n2316 , n51 , n2315 );
nand ( n2317 , n35 , n2316 );
not ( n2318 , n2317 );
and ( n2319 , n43 , n2318 );
nand ( n2320 , n67 , n2319 );
not ( n2321 , n2320 );
and ( n2322 , n63 , n2321 );
nand ( n2323 , n57 , n2322 );
nor ( n2324 , n996 , n2323 );
nand ( n2325 , n71 , n2324 );
nor ( n2326 , n2313 , n2325 );
or ( n2327 , n83 , n2326 );
nand ( n2328 , n83 , n2326 );
nand ( n2329 , n1725 , n2286 );
nand ( n2330 , n2329 , n2287 );
nor ( n2331 , n2330 , n2278 );
not ( n2332 , n2306 );
nor ( n2333 , n2332 , n2297 );
nand ( n2334 , n2331 , n158 , n2333 );
not ( n2335 , n2334 );
nand ( n2336 , n2327 , n2328 , n2335 );
nand ( n2337 , n2303 , n2312 , n2336 );
nor ( n2338 , n2289 , n2337 );
buf ( n2339 , n2329 );
not ( n2340 , n2339 );
not ( n2341 , n2340 );
not ( n2342 , n2341 );
nand ( n2343 , n1917 , n2342 );
nand ( n2344 , n2283 , n2338 , n2343 );
not ( n2345 , n2282 );
not ( n2346 , n1377 );
or ( n2347 , n2345 , n2346 );
buf ( n2348 , n1719 );
and ( n2349 , n2348 , n2342 );
nand ( n2350 , n1873 , n2288 );
and ( n2351 , n1520 , n2310 );
not ( n2352 , n2335 );
not ( n2353 , n2328 );
nor ( n2354 , n2353 , n77 );
not ( n2355 , n77 );
nor ( n2356 , n2355 , n2328 );
nor ( n2357 , n2352 , n2354 , n2356 );
nor ( n2358 , n2351 , n2357 );
not ( n2359 , n2298 );
and ( n2360 , n1527 , n2359 );
and ( n2361 , n77 , n2301 );
nor ( n2362 , n2360 , n2361 );
nand ( n2363 , n2350 , n2358 , n2362 );
nor ( n2364 , n2349 , n2363 );
nand ( n2365 , n2347 , n2364 );
not ( n2366 , n38 );
not ( n2367 , n1887 );
or ( n2368 , n2366 , n2367 );
not ( n2369 , n1286 );
not ( n2370 , n1278 );
not ( n2371 , n1270 );
not ( n2372 , n1234 );
nand ( n2373 , n2371 , n2372 );
nor ( n2374 , n2370 , n2373 );
not ( n2375 , n1292 );
not ( n2376 , n2375 );
nand ( n2377 , n2374 , n2376 );
nand ( n2378 , n2369 , n2377 );
not ( n2379 , n2377 );
and ( n2380 , n1286 , n2379 );
nor ( n2381 , n2380 , n2064 );
and ( n2382 , n2378 , n2381 );
not ( n2383 , n1373 );
not ( n2384 , n2370 );
and ( n2385 , n2383 , n2384 );
nor ( n2386 , n2382 , n2385 );
not ( n2387 , n2386 );
and ( n2388 , n1378 , n2387 );
not ( n2389 , n1835 );
not ( n2390 , n2389 );
nand ( n2391 , n2390 , n1863 );
not ( n2392 , n2391 );
not ( n2393 , n2392 );
not ( n2394 , n1859 );
not ( n2395 , n2394 );
or ( n2396 , n2393 , n2395 );
not ( n2397 , n2394 );
nand ( n2398 , n2391 , n2397 );
nand ( n2399 , n2396 , n2398 );
and ( n2400 , n1879 , n2399 );
nand ( n2401 , n1650 , n1625 );
not ( n2402 , n1646 );
and ( n2403 , n2401 , n2402 );
not ( n2404 , n2401 );
not ( n2405 , n2402 );
and ( n2406 , n2404 , n2405 );
nor ( n2407 , n2403 , n2406 );
and ( n2408 , n1727 , n2407 );
nor ( n2409 , n2400 , n2408 );
and ( n2410 , n1498 , n1474 );
not ( n2411 , n1498 );
and ( n2412 , n2411 , n1475 );
nor ( n2413 , n2410 , n2412 );
not ( n2414 , n2413 );
and ( n2415 , n1522 , n2414 );
and ( n2416 , n1526 , n1474 );
nor ( n2417 , n2415 , n2416 );
nand ( n2418 , n2409 , n2417 );
nor ( n2419 , n2388 , n2418 );
or ( n2420 , n2419 , n1887 );
nand ( n2421 , n2368 , n2420 );
not ( n2422 , n40 );
not ( n2423 , n744 );
or ( n2424 , n2422 , n2423 );
or ( n2425 , n2419 , n744 );
nand ( n2426 , n2424 , n2425 );
and ( n2427 , n744 , n966 );
not ( n2428 , n744 );
and ( n2429 , n2196 , n2116 );
not ( n2430 , n2196 );
not ( n2431 , n2116 );
and ( n2432 , n2430 , n2431 );
nor ( n2433 , n2429 , n2432 );
not ( n2434 , n2433 );
and ( n2435 , n1522 , n2434 );
nor ( n2436 , n1994 , n2116 );
nor ( n2437 , n2435 , n2436 );
not ( n2438 , n1973 );
not ( n2439 , n2438 );
not ( n2440 , n2439 );
nand ( n2441 , n2089 , n2086 );
not ( n2442 , n2441 );
or ( n2443 , n2440 , n2442 );
not ( n2444 , n2441 );
nand ( n2445 , n2438 , n2444 );
nand ( n2446 , n2443 , n2445 );
nand ( n2447 , n1879 , n2446 );
nand ( n2448 , n1567 , n1610 );
not ( n2449 , n2448 );
buf ( n2450 , n2128 );
not ( n2451 , n2450 );
or ( n2452 , n2449 , n2451 );
or ( n2453 , n2448 , n2450 );
nand ( n2454 , n2452 , n2453 );
nand ( n2455 , n1727 , n2454 );
nand ( n2456 , n2437 , n2447 , n2455 );
not ( n2457 , n2063 );
and ( n2458 , n2457 , n1250 );
not ( n2459 , n2457 );
buf ( n2460 , n1959 );
nor ( n2461 , n2460 , n2242 );
not ( n2462 , n2461 );
nand ( n2463 , n2462 , n2106 );
and ( n2464 , n2459 , n2463 );
or ( n2465 , n2458 , n2464 );
nor ( n2466 , n741 , n2465 );
nor ( n2467 , n2456 , n2466 );
and ( n2468 , n2428 , n2467 );
nor ( n2469 , n2427 , n2468 );
not ( n2470 , n1830 );
not ( n2471 , n1864 );
or ( n2472 , n2470 , n2471 );
not ( n2473 , n1813 );
nand ( n2474 , n2472 , n2473 );
not ( n2475 , n1818 );
and ( n2476 , n2474 , n2475 );
not ( n2477 , n1826 );
nor ( n2478 , n2476 , n2477 );
not ( n2479 , n2478 );
nor ( n2480 , n1866 , n1823 );
not ( n2481 , n2480 );
or ( n2482 , n2479 , n2481 );
or ( n2483 , n2478 , n2480 );
nand ( n2484 , n2482 , n2483 );
not ( n2485 , n2484 );
nor ( n2486 , n2166 , n2485 );
not ( n2487 , n1378 );
not ( n2488 , n2064 );
buf ( n2489 , n1301 );
not ( n2490 , n2489 );
or ( n2491 , n2488 , n2490 );
not ( n2492 , n2099 );
buf ( n2493 , n2372 );
nand ( n2494 , n1310 , n2493 );
nor ( n2495 , n2494 , n1250 );
not ( n2496 , n2495 );
not ( n2497 , n2496 );
or ( n2498 , n2492 , n2497 );
not ( n2499 , n2099 );
and ( n2500 , n2499 , n2495 );
nor ( n2501 , n2500 , n786 );
nand ( n2502 , n2498 , n2501 );
nand ( n2503 , n2491 , n2502 );
not ( n2504 , n2503 );
or ( n2505 , n2487 , n2504 );
not ( n2506 , n1690 );
not ( n2507 , n2506 );
not ( n2508 , n1668 );
not ( n2509 , n2508 );
or ( n2510 , n2507 , n2509 );
not ( n2511 , n1684 );
nand ( n2512 , n2510 , n2511 );
nand ( n2513 , n2512 , n1692 );
not ( n2514 , n1677 );
and ( n2515 , n1697 , n2514 );
and ( n2516 , n2513 , n2515 );
not ( n2517 , n2513 );
not ( n2518 , n2515 );
and ( n2519 , n2517 , n2518 );
nor ( n2520 , n2516 , n2519 );
and ( n2521 , n1728 , n2520 );
xor ( n2522 , n1460 , n1515 );
not ( n2523 , n2522 );
or ( n2524 , n2523 , n1523 );
or ( n2525 , n1994 , n1460 );
nand ( n2526 , n2524 , n2525 );
nor ( n2527 , n2521 , n2526 );
nand ( n2528 , n2505 , n2527 );
nor ( n2529 , n2486 , n2528 );
and ( n2530 , n745 , n2529 );
not ( n2531 , n745 );
and ( n2532 , n2531 , n928 );
nor ( n2533 , n2530 , n2532 );
nand ( n2534 , n2068 , n2282 );
nand ( n2535 , n2038 , n2342 );
and ( n2536 , n2054 , n2288 );
and ( n2537 , n1541 , n2299 );
and ( n2538 , n75 , n2301 );
nor ( n2539 , n2537 , n2538 );
not ( n2540 , n2308 );
not ( n2541 , n2076 );
nand ( n2542 , n2540 , n2541 );
not ( n2543 , n75 );
nand ( n2544 , n2543 , n2325 );
not ( n2545 , n2326 );
nand ( n2546 , n2544 , n2545 , n2335 );
nand ( n2547 , n2539 , n2542 , n2546 );
nor ( n2548 , n2536 , n2547 );
nand ( n2549 , n2534 , n2535 , n2548 );
and ( n2550 , n2016 , n2529 );
not ( n2551 , n2016 );
and ( n2552 , n2551 , n939 );
nor ( n2553 , n2550 , n2552 );
and ( n2554 , n1887 , n970 );
not ( n2555 , n1887 );
and ( n2556 , n2555 , n2467 );
nor ( n2557 , n2554 , n2556 );
nand ( n2558 , n2282 , n1971 );
nand ( n2559 , n2342 , n2009 );
buf ( n2560 , n1984 );
and ( n2561 , n2288 , n2560 );
not ( n2562 , n2298 );
and ( n2563 , n1995 , n2562 );
and ( n2564 , n71 , n2301 );
nor ( n2565 , n2563 , n2564 );
nand ( n2566 , n2540 , n1992 );
or ( n2567 , n71 , n2324 );
nand ( n2568 , n2567 , n2325 );
not ( n2569 , n2568 );
nand ( n2570 , n2569 , n2335 );
nand ( n2571 , n2565 , n2566 , n2570 );
nor ( n2572 , n2561 , n2571 );
nand ( n2573 , n2558 , n2559 , n2572 );
nand ( n2574 , n704 , n694 );
not ( n2575 , n2574 );
nand ( n2576 , n2575 , n679 );
not ( n2577 , n2576 );
nor ( n2578 , n730 , n741 );
nand ( n2579 , n2577 , n2578 );
not ( n2580 , n2579 );
nand ( n2581 , n2580 , n1971 );
not ( n2582 , n2576 );
nand ( n2583 , n2582 , n1726 );
not ( n2584 , n2583 );
not ( n2585 , n2584 );
not ( n2586 , n2585 );
nand ( n2587 , n2586 , n2009 );
not ( n2588 , n2576 );
buf ( n2589 , n2285 );
nand ( n2590 , n2588 , n2589 );
not ( n2591 , n2590 );
and ( n2592 , n2591 , n2560 );
not ( n2593 , n2576 );
nand ( n2594 , n2593 , n1526 );
not ( n2595 , n2594 );
and ( n2596 , n1995 , n2595 );
nor ( n2597 , n2568 , n2296 );
nor ( n2598 , n2596 , n2597 );
not ( n2599 , n2576 );
nand ( n2600 , n2599 , n1522 );
not ( n2601 , n2600 );
nand ( n2602 , n2601 , n1992 );
nor ( n2603 , n729 , n741 );
not ( n2604 , n2603 );
nand ( n2605 , n2294 , n695 );
nand ( n2606 , n2604 , n705 , n1885 , n2605 );
nand ( n2607 , n69 , n2606 );
nand ( n2608 , n2598 , n2602 , n2607 );
nor ( n2609 , n2592 , n2608 );
nand ( n2610 , n2581 , n2587 , n2609 );
nand ( n2611 , n2580 , n2164 );
not ( n2612 , n2178 );
and ( n2613 , n2591 , n2612 );
and ( n2614 , n53 , n2606 );
and ( n2615 , n996 , n2323 );
nor ( n2616 , n2615 , n2324 );
not ( n2617 , n2296 );
and ( n2618 , n2616 , n2617 );
nor ( n2619 , n2614 , n2618 );
nand ( n2620 , n2601 , n2204 );
not ( n2621 , n2207 );
nand ( n2622 , n2621 , n2595 );
nand ( n2623 , n2619 , n2620 , n2622 );
nor ( n2624 , n2613 , n2623 );
buf ( n2625 , n2194 );
nand ( n2626 , n2625 , n2586 );
nand ( n2627 , n2611 , n2624 , n2626 );
nand ( n2628 , n2282 , n2164 );
and ( n2629 , n2288 , n2612 );
and ( n2630 , n2621 , n2359 );
and ( n2631 , n55 , n2301 );
nor ( n2632 , n2630 , n2631 );
nand ( n2633 , n2310 , n2204 );
not ( n2634 , n2616 );
not ( n2635 , n2634 );
nand ( n2636 , n2635 , n2335 );
nand ( n2637 , n2632 , n2633 , n2636 );
nor ( n2638 , n2629 , n2637 );
nand ( n2639 , n2625 , n2342 );
nand ( n2640 , n2628 , n2638 , n2639 );
not ( n2641 , n2281 );
nand ( n2642 , n2641 , n2244 );
and ( n2643 , n2235 , n2288 );
not ( n2644 , n2308 );
and ( n2645 , n2250 , n2644 );
not ( n2646 , n57 );
nor ( n2647 , n2646 , n158 );
nor ( n2648 , n2645 , n2647 );
nand ( n2649 , n1580 , n2299 );
or ( n2650 , n57 , n2322 );
nand ( n2651 , n2650 , n2323 );
not ( n2652 , n2651 );
nand ( n2653 , n2652 , n2335 );
nand ( n2654 , n2648 , n2649 , n2653 );
nor ( n2655 , n2643 , n2654 );
nand ( n2656 , n2261 , n2342 );
nand ( n2657 , n2642 , n2655 , n2656 );
not ( n2658 , n788 );
not ( n2659 , n2371 );
or ( n2660 , n2658 , n2659 );
not ( n2661 , n2374 );
not ( n2662 , n2661 );
not ( n2663 , n2375 );
not ( n2664 , n2663 );
not ( n2665 , n2664 );
or ( n2666 , n2662 , n2665 );
and ( n2667 , n2374 , n2663 );
nor ( n2668 , n2667 , n1372 );
nand ( n2669 , n2666 , n2668 );
nand ( n2670 , n2660 , n2669 );
and ( n2671 , n1378 , n2670 );
not ( n2672 , n1879 );
and ( n2673 , n1836 , n1847 );
not ( n2674 , n1844 );
nor ( n2675 , n2673 , n2674 );
not ( n2676 , n2675 );
not ( n2677 , n1858 );
nor ( n2678 , n2677 , n1856 );
not ( n2679 , n2678 );
or ( n2680 , n2676 , n2679 );
or ( n2681 , n2675 , n2678 );
nand ( n2682 , n2680 , n2681 );
not ( n2683 , n2682 );
or ( n2684 , n2672 , n2683 );
not ( n2685 , n1643 );
nand ( n2686 , n2685 , n1645 );
not ( n2687 , n2686 );
not ( n2688 , n1634 );
not ( n2689 , n2688 );
or ( n2690 , n2687 , n2689 );
or ( n2691 , n2686 , n2688 );
nand ( n2692 , n2690 , n2691 );
and ( n2693 , n1726 , n2692 );
and ( n2694 , n1497 , n1484 );
not ( n2695 , n1497 );
and ( n2696 , n2695 , n1483 );
nor ( n2697 , n2694 , n2696 );
and ( n2698 , n1522 , n2697 );
and ( n2699 , n1526 , n1484 );
nor ( n2700 , n2693 , n2698 , n2699 );
nand ( n2701 , n2684 , n2700 );
nor ( n2702 , n2671 , n2701 );
or ( n2703 , n2702 , n1887 );
not ( n2704 , n157 );
or ( n2705 , n2704 , n2016 );
nand ( n2706 , n2703 , n2705 );
nand ( n2707 , n2580 , n2244 );
and ( n2708 , n2235 , n2591 );
and ( n2709 , n2250 , n2601 );
nor ( n2710 , n1445 , n2594 );
nor ( n2711 , n2709 , n2710 );
and ( n2712 , n58 , n2606 );
not ( n2713 , n2651 );
and ( n2714 , n2713 , n2617 );
nor ( n2715 , n2712 , n2714 );
nand ( n2716 , n2711 , n2715 );
nor ( n2717 , n2708 , n2716 );
nand ( n2718 , n2261 , n2586 );
nand ( n2719 , n2707 , n2717 , n2718 );
nand ( n2720 , n2114 , n2580 );
nand ( n2721 , n2586 , n2138 );
nand ( n2722 , n2591 , n2096 );
and ( n2723 , n2121 , n2601 );
or ( n2724 , n1437 , n2594 );
xor ( n2725 , n63 , n2321 );
not ( n2726 , n2725 );
or ( n2727 , n2726 , n2296 );
nand ( n2728 , n2724 , n2727 );
not ( n2729 , n61 );
not ( n2730 , n2606 );
nor ( n2731 , n2729 , n2730 );
nor ( n2732 , n2723 , n2728 , n2731 );
nand ( n2733 , n2720 , n2721 , n2722 , n2732 );
not ( n2734 , n787 );
not ( n2735 , n2734 );
not ( n2736 , n1286 );
or ( n2737 , n2735 , n2736 );
not ( n2738 , n2489 );
buf ( n2739 , n1308 );
buf ( n2740 , n1293 );
not ( n2741 , n2493 );
nor ( n2742 , n2740 , n2741 );
nand ( n2743 , n2739 , n2742 );
not ( n2744 , n2743 );
not ( n2745 , n2744 );
or ( n2746 , n2738 , n2745 );
not ( n2747 , n2489 );
and ( n2748 , n2747 , n2743 );
nor ( n2749 , n2748 , n2457 );
nand ( n2750 , n2746 , n2749 );
nand ( n2751 , n2737 , n2750 );
and ( n2752 , n1378 , n2751 );
not ( n2753 , n1879 );
not ( n2754 , n1829 );
not ( n2755 , n2754 );
not ( n2756 , n1864 );
or ( n2757 , n2755 , n2756 );
nand ( n2758 , n2757 , n1805 );
not ( n2759 , n1810 );
nand ( n2760 , n2759 , n1812 );
and ( n2761 , n2758 , n2760 );
not ( n2762 , n2758 );
not ( n2763 , n2760 );
and ( n2764 , n2762 , n2763 );
nor ( n2765 , n2761 , n2764 );
not ( n2766 , n2765 );
not ( n2767 , n2766 );
or ( n2768 , n2753 , n2767 );
buf ( n2769 , n1651 );
not ( n2770 , n2769 );
not ( n2771 , n1659 );
not ( n2772 , n2771 );
or ( n2773 , n2770 , n2772 );
nand ( n2774 , n2773 , n1687 );
not ( n2775 , n1666 );
nand ( n2776 , n2775 , n1689 );
and ( n2777 , n2774 , n2776 );
not ( n2778 , n2774 );
not ( n2779 , n2776 );
and ( n2780 , n2778 , n2779 );
nor ( n2781 , n2777 , n2780 );
not ( n2782 , n2781 );
and ( n2783 , n1728 , n2782 );
and ( n2784 , n1513 , n1499 );
and ( n2785 , n2784 , n1506 );
not ( n2786 , n2784 );
and ( n2787 , n2786 , n1507 );
nor ( n2788 , n2785 , n2787 );
or ( n2789 , n1523 , n2788 );
or ( n2790 , n1994 , n1507 );
nand ( n2791 , n2789 , n2790 );
nor ( n2792 , n2783 , n2791 );
nand ( n2793 , n2768 , n2792 );
nor ( n2794 , n2752 , n2793 );
or ( n2795 , n2794 , n1887 );
or ( n2796 , n904 , n2016 );
nand ( n2797 , n2795 , n2796 );
or ( n2798 , n2794 , n744 );
or ( n2799 , n910 , n745 );
nand ( n2800 , n2798 , n2799 );
or ( n2801 , n2702 , n744 );
not ( n2802 , n156 );
or ( n2803 , n2802 , n745 );
nand ( n2804 , n2801 , n2803 );
or ( n2805 , n2281 , n2386 );
not ( n2806 , n39 );
and ( n2807 , n2806 , n2335 );
and ( n2808 , n1474 , n2359 );
nor ( n2809 , n2807 , n2808 );
and ( n2810 , n2288 , n2399 );
and ( n2811 , n2407 , n2340 );
or ( n2812 , n2308 , n2413 );
or ( n2813 , n2806 , n158 );
nand ( n2814 , n2812 , n2813 );
nor ( n2815 , n2810 , n2811 , n2814 );
nand ( n2816 , n2805 , n2809 , n2815 );
buf ( n2817 , n2280 );
nand ( n2818 , n2114 , n2817 );
nand ( n2819 , n2342 , n2138 );
nand ( n2820 , n2288 , n2096 );
not ( n2821 , n2725 );
not ( n2822 , n2335 );
or ( n2823 , n2821 , n2822 );
nand ( n2824 , n1436 , n2299 );
nand ( n2825 , n2823 , n2824 );
not ( n2826 , n2121 );
or ( n2827 , n2826 , n2309 );
nand ( n2828 , n63 , n2301 );
nand ( n2829 , n2827 , n2828 );
nor ( n2830 , n2825 , n2829 );
nand ( n2831 , n2818 , n2819 , n2820 , n2830 );
not ( n2832 , n2503 );
or ( n2833 , n2579 , n2832 );
not ( n2834 , n2520 );
or ( n2835 , n2834 , n2585 );
and ( n2836 , n2484 , n2591 );
and ( n2837 , n42 , n2606 );
xor ( n2838 , n43 , n2318 );
and ( n2839 , n2838 , n2617 );
nor ( n2840 , n2837 , n2839 );
not ( n2841 , n1460 );
nand ( n2842 , n2841 , n2595 );
nand ( n2843 , n2522 , n2601 );
nand ( n2844 , n2840 , n2842 , n2843 );
nor ( n2845 , n2836 , n2844 );
nand ( n2846 , n2833 , n2835 , n2845 );
not ( n2847 , n2494 );
not ( n2848 , n2847 );
not ( n2849 , n1250 );
not ( n2850 , n2849 );
or ( n2851 , n2848 , n2850 );
and ( n2852 , n2494 , n1250 );
nor ( n2853 , n2852 , n786 );
nand ( n2854 , n2851 , n2853 );
nand ( n2855 , n786 , n2739 );
and ( n2856 , n2854 , n2855 );
nor ( n2857 , n741 , n2856 );
and ( n2858 , n1514 , n1468 );
not ( n2859 , n1514 );
not ( n2860 , n1468 );
and ( n2861 , n2859 , n2860 );
nor ( n2862 , n2858 , n2861 );
and ( n2863 , n1522 , n2862 );
not ( n2864 , n2860 );
and ( n2865 , n1526 , n2864 );
nor ( n2866 , n2863 , n2865 );
not ( n2867 , n1813 );
nand ( n2868 , n1863 , n2394 );
nand ( n2869 , n1835 , n1830 , n2868 );
nand ( n2870 , n2867 , n2869 );
nand ( n2871 , n1826 , n2475 );
not ( n2872 , n2871 );
and ( n2873 , n2870 , n2872 );
not ( n2874 , n2870 );
and ( n2875 , n2874 , n2871 );
nor ( n2876 , n2873 , n2875 );
nand ( n2877 , n1879 , n2876 );
nand ( n2878 , n1650 , n2402 );
nand ( n2879 , n1625 , n2878 , n1667 );
nand ( n2880 , n2506 , n2879 );
not ( n2881 , n2880 );
not ( n2882 , n2881 );
nand ( n2883 , n1692 , n2511 );
not ( n2884 , n2883 );
not ( n2885 , n2884 );
or ( n2886 , n2882 , n2885 );
nand ( n2887 , n2880 , n2883 );
nand ( n2888 , n2886 , n2887 );
nand ( n2889 , n1727 , n2888 );
nand ( n2890 , n2866 , n2877 , n2889 );
nor ( n2891 , n2857 , n2890 );
or ( n2892 , n2891 , n744 );
not ( n2893 , n36 );
or ( n2894 , n2893 , n745 );
nand ( n2895 , n2892 , n2894 );
or ( n2896 , n2891 , n1887 );
not ( n2897 , n34 );
or ( n2898 , n2897 , n2016 );
nand ( n2899 , n2896 , n2898 );
and ( n2900 , n2591 , n2766 );
nor ( n2901 , n2585 , n2781 );
nor ( n2902 , n2900 , n2901 );
nand ( n2903 , n2751 , n2580 );
and ( n2904 , n49 , n2606 );
and ( n2905 , n1506 , n2595 );
nor ( n2906 , n2904 , n2905 );
not ( n2907 , n2788 );
and ( n2908 , n2601 , n2907 );
xor ( n2909 , n51 , n2315 );
and ( n2910 , n2909 , n2617 );
nor ( n2911 , n2908 , n2910 );
nand ( n2912 , n2902 , n2903 , n2906 , n2911 );
nand ( n2913 , n2817 , n2503 );
and ( n2914 , n2838 , n2335 );
and ( n2915 , n2522 , n2540 );
nor ( n2916 , n2914 , n2915 );
and ( n2917 , n2841 , n2359 );
and ( n2918 , n43 , n2301 );
nor ( n2919 , n2917 , n2918 );
and ( n2920 , n2484 , n2288 );
and ( n2921 , n2520 , n2340 );
nor ( n2922 , n2920 , n2921 );
nand ( n2923 , n2913 , n2916 , n2919 , n2922 );
or ( n2924 , n2579 , n2386 );
not ( n2925 , n37 );
not ( n2926 , n2606 );
or ( n2927 , n2925 , n2926 );
or ( n2928 , n2600 , n2413 );
nand ( n2929 , n2927 , n2928 );
not ( n2930 , n2591 );
not ( n2931 , n2399 );
or ( n2932 , n2930 , n2931 );
nand ( n2933 , n2407 , n2584 );
nand ( n2934 , n2932 , n2933 );
or ( n2935 , n1475 , n2594 );
or ( n2936 , n39 , n2296 );
nand ( n2937 , n2935 , n2936 );
nor ( n2938 , n2929 , n2934 , n2937 );
nand ( n2939 , n2924 , n2938 );
not ( n2940 , n46 );
not ( n2941 , n1887 );
or ( n2942 , n2940 , n2941 );
or ( n2943 , n1373 , n2664 );
nor ( n2944 , n2739 , n2742 );
not ( n2945 , n2944 );
nand ( n2946 , n2945 , n787 , n2743 );
nand ( n2947 , n2943 , n2946 );
and ( n2948 , n1378 , n2947 );
and ( n2949 , n2771 , n1687 );
xor ( n2950 , n2949 , n2769 );
and ( n2951 , n2950 , n1727 );
not ( n2952 , n1513 );
not ( n2953 , n1499 );
nand ( n2954 , n2952 , n2953 );
not ( n2955 , n2954 );
nor ( n2956 , n2955 , n2784 );
not ( n2957 , n2956 );
or ( n2958 , n1523 , n2957 );
not ( n2959 , n2952 );
or ( n2960 , n1994 , n2959 );
nand ( n2961 , n2958 , n2960 );
nor ( n2962 , n2951 , n2961 );
nand ( n2963 , n1805 , n2754 );
not ( n2964 , n2963 );
and ( n2965 , n1864 , n2964 );
not ( n2966 , n1864 );
and ( n2967 , n2966 , n2963 );
nor ( n2968 , n2965 , n2967 );
nand ( n2969 , n2968 , n1879 );
nand ( n2970 , n2962 , n2969 );
nor ( n2971 , n2948 , n2970 );
or ( n2972 , n1887 , n2971 );
nand ( n2973 , n2942 , n2972 );
not ( n2974 , n2856 );
nand ( n2975 , n2280 , n2974 );
nand ( n2976 , n2876 , n2288 );
and ( n2977 , n2888 , n2340 );
not ( n2978 , n35 );
not ( n2979 , n2301 );
or ( n2980 , n2978 , n2979 );
not ( n2981 , n2307 );
not ( n2982 , n2862 );
or ( n2983 , n2981 , n2982 );
nand ( n2984 , n2980 , n2983 );
not ( n2985 , n2864 );
nor ( n2986 , n2985 , n2298 );
nor ( n2987 , n2977 , n2984 , n2986 );
or ( n2988 , n35 , n2316 );
nand ( n2989 , n2988 , n2317 );
not ( n2990 , n2989 );
nand ( n2991 , n2990 , n2335 );
nand ( n2992 , n2975 , n2976 , n2987 , n2991 );
not ( n2993 , n45 );
not ( n2994 , n744 );
or ( n2995 , n2993 , n2994 );
or ( n2996 , n744 , n2971 );
nand ( n2997 , n2995 , n2996 );
not ( n2998 , n2751 );
or ( n2999 , n2998 , n2281 );
not ( n3000 , n2909 );
not ( n3001 , n2335 );
or ( n3002 , n3000 , n3001 );
nor ( n3003 , n2339 , n2781 );
nor ( n3004 , n1507 , n2298 );
not ( n3005 , n51 );
nor ( n3006 , n3005 , n158 );
nor ( n3007 , n2981 , n2788 );
nor ( n3008 , n3003 , n3004 , n3006 , n3007 );
nand ( n3009 , n3002 , n3008 );
nor ( n3010 , n2287 , n2765 );
nor ( n3011 , n3009 , n3010 );
nand ( n3012 , n2999 , n3011 );
nand ( n3013 , n2817 , n2670 );
and ( n3014 , n2697 , n2540 );
and ( n3015 , n2288 , n2682 );
nor ( n3016 , n3014 , n3015 );
nor ( n3017 , n2301 , n2335 );
not ( n3018 , n3017 );
and ( n3019 , n154 , n3018 );
not ( n3020 , n2340 );
not ( n3021 , n2692 );
or ( n3022 , n3020 , n3021 );
or ( n3023 , n1483 , n2298 );
nand ( n3024 , n3022 , n3023 );
nor ( n3025 , n3019 , n3024 );
nand ( n3026 , n3013 , n3016 , n3025 );
not ( n3027 , n2465 );
nand ( n3028 , n3027 , n2817 );
or ( n3029 , n67 , n2319 );
nand ( n3030 , n3029 , n2320 );
not ( n3031 , n3030 );
not ( n3032 , n2334 );
and ( n3033 , n3031 , n3032 );
and ( n3034 , n2288 , n2446 );
nor ( n3035 , n3033 , n3034 );
not ( n3036 , n2341 );
and ( n3037 , n3036 , n2454 );
not ( n3038 , n2116 );
not ( n3039 , n3038 );
not ( n3040 , n2299 );
or ( n3041 , n3039 , n3040 );
not ( n3042 , n2308 );
and ( n3043 , n2434 , n3042 );
not ( n3044 , n67 );
nor ( n3045 , n3044 , n158 );
nor ( n3046 , n3043 , n3045 );
nand ( n3047 , n3041 , n3046 );
nor ( n3048 , n3037 , n3047 );
nand ( n3049 , n3028 , n3035 , n3048 );
not ( n3050 , n2661 );
and ( n3051 , n2370 , n2373 );
nor ( n3052 , n3051 , n786 );
not ( n3053 , n3052 );
or ( n3054 , n3050 , n3053 );
nand ( n3055 , n786 , n1233 );
nand ( n3056 , n3054 , n3055 );
and ( n3057 , n1378 , n3056 );
not ( n3058 , n1847 );
nor ( n3059 , n3058 , n2674 );
xnor ( n3060 , n1836 , n3059 );
or ( n3061 , n2166 , n3060 );
not ( n3062 , n2000 );
not ( n3063 , n1626 );
not ( n3064 , n1633 );
not ( n3065 , n3064 );
and ( n3066 , n3063 , n3065 );
and ( n3067 , n1626 , n3064 );
nor ( n3068 , n3066 , n3067 );
not ( n3069 , n3068 );
and ( n3070 , n3062 , n3069 );
not ( n3071 , n1850 );
and ( n3072 , n1490 , n3071 );
not ( n3073 , n1490 );
and ( n3074 , n3073 , n1850 );
nor ( n3075 , n3072 , n3074 );
or ( n3076 , n1523 , n3075 );
not ( n3077 , n3071 );
or ( n3078 , n1994 , n3077 );
nand ( n3079 , n3076 , n3078 );
nor ( n3080 , n3070 , n3079 );
nand ( n3081 , n3061 , n3080 );
nor ( n3082 , n3057 , n3081 );
or ( n3083 , n3082 , n1887 );
not ( n3084 , n152 );
or ( n3085 , n3084 , n2016 );
nand ( n3086 , n3083 , n3085 );
not ( n3087 , n48 );
not ( n3088 , n3087 );
not ( n3089 , n2730 );
and ( n3090 , n3088 , n3089 );
and ( n3091 , n2601 , n2956 );
nor ( n3092 , n3090 , n3091 );
or ( n3093 , n39 , n47 );
nand ( n3094 , n3093 , n2314 );
not ( n3095 , n3094 );
nand ( n3096 , n3095 , n2617 );
not ( n3097 , n2959 );
nand ( n3098 , n3097 , n2595 );
nand ( n3099 , n3092 , n3096 , n3098 );
not ( n3100 , n3099 );
and ( n3101 , n2968 , n2591 );
and ( n3102 , n2950 , n2584 );
nor ( n3103 , n3101 , n3102 );
nand ( n3104 , n2947 , n2580 );
nand ( n3105 , n3100 , n3103 , n3104 );
not ( n3106 , n2580 );
not ( n3107 , n2670 );
or ( n3108 , n3106 , n3107 );
nand ( n3109 , n1484 , n2595 );
nand ( n3110 , n155 , n2606 );
nand ( n3111 , n2697 , n2601 );
nand ( n3112 , n3109 , n3110 , n3111 );
not ( n3113 , n2591 );
not ( n3114 , n2682 );
or ( n3115 , n3113 , n3114 );
and ( n3116 , n2584 , n2692 );
and ( n3117 , n154 , n2617 );
nor ( n3118 , n3116 , n3117 );
nand ( n3119 , n3115 , n3118 );
nor ( n3120 , n3112 , n3119 );
nand ( n3121 , n3108 , n3120 );
or ( n3122 , n3082 , n744 );
not ( n3123 , n151 );
or ( n3124 , n3123 , n745 );
nand ( n3125 , n3122 , n3124 );
or ( n3126 , n2465 , n2579 );
not ( n3127 , n2454 );
or ( n3128 , n2585 , n3127 );
and ( n3129 , n2591 , n2446 );
or ( n3130 , n2433 , n2600 );
or ( n3131 , n2116 , n2594 );
and ( n3132 , n65 , n2606 );
nor ( n3133 , n3030 , n2296 );
nor ( n3134 , n3132 , n3133 );
nand ( n3135 , n3130 , n3131 , n3134 );
nor ( n3136 , n3129 , n3135 );
nand ( n3137 , n3126 , n3128 , n3136 );
or ( n3138 , n2579 , n2856 );
and ( n3139 , n2888 , n2584 );
not ( n3140 , n2876 );
nor ( n3141 , n3140 , n2590 );
nor ( n3142 , n3139 , n3141 );
not ( n3143 , n33 );
not ( n3144 , n2606 );
or ( n3145 , n3143 , n3144 );
or ( n3146 , n2989 , n2296 );
nand ( n3147 , n3145 , n3146 );
not ( n3148 , n2864 );
not ( n3149 , n2595 );
or ( n3150 , n3148 , n3149 );
nand ( n3151 , n2601 , n2862 );
nand ( n3152 , n3150 , n3151 );
nor ( n3153 , n3147 , n3152 );
nand ( n3154 , n3138 , n3142 , n3153 );
or ( n3155 , n3094 , n2334 );
not ( n3156 , n2950 );
not ( n3157 , n2340 );
or ( n3158 , n3156 , n3157 );
nand ( n3159 , n3155 , n3158 );
nand ( n3160 , n2968 , n2288 );
and ( n3161 , n3097 , n2562 );
not ( n3162 , n47 );
not ( n3163 , n2301 );
or ( n3164 , n3162 , n3163 );
nand ( n3165 , n2307 , n2956 );
nand ( n3166 , n3164 , n3165 );
nor ( n3167 , n3161 , n3166 );
nand ( n3168 , n3160 , n3167 );
nor ( n3169 , n3159 , n3168 );
nand ( n3170 , n2947 , n2817 );
nand ( n3171 , n3169 , n3170 );
not ( n3172 , n149 );
not ( n3173 , n744 );
or ( n3174 , n3172 , n3173 );
not ( n3175 , n2741 );
nor ( n3176 , n2371 , n3175 );
not ( n3177 , n3176 );
nand ( n3178 , n3177 , n2063 , n2373 );
not ( n3179 , n3178 );
and ( n3180 , n1378 , n3179 );
and ( n3181 , n1233 , n1490 );
not ( n3182 , n1233 );
and ( n3183 , n3182 , n1489 );
nor ( n3184 , n3181 , n3183 );
or ( n3185 , n2166 , n3184 );
or ( n3186 , n2000 , n3184 );
nor ( n3187 , n1526 , n1522 );
or ( n3188 , n1490 , n3187 );
nand ( n3189 , n3185 , n3186 , n3188 );
nor ( n3190 , n3180 , n3189 );
or ( n3191 , n3190 , n744 );
nand ( n3192 , n3174 , n3191 );
not ( n3193 , n148 );
not ( n3194 , n1887 );
or ( n3195 , n3193 , n3194 );
or ( n3196 , n3190 , n1887 );
nand ( n3197 , n3195 , n3196 );
nand ( n3198 , n3056 , n2580 );
not ( n3199 , n3075 );
not ( n3200 , n3199 );
not ( n3201 , n2601 );
or ( n3202 , n3200 , n3201 );
nand ( n3203 , n153 , n2606 );
nand ( n3204 , n3202 , n3203 );
not ( n3205 , n3071 );
nor ( n3206 , n3205 , n2594 );
nor ( n3207 , n3204 , n3206 );
or ( n3208 , n2583 , n3068 );
not ( n3209 , n150 );
or ( n3210 , n3209 , n2296 );
nand ( n3211 , n3208 , n3210 );
nor ( n3212 , n3060 , n2590 );
nor ( n3213 , n3211 , n3212 );
nand ( n3214 , n3198 , n3207 , n3213 );
or ( n3215 , n3209 , n3017 );
nand ( n3216 , n3056 , n2280 );
or ( n3217 , n3205 , n2298 );
or ( n3218 , n2339 , n3068 );
nand ( n3219 , n3217 , n3218 );
not ( n3220 , n3199 );
not ( n3221 , n2307 );
or ( n3222 , n3220 , n3221 );
or ( n3223 , n3060 , n2287 );
nand ( n3224 , n3222 , n3223 );
nor ( n3225 , n3219 , n3224 );
nand ( n3226 , n3215 , n3216 , n3225 );
not ( n3227 , n146 );
or ( n3228 , n3227 , n3017 );
not ( n3229 , n2279 );
and ( n3230 , n3229 , n3179 );
or ( n3231 , n1490 , n2333 );
not ( n3232 , n3184 );
nand ( n3233 , n2330 , n3232 );
nand ( n3234 , n3231 , n3233 );
nor ( n3235 , n3230 , n3234 );
nand ( n3236 , n3228 , n3235 );
nand ( n3237 , n2580 , n3179 );
nand ( n3238 , n146 , n2617 );
and ( n3239 , n2583 , n2590 );
nor ( n3240 , n3239 , n3184 );
and ( n3241 , n2594 , n2600 );
nor ( n3242 , n3241 , n1490 );
not ( n3243 , n147 );
nor ( n3244 , n3243 , n2730 );
nor ( n3245 , n3240 , n3242 , n3244 );
nand ( n3246 , n3237 , n3238 , n3245 );
and ( n3247 , n158 , n699 , n2275 );
not ( n3248 , n1225 );
and ( n3249 , n3247 , n3248 );
not ( n3250 , n3247 );
not ( n3251 , n178 );
and ( n3252 , n3250 , n3251 );
nor ( n3253 , n3249 , n3252 );
not ( n3254 , n1128 );
not ( n3255 , n1156 );
and ( n3256 , n1185 , n3255 );
not ( n3257 , n1105 );
and ( n3258 , n1192 , n1213 );
and ( n3259 , n3254 , n3256 , n3257 , n3258 );
and ( n3260 , n1199 , n1173 );
nand ( n3261 , n3259 , n3260 , n1134 , n1073 );
nor ( n3262 , n1178 , n3261 );
not ( n3263 , n1178 );
not ( n3264 , n3261 );
or ( n3265 , n3263 , n3264 );
nand ( n3266 , n3265 , n3247 );
or ( n3267 , n3262 , n3266 );
not ( n3268 , n179 );
or ( n3269 , n3268 , n3247 );
nand ( n3270 , n3267 , n3269 );
not ( n3271 , n161 );
not ( n3272 , n705 );
not ( n3273 , n3272 );
or ( n3274 , n3271 , n3273 );
nand ( n3275 , n3274 , n2574 );
endmodule
