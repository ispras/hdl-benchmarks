// IWLS benchmark module "clmB" printed on Wed May 29 22:05:54 2002
module clmB(\IN-i91 , \IN-i191 , \IN-i291 , \IN-i391 , \IN-i90 , \IN-i190 , \IN-i290 , \IN-i390 , \IN-i89 , \IN-i189 , \IN-i289 , \IN-i389 , \IN-i88 , \IN-i188 , \IN-i288 , \IN-i388 , \IN-i87 , \IN-i187 , \IN-i287 , \IN-i387 , \IN-i86 , \IN-i186 , \IN-i286 , \IN-i386 , \IN-i85 , \IN-i185 , \IN-i285 , \IN-i385 , \IN-i84 , \IN-i184 , \IN-i284 , \IN-i384 , \IN-i83 , \IN-i183 , \IN-i283 , \IN-i383 , \IN-i82 , \IN-i182 , \IN-i282 , \IN-i382 , \IN-i81 , \IN-i181 , \IN-i281 , \IN-i381 , \IN-i80 , \IN-i180 , \IN-i280 , \IN-i380 , \IN-i79 , \IN-i179 , \IN-i279 , \IN-i379 , \IN-i78 , \IN-i178 , \IN-i278 , \IN-i378 , \IN-i77 , \IN-i177 , \IN-i277 , \IN-i377 , \IN-i76 , \IN-i176 , \IN-i276 , \IN-i376 , \IN-i75 , \IN-i175 , \IN-i275 , \IN-i375 , \IN-i74 , \IN-i174 , \IN-i274 , \IN-i374 , \IN-i73 , \IN-i173 , \IN-i273 , \IN-i373 , \IN-i72 , \IN-i172 , \IN-i272 , \IN-i372 , \IN-i71 , \IN-i171 , \IN-i271 , \IN-i371 , \IN-i70 , \IN-i170 , \IN-i270 , \IN-i370 , \IN-i69 , \IN-i169 , \IN-i269 , \IN-i369 , \IN-i68 , \IN-i168 , \IN-i268 , \IN-i368 , \IN-i67 , \IN-i167 , \IN-i267 , \IN-i367 , \IN-i66 , \IN-i166 , \IN-i266 , \IN-i366 , \IN-i65 , \IN-i165 , \IN-i265 , \IN-i365 , \IN-i64 , \IN-i164 , \IN-i264 , \IN-i364 , \IN-i63 , \IN-i163 , \IN-i263 , \IN-i363 , \IN-i62 , \IN-i162 , \IN-i262 , \IN-i362 , \IN-i61 , \IN-i161 , \IN-i261 , \IN-i361 , \IN-i60 , \IN-i160 , \IN-i260 , \IN-i360 , \IN-i59 , \IN-i159 , \IN-i259 , \IN-i359 , \IN-i58 , \IN-i158 , \IN-i258 , \IN-i358 , \IN-i57 , \IN-i157 , \IN-i257 , \IN-i357 , \IN-i56 , \IN-i156 , \IN-i256 , \IN-i356 , \IN-i55 , \IN-i155 , \IN-i255 , \IN-i355 , \IN-i54 , \IN-i154 , \IN-i254 , \IN-i354 , \IN-i53 , \IN-i153 , \IN-i253 , \IN-i353 , \IN-i52 , \IN-i152 , \IN-i252 , \IN-i352 , \IN-i51 , \IN-i151 , \IN-i251 , \IN-i351 , \IN-i50 , \IN-i150 , \IN-i250 , \IN-i350 , \IN-i49 , \IN-i149 , \IN-i249 , \IN-i349 , \IN-i148 , \IN-i248 , \IN-i348 , \IN-i147 , \IN-i247 , \IN-i347 , \IN-i146 , \IN-i246 , \IN-i346 , \IN-i145 , \IN-i245 , \IN-i345 , \IN-i144 , \IN-i244 , \IN-i344 , \IN-i143 , \IN-i243 , \IN-i343 , \IN-i142 , \IN-i242 , \IN-i342 , \IN-i141 , \IN-i241 , \IN-i341 , \IN-i140 , \IN-i240 , \IN-i340 , \IN-i139 , \IN-i239 , \IN-i339 , \IN-i138 , \IN-i238 , \IN-i338 , \IN-i137 , \IN-i237 , \IN-i337 , \IN-i136 , \IN-i236 , \IN-i336 , \IN-i135 , \IN-i235 , \IN-i335 , \IN-i134 , \IN-i234 , \IN-i334 , \IN-i133 , \IN-i233 , \IN-i333 , \IN-i132 , \IN-i232 , \IN-i332 , \IN-i131 , \IN-i231 , \IN-i331 , \IN-i130 , \IN-i230 , \IN-i330 , \IN-i129 , \IN-i229 , \IN-i329 , \IN-i28 , \IN-i128 , \IN-i228 , \IN-i328 , i27, \IN-i127 , \IN-i227 , \IN-i327 , i26, \IN-i126 , \IN-i226 , \IN-i326 , i25, \IN-i125 , \IN-i225 , \IN-i325 , i24, \IN-i124 , \IN-i224 , \IN-i324 , i23, \IN-i123 , \IN-i223 , \IN-i323 , i22, \IN-i122 , \IN-i222 , \IN-i322 , i21, \IN-i121 , \IN-i221 , \IN-i321 , i20, \IN-i120 , \IN-i220 , \IN-i320 , i19, \IN-i119 , \IN-i219 , \IN-i319 , i18, \IN-i118 , \IN-i218 , \IN-i318 , i17, \IN-i117 , \IN-i217 , \IN-i317 , i16, \IN-i116 , \IN-i216 , \IN-i316 , \IN-i416 , i15, \IN-i115 , \IN-i215 , \IN-i315 , \IN-i415 , \IN-i114 , \IN-i214 , \IN-i314 , \IN-i414 , \IN-i113 , \IN-i213 , \IN-i313 , \IN-i413 , \IN-i112 , \IN-i212 , \IN-i312 , \IN-i412 , \IN-i111 , \IN-i211 , \IN-i311 , \IN-i411 , \IN-i110 , \IN-i210 , \IN-i310 , \IN-i410 , \IN-i109 , \IN-i209 , \IN-i309 , \IN-i409 , \IN-i108 , \IN-i208 , \IN-i308 , \IN-i408 , \IN-i107 , \IN-i207 , \IN-i307 , \IN-i407 , \IN-i106 , \IN-i206 , \IN-i306 , \IN-i406 , \IN-i105 , \IN-i205 , \IN-i305 , \IN-i405 , \IN-i104 , \IN-i204 , \IN-i304 , \IN-i404 , \IN-i103 , \IN-i203 , \IN-i303 , \IN-i403 , \IN-i102 , \IN-i202 , \IN-i302 , \IN-i402 , \IN-i101 , \IN-i201 , \IN-i301 , \IN-i401 , \IN-i100 , \IN-i200 , \IN-i300 , \IN-i400 , \IN-i99 , \IN-i199 , \IN-i299 , \IN-i399 , \IN-i98 , \IN-i198 , \IN-i298 , \IN-i398 , \IN-i97 , \IN-i197 , \IN-i297 , \IN-i397 , \IN-i96 , \IN-i196 , \IN-i296 , \IN-i396 , \IN-i95 , \IN-i195 , \IN-i295 , \IN-i395 , \IN-i94 , \IN-i194 , \IN-i294 , \IN-i394 , \IN-i93 , \IN-i193 , \IN-i293 , \IN-i393 , \IN-i92 , \IN-i192 , \IN-i292 , \IN-i392 , i91, i191, i291, i391, i90, i190, i290, i390, i89, i189, i289, i389, i88, i188, i288, i388, i87, i187, i287, i387, i86, i186, i286, i386, i85, i185, i285, i385, i84, i184, i284, i384, i83, i183, i283, i383, i82, i182, i282, i382, i81, i181, i281, i381, i80, i180, i280, i380, i79, i179, i279, i379, i78, i178, i278, i378, i77, i177, i277, i377, i76, i176, i276, i376, i75, i175, i275, i375, i74, i174, i274, i374, i73, i173, i273, i373, i72, i172, i272, i372, i71, i171, i271, i371, i70, i170, i270, i370, i69, i169, i269, i369, i68, i168, i268, i368, i67, i167, i267, i367, i66, i166, i266, i366, i65, i165, i265, i365, i64, i164, i264, i364, i63, i163, i263, i363, i62, i162, i262, i362, i61, i161, i261, i361, i60, i160, i260, i360, i59, i159, i259, i359, i58, i158, i258, i358, i57, i157, i257, i357, i56, i156, i256, i356, i55, i155, i255, i355, i54, i154, i254, i354, i53, i153, i253, i353, i52, i152, i252, i352, i51, i151, i251, i351, i50, i150, i250, i350, i49, i149, i249, i349, i148, i248, i348, i147, i247, i347, i146, i246, i346, i145, i245, i345, i144, i244, i344, i143, i243, i343, i142, i242, i342, i141, i241, i341, i140, i240, i340, i139, i239, i339, i138, i238, i338, i137, i237, i337, i136, i236, i336, i135, i235, i335, i134, i234, i334, i133, i233, i333, i132, i232, i332, i131, i231, i331, i130, i230, i330, i129, i229, i329, i28, i128, i228, i328, i127, i227, i327, i126, i226, i326, i125, i225, i325, i124, i224, i324, i123, i223, i323, i122, i222, i322, i121, i221, i321, i120, i220, i320, i119, i219, i319, i118, i218, i318, i117, i217, i317, i116, i216, i316, i416, i115, i215, i315, i415, i114, i214, i314, i414, i113, i213, i313, i413, i112, i212, i312, i412, i111, i211, i311, i411, i110, i210, i310, i410, i109, i209, i309, i409, i108, i208, i308, i408, i107, i207, i307, i407, i106, i206, i306, i406, i105, i205, i305, i405, i104, i204, i304, i404, i103, i203, i303, i403, i102, i202, i302, i402, i101, i201, i301, i401, i100, i200, i300, i400, i99, i199, i299, i399, i98, i198, i298, i398, i97, i197, i297, i397, i96, i196, i296, i396, i95, i195, i295, i395, i94, i194, i294, i394, i93, i193, i293, i393, i92, i192, i292, i392);
input
  i15,
  i16,
  i17,
  i18,
  i19,
  i20,
  i21,
  i22,
  i23,
  i24,
  i25,
  i26,
  i27,
  \IN-i28 ,
  \IN-i49 ,
  \IN-i50 ,
  \IN-i51 ,
  \IN-i52 ,
  \IN-i53 ,
  \IN-i54 ,
  \IN-i55 ,
  \IN-i56 ,
  \IN-i57 ,
  \IN-i58 ,
  \IN-i59 ,
  \IN-i60 ,
  \IN-i61 ,
  \IN-i62 ,
  \IN-i63 ,
  \IN-i64 ,
  \IN-i65 ,
  \IN-i66 ,
  \IN-i67 ,
  \IN-i68 ,
  \IN-i69 ,
  \IN-i70 ,
  \IN-i71 ,
  \IN-i72 ,
  \IN-i73 ,
  \IN-i74 ,
  \IN-i75 ,
  \IN-i76 ,
  \IN-i77 ,
  \IN-i78 ,
  \IN-i79 ,
  \IN-i80 ,
  \IN-i81 ,
  \IN-i82 ,
  \IN-i83 ,
  \IN-i84 ,
  \IN-i85 ,
  \IN-i86 ,
  \IN-i87 ,
  \IN-i88 ,
  \IN-i89 ,
  \IN-i90 ,
  \IN-i91 ,
  \IN-i92 ,
  \IN-i93 ,
  \IN-i94 ,
  \IN-i95 ,
  \IN-i96 ,
  \IN-i97 ,
  \IN-i98 ,
  \IN-i99 ,
  \IN-i110 ,
  \IN-i111 ,
  \IN-i112 ,
  \IN-i113 ,
  \IN-i114 ,
  \IN-i115 ,
  \IN-i116 ,
  \IN-i117 ,
  \IN-i118 ,
  \IN-i119 ,
  \IN-i120 ,
  \IN-i121 ,
  \IN-i122 ,
  \IN-i123 ,
  \IN-i124 ,
  \IN-i125 ,
  \IN-i126 ,
  \IN-i127 ,
  \IN-i128 ,
  \IN-i129 ,
  \IN-i130 ,
  \IN-i131 ,
  \IN-i132 ,
  \IN-i133 ,
  \IN-i134 ,
  \IN-i135 ,
  \IN-i136 ,
  \IN-i137 ,
  \IN-i138 ,
  \IN-i139 ,
  \IN-i140 ,
  \IN-i141 ,
  \IN-i142 ,
  \IN-i143 ,
  \IN-i144 ,
  \IN-i145 ,
  \IN-i146 ,
  \IN-i147 ,
  \IN-i148 ,
  \IN-i149 ,
  \IN-i100 ,
  \IN-i101 ,
  \IN-i102 ,
  \IN-i103 ,
  \IN-i104 ,
  \IN-i105 ,
  \IN-i106 ,
  \IN-i107 ,
  \IN-i108 ,
  \IN-i109 ,
  \IN-i190 ,
  \IN-i191 ,
  \IN-i192 ,
  \IN-i193 ,
  \IN-i194 ,
  \IN-i195 ,
  \IN-i196 ,
  \IN-i197 ,
  \IN-i198 ,
  \IN-i199 ,
  \IN-i150 ,
  \IN-i151 ,
  \IN-i152 ,
  \IN-i153 ,
  \IN-i154 ,
  \IN-i155 ,
  \IN-i156 ,
  \IN-i157 ,
  \IN-i158 ,
  \IN-i159 ,
  \IN-i160 ,
  \IN-i161 ,
  \IN-i162 ,
  \IN-i163 ,
  \IN-i164 ,
  \IN-i165 ,
  \IN-i166 ,
  \IN-i167 ,
  \IN-i168 ,
  \IN-i169 ,
  \IN-i170 ,
  \IN-i171 ,
  \IN-i172 ,
  \IN-i173 ,
  \IN-i174 ,
  \IN-i175 ,
  \IN-i176 ,
  \IN-i177 ,
  \IN-i178 ,
  \IN-i179 ,
  \IN-i180 ,
  \IN-i181 ,
  \IN-i182 ,
  \IN-i183 ,
  \IN-i184 ,
  \IN-i185 ,
  \IN-i186 ,
  \IN-i187 ,
  \IN-i188 ,
  \IN-i189 ,
  \IN-i210 ,
  \IN-i211 ,
  \IN-i212 ,
  \IN-i213 ,
  \IN-i214 ,
  \IN-i215 ,
  \IN-i216 ,
  \IN-i217 ,
  \IN-i218 ,
  \IN-i219 ,
  \IN-i220 ,
  \IN-i221 ,
  \IN-i222 ,
  \IN-i223 ,
  \IN-i224 ,
  \IN-i225 ,
  \IN-i226 ,
  \IN-i227 ,
  \IN-i228 ,
  \IN-i229 ,
  \IN-i230 ,
  \IN-i231 ,
  \IN-i232 ,
  \IN-i233 ,
  \IN-i234 ,
  \IN-i235 ,
  \IN-i236 ,
  \IN-i237 ,
  \IN-i238 ,
  \IN-i239 ,
  \IN-i240 ,
  \IN-i241 ,
  \IN-i242 ,
  \IN-i243 ,
  \IN-i244 ,
  \IN-i245 ,
  \IN-i246 ,
  \IN-i247 ,
  \IN-i248 ,
  \IN-i249 ,
  \IN-i200 ,
  \IN-i201 ,
  \IN-i202 ,
  \IN-i203 ,
  \IN-i204 ,
  \IN-i205 ,
  \IN-i206 ,
  \IN-i207 ,
  \IN-i208 ,
  \IN-i209 ,
  \IN-i290 ,
  \IN-i291 ,
  \IN-i292 ,
  \IN-i293 ,
  \IN-i294 ,
  \IN-i295 ,
  \IN-i296 ,
  \IN-i297 ,
  \IN-i298 ,
  \IN-i299 ,
  \IN-i250 ,
  \IN-i251 ,
  \IN-i252 ,
  \IN-i253 ,
  \IN-i254 ,
  \IN-i255 ,
  \IN-i256 ,
  \IN-i257 ,
  \IN-i258 ,
  \IN-i259 ,
  \IN-i260 ,
  \IN-i261 ,
  \IN-i262 ,
  \IN-i263 ,
  \IN-i264 ,
  \IN-i265 ,
  \IN-i266 ,
  \IN-i267 ,
  \IN-i268 ,
  \IN-i269 ,
  \IN-i270 ,
  \IN-i271 ,
  \IN-i272 ,
  \IN-i273 ,
  \IN-i274 ,
  \IN-i275 ,
  \IN-i276 ,
  \IN-i277 ,
  \IN-i278 ,
  \IN-i279 ,
  \IN-i280 ,
  \IN-i281 ,
  \IN-i282 ,
  \IN-i283 ,
  \IN-i284 ,
  \IN-i285 ,
  \IN-i286 ,
  \IN-i287 ,
  \IN-i288 ,
  \IN-i289 ,
  \IN-i310 ,
  \IN-i311 ,
  \IN-i312 ,
  \IN-i313 ,
  \IN-i314 ,
  \IN-i315 ,
  \IN-i316 ,
  \IN-i317 ,
  \IN-i318 ,
  \IN-i319 ,
  \IN-i320 ,
  \IN-i321 ,
  \IN-i322 ,
  \IN-i323 ,
  \IN-i324 ,
  \IN-i325 ,
  \IN-i326 ,
  \IN-i327 ,
  \IN-i328 ,
  \IN-i329 ,
  \IN-i330 ,
  \IN-i331 ,
  \IN-i332 ,
  \IN-i333 ,
  \IN-i334 ,
  \IN-i335 ,
  \IN-i336 ,
  \IN-i337 ,
  \IN-i338 ,
  \IN-i339 ,
  \IN-i340 ,
  \IN-i341 ,
  \IN-i342 ,
  \IN-i343 ,
  \IN-i344 ,
  \IN-i345 ,
  \IN-i346 ,
  \IN-i347 ,
  \IN-i348 ,
  \IN-i349 ,
  \IN-i300 ,
  \IN-i301 ,
  \IN-i302 ,
  \IN-i303 ,
  \IN-i304 ,
  \IN-i305 ,
  \IN-i306 ,
  \IN-i307 ,
  \IN-i308 ,
  \IN-i309 ,
  \IN-i390 ,
  \IN-i391 ,
  \IN-i392 ,
  \IN-i393 ,
  \IN-i394 ,
  \IN-i395 ,
  \IN-i396 ,
  \IN-i397 ,
  \IN-i398 ,
  \IN-i399 ,
  \IN-i350 ,
  \IN-i351 ,
  \IN-i352 ,
  \IN-i353 ,
  \IN-i354 ,
  \IN-i355 ,
  \IN-i356 ,
  \IN-i357 ,
  \IN-i358 ,
  \IN-i359 ,
  \IN-i360 ,
  \IN-i361 ,
  \IN-i362 ,
  \IN-i363 ,
  \IN-i364 ,
  \IN-i365 ,
  \IN-i366 ,
  \IN-i367 ,
  \IN-i368 ,
  \IN-i369 ,
  \IN-i370 ,
  \IN-i371 ,
  \IN-i372 ,
  \IN-i373 ,
  \IN-i374 ,
  \IN-i375 ,
  \IN-i376 ,
  \IN-i377 ,
  \IN-i378 ,
  \IN-i379 ,
  \IN-i380 ,
  \IN-i381 ,
  \IN-i382 ,
  \IN-i383 ,
  \IN-i384 ,
  \IN-i385 ,
  \IN-i386 ,
  \IN-i387 ,
  \IN-i388 ,
  \IN-i389 ,
  \IN-i410 ,
  \IN-i411 ,
  \IN-i412 ,
  \IN-i413 ,
  \IN-i414 ,
  \IN-i415 ,
  \IN-i416 ,
  \IN-i400 ,
  \IN-i401 ,
  \IN-i402 ,
  \IN-i403 ,
  \IN-i404 ,
  \IN-i405 ,
  \IN-i406 ,
  \IN-i407 ,
  \IN-i408 ,
  \IN-i409 ;
output
  i28,
  i49,
  i50,
  i51,
  i52,
  i53,
  i54,
  i55,
  i56,
  i57,
  i58,
  i59,
  i60,
  i61,
  i62,
  i63,
  i64,
  i65,
  i66,
  i67,
  i68,
  i69,
  i70,
  i71,
  i72,
  i73,
  i74,
  i75,
  i76,
  i77,
  i78,
  i79,
  i80,
  i81,
  i82,
  i83,
  i84,
  i85,
  i86,
  i87,
  i88,
  i89,
  i90,
  i91,
  i92,
  i93,
  i94,
  i95,
  i96,
  i97,
  i98,
  i99,
  i100,
  i101,
  i102,
  i103,
  i104,
  i105,
  i106,
  i107,
  i108,
  i109,
  i110,
  i111,
  i112,
  i113,
  i114,
  i115,
  i116,
  i117,
  i118,
  i119,
  i120,
  i121,
  i122,
  i123,
  i124,
  i125,
  i126,
  i127,
  i128,
  i129,
  i130,
  i131,
  i132,
  i133,
  i134,
  i135,
  i136,
  i137,
  i138,
  i139,
  i140,
  i141,
  i142,
  i143,
  i144,
  i145,
  i146,
  i147,
  i148,
  i149,
  i150,
  i151,
  i152,
  i153,
  i154,
  i155,
  i156,
  i157,
  i158,
  i159,
  i160,
  i161,
  i162,
  i163,
  i164,
  i165,
  i166,
  i167,
  i168,
  i169,
  i170,
  i171,
  i172,
  i173,
  i174,
  i175,
  i176,
  i177,
  i178,
  i179,
  i180,
  i181,
  i182,
  i183,
  i184,
  i185,
  i186,
  i187,
  i188,
  i189,
  i190,
  i191,
  i192,
  i193,
  i194,
  i195,
  i196,
  i197,
  i198,
  i199,
  i200,
  i201,
  i202,
  i203,
  i204,
  i205,
  i206,
  i207,
  i208,
  i209,
  i210,
  i211,
  i212,
  i213,
  i214,
  i215,
  i216,
  i217,
  i218,
  i219,
  i220,
  i221,
  i222,
  i223,
  i224,
  i225,
  i226,
  i227,
  i228,
  i229,
  i230,
  i231,
  i232,
  i233,
  i234,
  i235,
  i236,
  i237,
  i238,
  i239,
  i240,
  i241,
  i242,
  i243,
  i244,
  i245,
  i246,
  i247,
  i248,
  i249,
  i250,
  i251,
  i252,
  i253,
  i254,
  i255,
  i256,
  i257,
  i258,
  i259,
  i260,
  i261,
  i262,
  i263,
  i264,
  i265,
  i266,
  i267,
  i268,
  i269,
  i270,
  i271,
  i272,
  i273,
  i274,
  i275,
  i276,
  i277,
  i278,
  i279,
  i280,
  i281,
  i282,
  i283,
  i284,
  i285,
  i286,
  i287,
  i288,
  i289,
  i290,
  i291,
  i292,
  i293,
  i294,
  i295,
  i296,
  i297,
  i298,
  i299,
  i300,
  i301,
  i302,
  i303,
  i304,
  i305,
  i306,
  i307,
  i308,
  i309,
  i310,
  i311,
  i312,
  i313,
  i314,
  i315,
  i316,
  i317,
  i318,
  i319,
  i320,
  i321,
  i322,
  i323,
  i324,
  i325,
  i326,
  i327,
  i328,
  i329,
  i330,
  i331,
  i332,
  i333,
  i334,
  i335,
  i336,
  i337,
  i338,
  i339,
  i340,
  i341,
  i342,
  i343,
  i344,
  i345,
  i346,
  i347,
  i348,
  i349,
  i350,
  i351,
  i352,
  i353,
  i354,
  i355,
  i356,
  i357,
  i358,
  i359,
  i360,
  i361,
  i362,
  i363,
  i364,
  i365,
  i366,
  i367,
  i368,
  i369,
  i370,
  i371,
  i372,
  i373,
  i374,
  i375,
  i376,
  i377,
  i378,
  i379,
  i380,
  i381,
  i382,
  i383,
  i384,
  i385,
  i386,
  i387,
  i388,
  i389,
  i390,
  i391,
  i392,
  i393,
  i394,
  i395,
  i396,
  i397,
  i398,
  i399,
  i400,
  i401,
  i402,
  i403,
  i404,
  i405,
  i406,
  i407,
  i408,
  i409,
  i410,
  i411,
  i412,
  i413,
  i414,
  i415,
  i416;
assign
  i28 = \IN-i28 ,
  i49 = \IN-i49 ,
  i50 = \IN-i50 ,
  i51 = \IN-i51 ,
  i52 = \IN-i52 ,
  i53 = \IN-i53 ,
  i54 = \IN-i54 ,
  i55 = \IN-i55 ,
  i56 = \IN-i56 ,
  i57 = \IN-i57 ,
  i58 = \IN-i58 ,
  i59 = \IN-i59 ,
  i60 = \IN-i60 ,
  i61 = \IN-i61 ,
  i62 = \IN-i62 ,
  i63 = \IN-i63 ,
  i64 = \IN-i64 ,
  i65 = \IN-i65 ,
  i66 = \IN-i66 ,
  i67 = \IN-i67 ,
  i68 = \IN-i68 ,
  i69 = \IN-i69 ,
  i70 = \IN-i70 ,
  i71 = \IN-i71 ,
  i72 = \IN-i72 ,
  i73 = \IN-i73 ,
  i74 = \IN-i74 ,
  i75 = \IN-i75 ,
  i76 = \IN-i76 ,
  i77 = \IN-i77 ,
  i78 = \IN-i78 ,
  i79 = \IN-i79 ,
  i80 = \IN-i80 ,
  i81 = \IN-i81 ,
  i82 = \IN-i82 ,
  i83 = \IN-i83 ,
  i84 = \IN-i84 ,
  i85 = \IN-i85 ,
  i86 = \IN-i86 ,
  i87 = \IN-i87 ,
  i88 = \IN-i88 ,
  i89 = \IN-i89 ,
  i90 = \IN-i90 ,
  i91 = \IN-i91 ,
  i92 = \IN-i92 ,
  i93 = \IN-i93 ,
  i94 = \IN-i94 ,
  i95 = \IN-i95 ,
  i96 = \IN-i96 ,
  i97 = \IN-i97 ,
  i98 = \IN-i98 ,
  i99 = \IN-i99 ,
  i100 = \IN-i100 ,
  i101 = \IN-i101 ,
  i102 = \IN-i102 ,
  i103 = \IN-i103 ,
  i104 = \IN-i104 ,
  i105 = \IN-i105 ,
  i106 = \IN-i106 ,
  i107 = \IN-i107 ,
  i108 = \IN-i108 ,
  i109 = \IN-i109 ,
  i110 = \IN-i110 ,
  i111 = \IN-i111 ,
  i112 = \IN-i112 ,
  i113 = \IN-i113 ,
  i114 = \IN-i114 ,
  i115 = \IN-i115 ,
  i116 = \IN-i116 ,
  i117 = \IN-i117 ,
  i118 = \IN-i118 ,
  i119 = \IN-i119 ,
  i120 = \IN-i120 ,
  i121 = \IN-i121 ,
  i122 = \IN-i122 ,
  i123 = \IN-i123 ,
  i124 = \IN-i124 ,
  i125 = \IN-i125 ,
  i126 = \IN-i126 ,
  i127 = \IN-i127 ,
  i128 = \IN-i128 ,
  i129 = \IN-i129 ,
  i130 = \IN-i130 ,
  i131 = \IN-i131 ,
  i132 = \IN-i132 ,
  i133 = \IN-i133 ,
  i134 = \IN-i134 ,
  i135 = \IN-i135 ,
  i136 = \IN-i136 ,
  i137 = \IN-i137 ,
  i138 = \IN-i138 ,
  i139 = \IN-i139 ,
  i140 = \IN-i140 ,
  i141 = \IN-i141 ,
  i142 = \IN-i142 ,
  i143 = \IN-i143 ,
  i144 = \IN-i144 ,
  i145 = \IN-i145 ,
  i146 = \IN-i146 ,
  i147 = \IN-i147 ,
  i148 = \IN-i148 ,
  i149 = \IN-i149 ,
  i150 = \IN-i150 ,
  i151 = \IN-i151 ,
  i152 = \IN-i152 ,
  i153 = \IN-i153 ,
  i154 = \IN-i154 ,
  i155 = \IN-i155 ,
  i156 = \IN-i156 ,
  i157 = \IN-i157 ,
  i158 = \IN-i158 ,
  i159 = \IN-i159 ,
  i160 = \IN-i160 ,
  i161 = \IN-i161 ,
  i162 = \IN-i162 ,
  i163 = \IN-i163 ,
  i164 = \IN-i164 ,
  i165 = \IN-i165 ,
  i166 = \IN-i166 ,
  i167 = \IN-i167 ,
  i168 = \IN-i168 ,
  i169 = \IN-i169 ,
  i170 = \IN-i170 ,
  i171 = \IN-i171 ,
  i172 = \IN-i172 ,
  i173 = \IN-i173 ,
  i174 = \IN-i174 ,
  i175 = \IN-i175 ,
  i176 = \IN-i176 ,
  i177 = \IN-i177 ,
  i178 = \IN-i178 ,
  i179 = \IN-i179 ,
  i180 = \IN-i180 ,
  i181 = \IN-i181 ,
  i182 = \IN-i182 ,
  i183 = \IN-i183 ,
  i184 = \IN-i184 ,
  i185 = \IN-i185 ,
  i186 = \IN-i186 ,
  i187 = \IN-i187 ,
  i188 = \IN-i188 ,
  i189 = \IN-i189 ,
  i190 = \IN-i190 ,
  i191 = \IN-i191 ,
  i192 = \IN-i192 ,
  i193 = \IN-i193 ,
  i194 = \IN-i194 ,
  i195 = \IN-i195 ,
  i196 = \IN-i196 ,
  i197 = \IN-i197 ,
  i198 = \IN-i198 ,
  i199 = \IN-i199 ,
  i200 = \IN-i200 ,
  i201 = \IN-i201 ,
  i202 = \IN-i202 ,
  i203 = \IN-i203 ,
  i204 = \IN-i204 ,
  i205 = \IN-i205 ,
  i206 = \IN-i206 ,
  i207 = \IN-i207 ,
  i208 = \IN-i208 ,
  i209 = \IN-i209 ,
  i210 = \IN-i210 ,
  i211 = \IN-i211 ,
  i212 = \IN-i212 ,
  i213 = \IN-i213 ,
  i214 = \IN-i214 ,
  i215 = \IN-i215 ,
  i216 = \IN-i216 ,
  i217 = \IN-i217 ,
  i218 = \IN-i218 ,
  i219 = \IN-i219 ,
  i220 = \IN-i220 ,
  i221 = \IN-i221 ,
  i222 = \IN-i222 ,
  i223 = \IN-i223 ,
  i224 = \IN-i224 ,
  i225 = \IN-i225 ,
  i226 = \IN-i226 ,
  i227 = \IN-i227 ,
  i228 = \IN-i228 ,
  i229 = \IN-i229 ,
  i230 = \IN-i230 ,
  i231 = \IN-i231 ,
  i232 = \IN-i232 ,
  i233 = \IN-i233 ,
  i234 = \IN-i234 ,
  i235 = \IN-i235 ,
  i236 = \IN-i236 ,
  i237 = \IN-i237 ,
  i238 = \IN-i238 ,
  i239 = \IN-i239 ,
  i240 = \IN-i240 ,
  i241 = \IN-i241 ,
  i242 = \IN-i242 ,
  i243 = \IN-i243 ,
  i244 = \IN-i244 ,
  i245 = \IN-i245 ,
  i246 = \IN-i246 ,
  i247 = \IN-i247 ,
  i248 = \IN-i248 ,
  i249 = \IN-i249 ,
  i250 = \IN-i250 ,
  i251 = \IN-i251 ,
  i252 = \IN-i252 ,
  i253 = \IN-i253 ,
  i254 = \IN-i254 ,
  i255 = \IN-i255 ,
  i256 = \IN-i256 ,
  i257 = \IN-i257 ,
  i258 = \IN-i258 ,
  i259 = \IN-i259 ,
  i260 = \IN-i260 ,
  i261 = \IN-i261 ,
  i262 = \IN-i262 ,
  i263 = \IN-i263 ,
  i264 = \IN-i264 ,
  i265 = \IN-i265 ,
  i266 = \IN-i266 ,
  i267 = \IN-i267 ,
  i268 = \IN-i268 ,
  i269 = \IN-i269 ,
  i270 = \IN-i270 ,
  i271 = \IN-i271 ,
  i272 = \IN-i272 ,
  i273 = \IN-i273 ,
  i274 = \IN-i274 ,
  i275 = \IN-i275 ,
  i276 = \IN-i276 ,
  i277 = \IN-i277 ,
  i278 = \IN-i278 ,
  i279 = \IN-i279 ,
  i280 = \IN-i280 ,
  i281 = \IN-i281 ,
  i282 = \IN-i282 ,
  i283 = \IN-i283 ,
  i284 = \IN-i284 ,
  i285 = \IN-i285 ,
  i286 = \IN-i286 ,
  i287 = \IN-i287 ,
  i288 = \IN-i288 ,
  i289 = \IN-i289 ,
  i290 = \IN-i290 ,
  i291 = \IN-i291 ,
  i292 = \IN-i292 ,
  i293 = \IN-i293 ,
  i294 = \IN-i294 ,
  i295 = \IN-i295 ,
  i296 = \IN-i296 ,
  i297 = \IN-i297 ,
  i298 = \IN-i298 ,
  i299 = \IN-i299 ,
  i300 = \IN-i300 ,
  i301 = \IN-i301 ,
  i302 = \IN-i302 ,
  i303 = \IN-i303 ,
  i304 = \IN-i304 ,
  i305 = \IN-i305 ,
  i306 = \IN-i306 ,
  i307 = \IN-i307 ,
  i308 = \IN-i308 ,
  i309 = \IN-i309 ,
  i310 = \IN-i310 ,
  i311 = \IN-i311 ,
  i312 = \IN-i312 ,
  i313 = \IN-i313 ,
  i314 = \IN-i314 ,
  i315 = \IN-i315 ,
  i316 = \IN-i316 ,
  i317 = \IN-i317 ,
  i318 = \IN-i318 ,
  i319 = \IN-i319 ,
  i320 = \IN-i320 ,
  i321 = \IN-i321 ,
  i322 = \IN-i322 ,
  i323 = \IN-i323 ,
  i324 = \IN-i324 ,
  i325 = \IN-i325 ,
  i326 = \IN-i326 ,
  i327 = \IN-i327 ,
  i328 = \IN-i328 ,
  i329 = \IN-i329 ,
  i330 = \IN-i330 ,
  i331 = \IN-i331 ,
  i332 = \IN-i332 ,
  i333 = \IN-i333 ,
  i334 = \IN-i334 ,
  i335 = \IN-i335 ,
  i336 = \IN-i336 ,
  i337 = \IN-i337 ,
  i338 = \IN-i338 ,
  i339 = \IN-i339 ,
  i340 = \IN-i340 ,
  i341 = \IN-i341 ,
  i342 = \IN-i342 ,
  i343 = \IN-i343 ,
  i344 = \IN-i344 ,
  i345 = \IN-i345 ,
  i346 = \IN-i346 ,
  i347 = \IN-i347 ,
  i348 = \IN-i348 ,
  i349 = \IN-i349 ,
  i350 = \IN-i350 ,
  i351 = \IN-i351 ,
  i352 = \IN-i352 ,
  i353 = \IN-i353 ,
  i354 = \IN-i354 ,
  i355 = \IN-i355 ,
  i356 = \IN-i356 ,
  i357 = \IN-i357 ,
  i358 = \IN-i358 ,
  i359 = \IN-i359 ,
  i360 = \IN-i360 ,
  i361 = \IN-i361 ,
  i362 = \IN-i362 ,
  i363 = \IN-i363 ,
  i364 = \IN-i364 ,
  i365 = \IN-i365 ,
  i366 = \IN-i366 ,
  i367 = \IN-i367 ,
  i368 = \IN-i368 ,
  i369 = \IN-i369 ,
  i370 = \IN-i370 ,
  i371 = \IN-i371 ,
  i372 = \IN-i372 ,
  i373 = \IN-i373 ,
  i374 = \IN-i374 ,
  i375 = \IN-i375 ,
  i376 = \IN-i376 ,
  i377 = \IN-i377 ,
  i378 = \IN-i378 ,
  i379 = \IN-i379 ,
  i380 = \IN-i380 ,
  i381 = \IN-i381 ,
  i382 = \IN-i382 ,
  i383 = \IN-i383 ,
  i384 = \IN-i384 ,
  i385 = \IN-i385 ,
  i386 = \IN-i386 ,
  i387 = \IN-i387 ,
  i388 = \IN-i388 ,
  i389 = \IN-i389 ,
  i390 = \IN-i390 ,
  i391 = \IN-i391 ,
  i392 = \IN-i392 ,
  i393 = \IN-i393 ,
  i394 = \IN-i394 ,
  i395 = \IN-i395 ,
  i396 = \IN-i396 ,
  i397 = \IN-i397 ,
  i398 = \IN-i398 ,
  i399 = \IN-i399 ,
  i400 = \IN-i400 ,
  i401 = \IN-i401 ,
  i402 = \IN-i402 ,
  i403 = \IN-i403 ,
  i404 = \IN-i404 ,
  i405 = \IN-i405 ,
  i406 = \IN-i406 ,
  i407 = \IN-i407 ,
  i408 = \IN-i408 ,
  i409 = \IN-i409 ,
  i410 = \IN-i410 ,
  i411 = \IN-i411 ,
  i412 = \IN-i412 ,
  i413 = \IN-i413 ,
  i414 = \IN-i414 ,
  i415 = \IN-i415 ,
  i416 = \IN-i416 ;
endmodule

